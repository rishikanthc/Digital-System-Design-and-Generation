
module controlpath ( clk, reset, start, loadMatrix, loadVector, wr_en_x, 
        clear_acc, wr_en_y, done, addr_x, addr_y, .addr_a({\addr_a[31][5] , 
        \addr_a[31][4] , \addr_a[31][3] , \addr_a[31][2] , \addr_a[31][1] , 
        \addr_a[31][0] , \addr_a[30][5] , \addr_a[30][4] , \addr_a[30][3] , 
        \addr_a[30][2] , \addr_a[30][1] , \addr_a[30][0] , \addr_a[29][5] , 
        \addr_a[29][4] , \addr_a[29][3] , \addr_a[29][2] , \addr_a[29][1] , 
        \addr_a[29][0] , \addr_a[28][5] , \addr_a[28][4] , \addr_a[28][3] , 
        \addr_a[28][2] , \addr_a[28][1] , \addr_a[28][0] , \addr_a[27][5] , 
        \addr_a[27][4] , \addr_a[27][3] , \addr_a[27][2] , \addr_a[27][1] , 
        \addr_a[27][0] , \addr_a[26][5] , \addr_a[26][4] , \addr_a[26][3] , 
        \addr_a[26][2] , \addr_a[26][1] , \addr_a[26][0] , \addr_a[25][5] , 
        \addr_a[25][4] , \addr_a[25][3] , \addr_a[25][2] , \addr_a[25][1] , 
        \addr_a[25][0] , \addr_a[24][5] , \addr_a[24][4] , \addr_a[24][3] , 
        \addr_a[24][2] , \addr_a[24][1] , \addr_a[24][0] , \addr_a[23][5] , 
        \addr_a[23][4] , \addr_a[23][3] , \addr_a[23][2] , \addr_a[23][1] , 
        \addr_a[23][0] , \addr_a[22][5] , \addr_a[22][4] , \addr_a[22][3] , 
        \addr_a[22][2] , \addr_a[22][1] , \addr_a[22][0] , \addr_a[21][5] , 
        \addr_a[21][4] , \addr_a[21][3] , \addr_a[21][2] , \addr_a[21][1] , 
        \addr_a[21][0] , \addr_a[20][5] , \addr_a[20][4] , \addr_a[20][3] , 
        \addr_a[20][2] , \addr_a[20][1] , \addr_a[20][0] , \addr_a[19][5] , 
        \addr_a[19][4] , \addr_a[19][3] , \addr_a[19][2] , \addr_a[19][1] , 
        \addr_a[19][0] , \addr_a[18][5] , \addr_a[18][4] , \addr_a[18][3] , 
        \addr_a[18][2] , \addr_a[18][1] , \addr_a[18][0] , \addr_a[17][5] , 
        \addr_a[17][4] , \addr_a[17][3] , \addr_a[17][2] , \addr_a[17][1] , 
        \addr_a[17][0] , \addr_a[16][5] , \addr_a[16][4] , \addr_a[16][3] , 
        \addr_a[16][2] , \addr_a[16][1] , \addr_a[16][0] , \addr_a[15][5] , 
        \addr_a[15][4] , \addr_a[15][3] , \addr_a[15][2] , \addr_a[15][1] , 
        \addr_a[15][0] , \addr_a[14][5] , \addr_a[14][4] , \addr_a[14][3] , 
        \addr_a[14][2] , \addr_a[14][1] , \addr_a[14][0] , \addr_a[13][5] , 
        \addr_a[13][4] , \addr_a[13][3] , \addr_a[13][2] , \addr_a[13][1] , 
        \addr_a[13][0] , \addr_a[12][5] , \addr_a[12][4] , \addr_a[12][3] , 
        \addr_a[12][2] , \addr_a[12][1] , \addr_a[12][0] , \addr_a[11][5] , 
        \addr_a[11][4] , \addr_a[11][3] , \addr_a[11][2] , \addr_a[11][1] , 
        \addr_a[11][0] , \addr_a[10][5] , \addr_a[10][4] , \addr_a[10][3] , 
        \addr_a[10][2] , \addr_a[10][1] , \addr_a[10][0] , \addr_a[9][5] , 
        \addr_a[9][4] , \addr_a[9][3] , \addr_a[9][2] , \addr_a[9][1] , 
        \addr_a[9][0] , \addr_a[8][5] , \addr_a[8][4] , \addr_a[8][3] , 
        \addr_a[8][2] , \addr_a[8][1] , \addr_a[8][0] , \addr_a[7][5] , 
        \addr_a[7][4] , \addr_a[7][3] , \addr_a[7][2] , \addr_a[7][1] , 
        \addr_a[7][0] , \addr_a[6][5] , \addr_a[6][4] , \addr_a[6][3] , 
        \addr_a[6][2] , \addr_a[6][1] , \addr_a[6][0] , \addr_a[5][5] , 
        \addr_a[5][4] , \addr_a[5][3] , \addr_a[5][2] , \addr_a[5][1] , 
        \addr_a[5][0] , \addr_a[4][5] , \addr_a[4][4] , \addr_a[4][3] , 
        \addr_a[4][2] , \addr_a[4][1] , \addr_a[4][0] , \addr_a[3][5] , 
        \addr_a[3][4] , \addr_a[3][3] , \addr_a[3][2] , \addr_a[3][1] , 
        \addr_a[3][0] , \addr_a[2][5] , \addr_a[2][4] , \addr_a[2][3] , 
        \addr_a[2][2] , \addr_a[2][1] , \addr_a[2][0] , \addr_a[1][5] , 
        \addr_a[1][4] , \addr_a[1][3] , \addr_a[1][2] , \addr_a[1][1] , 
        \addr_a[1][0] , \addr_a[0][5] , \addr_a[0][4] , \addr_a[0][3] , 
        \addr_a[0][2] , \addr_a[0][1] , \addr_a[0][0] }), wr_en_a );
  output [5:0] addr_x;
  output [5:0] addr_y;
  output [31:0] wr_en_a;
  input clk, reset, start, loadMatrix, loadVector;
  output wr_en_x, clear_acc, wr_en_y, done, \addr_a[31][5] , \addr_a[31][4] ,
         \addr_a[31][3] , \addr_a[31][2] , \addr_a[31][1] , \addr_a[31][0] ,
         \addr_a[30][5] , \addr_a[30][4] , \addr_a[30][3] , \addr_a[30][2] ,
         \addr_a[30][1] , \addr_a[30][0] , \addr_a[29][5] , \addr_a[29][4] ,
         \addr_a[29][3] , \addr_a[29][2] , \addr_a[29][1] , \addr_a[29][0] ,
         \addr_a[28][5] , \addr_a[28][4] , \addr_a[28][3] , \addr_a[28][2] ,
         \addr_a[28][1] , \addr_a[28][0] , \addr_a[27][5] , \addr_a[27][4] ,
         \addr_a[27][3] , \addr_a[27][2] , \addr_a[27][1] , \addr_a[27][0] ,
         \addr_a[26][5] , \addr_a[26][4] , \addr_a[26][3] , \addr_a[26][2] ,
         \addr_a[26][1] , \addr_a[26][0] , \addr_a[25][5] , \addr_a[25][4] ,
         \addr_a[25][3] , \addr_a[25][2] , \addr_a[25][1] , \addr_a[25][0] ,
         \addr_a[24][5] , \addr_a[24][4] , \addr_a[24][3] , \addr_a[24][2] ,
         \addr_a[24][1] , \addr_a[24][0] , \addr_a[23][5] , \addr_a[23][4] ,
         \addr_a[23][3] , \addr_a[23][2] , \addr_a[23][1] , \addr_a[23][0] ,
         \addr_a[22][5] , \addr_a[22][4] , \addr_a[22][3] , \addr_a[22][2] ,
         \addr_a[22][1] , \addr_a[22][0] , \addr_a[21][5] , \addr_a[21][4] ,
         \addr_a[21][3] , \addr_a[21][2] , \addr_a[21][1] , \addr_a[21][0] ,
         \addr_a[20][5] , \addr_a[20][4] , \addr_a[20][3] , \addr_a[20][2] ,
         \addr_a[20][1] , \addr_a[20][0] , \addr_a[19][5] , \addr_a[19][4] ,
         \addr_a[19][3] , \addr_a[19][2] , \addr_a[19][1] , \addr_a[19][0] ,
         \addr_a[18][5] , \addr_a[18][4] , \addr_a[18][3] , \addr_a[18][2] ,
         \addr_a[18][1] , \addr_a[18][0] , \addr_a[17][5] , \addr_a[17][4] ,
         \addr_a[17][3] , \addr_a[17][2] , \addr_a[17][1] , \addr_a[17][0] ,
         \addr_a[16][5] , \addr_a[16][4] , \addr_a[16][3] , \addr_a[16][2] ,
         \addr_a[16][1] , \addr_a[16][0] , \addr_a[15][5] , \addr_a[15][4] ,
         \addr_a[15][3] , \addr_a[15][2] , \addr_a[15][1] , \addr_a[15][0] ,
         \addr_a[14][5] , \addr_a[14][4] , \addr_a[14][3] , \addr_a[14][2] ,
         \addr_a[14][1] , \addr_a[14][0] , \addr_a[13][5] , \addr_a[13][4] ,
         \addr_a[13][3] , \addr_a[13][2] , \addr_a[13][1] , \addr_a[13][0] ,
         \addr_a[12][5] , \addr_a[12][4] , \addr_a[12][3] , \addr_a[12][2] ,
         \addr_a[12][1] , \addr_a[12][0] , \addr_a[11][5] , \addr_a[11][4] ,
         \addr_a[11][3] , \addr_a[11][2] , \addr_a[11][1] , \addr_a[11][0] ,
         \addr_a[10][5] , \addr_a[10][4] , \addr_a[10][3] , \addr_a[10][2] ,
         \addr_a[10][1] , \addr_a[10][0] , \addr_a[9][5] , \addr_a[9][4] ,
         \addr_a[9][3] , \addr_a[9][2] , \addr_a[9][1] , \addr_a[9][0] ,
         \addr_a[8][5] , \addr_a[8][4] , \addr_a[8][3] , \addr_a[8][2] ,
         \addr_a[8][1] , \addr_a[8][0] , \addr_a[7][5] , \addr_a[7][4] ,
         \addr_a[7][3] , \addr_a[7][2] , \addr_a[7][1] , \addr_a[7][0] ,
         \addr_a[6][5] , \addr_a[6][4] , \addr_a[6][3] , \addr_a[6][2] ,
         \addr_a[6][1] , \addr_a[6][0] , \addr_a[5][5] , \addr_a[5][4] ,
         \addr_a[5][3] , \addr_a[5][2] , \addr_a[5][1] , \addr_a[5][0] ,
         \addr_a[4][5] , \addr_a[4][4] , \addr_a[4][3] , \addr_a[4][2] ,
         \addr_a[4][1] , \addr_a[4][0] , \addr_a[3][5] , \addr_a[3][4] ,
         \addr_a[3][3] , \addr_a[3][2] , \addr_a[3][1] , \addr_a[3][0] ,
         \addr_a[2][5] , \addr_a[2][4] , \addr_a[2][3] , \addr_a[2][2] ,
         \addr_a[2][1] , \addr_a[2][0] , \addr_a[1][5] , \addr_a[1][4] ,
         \addr_a[1][3] , \addr_a[1][2] , \addr_a[1][1] , \addr_a[1][0] ,
         \addr_a[0][5] , \addr_a[0][4] , \addr_a[0][3] , \addr_a[0][2] ,
         \addr_a[0][1] , \addr_a[0][0] ;
  wire   N173, N175, N176, N177, N178, N179, N180, N182, N183, N184, N185,
         N186, N200, N201, N202, N210, N211, N212, N213, N214, N215, N602,
         N603, N604, N605, N606, N607, N608, N1171, N1172, N1173, N1174, N1175,
         n13, n19, n20, n21, n28, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, \add_83/carry[5] , \add_83/carry[4] , \add_83/carry[3] ,
         \add_83/carry[2] , \add_80/carry[5] , \add_80/carry[4] ,
         \add_80/carry[3] , \add_80/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n14, n15, n16, n17, n18, n22, n23, n24, n25, n26,
         n27, n29, n30, n31, n32, n33, n34, n35, n36, n179, n180, n181, n182,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200;
  wire   [2:0] state;
  wire   [5:0] counter;
  wire   [5:0] counter2;
  assign \addr_a[0][5]  = 1'b0;
  assign \addr_a[1][5]  = 1'b0;
  assign \addr_a[2][5]  = 1'b0;
  assign \addr_a[3][5]  = 1'b0;
  assign \addr_a[4][5]  = 1'b0;
  assign \addr_a[5][5]  = 1'b0;
  assign \addr_a[6][5]  = 1'b0;
  assign \addr_a[7][5]  = 1'b0;
  assign \addr_a[8][5]  = 1'b0;
  assign \addr_a[9][5]  = 1'b0;
  assign \addr_a[10][5]  = 1'b0;
  assign \addr_a[11][5]  = 1'b0;
  assign \addr_a[12][5]  = 1'b0;
  assign \addr_a[13][5]  = 1'b0;
  assign \addr_a[14][5]  = 1'b0;
  assign \addr_a[15][5]  = 1'b0;
  assign \addr_a[16][5]  = 1'b0;
  assign \addr_a[17][5]  = 1'b0;
  assign \addr_a[18][5]  = 1'b0;
  assign \addr_a[19][5]  = 1'b0;
  assign \addr_a[20][5]  = 1'b0;
  assign \addr_a[21][5]  = 1'b0;
  assign \addr_a[22][5]  = 1'b0;
  assign \addr_a[23][5]  = 1'b0;
  assign \addr_a[24][5]  = 1'b0;
  assign \addr_a[25][5]  = 1'b0;
  assign \addr_a[26][5]  = 1'b0;
  assign \addr_a[27][5]  = 1'b0;
  assign \addr_a[28][5]  = 1'b0;
  assign \addr_a[29][5]  = 1'b0;
  assign \addr_a[30][5]  = 1'b0;
  assign \addr_a[31][5]  = 1'b0;
  assign addr_x[5] = 1'b0;

  OAI21_X2 U103 ( .B1(n192), .B2(n141), .A(n11), .ZN(addr_x[3]) );
  OAI21_X2 U108 ( .B1(n43), .B2(n6), .A(n11), .ZN(\addr_a[9][3] ) );
  OAI21_X2 U114 ( .B1(n48), .B2(n5), .A(n11), .ZN(\addr_a[8][3] ) );
  OAI21_X2 U120 ( .B1(n51), .B2(n150), .A(n11), .ZN(\addr_a[7][3] ) );
  OAI21_X2 U126 ( .B1(n55), .B2(n150), .A(n11), .ZN(\addr_a[6][3] ) );
  OAI21_X2 U132 ( .B1(n58), .B2(n150), .A(n11), .ZN(\addr_a[5][3] ) );
  OAI21_X2 U138 ( .B1(n61), .B2(n150), .A(n11), .ZN(\addr_a[4][3] ) );
  OAI21_X2 U144 ( .B1(n64), .B2(n150), .A(n11), .ZN(\addr_a[3][3] ) );
  OAI21_X2 U150 ( .B1(n67), .B2(n150), .A(n11), .ZN(\addr_a[31][3] ) );
  OAI21_X2 U156 ( .B1(n72), .B2(n6), .A(n10), .ZN(\addr_a[30][3] ) );
  OAI21_X2 U162 ( .B1(n74), .B2(n6), .A(n10), .ZN(\addr_a[2][3] ) );
  OAI21_X2 U167 ( .B1(n77), .B2(n6), .A(n10), .ZN(\addr_a[29][3] ) );
  OAI21_X2 U173 ( .B1(n79), .B2(n6), .A(n10), .ZN(\addr_a[28][3] ) );
  OAI21_X2 U179 ( .B1(n81), .B2(n6), .A(n10), .ZN(\addr_a[27][3] ) );
  OAI21_X2 U185 ( .B1(n83), .B2(n6), .A(n10), .ZN(\addr_a[26][3] ) );
  OAI21_X2 U191 ( .B1(n85), .B2(n6), .A(n10), .ZN(\addr_a[25][3] ) );
  OAI21_X2 U197 ( .B1(n87), .B2(n6), .A(n10), .ZN(\addr_a[24][3] ) );
  NOR3_X2 U202 ( .A1(n28), .A2(counter[5]), .A3(n25), .ZN(n163) );
  OAI21_X2 U204 ( .B1(n90), .B2(n6), .A(n10), .ZN(\addr_a[23][3] ) );
  OAI21_X2 U210 ( .B1(n93), .B2(n6), .A(n10), .ZN(\addr_a[22][3] ) );
  OAI21_X2 U216 ( .B1(n95), .B2(n6), .A(n10), .ZN(\addr_a[21][3] ) );
  OAI21_X2 U222 ( .B1(n97), .B2(n6), .A(n10), .ZN(\addr_a[20][3] ) );
  OAI21_X2 U228 ( .B1(n38), .B2(n5), .A(n142), .ZN(\addr_a[1][3] ) );
  OAI21_X2 U234 ( .B1(n100), .B2(n5), .A(n142), .ZN(\addr_a[19][3] ) );
  OAI21_X2 U240 ( .B1(n102), .B2(n5), .A(n142), .ZN(\addr_a[18][3] ) );
  OAI21_X2 U246 ( .B1(n104), .B2(n5), .A(n11), .ZN(\addr_a[17][3] ) );
  OAI21_X2 U253 ( .B1(n106), .B2(n5), .A(n142), .ZN(\addr_a[16][3] ) );
  NOR3_X2 U258 ( .A1(counter[3]), .A2(counter[5]), .A3(n25), .ZN(n165) );
  OAI21_X2 U260 ( .B1(n108), .B2(n5), .A(n142), .ZN(\addr_a[15][3] ) );
  OAI21_X2 U267 ( .B1(n110), .B2(n5), .A(n142), .ZN(\addr_a[14][3] ) );
  OAI21_X2 U274 ( .B1(n112), .B2(n5), .A(n142), .ZN(\addr_a[13][3] ) );
  OAI21_X2 U281 ( .B1(n114), .B2(n5), .A(n11), .ZN(\addr_a[12][3] ) );
  OAI21_X2 U288 ( .B1(n116), .B2(n5), .A(n142), .ZN(\addr_a[11][3] ) );
  OAI21_X2 U295 ( .B1(n118), .B2(n5), .A(n11), .ZN(\addr_a[10][3] ) );
  NOR3_X2 U300 ( .A1(counter[4]), .A2(counter[5]), .A3(n28), .ZN(n154) );
  OAI21_X2 U305 ( .B1(n40), .B2(n5), .A(n142), .ZN(\addr_a[0][3] ) );
  NOR3_X2 U342 ( .A1(counter[4]), .A2(counter[5]), .A3(counter[3]), .ZN(n158)
         );
  NAND3_X1 U367 ( .A1(N605), .A2(n88), .A3(N606), .ZN(n70) );
  NAND3_X1 U368 ( .A1(n194), .A2(n195), .A3(N602), .ZN(n45) );
  NAND3_X1 U369 ( .A1(n88), .A2(n18), .A3(N606), .ZN(n91) );
  NAND3_X1 U370 ( .A1(N603), .A2(N602), .A3(N604), .ZN(n53) );
  NAND3_X1 U371 ( .A1(N603), .A2(counter[0]), .A3(N604), .ZN(n56) );
  NAND3_X1 U372 ( .A1(N602), .A2(n194), .A3(N604), .ZN(n59) );
  NAND3_X1 U373 ( .A1(counter[0]), .A2(n194), .A3(N604), .ZN(n62) );
  NAND3_X1 U374 ( .A1(N602), .A2(n195), .A3(N603), .ZN(n65) );
  NAND3_X1 U375 ( .A1(counter[0]), .A2(n195), .A3(N603), .ZN(n75) );
  NAND3_X1 U376 ( .A1(n88), .A2(n196), .A3(N605), .ZN(n44) );
  NAND3_X1 U377 ( .A1(n18), .A2(n196), .A3(n88), .ZN(n52) );
  NAND3_X1 U378 ( .A1(n194), .A2(n195), .A3(counter[0]), .ZN(n49) );
  NAND3_X1 U379 ( .A1(n129), .A2(n130), .A3(N173), .ZN(n121) );
  NAND3_X1 U380 ( .A1(state[1]), .A2(n19), .A3(state[0]), .ZN(n131) );
  NAND3_X1 U382 ( .A1(n129), .A2(state[0]), .A3(n171), .ZN(n170) );
  NAND3_X1 U383 ( .A1(n20), .A2(n19), .A3(state[0]), .ZN(n120) );
  HA_X1 \add_83/U1_1_1  ( .A(counter[1]), .B(counter[0]), .CO(
        \add_83/carry[2] ), .S(N182) );
  HA_X1 \add_83/U1_1_2  ( .A(counter[2]), .B(\add_83/carry[2] ), .CO(
        \add_83/carry[3] ), .S(N183) );
  HA_X1 \add_83/U1_1_3  ( .A(counter[3]), .B(\add_83/carry[3] ), .CO(
        \add_83/carry[4] ), .S(N184) );
  HA_X1 \add_83/U1_1_4  ( .A(counter[4]), .B(\add_83/carry[4] ), .CO(
        \add_83/carry[5] ), .S(N185) );
  HA_X1 \add_80/U1_1_1  ( .A(counter2[1]), .B(counter2[0]), .CO(
        \add_80/carry[2] ), .S(N176) );
  HA_X1 \add_80/U1_1_2  ( .A(counter2[2]), .B(\add_80/carry[2] ), .CO(
        \add_80/carry[3] ), .S(N177) );
  HA_X1 \add_80/U1_1_3  ( .A(counter2[3]), .B(\add_80/carry[3] ), .CO(
        \add_80/carry[4] ), .S(N178) );
  HA_X1 \add_80/U1_1_4  ( .A(counter2[4]), .B(\add_80/carry[4] ), .CO(
        \add_80/carry[5] ), .S(N179) );
  DFF_X1 \state_reg[1]  ( .D(N201), .CK(clk), .Q(state[1]), .QN(n20) );
  DFF_X1 \counter2_reg[5]  ( .D(N215), .CK(clk), .Q(counter2[5]), .QN(n13) );
  DFF_X1 \state_reg[2]  ( .D(N202), .CK(clk), .Q(state[2]), .QN(n19) );
  DFF_X1 \counter_reg[5]  ( .D(n177), .CK(clk), .Q(counter[5]), .QN(n21) );
  DFF_X1 \counter_reg[4]  ( .D(n173), .CK(clk), .Q(counter[4]), .QN(n25) );
  DFF_X1 \counter_reg[3]  ( .D(n174), .CK(clk), .Q(counter[3]), .QN(n28) );
  DFF_X1 \counter_reg[2]  ( .D(n175), .CK(clk), .Q(counter[2]), .QN(n26) );
  DFF_X1 \counter_reg[1]  ( .D(n176), .CK(clk), .Q(counter[1]), .QN(n27) );
  DFF_X1 \counter_reg[0]  ( .D(n178), .CK(clk), .Q(counter[0]), .QN(N602) );
  DFF_X1 \counter2_reg[2]  ( .D(N212), .CK(clk), .Q(counter2[2]), .QN(n35) );
  DFF_X1 \counter2_reg[1]  ( .D(N211), .CK(clk), .Q(counter2[1]), .QN(n34) );
  DFF_X1 \counter2_reg[0]  ( .D(N210), .CK(clk), .Q(counter2[0]), .QN(N175) );
  DFF_X1 \counter2_reg[3]  ( .D(N213), .CK(clk), .Q(counter2[3]), .QN(n36) );
  DFF_X1 \counter2_reg[4]  ( .D(N214), .CK(clk), .Q(counter2[4]) );
  DFF_X1 \state_reg[0]  ( .D(N200), .CK(clk), .Q(state[0]) );
  NOR2_X1 U3 ( .A1(N608), .A2(N607), .ZN(n88) );
  OAI21_X1 U4 ( .B1(n38), .B2(n4), .A(n144), .ZN(\addr_a[1][2] ) );
  OAI21_X1 U5 ( .B1(n74), .B2(n4), .A(n144), .ZN(\addr_a[2][2] ) );
  OAI21_X1 U6 ( .B1(n64), .B2(n151), .A(n9), .ZN(\addr_a[3][2] ) );
  OAI21_X1 U7 ( .B1(n61), .B2(n151), .A(n9), .ZN(\addr_a[4][2] ) );
  OAI21_X1 U8 ( .B1(n58), .B2(n151), .A(n9), .ZN(\addr_a[5][2] ) );
  OAI21_X1 U9 ( .B1(n55), .B2(n151), .A(n9), .ZN(\addr_a[6][2] ) );
  OAI21_X1 U10 ( .B1(n51), .B2(n151), .A(n9), .ZN(\addr_a[7][2] ) );
  OAI21_X1 U11 ( .B1(n48), .B2(n151), .A(n9), .ZN(\addr_a[8][2] ) );
  OAI21_X1 U12 ( .B1(n43), .B2(n151), .A(n9), .ZN(\addr_a[9][2] ) );
  OAI21_X1 U13 ( .B1(n118), .B2(n4), .A(n144), .ZN(\addr_a[10][2] ) );
  OAI21_X1 U14 ( .B1(n116), .B2(n4), .A(n9), .ZN(\addr_a[11][2] ) );
  OAI21_X1 U15 ( .B1(n114), .B2(n4), .A(n9), .ZN(\addr_a[12][2] ) );
  OAI21_X1 U16 ( .B1(n112), .B2(n4), .A(n144), .ZN(\addr_a[13][2] ) );
  OAI21_X1 U17 ( .B1(n110), .B2(n4), .A(n144), .ZN(\addr_a[14][2] ) );
  OAI21_X1 U18 ( .B1(n108), .B2(n4), .A(n144), .ZN(\addr_a[15][2] ) );
  OAI21_X1 U19 ( .B1(n106), .B2(n4), .A(n144), .ZN(\addr_a[16][2] ) );
  OAI21_X1 U20 ( .B1(n104), .B2(n4), .A(n9), .ZN(\addr_a[17][2] ) );
  OAI21_X1 U21 ( .B1(n102), .B2(n4), .A(n9), .ZN(\addr_a[18][2] ) );
  OAI21_X1 U22 ( .B1(n100), .B2(n4), .A(n144), .ZN(\addr_a[19][2] ) );
  OAI21_X1 U23 ( .B1(n97), .B2(n151), .A(n144), .ZN(\addr_a[20][2] ) );
  OAI21_X1 U24 ( .B1(n95), .B2(n151), .A(n144), .ZN(\addr_a[21][2] ) );
  OAI21_X1 U25 ( .B1(n93), .B2(n151), .A(n144), .ZN(\addr_a[22][2] ) );
  OAI21_X1 U26 ( .B1(n90), .B2(n151), .A(n144), .ZN(\addr_a[23][2] ) );
  OAI21_X1 U27 ( .B1(n87), .B2(n151), .A(n144), .ZN(\addr_a[24][2] ) );
  OAI21_X1 U28 ( .B1(n85), .B2(n151), .A(n144), .ZN(\addr_a[25][2] ) );
  OAI21_X1 U29 ( .B1(n83), .B2(n151), .A(n144), .ZN(\addr_a[26][2] ) );
  OAI21_X1 U30 ( .B1(n81), .B2(n151), .A(n144), .ZN(\addr_a[27][2] ) );
  OAI21_X1 U31 ( .B1(n79), .B2(n4), .A(n144), .ZN(\addr_a[28][2] ) );
  OAI21_X1 U32 ( .B1(n77), .B2(n151), .A(n144), .ZN(\addr_a[29][2] ) );
  OAI21_X1 U33 ( .B1(n72), .B2(n151), .A(n144), .ZN(\addr_a[30][2] ) );
  OAI21_X1 U34 ( .B1(n67), .B2(n151), .A(n9), .ZN(\addr_a[31][2] ) );
  OAI21_X1 U35 ( .B1(n192), .B2(n143), .A(n9), .ZN(addr_x[2]) );
  OAI21_X1 U36 ( .B1(n40), .B2(n4), .A(n144), .ZN(\addr_a[0][2] ) );
  OAI21_X1 U37 ( .B1(n90), .B2(n7), .A(n140), .ZN(\addr_a[23][4] ) );
  OAI21_X1 U38 ( .B1(n72), .B2(n7), .A(n140), .ZN(\addr_a[30][4] ) );
  OAI21_X1 U39 ( .B1(n67), .B2(n7), .A(n12), .ZN(\addr_a[31][4] ) );
  OAI21_X1 U40 ( .B1(n40), .B2(n149), .A(n140), .ZN(\addr_a[0][4] ) );
  BUF_X1 U41 ( .A(n39), .Z(n16) );
  BUF_X1 U42 ( .A(n144), .Z(n9) );
  BUF_X1 U43 ( .A(n142), .Z(n11) );
  BUF_X1 U44 ( .A(n140), .Z(n12) );
  BUF_X1 U45 ( .A(n147), .Z(n8) );
  BUF_X1 U46 ( .A(n142), .Z(n10) );
  BUF_X1 U47 ( .A(n41), .Z(n15) );
  OAI21_X1 U48 ( .B1(n48), .B2(n149), .A(n12), .ZN(\addr_a[8][4] ) );
  OAI21_X1 U49 ( .B1(n43), .B2(n149), .A(n12), .ZN(\addr_a[9][4] ) );
  OAI21_X1 U50 ( .B1(n87), .B2(n7), .A(n140), .ZN(\addr_a[24][4] ) );
  OAI21_X1 U51 ( .B1(n85), .B2(n7), .A(n140), .ZN(\addr_a[25][4] ) );
  OAI21_X1 U52 ( .B1(n81), .B2(n7), .A(n140), .ZN(\addr_a[27][4] ) );
  OAI21_X1 U53 ( .B1(n79), .B2(n7), .A(n140), .ZN(\addr_a[28][4] ) );
  OAI21_X1 U54 ( .B1(n77), .B2(n7), .A(n140), .ZN(\addr_a[29][4] ) );
  OAI21_X1 U55 ( .B1(n106), .B2(n149), .A(n140), .ZN(\addr_a[16][4] ) );
  OAI21_X1 U56 ( .B1(n104), .B2(n149), .A(n12), .ZN(\addr_a[17][4] ) );
  OAI21_X1 U57 ( .B1(n102), .B2(n149), .A(n140), .ZN(\addr_a[18][4] ) );
  OAI21_X1 U58 ( .B1(n100), .B2(n149), .A(n140), .ZN(\addr_a[19][4] ) );
  OAI21_X1 U59 ( .B1(n97), .B2(n7), .A(n140), .ZN(\addr_a[20][4] ) );
  OAI21_X1 U60 ( .B1(n95), .B2(n7), .A(n140), .ZN(\addr_a[21][4] ) );
  OAI21_X1 U61 ( .B1(n93), .B2(n7), .A(n140), .ZN(\addr_a[22][4] ) );
  OAI21_X1 U62 ( .B1(n38), .B2(n149), .A(n140), .ZN(\addr_a[1][4] ) );
  OAI21_X1 U63 ( .B1(n74), .B2(n7), .A(n140), .ZN(\addr_a[2][4] ) );
  OAI21_X1 U64 ( .B1(n64), .B2(n149), .A(n12), .ZN(\addr_a[3][4] ) );
  OAI21_X1 U65 ( .B1(n61), .B2(n149), .A(n12), .ZN(\addr_a[4][4] ) );
  OAI21_X1 U66 ( .B1(n58), .B2(n149), .A(n12), .ZN(\addr_a[5][4] ) );
  OAI21_X1 U67 ( .B1(n55), .B2(n149), .A(n12), .ZN(\addr_a[6][4] ) );
  OAI21_X1 U68 ( .B1(n51), .B2(n149), .A(n12), .ZN(\addr_a[7][4] ) );
  OAI21_X1 U69 ( .B1(n118), .B2(n149), .A(n12), .ZN(\addr_a[10][4] ) );
  OAI21_X1 U70 ( .B1(n116), .B2(n7), .A(n140), .ZN(\addr_a[11][4] ) );
  OAI21_X1 U71 ( .B1(n114), .B2(n149), .A(n12), .ZN(\addr_a[12][4] ) );
  OAI21_X1 U72 ( .B1(n112), .B2(n149), .A(n140), .ZN(\addr_a[13][4] ) );
  OAI21_X1 U73 ( .B1(n110), .B2(n149), .A(n140), .ZN(\addr_a[14][4] ) );
  OAI21_X1 U74 ( .B1(n108), .B2(n149), .A(n140), .ZN(\addr_a[15][4] ) );
  OAI21_X1 U75 ( .B1(n83), .B2(n7), .A(n140), .ZN(\addr_a[26][4] ) );
  BUF_X1 U76 ( .A(n152), .Z(n3) );
  BUF_X1 U77 ( .A(n153), .Z(n2) );
  BUF_X1 U78 ( .A(n151), .Z(n4) );
  BUF_X1 U79 ( .A(n150), .Z(n6) );
  BUF_X1 U80 ( .A(n150), .Z(n5) );
  BUF_X1 U81 ( .A(n149), .Z(n7) );
  OAI21_X1 U82 ( .B1(n48), .B2(n3), .A(n39), .ZN(\addr_a[8][1] ) );
  OAI21_X1 U83 ( .B1(n48), .B2(n153), .A(n147), .ZN(\addr_a[8][0] ) );
  OAI21_X1 U84 ( .B1(n43), .B2(n152), .A(n39), .ZN(\addr_a[9][1] ) );
  OAI21_X1 U85 ( .B1(n43), .B2(n153), .A(n147), .ZN(\addr_a[9][0] ) );
  OAI21_X1 U86 ( .B1(n67), .B2(n152), .A(n39), .ZN(\addr_a[31][1] ) );
  OAI21_X1 U87 ( .B1(n67), .B2(n153), .A(n147), .ZN(\addr_a[31][0] ) );
  OAI21_X1 U88 ( .B1(n87), .B2(n3), .A(n16), .ZN(\addr_a[24][1] ) );
  OAI21_X1 U89 ( .B1(n87), .B2(n2), .A(n8), .ZN(\addr_a[24][0] ) );
  OAI21_X1 U90 ( .B1(n85), .B2(n3), .A(n16), .ZN(\addr_a[25][1] ) );
  OAI21_X1 U91 ( .B1(n85), .B2(n2), .A(n8), .ZN(\addr_a[25][0] ) );
  OAI21_X1 U92 ( .B1(n81), .B2(n3), .A(n16), .ZN(\addr_a[27][1] ) );
  OAI21_X1 U93 ( .B1(n81), .B2(n2), .A(n8), .ZN(\addr_a[27][0] ) );
  OAI21_X1 U94 ( .B1(n79), .B2(n3), .A(n16), .ZN(\addr_a[28][1] ) );
  OAI21_X1 U95 ( .B1(n79), .B2(n2), .A(n8), .ZN(\addr_a[28][0] ) );
  OAI21_X1 U96 ( .B1(n77), .B2(n3), .A(n39), .ZN(\addr_a[29][1] ) );
  OAI21_X1 U97 ( .B1(n77), .B2(n2), .A(n8), .ZN(\addr_a[29][0] ) );
  OAI21_X1 U98 ( .B1(n72), .B2(n3), .A(n39), .ZN(\addr_a[30][1] ) );
  OAI21_X1 U99 ( .B1(n72), .B2(n2), .A(n8), .ZN(\addr_a[30][0] ) );
  OAI21_X1 U100 ( .B1(n106), .B2(n152), .A(n39), .ZN(\addr_a[16][1] ) );
  OAI21_X1 U101 ( .B1(n106), .B2(n153), .A(n147), .ZN(\addr_a[16][0] ) );
  OAI21_X1 U102 ( .B1(n104), .B2(n152), .A(n16), .ZN(\addr_a[17][1] ) );
  OAI21_X1 U104 ( .B1(n104), .B2(n2), .A(n8), .ZN(\addr_a[17][0] ) );
  OAI21_X1 U105 ( .B1(n102), .B2(n152), .A(n16), .ZN(\addr_a[18][1] ) );
  OAI21_X1 U106 ( .B1(n102), .B2(n153), .A(n147), .ZN(\addr_a[18][0] ) );
  OAI21_X1 U107 ( .B1(n100), .B2(n152), .A(n16), .ZN(\addr_a[19][1] ) );
  OAI21_X1 U109 ( .B1(n100), .B2(n153), .A(n147), .ZN(\addr_a[19][0] ) );
  OAI21_X1 U110 ( .B1(n97), .B2(n3), .A(n16), .ZN(\addr_a[20][1] ) );
  OAI21_X1 U111 ( .B1(n97), .B2(n2), .A(n8), .ZN(\addr_a[20][0] ) );
  OAI21_X1 U112 ( .B1(n95), .B2(n3), .A(n16), .ZN(\addr_a[21][1] ) );
  OAI21_X1 U113 ( .B1(n95), .B2(n2), .A(n8), .ZN(\addr_a[21][0] ) );
  OAI21_X1 U115 ( .B1(n93), .B2(n3), .A(n16), .ZN(\addr_a[22][1] ) );
  OAI21_X1 U116 ( .B1(n93), .B2(n2), .A(n8), .ZN(\addr_a[22][0] ) );
  OAI21_X1 U117 ( .B1(n90), .B2(n3), .A(n16), .ZN(\addr_a[23][1] ) );
  OAI21_X1 U118 ( .B1(n90), .B2(n2), .A(n8), .ZN(\addr_a[23][0] ) );
  OAI21_X1 U119 ( .B1(n40), .B2(n3), .A(n39), .ZN(\addr_a[0][1] ) );
  OAI21_X1 U121 ( .B1(n40), .B2(n153), .A(n147), .ZN(\addr_a[0][0] ) );
  OAI21_X1 U122 ( .B1(n74), .B2(n3), .A(n39), .ZN(\addr_a[2][1] ) );
  OAI21_X1 U123 ( .B1(n74), .B2(n2), .A(n8), .ZN(\addr_a[2][0] ) );
  OAI21_X1 U124 ( .B1(n38), .B2(n152), .A(n16), .ZN(\addr_a[1][1] ) );
  OAI21_X1 U125 ( .B1(n38), .B2(n153), .A(n147), .ZN(\addr_a[1][0] ) );
  OAI21_X1 U127 ( .B1(n64), .B2(n152), .A(n39), .ZN(\addr_a[3][1] ) );
  OAI21_X1 U128 ( .B1(n64), .B2(n153), .A(n147), .ZN(\addr_a[3][0] ) );
  OAI21_X1 U129 ( .B1(n61), .B2(n152), .A(n39), .ZN(\addr_a[4][1] ) );
  OAI21_X1 U130 ( .B1(n61), .B2(n153), .A(n147), .ZN(\addr_a[4][0] ) );
  OAI21_X1 U131 ( .B1(n58), .B2(n152), .A(n39), .ZN(\addr_a[5][1] ) );
  OAI21_X1 U133 ( .B1(n58), .B2(n153), .A(n147), .ZN(\addr_a[5][0] ) );
  OAI21_X1 U134 ( .B1(n55), .B2(n152), .A(n16), .ZN(\addr_a[6][1] ) );
  OAI21_X1 U135 ( .B1(n55), .B2(n153), .A(n147), .ZN(\addr_a[6][0] ) );
  OAI21_X1 U136 ( .B1(n51), .B2(n152), .A(n39), .ZN(\addr_a[7][1] ) );
  OAI21_X1 U137 ( .B1(n51), .B2(n2), .A(n147), .ZN(\addr_a[7][0] ) );
  OAI21_X1 U139 ( .B1(n118), .B2(n152), .A(n39), .ZN(\addr_a[10][1] ) );
  OAI21_X1 U140 ( .B1(n118), .B2(n153), .A(n147), .ZN(\addr_a[10][0] ) );
  OAI21_X1 U141 ( .B1(n116), .B2(n152), .A(n39), .ZN(\addr_a[11][1] ) );
  OAI21_X1 U142 ( .B1(n116), .B2(n153), .A(n147), .ZN(\addr_a[11][0] ) );
  OAI21_X1 U143 ( .B1(n114), .B2(n152), .A(n39), .ZN(\addr_a[12][1] ) );
  OAI21_X1 U145 ( .B1(n114), .B2(n153), .A(n147), .ZN(\addr_a[12][0] ) );
  OAI21_X1 U146 ( .B1(n112), .B2(n152), .A(n39), .ZN(\addr_a[13][1] ) );
  OAI21_X1 U147 ( .B1(n112), .B2(n153), .A(n147), .ZN(\addr_a[13][0] ) );
  OAI21_X1 U148 ( .B1(n110), .B2(n152), .A(n39), .ZN(\addr_a[14][1] ) );
  OAI21_X1 U149 ( .B1(n110), .B2(n153), .A(n147), .ZN(\addr_a[14][0] ) );
  OAI21_X1 U151 ( .B1(n108), .B2(n152), .A(n39), .ZN(\addr_a[15][1] ) );
  OAI21_X1 U152 ( .B1(n108), .B2(n153), .A(n147), .ZN(\addr_a[15][0] ) );
  OAI21_X1 U153 ( .B1(n83), .B2(n3), .A(n16), .ZN(\addr_a[26][1] ) );
  OAI21_X1 U154 ( .B1(n83), .B2(n2), .A(n8), .ZN(\addr_a[26][0] ) );
  NAND2_X1 U155 ( .A1(n46), .A2(n184), .ZN(n41) );
  NAND2_X1 U157 ( .A1(n186), .A2(n190), .ZN(n39) );
  NAND2_X1 U158 ( .A1(n185), .A2(n190), .ZN(n147) );
  NAND2_X1 U159 ( .A1(n187), .A2(n190), .ZN(n144) );
  NAND2_X1 U160 ( .A1(n188), .A2(n190), .ZN(n142) );
  NAND2_X1 U161 ( .A1(n189), .A2(n190), .ZN(n140) );
  OR3_X1 U163 ( .A1(n70), .A2(n53), .A3(n184), .ZN(n69) );
  INV_X1 U164 ( .A(N606), .ZN(n196) );
  OAI21_X1 U165 ( .B1(n192), .B2(n139), .A(n12), .ZN(addr_x[4]) );
  NOR2_X1 U166 ( .A1(n198), .A2(N173), .ZN(n123) );
  NAND2_X1 U168 ( .A1(n154), .A2(n156), .ZN(n48) );
  NAND2_X1 U169 ( .A1(n154), .A2(n155), .ZN(n43) );
  NAND2_X1 U170 ( .A1(n163), .A2(n157), .ZN(n67) );
  NAND2_X1 U171 ( .A1(n163), .A2(n156), .ZN(n87) );
  NAND2_X1 U172 ( .A1(n163), .A2(n155), .ZN(n85) );
  NAND2_X1 U174 ( .A1(n163), .A2(n162), .ZN(n81) );
  NAND2_X1 U175 ( .A1(n163), .A2(n161), .ZN(n79) );
  NAND2_X1 U176 ( .A1(n163), .A2(n160), .ZN(n77) );
  NAND2_X1 U177 ( .A1(n163), .A2(n159), .ZN(n72) );
  NAND2_X1 U178 ( .A1(n165), .A2(n156), .ZN(n106) );
  NAND2_X1 U180 ( .A1(n165), .A2(n155), .ZN(n104) );
  NAND2_X1 U181 ( .A1(n165), .A2(n164), .ZN(n102) );
  NAND2_X1 U182 ( .A1(n165), .A2(n162), .ZN(n100) );
  NAND2_X1 U183 ( .A1(n165), .A2(n161), .ZN(n97) );
  NAND2_X1 U184 ( .A1(n165), .A2(n160), .ZN(n95) );
  NAND2_X1 U186 ( .A1(n165), .A2(n159), .ZN(n93) );
  NAND2_X1 U187 ( .A1(n165), .A2(n157), .ZN(n90) );
  NAND2_X1 U188 ( .A1(n156), .A2(n158), .ZN(n40) );
  NAND2_X1 U189 ( .A1(n164), .A2(n158), .ZN(n74) );
  NAND2_X1 U190 ( .A1(n155), .A2(n158), .ZN(n38) );
  BUF_X1 U192 ( .A(n46), .Z(n14) );
  NAND2_X1 U193 ( .A1(n162), .A2(n158), .ZN(n64) );
  NAND2_X1 U194 ( .A1(n161), .A2(n158), .ZN(n61) );
  NAND2_X1 U195 ( .A1(n160), .A2(n158), .ZN(n58) );
  NAND2_X1 U196 ( .A1(n159), .A2(n158), .ZN(n55) );
  NAND2_X1 U198 ( .A1(n157), .A2(n158), .ZN(n51) );
  NAND2_X1 U199 ( .A1(n164), .A2(n154), .ZN(n118) );
  NAND2_X1 U200 ( .A1(n162), .A2(n154), .ZN(n116) );
  NAND2_X1 U201 ( .A1(n161), .A2(n154), .ZN(n114) );
  NAND2_X1 U203 ( .A1(n160), .A2(n154), .ZN(n112) );
  NAND2_X1 U205 ( .A1(n159), .A2(n154), .ZN(n110) );
  NAND2_X1 U206 ( .A1(n157), .A2(n154), .ZN(n108) );
  NAND2_X1 U207 ( .A1(n164), .A2(n163), .ZN(n83) );
  INV_X1 U208 ( .A(n148), .ZN(n192) );
  NOR3_X1 U209 ( .A1(n184), .A2(n166), .A3(n74), .ZN(done) );
  INV_X1 U211 ( .A(n166), .ZN(n190) );
  NAND2_X1 U212 ( .A1(n68), .A2(n186), .ZN(n152) );
  OAI21_X1 U213 ( .B1(n192), .B2(n146), .A(n147), .ZN(addr_x[0]) );
  OAI21_X1 U214 ( .B1(n145), .B2(n192), .A(n39), .ZN(addr_x[1]) );
  AND2_X1 U215 ( .A1(N173), .A2(n129), .ZN(n167) );
  INV_X1 U217 ( .A(n138), .ZN(n184) );
  INV_X1 U218 ( .A(N604), .ZN(n195) );
  INV_X1 U219 ( .A(N603), .ZN(n194) );
  NAND2_X1 U220 ( .A1(n185), .A2(n68), .ZN(n153) );
  NAND2_X1 U221 ( .A1(n187), .A2(n68), .ZN(n151) );
  NAND2_X1 U223 ( .A1(n188), .A2(n68), .ZN(n150) );
  NAND2_X1 U224 ( .A1(n189), .A2(n68), .ZN(n149) );
  OR2_X1 U225 ( .A1(n198), .A2(n171), .ZN(n130) );
  INV_X1 U226 ( .A(n146), .ZN(n185) );
  INV_X1 U227 ( .A(n143), .ZN(n187) );
  INV_X1 U229 ( .A(n141), .ZN(n188) );
  INV_X1 U230 ( .A(n139), .ZN(n189) );
  INV_X1 U231 ( .A(n145), .ZN(n186) );
  INV_X1 U232 ( .A(n17), .ZN(n29) );
  AND2_X1 U233 ( .A1(N176), .A2(n167), .ZN(N211) );
  AND2_X1 U235 ( .A1(N177), .A2(n167), .ZN(N212) );
  AND2_X1 U236 ( .A1(N178), .A2(n167), .ZN(N213) );
  AND2_X1 U237 ( .A1(N179), .A2(n167), .ZN(N214) );
  INV_X1 U238 ( .A(n131), .ZN(n193) );
  NAND2_X1 U239 ( .A1(n193), .A2(n138), .ZN(n132) );
  INV_X1 U241 ( .A(n129), .ZN(n198) );
  NAND2_X1 U242 ( .A1(n132), .A2(n137), .ZN(addr_y[0]) );
  NAND2_X1 U243 ( .A1(N175), .A2(n193), .ZN(n137) );
  INV_X1 U244 ( .A(n30), .ZN(n179) );
  INV_X1 U245 ( .A(n32), .ZN(n181) );
  INV_X1 U247 ( .A(n31), .ZN(n180) );
  AND3_X1 U248 ( .A1(n193), .A2(n184), .A3(N1175), .ZN(addr_y[5]) );
  NOR3_X1 U249 ( .A1(counter[1]), .A2(counter[2]), .A3(counter[0]), .ZN(n156)
         );
  NOR3_X1 U250 ( .A1(counter[1]), .A2(counter[2]), .A3(N602), .ZN(n155) );
  NOR3_X1 U251 ( .A1(N602), .A2(counter[2]), .A3(n27), .ZN(n162) );
  NOR3_X1 U252 ( .A1(counter[0]), .A2(counter[1]), .A3(n26), .ZN(n161) );
  NOR3_X1 U254 ( .A1(N602), .A2(counter[1]), .A3(n26), .ZN(n160) );
  NOR3_X1 U255 ( .A1(n27), .A2(counter[0]), .A3(n26), .ZN(n159) );
  NOR3_X1 U256 ( .A1(n27), .A2(N602), .A3(n26), .ZN(n157) );
  NOR3_X1 U257 ( .A1(counter[0]), .A2(counter[2]), .A3(n27), .ZN(n164) );
  NOR4_X1 U259 ( .A1(counter2[1]), .A2(counter2[2]), .A3(counter2[0]), .A4(
        n172), .ZN(n138) );
  OR3_X1 U261 ( .A1(counter2[3]), .A2(counter2[5]), .A3(counter2[4]), .ZN(n172) );
  NOR2_X1 U262 ( .A1(n120), .A2(counter[5]), .ZN(n68) );
  NOR4_X1 U263 ( .A1(n37), .A2(n38), .A3(counter2[0]), .A4(n39), .ZN(wr_en_y)
         );
  OR3_X1 U264 ( .A1(counter2[3]), .A2(counter2[4]), .A3(counter2[2]), .ZN(n37)
         );
  AOI221_X1 U265 ( .B1(n40), .B2(n148), .C1(n191), .C2(counter[5]), .A(done), 
        .ZN(n171) );
  INV_X1 U266 ( .A(n120), .ZN(n191) );
  NOR3_X1 U268 ( .A1(state[1]), .A2(state[2]), .A3(state[0]), .ZN(n148) );
  OAI221_X1 U269 ( .B1(n168), .B2(n130), .C1(n198), .C2(n19), .A(n197), .ZN(
        N202) );
  OAI221_X1 U270 ( .B1(n166), .B2(n130), .C1(reset), .C2(n199), .A(n170), .ZN(
        N200) );
  INV_X1 U271 ( .A(n24), .ZN(N607) );
  INV_X1 U272 ( .A(n66), .ZN(wr_en_a[31]) );
  OAI211_X1 U273 ( .C1(n13), .C2(n67), .A(n68), .B(n69), .ZN(n66) );
  AOI21_X1 U275 ( .B1(n41), .B2(n98), .A(n38), .ZN(wr_en_a[1]) );
  OAI21_X1 U276 ( .B1(n45), .B2(n52), .A(n14), .ZN(n98) );
  AOI21_X1 U277 ( .B1(n15), .B2(n73), .A(n74), .ZN(wr_en_a[2]) );
  OAI21_X1 U278 ( .B1(n52), .B2(n75), .A(n46), .ZN(n73) );
  AOI21_X1 U279 ( .B1(n41), .B2(n63), .A(n64), .ZN(wr_en_a[3]) );
  OAI21_X1 U280 ( .B1(n52), .B2(n65), .A(n14), .ZN(n63) );
  AOI21_X1 U282 ( .B1(n41), .B2(n60), .A(n61), .ZN(wr_en_a[4]) );
  OAI21_X1 U283 ( .B1(n52), .B2(n62), .A(n14), .ZN(n60) );
  AOI21_X1 U284 ( .B1(n15), .B2(n57), .A(n58), .ZN(wr_en_a[5]) );
  OAI21_X1 U285 ( .B1(n52), .B2(n59), .A(n14), .ZN(n57) );
  AOI21_X1 U286 ( .B1(n41), .B2(n54), .A(n55), .ZN(wr_en_a[6]) );
  OAI21_X1 U287 ( .B1(n52), .B2(n56), .A(n14), .ZN(n54) );
  AOI21_X1 U289 ( .B1(n41), .B2(n50), .A(n51), .ZN(wr_en_a[7]) );
  OAI21_X1 U290 ( .B1(n52), .B2(n53), .A(n14), .ZN(n50) );
  AOI21_X1 U291 ( .B1(n41), .B2(n47), .A(n48), .ZN(wr_en_a[8]) );
  OAI21_X1 U292 ( .B1(n44), .B2(n49), .A(n14), .ZN(n47) );
  AOI21_X1 U293 ( .B1(n15), .B2(n42), .A(n43), .ZN(wr_en_a[9]) );
  OAI21_X1 U294 ( .B1(n44), .B2(n45), .A(n14), .ZN(n42) );
  AOI21_X1 U296 ( .B1(n41), .B2(n117), .A(n118), .ZN(wr_en_a[10]) );
  OAI21_X1 U297 ( .B1(n44), .B2(n75), .A(n46), .ZN(n117) );
  AOI21_X1 U298 ( .B1(n41), .B2(n115), .A(n116), .ZN(wr_en_a[11]) );
  OAI21_X1 U299 ( .B1(n44), .B2(n65), .A(n14), .ZN(n115) );
  AOI21_X1 U301 ( .B1(n41), .B2(n113), .A(n114), .ZN(wr_en_a[12]) );
  OAI21_X1 U302 ( .B1(n44), .B2(n62), .A(n46), .ZN(n113) );
  AOI21_X1 U303 ( .B1(n41), .B2(n111), .A(n112), .ZN(wr_en_a[13]) );
  OAI21_X1 U304 ( .B1(n44), .B2(n59), .A(n46), .ZN(n111) );
  AOI21_X1 U306 ( .B1(n41), .B2(n109), .A(n110), .ZN(wr_en_a[14]) );
  OAI21_X1 U307 ( .B1(n44), .B2(n56), .A(n46), .ZN(n109) );
  AOI21_X1 U308 ( .B1(n41), .B2(n107), .A(n108), .ZN(wr_en_a[15]) );
  OAI21_X1 U309 ( .B1(n44), .B2(n53), .A(n46), .ZN(n107) );
  AOI21_X1 U310 ( .B1(n41), .B2(n105), .A(n106), .ZN(wr_en_a[16]) );
  OAI21_X1 U311 ( .B1(n49), .B2(n91), .A(n14), .ZN(n105) );
  AOI21_X1 U312 ( .B1(n41), .B2(n103), .A(n104), .ZN(wr_en_a[17]) );
  OAI21_X1 U313 ( .B1(n45), .B2(n91), .A(n14), .ZN(n103) );
  AOI21_X1 U314 ( .B1(n41), .B2(n101), .A(n102), .ZN(wr_en_a[18]) );
  OAI21_X1 U315 ( .B1(n75), .B2(n91), .A(n14), .ZN(n101) );
  AOI21_X1 U316 ( .B1(n41), .B2(n99), .A(n100), .ZN(wr_en_a[19]) );
  OAI21_X1 U317 ( .B1(n65), .B2(n91), .A(n14), .ZN(n99) );
  AOI21_X1 U318 ( .B1(n15), .B2(n96), .A(n97), .ZN(wr_en_a[20]) );
  OAI21_X1 U319 ( .B1(n62), .B2(n91), .A(n14), .ZN(n96) );
  AOI21_X1 U320 ( .B1(n15), .B2(n94), .A(n95), .ZN(wr_en_a[21]) );
  OAI21_X1 U321 ( .B1(n59), .B2(n91), .A(n14), .ZN(n94) );
  AOI21_X1 U322 ( .B1(n15), .B2(n92), .A(n93), .ZN(wr_en_a[22]) );
  OAI21_X1 U323 ( .B1(n56), .B2(n91), .A(n14), .ZN(n92) );
  AOI21_X1 U324 ( .B1(n15), .B2(n89), .A(n90), .ZN(wr_en_a[23]) );
  OAI21_X1 U325 ( .B1(n53), .B2(n91), .A(n14), .ZN(n89) );
  AOI21_X1 U326 ( .B1(n15), .B2(n86), .A(n87), .ZN(wr_en_a[24]) );
  OAI21_X1 U327 ( .B1(n49), .B2(n70), .A(n14), .ZN(n86) );
  AOI21_X1 U328 ( .B1(n15), .B2(n84), .A(n85), .ZN(wr_en_a[25]) );
  OAI21_X1 U329 ( .B1(n45), .B2(n70), .A(n14), .ZN(n84) );
  AOI21_X1 U330 ( .B1(n15), .B2(n82), .A(n83), .ZN(wr_en_a[26]) );
  OAI21_X1 U331 ( .B1(n70), .B2(n75), .A(n14), .ZN(n82) );
  AOI21_X1 U332 ( .B1(n15), .B2(n80), .A(n81), .ZN(wr_en_a[27]) );
  OAI21_X1 U333 ( .B1(n65), .B2(n70), .A(n46), .ZN(n80) );
  AOI21_X1 U334 ( .B1(n15), .B2(n78), .A(n79), .ZN(wr_en_a[28]) );
  OAI21_X1 U335 ( .B1(n62), .B2(n70), .A(n46), .ZN(n78) );
  AOI21_X1 U336 ( .B1(n15), .B2(n76), .A(n77), .ZN(wr_en_a[29]) );
  OAI21_X1 U337 ( .B1(n59), .B2(n70), .A(n46), .ZN(n76) );
  AOI21_X1 U338 ( .B1(n15), .B2(n71), .A(n72), .ZN(wr_en_a[30]) );
  OAI21_X1 U339 ( .B1(n56), .B2(n70), .A(n46), .ZN(n71) );
  AOI21_X1 U340 ( .B1(n15), .B2(n119), .A(n40), .ZN(wr_en_a[0]) );
  OAI21_X1 U341 ( .B1(n49), .B2(n52), .A(n14), .ZN(n119) );
  NOR2_X1 U343 ( .A1(n40), .A2(n192), .ZN(wr_en_x) );
  NAND4_X1 U344 ( .A1(n131), .A2(n120), .A3(n192), .A4(n19), .ZN(clear_acc) );
  NOR2_X1 U345 ( .A1(n20), .A2(state[0]), .ZN(n168) );
  NOR2_X1 U346 ( .A1(n120), .A2(counter2[5]), .ZN(n46) );
  AND2_X1 U347 ( .A1(N180), .A2(n167), .ZN(N215) );
  NAND2_X1 U348 ( .A1(counter2[0]), .A2(n13), .ZN(n146) );
  OAI21_X1 U349 ( .B1(n25), .B2(n121), .A(n122), .ZN(n173) );
  NAND2_X1 U350 ( .A1(N185), .A2(n123), .ZN(n122) );
  OAI21_X1 U351 ( .B1(n28), .B2(n121), .A(n124), .ZN(n174) );
  NAND2_X1 U352 ( .A1(N184), .A2(n123), .ZN(n124) );
  OAI21_X1 U353 ( .B1(n26), .B2(n121), .A(n125), .ZN(n175) );
  NAND2_X1 U354 ( .A1(N183), .A2(n123), .ZN(n125) );
  OAI21_X1 U355 ( .B1(n27), .B2(n121), .A(n126), .ZN(n176) );
  NAND2_X1 U356 ( .A1(N182), .A2(n123), .ZN(n126) );
  OAI21_X1 U357 ( .B1(N602), .B2(n121), .A(n128), .ZN(n178) );
  NAND2_X1 U358 ( .A1(N602), .A2(n123), .ZN(n128) );
  OAI21_X1 U359 ( .B1(n21), .B2(n121), .A(n127), .ZN(n177) );
  NAND2_X1 U360 ( .A1(N186), .A2(n123), .ZN(n127) );
  NAND2_X1 U361 ( .A1(n168), .A2(n19), .ZN(n166) );
  NAND2_X1 U362 ( .A1(counter2[2]), .A2(n13), .ZN(n143) );
  NAND2_X1 U363 ( .A1(counter2[3]), .A2(n13), .ZN(n141) );
  NAND2_X1 U364 ( .A1(counter2[4]), .A2(n13), .ZN(n139) );
  NAND2_X1 U365 ( .A1(counter2[1]), .A2(n13), .ZN(n145) );
  INV_X1 U366 ( .A(n18), .ZN(N605) );
  OR2_X1 U384 ( .A1(n29), .A2(counter[2]), .ZN(n1) );
  AND2_X1 U385 ( .A1(N175), .A2(n167), .ZN(N210) );
  OAI21_X1 U386 ( .B1(n20), .B2(n198), .A(n169), .ZN(N201) );
  NAND4_X1 U387 ( .A1(start), .A2(n199), .A3(n200), .A4(n197), .ZN(n169) );
  INV_X1 U388 ( .A(loadVector), .ZN(n200) );
  NOR4_X1 U389 ( .A1(loadMatrix), .A2(loadVector), .A3(reset), .A4(start), 
        .ZN(n129) );
  NAND2_X1 U390 ( .A1(n132), .A2(n133), .ZN(addr_y[4]) );
  NAND2_X1 U391 ( .A1(N1174), .A2(n193), .ZN(n133) );
  NAND2_X1 U392 ( .A1(n132), .A2(n135), .ZN(addr_y[2]) );
  NAND2_X1 U393 ( .A1(N1172), .A2(n193), .ZN(n135) );
  NAND2_X1 U394 ( .A1(n132), .A2(n134), .ZN(addr_y[3]) );
  NAND2_X1 U395 ( .A1(N1173), .A2(n193), .ZN(n134) );
  INV_X1 U396 ( .A(reset), .ZN(n197) );
  NAND2_X1 U397 ( .A1(n132), .A2(n136), .ZN(addr_y[1]) );
  NAND2_X1 U398 ( .A1(N1171), .A2(n193), .ZN(n136) );
  INV_X1 U399 ( .A(loadMatrix), .ZN(n199) );
  XOR2_X1 U400 ( .A(\add_80/carry[5] ), .B(counter2[5]), .Z(N180) );
  XOR2_X1 U401 ( .A(\add_83/carry[5] ), .B(counter[5]), .Z(N186) );
  NOR2_X1 U402 ( .A1(counter[1]), .A2(counter[0]), .ZN(n17) );
  OAI21_X1 U403 ( .B1(N602), .B2(n27), .A(n29), .ZN(N603) );
  OAI21_X1 U404 ( .B1(n17), .B2(n26), .A(n1), .ZN(N604) );
  NOR2_X1 U405 ( .A1(n1), .A2(counter[3]), .ZN(n22) );
  AOI21_X1 U406 ( .B1(n1), .B2(counter[3]), .A(n22), .ZN(n18) );
  NAND2_X1 U407 ( .A1(n22), .A2(n25), .ZN(n23) );
  OAI21_X1 U408 ( .B1(n22), .B2(n25), .A(n23), .ZN(N606) );
  NOR2_X1 U409 ( .A1(n23), .A2(counter[5]), .ZN(N608) );
  AOI21_X1 U410 ( .B1(n23), .B2(counter[5]), .A(N608), .ZN(n24) );
  NOR2_X1 U411 ( .A1(counter2[1]), .A2(counter2[0]), .ZN(n30) );
  OAI21_X1 U412 ( .B1(N175), .B2(n34), .A(n179), .ZN(N1171) );
  NOR2_X1 U413 ( .A1(n179), .A2(counter2[2]), .ZN(n31) );
  OAI21_X1 U414 ( .B1(n30), .B2(n35), .A(n180), .ZN(N1172) );
  NOR2_X1 U415 ( .A1(n180), .A2(counter2[3]), .ZN(n32) );
  OAI21_X1 U416 ( .B1(n31), .B2(n36), .A(n181), .ZN(N1173) );
  XOR2_X1 U417 ( .A(counter2[4]), .B(n32), .Z(N1174) );
  NOR2_X1 U418 ( .A1(counter2[4]), .A2(n181), .ZN(n33) );
  XOR2_X1 U419 ( .A(counter2[5]), .B(n33), .Z(N1175) );
  AND4_X1 U420 ( .A1(counter2[3]), .A2(counter2[2]), .A3(counter2[1]), .A4(
        counter2[0]), .ZN(n182) );
  OAI22_X1 U421 ( .A1(counter2[5]), .A2(n182), .B1(counter2[5]), .B2(
        counter2[4]), .ZN(N173) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_32 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N18, N20, N21, N22,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n629), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n630), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n631), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n632), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n633), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n634), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n635), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n636), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n637), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n638), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n639), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n640), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n641), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n642), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n643), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n644), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n645), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n646), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n647), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n648), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n649), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n650), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n651), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n652), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n653), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n654), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n655), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n656), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n657), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n658), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n659), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n660), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n661), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n662), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n663), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n664), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n665), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n666), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n667), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n668), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n669), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n670), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n671), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n672), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n673), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n674), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n675), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n676), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n677), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n678), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n679), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n680), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n681), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n682), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n683), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n684), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n685), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n686), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n687), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n688), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n689), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n690), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n691), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n692), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n693), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n694), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n695), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n696), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n697), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n698), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n699), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n700), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n701), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n702), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n703), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n704), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n705), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n706), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n707), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n708), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n709), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n710), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n711), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n712), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n713), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n714), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n715), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n716), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n717), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n718), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n719), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n720), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n721), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n722), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n723), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n724), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n725), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n726), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n727), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n728), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n729), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n730), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n731), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n732), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n733), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n734), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n735), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n736), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n737), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n738), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n739), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n740), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n741), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n742), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n743), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n744), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n745), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n746), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n747), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n748), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n749), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n750), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n751), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n752), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n753), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n754), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n755), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n756), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n757), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n758), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n759), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n760), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n761), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n762), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n763), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n764), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n765), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n766), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n767), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n768), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n769), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n770), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n771), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n772), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n773), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n774), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n775), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n776), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n777), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n778), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n779), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n780), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n781), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n782), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n783), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n784), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n785), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n786), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n787), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n788), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n789), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n790), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n791), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n792), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n793), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n794), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n795), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n796), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n797), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n798), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n799), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n800), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n801), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n802), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n803), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n804), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n805), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n806), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n807), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n808), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n809), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n810), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n811), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n812), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n813), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n814), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n815), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n816), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n817), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n818), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n819), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n820), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n594), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n593), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n592), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n591), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n590), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n589), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n588), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n587), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n586), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n585), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n584), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n583), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n582), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n581), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n580), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n579), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n578), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n577), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n576), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n575), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n574), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n573), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n572), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n571), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n570), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n569), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n568), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n567), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n566), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n565), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n564), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n563), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n562), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n561), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n560), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n559), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n558), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n557), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n556), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n555), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n554), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n553), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n552), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n551), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n550), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n549), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n548), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n547), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n546), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n545), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n544), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n543), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n542), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n541), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n540), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n539), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n538), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n537), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n536), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n535), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n534), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n533), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n532), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n531), .CK(clk), .Q(\mem[0][0] ) );
  SDFF_X1 \data_out_reg[5]  ( .D(n182), .SI(n167), .SE(N14), .CK(clk), .Q(
        data_out[5]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n122), .SI(n107), .SE(N14), .CK(clk), .Q(
        data_out[3]) );
  NOR2_X1 U3 ( .A1(n845), .A2(addr[5]), .ZN(n311) );
  AND3_X1 U4 ( .A1(n846), .A2(n847), .A3(n311), .ZN(n240) );
  AND3_X1 U5 ( .A1(n311), .A2(n847), .A3(N13), .ZN(n321) );
  AND3_X1 U6 ( .A1(n311), .A2(n846), .A3(N14), .ZN(n394) );
  AND3_X1 U7 ( .A1(N13), .A2(n311), .A3(N14), .ZN(n467) );
  BUF_X1 U8 ( .A(n618), .Z(n615) );
  BUF_X1 U9 ( .A(n618), .Z(n616) );
  BUF_X1 U10 ( .A(n618), .Z(n617) );
  BUF_X1 U11 ( .A(n618), .Z(n613) );
  BUF_X1 U12 ( .A(N10), .Z(n614) );
  BUF_X1 U13 ( .A(N11), .Z(n611) );
  BUF_X1 U14 ( .A(N11), .Z(n612) );
  BUF_X1 U15 ( .A(N10), .Z(n618) );
  NOR3_X1 U16 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n239) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(n619), .ZN(n250) );
  NOR3_X1 U18 ( .A1(N10), .A2(N12), .A3(n620), .ZN(n260) );
  NOR3_X1 U19 ( .A1(n619), .A2(N12), .A3(n620), .ZN(n270) );
  INV_X1 U20 ( .A(n313), .ZN(n844) );
  INV_X1 U21 ( .A(n323), .ZN(n843) );
  INV_X1 U22 ( .A(n332), .ZN(n842) );
  INV_X1 U23 ( .A(n341), .ZN(n841) );
  INV_X1 U24 ( .A(n386), .ZN(n836) );
  INV_X1 U25 ( .A(n396), .ZN(n835) );
  INV_X1 U26 ( .A(n405), .ZN(n834) );
  INV_X1 U27 ( .A(n414), .ZN(n833) );
  INV_X1 U28 ( .A(n459), .ZN(n828) );
  INV_X1 U29 ( .A(n469), .ZN(n827) );
  INV_X1 U30 ( .A(n478), .ZN(n826) );
  INV_X1 U31 ( .A(n487), .ZN(n825) );
  INV_X1 U32 ( .A(n350), .ZN(n840) );
  INV_X1 U33 ( .A(n359), .ZN(n839) );
  INV_X1 U34 ( .A(n368), .ZN(n838) );
  INV_X1 U35 ( .A(n377), .ZN(n837) );
  INV_X1 U36 ( .A(n496), .ZN(n824) );
  INV_X1 U37 ( .A(n505), .ZN(n823) );
  INV_X1 U38 ( .A(n514), .ZN(n822) );
  INV_X1 U39 ( .A(n523), .ZN(n821) );
  INV_X1 U40 ( .A(n423), .ZN(n832) );
  INV_X1 U41 ( .A(n432), .ZN(n831) );
  INV_X1 U42 ( .A(n441), .ZN(n830) );
  INV_X1 U43 ( .A(n450), .ZN(n829) );
  BUF_X1 U44 ( .A(N12), .Z(n608) );
  BUF_X1 U45 ( .A(N12), .Z(n609) );
  INV_X1 U46 ( .A(N13), .ZN(n846) );
  AND3_X1 U47 ( .A1(n619), .A2(n620), .A3(N12), .ZN(n280) );
  AND3_X1 U48 ( .A1(N10), .A2(n620), .A3(N12), .ZN(n290) );
  AND3_X1 U49 ( .A1(N11), .A2(n619), .A3(N12), .ZN(n300) );
  AND3_X1 U50 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n310) );
  INV_X1 U51 ( .A(N14), .ZN(n847) );
  NAND2_X1 U52 ( .A1(n250), .A2(n240), .ZN(n241) );
  NAND2_X1 U53 ( .A1(n260), .A2(n240), .ZN(n251) );
  NAND2_X1 U54 ( .A1(n270), .A2(n240), .ZN(n261) );
  NAND2_X1 U55 ( .A1(n280), .A2(n240), .ZN(n271) );
  NAND2_X1 U56 ( .A1(n290), .A2(n240), .ZN(n281) );
  NAND2_X1 U57 ( .A1(n300), .A2(n240), .ZN(n291) );
  NAND2_X1 U58 ( .A1(n310), .A2(n240), .ZN(n301) );
  NAND2_X1 U59 ( .A1(n239), .A2(n240), .ZN(n230) );
  NAND2_X1 U60 ( .A1(n321), .A2(n239), .ZN(n313) );
  NAND2_X1 U61 ( .A1(n321), .A2(n250), .ZN(n323) );
  NAND2_X1 U62 ( .A1(n321), .A2(n260), .ZN(n332) );
  NAND2_X1 U63 ( .A1(n321), .A2(n270), .ZN(n341) );
  NAND2_X1 U64 ( .A1(n394), .A2(n239), .ZN(n386) );
  NAND2_X1 U65 ( .A1(n394), .A2(n250), .ZN(n396) );
  NAND2_X1 U66 ( .A1(n394), .A2(n260), .ZN(n405) );
  NAND2_X1 U67 ( .A1(n394), .A2(n270), .ZN(n414) );
  NAND2_X1 U68 ( .A1(n467), .A2(n239), .ZN(n459) );
  NAND2_X1 U69 ( .A1(n467), .A2(n250), .ZN(n469) );
  NAND2_X1 U70 ( .A1(n467), .A2(n260), .ZN(n478) );
  NAND2_X1 U71 ( .A1(n467), .A2(n270), .ZN(n487) );
  NAND2_X1 U72 ( .A1(n321), .A2(n280), .ZN(n350) );
  NAND2_X1 U73 ( .A1(n321), .A2(n290), .ZN(n359) );
  NAND2_X1 U74 ( .A1(n321), .A2(n300), .ZN(n368) );
  NAND2_X1 U75 ( .A1(n321), .A2(n310), .ZN(n377) );
  NAND2_X1 U76 ( .A1(n394), .A2(n280), .ZN(n423) );
  NAND2_X1 U77 ( .A1(n394), .A2(n290), .ZN(n432) );
  NAND2_X1 U78 ( .A1(n394), .A2(n300), .ZN(n441) );
  NAND2_X1 U79 ( .A1(n394), .A2(n310), .ZN(n450) );
  NAND2_X1 U80 ( .A1(n467), .A2(n280), .ZN(n496) );
  NAND2_X1 U81 ( .A1(n467), .A2(n290), .ZN(n505) );
  NAND2_X1 U82 ( .A1(n467), .A2(n300), .ZN(n514) );
  NAND2_X1 U83 ( .A1(n467), .A2(n310), .ZN(n523) );
  INV_X1 U84 ( .A(wr_en), .ZN(n845) );
  OAI21_X1 U85 ( .B1(n621), .B2(n271), .A(n272), .ZN(n563) );
  NAND2_X1 U86 ( .A1(\mem[4][0] ), .A2(n271), .ZN(n272) );
  OAI21_X1 U87 ( .B1(n622), .B2(n271), .A(n273), .ZN(n564) );
  NAND2_X1 U88 ( .A1(\mem[4][1] ), .A2(n271), .ZN(n273) );
  OAI21_X1 U89 ( .B1(n623), .B2(n271), .A(n274), .ZN(n565) );
  NAND2_X1 U90 ( .A1(\mem[4][2] ), .A2(n271), .ZN(n274) );
  OAI21_X1 U91 ( .B1(n624), .B2(n271), .A(n275), .ZN(n566) );
  NAND2_X1 U92 ( .A1(\mem[4][3] ), .A2(n271), .ZN(n275) );
  OAI21_X1 U93 ( .B1(n625), .B2(n271), .A(n276), .ZN(n567) );
  NAND2_X1 U94 ( .A1(\mem[4][4] ), .A2(n271), .ZN(n276) );
  OAI21_X1 U95 ( .B1(n626), .B2(n271), .A(n277), .ZN(n568) );
  NAND2_X1 U96 ( .A1(\mem[4][5] ), .A2(n271), .ZN(n277) );
  OAI21_X1 U97 ( .B1(n627), .B2(n271), .A(n278), .ZN(n569) );
  NAND2_X1 U98 ( .A1(\mem[4][6] ), .A2(n271), .ZN(n278) );
  OAI21_X1 U99 ( .B1(n628), .B2(n271), .A(n279), .ZN(n570) );
  NAND2_X1 U100 ( .A1(\mem[4][7] ), .A2(n271), .ZN(n279) );
  OAI21_X1 U101 ( .B1(n621), .B2(n291), .A(n292), .ZN(n579) );
  NAND2_X1 U102 ( .A1(\mem[6][0] ), .A2(n291), .ZN(n292) );
  OAI21_X1 U103 ( .B1(n622), .B2(n291), .A(n293), .ZN(n580) );
  NAND2_X1 U104 ( .A1(\mem[6][1] ), .A2(n291), .ZN(n293) );
  OAI21_X1 U105 ( .B1(n623), .B2(n291), .A(n294), .ZN(n581) );
  NAND2_X1 U106 ( .A1(\mem[6][2] ), .A2(n291), .ZN(n294) );
  OAI21_X1 U107 ( .B1(n624), .B2(n291), .A(n295), .ZN(n582) );
  NAND2_X1 U108 ( .A1(\mem[6][3] ), .A2(n291), .ZN(n295) );
  OAI21_X1 U109 ( .B1(n625), .B2(n291), .A(n296), .ZN(n583) );
  NAND2_X1 U110 ( .A1(\mem[6][4] ), .A2(n291), .ZN(n296) );
  OAI21_X1 U111 ( .B1(n626), .B2(n291), .A(n297), .ZN(n584) );
  NAND2_X1 U112 ( .A1(\mem[6][5] ), .A2(n291), .ZN(n297) );
  OAI21_X1 U113 ( .B1(n627), .B2(n291), .A(n298), .ZN(n585) );
  NAND2_X1 U114 ( .A1(\mem[6][6] ), .A2(n291), .ZN(n298) );
  OAI21_X1 U115 ( .B1(n628), .B2(n291), .A(n299), .ZN(n586) );
  NAND2_X1 U116 ( .A1(\mem[6][7] ), .A2(n291), .ZN(n299) );
  OAI21_X1 U117 ( .B1(n621), .B2(n301), .A(n302), .ZN(n587) );
  NAND2_X1 U118 ( .A1(\mem[7][0] ), .A2(n301), .ZN(n302) );
  OAI21_X1 U119 ( .B1(n622), .B2(n301), .A(n303), .ZN(n588) );
  NAND2_X1 U120 ( .A1(\mem[7][1] ), .A2(n301), .ZN(n303) );
  OAI21_X1 U121 ( .B1(n623), .B2(n301), .A(n304), .ZN(n589) );
  NAND2_X1 U122 ( .A1(\mem[7][2] ), .A2(n301), .ZN(n304) );
  OAI21_X1 U123 ( .B1(n624), .B2(n301), .A(n305), .ZN(n590) );
  NAND2_X1 U124 ( .A1(\mem[7][3] ), .A2(n301), .ZN(n305) );
  OAI21_X1 U125 ( .B1(n625), .B2(n301), .A(n306), .ZN(n591) );
  NAND2_X1 U126 ( .A1(\mem[7][4] ), .A2(n301), .ZN(n306) );
  OAI21_X1 U127 ( .B1(n626), .B2(n301), .A(n307), .ZN(n592) );
  NAND2_X1 U128 ( .A1(\mem[7][5] ), .A2(n301), .ZN(n307) );
  OAI21_X1 U129 ( .B1(n627), .B2(n301), .A(n308), .ZN(n593) );
  NAND2_X1 U130 ( .A1(\mem[7][6] ), .A2(n301), .ZN(n308) );
  OAI21_X1 U131 ( .B1(n628), .B2(n301), .A(n309), .ZN(n594) );
  NAND2_X1 U132 ( .A1(\mem[7][7] ), .A2(n301), .ZN(n309) );
  OAI21_X1 U133 ( .B1(n621), .B2(n241), .A(n242), .ZN(n539) );
  NAND2_X1 U134 ( .A1(\mem[1][0] ), .A2(n241), .ZN(n242) );
  OAI21_X1 U135 ( .B1(n622), .B2(n241), .A(n243), .ZN(n540) );
  NAND2_X1 U136 ( .A1(\mem[1][1] ), .A2(n241), .ZN(n243) );
  OAI21_X1 U137 ( .B1(n623), .B2(n241), .A(n244), .ZN(n541) );
  NAND2_X1 U138 ( .A1(\mem[1][2] ), .A2(n241), .ZN(n244) );
  OAI21_X1 U139 ( .B1(n624), .B2(n241), .A(n245), .ZN(n542) );
  NAND2_X1 U140 ( .A1(\mem[1][3] ), .A2(n241), .ZN(n245) );
  OAI21_X1 U141 ( .B1(n625), .B2(n241), .A(n246), .ZN(n543) );
  NAND2_X1 U142 ( .A1(\mem[1][4] ), .A2(n241), .ZN(n246) );
  OAI21_X1 U143 ( .B1(n626), .B2(n241), .A(n247), .ZN(n544) );
  NAND2_X1 U144 ( .A1(\mem[1][5] ), .A2(n241), .ZN(n247) );
  OAI21_X1 U145 ( .B1(n627), .B2(n241), .A(n248), .ZN(n545) );
  NAND2_X1 U146 ( .A1(\mem[1][6] ), .A2(n241), .ZN(n248) );
  OAI21_X1 U147 ( .B1(n628), .B2(n241), .A(n249), .ZN(n546) );
  NAND2_X1 U148 ( .A1(\mem[1][7] ), .A2(n241), .ZN(n249) );
  OAI21_X1 U149 ( .B1(n621), .B2(n251), .A(n252), .ZN(n547) );
  NAND2_X1 U150 ( .A1(\mem[2][0] ), .A2(n251), .ZN(n252) );
  OAI21_X1 U151 ( .B1(n622), .B2(n251), .A(n253), .ZN(n548) );
  NAND2_X1 U152 ( .A1(\mem[2][1] ), .A2(n251), .ZN(n253) );
  OAI21_X1 U153 ( .B1(n623), .B2(n251), .A(n254), .ZN(n549) );
  NAND2_X1 U154 ( .A1(\mem[2][2] ), .A2(n251), .ZN(n254) );
  OAI21_X1 U155 ( .B1(n624), .B2(n251), .A(n255), .ZN(n550) );
  NAND2_X1 U156 ( .A1(\mem[2][3] ), .A2(n251), .ZN(n255) );
  OAI21_X1 U157 ( .B1(n625), .B2(n251), .A(n256), .ZN(n551) );
  NAND2_X1 U158 ( .A1(\mem[2][4] ), .A2(n251), .ZN(n256) );
  OAI21_X1 U159 ( .B1(n626), .B2(n251), .A(n257), .ZN(n552) );
  NAND2_X1 U160 ( .A1(\mem[2][5] ), .A2(n251), .ZN(n257) );
  OAI21_X1 U161 ( .B1(n627), .B2(n251), .A(n258), .ZN(n553) );
  NAND2_X1 U162 ( .A1(\mem[2][6] ), .A2(n251), .ZN(n258) );
  OAI21_X1 U163 ( .B1(n628), .B2(n251), .A(n259), .ZN(n554) );
  NAND2_X1 U164 ( .A1(\mem[2][7] ), .A2(n251), .ZN(n259) );
  OAI21_X1 U165 ( .B1(n621), .B2(n261), .A(n262), .ZN(n555) );
  NAND2_X1 U166 ( .A1(\mem[3][0] ), .A2(n261), .ZN(n262) );
  OAI21_X1 U167 ( .B1(n622), .B2(n261), .A(n263), .ZN(n556) );
  NAND2_X1 U168 ( .A1(\mem[3][1] ), .A2(n261), .ZN(n263) );
  OAI21_X1 U169 ( .B1(n623), .B2(n261), .A(n264), .ZN(n557) );
  NAND2_X1 U170 ( .A1(\mem[3][2] ), .A2(n261), .ZN(n264) );
  OAI21_X1 U171 ( .B1(n624), .B2(n261), .A(n265), .ZN(n558) );
  NAND2_X1 U172 ( .A1(\mem[3][3] ), .A2(n261), .ZN(n265) );
  OAI21_X1 U173 ( .B1(n625), .B2(n261), .A(n266), .ZN(n559) );
  NAND2_X1 U174 ( .A1(\mem[3][4] ), .A2(n261), .ZN(n266) );
  OAI21_X1 U175 ( .B1(n626), .B2(n261), .A(n267), .ZN(n560) );
  NAND2_X1 U176 ( .A1(\mem[3][5] ), .A2(n261), .ZN(n267) );
  OAI21_X1 U177 ( .B1(n627), .B2(n261), .A(n268), .ZN(n561) );
  NAND2_X1 U178 ( .A1(\mem[3][6] ), .A2(n261), .ZN(n268) );
  OAI21_X1 U179 ( .B1(n628), .B2(n261), .A(n269), .ZN(n562) );
  NAND2_X1 U180 ( .A1(\mem[3][7] ), .A2(n261), .ZN(n269) );
  OAI21_X1 U181 ( .B1(n621), .B2(n281), .A(n282), .ZN(n571) );
  NAND2_X1 U182 ( .A1(\mem[5][0] ), .A2(n281), .ZN(n282) );
  OAI21_X1 U183 ( .B1(n622), .B2(n281), .A(n283), .ZN(n572) );
  NAND2_X1 U184 ( .A1(\mem[5][1] ), .A2(n281), .ZN(n283) );
  OAI21_X1 U185 ( .B1(n623), .B2(n281), .A(n284), .ZN(n573) );
  NAND2_X1 U186 ( .A1(\mem[5][2] ), .A2(n281), .ZN(n284) );
  OAI21_X1 U187 ( .B1(n624), .B2(n281), .A(n285), .ZN(n574) );
  NAND2_X1 U188 ( .A1(\mem[5][3] ), .A2(n281), .ZN(n285) );
  OAI21_X1 U189 ( .B1(n625), .B2(n281), .A(n286), .ZN(n575) );
  NAND2_X1 U190 ( .A1(\mem[5][4] ), .A2(n281), .ZN(n286) );
  OAI21_X1 U191 ( .B1(n626), .B2(n281), .A(n287), .ZN(n576) );
  NAND2_X1 U192 ( .A1(\mem[5][5] ), .A2(n281), .ZN(n287) );
  OAI21_X1 U193 ( .B1(n627), .B2(n281), .A(n288), .ZN(n577) );
  NAND2_X1 U194 ( .A1(\mem[5][6] ), .A2(n281), .ZN(n288) );
  OAI21_X1 U195 ( .B1(n628), .B2(n281), .A(n289), .ZN(n578) );
  NAND2_X1 U196 ( .A1(\mem[5][7] ), .A2(n281), .ZN(n289) );
  OAI21_X1 U197 ( .B1(n230), .B2(n621), .A(n231), .ZN(n531) );
  NAND2_X1 U198 ( .A1(\mem[0][0] ), .A2(n230), .ZN(n231) );
  OAI21_X1 U199 ( .B1(n230), .B2(n622), .A(n232), .ZN(n532) );
  NAND2_X1 U200 ( .A1(\mem[0][1] ), .A2(n230), .ZN(n232) );
  OAI21_X1 U201 ( .B1(n230), .B2(n623), .A(n233), .ZN(n533) );
  NAND2_X1 U202 ( .A1(\mem[0][2] ), .A2(n230), .ZN(n233) );
  OAI21_X1 U203 ( .B1(n230), .B2(n624), .A(n234), .ZN(n534) );
  NAND2_X1 U204 ( .A1(\mem[0][3] ), .A2(n230), .ZN(n234) );
  OAI21_X1 U205 ( .B1(n230), .B2(n625), .A(n235), .ZN(n535) );
  NAND2_X1 U206 ( .A1(\mem[0][4] ), .A2(n230), .ZN(n235) );
  OAI21_X1 U207 ( .B1(n230), .B2(n626), .A(n236), .ZN(n536) );
  NAND2_X1 U208 ( .A1(\mem[0][5] ), .A2(n230), .ZN(n236) );
  OAI21_X1 U209 ( .B1(n230), .B2(n627), .A(n237), .ZN(n537) );
  NAND2_X1 U210 ( .A1(\mem[0][6] ), .A2(n230), .ZN(n237) );
  OAI21_X1 U211 ( .B1(n230), .B2(n628), .A(n238), .ZN(n538) );
  NAND2_X1 U212 ( .A1(\mem[0][7] ), .A2(n230), .ZN(n238) );
  INV_X1 U213 ( .A(n312), .ZN(n820) );
  AOI22_X1 U214 ( .A1(data_in[0]), .A2(n844), .B1(n313), .B2(\mem[8][0] ), 
        .ZN(n312) );
  INV_X1 U215 ( .A(n314), .ZN(n819) );
  AOI22_X1 U216 ( .A1(data_in[1]), .A2(n844), .B1(n313), .B2(\mem[8][1] ), 
        .ZN(n314) );
  INV_X1 U217 ( .A(n315), .ZN(n818) );
  AOI22_X1 U218 ( .A1(data_in[2]), .A2(n844), .B1(n313), .B2(\mem[8][2] ), 
        .ZN(n315) );
  INV_X1 U219 ( .A(n316), .ZN(n817) );
  AOI22_X1 U220 ( .A1(data_in[3]), .A2(n844), .B1(n313), .B2(\mem[8][3] ), 
        .ZN(n316) );
  INV_X1 U221 ( .A(n317), .ZN(n816) );
  AOI22_X1 U222 ( .A1(data_in[4]), .A2(n844), .B1(n313), .B2(\mem[8][4] ), 
        .ZN(n317) );
  INV_X1 U223 ( .A(n318), .ZN(n815) );
  AOI22_X1 U224 ( .A1(data_in[5]), .A2(n844), .B1(n313), .B2(\mem[8][5] ), 
        .ZN(n318) );
  INV_X1 U225 ( .A(n319), .ZN(n814) );
  AOI22_X1 U226 ( .A1(data_in[6]), .A2(n844), .B1(n313), .B2(\mem[8][6] ), 
        .ZN(n319) );
  INV_X1 U227 ( .A(n320), .ZN(n813) );
  AOI22_X1 U228 ( .A1(data_in[7]), .A2(n844), .B1(n313), .B2(\mem[8][7] ), 
        .ZN(n320) );
  INV_X1 U229 ( .A(n322), .ZN(n812) );
  AOI22_X1 U230 ( .A1(data_in[0]), .A2(n843), .B1(n323), .B2(\mem[9][0] ), 
        .ZN(n322) );
  INV_X1 U231 ( .A(n324), .ZN(n811) );
  AOI22_X1 U232 ( .A1(data_in[1]), .A2(n843), .B1(n323), .B2(\mem[9][1] ), 
        .ZN(n324) );
  INV_X1 U233 ( .A(n325), .ZN(n810) );
  AOI22_X1 U234 ( .A1(data_in[2]), .A2(n843), .B1(n323), .B2(\mem[9][2] ), 
        .ZN(n325) );
  INV_X1 U235 ( .A(n326), .ZN(n809) );
  AOI22_X1 U236 ( .A1(data_in[3]), .A2(n843), .B1(n323), .B2(\mem[9][3] ), 
        .ZN(n326) );
  INV_X1 U237 ( .A(n327), .ZN(n808) );
  AOI22_X1 U238 ( .A1(data_in[4]), .A2(n843), .B1(n323), .B2(\mem[9][4] ), 
        .ZN(n327) );
  INV_X1 U239 ( .A(n328), .ZN(n807) );
  AOI22_X1 U240 ( .A1(data_in[5]), .A2(n843), .B1(n323), .B2(\mem[9][5] ), 
        .ZN(n328) );
  INV_X1 U241 ( .A(n329), .ZN(n806) );
  AOI22_X1 U242 ( .A1(data_in[6]), .A2(n843), .B1(n323), .B2(\mem[9][6] ), 
        .ZN(n329) );
  INV_X1 U243 ( .A(n330), .ZN(n805) );
  AOI22_X1 U244 ( .A1(data_in[7]), .A2(n843), .B1(n323), .B2(\mem[9][7] ), 
        .ZN(n330) );
  INV_X1 U245 ( .A(n331), .ZN(n804) );
  AOI22_X1 U246 ( .A1(data_in[0]), .A2(n842), .B1(n332), .B2(\mem[10][0] ), 
        .ZN(n331) );
  INV_X1 U247 ( .A(n333), .ZN(n803) );
  AOI22_X1 U248 ( .A1(data_in[1]), .A2(n842), .B1(n332), .B2(\mem[10][1] ), 
        .ZN(n333) );
  INV_X1 U249 ( .A(n334), .ZN(n802) );
  AOI22_X1 U250 ( .A1(data_in[2]), .A2(n842), .B1(n332), .B2(\mem[10][2] ), 
        .ZN(n334) );
  INV_X1 U251 ( .A(n335), .ZN(n801) );
  AOI22_X1 U252 ( .A1(data_in[3]), .A2(n842), .B1(n332), .B2(\mem[10][3] ), 
        .ZN(n335) );
  INV_X1 U253 ( .A(n336), .ZN(n800) );
  AOI22_X1 U254 ( .A1(data_in[4]), .A2(n842), .B1(n332), .B2(\mem[10][4] ), 
        .ZN(n336) );
  INV_X1 U255 ( .A(n337), .ZN(n799) );
  AOI22_X1 U256 ( .A1(data_in[5]), .A2(n842), .B1(n332), .B2(\mem[10][5] ), 
        .ZN(n337) );
  INV_X1 U257 ( .A(n338), .ZN(n798) );
  AOI22_X1 U258 ( .A1(data_in[6]), .A2(n842), .B1(n332), .B2(\mem[10][6] ), 
        .ZN(n338) );
  INV_X1 U259 ( .A(n339), .ZN(n797) );
  AOI22_X1 U260 ( .A1(data_in[7]), .A2(n842), .B1(n332), .B2(\mem[10][7] ), 
        .ZN(n339) );
  INV_X1 U261 ( .A(n340), .ZN(n796) );
  AOI22_X1 U262 ( .A1(data_in[0]), .A2(n841), .B1(n341), .B2(\mem[11][0] ), 
        .ZN(n340) );
  INV_X1 U263 ( .A(n342), .ZN(n795) );
  AOI22_X1 U264 ( .A1(data_in[1]), .A2(n841), .B1(n341), .B2(\mem[11][1] ), 
        .ZN(n342) );
  INV_X1 U265 ( .A(n343), .ZN(n794) );
  AOI22_X1 U266 ( .A1(data_in[2]), .A2(n841), .B1(n341), .B2(\mem[11][2] ), 
        .ZN(n343) );
  INV_X1 U267 ( .A(n344), .ZN(n793) );
  AOI22_X1 U268 ( .A1(data_in[3]), .A2(n841), .B1(n341), .B2(\mem[11][3] ), 
        .ZN(n344) );
  INV_X1 U269 ( .A(n345), .ZN(n792) );
  AOI22_X1 U270 ( .A1(data_in[4]), .A2(n841), .B1(n341), .B2(\mem[11][4] ), 
        .ZN(n345) );
  INV_X1 U271 ( .A(n346), .ZN(n791) );
  AOI22_X1 U272 ( .A1(data_in[5]), .A2(n841), .B1(n341), .B2(\mem[11][5] ), 
        .ZN(n346) );
  INV_X1 U273 ( .A(n347), .ZN(n790) );
  AOI22_X1 U274 ( .A1(data_in[6]), .A2(n841), .B1(n341), .B2(\mem[11][6] ), 
        .ZN(n347) );
  INV_X1 U275 ( .A(n348), .ZN(n789) );
  AOI22_X1 U276 ( .A1(data_in[7]), .A2(n841), .B1(n341), .B2(\mem[11][7] ), 
        .ZN(n348) );
  INV_X1 U277 ( .A(n349), .ZN(n788) );
  AOI22_X1 U278 ( .A1(data_in[0]), .A2(n840), .B1(n350), .B2(\mem[12][0] ), 
        .ZN(n349) );
  INV_X1 U279 ( .A(n351), .ZN(n787) );
  AOI22_X1 U280 ( .A1(data_in[1]), .A2(n840), .B1(n350), .B2(\mem[12][1] ), 
        .ZN(n351) );
  INV_X1 U281 ( .A(n352), .ZN(n786) );
  AOI22_X1 U282 ( .A1(data_in[2]), .A2(n840), .B1(n350), .B2(\mem[12][2] ), 
        .ZN(n352) );
  INV_X1 U283 ( .A(n353), .ZN(n785) );
  AOI22_X1 U284 ( .A1(data_in[3]), .A2(n840), .B1(n350), .B2(\mem[12][3] ), 
        .ZN(n353) );
  INV_X1 U285 ( .A(n354), .ZN(n784) );
  AOI22_X1 U286 ( .A1(data_in[4]), .A2(n840), .B1(n350), .B2(\mem[12][4] ), 
        .ZN(n354) );
  INV_X1 U287 ( .A(n355), .ZN(n783) );
  AOI22_X1 U288 ( .A1(data_in[5]), .A2(n840), .B1(n350), .B2(\mem[12][5] ), 
        .ZN(n355) );
  INV_X1 U289 ( .A(n356), .ZN(n782) );
  AOI22_X1 U290 ( .A1(data_in[6]), .A2(n840), .B1(n350), .B2(\mem[12][6] ), 
        .ZN(n356) );
  INV_X1 U291 ( .A(n357), .ZN(n781) );
  AOI22_X1 U292 ( .A1(data_in[7]), .A2(n840), .B1(n350), .B2(\mem[12][7] ), 
        .ZN(n357) );
  INV_X1 U293 ( .A(n358), .ZN(n780) );
  AOI22_X1 U294 ( .A1(data_in[0]), .A2(n839), .B1(n359), .B2(\mem[13][0] ), 
        .ZN(n358) );
  INV_X1 U295 ( .A(n360), .ZN(n779) );
  AOI22_X1 U296 ( .A1(data_in[1]), .A2(n839), .B1(n359), .B2(\mem[13][1] ), 
        .ZN(n360) );
  INV_X1 U297 ( .A(n361), .ZN(n778) );
  AOI22_X1 U298 ( .A1(data_in[2]), .A2(n839), .B1(n359), .B2(\mem[13][2] ), 
        .ZN(n361) );
  INV_X1 U299 ( .A(n362), .ZN(n777) );
  AOI22_X1 U300 ( .A1(data_in[3]), .A2(n839), .B1(n359), .B2(\mem[13][3] ), 
        .ZN(n362) );
  INV_X1 U301 ( .A(n363), .ZN(n776) );
  AOI22_X1 U302 ( .A1(data_in[4]), .A2(n839), .B1(n359), .B2(\mem[13][4] ), 
        .ZN(n363) );
  INV_X1 U303 ( .A(n364), .ZN(n775) );
  AOI22_X1 U304 ( .A1(data_in[5]), .A2(n839), .B1(n359), .B2(\mem[13][5] ), 
        .ZN(n364) );
  INV_X1 U305 ( .A(n365), .ZN(n774) );
  AOI22_X1 U306 ( .A1(data_in[6]), .A2(n839), .B1(n359), .B2(\mem[13][6] ), 
        .ZN(n365) );
  INV_X1 U307 ( .A(n366), .ZN(n773) );
  AOI22_X1 U308 ( .A1(data_in[7]), .A2(n839), .B1(n359), .B2(\mem[13][7] ), 
        .ZN(n366) );
  INV_X1 U309 ( .A(n367), .ZN(n772) );
  AOI22_X1 U310 ( .A1(data_in[0]), .A2(n838), .B1(n368), .B2(\mem[14][0] ), 
        .ZN(n367) );
  INV_X1 U311 ( .A(n369), .ZN(n771) );
  AOI22_X1 U312 ( .A1(data_in[1]), .A2(n838), .B1(n368), .B2(\mem[14][1] ), 
        .ZN(n369) );
  INV_X1 U313 ( .A(n370), .ZN(n770) );
  AOI22_X1 U314 ( .A1(data_in[2]), .A2(n838), .B1(n368), .B2(\mem[14][2] ), 
        .ZN(n370) );
  INV_X1 U315 ( .A(n371), .ZN(n769) );
  AOI22_X1 U316 ( .A1(data_in[3]), .A2(n838), .B1(n368), .B2(\mem[14][3] ), 
        .ZN(n371) );
  INV_X1 U317 ( .A(n372), .ZN(n768) );
  AOI22_X1 U318 ( .A1(data_in[4]), .A2(n838), .B1(n368), .B2(\mem[14][4] ), 
        .ZN(n372) );
  INV_X1 U319 ( .A(n373), .ZN(n767) );
  AOI22_X1 U320 ( .A1(data_in[5]), .A2(n838), .B1(n368), .B2(\mem[14][5] ), 
        .ZN(n373) );
  INV_X1 U321 ( .A(n374), .ZN(n766) );
  AOI22_X1 U322 ( .A1(data_in[6]), .A2(n838), .B1(n368), .B2(\mem[14][6] ), 
        .ZN(n374) );
  INV_X1 U323 ( .A(n375), .ZN(n765) );
  AOI22_X1 U324 ( .A1(data_in[7]), .A2(n838), .B1(n368), .B2(\mem[14][7] ), 
        .ZN(n375) );
  INV_X1 U325 ( .A(n376), .ZN(n764) );
  AOI22_X1 U326 ( .A1(data_in[0]), .A2(n837), .B1(n377), .B2(\mem[15][0] ), 
        .ZN(n376) );
  INV_X1 U327 ( .A(n378), .ZN(n763) );
  AOI22_X1 U328 ( .A1(data_in[1]), .A2(n837), .B1(n377), .B2(\mem[15][1] ), 
        .ZN(n378) );
  INV_X1 U329 ( .A(n379), .ZN(n762) );
  AOI22_X1 U330 ( .A1(data_in[2]), .A2(n837), .B1(n377), .B2(\mem[15][2] ), 
        .ZN(n379) );
  INV_X1 U331 ( .A(n380), .ZN(n761) );
  AOI22_X1 U332 ( .A1(data_in[3]), .A2(n837), .B1(n377), .B2(\mem[15][3] ), 
        .ZN(n380) );
  INV_X1 U333 ( .A(n381), .ZN(n760) );
  AOI22_X1 U334 ( .A1(data_in[4]), .A2(n837), .B1(n377), .B2(\mem[15][4] ), 
        .ZN(n381) );
  INV_X1 U335 ( .A(n382), .ZN(n759) );
  AOI22_X1 U336 ( .A1(data_in[5]), .A2(n837), .B1(n377), .B2(\mem[15][5] ), 
        .ZN(n382) );
  INV_X1 U337 ( .A(n383), .ZN(n758) );
  AOI22_X1 U338 ( .A1(data_in[6]), .A2(n837), .B1(n377), .B2(\mem[15][6] ), 
        .ZN(n383) );
  INV_X1 U339 ( .A(n384), .ZN(n757) );
  AOI22_X1 U340 ( .A1(data_in[7]), .A2(n837), .B1(n377), .B2(\mem[15][7] ), 
        .ZN(n384) );
  INV_X1 U341 ( .A(n385), .ZN(n756) );
  AOI22_X1 U342 ( .A1(data_in[0]), .A2(n836), .B1(n386), .B2(\mem[16][0] ), 
        .ZN(n385) );
  INV_X1 U343 ( .A(n387), .ZN(n755) );
  AOI22_X1 U344 ( .A1(data_in[1]), .A2(n836), .B1(n386), .B2(\mem[16][1] ), 
        .ZN(n387) );
  INV_X1 U345 ( .A(n388), .ZN(n754) );
  AOI22_X1 U346 ( .A1(data_in[2]), .A2(n836), .B1(n386), .B2(\mem[16][2] ), 
        .ZN(n388) );
  INV_X1 U347 ( .A(n389), .ZN(n753) );
  AOI22_X1 U348 ( .A1(data_in[3]), .A2(n836), .B1(n386), .B2(\mem[16][3] ), 
        .ZN(n389) );
  INV_X1 U349 ( .A(n390), .ZN(n752) );
  AOI22_X1 U350 ( .A1(data_in[4]), .A2(n836), .B1(n386), .B2(\mem[16][4] ), 
        .ZN(n390) );
  INV_X1 U351 ( .A(n391), .ZN(n751) );
  AOI22_X1 U352 ( .A1(data_in[5]), .A2(n836), .B1(n386), .B2(\mem[16][5] ), 
        .ZN(n391) );
  INV_X1 U353 ( .A(n392), .ZN(n750) );
  AOI22_X1 U354 ( .A1(data_in[6]), .A2(n836), .B1(n386), .B2(\mem[16][6] ), 
        .ZN(n392) );
  INV_X1 U355 ( .A(n393), .ZN(n749) );
  AOI22_X1 U356 ( .A1(data_in[7]), .A2(n836), .B1(n386), .B2(\mem[16][7] ), 
        .ZN(n393) );
  INV_X1 U357 ( .A(n395), .ZN(n748) );
  AOI22_X1 U358 ( .A1(data_in[0]), .A2(n835), .B1(n396), .B2(\mem[17][0] ), 
        .ZN(n395) );
  INV_X1 U359 ( .A(n397), .ZN(n747) );
  AOI22_X1 U360 ( .A1(data_in[1]), .A2(n835), .B1(n396), .B2(\mem[17][1] ), 
        .ZN(n397) );
  INV_X1 U361 ( .A(n398), .ZN(n746) );
  AOI22_X1 U362 ( .A1(data_in[2]), .A2(n835), .B1(n396), .B2(\mem[17][2] ), 
        .ZN(n398) );
  INV_X1 U363 ( .A(n399), .ZN(n745) );
  AOI22_X1 U364 ( .A1(data_in[3]), .A2(n835), .B1(n396), .B2(\mem[17][3] ), 
        .ZN(n399) );
  INV_X1 U365 ( .A(n400), .ZN(n744) );
  AOI22_X1 U366 ( .A1(data_in[4]), .A2(n835), .B1(n396), .B2(\mem[17][4] ), 
        .ZN(n400) );
  INV_X1 U367 ( .A(n401), .ZN(n743) );
  AOI22_X1 U368 ( .A1(data_in[5]), .A2(n835), .B1(n396), .B2(\mem[17][5] ), 
        .ZN(n401) );
  INV_X1 U369 ( .A(n402), .ZN(n742) );
  AOI22_X1 U370 ( .A1(data_in[6]), .A2(n835), .B1(n396), .B2(\mem[17][6] ), 
        .ZN(n402) );
  INV_X1 U371 ( .A(n403), .ZN(n741) );
  AOI22_X1 U372 ( .A1(data_in[7]), .A2(n835), .B1(n396), .B2(\mem[17][7] ), 
        .ZN(n403) );
  INV_X1 U373 ( .A(n404), .ZN(n740) );
  AOI22_X1 U374 ( .A1(data_in[0]), .A2(n834), .B1(n405), .B2(\mem[18][0] ), 
        .ZN(n404) );
  INV_X1 U375 ( .A(n406), .ZN(n739) );
  AOI22_X1 U376 ( .A1(data_in[1]), .A2(n834), .B1(n405), .B2(\mem[18][1] ), 
        .ZN(n406) );
  INV_X1 U377 ( .A(n407), .ZN(n738) );
  AOI22_X1 U378 ( .A1(data_in[2]), .A2(n834), .B1(n405), .B2(\mem[18][2] ), 
        .ZN(n407) );
  INV_X1 U379 ( .A(n408), .ZN(n737) );
  AOI22_X1 U380 ( .A1(data_in[3]), .A2(n834), .B1(n405), .B2(\mem[18][3] ), 
        .ZN(n408) );
  INV_X1 U381 ( .A(n409), .ZN(n736) );
  AOI22_X1 U382 ( .A1(data_in[4]), .A2(n834), .B1(n405), .B2(\mem[18][4] ), 
        .ZN(n409) );
  INV_X1 U383 ( .A(n410), .ZN(n735) );
  AOI22_X1 U384 ( .A1(data_in[5]), .A2(n834), .B1(n405), .B2(\mem[18][5] ), 
        .ZN(n410) );
  INV_X1 U385 ( .A(n411), .ZN(n734) );
  AOI22_X1 U386 ( .A1(data_in[6]), .A2(n834), .B1(n405), .B2(\mem[18][6] ), 
        .ZN(n411) );
  INV_X1 U387 ( .A(n412), .ZN(n733) );
  AOI22_X1 U388 ( .A1(data_in[7]), .A2(n834), .B1(n405), .B2(\mem[18][7] ), 
        .ZN(n412) );
  INV_X1 U389 ( .A(n413), .ZN(n732) );
  AOI22_X1 U390 ( .A1(data_in[0]), .A2(n833), .B1(n414), .B2(\mem[19][0] ), 
        .ZN(n413) );
  INV_X1 U391 ( .A(n415), .ZN(n731) );
  AOI22_X1 U392 ( .A1(data_in[1]), .A2(n833), .B1(n414), .B2(\mem[19][1] ), 
        .ZN(n415) );
  INV_X1 U393 ( .A(n416), .ZN(n730) );
  AOI22_X1 U394 ( .A1(data_in[2]), .A2(n833), .B1(n414), .B2(\mem[19][2] ), 
        .ZN(n416) );
  INV_X1 U395 ( .A(n417), .ZN(n729) );
  AOI22_X1 U396 ( .A1(data_in[3]), .A2(n833), .B1(n414), .B2(\mem[19][3] ), 
        .ZN(n417) );
  INV_X1 U397 ( .A(n418), .ZN(n728) );
  AOI22_X1 U398 ( .A1(data_in[4]), .A2(n833), .B1(n414), .B2(\mem[19][4] ), 
        .ZN(n418) );
  INV_X1 U399 ( .A(n419), .ZN(n727) );
  AOI22_X1 U400 ( .A1(data_in[5]), .A2(n833), .B1(n414), .B2(\mem[19][5] ), 
        .ZN(n419) );
  INV_X1 U401 ( .A(n420), .ZN(n726) );
  AOI22_X1 U402 ( .A1(data_in[6]), .A2(n833), .B1(n414), .B2(\mem[19][6] ), 
        .ZN(n420) );
  INV_X1 U403 ( .A(n421), .ZN(n725) );
  AOI22_X1 U404 ( .A1(data_in[7]), .A2(n833), .B1(n414), .B2(\mem[19][7] ), 
        .ZN(n421) );
  INV_X1 U405 ( .A(n422), .ZN(n724) );
  AOI22_X1 U406 ( .A1(data_in[0]), .A2(n832), .B1(n423), .B2(\mem[20][0] ), 
        .ZN(n422) );
  INV_X1 U407 ( .A(n424), .ZN(n723) );
  AOI22_X1 U408 ( .A1(data_in[1]), .A2(n832), .B1(n423), .B2(\mem[20][1] ), 
        .ZN(n424) );
  INV_X1 U409 ( .A(n425), .ZN(n722) );
  AOI22_X1 U410 ( .A1(data_in[2]), .A2(n832), .B1(n423), .B2(\mem[20][2] ), 
        .ZN(n425) );
  INV_X1 U411 ( .A(n426), .ZN(n721) );
  AOI22_X1 U412 ( .A1(data_in[3]), .A2(n832), .B1(n423), .B2(\mem[20][3] ), 
        .ZN(n426) );
  INV_X1 U413 ( .A(n427), .ZN(n720) );
  AOI22_X1 U414 ( .A1(data_in[4]), .A2(n832), .B1(n423), .B2(\mem[20][4] ), 
        .ZN(n427) );
  INV_X1 U415 ( .A(n428), .ZN(n719) );
  AOI22_X1 U416 ( .A1(data_in[5]), .A2(n832), .B1(n423), .B2(\mem[20][5] ), 
        .ZN(n428) );
  INV_X1 U417 ( .A(n429), .ZN(n718) );
  AOI22_X1 U418 ( .A1(data_in[6]), .A2(n832), .B1(n423), .B2(\mem[20][6] ), 
        .ZN(n429) );
  INV_X1 U419 ( .A(n430), .ZN(n717) );
  AOI22_X1 U420 ( .A1(data_in[7]), .A2(n832), .B1(n423), .B2(\mem[20][7] ), 
        .ZN(n430) );
  INV_X1 U421 ( .A(n431), .ZN(n716) );
  AOI22_X1 U422 ( .A1(data_in[0]), .A2(n831), .B1(n432), .B2(\mem[21][0] ), 
        .ZN(n431) );
  INV_X1 U423 ( .A(n433), .ZN(n715) );
  AOI22_X1 U424 ( .A1(data_in[1]), .A2(n831), .B1(n432), .B2(\mem[21][1] ), 
        .ZN(n433) );
  INV_X1 U425 ( .A(n434), .ZN(n714) );
  AOI22_X1 U426 ( .A1(data_in[2]), .A2(n831), .B1(n432), .B2(\mem[21][2] ), 
        .ZN(n434) );
  INV_X1 U427 ( .A(n435), .ZN(n713) );
  AOI22_X1 U428 ( .A1(data_in[3]), .A2(n831), .B1(n432), .B2(\mem[21][3] ), 
        .ZN(n435) );
  INV_X1 U429 ( .A(n436), .ZN(n712) );
  AOI22_X1 U430 ( .A1(data_in[4]), .A2(n831), .B1(n432), .B2(\mem[21][4] ), 
        .ZN(n436) );
  INV_X1 U431 ( .A(n437), .ZN(n711) );
  AOI22_X1 U432 ( .A1(data_in[5]), .A2(n831), .B1(n432), .B2(\mem[21][5] ), 
        .ZN(n437) );
  INV_X1 U433 ( .A(n438), .ZN(n710) );
  AOI22_X1 U434 ( .A1(data_in[6]), .A2(n831), .B1(n432), .B2(\mem[21][6] ), 
        .ZN(n438) );
  INV_X1 U435 ( .A(n439), .ZN(n709) );
  AOI22_X1 U436 ( .A1(data_in[7]), .A2(n831), .B1(n432), .B2(\mem[21][7] ), 
        .ZN(n439) );
  INV_X1 U437 ( .A(n440), .ZN(n708) );
  AOI22_X1 U438 ( .A1(data_in[0]), .A2(n830), .B1(n441), .B2(\mem[22][0] ), 
        .ZN(n440) );
  INV_X1 U439 ( .A(n442), .ZN(n707) );
  AOI22_X1 U440 ( .A1(data_in[1]), .A2(n830), .B1(n441), .B2(\mem[22][1] ), 
        .ZN(n442) );
  INV_X1 U441 ( .A(n443), .ZN(n706) );
  AOI22_X1 U442 ( .A1(data_in[2]), .A2(n830), .B1(n441), .B2(\mem[22][2] ), 
        .ZN(n443) );
  INV_X1 U443 ( .A(n444), .ZN(n705) );
  AOI22_X1 U444 ( .A1(data_in[3]), .A2(n830), .B1(n441), .B2(\mem[22][3] ), 
        .ZN(n444) );
  INV_X1 U445 ( .A(n445), .ZN(n704) );
  AOI22_X1 U446 ( .A1(data_in[4]), .A2(n830), .B1(n441), .B2(\mem[22][4] ), 
        .ZN(n445) );
  INV_X1 U447 ( .A(n446), .ZN(n703) );
  AOI22_X1 U448 ( .A1(data_in[5]), .A2(n830), .B1(n441), .B2(\mem[22][5] ), 
        .ZN(n446) );
  INV_X1 U449 ( .A(n447), .ZN(n702) );
  AOI22_X1 U450 ( .A1(data_in[6]), .A2(n830), .B1(n441), .B2(\mem[22][6] ), 
        .ZN(n447) );
  INV_X1 U451 ( .A(n448), .ZN(n701) );
  AOI22_X1 U452 ( .A1(data_in[7]), .A2(n830), .B1(n441), .B2(\mem[22][7] ), 
        .ZN(n448) );
  INV_X1 U453 ( .A(n449), .ZN(n700) );
  AOI22_X1 U454 ( .A1(data_in[0]), .A2(n829), .B1(n450), .B2(\mem[23][0] ), 
        .ZN(n449) );
  INV_X1 U455 ( .A(n451), .ZN(n699) );
  AOI22_X1 U456 ( .A1(data_in[1]), .A2(n829), .B1(n450), .B2(\mem[23][1] ), 
        .ZN(n451) );
  INV_X1 U457 ( .A(n452), .ZN(n698) );
  AOI22_X1 U458 ( .A1(data_in[2]), .A2(n829), .B1(n450), .B2(\mem[23][2] ), 
        .ZN(n452) );
  INV_X1 U459 ( .A(n453), .ZN(n697) );
  AOI22_X1 U460 ( .A1(data_in[3]), .A2(n829), .B1(n450), .B2(\mem[23][3] ), 
        .ZN(n453) );
  INV_X1 U461 ( .A(n454), .ZN(n696) );
  AOI22_X1 U462 ( .A1(data_in[4]), .A2(n829), .B1(n450), .B2(\mem[23][4] ), 
        .ZN(n454) );
  INV_X1 U463 ( .A(n455), .ZN(n695) );
  AOI22_X1 U464 ( .A1(data_in[5]), .A2(n829), .B1(n450), .B2(\mem[23][5] ), 
        .ZN(n455) );
  INV_X1 U465 ( .A(n456), .ZN(n694) );
  AOI22_X1 U466 ( .A1(data_in[6]), .A2(n829), .B1(n450), .B2(\mem[23][6] ), 
        .ZN(n456) );
  INV_X1 U467 ( .A(n457), .ZN(n693) );
  AOI22_X1 U468 ( .A1(data_in[7]), .A2(n829), .B1(n450), .B2(\mem[23][7] ), 
        .ZN(n457) );
  INV_X1 U469 ( .A(n458), .ZN(n692) );
  AOI22_X1 U470 ( .A1(data_in[0]), .A2(n828), .B1(n459), .B2(\mem[24][0] ), 
        .ZN(n458) );
  INV_X1 U471 ( .A(n460), .ZN(n691) );
  AOI22_X1 U472 ( .A1(data_in[1]), .A2(n828), .B1(n459), .B2(\mem[24][1] ), 
        .ZN(n460) );
  INV_X1 U473 ( .A(n461), .ZN(n690) );
  AOI22_X1 U474 ( .A1(data_in[2]), .A2(n828), .B1(n459), .B2(\mem[24][2] ), 
        .ZN(n461) );
  INV_X1 U475 ( .A(n462), .ZN(n689) );
  AOI22_X1 U476 ( .A1(data_in[3]), .A2(n828), .B1(n459), .B2(\mem[24][3] ), 
        .ZN(n462) );
  INV_X1 U477 ( .A(n463), .ZN(n688) );
  AOI22_X1 U478 ( .A1(data_in[4]), .A2(n828), .B1(n459), .B2(\mem[24][4] ), 
        .ZN(n463) );
  INV_X1 U479 ( .A(n464), .ZN(n687) );
  AOI22_X1 U480 ( .A1(data_in[5]), .A2(n828), .B1(n459), .B2(\mem[24][5] ), 
        .ZN(n464) );
  INV_X1 U481 ( .A(n465), .ZN(n686) );
  AOI22_X1 U482 ( .A1(data_in[6]), .A2(n828), .B1(n459), .B2(\mem[24][6] ), 
        .ZN(n465) );
  INV_X1 U483 ( .A(n466), .ZN(n685) );
  AOI22_X1 U484 ( .A1(data_in[7]), .A2(n828), .B1(n459), .B2(\mem[24][7] ), 
        .ZN(n466) );
  INV_X1 U485 ( .A(n468), .ZN(n684) );
  AOI22_X1 U486 ( .A1(data_in[0]), .A2(n827), .B1(n469), .B2(\mem[25][0] ), 
        .ZN(n468) );
  INV_X1 U487 ( .A(n470), .ZN(n683) );
  AOI22_X1 U488 ( .A1(data_in[1]), .A2(n827), .B1(n469), .B2(\mem[25][1] ), 
        .ZN(n470) );
  INV_X1 U489 ( .A(n471), .ZN(n682) );
  AOI22_X1 U490 ( .A1(data_in[2]), .A2(n827), .B1(n469), .B2(\mem[25][2] ), 
        .ZN(n471) );
  INV_X1 U491 ( .A(n472), .ZN(n681) );
  AOI22_X1 U492 ( .A1(data_in[3]), .A2(n827), .B1(n469), .B2(\mem[25][3] ), 
        .ZN(n472) );
  INV_X1 U493 ( .A(n473), .ZN(n680) );
  AOI22_X1 U494 ( .A1(data_in[4]), .A2(n827), .B1(n469), .B2(\mem[25][4] ), 
        .ZN(n473) );
  INV_X1 U495 ( .A(n474), .ZN(n679) );
  AOI22_X1 U496 ( .A1(data_in[5]), .A2(n827), .B1(n469), .B2(\mem[25][5] ), 
        .ZN(n474) );
  INV_X1 U497 ( .A(n475), .ZN(n678) );
  AOI22_X1 U498 ( .A1(data_in[6]), .A2(n827), .B1(n469), .B2(\mem[25][6] ), 
        .ZN(n475) );
  INV_X1 U499 ( .A(n476), .ZN(n677) );
  AOI22_X1 U500 ( .A1(data_in[7]), .A2(n827), .B1(n469), .B2(\mem[25][7] ), 
        .ZN(n476) );
  INV_X1 U501 ( .A(n477), .ZN(n676) );
  AOI22_X1 U502 ( .A1(data_in[0]), .A2(n826), .B1(n478), .B2(\mem[26][0] ), 
        .ZN(n477) );
  INV_X1 U503 ( .A(n479), .ZN(n675) );
  AOI22_X1 U504 ( .A1(data_in[1]), .A2(n826), .B1(n478), .B2(\mem[26][1] ), 
        .ZN(n479) );
  INV_X1 U505 ( .A(n480), .ZN(n674) );
  AOI22_X1 U506 ( .A1(data_in[2]), .A2(n826), .B1(n478), .B2(\mem[26][2] ), 
        .ZN(n480) );
  INV_X1 U507 ( .A(n481), .ZN(n673) );
  AOI22_X1 U508 ( .A1(data_in[3]), .A2(n826), .B1(n478), .B2(\mem[26][3] ), 
        .ZN(n481) );
  INV_X1 U509 ( .A(n482), .ZN(n672) );
  AOI22_X1 U510 ( .A1(data_in[4]), .A2(n826), .B1(n478), .B2(\mem[26][4] ), 
        .ZN(n482) );
  INV_X1 U511 ( .A(n483), .ZN(n671) );
  AOI22_X1 U512 ( .A1(data_in[5]), .A2(n826), .B1(n478), .B2(\mem[26][5] ), 
        .ZN(n483) );
  INV_X1 U513 ( .A(n484), .ZN(n670) );
  AOI22_X1 U514 ( .A1(data_in[6]), .A2(n826), .B1(n478), .B2(\mem[26][6] ), 
        .ZN(n484) );
  INV_X1 U515 ( .A(n485), .ZN(n669) );
  AOI22_X1 U516 ( .A1(data_in[7]), .A2(n826), .B1(n478), .B2(\mem[26][7] ), 
        .ZN(n485) );
  INV_X1 U517 ( .A(n486), .ZN(n668) );
  AOI22_X1 U518 ( .A1(data_in[0]), .A2(n825), .B1(n487), .B2(\mem[27][0] ), 
        .ZN(n486) );
  INV_X1 U519 ( .A(n488), .ZN(n667) );
  AOI22_X1 U520 ( .A1(data_in[1]), .A2(n825), .B1(n487), .B2(\mem[27][1] ), 
        .ZN(n488) );
  INV_X1 U521 ( .A(n489), .ZN(n666) );
  AOI22_X1 U522 ( .A1(data_in[2]), .A2(n825), .B1(n487), .B2(\mem[27][2] ), 
        .ZN(n489) );
  INV_X1 U523 ( .A(n490), .ZN(n665) );
  AOI22_X1 U524 ( .A1(data_in[3]), .A2(n825), .B1(n487), .B2(\mem[27][3] ), 
        .ZN(n490) );
  INV_X1 U525 ( .A(n491), .ZN(n664) );
  AOI22_X1 U526 ( .A1(data_in[4]), .A2(n825), .B1(n487), .B2(\mem[27][4] ), 
        .ZN(n491) );
  INV_X1 U527 ( .A(n492), .ZN(n663) );
  AOI22_X1 U528 ( .A1(data_in[5]), .A2(n825), .B1(n487), .B2(\mem[27][5] ), 
        .ZN(n492) );
  INV_X1 U529 ( .A(n493), .ZN(n662) );
  AOI22_X1 U530 ( .A1(data_in[6]), .A2(n825), .B1(n487), .B2(\mem[27][6] ), 
        .ZN(n493) );
  INV_X1 U531 ( .A(n494), .ZN(n661) );
  AOI22_X1 U532 ( .A1(data_in[7]), .A2(n825), .B1(n487), .B2(\mem[27][7] ), 
        .ZN(n494) );
  INV_X1 U533 ( .A(n495), .ZN(n660) );
  AOI22_X1 U534 ( .A1(data_in[0]), .A2(n824), .B1(n496), .B2(\mem[28][0] ), 
        .ZN(n495) );
  INV_X1 U535 ( .A(n497), .ZN(n659) );
  AOI22_X1 U536 ( .A1(data_in[1]), .A2(n824), .B1(n496), .B2(\mem[28][1] ), 
        .ZN(n497) );
  INV_X1 U537 ( .A(n498), .ZN(n658) );
  AOI22_X1 U538 ( .A1(data_in[2]), .A2(n824), .B1(n496), .B2(\mem[28][2] ), 
        .ZN(n498) );
  INV_X1 U539 ( .A(n499), .ZN(n657) );
  AOI22_X1 U540 ( .A1(data_in[3]), .A2(n824), .B1(n496), .B2(\mem[28][3] ), 
        .ZN(n499) );
  INV_X1 U541 ( .A(n500), .ZN(n656) );
  AOI22_X1 U542 ( .A1(data_in[4]), .A2(n824), .B1(n496), .B2(\mem[28][4] ), 
        .ZN(n500) );
  INV_X1 U543 ( .A(n501), .ZN(n655) );
  AOI22_X1 U544 ( .A1(data_in[5]), .A2(n824), .B1(n496), .B2(\mem[28][5] ), 
        .ZN(n501) );
  INV_X1 U545 ( .A(n502), .ZN(n654) );
  AOI22_X1 U546 ( .A1(data_in[6]), .A2(n824), .B1(n496), .B2(\mem[28][6] ), 
        .ZN(n502) );
  INV_X1 U547 ( .A(n503), .ZN(n653) );
  AOI22_X1 U548 ( .A1(data_in[7]), .A2(n824), .B1(n496), .B2(\mem[28][7] ), 
        .ZN(n503) );
  INV_X1 U549 ( .A(n504), .ZN(n652) );
  AOI22_X1 U550 ( .A1(data_in[0]), .A2(n823), .B1(n505), .B2(\mem[29][0] ), 
        .ZN(n504) );
  INV_X1 U551 ( .A(n506), .ZN(n651) );
  AOI22_X1 U552 ( .A1(data_in[1]), .A2(n823), .B1(n505), .B2(\mem[29][1] ), 
        .ZN(n506) );
  INV_X1 U553 ( .A(n507), .ZN(n650) );
  AOI22_X1 U554 ( .A1(data_in[2]), .A2(n823), .B1(n505), .B2(\mem[29][2] ), 
        .ZN(n507) );
  INV_X1 U555 ( .A(n508), .ZN(n649) );
  AOI22_X1 U556 ( .A1(data_in[3]), .A2(n823), .B1(n505), .B2(\mem[29][3] ), 
        .ZN(n508) );
  INV_X1 U557 ( .A(n509), .ZN(n648) );
  AOI22_X1 U558 ( .A1(data_in[4]), .A2(n823), .B1(n505), .B2(\mem[29][4] ), 
        .ZN(n509) );
  INV_X1 U559 ( .A(n510), .ZN(n647) );
  AOI22_X1 U560 ( .A1(data_in[5]), .A2(n823), .B1(n505), .B2(\mem[29][5] ), 
        .ZN(n510) );
  INV_X1 U561 ( .A(n511), .ZN(n646) );
  AOI22_X1 U562 ( .A1(data_in[6]), .A2(n823), .B1(n505), .B2(\mem[29][6] ), 
        .ZN(n511) );
  INV_X1 U563 ( .A(n512), .ZN(n645) );
  AOI22_X1 U564 ( .A1(data_in[7]), .A2(n823), .B1(n505), .B2(\mem[29][7] ), 
        .ZN(n512) );
  INV_X1 U565 ( .A(n513), .ZN(n644) );
  AOI22_X1 U566 ( .A1(data_in[0]), .A2(n822), .B1(n514), .B2(\mem[30][0] ), 
        .ZN(n513) );
  INV_X1 U567 ( .A(n515), .ZN(n643) );
  AOI22_X1 U568 ( .A1(data_in[1]), .A2(n822), .B1(n514), .B2(\mem[30][1] ), 
        .ZN(n515) );
  INV_X1 U569 ( .A(n516), .ZN(n642) );
  AOI22_X1 U570 ( .A1(data_in[2]), .A2(n822), .B1(n514), .B2(\mem[30][2] ), 
        .ZN(n516) );
  INV_X1 U571 ( .A(n517), .ZN(n641) );
  AOI22_X1 U572 ( .A1(data_in[3]), .A2(n822), .B1(n514), .B2(\mem[30][3] ), 
        .ZN(n517) );
  INV_X1 U573 ( .A(n518), .ZN(n640) );
  AOI22_X1 U574 ( .A1(data_in[4]), .A2(n822), .B1(n514), .B2(\mem[30][4] ), 
        .ZN(n518) );
  INV_X1 U575 ( .A(n519), .ZN(n639) );
  AOI22_X1 U576 ( .A1(data_in[5]), .A2(n822), .B1(n514), .B2(\mem[30][5] ), 
        .ZN(n519) );
  INV_X1 U577 ( .A(n520), .ZN(n638) );
  AOI22_X1 U578 ( .A1(data_in[6]), .A2(n822), .B1(n514), .B2(\mem[30][6] ), 
        .ZN(n520) );
  INV_X1 U579 ( .A(n521), .ZN(n637) );
  AOI22_X1 U580 ( .A1(data_in[7]), .A2(n822), .B1(n514), .B2(\mem[30][7] ), 
        .ZN(n521) );
  INV_X1 U581 ( .A(n522), .ZN(n636) );
  AOI22_X1 U582 ( .A1(data_in[0]), .A2(n821), .B1(n523), .B2(\mem[31][0] ), 
        .ZN(n522) );
  INV_X1 U583 ( .A(n524), .ZN(n635) );
  AOI22_X1 U584 ( .A1(data_in[1]), .A2(n821), .B1(n523), .B2(\mem[31][1] ), 
        .ZN(n524) );
  INV_X1 U585 ( .A(n525), .ZN(n634) );
  AOI22_X1 U586 ( .A1(data_in[2]), .A2(n821), .B1(n523), .B2(\mem[31][2] ), 
        .ZN(n525) );
  INV_X1 U587 ( .A(n526), .ZN(n633) );
  AOI22_X1 U588 ( .A1(data_in[3]), .A2(n821), .B1(n523), .B2(\mem[31][3] ), 
        .ZN(n526) );
  INV_X1 U589 ( .A(n527), .ZN(n632) );
  AOI22_X1 U590 ( .A1(data_in[4]), .A2(n821), .B1(n523), .B2(\mem[31][4] ), 
        .ZN(n527) );
  INV_X1 U591 ( .A(n528), .ZN(n631) );
  AOI22_X1 U592 ( .A1(data_in[5]), .A2(n821), .B1(n523), .B2(\mem[31][5] ), 
        .ZN(n528) );
  INV_X1 U593 ( .A(n529), .ZN(n630) );
  AOI22_X1 U594 ( .A1(data_in[6]), .A2(n821), .B1(n523), .B2(\mem[31][6] ), 
        .ZN(n529) );
  INV_X1 U595 ( .A(n530), .ZN(n629) );
  AOI22_X1 U596 ( .A1(data_in[7]), .A2(n821), .B1(n523), .B2(\mem[31][7] ), 
        .ZN(n530) );
  MUX2_X1 U597 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n613), .Z(n3) );
  MUX2_X1 U598 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n616), .Z(n4) );
  MUX2_X1 U599 ( .A(n4), .B(n3), .S(n610), .Z(n5) );
  MUX2_X1 U600 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n617), .Z(n6) );
  MUX2_X1 U601 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n613), .Z(n7) );
  MUX2_X1 U602 ( .A(n7), .B(n6), .S(n610), .Z(n8) );
  MUX2_X1 U603 ( .A(n8), .B(n5), .S(n608), .Z(n9) );
  MUX2_X1 U604 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n615), .Z(n10) );
  MUX2_X1 U605 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n616), .Z(n11) );
  MUX2_X1 U606 ( .A(n11), .B(n10), .S(n610), .Z(n12) );
  MUX2_X1 U607 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n617), .Z(n13) );
  MUX2_X1 U608 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n615), .Z(n14) );
  MUX2_X1 U609 ( .A(n14), .B(n13), .S(n610), .Z(n15) );
  MUX2_X1 U610 ( .A(n15), .B(n12), .S(N12), .Z(n16) );
  MUX2_X1 U611 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U612 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n613), .Z(n18) );
  MUX2_X1 U613 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n613), .Z(n19) );
  MUX2_X1 U614 ( .A(n19), .B(n18), .S(n612), .Z(n20) );
  MUX2_X1 U615 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n618), .Z(n21) );
  MUX2_X1 U616 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n22) );
  MUX2_X1 U617 ( .A(n22), .B(n21), .S(N11), .Z(n23) );
  MUX2_X1 U618 ( .A(n23), .B(n20), .S(N12), .Z(n24) );
  MUX2_X1 U619 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n614), .Z(n25) );
  MUX2_X1 U620 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n618), .Z(n26) );
  MUX2_X1 U621 ( .A(n26), .B(n25), .S(n612), .Z(n27) );
  MUX2_X1 U622 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n28) );
  MUX2_X1 U623 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n29) );
  MUX2_X1 U624 ( .A(n29), .B(n28), .S(N11), .Z(n30) );
  MUX2_X1 U625 ( .A(n30), .B(n27), .S(n609), .Z(n31) );
  MUX2_X1 U626 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U627 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U628 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n617), .Z(n33) );
  MUX2_X1 U629 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n617), .Z(n34) );
  MUX2_X1 U630 ( .A(n34), .B(n33), .S(n611), .Z(n35) );
  MUX2_X1 U631 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n616), .Z(n36) );
  MUX2_X1 U632 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n614), .Z(n37) );
  MUX2_X1 U633 ( .A(n37), .B(n36), .S(n612), .Z(n38) );
  MUX2_X1 U634 ( .A(n38), .B(n35), .S(n609), .Z(n39) );
  MUX2_X1 U635 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n614), .Z(n40) );
  MUX2_X1 U636 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n616), .Z(n41) );
  MUX2_X1 U637 ( .A(n41), .B(n40), .S(n610), .Z(n42) );
  MUX2_X1 U638 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n617), .Z(n43) );
  MUX2_X1 U639 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n618), .Z(n44) );
  MUX2_X1 U640 ( .A(n44), .B(n43), .S(N11), .Z(n45) );
  MUX2_X1 U641 ( .A(n45), .B(n42), .S(n608), .Z(n46) );
  MUX2_X1 U642 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U643 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n613), .Z(n48) );
  MUX2_X1 U644 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n615), .Z(n49) );
  MUX2_X1 U645 ( .A(n49), .B(n48), .S(n610), .Z(n50) );
  MUX2_X1 U646 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n616), .Z(n51) );
  MUX2_X1 U647 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(N10), .Z(n52) );
  MUX2_X1 U648 ( .A(n52), .B(n51), .S(N11), .Z(n53) );
  MUX2_X1 U649 ( .A(n53), .B(n50), .S(N12), .Z(n54) );
  MUX2_X1 U650 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n618), .Z(n55) );
  MUX2_X1 U651 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n618), .Z(n56) );
  MUX2_X1 U652 ( .A(n56), .B(n55), .S(n611), .Z(n57) );
  MUX2_X1 U653 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n617), .Z(n58) );
  MUX2_X1 U654 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(N10), .Z(n59) );
  MUX2_X1 U655 ( .A(n59), .B(n58), .S(n612), .Z(n60) );
  MUX2_X1 U656 ( .A(n60), .B(n57), .S(n608), .Z(n61) );
  MUX2_X1 U657 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U658 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U659 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n613), .Z(n63) );
  MUX2_X1 U660 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n613), .Z(n64) );
  MUX2_X1 U661 ( .A(n64), .B(n63), .S(n610), .Z(n65) );
  MUX2_X1 U662 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n613), .Z(n66) );
  MUX2_X1 U663 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n613), .Z(n67) );
  MUX2_X1 U664 ( .A(n67), .B(n66), .S(n610), .Z(n68) );
  MUX2_X1 U665 ( .A(n68), .B(n65), .S(n608), .Z(n69) );
  MUX2_X1 U666 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n613), .Z(n70) );
  MUX2_X1 U667 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n613), .Z(n71) );
  MUX2_X1 U668 ( .A(n71), .B(n70), .S(n610), .Z(n72) );
  MUX2_X1 U669 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n613), .Z(n73) );
  MUX2_X1 U670 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n613), .Z(n74) );
  MUX2_X1 U671 ( .A(n74), .B(n73), .S(n610), .Z(n75) );
  MUX2_X1 U672 ( .A(n75), .B(n72), .S(n608), .Z(n76) );
  MUX2_X1 U673 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U674 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n613), .Z(n78) );
  MUX2_X1 U675 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n613), .Z(n79) );
  MUX2_X1 U676 ( .A(n79), .B(n78), .S(n610), .Z(n80) );
  MUX2_X1 U677 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n613), .Z(n81) );
  MUX2_X1 U678 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n613), .Z(n82) );
  MUX2_X1 U679 ( .A(n82), .B(n81), .S(n610), .Z(n83) );
  MUX2_X1 U680 ( .A(n83), .B(n80), .S(n608), .Z(n84) );
  MUX2_X1 U681 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n614), .Z(n85) );
  MUX2_X1 U682 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n614), .Z(n86) );
  MUX2_X1 U683 ( .A(n86), .B(n85), .S(n610), .Z(n87) );
  MUX2_X1 U684 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n614), .Z(n88) );
  MUX2_X1 U685 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n614), .Z(n89) );
  MUX2_X1 U686 ( .A(n89), .B(n88), .S(n611), .Z(n90) );
  MUX2_X1 U687 ( .A(n90), .B(n87), .S(n608), .Z(n91) );
  MUX2_X1 U688 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U689 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U690 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n614), .Z(n93) );
  MUX2_X1 U691 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n614), .Z(n94) );
  MUX2_X1 U692 ( .A(n94), .B(n93), .S(n612), .Z(n95) );
  MUX2_X1 U693 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n614), .Z(n96) );
  MUX2_X1 U694 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n614), .Z(n97) );
  MUX2_X1 U695 ( .A(n97), .B(n96), .S(n612), .Z(n98) );
  MUX2_X1 U696 ( .A(n98), .B(n95), .S(n608), .Z(n99) );
  MUX2_X1 U697 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n614), .Z(n100) );
  MUX2_X1 U698 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n614), .Z(n101) );
  MUX2_X1 U699 ( .A(n101), .B(n100), .S(n610), .Z(n102) );
  MUX2_X1 U700 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n614), .Z(n103) );
  MUX2_X1 U701 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n614), .Z(n104) );
  MUX2_X1 U702 ( .A(n104), .B(n103), .S(n610), .Z(n105) );
  MUX2_X1 U703 ( .A(n105), .B(n102), .S(n608), .Z(n106) );
  MUX2_X1 U704 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U705 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n613), .Z(n108) );
  MUX2_X1 U706 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n618), .Z(n109) );
  MUX2_X1 U707 ( .A(n109), .B(n108), .S(n611), .Z(n110) );
  MUX2_X1 U708 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n618), .Z(n111) );
  MUX2_X1 U709 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n613), .Z(n112) );
  MUX2_X1 U710 ( .A(n112), .B(n111), .S(n611), .Z(n113) );
  MUX2_X1 U711 ( .A(n113), .B(n110), .S(n608), .Z(n114) );
  MUX2_X1 U712 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n618), .Z(n115) );
  MUX2_X1 U713 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n616), .Z(n116) );
  MUX2_X1 U714 ( .A(n116), .B(n115), .S(n611), .Z(n117) );
  MUX2_X1 U715 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n618), .Z(n118) );
  MUX2_X1 U716 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n615), .Z(n119) );
  MUX2_X1 U717 ( .A(n119), .B(n118), .S(n611), .Z(n120) );
  MUX2_X1 U718 ( .A(n120), .B(n117), .S(n608), .Z(n121) );
  MUX2_X1 U719 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U720 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n616), .Z(n123) );
  MUX2_X1 U721 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n617), .Z(n124) );
  MUX2_X1 U722 ( .A(n124), .B(n123), .S(n611), .Z(n125) );
  MUX2_X1 U723 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n615), .Z(n126) );
  MUX2_X1 U724 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n615), .Z(n127) );
  MUX2_X1 U725 ( .A(n127), .B(n126), .S(n611), .Z(n128) );
  MUX2_X1 U726 ( .A(n128), .B(n125), .S(n608), .Z(n129) );
  MUX2_X1 U727 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n618), .Z(n130) );
  MUX2_X1 U728 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n618), .Z(n131) );
  MUX2_X1 U729 ( .A(n131), .B(n130), .S(n611), .Z(n132) );
  MUX2_X1 U730 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n618), .Z(n133) );
  MUX2_X1 U731 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n618), .Z(n134) );
  MUX2_X1 U732 ( .A(n134), .B(n133), .S(n611), .Z(n135) );
  MUX2_X1 U733 ( .A(n135), .B(n132), .S(n608), .Z(n136) );
  MUX2_X1 U734 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U735 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n615), .Z(n138) );
  MUX2_X1 U736 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n618), .Z(n139) );
  MUX2_X1 U737 ( .A(n139), .B(n138), .S(n611), .Z(n140) );
  MUX2_X1 U738 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n618), .Z(n141) );
  MUX2_X1 U739 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n618), .Z(n142) );
  MUX2_X1 U740 ( .A(n142), .B(n141), .S(n611), .Z(n143) );
  MUX2_X1 U741 ( .A(n143), .B(n140), .S(n608), .Z(n144) );
  MUX2_X1 U742 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n618), .Z(n145) );
  MUX2_X1 U743 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n618), .Z(n146) );
  MUX2_X1 U744 ( .A(n146), .B(n145), .S(n611), .Z(n147) );
  MUX2_X1 U745 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n618), .Z(n148) );
  MUX2_X1 U746 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n618), .Z(n149) );
  MUX2_X1 U747 ( .A(n149), .B(n148), .S(n611), .Z(n150) );
  MUX2_X1 U748 ( .A(n150), .B(n147), .S(n608), .Z(n151) );
  MUX2_X1 U749 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U750 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U751 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n614), .Z(n153) );
  MUX2_X1 U752 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n614), .Z(n154) );
  MUX2_X1 U753 ( .A(n154), .B(n153), .S(n612), .Z(n155) );
  MUX2_X1 U754 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n614), .Z(n156) );
  MUX2_X1 U755 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n614), .Z(n157) );
  MUX2_X1 U756 ( .A(n157), .B(n156), .S(n612), .Z(n158) );
  MUX2_X1 U757 ( .A(n158), .B(n155), .S(n609), .Z(n159) );
  MUX2_X1 U758 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n614), .Z(n160) );
  MUX2_X1 U759 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n614), .Z(n161) );
  MUX2_X1 U760 ( .A(n161), .B(n160), .S(n612), .Z(n162) );
  MUX2_X1 U761 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n614), .Z(n163) );
  MUX2_X1 U762 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n614), .Z(n164) );
  MUX2_X1 U763 ( .A(n164), .B(n163), .S(n612), .Z(n165) );
  MUX2_X1 U764 ( .A(n165), .B(n162), .S(n609), .Z(n166) );
  MUX2_X1 U765 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U766 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n616), .Z(n168) );
  MUX2_X1 U767 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n617), .Z(n169) );
  MUX2_X1 U768 ( .A(n169), .B(n168), .S(n612), .Z(n170) );
  MUX2_X1 U769 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n615), .Z(n171) );
  MUX2_X1 U770 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n613), .Z(n172) );
  MUX2_X1 U771 ( .A(n172), .B(n171), .S(n612), .Z(n173) );
  MUX2_X1 U772 ( .A(n173), .B(n170), .S(n609), .Z(n174) );
  MUX2_X1 U773 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n615), .Z(n175) );
  MUX2_X1 U774 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n615), .Z(n176) );
  MUX2_X1 U775 ( .A(n176), .B(n175), .S(n612), .Z(n177) );
  MUX2_X1 U776 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n615), .Z(n178) );
  MUX2_X1 U777 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n615), .Z(n179) );
  MUX2_X1 U778 ( .A(n179), .B(n178), .S(n612), .Z(n180) );
  MUX2_X1 U779 ( .A(n180), .B(n177), .S(n609), .Z(n181) );
  MUX2_X1 U780 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U781 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n615), .Z(n183) );
  MUX2_X1 U782 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n615), .Z(n184) );
  MUX2_X1 U783 ( .A(n184), .B(n183), .S(n612), .Z(n185) );
  MUX2_X1 U784 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n615), .Z(n186) );
  MUX2_X1 U785 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n615), .Z(n187) );
  MUX2_X1 U786 ( .A(n187), .B(n186), .S(n612), .Z(n188) );
  MUX2_X1 U787 ( .A(n188), .B(n185), .S(n609), .Z(n189) );
  MUX2_X1 U788 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n615), .Z(n190) );
  MUX2_X1 U789 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n615), .Z(n191) );
  MUX2_X1 U790 ( .A(n191), .B(n190), .S(n612), .Z(n192) );
  MUX2_X1 U791 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n615), .Z(n193) );
  MUX2_X1 U792 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n615), .Z(n194) );
  MUX2_X1 U793 ( .A(n194), .B(n193), .S(n612), .Z(n195) );
  MUX2_X1 U794 ( .A(n195), .B(n192), .S(n609), .Z(n196) );
  MUX2_X1 U795 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U796 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n616), .Z(n198) );
  MUX2_X1 U797 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n616), .Z(n199) );
  MUX2_X1 U798 ( .A(n199), .B(n198), .S(n612), .Z(n200) );
  MUX2_X1 U799 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n616), .Z(n201) );
  MUX2_X1 U800 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n616), .Z(n202) );
  MUX2_X1 U801 ( .A(n202), .B(n201), .S(n612), .Z(n203) );
  MUX2_X1 U802 ( .A(n203), .B(n200), .S(n609), .Z(n204) );
  MUX2_X1 U803 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n616), .Z(n205) );
  MUX2_X1 U804 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n616), .Z(n206) );
  MUX2_X1 U805 ( .A(n206), .B(n205), .S(n611), .Z(n207) );
  MUX2_X1 U806 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n616), .Z(n208) );
  MUX2_X1 U807 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n616), .Z(n209) );
  MUX2_X1 U808 ( .A(n209), .B(n208), .S(n612), .Z(n210) );
  MUX2_X1 U809 ( .A(n210), .B(n207), .S(n609), .Z(n211) );
  MUX2_X1 U810 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U811 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U812 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n616), .Z(n213) );
  MUX2_X1 U813 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n616), .Z(n214) );
  MUX2_X1 U814 ( .A(n214), .B(n213), .S(n611), .Z(n215) );
  MUX2_X1 U815 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n616), .Z(n216) );
  MUX2_X1 U816 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n616), .Z(n217) );
  MUX2_X1 U817 ( .A(n217), .B(n216), .S(N11), .Z(n218) );
  MUX2_X1 U818 ( .A(n218), .B(n215), .S(n609), .Z(n219) );
  MUX2_X1 U819 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n617), .Z(n220) );
  MUX2_X1 U820 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n617), .Z(n221) );
  MUX2_X1 U821 ( .A(n221), .B(n220), .S(n610), .Z(n222) );
  MUX2_X1 U822 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n617), .Z(n223) );
  MUX2_X1 U823 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n617), .Z(n224) );
  MUX2_X1 U824 ( .A(n224), .B(n223), .S(n610), .Z(n225) );
  MUX2_X1 U825 ( .A(n225), .B(n222), .S(n609), .Z(n226) );
  MUX2_X1 U826 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U827 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n617), .Z(n228) );
  MUX2_X1 U828 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n617), .Z(n229) );
  MUX2_X1 U829 ( .A(n229), .B(n228), .S(n611), .Z(n595) );
  MUX2_X1 U830 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n617), .Z(n596) );
  MUX2_X1 U831 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n617), .Z(n597) );
  MUX2_X1 U832 ( .A(n597), .B(n596), .S(n611), .Z(n598) );
  MUX2_X1 U833 ( .A(n598), .B(n595), .S(n609), .Z(n599) );
  MUX2_X1 U834 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n617), .Z(n600) );
  MUX2_X1 U835 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n617), .Z(n601) );
  MUX2_X1 U836 ( .A(n601), .B(n600), .S(n610), .Z(n602) );
  MUX2_X1 U837 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n617), .Z(n603) );
  MUX2_X1 U838 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n617), .Z(n604) );
  MUX2_X1 U839 ( .A(n604), .B(n603), .S(n611), .Z(n605) );
  MUX2_X1 U840 ( .A(n605), .B(n602), .S(n609), .Z(n606) );
  MUX2_X1 U841 ( .A(n606), .B(n599), .S(N13), .Z(n607) );
  MUX2_X1 U842 ( .A(n607), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U843 ( .A(N11), .Z(n610) );
  INV_X1 U844 ( .A(N10), .ZN(n619) );
  INV_X1 U845 ( .A(N11), .ZN(n620) );
  INV_X1 U846 ( .A(data_in[0]), .ZN(n621) );
  INV_X1 U847 ( .A(data_in[1]), .ZN(n622) );
  INV_X1 U848 ( .A(data_in[2]), .ZN(n623) );
  INV_X1 U849 ( .A(data_in[3]), .ZN(n624) );
  INV_X1 U850 ( .A(data_in[4]), .ZN(n625) );
  INV_X1 U851 ( .A(data_in[5]), .ZN(n626) );
  INV_X1 U852 ( .A(data_in[6]), .ZN(n627) );
  INV_X1 U853 ( .A(data_in[7]), .ZN(n628) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_31 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n629), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n630), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n631), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n632), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n633), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n634), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n635), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n636), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n637), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n638), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n639), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n640), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n641), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n642), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n643), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n644), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n645), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n646), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n647), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n648), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n649), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n650), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n651), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n652), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n653), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n654), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n655), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n656), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n657), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n658), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n659), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n660), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n661), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n662), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n663), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n664), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n665), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n666), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n667), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n668), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n669), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n670), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n671), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n672), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n673), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n674), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n675), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n676), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n677), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n678), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n679), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n680), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n681), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n682), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n683), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n684), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n685), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n686), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n687), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n688), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n689), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n690), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n691), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n692), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n693), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n694), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n695), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n696), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n697), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n698), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n699), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n700), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n701), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n702), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n703), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n704), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n705), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n706), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n707), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n708), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n709), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n710), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n711), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n712), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n713), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n714), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n715), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n716), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n717), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n718), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n719), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n720), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n721), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n722), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n723), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n724), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n725), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n726), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n727), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n728), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n729), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n730), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n731), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n732), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n733), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n734), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n735), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n736), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n737), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n738), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n739), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n740), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n741), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n742), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n743), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n744), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n745), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n746), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n747), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n748), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n749), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n750), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n751), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n752), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n753), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n754), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n755), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n756), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n757), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n758), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n759), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n760), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n761), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n762), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n763), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n764), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n765), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n766), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n767), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n768), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n769), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n770), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n771), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n772), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n773), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n774), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n775), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n776), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n777), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n778), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n779), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n780), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n781), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n782), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n783), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n784), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n785), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n786), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n787), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n788), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n789), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n790), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n791), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n792), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n793), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n794), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n795), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n796), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n797), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n798), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n799), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n800), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n801), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n802), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n803), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n804), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n805), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n806), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n807), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n808), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n809), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n810), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n811), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n812), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n813), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n814), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n815), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n816), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n817), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n818), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n819), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n820), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n848), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n849), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n850), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n851), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n852), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n853), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n854), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n855), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n856), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n857), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n858), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n859), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n860), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n861), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n862), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n863), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n864), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n865), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n866), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n867), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n868), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n869), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n870), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n871), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n872), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n873), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n874), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n875), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n876), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n877), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n878), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n879), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n880), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n881), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n882), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n883), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n884), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n885), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n886), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n887), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n888), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n889), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n890), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n891), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n892), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n893), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n894), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n895), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n896), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n897), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n898), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n899), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n900), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n901), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n902), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n903), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n904), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n905), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n906), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n907), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n908), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n909), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n910), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n911), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n617), .Z(n613) );
  INV_X2 U4 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U5 ( .A(n617), .Z(n615) );
  BUF_X1 U6 ( .A(n617), .Z(n614) );
  BUF_X1 U7 ( .A(n617), .Z(n616) );
  BUF_X1 U8 ( .A(N11), .Z(n611) );
  BUF_X1 U9 ( .A(N11), .Z(n612) );
  BUF_X1 U10 ( .A(N10), .Z(n618) );
  BUF_X1 U11 ( .A(N10), .Z(n617) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1203) );
  NOR3_X1 U13 ( .A1(N11), .A2(N12), .A3(n619), .ZN(n1192) );
  NOR3_X1 U14 ( .A1(N10), .A2(N12), .A3(n620), .ZN(n1182) );
  NOR3_X1 U15 ( .A1(n619), .A2(N12), .A3(n620), .ZN(n1172) );
  INV_X1 U16 ( .A(n1129), .ZN(n844) );
  INV_X1 U17 ( .A(n1119), .ZN(n843) );
  INV_X1 U18 ( .A(n1110), .ZN(n842) );
  INV_X1 U19 ( .A(n1101), .ZN(n841) );
  INV_X1 U20 ( .A(n1056), .ZN(n836) );
  INV_X1 U21 ( .A(n1046), .ZN(n835) );
  INV_X1 U22 ( .A(n1037), .ZN(n834) );
  INV_X1 U23 ( .A(n1028), .ZN(n833) );
  INV_X1 U24 ( .A(n983), .ZN(n828) );
  INV_X1 U25 ( .A(n973), .ZN(n827) );
  INV_X1 U26 ( .A(n964), .ZN(n826) );
  INV_X1 U27 ( .A(n955), .ZN(n825) );
  INV_X1 U28 ( .A(n1092), .ZN(n840) );
  INV_X1 U29 ( .A(n1083), .ZN(n839) );
  INV_X1 U30 ( .A(n1074), .ZN(n838) );
  INV_X1 U31 ( .A(n1065), .ZN(n837) );
  INV_X1 U32 ( .A(n946), .ZN(n824) );
  INV_X1 U33 ( .A(n937), .ZN(n823) );
  INV_X1 U34 ( .A(n928), .ZN(n822) );
  INV_X1 U35 ( .A(n919), .ZN(n821) );
  INV_X1 U36 ( .A(n1019), .ZN(n832) );
  INV_X1 U37 ( .A(n1010), .ZN(n831) );
  INV_X1 U38 ( .A(n1001), .ZN(n830) );
  INV_X1 U39 ( .A(n992), .ZN(n829) );
  BUF_X1 U40 ( .A(N12), .Z(n609) );
  INV_X1 U41 ( .A(N13), .ZN(n846) );
  AND3_X1 U42 ( .A1(n619), .A2(n620), .A3(N12), .ZN(n1162) );
  AND3_X1 U43 ( .A1(N10), .A2(n620), .A3(N12), .ZN(n1152) );
  AND3_X1 U44 ( .A1(N11), .A2(n619), .A3(N12), .ZN(n1142) );
  AND3_X1 U45 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1132) );
  BUF_X1 U46 ( .A(N12), .Z(n608) );
  INV_X1 U47 ( .A(N14), .ZN(n847) );
  NAND2_X1 U48 ( .A1(n1192), .A2(n1202), .ZN(n1201) );
  NAND2_X1 U49 ( .A1(n1182), .A2(n1202), .ZN(n1191) );
  NAND2_X1 U50 ( .A1(n1172), .A2(n1202), .ZN(n1181) );
  NAND2_X1 U51 ( .A1(n1162), .A2(n1202), .ZN(n1171) );
  NAND2_X1 U52 ( .A1(n1152), .A2(n1202), .ZN(n1161) );
  NAND2_X1 U53 ( .A1(n1142), .A2(n1202), .ZN(n1151) );
  NAND2_X1 U54 ( .A1(n1132), .A2(n1202), .ZN(n1141) );
  NAND2_X1 U55 ( .A1(n1203), .A2(n1202), .ZN(n1212) );
  NAND2_X1 U56 ( .A1(n1121), .A2(n1203), .ZN(n1129) );
  NAND2_X1 U57 ( .A1(n1121), .A2(n1192), .ZN(n1119) );
  NAND2_X1 U58 ( .A1(n1121), .A2(n1182), .ZN(n1110) );
  NAND2_X1 U59 ( .A1(n1121), .A2(n1172), .ZN(n1101) );
  NAND2_X1 U60 ( .A1(n1048), .A2(n1203), .ZN(n1056) );
  NAND2_X1 U61 ( .A1(n1048), .A2(n1192), .ZN(n1046) );
  NAND2_X1 U62 ( .A1(n1048), .A2(n1182), .ZN(n1037) );
  NAND2_X1 U63 ( .A1(n1048), .A2(n1172), .ZN(n1028) );
  NAND2_X1 U64 ( .A1(n975), .A2(n1203), .ZN(n983) );
  NAND2_X1 U65 ( .A1(n975), .A2(n1192), .ZN(n973) );
  NAND2_X1 U66 ( .A1(n975), .A2(n1182), .ZN(n964) );
  NAND2_X1 U67 ( .A1(n975), .A2(n1172), .ZN(n955) );
  NAND2_X1 U68 ( .A1(n1121), .A2(n1162), .ZN(n1092) );
  NAND2_X1 U69 ( .A1(n1121), .A2(n1152), .ZN(n1083) );
  NAND2_X1 U70 ( .A1(n1121), .A2(n1142), .ZN(n1074) );
  NAND2_X1 U71 ( .A1(n1121), .A2(n1132), .ZN(n1065) );
  NAND2_X1 U72 ( .A1(n1048), .A2(n1162), .ZN(n1019) );
  NAND2_X1 U73 ( .A1(n1048), .A2(n1152), .ZN(n1010) );
  NAND2_X1 U74 ( .A1(n1048), .A2(n1142), .ZN(n1001) );
  NAND2_X1 U75 ( .A1(n1048), .A2(n1132), .ZN(n992) );
  NAND2_X1 U76 ( .A1(n975), .A2(n1162), .ZN(n946) );
  NAND2_X1 U77 ( .A1(n975), .A2(n1152), .ZN(n937) );
  NAND2_X1 U78 ( .A1(n975), .A2(n1142), .ZN(n928) );
  NAND2_X1 U79 ( .A1(n975), .A2(n1132), .ZN(n919) );
  AND3_X1 U80 ( .A1(n846), .A2(n847), .A3(n1131), .ZN(n1202) );
  AND3_X1 U81 ( .A1(N13), .A2(n1131), .A3(N14), .ZN(n975) );
  AND3_X1 U82 ( .A1(n1131), .A2(n847), .A3(N13), .ZN(n1121) );
  AND3_X1 U83 ( .A1(n1131), .A2(n846), .A3(N14), .ZN(n1048) );
  NOR2_X1 U84 ( .A1(n845), .A2(addr[5]), .ZN(n1131) );
  INV_X1 U85 ( .A(wr_en), .ZN(n845) );
  OAI21_X1 U86 ( .B1(n621), .B2(n1171), .A(n1170), .ZN(n879) );
  NAND2_X1 U87 ( .A1(\mem[4][0] ), .A2(n1171), .ZN(n1170) );
  OAI21_X1 U88 ( .B1(n622), .B2(n1171), .A(n1169), .ZN(n878) );
  NAND2_X1 U89 ( .A1(\mem[4][1] ), .A2(n1171), .ZN(n1169) );
  OAI21_X1 U90 ( .B1(n623), .B2(n1171), .A(n1168), .ZN(n877) );
  NAND2_X1 U91 ( .A1(\mem[4][2] ), .A2(n1171), .ZN(n1168) );
  OAI21_X1 U92 ( .B1(n624), .B2(n1171), .A(n1167), .ZN(n876) );
  NAND2_X1 U93 ( .A1(\mem[4][3] ), .A2(n1171), .ZN(n1167) );
  OAI21_X1 U94 ( .B1(n625), .B2(n1171), .A(n1166), .ZN(n875) );
  NAND2_X1 U95 ( .A1(\mem[4][4] ), .A2(n1171), .ZN(n1166) );
  OAI21_X1 U96 ( .B1(n626), .B2(n1171), .A(n1165), .ZN(n874) );
  NAND2_X1 U97 ( .A1(\mem[4][5] ), .A2(n1171), .ZN(n1165) );
  OAI21_X1 U98 ( .B1(n627), .B2(n1171), .A(n1164), .ZN(n873) );
  NAND2_X1 U99 ( .A1(\mem[4][6] ), .A2(n1171), .ZN(n1164) );
  OAI21_X1 U100 ( .B1(n628), .B2(n1171), .A(n1163), .ZN(n872) );
  NAND2_X1 U101 ( .A1(\mem[4][7] ), .A2(n1171), .ZN(n1163) );
  OAI21_X1 U102 ( .B1(n621), .B2(n1151), .A(n1150), .ZN(n863) );
  NAND2_X1 U103 ( .A1(\mem[6][0] ), .A2(n1151), .ZN(n1150) );
  OAI21_X1 U104 ( .B1(n622), .B2(n1151), .A(n1149), .ZN(n862) );
  NAND2_X1 U105 ( .A1(\mem[6][1] ), .A2(n1151), .ZN(n1149) );
  OAI21_X1 U106 ( .B1(n623), .B2(n1151), .A(n1148), .ZN(n861) );
  NAND2_X1 U107 ( .A1(\mem[6][2] ), .A2(n1151), .ZN(n1148) );
  OAI21_X1 U108 ( .B1(n624), .B2(n1151), .A(n1147), .ZN(n860) );
  NAND2_X1 U109 ( .A1(\mem[6][3] ), .A2(n1151), .ZN(n1147) );
  OAI21_X1 U110 ( .B1(n625), .B2(n1151), .A(n1146), .ZN(n859) );
  NAND2_X1 U111 ( .A1(\mem[6][4] ), .A2(n1151), .ZN(n1146) );
  OAI21_X1 U112 ( .B1(n626), .B2(n1151), .A(n1145), .ZN(n858) );
  NAND2_X1 U113 ( .A1(\mem[6][5] ), .A2(n1151), .ZN(n1145) );
  OAI21_X1 U114 ( .B1(n627), .B2(n1151), .A(n1144), .ZN(n857) );
  NAND2_X1 U115 ( .A1(\mem[6][6] ), .A2(n1151), .ZN(n1144) );
  OAI21_X1 U116 ( .B1(n628), .B2(n1151), .A(n1143), .ZN(n856) );
  NAND2_X1 U117 ( .A1(\mem[6][7] ), .A2(n1151), .ZN(n1143) );
  OAI21_X1 U118 ( .B1(n621), .B2(n1141), .A(n1140), .ZN(n855) );
  NAND2_X1 U119 ( .A1(\mem[7][0] ), .A2(n1141), .ZN(n1140) );
  OAI21_X1 U120 ( .B1(n622), .B2(n1141), .A(n1139), .ZN(n854) );
  NAND2_X1 U121 ( .A1(\mem[7][1] ), .A2(n1141), .ZN(n1139) );
  OAI21_X1 U122 ( .B1(n623), .B2(n1141), .A(n1138), .ZN(n853) );
  NAND2_X1 U123 ( .A1(\mem[7][2] ), .A2(n1141), .ZN(n1138) );
  OAI21_X1 U124 ( .B1(n624), .B2(n1141), .A(n1137), .ZN(n852) );
  NAND2_X1 U125 ( .A1(\mem[7][3] ), .A2(n1141), .ZN(n1137) );
  OAI21_X1 U126 ( .B1(n625), .B2(n1141), .A(n1136), .ZN(n851) );
  NAND2_X1 U127 ( .A1(\mem[7][4] ), .A2(n1141), .ZN(n1136) );
  OAI21_X1 U128 ( .B1(n626), .B2(n1141), .A(n1135), .ZN(n850) );
  NAND2_X1 U129 ( .A1(\mem[7][5] ), .A2(n1141), .ZN(n1135) );
  OAI21_X1 U130 ( .B1(n627), .B2(n1141), .A(n1134), .ZN(n849) );
  NAND2_X1 U131 ( .A1(\mem[7][6] ), .A2(n1141), .ZN(n1134) );
  OAI21_X1 U132 ( .B1(n628), .B2(n1141), .A(n1133), .ZN(n848) );
  NAND2_X1 U133 ( .A1(\mem[7][7] ), .A2(n1141), .ZN(n1133) );
  OAI21_X1 U134 ( .B1(n621), .B2(n1201), .A(n1200), .ZN(n903) );
  NAND2_X1 U135 ( .A1(\mem[1][0] ), .A2(n1201), .ZN(n1200) );
  OAI21_X1 U136 ( .B1(n622), .B2(n1201), .A(n1199), .ZN(n902) );
  NAND2_X1 U137 ( .A1(\mem[1][1] ), .A2(n1201), .ZN(n1199) );
  OAI21_X1 U138 ( .B1(n623), .B2(n1201), .A(n1198), .ZN(n901) );
  NAND2_X1 U139 ( .A1(\mem[1][2] ), .A2(n1201), .ZN(n1198) );
  OAI21_X1 U140 ( .B1(n624), .B2(n1201), .A(n1197), .ZN(n900) );
  NAND2_X1 U141 ( .A1(\mem[1][3] ), .A2(n1201), .ZN(n1197) );
  OAI21_X1 U142 ( .B1(n625), .B2(n1201), .A(n1196), .ZN(n899) );
  NAND2_X1 U143 ( .A1(\mem[1][4] ), .A2(n1201), .ZN(n1196) );
  OAI21_X1 U144 ( .B1(n626), .B2(n1201), .A(n1195), .ZN(n898) );
  NAND2_X1 U145 ( .A1(\mem[1][5] ), .A2(n1201), .ZN(n1195) );
  OAI21_X1 U146 ( .B1(n627), .B2(n1201), .A(n1194), .ZN(n897) );
  NAND2_X1 U147 ( .A1(\mem[1][6] ), .A2(n1201), .ZN(n1194) );
  OAI21_X1 U148 ( .B1(n628), .B2(n1201), .A(n1193), .ZN(n896) );
  NAND2_X1 U149 ( .A1(\mem[1][7] ), .A2(n1201), .ZN(n1193) );
  OAI21_X1 U150 ( .B1(n621), .B2(n1191), .A(n1190), .ZN(n895) );
  NAND2_X1 U151 ( .A1(\mem[2][0] ), .A2(n1191), .ZN(n1190) );
  OAI21_X1 U152 ( .B1(n622), .B2(n1191), .A(n1189), .ZN(n894) );
  NAND2_X1 U153 ( .A1(\mem[2][1] ), .A2(n1191), .ZN(n1189) );
  OAI21_X1 U154 ( .B1(n623), .B2(n1191), .A(n1188), .ZN(n893) );
  NAND2_X1 U155 ( .A1(\mem[2][2] ), .A2(n1191), .ZN(n1188) );
  OAI21_X1 U156 ( .B1(n624), .B2(n1191), .A(n1187), .ZN(n892) );
  NAND2_X1 U157 ( .A1(\mem[2][3] ), .A2(n1191), .ZN(n1187) );
  OAI21_X1 U158 ( .B1(n625), .B2(n1191), .A(n1186), .ZN(n891) );
  NAND2_X1 U159 ( .A1(\mem[2][4] ), .A2(n1191), .ZN(n1186) );
  OAI21_X1 U160 ( .B1(n626), .B2(n1191), .A(n1185), .ZN(n890) );
  NAND2_X1 U161 ( .A1(\mem[2][5] ), .A2(n1191), .ZN(n1185) );
  OAI21_X1 U162 ( .B1(n627), .B2(n1191), .A(n1184), .ZN(n889) );
  NAND2_X1 U163 ( .A1(\mem[2][6] ), .A2(n1191), .ZN(n1184) );
  OAI21_X1 U164 ( .B1(n628), .B2(n1191), .A(n1183), .ZN(n888) );
  NAND2_X1 U165 ( .A1(\mem[2][7] ), .A2(n1191), .ZN(n1183) );
  OAI21_X1 U166 ( .B1(n621), .B2(n1181), .A(n1180), .ZN(n887) );
  NAND2_X1 U167 ( .A1(\mem[3][0] ), .A2(n1181), .ZN(n1180) );
  OAI21_X1 U168 ( .B1(n622), .B2(n1181), .A(n1179), .ZN(n886) );
  NAND2_X1 U169 ( .A1(\mem[3][1] ), .A2(n1181), .ZN(n1179) );
  OAI21_X1 U170 ( .B1(n623), .B2(n1181), .A(n1178), .ZN(n885) );
  NAND2_X1 U171 ( .A1(\mem[3][2] ), .A2(n1181), .ZN(n1178) );
  OAI21_X1 U172 ( .B1(n624), .B2(n1181), .A(n1177), .ZN(n884) );
  NAND2_X1 U173 ( .A1(\mem[3][3] ), .A2(n1181), .ZN(n1177) );
  OAI21_X1 U174 ( .B1(n625), .B2(n1181), .A(n1176), .ZN(n883) );
  NAND2_X1 U175 ( .A1(\mem[3][4] ), .A2(n1181), .ZN(n1176) );
  OAI21_X1 U176 ( .B1(n626), .B2(n1181), .A(n1175), .ZN(n882) );
  NAND2_X1 U177 ( .A1(\mem[3][5] ), .A2(n1181), .ZN(n1175) );
  OAI21_X1 U178 ( .B1(n627), .B2(n1181), .A(n1174), .ZN(n881) );
  NAND2_X1 U179 ( .A1(\mem[3][6] ), .A2(n1181), .ZN(n1174) );
  OAI21_X1 U180 ( .B1(n628), .B2(n1181), .A(n1173), .ZN(n880) );
  NAND2_X1 U181 ( .A1(\mem[3][7] ), .A2(n1181), .ZN(n1173) );
  OAI21_X1 U182 ( .B1(n621), .B2(n1161), .A(n1160), .ZN(n871) );
  NAND2_X1 U183 ( .A1(\mem[5][0] ), .A2(n1161), .ZN(n1160) );
  OAI21_X1 U184 ( .B1(n622), .B2(n1161), .A(n1159), .ZN(n870) );
  NAND2_X1 U185 ( .A1(\mem[5][1] ), .A2(n1161), .ZN(n1159) );
  OAI21_X1 U186 ( .B1(n623), .B2(n1161), .A(n1158), .ZN(n869) );
  NAND2_X1 U187 ( .A1(\mem[5][2] ), .A2(n1161), .ZN(n1158) );
  OAI21_X1 U188 ( .B1(n624), .B2(n1161), .A(n1157), .ZN(n868) );
  NAND2_X1 U189 ( .A1(\mem[5][3] ), .A2(n1161), .ZN(n1157) );
  OAI21_X1 U190 ( .B1(n625), .B2(n1161), .A(n1156), .ZN(n867) );
  NAND2_X1 U191 ( .A1(\mem[5][4] ), .A2(n1161), .ZN(n1156) );
  OAI21_X1 U192 ( .B1(n626), .B2(n1161), .A(n1155), .ZN(n866) );
  NAND2_X1 U193 ( .A1(\mem[5][5] ), .A2(n1161), .ZN(n1155) );
  OAI21_X1 U194 ( .B1(n627), .B2(n1161), .A(n1154), .ZN(n865) );
  NAND2_X1 U195 ( .A1(\mem[5][6] ), .A2(n1161), .ZN(n1154) );
  OAI21_X1 U196 ( .B1(n628), .B2(n1161), .A(n1153), .ZN(n864) );
  NAND2_X1 U197 ( .A1(\mem[5][7] ), .A2(n1161), .ZN(n1153) );
  OAI21_X1 U198 ( .B1(n1212), .B2(n621), .A(n1211), .ZN(n911) );
  NAND2_X1 U199 ( .A1(\mem[0][0] ), .A2(n1212), .ZN(n1211) );
  OAI21_X1 U200 ( .B1(n1212), .B2(n622), .A(n1210), .ZN(n910) );
  NAND2_X1 U201 ( .A1(\mem[0][1] ), .A2(n1212), .ZN(n1210) );
  OAI21_X1 U202 ( .B1(n1212), .B2(n623), .A(n1209), .ZN(n909) );
  NAND2_X1 U203 ( .A1(\mem[0][2] ), .A2(n1212), .ZN(n1209) );
  OAI21_X1 U204 ( .B1(n1212), .B2(n624), .A(n1208), .ZN(n908) );
  NAND2_X1 U205 ( .A1(\mem[0][3] ), .A2(n1212), .ZN(n1208) );
  OAI21_X1 U206 ( .B1(n1212), .B2(n625), .A(n1207), .ZN(n907) );
  NAND2_X1 U207 ( .A1(\mem[0][4] ), .A2(n1212), .ZN(n1207) );
  OAI21_X1 U208 ( .B1(n1212), .B2(n626), .A(n1206), .ZN(n906) );
  NAND2_X1 U209 ( .A1(\mem[0][5] ), .A2(n1212), .ZN(n1206) );
  OAI21_X1 U210 ( .B1(n1212), .B2(n627), .A(n1205), .ZN(n905) );
  NAND2_X1 U211 ( .A1(\mem[0][6] ), .A2(n1212), .ZN(n1205) );
  OAI21_X1 U212 ( .B1(n1212), .B2(n628), .A(n1204), .ZN(n904) );
  NAND2_X1 U213 ( .A1(\mem[0][7] ), .A2(n1212), .ZN(n1204) );
  INV_X1 U214 ( .A(n1130), .ZN(n820) );
  AOI22_X1 U215 ( .A1(data_in[0]), .A2(n844), .B1(n1129), .B2(\mem[8][0] ), 
        .ZN(n1130) );
  INV_X1 U216 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U217 ( .A1(data_in[1]), .A2(n844), .B1(n1129), .B2(\mem[8][1] ), 
        .ZN(n1128) );
  INV_X1 U218 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U219 ( .A1(data_in[2]), .A2(n844), .B1(n1129), .B2(\mem[8][2] ), 
        .ZN(n1127) );
  INV_X1 U220 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U221 ( .A1(data_in[3]), .A2(n844), .B1(n1129), .B2(\mem[8][3] ), 
        .ZN(n1126) );
  INV_X1 U222 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U223 ( .A1(data_in[4]), .A2(n844), .B1(n1129), .B2(\mem[8][4] ), 
        .ZN(n1125) );
  INV_X1 U224 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U225 ( .A1(data_in[5]), .A2(n844), .B1(n1129), .B2(\mem[8][5] ), 
        .ZN(n1124) );
  INV_X1 U226 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U227 ( .A1(data_in[6]), .A2(n844), .B1(n1129), .B2(\mem[8][6] ), 
        .ZN(n1123) );
  INV_X1 U228 ( .A(n1122), .ZN(n813) );
  AOI22_X1 U229 ( .A1(data_in[7]), .A2(n844), .B1(n1129), .B2(\mem[8][7] ), 
        .ZN(n1122) );
  INV_X1 U230 ( .A(n1120), .ZN(n812) );
  AOI22_X1 U231 ( .A1(data_in[0]), .A2(n843), .B1(n1119), .B2(\mem[9][0] ), 
        .ZN(n1120) );
  INV_X1 U232 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U233 ( .A1(data_in[1]), .A2(n843), .B1(n1119), .B2(\mem[9][1] ), 
        .ZN(n1118) );
  INV_X1 U234 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U235 ( .A1(data_in[2]), .A2(n843), .B1(n1119), .B2(\mem[9][2] ), 
        .ZN(n1117) );
  INV_X1 U236 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U237 ( .A1(data_in[3]), .A2(n843), .B1(n1119), .B2(\mem[9][3] ), 
        .ZN(n1116) );
  INV_X1 U238 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U239 ( .A1(data_in[4]), .A2(n843), .B1(n1119), .B2(\mem[9][4] ), 
        .ZN(n1115) );
  INV_X1 U240 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U241 ( .A1(data_in[5]), .A2(n843), .B1(n1119), .B2(\mem[9][5] ), 
        .ZN(n1114) );
  INV_X1 U242 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U243 ( .A1(data_in[6]), .A2(n843), .B1(n1119), .B2(\mem[9][6] ), 
        .ZN(n1113) );
  INV_X1 U244 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U245 ( .A1(data_in[7]), .A2(n843), .B1(n1119), .B2(\mem[9][7] ), 
        .ZN(n1112) );
  INV_X1 U246 ( .A(n1111), .ZN(n804) );
  AOI22_X1 U247 ( .A1(data_in[0]), .A2(n842), .B1(n1110), .B2(\mem[10][0] ), 
        .ZN(n1111) );
  INV_X1 U248 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U249 ( .A1(data_in[1]), .A2(n842), .B1(n1110), .B2(\mem[10][1] ), 
        .ZN(n1109) );
  INV_X1 U250 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U251 ( .A1(data_in[2]), .A2(n842), .B1(n1110), .B2(\mem[10][2] ), 
        .ZN(n1108) );
  INV_X1 U252 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U253 ( .A1(data_in[3]), .A2(n842), .B1(n1110), .B2(\mem[10][3] ), 
        .ZN(n1107) );
  INV_X1 U254 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U255 ( .A1(data_in[4]), .A2(n842), .B1(n1110), .B2(\mem[10][4] ), 
        .ZN(n1106) );
  INV_X1 U256 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U257 ( .A1(data_in[5]), .A2(n842), .B1(n1110), .B2(\mem[10][5] ), 
        .ZN(n1105) );
  INV_X1 U258 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U259 ( .A1(data_in[6]), .A2(n842), .B1(n1110), .B2(\mem[10][6] ), 
        .ZN(n1104) );
  INV_X1 U260 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U261 ( .A1(data_in[7]), .A2(n842), .B1(n1110), .B2(\mem[10][7] ), 
        .ZN(n1103) );
  INV_X1 U262 ( .A(n1102), .ZN(n796) );
  AOI22_X1 U263 ( .A1(data_in[0]), .A2(n841), .B1(n1101), .B2(\mem[11][0] ), 
        .ZN(n1102) );
  INV_X1 U264 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U265 ( .A1(data_in[1]), .A2(n841), .B1(n1101), .B2(\mem[11][1] ), 
        .ZN(n1100) );
  INV_X1 U266 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U267 ( .A1(data_in[2]), .A2(n841), .B1(n1101), .B2(\mem[11][2] ), 
        .ZN(n1099) );
  INV_X1 U268 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U269 ( .A1(data_in[3]), .A2(n841), .B1(n1101), .B2(\mem[11][3] ), 
        .ZN(n1098) );
  INV_X1 U270 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U271 ( .A1(data_in[4]), .A2(n841), .B1(n1101), .B2(\mem[11][4] ), 
        .ZN(n1097) );
  INV_X1 U272 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U273 ( .A1(data_in[5]), .A2(n841), .B1(n1101), .B2(\mem[11][5] ), 
        .ZN(n1096) );
  INV_X1 U274 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U275 ( .A1(data_in[6]), .A2(n841), .B1(n1101), .B2(\mem[11][6] ), 
        .ZN(n1095) );
  INV_X1 U276 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U277 ( .A1(data_in[7]), .A2(n841), .B1(n1101), .B2(\mem[11][7] ), 
        .ZN(n1094) );
  INV_X1 U278 ( .A(n1093), .ZN(n788) );
  AOI22_X1 U279 ( .A1(data_in[0]), .A2(n840), .B1(n1092), .B2(\mem[12][0] ), 
        .ZN(n1093) );
  INV_X1 U280 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U281 ( .A1(data_in[1]), .A2(n840), .B1(n1092), .B2(\mem[12][1] ), 
        .ZN(n1091) );
  INV_X1 U282 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U283 ( .A1(data_in[2]), .A2(n840), .B1(n1092), .B2(\mem[12][2] ), 
        .ZN(n1090) );
  INV_X1 U284 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U285 ( .A1(data_in[3]), .A2(n840), .B1(n1092), .B2(\mem[12][3] ), 
        .ZN(n1089) );
  INV_X1 U286 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U287 ( .A1(data_in[4]), .A2(n840), .B1(n1092), .B2(\mem[12][4] ), 
        .ZN(n1088) );
  INV_X1 U288 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U289 ( .A1(data_in[5]), .A2(n840), .B1(n1092), .B2(\mem[12][5] ), 
        .ZN(n1087) );
  INV_X1 U290 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U291 ( .A1(data_in[6]), .A2(n840), .B1(n1092), .B2(\mem[12][6] ), 
        .ZN(n1086) );
  INV_X1 U292 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U293 ( .A1(data_in[7]), .A2(n840), .B1(n1092), .B2(\mem[12][7] ), 
        .ZN(n1085) );
  INV_X1 U294 ( .A(n1084), .ZN(n780) );
  AOI22_X1 U295 ( .A1(data_in[0]), .A2(n839), .B1(n1083), .B2(\mem[13][0] ), 
        .ZN(n1084) );
  INV_X1 U296 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U297 ( .A1(data_in[1]), .A2(n839), .B1(n1083), .B2(\mem[13][1] ), 
        .ZN(n1082) );
  INV_X1 U298 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U299 ( .A1(data_in[2]), .A2(n839), .B1(n1083), .B2(\mem[13][2] ), 
        .ZN(n1081) );
  INV_X1 U300 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U301 ( .A1(data_in[3]), .A2(n839), .B1(n1083), .B2(\mem[13][3] ), 
        .ZN(n1080) );
  INV_X1 U302 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U303 ( .A1(data_in[4]), .A2(n839), .B1(n1083), .B2(\mem[13][4] ), 
        .ZN(n1079) );
  INV_X1 U304 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U305 ( .A1(data_in[5]), .A2(n839), .B1(n1083), .B2(\mem[13][5] ), 
        .ZN(n1078) );
  INV_X1 U306 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U307 ( .A1(data_in[6]), .A2(n839), .B1(n1083), .B2(\mem[13][6] ), 
        .ZN(n1077) );
  INV_X1 U308 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U309 ( .A1(data_in[7]), .A2(n839), .B1(n1083), .B2(\mem[13][7] ), 
        .ZN(n1076) );
  INV_X1 U310 ( .A(n1075), .ZN(n772) );
  AOI22_X1 U311 ( .A1(data_in[0]), .A2(n838), .B1(n1074), .B2(\mem[14][0] ), 
        .ZN(n1075) );
  INV_X1 U312 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U313 ( .A1(data_in[1]), .A2(n838), .B1(n1074), .B2(\mem[14][1] ), 
        .ZN(n1073) );
  INV_X1 U314 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U315 ( .A1(data_in[2]), .A2(n838), .B1(n1074), .B2(\mem[14][2] ), 
        .ZN(n1072) );
  INV_X1 U316 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U317 ( .A1(data_in[3]), .A2(n838), .B1(n1074), .B2(\mem[14][3] ), 
        .ZN(n1071) );
  INV_X1 U318 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U319 ( .A1(data_in[4]), .A2(n838), .B1(n1074), .B2(\mem[14][4] ), 
        .ZN(n1070) );
  INV_X1 U320 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U321 ( .A1(data_in[5]), .A2(n838), .B1(n1074), .B2(\mem[14][5] ), 
        .ZN(n1069) );
  INV_X1 U322 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U323 ( .A1(data_in[6]), .A2(n838), .B1(n1074), .B2(\mem[14][6] ), 
        .ZN(n1068) );
  INV_X1 U324 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U325 ( .A1(data_in[7]), .A2(n838), .B1(n1074), .B2(\mem[14][7] ), 
        .ZN(n1067) );
  INV_X1 U326 ( .A(n1066), .ZN(n764) );
  AOI22_X1 U327 ( .A1(data_in[0]), .A2(n837), .B1(n1065), .B2(\mem[15][0] ), 
        .ZN(n1066) );
  INV_X1 U328 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U329 ( .A1(data_in[1]), .A2(n837), .B1(n1065), .B2(\mem[15][1] ), 
        .ZN(n1064) );
  INV_X1 U330 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U331 ( .A1(data_in[2]), .A2(n837), .B1(n1065), .B2(\mem[15][2] ), 
        .ZN(n1063) );
  INV_X1 U332 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U333 ( .A1(data_in[3]), .A2(n837), .B1(n1065), .B2(\mem[15][3] ), 
        .ZN(n1062) );
  INV_X1 U334 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U335 ( .A1(data_in[4]), .A2(n837), .B1(n1065), .B2(\mem[15][4] ), 
        .ZN(n1061) );
  INV_X1 U336 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U337 ( .A1(data_in[5]), .A2(n837), .B1(n1065), .B2(\mem[15][5] ), 
        .ZN(n1060) );
  INV_X1 U338 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U339 ( .A1(data_in[6]), .A2(n837), .B1(n1065), .B2(\mem[15][6] ), 
        .ZN(n1059) );
  INV_X1 U340 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U341 ( .A1(data_in[7]), .A2(n837), .B1(n1065), .B2(\mem[15][7] ), 
        .ZN(n1058) );
  INV_X1 U342 ( .A(n1057), .ZN(n756) );
  AOI22_X1 U343 ( .A1(data_in[0]), .A2(n836), .B1(n1056), .B2(\mem[16][0] ), 
        .ZN(n1057) );
  INV_X1 U344 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U345 ( .A1(data_in[1]), .A2(n836), .B1(n1056), .B2(\mem[16][1] ), 
        .ZN(n1055) );
  INV_X1 U346 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U347 ( .A1(data_in[2]), .A2(n836), .B1(n1056), .B2(\mem[16][2] ), 
        .ZN(n1054) );
  INV_X1 U348 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U349 ( .A1(data_in[3]), .A2(n836), .B1(n1056), .B2(\mem[16][3] ), 
        .ZN(n1053) );
  INV_X1 U350 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U351 ( .A1(data_in[4]), .A2(n836), .B1(n1056), .B2(\mem[16][4] ), 
        .ZN(n1052) );
  INV_X1 U352 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U353 ( .A1(data_in[5]), .A2(n836), .B1(n1056), .B2(\mem[16][5] ), 
        .ZN(n1051) );
  INV_X1 U354 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U355 ( .A1(data_in[6]), .A2(n836), .B1(n1056), .B2(\mem[16][6] ), 
        .ZN(n1050) );
  INV_X1 U356 ( .A(n1049), .ZN(n749) );
  AOI22_X1 U357 ( .A1(data_in[7]), .A2(n836), .B1(n1056), .B2(\mem[16][7] ), 
        .ZN(n1049) );
  INV_X1 U358 ( .A(n1047), .ZN(n748) );
  AOI22_X1 U359 ( .A1(data_in[0]), .A2(n835), .B1(n1046), .B2(\mem[17][0] ), 
        .ZN(n1047) );
  INV_X1 U360 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U361 ( .A1(data_in[1]), .A2(n835), .B1(n1046), .B2(\mem[17][1] ), 
        .ZN(n1045) );
  INV_X1 U362 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U363 ( .A1(data_in[2]), .A2(n835), .B1(n1046), .B2(\mem[17][2] ), 
        .ZN(n1044) );
  INV_X1 U364 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[3]), .A2(n835), .B1(n1046), .B2(\mem[17][3] ), 
        .ZN(n1043) );
  INV_X1 U366 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[4]), .A2(n835), .B1(n1046), .B2(\mem[17][4] ), 
        .ZN(n1042) );
  INV_X1 U368 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[5]), .A2(n835), .B1(n1046), .B2(\mem[17][5] ), 
        .ZN(n1041) );
  INV_X1 U370 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[6]), .A2(n835), .B1(n1046), .B2(\mem[17][6] ), 
        .ZN(n1040) );
  INV_X1 U372 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[7]), .A2(n835), .B1(n1046), .B2(\mem[17][7] ), 
        .ZN(n1039) );
  INV_X1 U374 ( .A(n1038), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[0]), .A2(n834), .B1(n1037), .B2(\mem[18][0] ), 
        .ZN(n1038) );
  INV_X1 U376 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[1]), .A2(n834), .B1(n1037), .B2(\mem[18][1] ), 
        .ZN(n1036) );
  INV_X1 U378 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[2]), .A2(n834), .B1(n1037), .B2(\mem[18][2] ), 
        .ZN(n1035) );
  INV_X1 U380 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U381 ( .A1(data_in[3]), .A2(n834), .B1(n1037), .B2(\mem[18][3] ), 
        .ZN(n1034) );
  INV_X1 U382 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U383 ( .A1(data_in[4]), .A2(n834), .B1(n1037), .B2(\mem[18][4] ), 
        .ZN(n1033) );
  INV_X1 U384 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U385 ( .A1(data_in[5]), .A2(n834), .B1(n1037), .B2(\mem[18][5] ), 
        .ZN(n1032) );
  INV_X1 U386 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U387 ( .A1(data_in[6]), .A2(n834), .B1(n1037), .B2(\mem[18][6] ), 
        .ZN(n1031) );
  INV_X1 U388 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U389 ( .A1(data_in[7]), .A2(n834), .B1(n1037), .B2(\mem[18][7] ), 
        .ZN(n1030) );
  INV_X1 U390 ( .A(n1029), .ZN(n732) );
  AOI22_X1 U391 ( .A1(data_in[0]), .A2(n833), .B1(n1028), .B2(\mem[19][0] ), 
        .ZN(n1029) );
  INV_X1 U392 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U393 ( .A1(data_in[1]), .A2(n833), .B1(n1028), .B2(\mem[19][1] ), 
        .ZN(n1027) );
  INV_X1 U394 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U395 ( .A1(data_in[2]), .A2(n833), .B1(n1028), .B2(\mem[19][2] ), 
        .ZN(n1026) );
  INV_X1 U396 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U397 ( .A1(data_in[3]), .A2(n833), .B1(n1028), .B2(\mem[19][3] ), 
        .ZN(n1025) );
  INV_X1 U398 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U399 ( .A1(data_in[4]), .A2(n833), .B1(n1028), .B2(\mem[19][4] ), 
        .ZN(n1024) );
  INV_X1 U400 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U401 ( .A1(data_in[5]), .A2(n833), .B1(n1028), .B2(\mem[19][5] ), 
        .ZN(n1023) );
  INV_X1 U402 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U403 ( .A1(data_in[6]), .A2(n833), .B1(n1028), .B2(\mem[19][6] ), 
        .ZN(n1022) );
  INV_X1 U404 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U405 ( .A1(data_in[7]), .A2(n833), .B1(n1028), .B2(\mem[19][7] ), 
        .ZN(n1021) );
  INV_X1 U406 ( .A(n1020), .ZN(n724) );
  AOI22_X1 U407 ( .A1(data_in[0]), .A2(n832), .B1(n1019), .B2(\mem[20][0] ), 
        .ZN(n1020) );
  INV_X1 U408 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U409 ( .A1(data_in[1]), .A2(n832), .B1(n1019), .B2(\mem[20][1] ), 
        .ZN(n1018) );
  INV_X1 U410 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U411 ( .A1(data_in[2]), .A2(n832), .B1(n1019), .B2(\mem[20][2] ), 
        .ZN(n1017) );
  INV_X1 U412 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U413 ( .A1(data_in[3]), .A2(n832), .B1(n1019), .B2(\mem[20][3] ), 
        .ZN(n1016) );
  INV_X1 U414 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U415 ( .A1(data_in[4]), .A2(n832), .B1(n1019), .B2(\mem[20][4] ), 
        .ZN(n1015) );
  INV_X1 U416 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U417 ( .A1(data_in[5]), .A2(n832), .B1(n1019), .B2(\mem[20][5] ), 
        .ZN(n1014) );
  INV_X1 U418 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U419 ( .A1(data_in[6]), .A2(n832), .B1(n1019), .B2(\mem[20][6] ), 
        .ZN(n1013) );
  INV_X1 U420 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U421 ( .A1(data_in[7]), .A2(n832), .B1(n1019), .B2(\mem[20][7] ), 
        .ZN(n1012) );
  INV_X1 U422 ( .A(n1011), .ZN(n716) );
  AOI22_X1 U423 ( .A1(data_in[0]), .A2(n831), .B1(n1010), .B2(\mem[21][0] ), 
        .ZN(n1011) );
  INV_X1 U424 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U425 ( .A1(data_in[1]), .A2(n831), .B1(n1010), .B2(\mem[21][1] ), 
        .ZN(n1009) );
  INV_X1 U426 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U427 ( .A1(data_in[2]), .A2(n831), .B1(n1010), .B2(\mem[21][2] ), 
        .ZN(n1008) );
  INV_X1 U428 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U429 ( .A1(data_in[3]), .A2(n831), .B1(n1010), .B2(\mem[21][3] ), 
        .ZN(n1007) );
  INV_X1 U430 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U431 ( .A1(data_in[4]), .A2(n831), .B1(n1010), .B2(\mem[21][4] ), 
        .ZN(n1006) );
  INV_X1 U432 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U433 ( .A1(data_in[5]), .A2(n831), .B1(n1010), .B2(\mem[21][5] ), 
        .ZN(n1005) );
  INV_X1 U434 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U435 ( .A1(data_in[6]), .A2(n831), .B1(n1010), .B2(\mem[21][6] ), 
        .ZN(n1004) );
  INV_X1 U436 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U437 ( .A1(data_in[7]), .A2(n831), .B1(n1010), .B2(\mem[21][7] ), 
        .ZN(n1003) );
  INV_X1 U438 ( .A(n1002), .ZN(n708) );
  AOI22_X1 U439 ( .A1(data_in[0]), .A2(n830), .B1(n1001), .B2(\mem[22][0] ), 
        .ZN(n1002) );
  INV_X1 U440 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U441 ( .A1(data_in[1]), .A2(n830), .B1(n1001), .B2(\mem[22][1] ), 
        .ZN(n1000) );
  INV_X1 U442 ( .A(n999), .ZN(n706) );
  AOI22_X1 U443 ( .A1(data_in[2]), .A2(n830), .B1(n1001), .B2(\mem[22][2] ), 
        .ZN(n999) );
  INV_X1 U444 ( .A(n998), .ZN(n705) );
  AOI22_X1 U445 ( .A1(data_in[3]), .A2(n830), .B1(n1001), .B2(\mem[22][3] ), 
        .ZN(n998) );
  INV_X1 U446 ( .A(n997), .ZN(n704) );
  AOI22_X1 U447 ( .A1(data_in[4]), .A2(n830), .B1(n1001), .B2(\mem[22][4] ), 
        .ZN(n997) );
  INV_X1 U448 ( .A(n996), .ZN(n703) );
  AOI22_X1 U449 ( .A1(data_in[5]), .A2(n830), .B1(n1001), .B2(\mem[22][5] ), 
        .ZN(n996) );
  INV_X1 U450 ( .A(n995), .ZN(n702) );
  AOI22_X1 U451 ( .A1(data_in[6]), .A2(n830), .B1(n1001), .B2(\mem[22][6] ), 
        .ZN(n995) );
  INV_X1 U452 ( .A(n994), .ZN(n701) );
  AOI22_X1 U453 ( .A1(data_in[7]), .A2(n830), .B1(n1001), .B2(\mem[22][7] ), 
        .ZN(n994) );
  INV_X1 U454 ( .A(n993), .ZN(n700) );
  AOI22_X1 U455 ( .A1(data_in[0]), .A2(n829), .B1(n992), .B2(\mem[23][0] ), 
        .ZN(n993) );
  INV_X1 U456 ( .A(n991), .ZN(n699) );
  AOI22_X1 U457 ( .A1(data_in[1]), .A2(n829), .B1(n992), .B2(\mem[23][1] ), 
        .ZN(n991) );
  INV_X1 U458 ( .A(n990), .ZN(n698) );
  AOI22_X1 U459 ( .A1(data_in[2]), .A2(n829), .B1(n992), .B2(\mem[23][2] ), 
        .ZN(n990) );
  INV_X1 U460 ( .A(n989), .ZN(n697) );
  AOI22_X1 U461 ( .A1(data_in[3]), .A2(n829), .B1(n992), .B2(\mem[23][3] ), 
        .ZN(n989) );
  INV_X1 U462 ( .A(n988), .ZN(n696) );
  AOI22_X1 U463 ( .A1(data_in[4]), .A2(n829), .B1(n992), .B2(\mem[23][4] ), 
        .ZN(n988) );
  INV_X1 U464 ( .A(n987), .ZN(n695) );
  AOI22_X1 U465 ( .A1(data_in[5]), .A2(n829), .B1(n992), .B2(\mem[23][5] ), 
        .ZN(n987) );
  INV_X1 U466 ( .A(n986), .ZN(n694) );
  AOI22_X1 U467 ( .A1(data_in[6]), .A2(n829), .B1(n992), .B2(\mem[23][6] ), 
        .ZN(n986) );
  INV_X1 U468 ( .A(n985), .ZN(n693) );
  AOI22_X1 U469 ( .A1(data_in[7]), .A2(n829), .B1(n992), .B2(\mem[23][7] ), 
        .ZN(n985) );
  INV_X1 U470 ( .A(n984), .ZN(n692) );
  AOI22_X1 U471 ( .A1(data_in[0]), .A2(n828), .B1(n983), .B2(\mem[24][0] ), 
        .ZN(n984) );
  INV_X1 U472 ( .A(n982), .ZN(n691) );
  AOI22_X1 U473 ( .A1(data_in[1]), .A2(n828), .B1(n983), .B2(\mem[24][1] ), 
        .ZN(n982) );
  INV_X1 U474 ( .A(n981), .ZN(n690) );
  AOI22_X1 U475 ( .A1(data_in[2]), .A2(n828), .B1(n983), .B2(\mem[24][2] ), 
        .ZN(n981) );
  INV_X1 U476 ( .A(n980), .ZN(n689) );
  AOI22_X1 U477 ( .A1(data_in[3]), .A2(n828), .B1(n983), .B2(\mem[24][3] ), 
        .ZN(n980) );
  INV_X1 U478 ( .A(n979), .ZN(n688) );
  AOI22_X1 U479 ( .A1(data_in[4]), .A2(n828), .B1(n983), .B2(\mem[24][4] ), 
        .ZN(n979) );
  INV_X1 U480 ( .A(n978), .ZN(n687) );
  AOI22_X1 U481 ( .A1(data_in[5]), .A2(n828), .B1(n983), .B2(\mem[24][5] ), 
        .ZN(n978) );
  INV_X1 U482 ( .A(n977), .ZN(n686) );
  AOI22_X1 U483 ( .A1(data_in[6]), .A2(n828), .B1(n983), .B2(\mem[24][6] ), 
        .ZN(n977) );
  INV_X1 U484 ( .A(n976), .ZN(n685) );
  AOI22_X1 U485 ( .A1(data_in[7]), .A2(n828), .B1(n983), .B2(\mem[24][7] ), 
        .ZN(n976) );
  INV_X1 U486 ( .A(n974), .ZN(n684) );
  AOI22_X1 U487 ( .A1(data_in[0]), .A2(n827), .B1(n973), .B2(\mem[25][0] ), 
        .ZN(n974) );
  INV_X1 U488 ( .A(n972), .ZN(n683) );
  AOI22_X1 U489 ( .A1(data_in[1]), .A2(n827), .B1(n973), .B2(\mem[25][1] ), 
        .ZN(n972) );
  INV_X1 U490 ( .A(n971), .ZN(n682) );
  AOI22_X1 U491 ( .A1(data_in[2]), .A2(n827), .B1(n973), .B2(\mem[25][2] ), 
        .ZN(n971) );
  INV_X1 U492 ( .A(n970), .ZN(n681) );
  AOI22_X1 U493 ( .A1(data_in[3]), .A2(n827), .B1(n973), .B2(\mem[25][3] ), 
        .ZN(n970) );
  INV_X1 U494 ( .A(n969), .ZN(n680) );
  AOI22_X1 U495 ( .A1(data_in[4]), .A2(n827), .B1(n973), .B2(\mem[25][4] ), 
        .ZN(n969) );
  INV_X1 U496 ( .A(n968), .ZN(n679) );
  AOI22_X1 U497 ( .A1(data_in[5]), .A2(n827), .B1(n973), .B2(\mem[25][5] ), 
        .ZN(n968) );
  INV_X1 U498 ( .A(n967), .ZN(n678) );
  AOI22_X1 U499 ( .A1(data_in[6]), .A2(n827), .B1(n973), .B2(\mem[25][6] ), 
        .ZN(n967) );
  INV_X1 U500 ( .A(n966), .ZN(n677) );
  AOI22_X1 U501 ( .A1(data_in[7]), .A2(n827), .B1(n973), .B2(\mem[25][7] ), 
        .ZN(n966) );
  INV_X1 U502 ( .A(n965), .ZN(n676) );
  AOI22_X1 U503 ( .A1(data_in[0]), .A2(n826), .B1(n964), .B2(\mem[26][0] ), 
        .ZN(n965) );
  INV_X1 U504 ( .A(n963), .ZN(n675) );
  AOI22_X1 U505 ( .A1(data_in[1]), .A2(n826), .B1(n964), .B2(\mem[26][1] ), 
        .ZN(n963) );
  INV_X1 U506 ( .A(n962), .ZN(n674) );
  AOI22_X1 U507 ( .A1(data_in[2]), .A2(n826), .B1(n964), .B2(\mem[26][2] ), 
        .ZN(n962) );
  INV_X1 U508 ( .A(n961), .ZN(n673) );
  AOI22_X1 U509 ( .A1(data_in[3]), .A2(n826), .B1(n964), .B2(\mem[26][3] ), 
        .ZN(n961) );
  INV_X1 U510 ( .A(n960), .ZN(n672) );
  AOI22_X1 U511 ( .A1(data_in[4]), .A2(n826), .B1(n964), .B2(\mem[26][4] ), 
        .ZN(n960) );
  INV_X1 U512 ( .A(n959), .ZN(n671) );
  AOI22_X1 U513 ( .A1(data_in[5]), .A2(n826), .B1(n964), .B2(\mem[26][5] ), 
        .ZN(n959) );
  INV_X1 U514 ( .A(n958), .ZN(n670) );
  AOI22_X1 U515 ( .A1(data_in[6]), .A2(n826), .B1(n964), .B2(\mem[26][6] ), 
        .ZN(n958) );
  INV_X1 U516 ( .A(n957), .ZN(n669) );
  AOI22_X1 U517 ( .A1(data_in[7]), .A2(n826), .B1(n964), .B2(\mem[26][7] ), 
        .ZN(n957) );
  INV_X1 U518 ( .A(n956), .ZN(n668) );
  AOI22_X1 U519 ( .A1(data_in[0]), .A2(n825), .B1(n955), .B2(\mem[27][0] ), 
        .ZN(n956) );
  INV_X1 U520 ( .A(n954), .ZN(n667) );
  AOI22_X1 U521 ( .A1(data_in[1]), .A2(n825), .B1(n955), .B2(\mem[27][1] ), 
        .ZN(n954) );
  INV_X1 U522 ( .A(n953), .ZN(n666) );
  AOI22_X1 U523 ( .A1(data_in[2]), .A2(n825), .B1(n955), .B2(\mem[27][2] ), 
        .ZN(n953) );
  INV_X1 U524 ( .A(n952), .ZN(n665) );
  AOI22_X1 U525 ( .A1(data_in[3]), .A2(n825), .B1(n955), .B2(\mem[27][3] ), 
        .ZN(n952) );
  INV_X1 U526 ( .A(n951), .ZN(n664) );
  AOI22_X1 U527 ( .A1(data_in[4]), .A2(n825), .B1(n955), .B2(\mem[27][4] ), 
        .ZN(n951) );
  INV_X1 U528 ( .A(n950), .ZN(n663) );
  AOI22_X1 U529 ( .A1(data_in[5]), .A2(n825), .B1(n955), .B2(\mem[27][5] ), 
        .ZN(n950) );
  INV_X1 U530 ( .A(n949), .ZN(n662) );
  AOI22_X1 U531 ( .A1(data_in[6]), .A2(n825), .B1(n955), .B2(\mem[27][6] ), 
        .ZN(n949) );
  INV_X1 U532 ( .A(n948), .ZN(n661) );
  AOI22_X1 U533 ( .A1(data_in[7]), .A2(n825), .B1(n955), .B2(\mem[27][7] ), 
        .ZN(n948) );
  INV_X1 U534 ( .A(n947), .ZN(n660) );
  AOI22_X1 U535 ( .A1(data_in[0]), .A2(n824), .B1(n946), .B2(\mem[28][0] ), 
        .ZN(n947) );
  INV_X1 U536 ( .A(n945), .ZN(n659) );
  AOI22_X1 U537 ( .A1(data_in[1]), .A2(n824), .B1(n946), .B2(\mem[28][1] ), 
        .ZN(n945) );
  INV_X1 U538 ( .A(n944), .ZN(n658) );
  AOI22_X1 U539 ( .A1(data_in[2]), .A2(n824), .B1(n946), .B2(\mem[28][2] ), 
        .ZN(n944) );
  INV_X1 U540 ( .A(n943), .ZN(n657) );
  AOI22_X1 U541 ( .A1(data_in[3]), .A2(n824), .B1(n946), .B2(\mem[28][3] ), 
        .ZN(n943) );
  INV_X1 U542 ( .A(n942), .ZN(n656) );
  AOI22_X1 U543 ( .A1(data_in[4]), .A2(n824), .B1(n946), .B2(\mem[28][4] ), 
        .ZN(n942) );
  INV_X1 U544 ( .A(n941), .ZN(n655) );
  AOI22_X1 U545 ( .A1(data_in[5]), .A2(n824), .B1(n946), .B2(\mem[28][5] ), 
        .ZN(n941) );
  INV_X1 U546 ( .A(n940), .ZN(n654) );
  AOI22_X1 U547 ( .A1(data_in[6]), .A2(n824), .B1(n946), .B2(\mem[28][6] ), 
        .ZN(n940) );
  INV_X1 U548 ( .A(n939), .ZN(n653) );
  AOI22_X1 U549 ( .A1(data_in[7]), .A2(n824), .B1(n946), .B2(\mem[28][7] ), 
        .ZN(n939) );
  INV_X1 U550 ( .A(n938), .ZN(n652) );
  AOI22_X1 U551 ( .A1(data_in[0]), .A2(n823), .B1(n937), .B2(\mem[29][0] ), 
        .ZN(n938) );
  INV_X1 U552 ( .A(n936), .ZN(n651) );
  AOI22_X1 U553 ( .A1(data_in[1]), .A2(n823), .B1(n937), .B2(\mem[29][1] ), 
        .ZN(n936) );
  INV_X1 U554 ( .A(n935), .ZN(n650) );
  AOI22_X1 U555 ( .A1(data_in[2]), .A2(n823), .B1(n937), .B2(\mem[29][2] ), 
        .ZN(n935) );
  INV_X1 U556 ( .A(n934), .ZN(n649) );
  AOI22_X1 U557 ( .A1(data_in[3]), .A2(n823), .B1(n937), .B2(\mem[29][3] ), 
        .ZN(n934) );
  INV_X1 U558 ( .A(n933), .ZN(n648) );
  AOI22_X1 U559 ( .A1(data_in[4]), .A2(n823), .B1(n937), .B2(\mem[29][4] ), 
        .ZN(n933) );
  INV_X1 U560 ( .A(n932), .ZN(n647) );
  AOI22_X1 U561 ( .A1(data_in[5]), .A2(n823), .B1(n937), .B2(\mem[29][5] ), 
        .ZN(n932) );
  INV_X1 U562 ( .A(n931), .ZN(n646) );
  AOI22_X1 U563 ( .A1(data_in[6]), .A2(n823), .B1(n937), .B2(\mem[29][6] ), 
        .ZN(n931) );
  INV_X1 U564 ( .A(n930), .ZN(n645) );
  AOI22_X1 U565 ( .A1(data_in[7]), .A2(n823), .B1(n937), .B2(\mem[29][7] ), 
        .ZN(n930) );
  INV_X1 U566 ( .A(n929), .ZN(n644) );
  AOI22_X1 U567 ( .A1(data_in[0]), .A2(n822), .B1(n928), .B2(\mem[30][0] ), 
        .ZN(n929) );
  INV_X1 U568 ( .A(n927), .ZN(n643) );
  AOI22_X1 U569 ( .A1(data_in[1]), .A2(n822), .B1(n928), .B2(\mem[30][1] ), 
        .ZN(n927) );
  INV_X1 U570 ( .A(n926), .ZN(n642) );
  AOI22_X1 U571 ( .A1(data_in[2]), .A2(n822), .B1(n928), .B2(\mem[30][2] ), 
        .ZN(n926) );
  INV_X1 U572 ( .A(n925), .ZN(n641) );
  AOI22_X1 U573 ( .A1(data_in[3]), .A2(n822), .B1(n928), .B2(\mem[30][3] ), 
        .ZN(n925) );
  INV_X1 U574 ( .A(n924), .ZN(n640) );
  AOI22_X1 U575 ( .A1(data_in[4]), .A2(n822), .B1(n928), .B2(\mem[30][4] ), 
        .ZN(n924) );
  INV_X1 U576 ( .A(n923), .ZN(n639) );
  AOI22_X1 U577 ( .A1(data_in[5]), .A2(n822), .B1(n928), .B2(\mem[30][5] ), 
        .ZN(n923) );
  INV_X1 U578 ( .A(n922), .ZN(n638) );
  AOI22_X1 U579 ( .A1(data_in[6]), .A2(n822), .B1(n928), .B2(\mem[30][6] ), 
        .ZN(n922) );
  INV_X1 U580 ( .A(n921), .ZN(n637) );
  AOI22_X1 U581 ( .A1(data_in[7]), .A2(n822), .B1(n928), .B2(\mem[30][7] ), 
        .ZN(n921) );
  INV_X1 U582 ( .A(n920), .ZN(n636) );
  AOI22_X1 U583 ( .A1(data_in[0]), .A2(n821), .B1(n919), .B2(\mem[31][0] ), 
        .ZN(n920) );
  INV_X1 U584 ( .A(n918), .ZN(n635) );
  AOI22_X1 U585 ( .A1(data_in[1]), .A2(n821), .B1(n919), .B2(\mem[31][1] ), 
        .ZN(n918) );
  INV_X1 U586 ( .A(n917), .ZN(n634) );
  AOI22_X1 U587 ( .A1(data_in[2]), .A2(n821), .B1(n919), .B2(\mem[31][2] ), 
        .ZN(n917) );
  INV_X1 U588 ( .A(n916), .ZN(n633) );
  AOI22_X1 U589 ( .A1(data_in[3]), .A2(n821), .B1(n919), .B2(\mem[31][3] ), 
        .ZN(n916) );
  INV_X1 U590 ( .A(n915), .ZN(n632) );
  AOI22_X1 U591 ( .A1(data_in[4]), .A2(n821), .B1(n919), .B2(\mem[31][4] ), 
        .ZN(n915) );
  INV_X1 U592 ( .A(n914), .ZN(n631) );
  AOI22_X1 U593 ( .A1(data_in[5]), .A2(n821), .B1(n919), .B2(\mem[31][5] ), 
        .ZN(n914) );
  INV_X1 U594 ( .A(n913), .ZN(n630) );
  AOI22_X1 U595 ( .A1(data_in[6]), .A2(n821), .B1(n919), .B2(\mem[31][6] ), 
        .ZN(n913) );
  INV_X1 U596 ( .A(n912), .ZN(n629) );
  AOI22_X1 U597 ( .A1(data_in[7]), .A2(n821), .B1(n919), .B2(\mem[31][7] ), 
        .ZN(n912) );
  MUX2_X1 U598 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n613), .Z(n3) );
  MUX2_X1 U599 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n613), .Z(n4) );
  MUX2_X1 U600 ( .A(n4), .B(n3), .S(n610), .Z(n5) );
  MUX2_X1 U601 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n613), .Z(n6) );
  MUX2_X1 U602 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n613), .Z(n7) );
  MUX2_X1 U603 ( .A(n7), .B(n6), .S(n610), .Z(n8) );
  MUX2_X1 U604 ( .A(n8), .B(n5), .S(n608), .Z(n9) );
  MUX2_X1 U605 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n613), .Z(n10) );
  MUX2_X1 U606 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n613), .Z(n11) );
  MUX2_X1 U607 ( .A(n11), .B(n10), .S(n610), .Z(n12) );
  MUX2_X1 U608 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n613), .Z(n13) );
  MUX2_X1 U609 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n613), .Z(n14) );
  MUX2_X1 U610 ( .A(n14), .B(n13), .S(n610), .Z(n15) );
  MUX2_X1 U611 ( .A(n15), .B(n12), .S(n608), .Z(n16) );
  MUX2_X1 U612 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U613 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n614), .Z(n18) );
  MUX2_X1 U614 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n614), .Z(n19) );
  MUX2_X1 U615 ( .A(n19), .B(n18), .S(n611), .Z(n20) );
  MUX2_X1 U616 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n614), .Z(n21) );
  MUX2_X1 U617 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n614), .Z(n22) );
  MUX2_X1 U618 ( .A(n22), .B(n21), .S(n611), .Z(n23) );
  MUX2_X1 U619 ( .A(n23), .B(n20), .S(n608), .Z(n24) );
  MUX2_X1 U620 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n614), .Z(n25) );
  MUX2_X1 U621 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n614), .Z(n26) );
  MUX2_X1 U622 ( .A(n26), .B(n25), .S(n611), .Z(n27) );
  MUX2_X1 U623 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n614), .Z(n28) );
  MUX2_X1 U624 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n614), .Z(n29) );
  MUX2_X1 U625 ( .A(n29), .B(n28), .S(n611), .Z(n30) );
  MUX2_X1 U626 ( .A(n30), .B(n27), .S(n608), .Z(n31) );
  MUX2_X1 U627 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U628 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U629 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n614), .Z(n33) );
  MUX2_X1 U630 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n614), .Z(n34) );
  MUX2_X1 U631 ( .A(n34), .B(n33), .S(n611), .Z(n35) );
  MUX2_X1 U632 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n614), .Z(n36) );
  MUX2_X1 U633 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n614), .Z(n37) );
  MUX2_X1 U634 ( .A(n37), .B(n36), .S(n611), .Z(n38) );
  MUX2_X1 U635 ( .A(n38), .B(n35), .S(n608), .Z(n39) );
  MUX2_X1 U636 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n615), .Z(n40) );
  MUX2_X1 U637 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n615), .Z(n41) );
  MUX2_X1 U638 ( .A(n41), .B(n40), .S(n611), .Z(n42) );
  MUX2_X1 U639 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n615), .Z(n43) );
  MUX2_X1 U640 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n615), .Z(n44) );
  MUX2_X1 U641 ( .A(n44), .B(n43), .S(n611), .Z(n45) );
  MUX2_X1 U642 ( .A(n45), .B(n42), .S(n608), .Z(n46) );
  MUX2_X1 U643 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U644 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n615), .Z(n48) );
  MUX2_X1 U645 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n615), .Z(n49) );
  MUX2_X1 U646 ( .A(n49), .B(n48), .S(n611), .Z(n50) );
  MUX2_X1 U647 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n615), .Z(n51) );
  MUX2_X1 U648 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n615), .Z(n52) );
  MUX2_X1 U649 ( .A(n52), .B(n51), .S(n611), .Z(n53) );
  MUX2_X1 U650 ( .A(n53), .B(n50), .S(n608), .Z(n54) );
  MUX2_X1 U651 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n615), .Z(n55) );
  MUX2_X1 U652 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n615), .Z(n56) );
  MUX2_X1 U653 ( .A(n56), .B(n55), .S(n611), .Z(n57) );
  MUX2_X1 U654 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n615), .Z(n58) );
  MUX2_X1 U655 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n615), .Z(n59) );
  MUX2_X1 U656 ( .A(n59), .B(n58), .S(n611), .Z(n60) );
  MUX2_X1 U657 ( .A(n60), .B(n57), .S(n608), .Z(n61) );
  MUX2_X1 U658 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U659 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U660 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n616), .Z(n63) );
  MUX2_X1 U661 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n616), .Z(n64) );
  MUX2_X1 U662 ( .A(n64), .B(n63), .S(n612), .Z(n65) );
  MUX2_X1 U663 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n616), .Z(n66) );
  MUX2_X1 U664 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n616), .Z(n67) );
  MUX2_X1 U665 ( .A(n67), .B(n66), .S(n612), .Z(n68) );
  MUX2_X1 U666 ( .A(n68), .B(n65), .S(n609), .Z(n69) );
  MUX2_X1 U667 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n616), .Z(n70) );
  MUX2_X1 U668 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n616), .Z(n71) );
  MUX2_X1 U669 ( .A(n71), .B(n70), .S(n612), .Z(n72) );
  MUX2_X1 U670 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n616), .Z(n73) );
  MUX2_X1 U671 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n616), .Z(n74) );
  MUX2_X1 U672 ( .A(n74), .B(n73), .S(n612), .Z(n75) );
  MUX2_X1 U673 ( .A(n75), .B(n72), .S(n609), .Z(n76) );
  MUX2_X1 U674 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U675 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n616), .Z(n78) );
  MUX2_X1 U676 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n616), .Z(n79) );
  MUX2_X1 U677 ( .A(n79), .B(n78), .S(n612), .Z(n80) );
  MUX2_X1 U678 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n616), .Z(n81) );
  MUX2_X1 U679 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n616), .Z(n82) );
  MUX2_X1 U680 ( .A(n82), .B(n81), .S(n612), .Z(n83) );
  MUX2_X1 U681 ( .A(n83), .B(n80), .S(n609), .Z(n84) );
  MUX2_X1 U682 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n614), .Z(n85) );
  MUX2_X1 U683 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n615), .Z(n86) );
  MUX2_X1 U684 ( .A(n86), .B(n85), .S(n612), .Z(n87) );
  MUX2_X1 U685 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n613), .Z(n88) );
  MUX2_X1 U686 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n613), .Z(n89) );
  MUX2_X1 U687 ( .A(n89), .B(n88), .S(n612), .Z(n90) );
  MUX2_X1 U688 ( .A(n90), .B(n87), .S(n609), .Z(n91) );
  MUX2_X1 U689 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U690 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U691 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n616), .Z(n93) );
  MUX2_X1 U692 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n615), .Z(n94) );
  MUX2_X1 U693 ( .A(n94), .B(n93), .S(n612), .Z(n95) );
  MUX2_X1 U694 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n614), .Z(n96) );
  MUX2_X1 U695 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n615), .Z(n97) );
  MUX2_X1 U696 ( .A(n97), .B(n96), .S(n612), .Z(n98) );
  MUX2_X1 U697 ( .A(n98), .B(n95), .S(n609), .Z(n99) );
  MUX2_X1 U698 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n613), .Z(n100) );
  MUX2_X1 U699 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n616), .Z(n101) );
  MUX2_X1 U700 ( .A(n101), .B(n100), .S(n612), .Z(n102) );
  MUX2_X1 U701 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n613), .Z(n103) );
  MUX2_X1 U702 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n616), .Z(n104) );
  MUX2_X1 U703 ( .A(n104), .B(n103), .S(n612), .Z(n105) );
  MUX2_X1 U704 ( .A(n105), .B(n102), .S(n609), .Z(n106) );
  MUX2_X1 U705 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U706 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n615), .Z(n108) );
  MUX2_X1 U707 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n618), .Z(n109) );
  MUX2_X1 U708 ( .A(n109), .B(n108), .S(n611), .Z(n110) );
  MUX2_X1 U709 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n617), .Z(n111) );
  MUX2_X1 U710 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n617), .Z(n112) );
  MUX2_X1 U711 ( .A(n112), .B(n111), .S(n611), .Z(n113) );
  MUX2_X1 U712 ( .A(n113), .B(n110), .S(n609), .Z(n114) );
  MUX2_X1 U713 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n618), .Z(n115) );
  MUX2_X1 U714 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n618), .Z(n116) );
  MUX2_X1 U715 ( .A(n116), .B(n115), .S(n612), .Z(n117) );
  MUX2_X1 U716 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n614), .Z(n118) );
  MUX2_X1 U717 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n616), .Z(n119) );
  MUX2_X1 U718 ( .A(n119), .B(n118), .S(n610), .Z(n120) );
  MUX2_X1 U719 ( .A(n120), .B(n117), .S(n609), .Z(n121) );
  MUX2_X1 U720 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U721 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U722 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n618), .Z(n123) );
  MUX2_X1 U723 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n618), .Z(n124) );
  MUX2_X1 U724 ( .A(n124), .B(n123), .S(n610), .Z(n125) );
  MUX2_X1 U725 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n615), .Z(n126) );
  MUX2_X1 U726 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n617), .Z(n127) );
  MUX2_X1 U727 ( .A(n127), .B(n126), .S(n611), .Z(n128) );
  MUX2_X1 U728 ( .A(n128), .B(n125), .S(n609), .Z(n129) );
  MUX2_X1 U729 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n618), .Z(n130) );
  MUX2_X1 U730 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n617), .Z(n131) );
  MUX2_X1 U731 ( .A(n131), .B(n130), .S(n610), .Z(n132) );
  MUX2_X1 U732 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n617), .Z(n133) );
  MUX2_X1 U733 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n618), .Z(n134) );
  MUX2_X1 U734 ( .A(n134), .B(n133), .S(n610), .Z(n135) );
  MUX2_X1 U735 ( .A(n135), .B(n132), .S(n609), .Z(n136) );
  MUX2_X1 U736 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U737 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n618), .Z(n138) );
  MUX2_X1 U738 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n618), .Z(n139) );
  MUX2_X1 U739 ( .A(n139), .B(n138), .S(n612), .Z(n140) );
  MUX2_X1 U740 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n617), .Z(n141) );
  MUX2_X1 U741 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n618), .Z(n142) );
  MUX2_X1 U742 ( .A(n142), .B(n141), .S(n612), .Z(n143) );
  MUX2_X1 U743 ( .A(n143), .B(n140), .S(n609), .Z(n144) );
  MUX2_X1 U744 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n618), .Z(n145) );
  MUX2_X1 U745 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n617), .Z(n146) );
  MUX2_X1 U746 ( .A(n146), .B(n145), .S(n610), .Z(n147) );
  MUX2_X1 U747 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n617), .Z(n148) );
  MUX2_X1 U748 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n617), .Z(n149) );
  MUX2_X1 U749 ( .A(n149), .B(n148), .S(n611), .Z(n150) );
  MUX2_X1 U750 ( .A(n150), .B(n147), .S(n609), .Z(n151) );
  MUX2_X1 U751 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U752 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U753 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n613), .Z(n153) );
  MUX2_X1 U754 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n617), .Z(n154) );
  MUX2_X1 U755 ( .A(n154), .B(n153), .S(n611), .Z(n155) );
  MUX2_X1 U756 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n618), .Z(n156) );
  MUX2_X1 U757 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(N10), .Z(n157) );
  MUX2_X1 U758 ( .A(n157), .B(n156), .S(n611), .Z(n158) );
  MUX2_X1 U759 ( .A(n158), .B(n155), .S(n608), .Z(n159) );
  MUX2_X1 U760 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n617), .Z(n160) );
  MUX2_X1 U761 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(N10), .Z(n161) );
  MUX2_X1 U762 ( .A(n161), .B(n160), .S(N11), .Z(n162) );
  MUX2_X1 U763 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(N10), .Z(n163) );
  MUX2_X1 U764 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(N10), .Z(n164) );
  MUX2_X1 U765 ( .A(n164), .B(n163), .S(N11), .Z(n165) );
  MUX2_X1 U766 ( .A(n165), .B(n162), .S(N12), .Z(n166) );
  MUX2_X1 U767 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U768 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n613), .Z(n168) );
  MUX2_X1 U769 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n613), .Z(n169) );
  MUX2_X1 U770 ( .A(n169), .B(n168), .S(n610), .Z(n170) );
  MUX2_X1 U771 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n618), .Z(n171) );
  MUX2_X1 U772 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(N10), .Z(n172) );
  MUX2_X1 U773 ( .A(n172), .B(n171), .S(N11), .Z(n173) );
  MUX2_X1 U774 ( .A(n173), .B(n170), .S(n608), .Z(n174) );
  MUX2_X1 U775 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n613), .Z(n175) );
  MUX2_X1 U776 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n614), .Z(n176) );
  MUX2_X1 U777 ( .A(n176), .B(n175), .S(n612), .Z(n177) );
  MUX2_X1 U778 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n616), .Z(n178) );
  MUX2_X1 U779 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n613), .Z(n179) );
  MUX2_X1 U780 ( .A(n179), .B(n178), .S(n612), .Z(n180) );
  MUX2_X1 U781 ( .A(n180), .B(n177), .S(n609), .Z(n181) );
  MUX2_X1 U782 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U783 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U784 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n616), .Z(n183) );
  MUX2_X1 U785 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n615), .Z(n184) );
  MUX2_X1 U786 ( .A(n184), .B(n183), .S(n612), .Z(n185) );
  MUX2_X1 U787 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n614), .Z(n186) );
  MUX2_X1 U788 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n616), .Z(n187) );
  MUX2_X1 U789 ( .A(n187), .B(n186), .S(N11), .Z(n188) );
  MUX2_X1 U790 ( .A(n188), .B(n185), .S(n608), .Z(n189) );
  MUX2_X1 U791 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n613), .Z(n190) );
  MUX2_X1 U792 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n616), .Z(n191) );
  MUX2_X1 U793 ( .A(n191), .B(n190), .S(N11), .Z(n192) );
  MUX2_X1 U794 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n614), .Z(n193) );
  MUX2_X1 U795 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n614), .Z(n194) );
  MUX2_X1 U796 ( .A(n194), .B(n193), .S(n611), .Z(n195) );
  MUX2_X1 U797 ( .A(n195), .B(n192), .S(N12), .Z(n196) );
  MUX2_X1 U798 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U799 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n617), .Z(n198) );
  MUX2_X1 U800 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n617), .Z(n199) );
  MUX2_X1 U801 ( .A(n199), .B(n198), .S(n610), .Z(n200) );
  MUX2_X1 U802 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n617), .Z(n201) );
  MUX2_X1 U803 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n615), .Z(n202) );
  MUX2_X1 U804 ( .A(n202), .B(n201), .S(n611), .Z(n203) );
  MUX2_X1 U805 ( .A(n203), .B(n200), .S(n608), .Z(n204) );
  MUX2_X1 U806 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n617), .Z(n205) );
  MUX2_X1 U807 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n618), .Z(n206) );
  MUX2_X1 U808 ( .A(n206), .B(n205), .S(n610), .Z(n207) );
  MUX2_X1 U809 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n615), .Z(n208) );
  MUX2_X1 U810 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n614), .Z(n209) );
  MUX2_X1 U811 ( .A(n209), .B(n208), .S(n611), .Z(n210) );
  MUX2_X1 U812 ( .A(n210), .B(n207), .S(n609), .Z(n211) );
  MUX2_X1 U813 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U814 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U815 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n618), .Z(n213) );
  MUX2_X1 U816 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n618), .Z(n214) );
  MUX2_X1 U817 ( .A(n214), .B(n213), .S(n610), .Z(n215) );
  MUX2_X1 U818 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n613), .Z(n216) );
  MUX2_X1 U819 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n618), .Z(n217) );
  MUX2_X1 U820 ( .A(n217), .B(n216), .S(n610), .Z(n218) );
  MUX2_X1 U821 ( .A(n218), .B(n215), .S(n608), .Z(n219) );
  MUX2_X1 U822 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n618), .Z(n220) );
  MUX2_X1 U823 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n618), .Z(n221) );
  MUX2_X1 U824 ( .A(n221), .B(n220), .S(n610), .Z(n222) );
  MUX2_X1 U825 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n617), .Z(n223) );
  MUX2_X1 U826 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n617), .Z(n224) );
  MUX2_X1 U827 ( .A(n224), .B(n223), .S(n612), .Z(n225) );
  MUX2_X1 U828 ( .A(n225), .B(n222), .S(N12), .Z(n226) );
  MUX2_X1 U829 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U830 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n618), .Z(n228) );
  MUX2_X1 U831 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n617), .Z(n229) );
  MUX2_X1 U832 ( .A(n229), .B(n228), .S(n610), .Z(n595) );
  MUX2_X1 U833 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n618), .Z(n596) );
  MUX2_X1 U834 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n618), .Z(n597) );
  MUX2_X1 U835 ( .A(n597), .B(n596), .S(n612), .Z(n598) );
  MUX2_X1 U836 ( .A(n598), .B(n595), .S(n609), .Z(n599) );
  MUX2_X1 U837 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n613), .Z(n600) );
  MUX2_X1 U838 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n618), .Z(n601) );
  MUX2_X1 U839 ( .A(n601), .B(n600), .S(n610), .Z(n602) );
  MUX2_X1 U840 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n617), .Z(n603) );
  MUX2_X1 U841 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n617), .Z(n604) );
  MUX2_X1 U842 ( .A(n604), .B(n603), .S(n610), .Z(n605) );
  MUX2_X1 U843 ( .A(n605), .B(n602), .S(n608), .Z(n606) );
  MUX2_X1 U844 ( .A(n606), .B(n599), .S(N13), .Z(n607) );
  MUX2_X1 U845 ( .A(n607), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U846 ( .A(N11), .Z(n610) );
  INV_X1 U847 ( .A(N10), .ZN(n619) );
  INV_X1 U848 ( .A(N11), .ZN(n620) );
  INV_X1 U849 ( .A(data_in[0]), .ZN(n621) );
  INV_X1 U850 ( .A(data_in[1]), .ZN(n622) );
  INV_X1 U851 ( .A(data_in[2]), .ZN(n623) );
  INV_X1 U852 ( .A(data_in[3]), .ZN(n624) );
  INV_X1 U853 ( .A(data_in[4]), .ZN(n625) );
  INV_X1 U854 ( .A(data_in[5]), .ZN(n626) );
  INV_X1 U855 ( .A(data_in[6]), .ZN(n627) );
  INV_X1 U856 ( .A(data_in[7]), .ZN(n628) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_30 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n630), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n631), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n632), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n633), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n634), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n635), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n636), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n637), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n638), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n639), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n640), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n641), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n642), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n643), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n644), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n645), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n646), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n647), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n648), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n649), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n650), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n651), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n652), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n653), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n654), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n655), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n656), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n657), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n658), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n659), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n660), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n661), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n662), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n663), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n664), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n665), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n666), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n667), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n668), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n669), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n670), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n671), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n672), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n673), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n674), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n675), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n676), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n677), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n678), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n679), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n680), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n681), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n682), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n683), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n684), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n685), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n686), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n687), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n688), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n689), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n690), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n691), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n692), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n693), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n694), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n695), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n696), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n697), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n698), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n699), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n700), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n701), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n702), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n703), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n704), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n705), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n706), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n707), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n708), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n709), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n710), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n711), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n712), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n713), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n714), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n715), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n716), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n717), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n718), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n719), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n720), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n721), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n722), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n723), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n724), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n725), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n726), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n727), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n728), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n729), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n730), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n731), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n732), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n733), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n734), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n735), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n736), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n737), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n738), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n739), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n740), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n741), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n742), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n743), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n744), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n745), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n746), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n747), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n748), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n749), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n750), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n751), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n752), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n753), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n754), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n755), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n756), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n757), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n758), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n759), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n760), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n761), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n762), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n763), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n764), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n765), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n766), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n767), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n768), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n769), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n770), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n771), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n772), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n773), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n774), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n775), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n776), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n777), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n778), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n779), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n780), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n781), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n782), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n783), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n784), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n785), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n786), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n787), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n788), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n789), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n790), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n791), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n792), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n793), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n794), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n795), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n796), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n797), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n798), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n799), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n800), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n801), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n802), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n803), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n804), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n805), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n806), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n807), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n808), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n809), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n810), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n811), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n812), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n813), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n814), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n815), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n816), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n817), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n818), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n819), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n820), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n821), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n849), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n850), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n851), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n852), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n853), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n854), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n855), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n856), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n857), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n858), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n859), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n860), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n861), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n862), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n863), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n864), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n865), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n866), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n867), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n868), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n869), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n870), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n871), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n872), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n873), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n874), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n875), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n876), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n877), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n878), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n879), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n880), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n881), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n882), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n883), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n884), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n885), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n886), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n887), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n888), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n889), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n890), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n891), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n892), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n893), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n894), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n895), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n896), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n897), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n898), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n899), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n900), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n901), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n902), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n903), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n904), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n905), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n906), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n907), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n908), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n909), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n910), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n911), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n912), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n619), .Z(n611) );
  CLKBUF_X1 U4 ( .A(N11), .Z(n610) );
  BUF_X1 U5 ( .A(n619), .Z(n616) );
  BUF_X1 U6 ( .A(n619), .Z(n617) );
  BUF_X1 U7 ( .A(n619), .Z(n618) );
  BUF_X1 U8 ( .A(n619), .Z(n614) );
  BUF_X1 U9 ( .A(n619), .Z(n615) );
  BUF_X1 U10 ( .A(n619), .Z(n612) );
  BUF_X1 U11 ( .A(n619), .Z(n613) );
  BUF_X1 U12 ( .A(N11), .Z(n609) );
  BUF_X1 U13 ( .A(N10), .Z(n619) );
  NOR3_X1 U14 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1204) );
  NOR3_X1 U15 ( .A1(N11), .A2(N12), .A3(n620), .ZN(n1193) );
  NOR3_X1 U16 ( .A1(N10), .A2(N12), .A3(n621), .ZN(n1183) );
  NOR3_X1 U17 ( .A1(n620), .A2(N12), .A3(n621), .ZN(n1173) );
  INV_X1 U18 ( .A(n1130), .ZN(n845) );
  INV_X1 U19 ( .A(n1120), .ZN(n844) );
  INV_X1 U20 ( .A(n1111), .ZN(n843) );
  INV_X1 U21 ( .A(n1102), .ZN(n842) );
  INV_X1 U22 ( .A(n1057), .ZN(n837) );
  INV_X1 U23 ( .A(n1047), .ZN(n836) );
  INV_X1 U24 ( .A(n1038), .ZN(n835) );
  INV_X1 U25 ( .A(n1029), .ZN(n834) );
  INV_X1 U26 ( .A(n984), .ZN(n829) );
  INV_X1 U27 ( .A(n974), .ZN(n828) );
  INV_X1 U28 ( .A(n965), .ZN(n827) );
  INV_X1 U29 ( .A(n956), .ZN(n826) );
  INV_X1 U30 ( .A(n1093), .ZN(n841) );
  INV_X1 U31 ( .A(n1084), .ZN(n840) );
  INV_X1 U32 ( .A(n1075), .ZN(n839) );
  INV_X1 U33 ( .A(n1066), .ZN(n838) );
  INV_X1 U34 ( .A(n947), .ZN(n825) );
  INV_X1 U35 ( .A(n938), .ZN(n824) );
  INV_X1 U36 ( .A(n929), .ZN(n823) );
  INV_X1 U37 ( .A(n920), .ZN(n822) );
  INV_X1 U38 ( .A(n1020), .ZN(n833) );
  INV_X1 U39 ( .A(n1011), .ZN(n832) );
  INV_X1 U40 ( .A(n1002), .ZN(n831) );
  INV_X1 U41 ( .A(n993), .ZN(n830) );
  BUF_X1 U42 ( .A(N12), .Z(n607) );
  INV_X1 U43 ( .A(N13), .ZN(n847) );
  AND3_X1 U44 ( .A1(n620), .A2(n621), .A3(N12), .ZN(n1163) );
  AND3_X1 U45 ( .A1(N10), .A2(n621), .A3(N12), .ZN(n1153) );
  AND3_X1 U46 ( .A1(N11), .A2(n620), .A3(N12), .ZN(n1143) );
  AND3_X1 U47 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1133) );
  BUF_X1 U48 ( .A(N12), .Z(n606) );
  INV_X1 U49 ( .A(N14), .ZN(n848) );
  NAND2_X1 U50 ( .A1(n1193), .A2(n1203), .ZN(n1202) );
  NAND2_X1 U51 ( .A1(n1183), .A2(n1203), .ZN(n1192) );
  NAND2_X1 U52 ( .A1(n1173), .A2(n1203), .ZN(n1182) );
  NAND2_X1 U53 ( .A1(n1163), .A2(n1203), .ZN(n1172) );
  NAND2_X1 U54 ( .A1(n1153), .A2(n1203), .ZN(n1162) );
  NAND2_X1 U55 ( .A1(n1143), .A2(n1203), .ZN(n1152) );
  NAND2_X1 U56 ( .A1(n1133), .A2(n1203), .ZN(n1142) );
  NAND2_X1 U57 ( .A1(n1204), .A2(n1203), .ZN(n1213) );
  NAND2_X1 U58 ( .A1(n1122), .A2(n1204), .ZN(n1130) );
  NAND2_X1 U59 ( .A1(n1122), .A2(n1193), .ZN(n1120) );
  NAND2_X1 U60 ( .A1(n1122), .A2(n1183), .ZN(n1111) );
  NAND2_X1 U61 ( .A1(n1122), .A2(n1173), .ZN(n1102) );
  NAND2_X1 U62 ( .A1(n1049), .A2(n1204), .ZN(n1057) );
  NAND2_X1 U63 ( .A1(n1049), .A2(n1193), .ZN(n1047) );
  NAND2_X1 U64 ( .A1(n1049), .A2(n1183), .ZN(n1038) );
  NAND2_X1 U65 ( .A1(n1049), .A2(n1173), .ZN(n1029) );
  NAND2_X1 U66 ( .A1(n976), .A2(n1204), .ZN(n984) );
  NAND2_X1 U67 ( .A1(n976), .A2(n1193), .ZN(n974) );
  NAND2_X1 U68 ( .A1(n976), .A2(n1183), .ZN(n965) );
  NAND2_X1 U69 ( .A1(n976), .A2(n1173), .ZN(n956) );
  NAND2_X1 U70 ( .A1(n1122), .A2(n1163), .ZN(n1093) );
  NAND2_X1 U71 ( .A1(n1122), .A2(n1153), .ZN(n1084) );
  NAND2_X1 U72 ( .A1(n1122), .A2(n1143), .ZN(n1075) );
  NAND2_X1 U73 ( .A1(n1122), .A2(n1133), .ZN(n1066) );
  NAND2_X1 U74 ( .A1(n1049), .A2(n1163), .ZN(n1020) );
  NAND2_X1 U75 ( .A1(n1049), .A2(n1153), .ZN(n1011) );
  NAND2_X1 U76 ( .A1(n1049), .A2(n1143), .ZN(n1002) );
  NAND2_X1 U77 ( .A1(n1049), .A2(n1133), .ZN(n993) );
  NAND2_X1 U78 ( .A1(n976), .A2(n1163), .ZN(n947) );
  NAND2_X1 U79 ( .A1(n976), .A2(n1153), .ZN(n938) );
  NAND2_X1 U80 ( .A1(n976), .A2(n1143), .ZN(n929) );
  NAND2_X1 U81 ( .A1(n976), .A2(n1133), .ZN(n920) );
  AND3_X1 U82 ( .A1(n847), .A2(n848), .A3(n1132), .ZN(n1203) );
  AND3_X1 U83 ( .A1(N13), .A2(n1132), .A3(N14), .ZN(n976) );
  AND3_X1 U84 ( .A1(n1132), .A2(n848), .A3(N13), .ZN(n1122) );
  AND3_X1 U85 ( .A1(n1132), .A2(n847), .A3(N14), .ZN(n1049) );
  NOR2_X1 U86 ( .A1(n846), .A2(addr[5]), .ZN(n1132) );
  INV_X1 U87 ( .A(wr_en), .ZN(n846) );
  OAI21_X1 U88 ( .B1(n622), .B2(n1172), .A(n1171), .ZN(n880) );
  NAND2_X1 U89 ( .A1(\mem[4][0] ), .A2(n1172), .ZN(n1171) );
  OAI21_X1 U90 ( .B1(n623), .B2(n1172), .A(n1170), .ZN(n879) );
  NAND2_X1 U91 ( .A1(\mem[4][1] ), .A2(n1172), .ZN(n1170) );
  OAI21_X1 U92 ( .B1(n624), .B2(n1172), .A(n1169), .ZN(n878) );
  NAND2_X1 U93 ( .A1(\mem[4][2] ), .A2(n1172), .ZN(n1169) );
  OAI21_X1 U94 ( .B1(n625), .B2(n1172), .A(n1168), .ZN(n877) );
  NAND2_X1 U95 ( .A1(\mem[4][3] ), .A2(n1172), .ZN(n1168) );
  OAI21_X1 U96 ( .B1(n626), .B2(n1172), .A(n1167), .ZN(n876) );
  NAND2_X1 U97 ( .A1(\mem[4][4] ), .A2(n1172), .ZN(n1167) );
  OAI21_X1 U98 ( .B1(n627), .B2(n1172), .A(n1166), .ZN(n875) );
  NAND2_X1 U99 ( .A1(\mem[4][5] ), .A2(n1172), .ZN(n1166) );
  OAI21_X1 U100 ( .B1(n628), .B2(n1172), .A(n1165), .ZN(n874) );
  NAND2_X1 U101 ( .A1(\mem[4][6] ), .A2(n1172), .ZN(n1165) );
  OAI21_X1 U102 ( .B1(n629), .B2(n1172), .A(n1164), .ZN(n873) );
  NAND2_X1 U103 ( .A1(\mem[4][7] ), .A2(n1172), .ZN(n1164) );
  OAI21_X1 U104 ( .B1(n622), .B2(n1152), .A(n1151), .ZN(n864) );
  NAND2_X1 U105 ( .A1(\mem[6][0] ), .A2(n1152), .ZN(n1151) );
  OAI21_X1 U106 ( .B1(n623), .B2(n1152), .A(n1150), .ZN(n863) );
  NAND2_X1 U107 ( .A1(\mem[6][1] ), .A2(n1152), .ZN(n1150) );
  OAI21_X1 U108 ( .B1(n624), .B2(n1152), .A(n1149), .ZN(n862) );
  NAND2_X1 U109 ( .A1(\mem[6][2] ), .A2(n1152), .ZN(n1149) );
  OAI21_X1 U110 ( .B1(n625), .B2(n1152), .A(n1148), .ZN(n861) );
  NAND2_X1 U111 ( .A1(\mem[6][3] ), .A2(n1152), .ZN(n1148) );
  OAI21_X1 U112 ( .B1(n626), .B2(n1152), .A(n1147), .ZN(n860) );
  NAND2_X1 U113 ( .A1(\mem[6][4] ), .A2(n1152), .ZN(n1147) );
  OAI21_X1 U114 ( .B1(n627), .B2(n1152), .A(n1146), .ZN(n859) );
  NAND2_X1 U115 ( .A1(\mem[6][5] ), .A2(n1152), .ZN(n1146) );
  OAI21_X1 U116 ( .B1(n628), .B2(n1152), .A(n1145), .ZN(n858) );
  NAND2_X1 U117 ( .A1(\mem[6][6] ), .A2(n1152), .ZN(n1145) );
  OAI21_X1 U118 ( .B1(n629), .B2(n1152), .A(n1144), .ZN(n857) );
  NAND2_X1 U119 ( .A1(\mem[6][7] ), .A2(n1152), .ZN(n1144) );
  OAI21_X1 U120 ( .B1(n622), .B2(n1142), .A(n1141), .ZN(n856) );
  NAND2_X1 U121 ( .A1(\mem[7][0] ), .A2(n1142), .ZN(n1141) );
  OAI21_X1 U122 ( .B1(n623), .B2(n1142), .A(n1140), .ZN(n855) );
  NAND2_X1 U123 ( .A1(\mem[7][1] ), .A2(n1142), .ZN(n1140) );
  OAI21_X1 U124 ( .B1(n624), .B2(n1142), .A(n1139), .ZN(n854) );
  NAND2_X1 U125 ( .A1(\mem[7][2] ), .A2(n1142), .ZN(n1139) );
  OAI21_X1 U126 ( .B1(n625), .B2(n1142), .A(n1138), .ZN(n853) );
  NAND2_X1 U127 ( .A1(\mem[7][3] ), .A2(n1142), .ZN(n1138) );
  OAI21_X1 U128 ( .B1(n626), .B2(n1142), .A(n1137), .ZN(n852) );
  NAND2_X1 U129 ( .A1(\mem[7][4] ), .A2(n1142), .ZN(n1137) );
  OAI21_X1 U130 ( .B1(n627), .B2(n1142), .A(n1136), .ZN(n851) );
  NAND2_X1 U131 ( .A1(\mem[7][5] ), .A2(n1142), .ZN(n1136) );
  OAI21_X1 U132 ( .B1(n628), .B2(n1142), .A(n1135), .ZN(n850) );
  NAND2_X1 U133 ( .A1(\mem[7][6] ), .A2(n1142), .ZN(n1135) );
  OAI21_X1 U134 ( .B1(n629), .B2(n1142), .A(n1134), .ZN(n849) );
  NAND2_X1 U135 ( .A1(\mem[7][7] ), .A2(n1142), .ZN(n1134) );
  OAI21_X1 U136 ( .B1(n622), .B2(n1202), .A(n1201), .ZN(n904) );
  NAND2_X1 U137 ( .A1(\mem[1][0] ), .A2(n1202), .ZN(n1201) );
  OAI21_X1 U138 ( .B1(n623), .B2(n1202), .A(n1200), .ZN(n903) );
  NAND2_X1 U139 ( .A1(\mem[1][1] ), .A2(n1202), .ZN(n1200) );
  OAI21_X1 U140 ( .B1(n624), .B2(n1202), .A(n1199), .ZN(n902) );
  NAND2_X1 U141 ( .A1(\mem[1][2] ), .A2(n1202), .ZN(n1199) );
  OAI21_X1 U142 ( .B1(n625), .B2(n1202), .A(n1198), .ZN(n901) );
  NAND2_X1 U143 ( .A1(\mem[1][3] ), .A2(n1202), .ZN(n1198) );
  OAI21_X1 U144 ( .B1(n626), .B2(n1202), .A(n1197), .ZN(n900) );
  NAND2_X1 U145 ( .A1(\mem[1][4] ), .A2(n1202), .ZN(n1197) );
  OAI21_X1 U146 ( .B1(n627), .B2(n1202), .A(n1196), .ZN(n899) );
  NAND2_X1 U147 ( .A1(\mem[1][5] ), .A2(n1202), .ZN(n1196) );
  OAI21_X1 U148 ( .B1(n628), .B2(n1202), .A(n1195), .ZN(n898) );
  NAND2_X1 U149 ( .A1(\mem[1][6] ), .A2(n1202), .ZN(n1195) );
  OAI21_X1 U150 ( .B1(n629), .B2(n1202), .A(n1194), .ZN(n897) );
  NAND2_X1 U151 ( .A1(\mem[1][7] ), .A2(n1202), .ZN(n1194) );
  OAI21_X1 U152 ( .B1(n622), .B2(n1192), .A(n1191), .ZN(n896) );
  NAND2_X1 U153 ( .A1(\mem[2][0] ), .A2(n1192), .ZN(n1191) );
  OAI21_X1 U154 ( .B1(n623), .B2(n1192), .A(n1190), .ZN(n895) );
  NAND2_X1 U155 ( .A1(\mem[2][1] ), .A2(n1192), .ZN(n1190) );
  OAI21_X1 U156 ( .B1(n624), .B2(n1192), .A(n1189), .ZN(n894) );
  NAND2_X1 U157 ( .A1(\mem[2][2] ), .A2(n1192), .ZN(n1189) );
  OAI21_X1 U158 ( .B1(n625), .B2(n1192), .A(n1188), .ZN(n893) );
  NAND2_X1 U159 ( .A1(\mem[2][3] ), .A2(n1192), .ZN(n1188) );
  OAI21_X1 U160 ( .B1(n626), .B2(n1192), .A(n1187), .ZN(n892) );
  NAND2_X1 U161 ( .A1(\mem[2][4] ), .A2(n1192), .ZN(n1187) );
  OAI21_X1 U162 ( .B1(n627), .B2(n1192), .A(n1186), .ZN(n891) );
  NAND2_X1 U163 ( .A1(\mem[2][5] ), .A2(n1192), .ZN(n1186) );
  OAI21_X1 U164 ( .B1(n628), .B2(n1192), .A(n1185), .ZN(n890) );
  NAND2_X1 U165 ( .A1(\mem[2][6] ), .A2(n1192), .ZN(n1185) );
  OAI21_X1 U166 ( .B1(n629), .B2(n1192), .A(n1184), .ZN(n889) );
  NAND2_X1 U167 ( .A1(\mem[2][7] ), .A2(n1192), .ZN(n1184) );
  OAI21_X1 U168 ( .B1(n622), .B2(n1182), .A(n1181), .ZN(n888) );
  NAND2_X1 U169 ( .A1(\mem[3][0] ), .A2(n1182), .ZN(n1181) );
  OAI21_X1 U170 ( .B1(n623), .B2(n1182), .A(n1180), .ZN(n887) );
  NAND2_X1 U171 ( .A1(\mem[3][1] ), .A2(n1182), .ZN(n1180) );
  OAI21_X1 U172 ( .B1(n624), .B2(n1182), .A(n1179), .ZN(n886) );
  NAND2_X1 U173 ( .A1(\mem[3][2] ), .A2(n1182), .ZN(n1179) );
  OAI21_X1 U174 ( .B1(n625), .B2(n1182), .A(n1178), .ZN(n885) );
  NAND2_X1 U175 ( .A1(\mem[3][3] ), .A2(n1182), .ZN(n1178) );
  OAI21_X1 U176 ( .B1(n626), .B2(n1182), .A(n1177), .ZN(n884) );
  NAND2_X1 U177 ( .A1(\mem[3][4] ), .A2(n1182), .ZN(n1177) );
  OAI21_X1 U178 ( .B1(n627), .B2(n1182), .A(n1176), .ZN(n883) );
  NAND2_X1 U179 ( .A1(\mem[3][5] ), .A2(n1182), .ZN(n1176) );
  OAI21_X1 U180 ( .B1(n628), .B2(n1182), .A(n1175), .ZN(n882) );
  NAND2_X1 U181 ( .A1(\mem[3][6] ), .A2(n1182), .ZN(n1175) );
  OAI21_X1 U182 ( .B1(n629), .B2(n1182), .A(n1174), .ZN(n881) );
  NAND2_X1 U183 ( .A1(\mem[3][7] ), .A2(n1182), .ZN(n1174) );
  OAI21_X1 U184 ( .B1(n622), .B2(n1162), .A(n1161), .ZN(n872) );
  NAND2_X1 U185 ( .A1(\mem[5][0] ), .A2(n1162), .ZN(n1161) );
  OAI21_X1 U186 ( .B1(n623), .B2(n1162), .A(n1160), .ZN(n871) );
  NAND2_X1 U187 ( .A1(\mem[5][1] ), .A2(n1162), .ZN(n1160) );
  OAI21_X1 U188 ( .B1(n624), .B2(n1162), .A(n1159), .ZN(n870) );
  NAND2_X1 U189 ( .A1(\mem[5][2] ), .A2(n1162), .ZN(n1159) );
  OAI21_X1 U190 ( .B1(n625), .B2(n1162), .A(n1158), .ZN(n869) );
  NAND2_X1 U191 ( .A1(\mem[5][3] ), .A2(n1162), .ZN(n1158) );
  OAI21_X1 U192 ( .B1(n626), .B2(n1162), .A(n1157), .ZN(n868) );
  NAND2_X1 U193 ( .A1(\mem[5][4] ), .A2(n1162), .ZN(n1157) );
  OAI21_X1 U194 ( .B1(n627), .B2(n1162), .A(n1156), .ZN(n867) );
  NAND2_X1 U195 ( .A1(\mem[5][5] ), .A2(n1162), .ZN(n1156) );
  OAI21_X1 U196 ( .B1(n628), .B2(n1162), .A(n1155), .ZN(n866) );
  NAND2_X1 U197 ( .A1(\mem[5][6] ), .A2(n1162), .ZN(n1155) );
  OAI21_X1 U198 ( .B1(n629), .B2(n1162), .A(n1154), .ZN(n865) );
  NAND2_X1 U199 ( .A1(\mem[5][7] ), .A2(n1162), .ZN(n1154) );
  OAI21_X1 U200 ( .B1(n1213), .B2(n622), .A(n1212), .ZN(n912) );
  NAND2_X1 U201 ( .A1(\mem[0][0] ), .A2(n1213), .ZN(n1212) );
  OAI21_X1 U202 ( .B1(n1213), .B2(n623), .A(n1211), .ZN(n911) );
  NAND2_X1 U203 ( .A1(\mem[0][1] ), .A2(n1213), .ZN(n1211) );
  OAI21_X1 U204 ( .B1(n1213), .B2(n624), .A(n1210), .ZN(n910) );
  NAND2_X1 U205 ( .A1(\mem[0][2] ), .A2(n1213), .ZN(n1210) );
  OAI21_X1 U206 ( .B1(n1213), .B2(n625), .A(n1209), .ZN(n909) );
  NAND2_X1 U207 ( .A1(\mem[0][3] ), .A2(n1213), .ZN(n1209) );
  OAI21_X1 U208 ( .B1(n1213), .B2(n626), .A(n1208), .ZN(n908) );
  NAND2_X1 U209 ( .A1(\mem[0][4] ), .A2(n1213), .ZN(n1208) );
  OAI21_X1 U210 ( .B1(n1213), .B2(n627), .A(n1207), .ZN(n907) );
  NAND2_X1 U211 ( .A1(\mem[0][5] ), .A2(n1213), .ZN(n1207) );
  OAI21_X1 U212 ( .B1(n1213), .B2(n628), .A(n1206), .ZN(n906) );
  NAND2_X1 U213 ( .A1(\mem[0][6] ), .A2(n1213), .ZN(n1206) );
  OAI21_X1 U214 ( .B1(n1213), .B2(n629), .A(n1205), .ZN(n905) );
  NAND2_X1 U215 ( .A1(\mem[0][7] ), .A2(n1213), .ZN(n1205) );
  INV_X1 U216 ( .A(n1131), .ZN(n821) );
  AOI22_X1 U217 ( .A1(data_in[0]), .A2(n845), .B1(n1130), .B2(\mem[8][0] ), 
        .ZN(n1131) );
  INV_X1 U218 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U219 ( .A1(data_in[1]), .A2(n845), .B1(n1130), .B2(\mem[8][1] ), 
        .ZN(n1129) );
  INV_X1 U220 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U221 ( .A1(data_in[2]), .A2(n845), .B1(n1130), .B2(\mem[8][2] ), 
        .ZN(n1128) );
  INV_X1 U222 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U223 ( .A1(data_in[3]), .A2(n845), .B1(n1130), .B2(\mem[8][3] ), 
        .ZN(n1127) );
  INV_X1 U224 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U225 ( .A1(data_in[4]), .A2(n845), .B1(n1130), .B2(\mem[8][4] ), 
        .ZN(n1126) );
  INV_X1 U226 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U227 ( .A1(data_in[5]), .A2(n845), .B1(n1130), .B2(\mem[8][5] ), 
        .ZN(n1125) );
  INV_X1 U228 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U229 ( .A1(data_in[6]), .A2(n845), .B1(n1130), .B2(\mem[8][6] ), 
        .ZN(n1124) );
  INV_X1 U230 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U231 ( .A1(data_in[7]), .A2(n845), .B1(n1130), .B2(\mem[8][7] ), 
        .ZN(n1123) );
  INV_X1 U232 ( .A(n1121), .ZN(n813) );
  AOI22_X1 U233 ( .A1(data_in[0]), .A2(n844), .B1(n1120), .B2(\mem[9][0] ), 
        .ZN(n1121) );
  INV_X1 U234 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U235 ( .A1(data_in[1]), .A2(n844), .B1(n1120), .B2(\mem[9][1] ), 
        .ZN(n1119) );
  INV_X1 U236 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U237 ( .A1(data_in[2]), .A2(n844), .B1(n1120), .B2(\mem[9][2] ), 
        .ZN(n1118) );
  INV_X1 U238 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U239 ( .A1(data_in[3]), .A2(n844), .B1(n1120), .B2(\mem[9][3] ), 
        .ZN(n1117) );
  INV_X1 U240 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U241 ( .A1(data_in[4]), .A2(n844), .B1(n1120), .B2(\mem[9][4] ), 
        .ZN(n1116) );
  INV_X1 U242 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U243 ( .A1(data_in[5]), .A2(n844), .B1(n1120), .B2(\mem[9][5] ), 
        .ZN(n1115) );
  INV_X1 U244 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U245 ( .A1(data_in[6]), .A2(n844), .B1(n1120), .B2(\mem[9][6] ), 
        .ZN(n1114) );
  INV_X1 U246 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U247 ( .A1(data_in[7]), .A2(n844), .B1(n1120), .B2(\mem[9][7] ), 
        .ZN(n1113) );
  INV_X1 U248 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U249 ( .A1(data_in[0]), .A2(n843), .B1(n1111), .B2(\mem[10][0] ), 
        .ZN(n1112) );
  INV_X1 U250 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U251 ( .A1(data_in[1]), .A2(n843), .B1(n1111), .B2(\mem[10][1] ), 
        .ZN(n1110) );
  INV_X1 U252 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U253 ( .A1(data_in[2]), .A2(n843), .B1(n1111), .B2(\mem[10][2] ), 
        .ZN(n1109) );
  INV_X1 U254 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U255 ( .A1(data_in[3]), .A2(n843), .B1(n1111), .B2(\mem[10][3] ), 
        .ZN(n1108) );
  INV_X1 U256 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U257 ( .A1(data_in[4]), .A2(n843), .B1(n1111), .B2(\mem[10][4] ), 
        .ZN(n1107) );
  INV_X1 U258 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U259 ( .A1(data_in[5]), .A2(n843), .B1(n1111), .B2(\mem[10][5] ), 
        .ZN(n1106) );
  INV_X1 U260 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U261 ( .A1(data_in[6]), .A2(n843), .B1(n1111), .B2(\mem[10][6] ), 
        .ZN(n1105) );
  INV_X1 U262 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U263 ( .A1(data_in[7]), .A2(n843), .B1(n1111), .B2(\mem[10][7] ), 
        .ZN(n1104) );
  INV_X1 U264 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U265 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[11][0] ), 
        .ZN(n1103) );
  INV_X1 U266 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U267 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[11][1] ), 
        .ZN(n1101) );
  INV_X1 U268 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U269 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[11][2] ), 
        .ZN(n1100) );
  INV_X1 U270 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U271 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[11][3] ), 
        .ZN(n1099) );
  INV_X1 U272 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U273 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[11][4] ), 
        .ZN(n1098) );
  INV_X1 U274 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U275 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[11][5] ), 
        .ZN(n1097) );
  INV_X1 U276 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U277 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[11][6] ), 
        .ZN(n1096) );
  INV_X1 U278 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U279 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[11][7] ), 
        .ZN(n1095) );
  INV_X1 U280 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U281 ( .A1(data_in[0]), .A2(n841), .B1(n1093), .B2(\mem[12][0] ), 
        .ZN(n1094) );
  INV_X1 U282 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U283 ( .A1(data_in[1]), .A2(n841), .B1(n1093), .B2(\mem[12][1] ), 
        .ZN(n1092) );
  INV_X1 U284 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U285 ( .A1(data_in[2]), .A2(n841), .B1(n1093), .B2(\mem[12][2] ), 
        .ZN(n1091) );
  INV_X1 U286 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U287 ( .A1(data_in[3]), .A2(n841), .B1(n1093), .B2(\mem[12][3] ), 
        .ZN(n1090) );
  INV_X1 U288 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U289 ( .A1(data_in[4]), .A2(n841), .B1(n1093), .B2(\mem[12][4] ), 
        .ZN(n1089) );
  INV_X1 U290 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U291 ( .A1(data_in[5]), .A2(n841), .B1(n1093), .B2(\mem[12][5] ), 
        .ZN(n1088) );
  INV_X1 U292 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U293 ( .A1(data_in[6]), .A2(n841), .B1(n1093), .B2(\mem[12][6] ), 
        .ZN(n1087) );
  INV_X1 U294 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U295 ( .A1(data_in[7]), .A2(n841), .B1(n1093), .B2(\mem[12][7] ), 
        .ZN(n1086) );
  INV_X1 U296 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U297 ( .A1(data_in[0]), .A2(n840), .B1(n1084), .B2(\mem[13][0] ), 
        .ZN(n1085) );
  INV_X1 U298 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U299 ( .A1(data_in[1]), .A2(n840), .B1(n1084), .B2(\mem[13][1] ), 
        .ZN(n1083) );
  INV_X1 U300 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U301 ( .A1(data_in[2]), .A2(n840), .B1(n1084), .B2(\mem[13][2] ), 
        .ZN(n1082) );
  INV_X1 U302 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U303 ( .A1(data_in[3]), .A2(n840), .B1(n1084), .B2(\mem[13][3] ), 
        .ZN(n1081) );
  INV_X1 U304 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U305 ( .A1(data_in[4]), .A2(n840), .B1(n1084), .B2(\mem[13][4] ), 
        .ZN(n1080) );
  INV_X1 U306 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U307 ( .A1(data_in[5]), .A2(n840), .B1(n1084), .B2(\mem[13][5] ), 
        .ZN(n1079) );
  INV_X1 U308 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U309 ( .A1(data_in[6]), .A2(n840), .B1(n1084), .B2(\mem[13][6] ), 
        .ZN(n1078) );
  INV_X1 U310 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U311 ( .A1(data_in[7]), .A2(n840), .B1(n1084), .B2(\mem[13][7] ), 
        .ZN(n1077) );
  INV_X1 U312 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U313 ( .A1(data_in[0]), .A2(n839), .B1(n1075), .B2(\mem[14][0] ), 
        .ZN(n1076) );
  INV_X1 U314 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U315 ( .A1(data_in[1]), .A2(n839), .B1(n1075), .B2(\mem[14][1] ), 
        .ZN(n1074) );
  INV_X1 U316 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U317 ( .A1(data_in[2]), .A2(n839), .B1(n1075), .B2(\mem[14][2] ), 
        .ZN(n1073) );
  INV_X1 U318 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U319 ( .A1(data_in[3]), .A2(n839), .B1(n1075), .B2(\mem[14][3] ), 
        .ZN(n1072) );
  INV_X1 U320 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U321 ( .A1(data_in[4]), .A2(n839), .B1(n1075), .B2(\mem[14][4] ), 
        .ZN(n1071) );
  INV_X1 U322 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U323 ( .A1(data_in[5]), .A2(n839), .B1(n1075), .B2(\mem[14][5] ), 
        .ZN(n1070) );
  INV_X1 U324 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U325 ( .A1(data_in[6]), .A2(n839), .B1(n1075), .B2(\mem[14][6] ), 
        .ZN(n1069) );
  INV_X1 U326 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U327 ( .A1(data_in[7]), .A2(n839), .B1(n1075), .B2(\mem[14][7] ), 
        .ZN(n1068) );
  INV_X1 U328 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U329 ( .A1(data_in[0]), .A2(n838), .B1(n1066), .B2(\mem[15][0] ), 
        .ZN(n1067) );
  INV_X1 U330 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U331 ( .A1(data_in[1]), .A2(n838), .B1(n1066), .B2(\mem[15][1] ), 
        .ZN(n1065) );
  INV_X1 U332 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U333 ( .A1(data_in[2]), .A2(n838), .B1(n1066), .B2(\mem[15][2] ), 
        .ZN(n1064) );
  INV_X1 U334 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U335 ( .A1(data_in[3]), .A2(n838), .B1(n1066), .B2(\mem[15][3] ), 
        .ZN(n1063) );
  INV_X1 U336 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U337 ( .A1(data_in[4]), .A2(n838), .B1(n1066), .B2(\mem[15][4] ), 
        .ZN(n1062) );
  INV_X1 U338 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U339 ( .A1(data_in[5]), .A2(n838), .B1(n1066), .B2(\mem[15][5] ), 
        .ZN(n1061) );
  INV_X1 U340 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U341 ( .A1(data_in[6]), .A2(n838), .B1(n1066), .B2(\mem[15][6] ), 
        .ZN(n1060) );
  INV_X1 U342 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U343 ( .A1(data_in[7]), .A2(n838), .B1(n1066), .B2(\mem[15][7] ), 
        .ZN(n1059) );
  INV_X1 U344 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U345 ( .A1(data_in[0]), .A2(n837), .B1(n1057), .B2(\mem[16][0] ), 
        .ZN(n1058) );
  INV_X1 U346 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U347 ( .A1(data_in[1]), .A2(n837), .B1(n1057), .B2(\mem[16][1] ), 
        .ZN(n1056) );
  INV_X1 U348 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U349 ( .A1(data_in[2]), .A2(n837), .B1(n1057), .B2(\mem[16][2] ), 
        .ZN(n1055) );
  INV_X1 U350 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U351 ( .A1(data_in[3]), .A2(n837), .B1(n1057), .B2(\mem[16][3] ), 
        .ZN(n1054) );
  INV_X1 U352 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U353 ( .A1(data_in[4]), .A2(n837), .B1(n1057), .B2(\mem[16][4] ), 
        .ZN(n1053) );
  INV_X1 U354 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U355 ( .A1(data_in[5]), .A2(n837), .B1(n1057), .B2(\mem[16][5] ), 
        .ZN(n1052) );
  INV_X1 U356 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U357 ( .A1(data_in[6]), .A2(n837), .B1(n1057), .B2(\mem[16][6] ), 
        .ZN(n1051) );
  INV_X1 U358 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U359 ( .A1(data_in[7]), .A2(n837), .B1(n1057), .B2(\mem[16][7] ), 
        .ZN(n1050) );
  INV_X1 U360 ( .A(n1048), .ZN(n749) );
  AOI22_X1 U361 ( .A1(data_in[0]), .A2(n836), .B1(n1047), .B2(\mem[17][0] ), 
        .ZN(n1048) );
  INV_X1 U362 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U363 ( .A1(data_in[1]), .A2(n836), .B1(n1047), .B2(\mem[17][1] ), 
        .ZN(n1046) );
  INV_X1 U364 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U365 ( .A1(data_in[2]), .A2(n836), .B1(n1047), .B2(\mem[17][2] ), 
        .ZN(n1045) );
  INV_X1 U366 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U367 ( .A1(data_in[3]), .A2(n836), .B1(n1047), .B2(\mem[17][3] ), 
        .ZN(n1044) );
  INV_X1 U368 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U369 ( .A1(data_in[4]), .A2(n836), .B1(n1047), .B2(\mem[17][4] ), 
        .ZN(n1043) );
  INV_X1 U370 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U371 ( .A1(data_in[5]), .A2(n836), .B1(n1047), .B2(\mem[17][5] ), 
        .ZN(n1042) );
  INV_X1 U372 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U373 ( .A1(data_in[6]), .A2(n836), .B1(n1047), .B2(\mem[17][6] ), 
        .ZN(n1041) );
  INV_X1 U374 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U375 ( .A1(data_in[7]), .A2(n836), .B1(n1047), .B2(\mem[17][7] ), 
        .ZN(n1040) );
  INV_X1 U376 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U377 ( .A1(data_in[0]), .A2(n835), .B1(n1038), .B2(\mem[18][0] ), 
        .ZN(n1039) );
  INV_X1 U378 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U379 ( .A1(data_in[1]), .A2(n835), .B1(n1038), .B2(\mem[18][1] ), 
        .ZN(n1037) );
  INV_X1 U380 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U381 ( .A1(data_in[2]), .A2(n835), .B1(n1038), .B2(\mem[18][2] ), 
        .ZN(n1036) );
  INV_X1 U382 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U383 ( .A1(data_in[3]), .A2(n835), .B1(n1038), .B2(\mem[18][3] ), 
        .ZN(n1035) );
  INV_X1 U384 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U385 ( .A1(data_in[4]), .A2(n835), .B1(n1038), .B2(\mem[18][4] ), 
        .ZN(n1034) );
  INV_X1 U386 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U387 ( .A1(data_in[5]), .A2(n835), .B1(n1038), .B2(\mem[18][5] ), 
        .ZN(n1033) );
  INV_X1 U388 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U389 ( .A1(data_in[6]), .A2(n835), .B1(n1038), .B2(\mem[18][6] ), 
        .ZN(n1032) );
  INV_X1 U390 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U391 ( .A1(data_in[7]), .A2(n835), .B1(n1038), .B2(\mem[18][7] ), 
        .ZN(n1031) );
  INV_X1 U392 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U393 ( .A1(data_in[0]), .A2(n834), .B1(n1029), .B2(\mem[19][0] ), 
        .ZN(n1030) );
  INV_X1 U394 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U395 ( .A1(data_in[1]), .A2(n834), .B1(n1029), .B2(\mem[19][1] ), 
        .ZN(n1028) );
  INV_X1 U396 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U397 ( .A1(data_in[2]), .A2(n834), .B1(n1029), .B2(\mem[19][2] ), 
        .ZN(n1027) );
  INV_X1 U398 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U399 ( .A1(data_in[3]), .A2(n834), .B1(n1029), .B2(\mem[19][3] ), 
        .ZN(n1026) );
  INV_X1 U400 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U401 ( .A1(data_in[4]), .A2(n834), .B1(n1029), .B2(\mem[19][4] ), 
        .ZN(n1025) );
  INV_X1 U402 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U403 ( .A1(data_in[5]), .A2(n834), .B1(n1029), .B2(\mem[19][5] ), 
        .ZN(n1024) );
  INV_X1 U404 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U405 ( .A1(data_in[6]), .A2(n834), .B1(n1029), .B2(\mem[19][6] ), 
        .ZN(n1023) );
  INV_X1 U406 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U407 ( .A1(data_in[7]), .A2(n834), .B1(n1029), .B2(\mem[19][7] ), 
        .ZN(n1022) );
  INV_X1 U408 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U409 ( .A1(data_in[0]), .A2(n833), .B1(n1020), .B2(\mem[20][0] ), 
        .ZN(n1021) );
  INV_X1 U410 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U411 ( .A1(data_in[1]), .A2(n833), .B1(n1020), .B2(\mem[20][1] ), 
        .ZN(n1019) );
  INV_X1 U412 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U413 ( .A1(data_in[2]), .A2(n833), .B1(n1020), .B2(\mem[20][2] ), 
        .ZN(n1018) );
  INV_X1 U414 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U415 ( .A1(data_in[3]), .A2(n833), .B1(n1020), .B2(\mem[20][3] ), 
        .ZN(n1017) );
  INV_X1 U416 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U417 ( .A1(data_in[4]), .A2(n833), .B1(n1020), .B2(\mem[20][4] ), 
        .ZN(n1016) );
  INV_X1 U418 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U419 ( .A1(data_in[5]), .A2(n833), .B1(n1020), .B2(\mem[20][5] ), 
        .ZN(n1015) );
  INV_X1 U420 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U421 ( .A1(data_in[6]), .A2(n833), .B1(n1020), .B2(\mem[20][6] ), 
        .ZN(n1014) );
  INV_X1 U422 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U423 ( .A1(data_in[7]), .A2(n833), .B1(n1020), .B2(\mem[20][7] ), 
        .ZN(n1013) );
  INV_X1 U424 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U425 ( .A1(data_in[0]), .A2(n832), .B1(n1011), .B2(\mem[21][0] ), 
        .ZN(n1012) );
  INV_X1 U426 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U427 ( .A1(data_in[1]), .A2(n832), .B1(n1011), .B2(\mem[21][1] ), 
        .ZN(n1010) );
  INV_X1 U428 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U429 ( .A1(data_in[2]), .A2(n832), .B1(n1011), .B2(\mem[21][2] ), 
        .ZN(n1009) );
  INV_X1 U430 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U431 ( .A1(data_in[3]), .A2(n832), .B1(n1011), .B2(\mem[21][3] ), 
        .ZN(n1008) );
  INV_X1 U432 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U433 ( .A1(data_in[4]), .A2(n832), .B1(n1011), .B2(\mem[21][4] ), 
        .ZN(n1007) );
  INV_X1 U434 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U435 ( .A1(data_in[5]), .A2(n832), .B1(n1011), .B2(\mem[21][5] ), 
        .ZN(n1006) );
  INV_X1 U436 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U437 ( .A1(data_in[6]), .A2(n832), .B1(n1011), .B2(\mem[21][6] ), 
        .ZN(n1005) );
  INV_X1 U438 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U439 ( .A1(data_in[7]), .A2(n832), .B1(n1011), .B2(\mem[21][7] ), 
        .ZN(n1004) );
  INV_X1 U440 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U441 ( .A1(data_in[0]), .A2(n831), .B1(n1002), .B2(\mem[22][0] ), 
        .ZN(n1003) );
  INV_X1 U442 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U443 ( .A1(data_in[1]), .A2(n831), .B1(n1002), .B2(\mem[22][1] ), 
        .ZN(n1001) );
  INV_X1 U444 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U445 ( .A1(data_in[2]), .A2(n831), .B1(n1002), .B2(\mem[22][2] ), 
        .ZN(n1000) );
  INV_X1 U446 ( .A(n999), .ZN(n706) );
  AOI22_X1 U447 ( .A1(data_in[3]), .A2(n831), .B1(n1002), .B2(\mem[22][3] ), 
        .ZN(n999) );
  INV_X1 U448 ( .A(n998), .ZN(n705) );
  AOI22_X1 U449 ( .A1(data_in[4]), .A2(n831), .B1(n1002), .B2(\mem[22][4] ), 
        .ZN(n998) );
  INV_X1 U450 ( .A(n997), .ZN(n704) );
  AOI22_X1 U451 ( .A1(data_in[5]), .A2(n831), .B1(n1002), .B2(\mem[22][5] ), 
        .ZN(n997) );
  INV_X1 U452 ( .A(n996), .ZN(n703) );
  AOI22_X1 U453 ( .A1(data_in[6]), .A2(n831), .B1(n1002), .B2(\mem[22][6] ), 
        .ZN(n996) );
  INV_X1 U454 ( .A(n995), .ZN(n702) );
  AOI22_X1 U455 ( .A1(data_in[7]), .A2(n831), .B1(n1002), .B2(\mem[22][7] ), 
        .ZN(n995) );
  INV_X1 U456 ( .A(n994), .ZN(n701) );
  AOI22_X1 U457 ( .A1(data_in[0]), .A2(n830), .B1(n993), .B2(\mem[23][0] ), 
        .ZN(n994) );
  INV_X1 U458 ( .A(n992), .ZN(n700) );
  AOI22_X1 U459 ( .A1(data_in[1]), .A2(n830), .B1(n993), .B2(\mem[23][1] ), 
        .ZN(n992) );
  INV_X1 U460 ( .A(n991), .ZN(n699) );
  AOI22_X1 U461 ( .A1(data_in[2]), .A2(n830), .B1(n993), .B2(\mem[23][2] ), 
        .ZN(n991) );
  INV_X1 U462 ( .A(n990), .ZN(n698) );
  AOI22_X1 U463 ( .A1(data_in[3]), .A2(n830), .B1(n993), .B2(\mem[23][3] ), 
        .ZN(n990) );
  INV_X1 U464 ( .A(n989), .ZN(n697) );
  AOI22_X1 U465 ( .A1(data_in[4]), .A2(n830), .B1(n993), .B2(\mem[23][4] ), 
        .ZN(n989) );
  INV_X1 U466 ( .A(n988), .ZN(n696) );
  AOI22_X1 U467 ( .A1(data_in[5]), .A2(n830), .B1(n993), .B2(\mem[23][5] ), 
        .ZN(n988) );
  INV_X1 U468 ( .A(n987), .ZN(n695) );
  AOI22_X1 U469 ( .A1(data_in[6]), .A2(n830), .B1(n993), .B2(\mem[23][6] ), 
        .ZN(n987) );
  INV_X1 U470 ( .A(n986), .ZN(n694) );
  AOI22_X1 U471 ( .A1(data_in[7]), .A2(n830), .B1(n993), .B2(\mem[23][7] ), 
        .ZN(n986) );
  INV_X1 U472 ( .A(n985), .ZN(n693) );
  AOI22_X1 U473 ( .A1(data_in[0]), .A2(n829), .B1(n984), .B2(\mem[24][0] ), 
        .ZN(n985) );
  INV_X1 U474 ( .A(n983), .ZN(n692) );
  AOI22_X1 U475 ( .A1(data_in[1]), .A2(n829), .B1(n984), .B2(\mem[24][1] ), 
        .ZN(n983) );
  INV_X1 U476 ( .A(n982), .ZN(n691) );
  AOI22_X1 U477 ( .A1(data_in[2]), .A2(n829), .B1(n984), .B2(\mem[24][2] ), 
        .ZN(n982) );
  INV_X1 U478 ( .A(n981), .ZN(n690) );
  AOI22_X1 U479 ( .A1(data_in[3]), .A2(n829), .B1(n984), .B2(\mem[24][3] ), 
        .ZN(n981) );
  INV_X1 U480 ( .A(n980), .ZN(n689) );
  AOI22_X1 U481 ( .A1(data_in[4]), .A2(n829), .B1(n984), .B2(\mem[24][4] ), 
        .ZN(n980) );
  INV_X1 U482 ( .A(n979), .ZN(n688) );
  AOI22_X1 U483 ( .A1(data_in[5]), .A2(n829), .B1(n984), .B2(\mem[24][5] ), 
        .ZN(n979) );
  INV_X1 U484 ( .A(n978), .ZN(n687) );
  AOI22_X1 U485 ( .A1(data_in[6]), .A2(n829), .B1(n984), .B2(\mem[24][6] ), 
        .ZN(n978) );
  INV_X1 U486 ( .A(n977), .ZN(n686) );
  AOI22_X1 U487 ( .A1(data_in[7]), .A2(n829), .B1(n984), .B2(\mem[24][7] ), 
        .ZN(n977) );
  INV_X1 U488 ( .A(n975), .ZN(n685) );
  AOI22_X1 U489 ( .A1(data_in[0]), .A2(n828), .B1(n974), .B2(\mem[25][0] ), 
        .ZN(n975) );
  INV_X1 U490 ( .A(n973), .ZN(n684) );
  AOI22_X1 U491 ( .A1(data_in[1]), .A2(n828), .B1(n974), .B2(\mem[25][1] ), 
        .ZN(n973) );
  INV_X1 U492 ( .A(n972), .ZN(n683) );
  AOI22_X1 U493 ( .A1(data_in[2]), .A2(n828), .B1(n974), .B2(\mem[25][2] ), 
        .ZN(n972) );
  INV_X1 U494 ( .A(n971), .ZN(n682) );
  AOI22_X1 U495 ( .A1(data_in[3]), .A2(n828), .B1(n974), .B2(\mem[25][3] ), 
        .ZN(n971) );
  INV_X1 U496 ( .A(n970), .ZN(n681) );
  AOI22_X1 U497 ( .A1(data_in[4]), .A2(n828), .B1(n974), .B2(\mem[25][4] ), 
        .ZN(n970) );
  INV_X1 U498 ( .A(n969), .ZN(n680) );
  AOI22_X1 U499 ( .A1(data_in[5]), .A2(n828), .B1(n974), .B2(\mem[25][5] ), 
        .ZN(n969) );
  INV_X1 U500 ( .A(n968), .ZN(n679) );
  AOI22_X1 U501 ( .A1(data_in[6]), .A2(n828), .B1(n974), .B2(\mem[25][6] ), 
        .ZN(n968) );
  INV_X1 U502 ( .A(n967), .ZN(n678) );
  AOI22_X1 U503 ( .A1(data_in[7]), .A2(n828), .B1(n974), .B2(\mem[25][7] ), 
        .ZN(n967) );
  INV_X1 U504 ( .A(n966), .ZN(n677) );
  AOI22_X1 U505 ( .A1(data_in[0]), .A2(n827), .B1(n965), .B2(\mem[26][0] ), 
        .ZN(n966) );
  INV_X1 U506 ( .A(n964), .ZN(n676) );
  AOI22_X1 U507 ( .A1(data_in[1]), .A2(n827), .B1(n965), .B2(\mem[26][1] ), 
        .ZN(n964) );
  INV_X1 U508 ( .A(n963), .ZN(n675) );
  AOI22_X1 U509 ( .A1(data_in[2]), .A2(n827), .B1(n965), .B2(\mem[26][2] ), 
        .ZN(n963) );
  INV_X1 U510 ( .A(n962), .ZN(n674) );
  AOI22_X1 U511 ( .A1(data_in[3]), .A2(n827), .B1(n965), .B2(\mem[26][3] ), 
        .ZN(n962) );
  INV_X1 U512 ( .A(n961), .ZN(n673) );
  AOI22_X1 U513 ( .A1(data_in[4]), .A2(n827), .B1(n965), .B2(\mem[26][4] ), 
        .ZN(n961) );
  INV_X1 U514 ( .A(n960), .ZN(n672) );
  AOI22_X1 U515 ( .A1(data_in[5]), .A2(n827), .B1(n965), .B2(\mem[26][5] ), 
        .ZN(n960) );
  INV_X1 U516 ( .A(n959), .ZN(n671) );
  AOI22_X1 U517 ( .A1(data_in[6]), .A2(n827), .B1(n965), .B2(\mem[26][6] ), 
        .ZN(n959) );
  INV_X1 U518 ( .A(n958), .ZN(n670) );
  AOI22_X1 U519 ( .A1(data_in[7]), .A2(n827), .B1(n965), .B2(\mem[26][7] ), 
        .ZN(n958) );
  INV_X1 U520 ( .A(n957), .ZN(n669) );
  AOI22_X1 U521 ( .A1(data_in[0]), .A2(n826), .B1(n956), .B2(\mem[27][0] ), 
        .ZN(n957) );
  INV_X1 U522 ( .A(n955), .ZN(n668) );
  AOI22_X1 U523 ( .A1(data_in[1]), .A2(n826), .B1(n956), .B2(\mem[27][1] ), 
        .ZN(n955) );
  INV_X1 U524 ( .A(n954), .ZN(n667) );
  AOI22_X1 U525 ( .A1(data_in[2]), .A2(n826), .B1(n956), .B2(\mem[27][2] ), 
        .ZN(n954) );
  INV_X1 U526 ( .A(n953), .ZN(n666) );
  AOI22_X1 U527 ( .A1(data_in[3]), .A2(n826), .B1(n956), .B2(\mem[27][3] ), 
        .ZN(n953) );
  INV_X1 U528 ( .A(n952), .ZN(n665) );
  AOI22_X1 U529 ( .A1(data_in[4]), .A2(n826), .B1(n956), .B2(\mem[27][4] ), 
        .ZN(n952) );
  INV_X1 U530 ( .A(n951), .ZN(n664) );
  AOI22_X1 U531 ( .A1(data_in[5]), .A2(n826), .B1(n956), .B2(\mem[27][5] ), 
        .ZN(n951) );
  INV_X1 U532 ( .A(n950), .ZN(n663) );
  AOI22_X1 U533 ( .A1(data_in[6]), .A2(n826), .B1(n956), .B2(\mem[27][6] ), 
        .ZN(n950) );
  INV_X1 U534 ( .A(n949), .ZN(n662) );
  AOI22_X1 U535 ( .A1(data_in[7]), .A2(n826), .B1(n956), .B2(\mem[27][7] ), 
        .ZN(n949) );
  INV_X1 U536 ( .A(n948), .ZN(n661) );
  AOI22_X1 U537 ( .A1(data_in[0]), .A2(n825), .B1(n947), .B2(\mem[28][0] ), 
        .ZN(n948) );
  INV_X1 U538 ( .A(n946), .ZN(n660) );
  AOI22_X1 U539 ( .A1(data_in[1]), .A2(n825), .B1(n947), .B2(\mem[28][1] ), 
        .ZN(n946) );
  INV_X1 U540 ( .A(n945), .ZN(n659) );
  AOI22_X1 U541 ( .A1(data_in[2]), .A2(n825), .B1(n947), .B2(\mem[28][2] ), 
        .ZN(n945) );
  INV_X1 U542 ( .A(n944), .ZN(n658) );
  AOI22_X1 U543 ( .A1(data_in[3]), .A2(n825), .B1(n947), .B2(\mem[28][3] ), 
        .ZN(n944) );
  INV_X1 U544 ( .A(n943), .ZN(n657) );
  AOI22_X1 U545 ( .A1(data_in[4]), .A2(n825), .B1(n947), .B2(\mem[28][4] ), 
        .ZN(n943) );
  INV_X1 U546 ( .A(n942), .ZN(n656) );
  AOI22_X1 U547 ( .A1(data_in[5]), .A2(n825), .B1(n947), .B2(\mem[28][5] ), 
        .ZN(n942) );
  INV_X1 U548 ( .A(n941), .ZN(n655) );
  AOI22_X1 U549 ( .A1(data_in[6]), .A2(n825), .B1(n947), .B2(\mem[28][6] ), 
        .ZN(n941) );
  INV_X1 U550 ( .A(n940), .ZN(n654) );
  AOI22_X1 U551 ( .A1(data_in[7]), .A2(n825), .B1(n947), .B2(\mem[28][7] ), 
        .ZN(n940) );
  INV_X1 U552 ( .A(n939), .ZN(n653) );
  AOI22_X1 U553 ( .A1(data_in[0]), .A2(n824), .B1(n938), .B2(\mem[29][0] ), 
        .ZN(n939) );
  INV_X1 U554 ( .A(n937), .ZN(n652) );
  AOI22_X1 U555 ( .A1(data_in[1]), .A2(n824), .B1(n938), .B2(\mem[29][1] ), 
        .ZN(n937) );
  INV_X1 U556 ( .A(n936), .ZN(n651) );
  AOI22_X1 U557 ( .A1(data_in[2]), .A2(n824), .B1(n938), .B2(\mem[29][2] ), 
        .ZN(n936) );
  INV_X1 U558 ( .A(n935), .ZN(n650) );
  AOI22_X1 U559 ( .A1(data_in[3]), .A2(n824), .B1(n938), .B2(\mem[29][3] ), 
        .ZN(n935) );
  INV_X1 U560 ( .A(n934), .ZN(n649) );
  AOI22_X1 U561 ( .A1(data_in[4]), .A2(n824), .B1(n938), .B2(\mem[29][4] ), 
        .ZN(n934) );
  INV_X1 U562 ( .A(n933), .ZN(n648) );
  AOI22_X1 U563 ( .A1(data_in[5]), .A2(n824), .B1(n938), .B2(\mem[29][5] ), 
        .ZN(n933) );
  INV_X1 U564 ( .A(n932), .ZN(n647) );
  AOI22_X1 U565 ( .A1(data_in[6]), .A2(n824), .B1(n938), .B2(\mem[29][6] ), 
        .ZN(n932) );
  INV_X1 U566 ( .A(n931), .ZN(n646) );
  AOI22_X1 U567 ( .A1(data_in[7]), .A2(n824), .B1(n938), .B2(\mem[29][7] ), 
        .ZN(n931) );
  INV_X1 U568 ( .A(n930), .ZN(n645) );
  AOI22_X1 U569 ( .A1(data_in[0]), .A2(n823), .B1(n929), .B2(\mem[30][0] ), 
        .ZN(n930) );
  INV_X1 U570 ( .A(n928), .ZN(n644) );
  AOI22_X1 U571 ( .A1(data_in[1]), .A2(n823), .B1(n929), .B2(\mem[30][1] ), 
        .ZN(n928) );
  INV_X1 U572 ( .A(n927), .ZN(n643) );
  AOI22_X1 U573 ( .A1(data_in[2]), .A2(n823), .B1(n929), .B2(\mem[30][2] ), 
        .ZN(n927) );
  INV_X1 U574 ( .A(n926), .ZN(n642) );
  AOI22_X1 U575 ( .A1(data_in[3]), .A2(n823), .B1(n929), .B2(\mem[30][3] ), 
        .ZN(n926) );
  INV_X1 U576 ( .A(n925), .ZN(n641) );
  AOI22_X1 U577 ( .A1(data_in[4]), .A2(n823), .B1(n929), .B2(\mem[30][4] ), 
        .ZN(n925) );
  INV_X1 U578 ( .A(n924), .ZN(n640) );
  AOI22_X1 U579 ( .A1(data_in[5]), .A2(n823), .B1(n929), .B2(\mem[30][5] ), 
        .ZN(n924) );
  INV_X1 U580 ( .A(n923), .ZN(n639) );
  AOI22_X1 U581 ( .A1(data_in[6]), .A2(n823), .B1(n929), .B2(\mem[30][6] ), 
        .ZN(n923) );
  INV_X1 U582 ( .A(n922), .ZN(n638) );
  AOI22_X1 U583 ( .A1(data_in[7]), .A2(n823), .B1(n929), .B2(\mem[30][7] ), 
        .ZN(n922) );
  INV_X1 U584 ( .A(n921), .ZN(n637) );
  AOI22_X1 U585 ( .A1(data_in[0]), .A2(n822), .B1(n920), .B2(\mem[31][0] ), 
        .ZN(n921) );
  INV_X1 U586 ( .A(n919), .ZN(n636) );
  AOI22_X1 U587 ( .A1(data_in[1]), .A2(n822), .B1(n920), .B2(\mem[31][1] ), 
        .ZN(n919) );
  INV_X1 U588 ( .A(n918), .ZN(n635) );
  AOI22_X1 U589 ( .A1(data_in[2]), .A2(n822), .B1(n920), .B2(\mem[31][2] ), 
        .ZN(n918) );
  INV_X1 U590 ( .A(n917), .ZN(n634) );
  AOI22_X1 U591 ( .A1(data_in[3]), .A2(n822), .B1(n920), .B2(\mem[31][3] ), 
        .ZN(n917) );
  INV_X1 U592 ( .A(n916), .ZN(n633) );
  AOI22_X1 U593 ( .A1(data_in[4]), .A2(n822), .B1(n920), .B2(\mem[31][4] ), 
        .ZN(n916) );
  INV_X1 U594 ( .A(n915), .ZN(n632) );
  AOI22_X1 U595 ( .A1(data_in[5]), .A2(n822), .B1(n920), .B2(\mem[31][5] ), 
        .ZN(n915) );
  INV_X1 U596 ( .A(n914), .ZN(n631) );
  AOI22_X1 U597 ( .A1(data_in[6]), .A2(n822), .B1(n920), .B2(\mem[31][6] ), 
        .ZN(n914) );
  INV_X1 U598 ( .A(n913), .ZN(n630) );
  AOI22_X1 U599 ( .A1(data_in[7]), .A2(n822), .B1(n920), .B2(\mem[31][7] ), 
        .ZN(n913) );
  MUX2_X1 U600 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n611), .Z(n1) );
  MUX2_X1 U601 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n611), .Z(n2) );
  MUX2_X1 U602 ( .A(n2), .B(n1), .S(n608), .Z(n3) );
  MUX2_X1 U603 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n611), .Z(n4) );
  MUX2_X1 U604 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n611), .Z(n5) );
  MUX2_X1 U605 ( .A(n5), .B(n4), .S(n608), .Z(n6) );
  MUX2_X1 U606 ( .A(n6), .B(n3), .S(n606), .Z(n7) );
  MUX2_X1 U607 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n611), .Z(n8) );
  MUX2_X1 U608 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n611), .Z(n9) );
  MUX2_X1 U609 ( .A(n9), .B(n8), .S(n608), .Z(n10) );
  MUX2_X1 U610 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n611), .Z(n11) );
  MUX2_X1 U611 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n611), .Z(n12) );
  MUX2_X1 U612 ( .A(n12), .B(n11), .S(n608), .Z(n13) );
  MUX2_X1 U613 ( .A(n13), .B(n10), .S(n606), .Z(n14) );
  MUX2_X1 U614 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U615 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n619), .Z(n16) );
  MUX2_X1 U616 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(N10), .Z(n17) );
  MUX2_X1 U617 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U618 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n619), .Z(n19) );
  MUX2_X1 U619 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n20) );
  MUX2_X1 U620 ( .A(n20), .B(n19), .S(n609), .Z(n21) );
  MUX2_X1 U621 ( .A(n21), .B(n18), .S(n606), .Z(n22) );
  MUX2_X1 U622 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n619), .Z(n23) );
  MUX2_X1 U623 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n24) );
  MUX2_X1 U624 ( .A(n24), .B(n23), .S(n609), .Z(n25) );
  MUX2_X1 U625 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n26) );
  MUX2_X1 U626 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n27) );
  MUX2_X1 U627 ( .A(n27), .B(n26), .S(N11), .Z(n28) );
  MUX2_X1 U628 ( .A(n28), .B(n25), .S(n606), .Z(n29) );
  MUX2_X1 U629 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U630 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U631 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(N10), .Z(n31) );
  MUX2_X1 U632 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n616), .Z(n32) );
  MUX2_X1 U633 ( .A(n32), .B(n31), .S(n608), .Z(n33) );
  MUX2_X1 U634 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n619), .Z(n34) );
  MUX2_X1 U635 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n617), .Z(n35) );
  MUX2_X1 U636 ( .A(n35), .B(n34), .S(n609), .Z(n36) );
  MUX2_X1 U637 ( .A(n36), .B(n33), .S(n606), .Z(n37) );
  MUX2_X1 U638 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n611), .Z(n38) );
  MUX2_X1 U639 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n611), .Z(n39) );
  MUX2_X1 U640 ( .A(n39), .B(n38), .S(n608), .Z(n40) );
  MUX2_X1 U641 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n611), .Z(n41) );
  MUX2_X1 U642 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n618), .Z(n42) );
  MUX2_X1 U643 ( .A(n42), .B(n41), .S(n608), .Z(n43) );
  MUX2_X1 U644 ( .A(n43), .B(n40), .S(n606), .Z(n44) );
  MUX2_X1 U645 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U646 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n614), .Z(n46) );
  MUX2_X1 U647 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n618), .Z(n47) );
  MUX2_X1 U648 ( .A(n47), .B(n46), .S(n609), .Z(n48) );
  MUX2_X1 U649 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n611), .Z(n49) );
  MUX2_X1 U650 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n615), .Z(n50) );
  MUX2_X1 U651 ( .A(n50), .B(n49), .S(n610), .Z(n51) );
  MUX2_X1 U652 ( .A(n51), .B(n48), .S(n606), .Z(n52) );
  MUX2_X1 U653 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n617), .Z(n53) );
  MUX2_X1 U654 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n615), .Z(n54) );
  MUX2_X1 U655 ( .A(n54), .B(n53), .S(n609), .Z(n55) );
  MUX2_X1 U656 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n619), .Z(n56) );
  MUX2_X1 U657 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n619), .Z(n57) );
  MUX2_X1 U658 ( .A(n57), .B(n56), .S(N11), .Z(n58) );
  MUX2_X1 U659 ( .A(n58), .B(n55), .S(n606), .Z(n59) );
  MUX2_X1 U660 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U661 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U662 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n612), .Z(n61) );
  MUX2_X1 U663 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n612), .Z(n62) );
  MUX2_X1 U664 ( .A(n62), .B(n61), .S(n608), .Z(n63) );
  MUX2_X1 U665 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n612), .Z(n64) );
  MUX2_X1 U666 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n612), .Z(n65) );
  MUX2_X1 U667 ( .A(n65), .B(n64), .S(n608), .Z(n66) );
  MUX2_X1 U668 ( .A(n66), .B(n63), .S(n607), .Z(n67) );
  MUX2_X1 U669 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n612), .Z(n68) );
  MUX2_X1 U670 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n612), .Z(n69) );
  MUX2_X1 U671 ( .A(n69), .B(n68), .S(N11), .Z(n70) );
  MUX2_X1 U672 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n612), .Z(n71) );
  MUX2_X1 U673 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n612), .Z(n72) );
  MUX2_X1 U674 ( .A(n72), .B(n71), .S(N11), .Z(n73) );
  MUX2_X1 U675 ( .A(n73), .B(n70), .S(n607), .Z(n74) );
  MUX2_X1 U676 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U677 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n612), .Z(n76) );
  MUX2_X1 U678 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n612), .Z(n77) );
  MUX2_X1 U679 ( .A(n77), .B(n76), .S(n608), .Z(n78) );
  MUX2_X1 U680 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n612), .Z(n79) );
  MUX2_X1 U681 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n612), .Z(n80) );
  MUX2_X1 U682 ( .A(n80), .B(n79), .S(n610), .Z(n81) );
  MUX2_X1 U683 ( .A(n81), .B(n78), .S(n607), .Z(n82) );
  MUX2_X1 U684 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n613), .Z(n83) );
  MUX2_X1 U685 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n613), .Z(n84) );
  MUX2_X1 U686 ( .A(n84), .B(n83), .S(n609), .Z(n85) );
  MUX2_X1 U687 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n613), .Z(n86) );
  MUX2_X1 U688 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n613), .Z(n87) );
  MUX2_X1 U689 ( .A(n87), .B(n86), .S(n609), .Z(n88) );
  MUX2_X1 U690 ( .A(n88), .B(n85), .S(n607), .Z(n89) );
  MUX2_X1 U691 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U692 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U693 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n613), .Z(n91) );
  MUX2_X1 U694 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n613), .Z(n92) );
  MUX2_X1 U695 ( .A(n92), .B(n91), .S(n608), .Z(n93) );
  MUX2_X1 U696 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n613), .Z(n94) );
  MUX2_X1 U697 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n613), .Z(n95) );
  MUX2_X1 U698 ( .A(n95), .B(n94), .S(n608), .Z(n96) );
  MUX2_X1 U699 ( .A(n96), .B(n93), .S(n607), .Z(n97) );
  MUX2_X1 U700 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n613), .Z(n98) );
  MUX2_X1 U701 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n613), .Z(n99) );
  MUX2_X1 U702 ( .A(n99), .B(n98), .S(n608), .Z(n100) );
  MUX2_X1 U703 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n613), .Z(n101) );
  MUX2_X1 U704 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n613), .Z(n102) );
  MUX2_X1 U705 ( .A(n102), .B(n101), .S(n608), .Z(n103) );
  MUX2_X1 U706 ( .A(n103), .B(n100), .S(n607), .Z(n104) );
  MUX2_X1 U707 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U708 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n614), .Z(n106) );
  MUX2_X1 U709 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n614), .Z(n107) );
  MUX2_X1 U710 ( .A(n107), .B(n106), .S(n609), .Z(n108) );
  MUX2_X1 U711 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n614), .Z(n109) );
  MUX2_X1 U712 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n614), .Z(n110) );
  MUX2_X1 U713 ( .A(n110), .B(n109), .S(n609), .Z(n111) );
  MUX2_X1 U714 ( .A(n111), .B(n108), .S(n607), .Z(n112) );
  MUX2_X1 U715 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n614), .Z(n113) );
  MUX2_X1 U716 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n614), .Z(n114) );
  MUX2_X1 U717 ( .A(n114), .B(n113), .S(n609), .Z(n115) );
  MUX2_X1 U718 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n614), .Z(n116) );
  MUX2_X1 U719 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n614), .Z(n117) );
  MUX2_X1 U720 ( .A(n117), .B(n116), .S(n609), .Z(n118) );
  MUX2_X1 U721 ( .A(n118), .B(n115), .S(n607), .Z(n119) );
  MUX2_X1 U722 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U723 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U724 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n614), .Z(n121) );
  MUX2_X1 U725 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n614), .Z(n122) );
  MUX2_X1 U726 ( .A(n122), .B(n121), .S(n609), .Z(n123) );
  MUX2_X1 U727 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n614), .Z(n124) );
  MUX2_X1 U728 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n614), .Z(n125) );
  MUX2_X1 U729 ( .A(n125), .B(n124), .S(n609), .Z(n126) );
  MUX2_X1 U730 ( .A(n126), .B(n123), .S(n607), .Z(n127) );
  MUX2_X1 U731 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n615), .Z(n128) );
  MUX2_X1 U732 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n615), .Z(n129) );
  MUX2_X1 U733 ( .A(n129), .B(n128), .S(n609), .Z(n130) );
  MUX2_X1 U734 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n615), .Z(n131) );
  MUX2_X1 U735 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n615), .Z(n132) );
  MUX2_X1 U736 ( .A(n132), .B(n131), .S(n609), .Z(n133) );
  MUX2_X1 U737 ( .A(n133), .B(n130), .S(n607), .Z(n134) );
  MUX2_X1 U738 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U739 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n615), .Z(n136) );
  MUX2_X1 U740 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n615), .Z(n137) );
  MUX2_X1 U741 ( .A(n137), .B(n136), .S(n609), .Z(n138) );
  MUX2_X1 U742 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n615), .Z(n139) );
  MUX2_X1 U743 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n615), .Z(n140) );
  MUX2_X1 U744 ( .A(n140), .B(n139), .S(n609), .Z(n141) );
  MUX2_X1 U745 ( .A(n141), .B(n138), .S(n607), .Z(n142) );
  MUX2_X1 U746 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n615), .Z(n143) );
  MUX2_X1 U747 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n615), .Z(n144) );
  MUX2_X1 U748 ( .A(n144), .B(n143), .S(n609), .Z(n145) );
  MUX2_X1 U749 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n615), .Z(n146) );
  MUX2_X1 U750 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n615), .Z(n147) );
  MUX2_X1 U751 ( .A(n147), .B(n146), .S(n609), .Z(n148) );
  MUX2_X1 U752 ( .A(n148), .B(n145), .S(n607), .Z(n149) );
  MUX2_X1 U753 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U754 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U755 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n611), .Z(n151) );
  MUX2_X1 U756 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n614), .Z(n152) );
  MUX2_X1 U757 ( .A(n152), .B(n151), .S(n610), .Z(n153) );
  MUX2_X1 U758 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n613), .Z(n154) );
  MUX2_X1 U759 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n611), .Z(n155) );
  MUX2_X1 U760 ( .A(n155), .B(n154), .S(n610), .Z(n156) );
  MUX2_X1 U761 ( .A(n156), .B(n153), .S(n606), .Z(n157) );
  MUX2_X1 U762 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n616), .Z(n158) );
  MUX2_X1 U763 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n619), .Z(n159) );
  MUX2_X1 U764 ( .A(n159), .B(n158), .S(n610), .Z(n160) );
  MUX2_X1 U765 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n613), .Z(n161) );
  MUX2_X1 U766 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n619), .Z(n162) );
  MUX2_X1 U767 ( .A(n162), .B(n161), .S(n610), .Z(n163) );
  MUX2_X1 U768 ( .A(n163), .B(n160), .S(n606), .Z(n164) );
  MUX2_X1 U769 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U770 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n612), .Z(n166) );
  MUX2_X1 U771 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n619), .Z(n167) );
  MUX2_X1 U772 ( .A(n167), .B(n166), .S(n610), .Z(n168) );
  MUX2_X1 U773 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n612), .Z(n169) );
  MUX2_X1 U774 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n619), .Z(n170) );
  MUX2_X1 U775 ( .A(n170), .B(n169), .S(n610), .Z(n171) );
  MUX2_X1 U776 ( .A(n171), .B(n168), .S(n606), .Z(n172) );
  MUX2_X1 U777 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n616), .Z(n173) );
  MUX2_X1 U778 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n616), .Z(n174) );
  MUX2_X1 U779 ( .A(n174), .B(n173), .S(n610), .Z(n175) );
  MUX2_X1 U780 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n616), .Z(n176) );
  MUX2_X1 U781 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n616), .Z(n177) );
  MUX2_X1 U782 ( .A(n177), .B(n176), .S(n610), .Z(n178) );
  MUX2_X1 U783 ( .A(n178), .B(n175), .S(n606), .Z(n179) );
  MUX2_X1 U784 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U785 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U786 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n616), .Z(n181) );
  MUX2_X1 U787 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n616), .Z(n182) );
  MUX2_X1 U788 ( .A(n182), .B(n181), .S(n610), .Z(n183) );
  MUX2_X1 U789 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n616), .Z(n184) );
  MUX2_X1 U790 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n616), .Z(n185) );
  MUX2_X1 U791 ( .A(n185), .B(n184), .S(n610), .Z(n186) );
  MUX2_X1 U792 ( .A(n186), .B(n183), .S(n607), .Z(n187) );
  MUX2_X1 U793 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n616), .Z(n188) );
  MUX2_X1 U794 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n616), .Z(n189) );
  MUX2_X1 U795 ( .A(n189), .B(n188), .S(n610), .Z(n190) );
  MUX2_X1 U796 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n616), .Z(n191) );
  MUX2_X1 U797 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n616), .Z(n192) );
  MUX2_X1 U798 ( .A(n192), .B(n191), .S(n610), .Z(n193) );
  MUX2_X1 U799 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U800 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U801 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n617), .Z(n196) );
  MUX2_X1 U802 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n617), .Z(n197) );
  MUX2_X1 U803 ( .A(n197), .B(n196), .S(n608), .Z(n198) );
  MUX2_X1 U804 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n617), .Z(n199) );
  MUX2_X1 U805 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n617), .Z(n200) );
  MUX2_X1 U806 ( .A(n200), .B(n199), .S(n609), .Z(n201) );
  MUX2_X1 U807 ( .A(n201), .B(n198), .S(N12), .Z(n202) );
  MUX2_X1 U808 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n617), .Z(n203) );
  MUX2_X1 U809 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n617), .Z(n204) );
  MUX2_X1 U810 ( .A(n204), .B(n203), .S(n610), .Z(n205) );
  MUX2_X1 U811 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n617), .Z(n206) );
  MUX2_X1 U812 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n617), .Z(n207) );
  MUX2_X1 U813 ( .A(n207), .B(n206), .S(n610), .Z(n208) );
  MUX2_X1 U814 ( .A(n208), .B(n205), .S(n606), .Z(n209) );
  MUX2_X1 U815 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U816 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U817 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n617), .Z(n211) );
  MUX2_X1 U818 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n617), .Z(n212) );
  MUX2_X1 U819 ( .A(n212), .B(n211), .S(n610), .Z(n213) );
  MUX2_X1 U820 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n617), .Z(n214) );
  MUX2_X1 U821 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n617), .Z(n215) );
  MUX2_X1 U822 ( .A(n215), .B(n214), .S(n608), .Z(n216) );
  MUX2_X1 U823 ( .A(n216), .B(n213), .S(n606), .Z(n217) );
  MUX2_X1 U824 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n618), .Z(n218) );
  MUX2_X1 U825 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n618), .Z(n219) );
  MUX2_X1 U826 ( .A(n219), .B(n218), .S(n610), .Z(n220) );
  MUX2_X1 U827 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n618), .Z(n221) );
  MUX2_X1 U828 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n618), .Z(n222) );
  MUX2_X1 U829 ( .A(n222), .B(n221), .S(n608), .Z(n223) );
  MUX2_X1 U830 ( .A(n223), .B(n220), .S(n607), .Z(n224) );
  MUX2_X1 U831 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U832 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n618), .Z(n226) );
  MUX2_X1 U833 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n618), .Z(n227) );
  MUX2_X1 U834 ( .A(n227), .B(n226), .S(n609), .Z(n228) );
  MUX2_X1 U835 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n618), .Z(n229) );
  MUX2_X1 U836 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n618), .Z(n595) );
  MUX2_X1 U837 ( .A(n595), .B(n229), .S(n610), .Z(n596) );
  MUX2_X1 U838 ( .A(n596), .B(n228), .S(N12), .Z(n597) );
  MUX2_X1 U839 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n618), .Z(n598) );
  MUX2_X1 U840 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n618), .Z(n599) );
  MUX2_X1 U841 ( .A(n599), .B(n598), .S(n608), .Z(n600) );
  MUX2_X1 U842 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n618), .Z(n601) );
  MUX2_X1 U843 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n618), .Z(n602) );
  MUX2_X1 U844 ( .A(n602), .B(n601), .S(n608), .Z(n603) );
  MUX2_X1 U845 ( .A(n603), .B(n600), .S(n607), .Z(n604) );
  MUX2_X1 U846 ( .A(n604), .B(n597), .S(N13), .Z(n605) );
  MUX2_X1 U847 ( .A(n605), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U848 ( .A(N11), .Z(n608) );
  INV_X1 U849 ( .A(N10), .ZN(n620) );
  INV_X1 U850 ( .A(N11), .ZN(n621) );
  INV_X1 U851 ( .A(data_in[0]), .ZN(n622) );
  INV_X1 U852 ( .A(data_in[1]), .ZN(n623) );
  INV_X1 U853 ( .A(data_in[2]), .ZN(n624) );
  INV_X1 U854 ( .A(data_in[3]), .ZN(n625) );
  INV_X1 U855 ( .A(data_in[4]), .ZN(n626) );
  INV_X1 U856 ( .A(data_in[5]), .ZN(n627) );
  INV_X1 U857 ( .A(data_in[6]), .ZN(n628) );
  INV_X1 U858 ( .A(data_in[7]), .ZN(n629) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_29 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n629), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n630), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n631), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n632), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n633), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n634), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n635), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n636), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n637), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n638), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n639), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n640), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n641), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n642), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n643), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n644), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n645), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n646), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n647), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n648), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n649), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n650), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n651), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n652), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n653), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n654), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n655), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n656), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n657), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n658), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n659), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n660), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n661), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n662), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n663), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n664), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n665), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n666), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n667), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n668), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n669), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n670), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n671), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n672), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n673), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n674), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n675), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n676), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n677), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n678), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n679), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n680), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n681), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n682), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n683), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n684), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n685), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n686), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n687), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n688), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n689), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n690), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n691), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n692), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n693), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n694), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n695), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n696), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n697), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n698), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n699), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n700), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n701), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n702), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n703), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n704), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n705), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n706), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n707), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n708), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n709), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n710), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n711), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n712), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n713), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n714), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n715), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n716), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n717), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n718), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n719), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n720), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n721), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n722), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n723), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n724), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n725), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n726), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n727), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n728), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n729), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n730), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n731), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n732), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n733), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n734), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n735), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n736), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n737), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n738), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n739), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n740), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n741), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n742), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n743), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n744), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n745), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n746), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n747), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n748), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n749), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n750), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n751), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n752), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n753), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n754), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n755), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n756), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n757), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n758), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n759), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n760), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n761), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n762), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n763), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n764), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n765), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n766), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n767), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n768), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n769), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n770), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n771), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n772), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n773), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n774), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n775), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n776), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n777), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n778), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n779), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n780), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n781), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n782), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n783), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n784), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n785), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n786), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n787), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n788), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n789), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n790), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n791), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n792), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n793), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n794), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n795), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n796), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n797), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n798), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n799), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n800), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n801), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n802), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n803), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n804), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n805), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n806), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n807), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n808), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n809), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n810), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n811), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n812), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n813), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n814), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n815), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n816), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n817), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n818), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n819), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n820), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n848), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n849), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n850), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n851), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n852), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n853), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n854), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n855), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n856), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n857), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n858), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n859), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n860), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n861), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n862), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n863), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n864), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n865), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n866), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n867), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n868), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n869), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n870), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n871), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n872), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n873), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n874), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n875), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n876), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n877), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n878), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n879), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n880), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n881), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n882), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n883), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n884), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n885), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n886), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n887), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n888), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n889), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n890), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n891), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n892), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n893), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n894), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n895), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n896), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n897), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n898), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n899), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n900), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n901), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n902), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n903), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n904), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n905), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n906), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n907), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n908), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n909), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n910), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n911), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(n618), .Z(n616) );
  BUF_X1 U5 ( .A(n618), .Z(n617) );
  BUF_X1 U6 ( .A(N10), .Z(n614) );
  BUF_X1 U7 ( .A(n618), .Z(n615) );
  BUF_X1 U8 ( .A(N11), .Z(n611) );
  BUF_X1 U9 ( .A(N11), .Z(n612) );
  BUF_X1 U10 ( .A(N10), .Z(n618) );
  NOR3_X1 U11 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1203) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(n619), .ZN(n1192) );
  NOR3_X1 U13 ( .A1(N10), .A2(N12), .A3(n620), .ZN(n1182) );
  NOR3_X1 U14 ( .A1(n619), .A2(N12), .A3(n620), .ZN(n1172) );
  INV_X1 U15 ( .A(n1129), .ZN(n844) );
  INV_X1 U16 ( .A(n1119), .ZN(n843) );
  INV_X1 U17 ( .A(n1110), .ZN(n842) );
  INV_X1 U18 ( .A(n1101), .ZN(n841) );
  INV_X1 U19 ( .A(n1056), .ZN(n836) );
  INV_X1 U20 ( .A(n1046), .ZN(n835) );
  INV_X1 U21 ( .A(n1037), .ZN(n834) );
  INV_X1 U22 ( .A(n1028), .ZN(n833) );
  INV_X1 U23 ( .A(n983), .ZN(n828) );
  INV_X1 U24 ( .A(n973), .ZN(n827) );
  INV_X1 U25 ( .A(n964), .ZN(n826) );
  INV_X1 U26 ( .A(n955), .ZN(n825) );
  INV_X1 U27 ( .A(n1092), .ZN(n840) );
  INV_X1 U28 ( .A(n1083), .ZN(n839) );
  INV_X1 U29 ( .A(n1074), .ZN(n838) );
  INV_X1 U30 ( .A(n1065), .ZN(n837) );
  INV_X1 U31 ( .A(n946), .ZN(n824) );
  INV_X1 U32 ( .A(n937), .ZN(n823) );
  INV_X1 U33 ( .A(n928), .ZN(n822) );
  INV_X1 U34 ( .A(n919), .ZN(n821) );
  INV_X1 U35 ( .A(n1019), .ZN(n832) );
  INV_X1 U36 ( .A(n1010), .ZN(n831) );
  INV_X1 U37 ( .A(n1001), .ZN(n830) );
  INV_X1 U38 ( .A(n992), .ZN(n829) );
  BUF_X1 U39 ( .A(N12), .Z(n608) );
  BUF_X1 U40 ( .A(N12), .Z(n609) );
  INV_X1 U41 ( .A(N13), .ZN(n846) );
  AND3_X1 U42 ( .A1(n619), .A2(n620), .A3(N12), .ZN(n1162) );
  AND3_X1 U43 ( .A1(N10), .A2(n620), .A3(N12), .ZN(n1152) );
  AND3_X1 U44 ( .A1(N11), .A2(n619), .A3(N12), .ZN(n1142) );
  AND3_X1 U45 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1132) );
  INV_X1 U46 ( .A(N14), .ZN(n847) );
  NAND2_X1 U47 ( .A1(n1192), .A2(n1202), .ZN(n1201) );
  NAND2_X1 U48 ( .A1(n1182), .A2(n1202), .ZN(n1191) );
  NAND2_X1 U49 ( .A1(n1172), .A2(n1202), .ZN(n1181) );
  NAND2_X1 U50 ( .A1(n1162), .A2(n1202), .ZN(n1171) );
  NAND2_X1 U51 ( .A1(n1152), .A2(n1202), .ZN(n1161) );
  NAND2_X1 U52 ( .A1(n1142), .A2(n1202), .ZN(n1151) );
  NAND2_X1 U53 ( .A1(n1132), .A2(n1202), .ZN(n1141) );
  NAND2_X1 U54 ( .A1(n1203), .A2(n1202), .ZN(n1212) );
  NAND2_X1 U55 ( .A1(n1121), .A2(n1203), .ZN(n1129) );
  NAND2_X1 U56 ( .A1(n1121), .A2(n1192), .ZN(n1119) );
  NAND2_X1 U57 ( .A1(n1121), .A2(n1182), .ZN(n1110) );
  NAND2_X1 U58 ( .A1(n1121), .A2(n1172), .ZN(n1101) );
  NAND2_X1 U59 ( .A1(n1048), .A2(n1203), .ZN(n1056) );
  NAND2_X1 U60 ( .A1(n1048), .A2(n1192), .ZN(n1046) );
  NAND2_X1 U61 ( .A1(n1048), .A2(n1182), .ZN(n1037) );
  NAND2_X1 U62 ( .A1(n1048), .A2(n1172), .ZN(n1028) );
  NAND2_X1 U63 ( .A1(n975), .A2(n1203), .ZN(n983) );
  NAND2_X1 U64 ( .A1(n975), .A2(n1192), .ZN(n973) );
  NAND2_X1 U65 ( .A1(n975), .A2(n1182), .ZN(n964) );
  NAND2_X1 U66 ( .A1(n975), .A2(n1172), .ZN(n955) );
  NAND2_X1 U67 ( .A1(n1121), .A2(n1162), .ZN(n1092) );
  NAND2_X1 U68 ( .A1(n1121), .A2(n1152), .ZN(n1083) );
  NAND2_X1 U69 ( .A1(n1121), .A2(n1142), .ZN(n1074) );
  NAND2_X1 U70 ( .A1(n1121), .A2(n1132), .ZN(n1065) );
  NAND2_X1 U71 ( .A1(n1048), .A2(n1162), .ZN(n1019) );
  NAND2_X1 U72 ( .A1(n1048), .A2(n1152), .ZN(n1010) );
  NAND2_X1 U73 ( .A1(n1048), .A2(n1142), .ZN(n1001) );
  NAND2_X1 U74 ( .A1(n1048), .A2(n1132), .ZN(n992) );
  NAND2_X1 U75 ( .A1(n975), .A2(n1162), .ZN(n946) );
  NAND2_X1 U76 ( .A1(n975), .A2(n1152), .ZN(n937) );
  NAND2_X1 U77 ( .A1(n975), .A2(n1142), .ZN(n928) );
  NAND2_X1 U78 ( .A1(n975), .A2(n1132), .ZN(n919) );
  AND3_X1 U79 ( .A1(n846), .A2(n847), .A3(n1131), .ZN(n1202) );
  AND3_X1 U80 ( .A1(N13), .A2(n1131), .A3(N14), .ZN(n975) );
  AND3_X1 U81 ( .A1(n1131), .A2(n847), .A3(N13), .ZN(n1121) );
  AND3_X1 U82 ( .A1(n1131), .A2(n846), .A3(N14), .ZN(n1048) );
  NOR2_X1 U83 ( .A1(n845), .A2(addr[5]), .ZN(n1131) );
  INV_X1 U84 ( .A(wr_en), .ZN(n845) );
  OAI21_X1 U85 ( .B1(n621), .B2(n1171), .A(n1170), .ZN(n879) );
  NAND2_X1 U86 ( .A1(\mem[4][0] ), .A2(n1171), .ZN(n1170) );
  OAI21_X1 U87 ( .B1(n622), .B2(n1171), .A(n1169), .ZN(n878) );
  NAND2_X1 U88 ( .A1(\mem[4][1] ), .A2(n1171), .ZN(n1169) );
  OAI21_X1 U89 ( .B1(n623), .B2(n1171), .A(n1168), .ZN(n877) );
  NAND2_X1 U90 ( .A1(\mem[4][2] ), .A2(n1171), .ZN(n1168) );
  OAI21_X1 U91 ( .B1(n624), .B2(n1171), .A(n1167), .ZN(n876) );
  NAND2_X1 U92 ( .A1(\mem[4][3] ), .A2(n1171), .ZN(n1167) );
  OAI21_X1 U93 ( .B1(n625), .B2(n1171), .A(n1166), .ZN(n875) );
  NAND2_X1 U94 ( .A1(\mem[4][4] ), .A2(n1171), .ZN(n1166) );
  OAI21_X1 U95 ( .B1(n626), .B2(n1171), .A(n1165), .ZN(n874) );
  NAND2_X1 U96 ( .A1(\mem[4][5] ), .A2(n1171), .ZN(n1165) );
  OAI21_X1 U97 ( .B1(n627), .B2(n1171), .A(n1164), .ZN(n873) );
  NAND2_X1 U98 ( .A1(\mem[4][6] ), .A2(n1171), .ZN(n1164) );
  OAI21_X1 U99 ( .B1(n628), .B2(n1171), .A(n1163), .ZN(n872) );
  NAND2_X1 U100 ( .A1(\mem[4][7] ), .A2(n1171), .ZN(n1163) );
  OAI21_X1 U101 ( .B1(n621), .B2(n1151), .A(n1150), .ZN(n863) );
  NAND2_X1 U102 ( .A1(\mem[6][0] ), .A2(n1151), .ZN(n1150) );
  OAI21_X1 U103 ( .B1(n622), .B2(n1151), .A(n1149), .ZN(n862) );
  NAND2_X1 U104 ( .A1(\mem[6][1] ), .A2(n1151), .ZN(n1149) );
  OAI21_X1 U105 ( .B1(n623), .B2(n1151), .A(n1148), .ZN(n861) );
  NAND2_X1 U106 ( .A1(\mem[6][2] ), .A2(n1151), .ZN(n1148) );
  OAI21_X1 U107 ( .B1(n624), .B2(n1151), .A(n1147), .ZN(n860) );
  NAND2_X1 U108 ( .A1(\mem[6][3] ), .A2(n1151), .ZN(n1147) );
  OAI21_X1 U109 ( .B1(n625), .B2(n1151), .A(n1146), .ZN(n859) );
  NAND2_X1 U110 ( .A1(\mem[6][4] ), .A2(n1151), .ZN(n1146) );
  OAI21_X1 U111 ( .B1(n626), .B2(n1151), .A(n1145), .ZN(n858) );
  NAND2_X1 U112 ( .A1(\mem[6][5] ), .A2(n1151), .ZN(n1145) );
  OAI21_X1 U113 ( .B1(n627), .B2(n1151), .A(n1144), .ZN(n857) );
  NAND2_X1 U114 ( .A1(\mem[6][6] ), .A2(n1151), .ZN(n1144) );
  OAI21_X1 U115 ( .B1(n628), .B2(n1151), .A(n1143), .ZN(n856) );
  NAND2_X1 U116 ( .A1(\mem[6][7] ), .A2(n1151), .ZN(n1143) );
  OAI21_X1 U117 ( .B1(n621), .B2(n1141), .A(n1140), .ZN(n855) );
  NAND2_X1 U118 ( .A1(\mem[7][0] ), .A2(n1141), .ZN(n1140) );
  OAI21_X1 U119 ( .B1(n622), .B2(n1141), .A(n1139), .ZN(n854) );
  NAND2_X1 U120 ( .A1(\mem[7][1] ), .A2(n1141), .ZN(n1139) );
  OAI21_X1 U121 ( .B1(n623), .B2(n1141), .A(n1138), .ZN(n853) );
  NAND2_X1 U122 ( .A1(\mem[7][2] ), .A2(n1141), .ZN(n1138) );
  OAI21_X1 U123 ( .B1(n624), .B2(n1141), .A(n1137), .ZN(n852) );
  NAND2_X1 U124 ( .A1(\mem[7][3] ), .A2(n1141), .ZN(n1137) );
  OAI21_X1 U125 ( .B1(n625), .B2(n1141), .A(n1136), .ZN(n851) );
  NAND2_X1 U126 ( .A1(\mem[7][4] ), .A2(n1141), .ZN(n1136) );
  OAI21_X1 U127 ( .B1(n626), .B2(n1141), .A(n1135), .ZN(n850) );
  NAND2_X1 U128 ( .A1(\mem[7][5] ), .A2(n1141), .ZN(n1135) );
  OAI21_X1 U129 ( .B1(n627), .B2(n1141), .A(n1134), .ZN(n849) );
  NAND2_X1 U130 ( .A1(\mem[7][6] ), .A2(n1141), .ZN(n1134) );
  OAI21_X1 U131 ( .B1(n628), .B2(n1141), .A(n1133), .ZN(n848) );
  NAND2_X1 U132 ( .A1(\mem[7][7] ), .A2(n1141), .ZN(n1133) );
  OAI21_X1 U133 ( .B1(n621), .B2(n1201), .A(n1200), .ZN(n903) );
  NAND2_X1 U134 ( .A1(\mem[1][0] ), .A2(n1201), .ZN(n1200) );
  OAI21_X1 U135 ( .B1(n622), .B2(n1201), .A(n1199), .ZN(n902) );
  NAND2_X1 U136 ( .A1(\mem[1][1] ), .A2(n1201), .ZN(n1199) );
  OAI21_X1 U137 ( .B1(n623), .B2(n1201), .A(n1198), .ZN(n901) );
  NAND2_X1 U138 ( .A1(\mem[1][2] ), .A2(n1201), .ZN(n1198) );
  OAI21_X1 U139 ( .B1(n624), .B2(n1201), .A(n1197), .ZN(n900) );
  NAND2_X1 U140 ( .A1(\mem[1][3] ), .A2(n1201), .ZN(n1197) );
  OAI21_X1 U141 ( .B1(n625), .B2(n1201), .A(n1196), .ZN(n899) );
  NAND2_X1 U142 ( .A1(\mem[1][4] ), .A2(n1201), .ZN(n1196) );
  OAI21_X1 U143 ( .B1(n626), .B2(n1201), .A(n1195), .ZN(n898) );
  NAND2_X1 U144 ( .A1(\mem[1][5] ), .A2(n1201), .ZN(n1195) );
  OAI21_X1 U145 ( .B1(n627), .B2(n1201), .A(n1194), .ZN(n897) );
  NAND2_X1 U146 ( .A1(\mem[1][6] ), .A2(n1201), .ZN(n1194) );
  OAI21_X1 U147 ( .B1(n628), .B2(n1201), .A(n1193), .ZN(n896) );
  NAND2_X1 U148 ( .A1(\mem[1][7] ), .A2(n1201), .ZN(n1193) );
  OAI21_X1 U149 ( .B1(n621), .B2(n1191), .A(n1190), .ZN(n895) );
  NAND2_X1 U150 ( .A1(\mem[2][0] ), .A2(n1191), .ZN(n1190) );
  OAI21_X1 U151 ( .B1(n622), .B2(n1191), .A(n1189), .ZN(n894) );
  NAND2_X1 U152 ( .A1(\mem[2][1] ), .A2(n1191), .ZN(n1189) );
  OAI21_X1 U153 ( .B1(n623), .B2(n1191), .A(n1188), .ZN(n893) );
  NAND2_X1 U154 ( .A1(\mem[2][2] ), .A2(n1191), .ZN(n1188) );
  OAI21_X1 U155 ( .B1(n624), .B2(n1191), .A(n1187), .ZN(n892) );
  NAND2_X1 U156 ( .A1(\mem[2][3] ), .A2(n1191), .ZN(n1187) );
  OAI21_X1 U157 ( .B1(n625), .B2(n1191), .A(n1186), .ZN(n891) );
  NAND2_X1 U158 ( .A1(\mem[2][4] ), .A2(n1191), .ZN(n1186) );
  OAI21_X1 U159 ( .B1(n626), .B2(n1191), .A(n1185), .ZN(n890) );
  NAND2_X1 U160 ( .A1(\mem[2][5] ), .A2(n1191), .ZN(n1185) );
  OAI21_X1 U161 ( .B1(n627), .B2(n1191), .A(n1184), .ZN(n889) );
  NAND2_X1 U162 ( .A1(\mem[2][6] ), .A2(n1191), .ZN(n1184) );
  OAI21_X1 U163 ( .B1(n628), .B2(n1191), .A(n1183), .ZN(n888) );
  NAND2_X1 U164 ( .A1(\mem[2][7] ), .A2(n1191), .ZN(n1183) );
  OAI21_X1 U165 ( .B1(n621), .B2(n1181), .A(n1180), .ZN(n887) );
  NAND2_X1 U166 ( .A1(\mem[3][0] ), .A2(n1181), .ZN(n1180) );
  OAI21_X1 U167 ( .B1(n622), .B2(n1181), .A(n1179), .ZN(n886) );
  NAND2_X1 U168 ( .A1(\mem[3][1] ), .A2(n1181), .ZN(n1179) );
  OAI21_X1 U169 ( .B1(n623), .B2(n1181), .A(n1178), .ZN(n885) );
  NAND2_X1 U170 ( .A1(\mem[3][2] ), .A2(n1181), .ZN(n1178) );
  OAI21_X1 U171 ( .B1(n624), .B2(n1181), .A(n1177), .ZN(n884) );
  NAND2_X1 U172 ( .A1(\mem[3][3] ), .A2(n1181), .ZN(n1177) );
  OAI21_X1 U173 ( .B1(n625), .B2(n1181), .A(n1176), .ZN(n883) );
  NAND2_X1 U174 ( .A1(\mem[3][4] ), .A2(n1181), .ZN(n1176) );
  OAI21_X1 U175 ( .B1(n626), .B2(n1181), .A(n1175), .ZN(n882) );
  NAND2_X1 U176 ( .A1(\mem[3][5] ), .A2(n1181), .ZN(n1175) );
  OAI21_X1 U177 ( .B1(n627), .B2(n1181), .A(n1174), .ZN(n881) );
  NAND2_X1 U178 ( .A1(\mem[3][6] ), .A2(n1181), .ZN(n1174) );
  OAI21_X1 U179 ( .B1(n628), .B2(n1181), .A(n1173), .ZN(n880) );
  NAND2_X1 U180 ( .A1(\mem[3][7] ), .A2(n1181), .ZN(n1173) );
  OAI21_X1 U181 ( .B1(n621), .B2(n1161), .A(n1160), .ZN(n871) );
  NAND2_X1 U182 ( .A1(\mem[5][0] ), .A2(n1161), .ZN(n1160) );
  OAI21_X1 U183 ( .B1(n622), .B2(n1161), .A(n1159), .ZN(n870) );
  NAND2_X1 U184 ( .A1(\mem[5][1] ), .A2(n1161), .ZN(n1159) );
  OAI21_X1 U185 ( .B1(n623), .B2(n1161), .A(n1158), .ZN(n869) );
  NAND2_X1 U186 ( .A1(\mem[5][2] ), .A2(n1161), .ZN(n1158) );
  OAI21_X1 U187 ( .B1(n624), .B2(n1161), .A(n1157), .ZN(n868) );
  NAND2_X1 U188 ( .A1(\mem[5][3] ), .A2(n1161), .ZN(n1157) );
  OAI21_X1 U189 ( .B1(n625), .B2(n1161), .A(n1156), .ZN(n867) );
  NAND2_X1 U190 ( .A1(\mem[5][4] ), .A2(n1161), .ZN(n1156) );
  OAI21_X1 U191 ( .B1(n626), .B2(n1161), .A(n1155), .ZN(n866) );
  NAND2_X1 U192 ( .A1(\mem[5][5] ), .A2(n1161), .ZN(n1155) );
  OAI21_X1 U193 ( .B1(n627), .B2(n1161), .A(n1154), .ZN(n865) );
  NAND2_X1 U194 ( .A1(\mem[5][6] ), .A2(n1161), .ZN(n1154) );
  OAI21_X1 U195 ( .B1(n628), .B2(n1161), .A(n1153), .ZN(n864) );
  NAND2_X1 U196 ( .A1(\mem[5][7] ), .A2(n1161), .ZN(n1153) );
  OAI21_X1 U197 ( .B1(n1212), .B2(n621), .A(n1211), .ZN(n911) );
  NAND2_X1 U198 ( .A1(\mem[0][0] ), .A2(n1212), .ZN(n1211) );
  OAI21_X1 U199 ( .B1(n1212), .B2(n622), .A(n1210), .ZN(n910) );
  NAND2_X1 U200 ( .A1(\mem[0][1] ), .A2(n1212), .ZN(n1210) );
  OAI21_X1 U201 ( .B1(n1212), .B2(n623), .A(n1209), .ZN(n909) );
  NAND2_X1 U202 ( .A1(\mem[0][2] ), .A2(n1212), .ZN(n1209) );
  OAI21_X1 U203 ( .B1(n1212), .B2(n624), .A(n1208), .ZN(n908) );
  NAND2_X1 U204 ( .A1(\mem[0][3] ), .A2(n1212), .ZN(n1208) );
  OAI21_X1 U205 ( .B1(n1212), .B2(n625), .A(n1207), .ZN(n907) );
  NAND2_X1 U206 ( .A1(\mem[0][4] ), .A2(n1212), .ZN(n1207) );
  OAI21_X1 U207 ( .B1(n1212), .B2(n626), .A(n1206), .ZN(n906) );
  NAND2_X1 U208 ( .A1(\mem[0][5] ), .A2(n1212), .ZN(n1206) );
  OAI21_X1 U209 ( .B1(n1212), .B2(n627), .A(n1205), .ZN(n905) );
  NAND2_X1 U210 ( .A1(\mem[0][6] ), .A2(n1212), .ZN(n1205) );
  OAI21_X1 U211 ( .B1(n1212), .B2(n628), .A(n1204), .ZN(n904) );
  NAND2_X1 U212 ( .A1(\mem[0][7] ), .A2(n1212), .ZN(n1204) );
  INV_X1 U213 ( .A(n1130), .ZN(n820) );
  AOI22_X1 U214 ( .A1(data_in[0]), .A2(n844), .B1(n1129), .B2(\mem[8][0] ), 
        .ZN(n1130) );
  INV_X1 U215 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U216 ( .A1(data_in[1]), .A2(n844), .B1(n1129), .B2(\mem[8][1] ), 
        .ZN(n1128) );
  INV_X1 U217 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U218 ( .A1(data_in[2]), .A2(n844), .B1(n1129), .B2(\mem[8][2] ), 
        .ZN(n1127) );
  INV_X1 U219 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U220 ( .A1(data_in[3]), .A2(n844), .B1(n1129), .B2(\mem[8][3] ), 
        .ZN(n1126) );
  INV_X1 U221 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U222 ( .A1(data_in[4]), .A2(n844), .B1(n1129), .B2(\mem[8][4] ), 
        .ZN(n1125) );
  INV_X1 U223 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U224 ( .A1(data_in[5]), .A2(n844), .B1(n1129), .B2(\mem[8][5] ), 
        .ZN(n1124) );
  INV_X1 U225 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U226 ( .A1(data_in[6]), .A2(n844), .B1(n1129), .B2(\mem[8][6] ), 
        .ZN(n1123) );
  INV_X1 U227 ( .A(n1122), .ZN(n813) );
  AOI22_X1 U228 ( .A1(data_in[7]), .A2(n844), .B1(n1129), .B2(\mem[8][7] ), 
        .ZN(n1122) );
  INV_X1 U229 ( .A(n1120), .ZN(n812) );
  AOI22_X1 U230 ( .A1(data_in[0]), .A2(n843), .B1(n1119), .B2(\mem[9][0] ), 
        .ZN(n1120) );
  INV_X1 U231 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U232 ( .A1(data_in[1]), .A2(n843), .B1(n1119), .B2(\mem[9][1] ), 
        .ZN(n1118) );
  INV_X1 U233 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U234 ( .A1(data_in[2]), .A2(n843), .B1(n1119), .B2(\mem[9][2] ), 
        .ZN(n1117) );
  INV_X1 U235 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U236 ( .A1(data_in[3]), .A2(n843), .B1(n1119), .B2(\mem[9][3] ), 
        .ZN(n1116) );
  INV_X1 U237 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U238 ( .A1(data_in[4]), .A2(n843), .B1(n1119), .B2(\mem[9][4] ), 
        .ZN(n1115) );
  INV_X1 U239 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U240 ( .A1(data_in[5]), .A2(n843), .B1(n1119), .B2(\mem[9][5] ), 
        .ZN(n1114) );
  INV_X1 U241 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U242 ( .A1(data_in[6]), .A2(n843), .B1(n1119), .B2(\mem[9][6] ), 
        .ZN(n1113) );
  INV_X1 U243 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U244 ( .A1(data_in[7]), .A2(n843), .B1(n1119), .B2(\mem[9][7] ), 
        .ZN(n1112) );
  INV_X1 U245 ( .A(n1111), .ZN(n804) );
  AOI22_X1 U246 ( .A1(data_in[0]), .A2(n842), .B1(n1110), .B2(\mem[10][0] ), 
        .ZN(n1111) );
  INV_X1 U247 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U248 ( .A1(data_in[1]), .A2(n842), .B1(n1110), .B2(\mem[10][1] ), 
        .ZN(n1109) );
  INV_X1 U249 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U250 ( .A1(data_in[2]), .A2(n842), .B1(n1110), .B2(\mem[10][2] ), 
        .ZN(n1108) );
  INV_X1 U251 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U252 ( .A1(data_in[3]), .A2(n842), .B1(n1110), .B2(\mem[10][3] ), 
        .ZN(n1107) );
  INV_X1 U253 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U254 ( .A1(data_in[4]), .A2(n842), .B1(n1110), .B2(\mem[10][4] ), 
        .ZN(n1106) );
  INV_X1 U255 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U256 ( .A1(data_in[5]), .A2(n842), .B1(n1110), .B2(\mem[10][5] ), 
        .ZN(n1105) );
  INV_X1 U257 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U258 ( .A1(data_in[6]), .A2(n842), .B1(n1110), .B2(\mem[10][6] ), 
        .ZN(n1104) );
  INV_X1 U259 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U260 ( .A1(data_in[7]), .A2(n842), .B1(n1110), .B2(\mem[10][7] ), 
        .ZN(n1103) );
  INV_X1 U261 ( .A(n1102), .ZN(n796) );
  AOI22_X1 U262 ( .A1(data_in[0]), .A2(n841), .B1(n1101), .B2(\mem[11][0] ), 
        .ZN(n1102) );
  INV_X1 U263 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U264 ( .A1(data_in[1]), .A2(n841), .B1(n1101), .B2(\mem[11][1] ), 
        .ZN(n1100) );
  INV_X1 U265 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U266 ( .A1(data_in[2]), .A2(n841), .B1(n1101), .B2(\mem[11][2] ), 
        .ZN(n1099) );
  INV_X1 U267 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U268 ( .A1(data_in[3]), .A2(n841), .B1(n1101), .B2(\mem[11][3] ), 
        .ZN(n1098) );
  INV_X1 U269 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U270 ( .A1(data_in[4]), .A2(n841), .B1(n1101), .B2(\mem[11][4] ), 
        .ZN(n1097) );
  INV_X1 U271 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U272 ( .A1(data_in[5]), .A2(n841), .B1(n1101), .B2(\mem[11][5] ), 
        .ZN(n1096) );
  INV_X1 U273 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U274 ( .A1(data_in[6]), .A2(n841), .B1(n1101), .B2(\mem[11][6] ), 
        .ZN(n1095) );
  INV_X1 U275 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U276 ( .A1(data_in[7]), .A2(n841), .B1(n1101), .B2(\mem[11][7] ), 
        .ZN(n1094) );
  INV_X1 U277 ( .A(n1093), .ZN(n788) );
  AOI22_X1 U278 ( .A1(data_in[0]), .A2(n840), .B1(n1092), .B2(\mem[12][0] ), 
        .ZN(n1093) );
  INV_X1 U279 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U280 ( .A1(data_in[1]), .A2(n840), .B1(n1092), .B2(\mem[12][1] ), 
        .ZN(n1091) );
  INV_X1 U281 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U282 ( .A1(data_in[2]), .A2(n840), .B1(n1092), .B2(\mem[12][2] ), 
        .ZN(n1090) );
  INV_X1 U283 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U284 ( .A1(data_in[3]), .A2(n840), .B1(n1092), .B2(\mem[12][3] ), 
        .ZN(n1089) );
  INV_X1 U285 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U286 ( .A1(data_in[4]), .A2(n840), .B1(n1092), .B2(\mem[12][4] ), 
        .ZN(n1088) );
  INV_X1 U287 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U288 ( .A1(data_in[5]), .A2(n840), .B1(n1092), .B2(\mem[12][5] ), 
        .ZN(n1087) );
  INV_X1 U289 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U290 ( .A1(data_in[6]), .A2(n840), .B1(n1092), .B2(\mem[12][6] ), 
        .ZN(n1086) );
  INV_X1 U291 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U292 ( .A1(data_in[7]), .A2(n840), .B1(n1092), .B2(\mem[12][7] ), 
        .ZN(n1085) );
  INV_X1 U293 ( .A(n1084), .ZN(n780) );
  AOI22_X1 U294 ( .A1(data_in[0]), .A2(n839), .B1(n1083), .B2(\mem[13][0] ), 
        .ZN(n1084) );
  INV_X1 U295 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U296 ( .A1(data_in[1]), .A2(n839), .B1(n1083), .B2(\mem[13][1] ), 
        .ZN(n1082) );
  INV_X1 U297 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U298 ( .A1(data_in[2]), .A2(n839), .B1(n1083), .B2(\mem[13][2] ), 
        .ZN(n1081) );
  INV_X1 U299 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U300 ( .A1(data_in[3]), .A2(n839), .B1(n1083), .B2(\mem[13][3] ), 
        .ZN(n1080) );
  INV_X1 U301 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U302 ( .A1(data_in[4]), .A2(n839), .B1(n1083), .B2(\mem[13][4] ), 
        .ZN(n1079) );
  INV_X1 U303 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U304 ( .A1(data_in[5]), .A2(n839), .B1(n1083), .B2(\mem[13][5] ), 
        .ZN(n1078) );
  INV_X1 U305 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U306 ( .A1(data_in[6]), .A2(n839), .B1(n1083), .B2(\mem[13][6] ), 
        .ZN(n1077) );
  INV_X1 U307 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U308 ( .A1(data_in[7]), .A2(n839), .B1(n1083), .B2(\mem[13][7] ), 
        .ZN(n1076) );
  INV_X1 U309 ( .A(n1075), .ZN(n772) );
  AOI22_X1 U310 ( .A1(data_in[0]), .A2(n838), .B1(n1074), .B2(\mem[14][0] ), 
        .ZN(n1075) );
  INV_X1 U311 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U312 ( .A1(data_in[1]), .A2(n838), .B1(n1074), .B2(\mem[14][1] ), 
        .ZN(n1073) );
  INV_X1 U313 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U314 ( .A1(data_in[2]), .A2(n838), .B1(n1074), .B2(\mem[14][2] ), 
        .ZN(n1072) );
  INV_X1 U315 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U316 ( .A1(data_in[3]), .A2(n838), .B1(n1074), .B2(\mem[14][3] ), 
        .ZN(n1071) );
  INV_X1 U317 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U318 ( .A1(data_in[4]), .A2(n838), .B1(n1074), .B2(\mem[14][4] ), 
        .ZN(n1070) );
  INV_X1 U319 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U320 ( .A1(data_in[5]), .A2(n838), .B1(n1074), .B2(\mem[14][5] ), 
        .ZN(n1069) );
  INV_X1 U321 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U322 ( .A1(data_in[6]), .A2(n838), .B1(n1074), .B2(\mem[14][6] ), 
        .ZN(n1068) );
  INV_X1 U323 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U324 ( .A1(data_in[7]), .A2(n838), .B1(n1074), .B2(\mem[14][7] ), 
        .ZN(n1067) );
  INV_X1 U325 ( .A(n1066), .ZN(n764) );
  AOI22_X1 U326 ( .A1(data_in[0]), .A2(n837), .B1(n1065), .B2(\mem[15][0] ), 
        .ZN(n1066) );
  INV_X1 U327 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U328 ( .A1(data_in[1]), .A2(n837), .B1(n1065), .B2(\mem[15][1] ), 
        .ZN(n1064) );
  INV_X1 U329 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U330 ( .A1(data_in[2]), .A2(n837), .B1(n1065), .B2(\mem[15][2] ), 
        .ZN(n1063) );
  INV_X1 U331 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U332 ( .A1(data_in[3]), .A2(n837), .B1(n1065), .B2(\mem[15][3] ), 
        .ZN(n1062) );
  INV_X1 U333 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U334 ( .A1(data_in[4]), .A2(n837), .B1(n1065), .B2(\mem[15][4] ), 
        .ZN(n1061) );
  INV_X1 U335 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U336 ( .A1(data_in[5]), .A2(n837), .B1(n1065), .B2(\mem[15][5] ), 
        .ZN(n1060) );
  INV_X1 U337 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U338 ( .A1(data_in[6]), .A2(n837), .B1(n1065), .B2(\mem[15][6] ), 
        .ZN(n1059) );
  INV_X1 U339 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U340 ( .A1(data_in[7]), .A2(n837), .B1(n1065), .B2(\mem[15][7] ), 
        .ZN(n1058) );
  INV_X1 U341 ( .A(n1057), .ZN(n756) );
  AOI22_X1 U342 ( .A1(data_in[0]), .A2(n836), .B1(n1056), .B2(\mem[16][0] ), 
        .ZN(n1057) );
  INV_X1 U343 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U344 ( .A1(data_in[1]), .A2(n836), .B1(n1056), .B2(\mem[16][1] ), 
        .ZN(n1055) );
  INV_X1 U345 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U346 ( .A1(data_in[2]), .A2(n836), .B1(n1056), .B2(\mem[16][2] ), 
        .ZN(n1054) );
  INV_X1 U347 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U348 ( .A1(data_in[3]), .A2(n836), .B1(n1056), .B2(\mem[16][3] ), 
        .ZN(n1053) );
  INV_X1 U349 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U350 ( .A1(data_in[4]), .A2(n836), .B1(n1056), .B2(\mem[16][4] ), 
        .ZN(n1052) );
  INV_X1 U351 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U352 ( .A1(data_in[5]), .A2(n836), .B1(n1056), .B2(\mem[16][5] ), 
        .ZN(n1051) );
  INV_X1 U353 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U354 ( .A1(data_in[6]), .A2(n836), .B1(n1056), .B2(\mem[16][6] ), 
        .ZN(n1050) );
  INV_X1 U355 ( .A(n1049), .ZN(n749) );
  AOI22_X1 U356 ( .A1(data_in[7]), .A2(n836), .B1(n1056), .B2(\mem[16][7] ), 
        .ZN(n1049) );
  INV_X1 U357 ( .A(n1047), .ZN(n748) );
  AOI22_X1 U358 ( .A1(data_in[0]), .A2(n835), .B1(n1046), .B2(\mem[17][0] ), 
        .ZN(n1047) );
  INV_X1 U359 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U360 ( .A1(data_in[1]), .A2(n835), .B1(n1046), .B2(\mem[17][1] ), 
        .ZN(n1045) );
  INV_X1 U361 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U362 ( .A1(data_in[2]), .A2(n835), .B1(n1046), .B2(\mem[17][2] ), 
        .ZN(n1044) );
  INV_X1 U363 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U364 ( .A1(data_in[3]), .A2(n835), .B1(n1046), .B2(\mem[17][3] ), 
        .ZN(n1043) );
  INV_X1 U365 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U366 ( .A1(data_in[4]), .A2(n835), .B1(n1046), .B2(\mem[17][4] ), 
        .ZN(n1042) );
  INV_X1 U367 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U368 ( .A1(data_in[5]), .A2(n835), .B1(n1046), .B2(\mem[17][5] ), 
        .ZN(n1041) );
  INV_X1 U369 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U370 ( .A1(data_in[6]), .A2(n835), .B1(n1046), .B2(\mem[17][6] ), 
        .ZN(n1040) );
  INV_X1 U371 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U372 ( .A1(data_in[7]), .A2(n835), .B1(n1046), .B2(\mem[17][7] ), 
        .ZN(n1039) );
  INV_X1 U373 ( .A(n1038), .ZN(n740) );
  AOI22_X1 U374 ( .A1(data_in[0]), .A2(n834), .B1(n1037), .B2(\mem[18][0] ), 
        .ZN(n1038) );
  INV_X1 U375 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U376 ( .A1(data_in[1]), .A2(n834), .B1(n1037), .B2(\mem[18][1] ), 
        .ZN(n1036) );
  INV_X1 U377 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U378 ( .A1(data_in[2]), .A2(n834), .B1(n1037), .B2(\mem[18][2] ), 
        .ZN(n1035) );
  INV_X1 U379 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U380 ( .A1(data_in[3]), .A2(n834), .B1(n1037), .B2(\mem[18][3] ), 
        .ZN(n1034) );
  INV_X1 U381 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U382 ( .A1(data_in[4]), .A2(n834), .B1(n1037), .B2(\mem[18][4] ), 
        .ZN(n1033) );
  INV_X1 U383 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U384 ( .A1(data_in[5]), .A2(n834), .B1(n1037), .B2(\mem[18][5] ), 
        .ZN(n1032) );
  INV_X1 U385 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U386 ( .A1(data_in[6]), .A2(n834), .B1(n1037), .B2(\mem[18][6] ), 
        .ZN(n1031) );
  INV_X1 U387 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U388 ( .A1(data_in[7]), .A2(n834), .B1(n1037), .B2(\mem[18][7] ), 
        .ZN(n1030) );
  INV_X1 U389 ( .A(n1029), .ZN(n732) );
  AOI22_X1 U390 ( .A1(data_in[0]), .A2(n833), .B1(n1028), .B2(\mem[19][0] ), 
        .ZN(n1029) );
  INV_X1 U391 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U392 ( .A1(data_in[1]), .A2(n833), .B1(n1028), .B2(\mem[19][1] ), 
        .ZN(n1027) );
  INV_X1 U393 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U394 ( .A1(data_in[2]), .A2(n833), .B1(n1028), .B2(\mem[19][2] ), 
        .ZN(n1026) );
  INV_X1 U395 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U396 ( .A1(data_in[3]), .A2(n833), .B1(n1028), .B2(\mem[19][3] ), 
        .ZN(n1025) );
  INV_X1 U397 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U398 ( .A1(data_in[4]), .A2(n833), .B1(n1028), .B2(\mem[19][4] ), 
        .ZN(n1024) );
  INV_X1 U399 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U400 ( .A1(data_in[5]), .A2(n833), .B1(n1028), .B2(\mem[19][5] ), 
        .ZN(n1023) );
  INV_X1 U401 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U402 ( .A1(data_in[6]), .A2(n833), .B1(n1028), .B2(\mem[19][6] ), 
        .ZN(n1022) );
  INV_X1 U403 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U404 ( .A1(data_in[7]), .A2(n833), .B1(n1028), .B2(\mem[19][7] ), 
        .ZN(n1021) );
  INV_X1 U405 ( .A(n1020), .ZN(n724) );
  AOI22_X1 U406 ( .A1(data_in[0]), .A2(n832), .B1(n1019), .B2(\mem[20][0] ), 
        .ZN(n1020) );
  INV_X1 U407 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U408 ( .A1(data_in[1]), .A2(n832), .B1(n1019), .B2(\mem[20][1] ), 
        .ZN(n1018) );
  INV_X1 U409 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U410 ( .A1(data_in[2]), .A2(n832), .B1(n1019), .B2(\mem[20][2] ), 
        .ZN(n1017) );
  INV_X1 U411 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U412 ( .A1(data_in[3]), .A2(n832), .B1(n1019), .B2(\mem[20][3] ), 
        .ZN(n1016) );
  INV_X1 U413 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U414 ( .A1(data_in[4]), .A2(n832), .B1(n1019), .B2(\mem[20][4] ), 
        .ZN(n1015) );
  INV_X1 U415 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U416 ( .A1(data_in[5]), .A2(n832), .B1(n1019), .B2(\mem[20][5] ), 
        .ZN(n1014) );
  INV_X1 U417 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U418 ( .A1(data_in[6]), .A2(n832), .B1(n1019), .B2(\mem[20][6] ), 
        .ZN(n1013) );
  INV_X1 U419 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U420 ( .A1(data_in[7]), .A2(n832), .B1(n1019), .B2(\mem[20][7] ), 
        .ZN(n1012) );
  INV_X1 U421 ( .A(n1011), .ZN(n716) );
  AOI22_X1 U422 ( .A1(data_in[0]), .A2(n831), .B1(n1010), .B2(\mem[21][0] ), 
        .ZN(n1011) );
  INV_X1 U423 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U424 ( .A1(data_in[1]), .A2(n831), .B1(n1010), .B2(\mem[21][1] ), 
        .ZN(n1009) );
  INV_X1 U425 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U426 ( .A1(data_in[2]), .A2(n831), .B1(n1010), .B2(\mem[21][2] ), 
        .ZN(n1008) );
  INV_X1 U427 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U428 ( .A1(data_in[3]), .A2(n831), .B1(n1010), .B2(\mem[21][3] ), 
        .ZN(n1007) );
  INV_X1 U429 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U430 ( .A1(data_in[4]), .A2(n831), .B1(n1010), .B2(\mem[21][4] ), 
        .ZN(n1006) );
  INV_X1 U431 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U432 ( .A1(data_in[5]), .A2(n831), .B1(n1010), .B2(\mem[21][5] ), 
        .ZN(n1005) );
  INV_X1 U433 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U434 ( .A1(data_in[6]), .A2(n831), .B1(n1010), .B2(\mem[21][6] ), 
        .ZN(n1004) );
  INV_X1 U435 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U436 ( .A1(data_in[7]), .A2(n831), .B1(n1010), .B2(\mem[21][7] ), 
        .ZN(n1003) );
  INV_X1 U437 ( .A(n1002), .ZN(n708) );
  AOI22_X1 U438 ( .A1(data_in[0]), .A2(n830), .B1(n1001), .B2(\mem[22][0] ), 
        .ZN(n1002) );
  INV_X1 U439 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U440 ( .A1(data_in[1]), .A2(n830), .B1(n1001), .B2(\mem[22][1] ), 
        .ZN(n1000) );
  INV_X1 U441 ( .A(n999), .ZN(n706) );
  AOI22_X1 U442 ( .A1(data_in[2]), .A2(n830), .B1(n1001), .B2(\mem[22][2] ), 
        .ZN(n999) );
  INV_X1 U443 ( .A(n998), .ZN(n705) );
  AOI22_X1 U444 ( .A1(data_in[3]), .A2(n830), .B1(n1001), .B2(\mem[22][3] ), 
        .ZN(n998) );
  INV_X1 U445 ( .A(n997), .ZN(n704) );
  AOI22_X1 U446 ( .A1(data_in[4]), .A2(n830), .B1(n1001), .B2(\mem[22][4] ), 
        .ZN(n997) );
  INV_X1 U447 ( .A(n996), .ZN(n703) );
  AOI22_X1 U448 ( .A1(data_in[5]), .A2(n830), .B1(n1001), .B2(\mem[22][5] ), 
        .ZN(n996) );
  INV_X1 U449 ( .A(n995), .ZN(n702) );
  AOI22_X1 U450 ( .A1(data_in[6]), .A2(n830), .B1(n1001), .B2(\mem[22][6] ), 
        .ZN(n995) );
  INV_X1 U451 ( .A(n994), .ZN(n701) );
  AOI22_X1 U452 ( .A1(data_in[7]), .A2(n830), .B1(n1001), .B2(\mem[22][7] ), 
        .ZN(n994) );
  INV_X1 U453 ( .A(n993), .ZN(n700) );
  AOI22_X1 U454 ( .A1(data_in[0]), .A2(n829), .B1(n992), .B2(\mem[23][0] ), 
        .ZN(n993) );
  INV_X1 U455 ( .A(n991), .ZN(n699) );
  AOI22_X1 U456 ( .A1(data_in[1]), .A2(n829), .B1(n992), .B2(\mem[23][1] ), 
        .ZN(n991) );
  INV_X1 U457 ( .A(n990), .ZN(n698) );
  AOI22_X1 U458 ( .A1(data_in[2]), .A2(n829), .B1(n992), .B2(\mem[23][2] ), 
        .ZN(n990) );
  INV_X1 U459 ( .A(n989), .ZN(n697) );
  AOI22_X1 U460 ( .A1(data_in[3]), .A2(n829), .B1(n992), .B2(\mem[23][3] ), 
        .ZN(n989) );
  INV_X1 U461 ( .A(n988), .ZN(n696) );
  AOI22_X1 U462 ( .A1(data_in[4]), .A2(n829), .B1(n992), .B2(\mem[23][4] ), 
        .ZN(n988) );
  INV_X1 U463 ( .A(n987), .ZN(n695) );
  AOI22_X1 U464 ( .A1(data_in[5]), .A2(n829), .B1(n992), .B2(\mem[23][5] ), 
        .ZN(n987) );
  INV_X1 U465 ( .A(n986), .ZN(n694) );
  AOI22_X1 U466 ( .A1(data_in[6]), .A2(n829), .B1(n992), .B2(\mem[23][6] ), 
        .ZN(n986) );
  INV_X1 U467 ( .A(n985), .ZN(n693) );
  AOI22_X1 U468 ( .A1(data_in[7]), .A2(n829), .B1(n992), .B2(\mem[23][7] ), 
        .ZN(n985) );
  INV_X1 U469 ( .A(n984), .ZN(n692) );
  AOI22_X1 U470 ( .A1(data_in[0]), .A2(n828), .B1(n983), .B2(\mem[24][0] ), 
        .ZN(n984) );
  INV_X1 U471 ( .A(n982), .ZN(n691) );
  AOI22_X1 U472 ( .A1(data_in[1]), .A2(n828), .B1(n983), .B2(\mem[24][1] ), 
        .ZN(n982) );
  INV_X1 U473 ( .A(n981), .ZN(n690) );
  AOI22_X1 U474 ( .A1(data_in[2]), .A2(n828), .B1(n983), .B2(\mem[24][2] ), 
        .ZN(n981) );
  INV_X1 U475 ( .A(n980), .ZN(n689) );
  AOI22_X1 U476 ( .A1(data_in[3]), .A2(n828), .B1(n983), .B2(\mem[24][3] ), 
        .ZN(n980) );
  INV_X1 U477 ( .A(n979), .ZN(n688) );
  AOI22_X1 U478 ( .A1(data_in[4]), .A2(n828), .B1(n983), .B2(\mem[24][4] ), 
        .ZN(n979) );
  INV_X1 U479 ( .A(n978), .ZN(n687) );
  AOI22_X1 U480 ( .A1(data_in[5]), .A2(n828), .B1(n983), .B2(\mem[24][5] ), 
        .ZN(n978) );
  INV_X1 U481 ( .A(n977), .ZN(n686) );
  AOI22_X1 U482 ( .A1(data_in[6]), .A2(n828), .B1(n983), .B2(\mem[24][6] ), 
        .ZN(n977) );
  INV_X1 U483 ( .A(n976), .ZN(n685) );
  AOI22_X1 U484 ( .A1(data_in[7]), .A2(n828), .B1(n983), .B2(\mem[24][7] ), 
        .ZN(n976) );
  INV_X1 U485 ( .A(n974), .ZN(n684) );
  AOI22_X1 U486 ( .A1(data_in[0]), .A2(n827), .B1(n973), .B2(\mem[25][0] ), 
        .ZN(n974) );
  INV_X1 U487 ( .A(n972), .ZN(n683) );
  AOI22_X1 U488 ( .A1(data_in[1]), .A2(n827), .B1(n973), .B2(\mem[25][1] ), 
        .ZN(n972) );
  INV_X1 U489 ( .A(n971), .ZN(n682) );
  AOI22_X1 U490 ( .A1(data_in[2]), .A2(n827), .B1(n973), .B2(\mem[25][2] ), 
        .ZN(n971) );
  INV_X1 U491 ( .A(n970), .ZN(n681) );
  AOI22_X1 U492 ( .A1(data_in[3]), .A2(n827), .B1(n973), .B2(\mem[25][3] ), 
        .ZN(n970) );
  INV_X1 U493 ( .A(n969), .ZN(n680) );
  AOI22_X1 U494 ( .A1(data_in[4]), .A2(n827), .B1(n973), .B2(\mem[25][4] ), 
        .ZN(n969) );
  INV_X1 U495 ( .A(n968), .ZN(n679) );
  AOI22_X1 U496 ( .A1(data_in[5]), .A2(n827), .B1(n973), .B2(\mem[25][5] ), 
        .ZN(n968) );
  INV_X1 U497 ( .A(n967), .ZN(n678) );
  AOI22_X1 U498 ( .A1(data_in[6]), .A2(n827), .B1(n973), .B2(\mem[25][6] ), 
        .ZN(n967) );
  INV_X1 U499 ( .A(n966), .ZN(n677) );
  AOI22_X1 U500 ( .A1(data_in[7]), .A2(n827), .B1(n973), .B2(\mem[25][7] ), 
        .ZN(n966) );
  INV_X1 U501 ( .A(n965), .ZN(n676) );
  AOI22_X1 U502 ( .A1(data_in[0]), .A2(n826), .B1(n964), .B2(\mem[26][0] ), 
        .ZN(n965) );
  INV_X1 U503 ( .A(n963), .ZN(n675) );
  AOI22_X1 U504 ( .A1(data_in[1]), .A2(n826), .B1(n964), .B2(\mem[26][1] ), 
        .ZN(n963) );
  INV_X1 U505 ( .A(n962), .ZN(n674) );
  AOI22_X1 U506 ( .A1(data_in[2]), .A2(n826), .B1(n964), .B2(\mem[26][2] ), 
        .ZN(n962) );
  INV_X1 U507 ( .A(n961), .ZN(n673) );
  AOI22_X1 U508 ( .A1(data_in[3]), .A2(n826), .B1(n964), .B2(\mem[26][3] ), 
        .ZN(n961) );
  INV_X1 U509 ( .A(n960), .ZN(n672) );
  AOI22_X1 U510 ( .A1(data_in[4]), .A2(n826), .B1(n964), .B2(\mem[26][4] ), 
        .ZN(n960) );
  INV_X1 U511 ( .A(n959), .ZN(n671) );
  AOI22_X1 U512 ( .A1(data_in[5]), .A2(n826), .B1(n964), .B2(\mem[26][5] ), 
        .ZN(n959) );
  INV_X1 U513 ( .A(n958), .ZN(n670) );
  AOI22_X1 U514 ( .A1(data_in[6]), .A2(n826), .B1(n964), .B2(\mem[26][6] ), 
        .ZN(n958) );
  INV_X1 U515 ( .A(n957), .ZN(n669) );
  AOI22_X1 U516 ( .A1(data_in[7]), .A2(n826), .B1(n964), .B2(\mem[26][7] ), 
        .ZN(n957) );
  INV_X1 U517 ( .A(n956), .ZN(n668) );
  AOI22_X1 U518 ( .A1(data_in[0]), .A2(n825), .B1(n955), .B2(\mem[27][0] ), 
        .ZN(n956) );
  INV_X1 U519 ( .A(n954), .ZN(n667) );
  AOI22_X1 U520 ( .A1(data_in[1]), .A2(n825), .B1(n955), .B2(\mem[27][1] ), 
        .ZN(n954) );
  INV_X1 U521 ( .A(n953), .ZN(n666) );
  AOI22_X1 U522 ( .A1(data_in[2]), .A2(n825), .B1(n955), .B2(\mem[27][2] ), 
        .ZN(n953) );
  INV_X1 U523 ( .A(n952), .ZN(n665) );
  AOI22_X1 U524 ( .A1(data_in[3]), .A2(n825), .B1(n955), .B2(\mem[27][3] ), 
        .ZN(n952) );
  INV_X1 U525 ( .A(n951), .ZN(n664) );
  AOI22_X1 U526 ( .A1(data_in[4]), .A2(n825), .B1(n955), .B2(\mem[27][4] ), 
        .ZN(n951) );
  INV_X1 U527 ( .A(n950), .ZN(n663) );
  AOI22_X1 U528 ( .A1(data_in[5]), .A2(n825), .B1(n955), .B2(\mem[27][5] ), 
        .ZN(n950) );
  INV_X1 U529 ( .A(n949), .ZN(n662) );
  AOI22_X1 U530 ( .A1(data_in[6]), .A2(n825), .B1(n955), .B2(\mem[27][6] ), 
        .ZN(n949) );
  INV_X1 U531 ( .A(n948), .ZN(n661) );
  AOI22_X1 U532 ( .A1(data_in[7]), .A2(n825), .B1(n955), .B2(\mem[27][7] ), 
        .ZN(n948) );
  INV_X1 U533 ( .A(n947), .ZN(n660) );
  AOI22_X1 U534 ( .A1(data_in[0]), .A2(n824), .B1(n946), .B2(\mem[28][0] ), 
        .ZN(n947) );
  INV_X1 U535 ( .A(n945), .ZN(n659) );
  AOI22_X1 U536 ( .A1(data_in[1]), .A2(n824), .B1(n946), .B2(\mem[28][1] ), 
        .ZN(n945) );
  INV_X1 U537 ( .A(n944), .ZN(n658) );
  AOI22_X1 U538 ( .A1(data_in[2]), .A2(n824), .B1(n946), .B2(\mem[28][2] ), 
        .ZN(n944) );
  INV_X1 U539 ( .A(n943), .ZN(n657) );
  AOI22_X1 U540 ( .A1(data_in[3]), .A2(n824), .B1(n946), .B2(\mem[28][3] ), 
        .ZN(n943) );
  INV_X1 U541 ( .A(n942), .ZN(n656) );
  AOI22_X1 U542 ( .A1(data_in[4]), .A2(n824), .B1(n946), .B2(\mem[28][4] ), 
        .ZN(n942) );
  INV_X1 U543 ( .A(n941), .ZN(n655) );
  AOI22_X1 U544 ( .A1(data_in[5]), .A2(n824), .B1(n946), .B2(\mem[28][5] ), 
        .ZN(n941) );
  INV_X1 U545 ( .A(n940), .ZN(n654) );
  AOI22_X1 U546 ( .A1(data_in[6]), .A2(n824), .B1(n946), .B2(\mem[28][6] ), 
        .ZN(n940) );
  INV_X1 U547 ( .A(n939), .ZN(n653) );
  AOI22_X1 U548 ( .A1(data_in[7]), .A2(n824), .B1(n946), .B2(\mem[28][7] ), 
        .ZN(n939) );
  INV_X1 U549 ( .A(n938), .ZN(n652) );
  AOI22_X1 U550 ( .A1(data_in[0]), .A2(n823), .B1(n937), .B2(\mem[29][0] ), 
        .ZN(n938) );
  INV_X1 U551 ( .A(n936), .ZN(n651) );
  AOI22_X1 U552 ( .A1(data_in[1]), .A2(n823), .B1(n937), .B2(\mem[29][1] ), 
        .ZN(n936) );
  INV_X1 U553 ( .A(n935), .ZN(n650) );
  AOI22_X1 U554 ( .A1(data_in[2]), .A2(n823), .B1(n937), .B2(\mem[29][2] ), 
        .ZN(n935) );
  INV_X1 U555 ( .A(n934), .ZN(n649) );
  AOI22_X1 U556 ( .A1(data_in[3]), .A2(n823), .B1(n937), .B2(\mem[29][3] ), 
        .ZN(n934) );
  INV_X1 U557 ( .A(n933), .ZN(n648) );
  AOI22_X1 U558 ( .A1(data_in[4]), .A2(n823), .B1(n937), .B2(\mem[29][4] ), 
        .ZN(n933) );
  INV_X1 U559 ( .A(n932), .ZN(n647) );
  AOI22_X1 U560 ( .A1(data_in[5]), .A2(n823), .B1(n937), .B2(\mem[29][5] ), 
        .ZN(n932) );
  INV_X1 U561 ( .A(n931), .ZN(n646) );
  AOI22_X1 U562 ( .A1(data_in[6]), .A2(n823), .B1(n937), .B2(\mem[29][6] ), 
        .ZN(n931) );
  INV_X1 U563 ( .A(n930), .ZN(n645) );
  AOI22_X1 U564 ( .A1(data_in[7]), .A2(n823), .B1(n937), .B2(\mem[29][7] ), 
        .ZN(n930) );
  INV_X1 U565 ( .A(n929), .ZN(n644) );
  AOI22_X1 U566 ( .A1(data_in[0]), .A2(n822), .B1(n928), .B2(\mem[30][0] ), 
        .ZN(n929) );
  INV_X1 U567 ( .A(n927), .ZN(n643) );
  AOI22_X1 U568 ( .A1(data_in[1]), .A2(n822), .B1(n928), .B2(\mem[30][1] ), 
        .ZN(n927) );
  INV_X1 U569 ( .A(n926), .ZN(n642) );
  AOI22_X1 U570 ( .A1(data_in[2]), .A2(n822), .B1(n928), .B2(\mem[30][2] ), 
        .ZN(n926) );
  INV_X1 U571 ( .A(n925), .ZN(n641) );
  AOI22_X1 U572 ( .A1(data_in[3]), .A2(n822), .B1(n928), .B2(\mem[30][3] ), 
        .ZN(n925) );
  INV_X1 U573 ( .A(n924), .ZN(n640) );
  AOI22_X1 U574 ( .A1(data_in[4]), .A2(n822), .B1(n928), .B2(\mem[30][4] ), 
        .ZN(n924) );
  INV_X1 U575 ( .A(n923), .ZN(n639) );
  AOI22_X1 U576 ( .A1(data_in[5]), .A2(n822), .B1(n928), .B2(\mem[30][5] ), 
        .ZN(n923) );
  INV_X1 U577 ( .A(n922), .ZN(n638) );
  AOI22_X1 U578 ( .A1(data_in[6]), .A2(n822), .B1(n928), .B2(\mem[30][6] ), 
        .ZN(n922) );
  INV_X1 U579 ( .A(n921), .ZN(n637) );
  AOI22_X1 U580 ( .A1(data_in[7]), .A2(n822), .B1(n928), .B2(\mem[30][7] ), 
        .ZN(n921) );
  INV_X1 U581 ( .A(n920), .ZN(n636) );
  AOI22_X1 U582 ( .A1(data_in[0]), .A2(n821), .B1(n919), .B2(\mem[31][0] ), 
        .ZN(n920) );
  INV_X1 U583 ( .A(n918), .ZN(n635) );
  AOI22_X1 U584 ( .A1(data_in[1]), .A2(n821), .B1(n919), .B2(\mem[31][1] ), 
        .ZN(n918) );
  INV_X1 U585 ( .A(n917), .ZN(n634) );
  AOI22_X1 U586 ( .A1(data_in[2]), .A2(n821), .B1(n919), .B2(\mem[31][2] ), 
        .ZN(n917) );
  INV_X1 U587 ( .A(n916), .ZN(n633) );
  AOI22_X1 U588 ( .A1(data_in[3]), .A2(n821), .B1(n919), .B2(\mem[31][3] ), 
        .ZN(n916) );
  INV_X1 U589 ( .A(n915), .ZN(n632) );
  AOI22_X1 U590 ( .A1(data_in[4]), .A2(n821), .B1(n919), .B2(\mem[31][4] ), 
        .ZN(n915) );
  INV_X1 U591 ( .A(n914), .ZN(n631) );
  AOI22_X1 U592 ( .A1(data_in[5]), .A2(n821), .B1(n919), .B2(\mem[31][5] ), 
        .ZN(n914) );
  INV_X1 U593 ( .A(n913), .ZN(n630) );
  AOI22_X1 U594 ( .A1(data_in[6]), .A2(n821), .B1(n919), .B2(\mem[31][6] ), 
        .ZN(n913) );
  INV_X1 U595 ( .A(n912), .ZN(n629) );
  AOI22_X1 U596 ( .A1(data_in[7]), .A2(n821), .B1(n919), .B2(\mem[31][7] ), 
        .ZN(n912) );
  MUX2_X1 U597 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n613), .Z(n3) );
  MUX2_X1 U598 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n613), .Z(n4) );
  MUX2_X1 U599 ( .A(n4), .B(n3), .S(n610), .Z(n5) );
  MUX2_X1 U600 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n613), .Z(n6) );
  MUX2_X1 U601 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n613), .Z(n7) );
  MUX2_X1 U602 ( .A(n7), .B(n6), .S(n610), .Z(n8) );
  MUX2_X1 U603 ( .A(n8), .B(n5), .S(N12), .Z(n9) );
  MUX2_X1 U604 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n613), .Z(n10) );
  MUX2_X1 U605 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n613), .Z(n11) );
  MUX2_X1 U606 ( .A(n11), .B(n10), .S(n610), .Z(n12) );
  MUX2_X1 U607 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n613), .Z(n13) );
  MUX2_X1 U608 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n613), .Z(n14) );
  MUX2_X1 U609 ( .A(n14), .B(n13), .S(n610), .Z(n15) );
  MUX2_X1 U610 ( .A(n15), .B(n12), .S(n608), .Z(n16) );
  MUX2_X1 U611 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U612 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n614), .Z(n18) );
  MUX2_X1 U613 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n615), .Z(n19) );
  MUX2_X1 U614 ( .A(n19), .B(n18), .S(n610), .Z(n20) );
  MUX2_X1 U615 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n618), .Z(n21) );
  MUX2_X1 U616 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n22) );
  MUX2_X1 U617 ( .A(n22), .B(n21), .S(N11), .Z(n23) );
  MUX2_X1 U618 ( .A(n23), .B(n20), .S(n609), .Z(n24) );
  MUX2_X1 U619 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n613), .Z(n25) );
  MUX2_X1 U620 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n26) );
  MUX2_X1 U621 ( .A(n26), .B(n25), .S(N11), .Z(n27) );
  MUX2_X1 U622 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n28) );
  MUX2_X1 U623 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n29) );
  MUX2_X1 U624 ( .A(n29), .B(n28), .S(n612), .Z(n30) );
  MUX2_X1 U625 ( .A(n30), .B(n27), .S(n609), .Z(n31) );
  MUX2_X1 U626 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U627 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U628 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n613), .Z(n33) );
  MUX2_X1 U629 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n613), .Z(n34) );
  MUX2_X1 U630 ( .A(n34), .B(n33), .S(n611), .Z(n35) );
  MUX2_X1 U631 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n613), .Z(n36) );
  MUX2_X1 U632 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n613), .Z(n37) );
  MUX2_X1 U633 ( .A(n37), .B(n36), .S(N11), .Z(n38) );
  MUX2_X1 U634 ( .A(n38), .B(n35), .S(N12), .Z(n39) );
  MUX2_X1 U635 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n618), .Z(n40) );
  MUX2_X1 U636 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n616), .Z(n41) );
  MUX2_X1 U637 ( .A(n41), .B(n40), .S(n611), .Z(n42) );
  MUX2_X1 U638 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n618), .Z(n43) );
  MUX2_X1 U639 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n614), .Z(n44) );
  MUX2_X1 U640 ( .A(n44), .B(n43), .S(n610), .Z(n45) );
  MUX2_X1 U641 ( .A(n45), .B(n42), .S(n609), .Z(n46) );
  MUX2_X1 U642 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U643 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n615), .Z(n48) );
  MUX2_X1 U644 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n618), .Z(n49) );
  MUX2_X1 U645 ( .A(n49), .B(n48), .S(n612), .Z(n50) );
  MUX2_X1 U646 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n618), .Z(n51) );
  MUX2_X1 U647 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n618), .Z(n52) );
  MUX2_X1 U648 ( .A(n52), .B(n51), .S(n612), .Z(n53) );
  MUX2_X1 U649 ( .A(n53), .B(n50), .S(n608), .Z(n54) );
  MUX2_X1 U650 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n617), .Z(n55) );
  MUX2_X1 U651 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n56) );
  MUX2_X1 U652 ( .A(n56), .B(n55), .S(N11), .Z(n57) );
  MUX2_X1 U653 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n614), .Z(n58) );
  MUX2_X1 U654 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n617), .Z(n59) );
  MUX2_X1 U655 ( .A(n59), .B(n58), .S(n611), .Z(n60) );
  MUX2_X1 U656 ( .A(n60), .B(n57), .S(N12), .Z(n61) );
  MUX2_X1 U657 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U658 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U659 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n614), .Z(n63) );
  MUX2_X1 U660 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n614), .Z(n64) );
  MUX2_X1 U661 ( .A(n64), .B(n63), .S(n610), .Z(n65) );
  MUX2_X1 U662 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n614), .Z(n66) );
  MUX2_X1 U663 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n614), .Z(n67) );
  MUX2_X1 U664 ( .A(n67), .B(n66), .S(n610), .Z(n68) );
  MUX2_X1 U665 ( .A(n68), .B(n65), .S(n608), .Z(n69) );
  MUX2_X1 U666 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n614), .Z(n70) );
  MUX2_X1 U667 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n614), .Z(n71) );
  MUX2_X1 U668 ( .A(n71), .B(n70), .S(n610), .Z(n72) );
  MUX2_X1 U669 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n614), .Z(n73) );
  MUX2_X1 U670 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n614), .Z(n74) );
  MUX2_X1 U671 ( .A(n74), .B(n73), .S(n610), .Z(n75) );
  MUX2_X1 U672 ( .A(n75), .B(n72), .S(n608), .Z(n76) );
  MUX2_X1 U673 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U674 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n614), .Z(n78) );
  MUX2_X1 U675 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n614), .Z(n79) );
  MUX2_X1 U676 ( .A(n79), .B(n78), .S(n610), .Z(n80) );
  MUX2_X1 U677 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n614), .Z(n81) );
  MUX2_X1 U678 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n614), .Z(n82) );
  MUX2_X1 U679 ( .A(n82), .B(n81), .S(n612), .Z(n83) );
  MUX2_X1 U680 ( .A(n83), .B(n80), .S(n608), .Z(n84) );
  MUX2_X1 U681 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n615), .Z(n85) );
  MUX2_X1 U682 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n615), .Z(n86) );
  MUX2_X1 U683 ( .A(n86), .B(n85), .S(n611), .Z(n87) );
  MUX2_X1 U684 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n615), .Z(n88) );
  MUX2_X1 U685 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n615), .Z(n89) );
  MUX2_X1 U686 ( .A(n89), .B(n88), .S(n610), .Z(n90) );
  MUX2_X1 U687 ( .A(n90), .B(n87), .S(n608), .Z(n91) );
  MUX2_X1 U688 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U689 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U690 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n615), .Z(n93) );
  MUX2_X1 U691 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n615), .Z(n94) );
  MUX2_X1 U692 ( .A(n94), .B(n93), .S(n610), .Z(n95) );
  MUX2_X1 U693 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n615), .Z(n96) );
  MUX2_X1 U694 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n615), .Z(n97) );
  MUX2_X1 U695 ( .A(n97), .B(n96), .S(n610), .Z(n98) );
  MUX2_X1 U696 ( .A(n98), .B(n95), .S(n608), .Z(n99) );
  MUX2_X1 U697 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n615), .Z(n100) );
  MUX2_X1 U698 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n615), .Z(n101) );
  MUX2_X1 U699 ( .A(n101), .B(n100), .S(n610), .Z(n102) );
  MUX2_X1 U700 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n615), .Z(n103) );
  MUX2_X1 U701 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n615), .Z(n104) );
  MUX2_X1 U702 ( .A(n104), .B(n103), .S(n612), .Z(n105) );
  MUX2_X1 U703 ( .A(n105), .B(n102), .S(n608), .Z(n106) );
  MUX2_X1 U704 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U705 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n618), .Z(n108) );
  MUX2_X1 U706 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n618), .Z(n109) );
  MUX2_X1 U707 ( .A(n109), .B(n108), .S(n611), .Z(n110) );
  MUX2_X1 U708 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n618), .Z(n111) );
  MUX2_X1 U709 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n618), .Z(n112) );
  MUX2_X1 U710 ( .A(n112), .B(n111), .S(n611), .Z(n113) );
  MUX2_X1 U711 ( .A(n113), .B(n110), .S(n608), .Z(n114) );
  MUX2_X1 U712 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n618), .Z(n115) );
  MUX2_X1 U713 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n618), .Z(n116) );
  MUX2_X1 U714 ( .A(n116), .B(n115), .S(n611), .Z(n117) );
  MUX2_X1 U715 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n618), .Z(n118) );
  MUX2_X1 U716 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n618), .Z(n119) );
  MUX2_X1 U717 ( .A(n119), .B(n118), .S(n611), .Z(n120) );
  MUX2_X1 U718 ( .A(n120), .B(n117), .S(n608), .Z(n121) );
  MUX2_X1 U719 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U720 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U721 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n615), .Z(n123) );
  MUX2_X1 U722 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n618), .Z(n124) );
  MUX2_X1 U723 ( .A(n124), .B(n123), .S(n611), .Z(n125) );
  MUX2_X1 U724 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n615), .Z(n126) );
  MUX2_X1 U725 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n618), .Z(n127) );
  MUX2_X1 U726 ( .A(n127), .B(n126), .S(n611), .Z(n128) );
  MUX2_X1 U727 ( .A(n128), .B(n125), .S(n608), .Z(n129) );
  MUX2_X1 U728 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n614), .Z(n130) );
  MUX2_X1 U729 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n618), .Z(n131) );
  MUX2_X1 U730 ( .A(n131), .B(n130), .S(n611), .Z(n132) );
  MUX2_X1 U731 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n613), .Z(n133) );
  MUX2_X1 U732 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n613), .Z(n134) );
  MUX2_X1 U733 ( .A(n134), .B(n133), .S(n611), .Z(n135) );
  MUX2_X1 U734 ( .A(n135), .B(n132), .S(n608), .Z(n136) );
  MUX2_X1 U735 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U736 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n613), .Z(n138) );
  MUX2_X1 U737 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n616), .Z(n139) );
  MUX2_X1 U738 ( .A(n139), .B(n138), .S(n611), .Z(n140) );
  MUX2_X1 U739 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n614), .Z(n141) );
  MUX2_X1 U740 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n618), .Z(n142) );
  MUX2_X1 U741 ( .A(n142), .B(n141), .S(n611), .Z(n143) );
  MUX2_X1 U742 ( .A(n143), .B(n140), .S(n608), .Z(n144) );
  MUX2_X1 U743 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n613), .Z(n145) );
  MUX2_X1 U744 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n618), .Z(n146) );
  MUX2_X1 U745 ( .A(n146), .B(n145), .S(n611), .Z(n147) );
  MUX2_X1 U746 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n616), .Z(n148) );
  MUX2_X1 U747 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n618), .Z(n149) );
  MUX2_X1 U748 ( .A(n149), .B(n148), .S(n611), .Z(n150) );
  MUX2_X1 U749 ( .A(n150), .B(n147), .S(n608), .Z(n151) );
  MUX2_X1 U750 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U751 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U752 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n614), .Z(n153) );
  MUX2_X1 U753 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n614), .Z(n154) );
  MUX2_X1 U754 ( .A(n154), .B(n153), .S(n612), .Z(n155) );
  MUX2_X1 U755 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n613), .Z(n156) );
  MUX2_X1 U756 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n613), .Z(n157) );
  MUX2_X1 U757 ( .A(n157), .B(n156), .S(n612), .Z(n158) );
  MUX2_X1 U758 ( .A(n158), .B(n155), .S(n609), .Z(n159) );
  MUX2_X1 U759 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n613), .Z(n160) );
  MUX2_X1 U760 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n613), .Z(n161) );
  MUX2_X1 U761 ( .A(n161), .B(n160), .S(n612), .Z(n162) );
  MUX2_X1 U762 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n614), .Z(n163) );
  MUX2_X1 U763 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n613), .Z(n164) );
  MUX2_X1 U764 ( .A(n164), .B(n163), .S(n612), .Z(n165) );
  MUX2_X1 U765 ( .A(n165), .B(n162), .S(n609), .Z(n166) );
  MUX2_X1 U766 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U767 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n614), .Z(n168) );
  MUX2_X1 U768 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n614), .Z(n169) );
  MUX2_X1 U769 ( .A(n169), .B(n168), .S(n612), .Z(n170) );
  MUX2_X1 U770 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n613), .Z(n171) );
  MUX2_X1 U771 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n614), .Z(n172) );
  MUX2_X1 U772 ( .A(n172), .B(n171), .S(n612), .Z(n173) );
  MUX2_X1 U773 ( .A(n173), .B(n170), .S(n609), .Z(n174) );
  MUX2_X1 U774 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n616), .Z(n175) );
  MUX2_X1 U775 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n616), .Z(n176) );
  MUX2_X1 U776 ( .A(n176), .B(n175), .S(n612), .Z(n177) );
  MUX2_X1 U777 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n616), .Z(n178) );
  MUX2_X1 U778 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n616), .Z(n179) );
  MUX2_X1 U779 ( .A(n179), .B(n178), .S(n612), .Z(n180) );
  MUX2_X1 U780 ( .A(n180), .B(n177), .S(n609), .Z(n181) );
  MUX2_X1 U781 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U782 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U783 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n616), .Z(n183) );
  MUX2_X1 U784 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n616), .Z(n184) );
  MUX2_X1 U785 ( .A(n184), .B(n183), .S(n612), .Z(n185) );
  MUX2_X1 U786 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n616), .Z(n186) );
  MUX2_X1 U787 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n616), .Z(n187) );
  MUX2_X1 U788 ( .A(n187), .B(n186), .S(n612), .Z(n188) );
  MUX2_X1 U789 ( .A(n188), .B(n185), .S(n609), .Z(n189) );
  MUX2_X1 U790 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n616), .Z(n190) );
  MUX2_X1 U791 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n616), .Z(n191) );
  MUX2_X1 U792 ( .A(n191), .B(n190), .S(n612), .Z(n192) );
  MUX2_X1 U793 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n616), .Z(n193) );
  MUX2_X1 U794 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n616), .Z(n194) );
  MUX2_X1 U795 ( .A(n194), .B(n193), .S(n612), .Z(n195) );
  MUX2_X1 U796 ( .A(n195), .B(n192), .S(n609), .Z(n196) );
  MUX2_X1 U797 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U798 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n617), .Z(n198) );
  MUX2_X1 U799 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n617), .Z(n199) );
  MUX2_X1 U800 ( .A(n199), .B(n198), .S(n611), .Z(n200) );
  MUX2_X1 U801 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n617), .Z(n201) );
  MUX2_X1 U802 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n617), .Z(n202) );
  MUX2_X1 U803 ( .A(n202), .B(n201), .S(n612), .Z(n203) );
  MUX2_X1 U804 ( .A(n203), .B(n200), .S(n609), .Z(n204) );
  MUX2_X1 U805 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n617), .Z(n205) );
  MUX2_X1 U806 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n617), .Z(n206) );
  MUX2_X1 U807 ( .A(n206), .B(n205), .S(n611), .Z(n207) );
  MUX2_X1 U808 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n617), .Z(n208) );
  MUX2_X1 U809 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n617), .Z(n209) );
  MUX2_X1 U810 ( .A(n209), .B(n208), .S(n610), .Z(n210) );
  MUX2_X1 U811 ( .A(n210), .B(n207), .S(n609), .Z(n211) );
  MUX2_X1 U812 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U813 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U814 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n617), .Z(n213) );
  MUX2_X1 U815 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n617), .Z(n214) );
  MUX2_X1 U816 ( .A(n214), .B(n213), .S(n612), .Z(n215) );
  MUX2_X1 U817 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n617), .Z(n216) );
  MUX2_X1 U818 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n617), .Z(n217) );
  MUX2_X1 U819 ( .A(n217), .B(n216), .S(n612), .Z(n218) );
  MUX2_X1 U820 ( .A(n218), .B(n215), .S(n609), .Z(n219) );
  MUX2_X1 U821 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n617), .Z(n220) );
  MUX2_X1 U822 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n616), .Z(n221) );
  MUX2_X1 U823 ( .A(n221), .B(n220), .S(N11), .Z(n222) );
  MUX2_X1 U824 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n615), .Z(n223) );
  MUX2_X1 U825 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n616), .Z(n224) );
  MUX2_X1 U826 ( .A(n224), .B(n223), .S(n611), .Z(n225) );
  MUX2_X1 U827 ( .A(n225), .B(n222), .S(n609), .Z(n226) );
  MUX2_X1 U828 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U829 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n618), .Z(n228) );
  MUX2_X1 U830 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n617), .Z(n229) );
  MUX2_X1 U831 ( .A(n229), .B(n228), .S(n610), .Z(n595) );
  MUX2_X1 U832 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n617), .Z(n596) );
  MUX2_X1 U833 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n615), .Z(n597) );
  MUX2_X1 U834 ( .A(n597), .B(n596), .S(n611), .Z(n598) );
  MUX2_X1 U835 ( .A(n598), .B(n595), .S(n609), .Z(n599) );
  MUX2_X1 U836 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n616), .Z(n600) );
  MUX2_X1 U837 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n616), .Z(n601) );
  MUX2_X1 U838 ( .A(n601), .B(n600), .S(n610), .Z(n602) );
  MUX2_X1 U839 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n617), .Z(n603) );
  MUX2_X1 U840 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n617), .Z(n604) );
  MUX2_X1 U841 ( .A(n604), .B(n603), .S(n612), .Z(n605) );
  MUX2_X1 U842 ( .A(n605), .B(n602), .S(n609), .Z(n606) );
  MUX2_X1 U843 ( .A(n606), .B(n599), .S(N13), .Z(n607) );
  MUX2_X1 U844 ( .A(n607), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U845 ( .A(N11), .Z(n610) );
  CLKBUF_X1 U846 ( .A(N10), .Z(n613) );
  INV_X1 U847 ( .A(N10), .ZN(n619) );
  INV_X1 U848 ( .A(N11), .ZN(n620) );
  INV_X1 U849 ( .A(data_in[0]), .ZN(n621) );
  INV_X1 U850 ( .A(data_in[1]), .ZN(n622) );
  INV_X1 U851 ( .A(data_in[2]), .ZN(n623) );
  INV_X1 U852 ( .A(data_in[3]), .ZN(n624) );
  INV_X1 U853 ( .A(data_in[4]), .ZN(n625) );
  INV_X1 U854 ( .A(data_in[5]), .ZN(n626) );
  INV_X1 U855 ( .A(data_in[6]), .ZN(n627) );
  INV_X1 U856 ( .A(data_in[7]), .ZN(n628) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_28 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n628), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n629), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n630), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n631), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n632), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n633), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n634), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n635), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n636), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n637), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n638), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n639), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n640), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n641), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n642), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n643), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n644), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n645), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n646), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n647), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n648), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n649), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n650), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n651), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n652), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n653), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n654), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n655), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n656), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n657), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n658), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n659), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n660), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n661), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n662), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n663), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n664), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n665), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n666), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n667), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n668), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n669), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n670), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n671), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n672), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n673), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n674), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n675), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n676), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n677), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n678), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n679), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n680), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n681), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n682), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n683), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n684), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n685), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n686), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n687), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n688), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n689), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n690), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n691), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n692), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n693), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n694), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n695), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n696), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n697), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n698), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n699), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n700), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n701), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n702), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n703), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n704), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n705), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n706), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n707), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n708), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n709), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n710), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n711), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n712), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n713), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n714), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n715), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n716), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n717), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n718), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n719), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n720), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n721), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n722), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n723), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n724), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n725), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n726), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n727), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n728), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n729), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n730), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n731), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n732), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n733), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n734), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n735), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n736), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n737), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n738), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n739), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n740), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n741), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n742), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n743), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n744), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n745), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n746), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n747), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n748), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n749), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n750), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n751), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n752), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n753), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n754), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n755), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n756), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n757), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n758), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n759), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n760), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n761), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n762), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n763), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n764), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n765), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n766), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n767), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n768), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n769), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n770), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n771), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n772), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n773), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n774), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n775), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n776), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n777), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n778), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n779), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n780), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n781), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n782), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n783), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n784), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n785), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n786), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n787), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n788), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n789), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n790), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n791), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n792), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n793), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n794), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n795), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n796), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n797), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n798), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n799), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n800), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n801), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n802), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n803), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n804), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n805), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n806), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n807), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n808), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n809), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n810), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n811), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n812), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n813), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n814), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n815), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n816), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n817), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n818), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n819), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n847), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n848), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n849), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n850), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n851), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n852), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n853), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n854), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n855), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n856), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n857), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n858), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n859), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n860), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n861), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n862), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n863), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n864), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n865), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n866), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n867), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n868), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n869), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n870), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n871), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n872), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n873), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n874), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n875), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n876), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n877), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n878), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n879), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n880), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n881), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n882), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n883), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n884), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n885), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n886), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n887), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n888), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n889), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n890), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n891), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n892), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n893), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n894), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n895), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n896), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n897), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n898), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n899), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n900), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n901), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n902), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n903), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n904), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n905), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n906), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n907), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n908), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n909), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n910), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n617), .Z(n615) );
  BUF_X1 U4 ( .A(n617), .Z(n616) );
  BUF_X1 U5 ( .A(N10), .Z(n612) );
  BUF_X1 U6 ( .A(N10), .Z(n613) );
  BUF_X1 U7 ( .A(n617), .Z(n614) );
  BUF_X1 U8 ( .A(N11), .Z(n609) );
  BUF_X1 U9 ( .A(N11), .Z(n610) );
  BUF_X1 U10 ( .A(N10), .Z(n617) );
  NOR3_X1 U11 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1202) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(n618), .ZN(n1191) );
  NOR3_X1 U13 ( .A1(N10), .A2(N12), .A3(n619), .ZN(n1181) );
  NOR3_X1 U14 ( .A1(n618), .A2(N12), .A3(n619), .ZN(n1171) );
  INV_X1 U15 ( .A(n1128), .ZN(n843) );
  INV_X1 U16 ( .A(n1118), .ZN(n842) );
  INV_X1 U17 ( .A(n1109), .ZN(n841) );
  INV_X1 U18 ( .A(n1100), .ZN(n840) );
  INV_X1 U19 ( .A(n1055), .ZN(n835) );
  INV_X1 U20 ( .A(n1045), .ZN(n834) );
  INV_X1 U21 ( .A(n1036), .ZN(n833) );
  INV_X1 U22 ( .A(n1027), .ZN(n832) );
  INV_X1 U23 ( .A(n982), .ZN(n827) );
  INV_X1 U24 ( .A(n972), .ZN(n826) );
  INV_X1 U25 ( .A(n963), .ZN(n825) );
  INV_X1 U26 ( .A(n954), .ZN(n824) );
  INV_X1 U27 ( .A(n1091), .ZN(n839) );
  INV_X1 U28 ( .A(n1082), .ZN(n838) );
  INV_X1 U29 ( .A(n1073), .ZN(n837) );
  INV_X1 U30 ( .A(n1064), .ZN(n836) );
  INV_X1 U31 ( .A(n945), .ZN(n823) );
  INV_X1 U32 ( .A(n936), .ZN(n822) );
  INV_X1 U33 ( .A(n927), .ZN(n821) );
  INV_X1 U34 ( .A(n918), .ZN(n820) );
  INV_X1 U35 ( .A(n1018), .ZN(n831) );
  INV_X1 U36 ( .A(n1009), .ZN(n830) );
  INV_X1 U37 ( .A(n1000), .ZN(n829) );
  INV_X1 U38 ( .A(n991), .ZN(n828) );
  BUF_X1 U39 ( .A(N12), .Z(n606) );
  BUF_X1 U40 ( .A(N12), .Z(n607) );
  INV_X1 U41 ( .A(N13), .ZN(n845) );
  AND3_X1 U42 ( .A1(n618), .A2(n619), .A3(N12), .ZN(n1161) );
  AND3_X1 U43 ( .A1(N10), .A2(n619), .A3(N12), .ZN(n1151) );
  AND3_X1 U44 ( .A1(N11), .A2(n618), .A3(N12), .ZN(n1141) );
  AND3_X1 U45 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1131) );
  INV_X1 U46 ( .A(N14), .ZN(n846) );
  NAND2_X1 U47 ( .A1(n1191), .A2(n1201), .ZN(n1200) );
  NAND2_X1 U48 ( .A1(n1181), .A2(n1201), .ZN(n1190) );
  NAND2_X1 U49 ( .A1(n1171), .A2(n1201), .ZN(n1180) );
  NAND2_X1 U50 ( .A1(n1161), .A2(n1201), .ZN(n1170) );
  NAND2_X1 U51 ( .A1(n1151), .A2(n1201), .ZN(n1160) );
  NAND2_X1 U52 ( .A1(n1141), .A2(n1201), .ZN(n1150) );
  NAND2_X1 U53 ( .A1(n1131), .A2(n1201), .ZN(n1140) );
  NAND2_X1 U54 ( .A1(n1202), .A2(n1201), .ZN(n1211) );
  NAND2_X1 U55 ( .A1(n1120), .A2(n1202), .ZN(n1128) );
  NAND2_X1 U56 ( .A1(n1120), .A2(n1191), .ZN(n1118) );
  NAND2_X1 U57 ( .A1(n1120), .A2(n1181), .ZN(n1109) );
  NAND2_X1 U58 ( .A1(n1120), .A2(n1171), .ZN(n1100) );
  NAND2_X1 U59 ( .A1(n1047), .A2(n1202), .ZN(n1055) );
  NAND2_X1 U60 ( .A1(n1047), .A2(n1191), .ZN(n1045) );
  NAND2_X1 U61 ( .A1(n1047), .A2(n1181), .ZN(n1036) );
  NAND2_X1 U62 ( .A1(n1047), .A2(n1171), .ZN(n1027) );
  NAND2_X1 U63 ( .A1(n974), .A2(n1202), .ZN(n982) );
  NAND2_X1 U64 ( .A1(n974), .A2(n1191), .ZN(n972) );
  NAND2_X1 U65 ( .A1(n974), .A2(n1181), .ZN(n963) );
  NAND2_X1 U66 ( .A1(n974), .A2(n1171), .ZN(n954) );
  NAND2_X1 U67 ( .A1(n1120), .A2(n1161), .ZN(n1091) );
  NAND2_X1 U68 ( .A1(n1120), .A2(n1151), .ZN(n1082) );
  NAND2_X1 U69 ( .A1(n1120), .A2(n1141), .ZN(n1073) );
  NAND2_X1 U70 ( .A1(n1120), .A2(n1131), .ZN(n1064) );
  NAND2_X1 U71 ( .A1(n1047), .A2(n1161), .ZN(n1018) );
  NAND2_X1 U72 ( .A1(n1047), .A2(n1151), .ZN(n1009) );
  NAND2_X1 U73 ( .A1(n1047), .A2(n1141), .ZN(n1000) );
  NAND2_X1 U74 ( .A1(n1047), .A2(n1131), .ZN(n991) );
  NAND2_X1 U75 ( .A1(n974), .A2(n1161), .ZN(n945) );
  NAND2_X1 U76 ( .A1(n974), .A2(n1151), .ZN(n936) );
  NAND2_X1 U77 ( .A1(n974), .A2(n1141), .ZN(n927) );
  NAND2_X1 U78 ( .A1(n974), .A2(n1131), .ZN(n918) );
  AND3_X1 U79 ( .A1(n845), .A2(n846), .A3(n1130), .ZN(n1201) );
  AND3_X1 U80 ( .A1(N13), .A2(n1130), .A3(N14), .ZN(n974) );
  AND3_X1 U81 ( .A1(n1130), .A2(n846), .A3(N13), .ZN(n1120) );
  AND3_X1 U82 ( .A1(n1130), .A2(n845), .A3(N14), .ZN(n1047) );
  NOR2_X1 U83 ( .A1(n844), .A2(addr[5]), .ZN(n1130) );
  INV_X1 U84 ( .A(wr_en), .ZN(n844) );
  OAI21_X1 U85 ( .B1(n620), .B2(n1170), .A(n1169), .ZN(n878) );
  NAND2_X1 U86 ( .A1(\mem[4][0] ), .A2(n1170), .ZN(n1169) );
  OAI21_X1 U87 ( .B1(n621), .B2(n1170), .A(n1168), .ZN(n877) );
  NAND2_X1 U88 ( .A1(\mem[4][1] ), .A2(n1170), .ZN(n1168) );
  OAI21_X1 U89 ( .B1(n622), .B2(n1170), .A(n1167), .ZN(n876) );
  NAND2_X1 U90 ( .A1(\mem[4][2] ), .A2(n1170), .ZN(n1167) );
  OAI21_X1 U91 ( .B1(n623), .B2(n1170), .A(n1166), .ZN(n875) );
  NAND2_X1 U92 ( .A1(\mem[4][3] ), .A2(n1170), .ZN(n1166) );
  OAI21_X1 U93 ( .B1(n624), .B2(n1170), .A(n1165), .ZN(n874) );
  NAND2_X1 U94 ( .A1(\mem[4][4] ), .A2(n1170), .ZN(n1165) );
  OAI21_X1 U95 ( .B1(n625), .B2(n1170), .A(n1164), .ZN(n873) );
  NAND2_X1 U96 ( .A1(\mem[4][5] ), .A2(n1170), .ZN(n1164) );
  OAI21_X1 U97 ( .B1(n626), .B2(n1170), .A(n1163), .ZN(n872) );
  NAND2_X1 U98 ( .A1(\mem[4][6] ), .A2(n1170), .ZN(n1163) );
  OAI21_X1 U99 ( .B1(n627), .B2(n1170), .A(n1162), .ZN(n871) );
  NAND2_X1 U100 ( .A1(\mem[4][7] ), .A2(n1170), .ZN(n1162) );
  OAI21_X1 U101 ( .B1(n620), .B2(n1150), .A(n1149), .ZN(n862) );
  NAND2_X1 U102 ( .A1(\mem[6][0] ), .A2(n1150), .ZN(n1149) );
  OAI21_X1 U103 ( .B1(n621), .B2(n1150), .A(n1148), .ZN(n861) );
  NAND2_X1 U104 ( .A1(\mem[6][1] ), .A2(n1150), .ZN(n1148) );
  OAI21_X1 U105 ( .B1(n622), .B2(n1150), .A(n1147), .ZN(n860) );
  NAND2_X1 U106 ( .A1(\mem[6][2] ), .A2(n1150), .ZN(n1147) );
  OAI21_X1 U107 ( .B1(n623), .B2(n1150), .A(n1146), .ZN(n859) );
  NAND2_X1 U108 ( .A1(\mem[6][3] ), .A2(n1150), .ZN(n1146) );
  OAI21_X1 U109 ( .B1(n624), .B2(n1150), .A(n1145), .ZN(n858) );
  NAND2_X1 U110 ( .A1(\mem[6][4] ), .A2(n1150), .ZN(n1145) );
  OAI21_X1 U111 ( .B1(n625), .B2(n1150), .A(n1144), .ZN(n857) );
  NAND2_X1 U112 ( .A1(\mem[6][5] ), .A2(n1150), .ZN(n1144) );
  OAI21_X1 U113 ( .B1(n626), .B2(n1150), .A(n1143), .ZN(n856) );
  NAND2_X1 U114 ( .A1(\mem[6][6] ), .A2(n1150), .ZN(n1143) );
  OAI21_X1 U115 ( .B1(n627), .B2(n1150), .A(n1142), .ZN(n855) );
  NAND2_X1 U116 ( .A1(\mem[6][7] ), .A2(n1150), .ZN(n1142) );
  OAI21_X1 U117 ( .B1(n620), .B2(n1140), .A(n1139), .ZN(n854) );
  NAND2_X1 U118 ( .A1(\mem[7][0] ), .A2(n1140), .ZN(n1139) );
  OAI21_X1 U119 ( .B1(n621), .B2(n1140), .A(n1138), .ZN(n853) );
  NAND2_X1 U120 ( .A1(\mem[7][1] ), .A2(n1140), .ZN(n1138) );
  OAI21_X1 U121 ( .B1(n622), .B2(n1140), .A(n1137), .ZN(n852) );
  NAND2_X1 U122 ( .A1(\mem[7][2] ), .A2(n1140), .ZN(n1137) );
  OAI21_X1 U123 ( .B1(n623), .B2(n1140), .A(n1136), .ZN(n851) );
  NAND2_X1 U124 ( .A1(\mem[7][3] ), .A2(n1140), .ZN(n1136) );
  OAI21_X1 U125 ( .B1(n624), .B2(n1140), .A(n1135), .ZN(n850) );
  NAND2_X1 U126 ( .A1(\mem[7][4] ), .A2(n1140), .ZN(n1135) );
  OAI21_X1 U127 ( .B1(n625), .B2(n1140), .A(n1134), .ZN(n849) );
  NAND2_X1 U128 ( .A1(\mem[7][5] ), .A2(n1140), .ZN(n1134) );
  OAI21_X1 U129 ( .B1(n626), .B2(n1140), .A(n1133), .ZN(n848) );
  NAND2_X1 U130 ( .A1(\mem[7][6] ), .A2(n1140), .ZN(n1133) );
  OAI21_X1 U131 ( .B1(n627), .B2(n1140), .A(n1132), .ZN(n847) );
  NAND2_X1 U132 ( .A1(\mem[7][7] ), .A2(n1140), .ZN(n1132) );
  OAI21_X1 U133 ( .B1(n620), .B2(n1200), .A(n1199), .ZN(n902) );
  NAND2_X1 U134 ( .A1(\mem[1][0] ), .A2(n1200), .ZN(n1199) );
  OAI21_X1 U135 ( .B1(n621), .B2(n1200), .A(n1198), .ZN(n901) );
  NAND2_X1 U136 ( .A1(\mem[1][1] ), .A2(n1200), .ZN(n1198) );
  OAI21_X1 U137 ( .B1(n622), .B2(n1200), .A(n1197), .ZN(n900) );
  NAND2_X1 U138 ( .A1(\mem[1][2] ), .A2(n1200), .ZN(n1197) );
  OAI21_X1 U139 ( .B1(n623), .B2(n1200), .A(n1196), .ZN(n899) );
  NAND2_X1 U140 ( .A1(\mem[1][3] ), .A2(n1200), .ZN(n1196) );
  OAI21_X1 U141 ( .B1(n624), .B2(n1200), .A(n1195), .ZN(n898) );
  NAND2_X1 U142 ( .A1(\mem[1][4] ), .A2(n1200), .ZN(n1195) );
  OAI21_X1 U143 ( .B1(n625), .B2(n1200), .A(n1194), .ZN(n897) );
  NAND2_X1 U144 ( .A1(\mem[1][5] ), .A2(n1200), .ZN(n1194) );
  OAI21_X1 U145 ( .B1(n626), .B2(n1200), .A(n1193), .ZN(n896) );
  NAND2_X1 U146 ( .A1(\mem[1][6] ), .A2(n1200), .ZN(n1193) );
  OAI21_X1 U147 ( .B1(n627), .B2(n1200), .A(n1192), .ZN(n895) );
  NAND2_X1 U148 ( .A1(\mem[1][7] ), .A2(n1200), .ZN(n1192) );
  OAI21_X1 U149 ( .B1(n620), .B2(n1190), .A(n1189), .ZN(n894) );
  NAND2_X1 U150 ( .A1(\mem[2][0] ), .A2(n1190), .ZN(n1189) );
  OAI21_X1 U151 ( .B1(n621), .B2(n1190), .A(n1188), .ZN(n893) );
  NAND2_X1 U152 ( .A1(\mem[2][1] ), .A2(n1190), .ZN(n1188) );
  OAI21_X1 U153 ( .B1(n622), .B2(n1190), .A(n1187), .ZN(n892) );
  NAND2_X1 U154 ( .A1(\mem[2][2] ), .A2(n1190), .ZN(n1187) );
  OAI21_X1 U155 ( .B1(n623), .B2(n1190), .A(n1186), .ZN(n891) );
  NAND2_X1 U156 ( .A1(\mem[2][3] ), .A2(n1190), .ZN(n1186) );
  OAI21_X1 U157 ( .B1(n624), .B2(n1190), .A(n1185), .ZN(n890) );
  NAND2_X1 U158 ( .A1(\mem[2][4] ), .A2(n1190), .ZN(n1185) );
  OAI21_X1 U159 ( .B1(n625), .B2(n1190), .A(n1184), .ZN(n889) );
  NAND2_X1 U160 ( .A1(\mem[2][5] ), .A2(n1190), .ZN(n1184) );
  OAI21_X1 U161 ( .B1(n626), .B2(n1190), .A(n1183), .ZN(n888) );
  NAND2_X1 U162 ( .A1(\mem[2][6] ), .A2(n1190), .ZN(n1183) );
  OAI21_X1 U163 ( .B1(n627), .B2(n1190), .A(n1182), .ZN(n887) );
  NAND2_X1 U164 ( .A1(\mem[2][7] ), .A2(n1190), .ZN(n1182) );
  OAI21_X1 U165 ( .B1(n620), .B2(n1180), .A(n1179), .ZN(n886) );
  NAND2_X1 U166 ( .A1(\mem[3][0] ), .A2(n1180), .ZN(n1179) );
  OAI21_X1 U167 ( .B1(n621), .B2(n1180), .A(n1178), .ZN(n885) );
  NAND2_X1 U168 ( .A1(\mem[3][1] ), .A2(n1180), .ZN(n1178) );
  OAI21_X1 U169 ( .B1(n622), .B2(n1180), .A(n1177), .ZN(n884) );
  NAND2_X1 U170 ( .A1(\mem[3][2] ), .A2(n1180), .ZN(n1177) );
  OAI21_X1 U171 ( .B1(n623), .B2(n1180), .A(n1176), .ZN(n883) );
  NAND2_X1 U172 ( .A1(\mem[3][3] ), .A2(n1180), .ZN(n1176) );
  OAI21_X1 U173 ( .B1(n624), .B2(n1180), .A(n1175), .ZN(n882) );
  NAND2_X1 U174 ( .A1(\mem[3][4] ), .A2(n1180), .ZN(n1175) );
  OAI21_X1 U175 ( .B1(n625), .B2(n1180), .A(n1174), .ZN(n881) );
  NAND2_X1 U176 ( .A1(\mem[3][5] ), .A2(n1180), .ZN(n1174) );
  OAI21_X1 U177 ( .B1(n626), .B2(n1180), .A(n1173), .ZN(n880) );
  NAND2_X1 U178 ( .A1(\mem[3][6] ), .A2(n1180), .ZN(n1173) );
  OAI21_X1 U179 ( .B1(n627), .B2(n1180), .A(n1172), .ZN(n879) );
  NAND2_X1 U180 ( .A1(\mem[3][7] ), .A2(n1180), .ZN(n1172) );
  OAI21_X1 U181 ( .B1(n620), .B2(n1160), .A(n1159), .ZN(n870) );
  NAND2_X1 U182 ( .A1(\mem[5][0] ), .A2(n1160), .ZN(n1159) );
  OAI21_X1 U183 ( .B1(n621), .B2(n1160), .A(n1158), .ZN(n869) );
  NAND2_X1 U184 ( .A1(\mem[5][1] ), .A2(n1160), .ZN(n1158) );
  OAI21_X1 U185 ( .B1(n622), .B2(n1160), .A(n1157), .ZN(n868) );
  NAND2_X1 U186 ( .A1(\mem[5][2] ), .A2(n1160), .ZN(n1157) );
  OAI21_X1 U187 ( .B1(n623), .B2(n1160), .A(n1156), .ZN(n867) );
  NAND2_X1 U188 ( .A1(\mem[5][3] ), .A2(n1160), .ZN(n1156) );
  OAI21_X1 U189 ( .B1(n624), .B2(n1160), .A(n1155), .ZN(n866) );
  NAND2_X1 U190 ( .A1(\mem[5][4] ), .A2(n1160), .ZN(n1155) );
  OAI21_X1 U191 ( .B1(n625), .B2(n1160), .A(n1154), .ZN(n865) );
  NAND2_X1 U192 ( .A1(\mem[5][5] ), .A2(n1160), .ZN(n1154) );
  OAI21_X1 U193 ( .B1(n626), .B2(n1160), .A(n1153), .ZN(n864) );
  NAND2_X1 U194 ( .A1(\mem[5][6] ), .A2(n1160), .ZN(n1153) );
  OAI21_X1 U195 ( .B1(n627), .B2(n1160), .A(n1152), .ZN(n863) );
  NAND2_X1 U196 ( .A1(\mem[5][7] ), .A2(n1160), .ZN(n1152) );
  OAI21_X1 U197 ( .B1(n1211), .B2(n620), .A(n1210), .ZN(n910) );
  NAND2_X1 U198 ( .A1(\mem[0][0] ), .A2(n1211), .ZN(n1210) );
  OAI21_X1 U199 ( .B1(n1211), .B2(n621), .A(n1209), .ZN(n909) );
  NAND2_X1 U200 ( .A1(\mem[0][1] ), .A2(n1211), .ZN(n1209) );
  OAI21_X1 U201 ( .B1(n1211), .B2(n622), .A(n1208), .ZN(n908) );
  NAND2_X1 U202 ( .A1(\mem[0][2] ), .A2(n1211), .ZN(n1208) );
  OAI21_X1 U203 ( .B1(n1211), .B2(n623), .A(n1207), .ZN(n907) );
  NAND2_X1 U204 ( .A1(\mem[0][3] ), .A2(n1211), .ZN(n1207) );
  OAI21_X1 U205 ( .B1(n1211), .B2(n624), .A(n1206), .ZN(n906) );
  NAND2_X1 U206 ( .A1(\mem[0][4] ), .A2(n1211), .ZN(n1206) );
  OAI21_X1 U207 ( .B1(n1211), .B2(n625), .A(n1205), .ZN(n905) );
  NAND2_X1 U208 ( .A1(\mem[0][5] ), .A2(n1211), .ZN(n1205) );
  OAI21_X1 U209 ( .B1(n1211), .B2(n626), .A(n1204), .ZN(n904) );
  NAND2_X1 U210 ( .A1(\mem[0][6] ), .A2(n1211), .ZN(n1204) );
  OAI21_X1 U211 ( .B1(n1211), .B2(n627), .A(n1203), .ZN(n903) );
  NAND2_X1 U212 ( .A1(\mem[0][7] ), .A2(n1211), .ZN(n1203) );
  INV_X1 U213 ( .A(n1129), .ZN(n819) );
  AOI22_X1 U214 ( .A1(data_in[0]), .A2(n843), .B1(n1128), .B2(\mem[8][0] ), 
        .ZN(n1129) );
  INV_X1 U215 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U216 ( .A1(data_in[1]), .A2(n843), .B1(n1128), .B2(\mem[8][1] ), 
        .ZN(n1127) );
  INV_X1 U217 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U218 ( .A1(data_in[2]), .A2(n843), .B1(n1128), .B2(\mem[8][2] ), 
        .ZN(n1126) );
  INV_X1 U219 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U220 ( .A1(data_in[3]), .A2(n843), .B1(n1128), .B2(\mem[8][3] ), 
        .ZN(n1125) );
  INV_X1 U221 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U222 ( .A1(data_in[4]), .A2(n843), .B1(n1128), .B2(\mem[8][4] ), 
        .ZN(n1124) );
  INV_X1 U223 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U224 ( .A1(data_in[5]), .A2(n843), .B1(n1128), .B2(\mem[8][5] ), 
        .ZN(n1123) );
  INV_X1 U225 ( .A(n1122), .ZN(n813) );
  AOI22_X1 U226 ( .A1(data_in[6]), .A2(n843), .B1(n1128), .B2(\mem[8][6] ), 
        .ZN(n1122) );
  INV_X1 U227 ( .A(n1121), .ZN(n812) );
  AOI22_X1 U228 ( .A1(data_in[7]), .A2(n843), .B1(n1128), .B2(\mem[8][7] ), 
        .ZN(n1121) );
  INV_X1 U229 ( .A(n1119), .ZN(n811) );
  AOI22_X1 U230 ( .A1(data_in[0]), .A2(n842), .B1(n1118), .B2(\mem[9][0] ), 
        .ZN(n1119) );
  INV_X1 U231 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U232 ( .A1(data_in[1]), .A2(n842), .B1(n1118), .B2(\mem[9][1] ), 
        .ZN(n1117) );
  INV_X1 U233 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U234 ( .A1(data_in[2]), .A2(n842), .B1(n1118), .B2(\mem[9][2] ), 
        .ZN(n1116) );
  INV_X1 U235 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U236 ( .A1(data_in[3]), .A2(n842), .B1(n1118), .B2(\mem[9][3] ), 
        .ZN(n1115) );
  INV_X1 U237 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U238 ( .A1(data_in[4]), .A2(n842), .B1(n1118), .B2(\mem[9][4] ), 
        .ZN(n1114) );
  INV_X1 U239 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U240 ( .A1(data_in[5]), .A2(n842), .B1(n1118), .B2(\mem[9][5] ), 
        .ZN(n1113) );
  INV_X1 U241 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U242 ( .A1(data_in[6]), .A2(n842), .B1(n1118), .B2(\mem[9][6] ), 
        .ZN(n1112) );
  INV_X1 U243 ( .A(n1111), .ZN(n804) );
  AOI22_X1 U244 ( .A1(data_in[7]), .A2(n842), .B1(n1118), .B2(\mem[9][7] ), 
        .ZN(n1111) );
  INV_X1 U245 ( .A(n1110), .ZN(n803) );
  AOI22_X1 U246 ( .A1(data_in[0]), .A2(n841), .B1(n1109), .B2(\mem[10][0] ), 
        .ZN(n1110) );
  INV_X1 U247 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U248 ( .A1(data_in[1]), .A2(n841), .B1(n1109), .B2(\mem[10][1] ), 
        .ZN(n1108) );
  INV_X1 U249 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U250 ( .A1(data_in[2]), .A2(n841), .B1(n1109), .B2(\mem[10][2] ), 
        .ZN(n1107) );
  INV_X1 U251 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U252 ( .A1(data_in[3]), .A2(n841), .B1(n1109), .B2(\mem[10][3] ), 
        .ZN(n1106) );
  INV_X1 U253 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U254 ( .A1(data_in[4]), .A2(n841), .B1(n1109), .B2(\mem[10][4] ), 
        .ZN(n1105) );
  INV_X1 U255 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U256 ( .A1(data_in[5]), .A2(n841), .B1(n1109), .B2(\mem[10][5] ), 
        .ZN(n1104) );
  INV_X1 U257 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U258 ( .A1(data_in[6]), .A2(n841), .B1(n1109), .B2(\mem[10][6] ), 
        .ZN(n1103) );
  INV_X1 U259 ( .A(n1102), .ZN(n796) );
  AOI22_X1 U260 ( .A1(data_in[7]), .A2(n841), .B1(n1109), .B2(\mem[10][7] ), 
        .ZN(n1102) );
  INV_X1 U261 ( .A(n1101), .ZN(n795) );
  AOI22_X1 U262 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[11][0] ), 
        .ZN(n1101) );
  INV_X1 U263 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U264 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[11][1] ), 
        .ZN(n1099) );
  INV_X1 U265 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U266 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[11][2] ), 
        .ZN(n1098) );
  INV_X1 U267 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U268 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[11][3] ), 
        .ZN(n1097) );
  INV_X1 U269 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U270 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[11][4] ), 
        .ZN(n1096) );
  INV_X1 U271 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U272 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[11][5] ), 
        .ZN(n1095) );
  INV_X1 U273 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U274 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[11][6] ), 
        .ZN(n1094) );
  INV_X1 U275 ( .A(n1093), .ZN(n788) );
  AOI22_X1 U276 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[11][7] ), 
        .ZN(n1093) );
  INV_X1 U277 ( .A(n1092), .ZN(n787) );
  AOI22_X1 U278 ( .A1(data_in[0]), .A2(n839), .B1(n1091), .B2(\mem[12][0] ), 
        .ZN(n1092) );
  INV_X1 U279 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U280 ( .A1(data_in[1]), .A2(n839), .B1(n1091), .B2(\mem[12][1] ), 
        .ZN(n1090) );
  INV_X1 U281 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U282 ( .A1(data_in[2]), .A2(n839), .B1(n1091), .B2(\mem[12][2] ), 
        .ZN(n1089) );
  INV_X1 U283 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U284 ( .A1(data_in[3]), .A2(n839), .B1(n1091), .B2(\mem[12][3] ), 
        .ZN(n1088) );
  INV_X1 U285 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U286 ( .A1(data_in[4]), .A2(n839), .B1(n1091), .B2(\mem[12][4] ), 
        .ZN(n1087) );
  INV_X1 U287 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U288 ( .A1(data_in[5]), .A2(n839), .B1(n1091), .B2(\mem[12][5] ), 
        .ZN(n1086) );
  INV_X1 U289 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U290 ( .A1(data_in[6]), .A2(n839), .B1(n1091), .B2(\mem[12][6] ), 
        .ZN(n1085) );
  INV_X1 U291 ( .A(n1084), .ZN(n780) );
  AOI22_X1 U292 ( .A1(data_in[7]), .A2(n839), .B1(n1091), .B2(\mem[12][7] ), 
        .ZN(n1084) );
  INV_X1 U293 ( .A(n1083), .ZN(n779) );
  AOI22_X1 U294 ( .A1(data_in[0]), .A2(n838), .B1(n1082), .B2(\mem[13][0] ), 
        .ZN(n1083) );
  INV_X1 U295 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U296 ( .A1(data_in[1]), .A2(n838), .B1(n1082), .B2(\mem[13][1] ), 
        .ZN(n1081) );
  INV_X1 U297 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U298 ( .A1(data_in[2]), .A2(n838), .B1(n1082), .B2(\mem[13][2] ), 
        .ZN(n1080) );
  INV_X1 U299 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U300 ( .A1(data_in[3]), .A2(n838), .B1(n1082), .B2(\mem[13][3] ), 
        .ZN(n1079) );
  INV_X1 U301 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U302 ( .A1(data_in[4]), .A2(n838), .B1(n1082), .B2(\mem[13][4] ), 
        .ZN(n1078) );
  INV_X1 U303 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U304 ( .A1(data_in[5]), .A2(n838), .B1(n1082), .B2(\mem[13][5] ), 
        .ZN(n1077) );
  INV_X1 U305 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U306 ( .A1(data_in[6]), .A2(n838), .B1(n1082), .B2(\mem[13][6] ), 
        .ZN(n1076) );
  INV_X1 U307 ( .A(n1075), .ZN(n772) );
  AOI22_X1 U308 ( .A1(data_in[7]), .A2(n838), .B1(n1082), .B2(\mem[13][7] ), 
        .ZN(n1075) );
  INV_X1 U309 ( .A(n1074), .ZN(n771) );
  AOI22_X1 U310 ( .A1(data_in[0]), .A2(n837), .B1(n1073), .B2(\mem[14][0] ), 
        .ZN(n1074) );
  INV_X1 U311 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U312 ( .A1(data_in[1]), .A2(n837), .B1(n1073), .B2(\mem[14][1] ), 
        .ZN(n1072) );
  INV_X1 U313 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U314 ( .A1(data_in[2]), .A2(n837), .B1(n1073), .B2(\mem[14][2] ), 
        .ZN(n1071) );
  INV_X1 U315 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U316 ( .A1(data_in[3]), .A2(n837), .B1(n1073), .B2(\mem[14][3] ), 
        .ZN(n1070) );
  INV_X1 U317 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U318 ( .A1(data_in[4]), .A2(n837), .B1(n1073), .B2(\mem[14][4] ), 
        .ZN(n1069) );
  INV_X1 U319 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U320 ( .A1(data_in[5]), .A2(n837), .B1(n1073), .B2(\mem[14][5] ), 
        .ZN(n1068) );
  INV_X1 U321 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U322 ( .A1(data_in[6]), .A2(n837), .B1(n1073), .B2(\mem[14][6] ), 
        .ZN(n1067) );
  INV_X1 U323 ( .A(n1066), .ZN(n764) );
  AOI22_X1 U324 ( .A1(data_in[7]), .A2(n837), .B1(n1073), .B2(\mem[14][7] ), 
        .ZN(n1066) );
  INV_X1 U325 ( .A(n1065), .ZN(n763) );
  AOI22_X1 U326 ( .A1(data_in[0]), .A2(n836), .B1(n1064), .B2(\mem[15][0] ), 
        .ZN(n1065) );
  INV_X1 U327 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U328 ( .A1(data_in[1]), .A2(n836), .B1(n1064), .B2(\mem[15][1] ), 
        .ZN(n1063) );
  INV_X1 U329 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U330 ( .A1(data_in[2]), .A2(n836), .B1(n1064), .B2(\mem[15][2] ), 
        .ZN(n1062) );
  INV_X1 U331 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U332 ( .A1(data_in[3]), .A2(n836), .B1(n1064), .B2(\mem[15][3] ), 
        .ZN(n1061) );
  INV_X1 U333 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U334 ( .A1(data_in[4]), .A2(n836), .B1(n1064), .B2(\mem[15][4] ), 
        .ZN(n1060) );
  INV_X1 U335 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U336 ( .A1(data_in[5]), .A2(n836), .B1(n1064), .B2(\mem[15][5] ), 
        .ZN(n1059) );
  INV_X1 U337 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U338 ( .A1(data_in[6]), .A2(n836), .B1(n1064), .B2(\mem[15][6] ), 
        .ZN(n1058) );
  INV_X1 U339 ( .A(n1057), .ZN(n756) );
  AOI22_X1 U340 ( .A1(data_in[7]), .A2(n836), .B1(n1064), .B2(\mem[15][7] ), 
        .ZN(n1057) );
  INV_X1 U341 ( .A(n1056), .ZN(n755) );
  AOI22_X1 U342 ( .A1(data_in[0]), .A2(n835), .B1(n1055), .B2(\mem[16][0] ), 
        .ZN(n1056) );
  INV_X1 U343 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U344 ( .A1(data_in[1]), .A2(n835), .B1(n1055), .B2(\mem[16][1] ), 
        .ZN(n1054) );
  INV_X1 U345 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U346 ( .A1(data_in[2]), .A2(n835), .B1(n1055), .B2(\mem[16][2] ), 
        .ZN(n1053) );
  INV_X1 U347 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U348 ( .A1(data_in[3]), .A2(n835), .B1(n1055), .B2(\mem[16][3] ), 
        .ZN(n1052) );
  INV_X1 U349 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U350 ( .A1(data_in[4]), .A2(n835), .B1(n1055), .B2(\mem[16][4] ), 
        .ZN(n1051) );
  INV_X1 U351 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U352 ( .A1(data_in[5]), .A2(n835), .B1(n1055), .B2(\mem[16][5] ), 
        .ZN(n1050) );
  INV_X1 U353 ( .A(n1049), .ZN(n749) );
  AOI22_X1 U354 ( .A1(data_in[6]), .A2(n835), .B1(n1055), .B2(\mem[16][6] ), 
        .ZN(n1049) );
  INV_X1 U355 ( .A(n1048), .ZN(n748) );
  AOI22_X1 U356 ( .A1(data_in[7]), .A2(n835), .B1(n1055), .B2(\mem[16][7] ), 
        .ZN(n1048) );
  INV_X1 U357 ( .A(n1046), .ZN(n747) );
  AOI22_X1 U358 ( .A1(data_in[0]), .A2(n834), .B1(n1045), .B2(\mem[17][0] ), 
        .ZN(n1046) );
  INV_X1 U359 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U360 ( .A1(data_in[1]), .A2(n834), .B1(n1045), .B2(\mem[17][1] ), 
        .ZN(n1044) );
  INV_X1 U361 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U362 ( .A1(data_in[2]), .A2(n834), .B1(n1045), .B2(\mem[17][2] ), 
        .ZN(n1043) );
  INV_X1 U363 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U364 ( .A1(data_in[3]), .A2(n834), .B1(n1045), .B2(\mem[17][3] ), 
        .ZN(n1042) );
  INV_X1 U365 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U366 ( .A1(data_in[4]), .A2(n834), .B1(n1045), .B2(\mem[17][4] ), 
        .ZN(n1041) );
  INV_X1 U367 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U368 ( .A1(data_in[5]), .A2(n834), .B1(n1045), .B2(\mem[17][5] ), 
        .ZN(n1040) );
  INV_X1 U369 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U370 ( .A1(data_in[6]), .A2(n834), .B1(n1045), .B2(\mem[17][6] ), 
        .ZN(n1039) );
  INV_X1 U371 ( .A(n1038), .ZN(n740) );
  AOI22_X1 U372 ( .A1(data_in[7]), .A2(n834), .B1(n1045), .B2(\mem[17][7] ), 
        .ZN(n1038) );
  INV_X1 U373 ( .A(n1037), .ZN(n739) );
  AOI22_X1 U374 ( .A1(data_in[0]), .A2(n833), .B1(n1036), .B2(\mem[18][0] ), 
        .ZN(n1037) );
  INV_X1 U375 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U376 ( .A1(data_in[1]), .A2(n833), .B1(n1036), .B2(\mem[18][1] ), 
        .ZN(n1035) );
  INV_X1 U377 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U378 ( .A1(data_in[2]), .A2(n833), .B1(n1036), .B2(\mem[18][2] ), 
        .ZN(n1034) );
  INV_X1 U379 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U380 ( .A1(data_in[3]), .A2(n833), .B1(n1036), .B2(\mem[18][3] ), 
        .ZN(n1033) );
  INV_X1 U381 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U382 ( .A1(data_in[4]), .A2(n833), .B1(n1036), .B2(\mem[18][4] ), 
        .ZN(n1032) );
  INV_X1 U383 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U384 ( .A1(data_in[5]), .A2(n833), .B1(n1036), .B2(\mem[18][5] ), 
        .ZN(n1031) );
  INV_X1 U385 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U386 ( .A1(data_in[6]), .A2(n833), .B1(n1036), .B2(\mem[18][6] ), 
        .ZN(n1030) );
  INV_X1 U387 ( .A(n1029), .ZN(n732) );
  AOI22_X1 U388 ( .A1(data_in[7]), .A2(n833), .B1(n1036), .B2(\mem[18][7] ), 
        .ZN(n1029) );
  INV_X1 U389 ( .A(n1028), .ZN(n731) );
  AOI22_X1 U390 ( .A1(data_in[0]), .A2(n832), .B1(n1027), .B2(\mem[19][0] ), 
        .ZN(n1028) );
  INV_X1 U391 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U392 ( .A1(data_in[1]), .A2(n832), .B1(n1027), .B2(\mem[19][1] ), 
        .ZN(n1026) );
  INV_X1 U393 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U394 ( .A1(data_in[2]), .A2(n832), .B1(n1027), .B2(\mem[19][2] ), 
        .ZN(n1025) );
  INV_X1 U395 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U396 ( .A1(data_in[3]), .A2(n832), .B1(n1027), .B2(\mem[19][3] ), 
        .ZN(n1024) );
  INV_X1 U397 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U398 ( .A1(data_in[4]), .A2(n832), .B1(n1027), .B2(\mem[19][4] ), 
        .ZN(n1023) );
  INV_X1 U399 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U400 ( .A1(data_in[5]), .A2(n832), .B1(n1027), .B2(\mem[19][5] ), 
        .ZN(n1022) );
  INV_X1 U401 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U402 ( .A1(data_in[6]), .A2(n832), .B1(n1027), .B2(\mem[19][6] ), 
        .ZN(n1021) );
  INV_X1 U403 ( .A(n1020), .ZN(n724) );
  AOI22_X1 U404 ( .A1(data_in[7]), .A2(n832), .B1(n1027), .B2(\mem[19][7] ), 
        .ZN(n1020) );
  INV_X1 U405 ( .A(n1019), .ZN(n723) );
  AOI22_X1 U406 ( .A1(data_in[0]), .A2(n831), .B1(n1018), .B2(\mem[20][0] ), 
        .ZN(n1019) );
  INV_X1 U407 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U408 ( .A1(data_in[1]), .A2(n831), .B1(n1018), .B2(\mem[20][1] ), 
        .ZN(n1017) );
  INV_X1 U409 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U410 ( .A1(data_in[2]), .A2(n831), .B1(n1018), .B2(\mem[20][2] ), 
        .ZN(n1016) );
  INV_X1 U411 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U412 ( .A1(data_in[3]), .A2(n831), .B1(n1018), .B2(\mem[20][3] ), 
        .ZN(n1015) );
  INV_X1 U413 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U414 ( .A1(data_in[4]), .A2(n831), .B1(n1018), .B2(\mem[20][4] ), 
        .ZN(n1014) );
  INV_X1 U415 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U416 ( .A1(data_in[5]), .A2(n831), .B1(n1018), .B2(\mem[20][5] ), 
        .ZN(n1013) );
  INV_X1 U417 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U418 ( .A1(data_in[6]), .A2(n831), .B1(n1018), .B2(\mem[20][6] ), 
        .ZN(n1012) );
  INV_X1 U419 ( .A(n1011), .ZN(n716) );
  AOI22_X1 U420 ( .A1(data_in[7]), .A2(n831), .B1(n1018), .B2(\mem[20][7] ), 
        .ZN(n1011) );
  INV_X1 U421 ( .A(n1010), .ZN(n715) );
  AOI22_X1 U422 ( .A1(data_in[0]), .A2(n830), .B1(n1009), .B2(\mem[21][0] ), 
        .ZN(n1010) );
  INV_X1 U423 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U424 ( .A1(data_in[1]), .A2(n830), .B1(n1009), .B2(\mem[21][1] ), 
        .ZN(n1008) );
  INV_X1 U425 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U426 ( .A1(data_in[2]), .A2(n830), .B1(n1009), .B2(\mem[21][2] ), 
        .ZN(n1007) );
  INV_X1 U427 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U428 ( .A1(data_in[3]), .A2(n830), .B1(n1009), .B2(\mem[21][3] ), 
        .ZN(n1006) );
  INV_X1 U429 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U430 ( .A1(data_in[4]), .A2(n830), .B1(n1009), .B2(\mem[21][4] ), 
        .ZN(n1005) );
  INV_X1 U431 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U432 ( .A1(data_in[5]), .A2(n830), .B1(n1009), .B2(\mem[21][5] ), 
        .ZN(n1004) );
  INV_X1 U433 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U434 ( .A1(data_in[6]), .A2(n830), .B1(n1009), .B2(\mem[21][6] ), 
        .ZN(n1003) );
  INV_X1 U435 ( .A(n1002), .ZN(n708) );
  AOI22_X1 U436 ( .A1(data_in[7]), .A2(n830), .B1(n1009), .B2(\mem[21][7] ), 
        .ZN(n1002) );
  INV_X1 U437 ( .A(n1001), .ZN(n707) );
  AOI22_X1 U438 ( .A1(data_in[0]), .A2(n829), .B1(n1000), .B2(\mem[22][0] ), 
        .ZN(n1001) );
  INV_X1 U439 ( .A(n999), .ZN(n706) );
  AOI22_X1 U440 ( .A1(data_in[1]), .A2(n829), .B1(n1000), .B2(\mem[22][1] ), 
        .ZN(n999) );
  INV_X1 U441 ( .A(n998), .ZN(n705) );
  AOI22_X1 U442 ( .A1(data_in[2]), .A2(n829), .B1(n1000), .B2(\mem[22][2] ), 
        .ZN(n998) );
  INV_X1 U443 ( .A(n997), .ZN(n704) );
  AOI22_X1 U444 ( .A1(data_in[3]), .A2(n829), .B1(n1000), .B2(\mem[22][3] ), 
        .ZN(n997) );
  INV_X1 U445 ( .A(n996), .ZN(n703) );
  AOI22_X1 U446 ( .A1(data_in[4]), .A2(n829), .B1(n1000), .B2(\mem[22][4] ), 
        .ZN(n996) );
  INV_X1 U447 ( .A(n995), .ZN(n702) );
  AOI22_X1 U448 ( .A1(data_in[5]), .A2(n829), .B1(n1000), .B2(\mem[22][5] ), 
        .ZN(n995) );
  INV_X1 U449 ( .A(n994), .ZN(n701) );
  AOI22_X1 U450 ( .A1(data_in[6]), .A2(n829), .B1(n1000), .B2(\mem[22][6] ), 
        .ZN(n994) );
  INV_X1 U451 ( .A(n993), .ZN(n700) );
  AOI22_X1 U452 ( .A1(data_in[7]), .A2(n829), .B1(n1000), .B2(\mem[22][7] ), 
        .ZN(n993) );
  INV_X1 U453 ( .A(n992), .ZN(n699) );
  AOI22_X1 U454 ( .A1(data_in[0]), .A2(n828), .B1(n991), .B2(\mem[23][0] ), 
        .ZN(n992) );
  INV_X1 U455 ( .A(n990), .ZN(n698) );
  AOI22_X1 U456 ( .A1(data_in[1]), .A2(n828), .B1(n991), .B2(\mem[23][1] ), 
        .ZN(n990) );
  INV_X1 U457 ( .A(n989), .ZN(n697) );
  AOI22_X1 U458 ( .A1(data_in[2]), .A2(n828), .B1(n991), .B2(\mem[23][2] ), 
        .ZN(n989) );
  INV_X1 U459 ( .A(n988), .ZN(n696) );
  AOI22_X1 U460 ( .A1(data_in[3]), .A2(n828), .B1(n991), .B2(\mem[23][3] ), 
        .ZN(n988) );
  INV_X1 U461 ( .A(n987), .ZN(n695) );
  AOI22_X1 U462 ( .A1(data_in[4]), .A2(n828), .B1(n991), .B2(\mem[23][4] ), 
        .ZN(n987) );
  INV_X1 U463 ( .A(n986), .ZN(n694) );
  AOI22_X1 U464 ( .A1(data_in[5]), .A2(n828), .B1(n991), .B2(\mem[23][5] ), 
        .ZN(n986) );
  INV_X1 U465 ( .A(n985), .ZN(n693) );
  AOI22_X1 U466 ( .A1(data_in[6]), .A2(n828), .B1(n991), .B2(\mem[23][6] ), 
        .ZN(n985) );
  INV_X1 U467 ( .A(n984), .ZN(n692) );
  AOI22_X1 U468 ( .A1(data_in[7]), .A2(n828), .B1(n991), .B2(\mem[23][7] ), 
        .ZN(n984) );
  INV_X1 U469 ( .A(n983), .ZN(n691) );
  AOI22_X1 U470 ( .A1(data_in[0]), .A2(n827), .B1(n982), .B2(\mem[24][0] ), 
        .ZN(n983) );
  INV_X1 U471 ( .A(n981), .ZN(n690) );
  AOI22_X1 U472 ( .A1(data_in[1]), .A2(n827), .B1(n982), .B2(\mem[24][1] ), 
        .ZN(n981) );
  INV_X1 U473 ( .A(n980), .ZN(n689) );
  AOI22_X1 U474 ( .A1(data_in[2]), .A2(n827), .B1(n982), .B2(\mem[24][2] ), 
        .ZN(n980) );
  INV_X1 U475 ( .A(n979), .ZN(n688) );
  AOI22_X1 U476 ( .A1(data_in[3]), .A2(n827), .B1(n982), .B2(\mem[24][3] ), 
        .ZN(n979) );
  INV_X1 U477 ( .A(n978), .ZN(n687) );
  AOI22_X1 U478 ( .A1(data_in[4]), .A2(n827), .B1(n982), .B2(\mem[24][4] ), 
        .ZN(n978) );
  INV_X1 U479 ( .A(n977), .ZN(n686) );
  AOI22_X1 U480 ( .A1(data_in[5]), .A2(n827), .B1(n982), .B2(\mem[24][5] ), 
        .ZN(n977) );
  INV_X1 U481 ( .A(n976), .ZN(n685) );
  AOI22_X1 U482 ( .A1(data_in[6]), .A2(n827), .B1(n982), .B2(\mem[24][6] ), 
        .ZN(n976) );
  INV_X1 U483 ( .A(n975), .ZN(n684) );
  AOI22_X1 U484 ( .A1(data_in[7]), .A2(n827), .B1(n982), .B2(\mem[24][7] ), 
        .ZN(n975) );
  INV_X1 U485 ( .A(n973), .ZN(n683) );
  AOI22_X1 U486 ( .A1(data_in[0]), .A2(n826), .B1(n972), .B2(\mem[25][0] ), 
        .ZN(n973) );
  INV_X1 U487 ( .A(n971), .ZN(n682) );
  AOI22_X1 U488 ( .A1(data_in[1]), .A2(n826), .B1(n972), .B2(\mem[25][1] ), 
        .ZN(n971) );
  INV_X1 U489 ( .A(n970), .ZN(n681) );
  AOI22_X1 U490 ( .A1(data_in[2]), .A2(n826), .B1(n972), .B2(\mem[25][2] ), 
        .ZN(n970) );
  INV_X1 U491 ( .A(n969), .ZN(n680) );
  AOI22_X1 U492 ( .A1(data_in[3]), .A2(n826), .B1(n972), .B2(\mem[25][3] ), 
        .ZN(n969) );
  INV_X1 U493 ( .A(n968), .ZN(n679) );
  AOI22_X1 U494 ( .A1(data_in[4]), .A2(n826), .B1(n972), .B2(\mem[25][4] ), 
        .ZN(n968) );
  INV_X1 U495 ( .A(n967), .ZN(n678) );
  AOI22_X1 U496 ( .A1(data_in[5]), .A2(n826), .B1(n972), .B2(\mem[25][5] ), 
        .ZN(n967) );
  INV_X1 U497 ( .A(n966), .ZN(n677) );
  AOI22_X1 U498 ( .A1(data_in[6]), .A2(n826), .B1(n972), .B2(\mem[25][6] ), 
        .ZN(n966) );
  INV_X1 U499 ( .A(n965), .ZN(n676) );
  AOI22_X1 U500 ( .A1(data_in[7]), .A2(n826), .B1(n972), .B2(\mem[25][7] ), 
        .ZN(n965) );
  INV_X1 U501 ( .A(n964), .ZN(n675) );
  AOI22_X1 U502 ( .A1(data_in[0]), .A2(n825), .B1(n963), .B2(\mem[26][0] ), 
        .ZN(n964) );
  INV_X1 U503 ( .A(n962), .ZN(n674) );
  AOI22_X1 U504 ( .A1(data_in[1]), .A2(n825), .B1(n963), .B2(\mem[26][1] ), 
        .ZN(n962) );
  INV_X1 U505 ( .A(n961), .ZN(n673) );
  AOI22_X1 U506 ( .A1(data_in[2]), .A2(n825), .B1(n963), .B2(\mem[26][2] ), 
        .ZN(n961) );
  INV_X1 U507 ( .A(n960), .ZN(n672) );
  AOI22_X1 U508 ( .A1(data_in[3]), .A2(n825), .B1(n963), .B2(\mem[26][3] ), 
        .ZN(n960) );
  INV_X1 U509 ( .A(n959), .ZN(n671) );
  AOI22_X1 U510 ( .A1(data_in[4]), .A2(n825), .B1(n963), .B2(\mem[26][4] ), 
        .ZN(n959) );
  INV_X1 U511 ( .A(n958), .ZN(n670) );
  AOI22_X1 U512 ( .A1(data_in[5]), .A2(n825), .B1(n963), .B2(\mem[26][5] ), 
        .ZN(n958) );
  INV_X1 U513 ( .A(n957), .ZN(n669) );
  AOI22_X1 U514 ( .A1(data_in[6]), .A2(n825), .B1(n963), .B2(\mem[26][6] ), 
        .ZN(n957) );
  INV_X1 U515 ( .A(n956), .ZN(n668) );
  AOI22_X1 U516 ( .A1(data_in[7]), .A2(n825), .B1(n963), .B2(\mem[26][7] ), 
        .ZN(n956) );
  INV_X1 U517 ( .A(n955), .ZN(n667) );
  AOI22_X1 U518 ( .A1(data_in[0]), .A2(n824), .B1(n954), .B2(\mem[27][0] ), 
        .ZN(n955) );
  INV_X1 U519 ( .A(n953), .ZN(n666) );
  AOI22_X1 U520 ( .A1(data_in[1]), .A2(n824), .B1(n954), .B2(\mem[27][1] ), 
        .ZN(n953) );
  INV_X1 U521 ( .A(n952), .ZN(n665) );
  AOI22_X1 U522 ( .A1(data_in[2]), .A2(n824), .B1(n954), .B2(\mem[27][2] ), 
        .ZN(n952) );
  INV_X1 U523 ( .A(n951), .ZN(n664) );
  AOI22_X1 U524 ( .A1(data_in[3]), .A2(n824), .B1(n954), .B2(\mem[27][3] ), 
        .ZN(n951) );
  INV_X1 U525 ( .A(n950), .ZN(n663) );
  AOI22_X1 U526 ( .A1(data_in[4]), .A2(n824), .B1(n954), .B2(\mem[27][4] ), 
        .ZN(n950) );
  INV_X1 U527 ( .A(n949), .ZN(n662) );
  AOI22_X1 U528 ( .A1(data_in[5]), .A2(n824), .B1(n954), .B2(\mem[27][5] ), 
        .ZN(n949) );
  INV_X1 U529 ( .A(n948), .ZN(n661) );
  AOI22_X1 U530 ( .A1(data_in[6]), .A2(n824), .B1(n954), .B2(\mem[27][6] ), 
        .ZN(n948) );
  INV_X1 U531 ( .A(n947), .ZN(n660) );
  AOI22_X1 U532 ( .A1(data_in[7]), .A2(n824), .B1(n954), .B2(\mem[27][7] ), 
        .ZN(n947) );
  INV_X1 U533 ( .A(n946), .ZN(n659) );
  AOI22_X1 U534 ( .A1(data_in[0]), .A2(n823), .B1(n945), .B2(\mem[28][0] ), 
        .ZN(n946) );
  INV_X1 U535 ( .A(n944), .ZN(n658) );
  AOI22_X1 U536 ( .A1(data_in[1]), .A2(n823), .B1(n945), .B2(\mem[28][1] ), 
        .ZN(n944) );
  INV_X1 U537 ( .A(n943), .ZN(n657) );
  AOI22_X1 U538 ( .A1(data_in[2]), .A2(n823), .B1(n945), .B2(\mem[28][2] ), 
        .ZN(n943) );
  INV_X1 U539 ( .A(n942), .ZN(n656) );
  AOI22_X1 U540 ( .A1(data_in[3]), .A2(n823), .B1(n945), .B2(\mem[28][3] ), 
        .ZN(n942) );
  INV_X1 U541 ( .A(n941), .ZN(n655) );
  AOI22_X1 U542 ( .A1(data_in[4]), .A2(n823), .B1(n945), .B2(\mem[28][4] ), 
        .ZN(n941) );
  INV_X1 U543 ( .A(n940), .ZN(n654) );
  AOI22_X1 U544 ( .A1(data_in[5]), .A2(n823), .B1(n945), .B2(\mem[28][5] ), 
        .ZN(n940) );
  INV_X1 U545 ( .A(n939), .ZN(n653) );
  AOI22_X1 U546 ( .A1(data_in[6]), .A2(n823), .B1(n945), .B2(\mem[28][6] ), 
        .ZN(n939) );
  INV_X1 U547 ( .A(n938), .ZN(n652) );
  AOI22_X1 U548 ( .A1(data_in[7]), .A2(n823), .B1(n945), .B2(\mem[28][7] ), 
        .ZN(n938) );
  INV_X1 U549 ( .A(n937), .ZN(n651) );
  AOI22_X1 U550 ( .A1(data_in[0]), .A2(n822), .B1(n936), .B2(\mem[29][0] ), 
        .ZN(n937) );
  INV_X1 U551 ( .A(n935), .ZN(n650) );
  AOI22_X1 U552 ( .A1(data_in[1]), .A2(n822), .B1(n936), .B2(\mem[29][1] ), 
        .ZN(n935) );
  INV_X1 U553 ( .A(n934), .ZN(n649) );
  AOI22_X1 U554 ( .A1(data_in[2]), .A2(n822), .B1(n936), .B2(\mem[29][2] ), 
        .ZN(n934) );
  INV_X1 U555 ( .A(n933), .ZN(n648) );
  AOI22_X1 U556 ( .A1(data_in[3]), .A2(n822), .B1(n936), .B2(\mem[29][3] ), 
        .ZN(n933) );
  INV_X1 U557 ( .A(n932), .ZN(n647) );
  AOI22_X1 U558 ( .A1(data_in[4]), .A2(n822), .B1(n936), .B2(\mem[29][4] ), 
        .ZN(n932) );
  INV_X1 U559 ( .A(n931), .ZN(n646) );
  AOI22_X1 U560 ( .A1(data_in[5]), .A2(n822), .B1(n936), .B2(\mem[29][5] ), 
        .ZN(n931) );
  INV_X1 U561 ( .A(n930), .ZN(n645) );
  AOI22_X1 U562 ( .A1(data_in[6]), .A2(n822), .B1(n936), .B2(\mem[29][6] ), 
        .ZN(n930) );
  INV_X1 U563 ( .A(n929), .ZN(n644) );
  AOI22_X1 U564 ( .A1(data_in[7]), .A2(n822), .B1(n936), .B2(\mem[29][7] ), 
        .ZN(n929) );
  INV_X1 U565 ( .A(n928), .ZN(n643) );
  AOI22_X1 U566 ( .A1(data_in[0]), .A2(n821), .B1(n927), .B2(\mem[30][0] ), 
        .ZN(n928) );
  INV_X1 U567 ( .A(n926), .ZN(n642) );
  AOI22_X1 U568 ( .A1(data_in[1]), .A2(n821), .B1(n927), .B2(\mem[30][1] ), 
        .ZN(n926) );
  INV_X1 U569 ( .A(n925), .ZN(n641) );
  AOI22_X1 U570 ( .A1(data_in[2]), .A2(n821), .B1(n927), .B2(\mem[30][2] ), 
        .ZN(n925) );
  INV_X1 U571 ( .A(n924), .ZN(n640) );
  AOI22_X1 U572 ( .A1(data_in[3]), .A2(n821), .B1(n927), .B2(\mem[30][3] ), 
        .ZN(n924) );
  INV_X1 U573 ( .A(n923), .ZN(n639) );
  AOI22_X1 U574 ( .A1(data_in[4]), .A2(n821), .B1(n927), .B2(\mem[30][4] ), 
        .ZN(n923) );
  INV_X1 U575 ( .A(n922), .ZN(n638) );
  AOI22_X1 U576 ( .A1(data_in[5]), .A2(n821), .B1(n927), .B2(\mem[30][5] ), 
        .ZN(n922) );
  INV_X1 U577 ( .A(n921), .ZN(n637) );
  AOI22_X1 U578 ( .A1(data_in[6]), .A2(n821), .B1(n927), .B2(\mem[30][6] ), 
        .ZN(n921) );
  INV_X1 U579 ( .A(n920), .ZN(n636) );
  AOI22_X1 U580 ( .A1(data_in[7]), .A2(n821), .B1(n927), .B2(\mem[30][7] ), 
        .ZN(n920) );
  INV_X1 U581 ( .A(n919), .ZN(n635) );
  AOI22_X1 U582 ( .A1(data_in[0]), .A2(n820), .B1(n918), .B2(\mem[31][0] ), 
        .ZN(n919) );
  INV_X1 U583 ( .A(n917), .ZN(n634) );
  AOI22_X1 U584 ( .A1(data_in[1]), .A2(n820), .B1(n918), .B2(\mem[31][1] ), 
        .ZN(n917) );
  INV_X1 U585 ( .A(n916), .ZN(n633) );
  AOI22_X1 U586 ( .A1(data_in[2]), .A2(n820), .B1(n918), .B2(\mem[31][2] ), 
        .ZN(n916) );
  INV_X1 U587 ( .A(n915), .ZN(n632) );
  AOI22_X1 U588 ( .A1(data_in[3]), .A2(n820), .B1(n918), .B2(\mem[31][3] ), 
        .ZN(n915) );
  INV_X1 U589 ( .A(n914), .ZN(n631) );
  AOI22_X1 U590 ( .A1(data_in[4]), .A2(n820), .B1(n918), .B2(\mem[31][4] ), 
        .ZN(n914) );
  INV_X1 U591 ( .A(n913), .ZN(n630) );
  AOI22_X1 U592 ( .A1(data_in[5]), .A2(n820), .B1(n918), .B2(\mem[31][5] ), 
        .ZN(n913) );
  INV_X1 U593 ( .A(n912), .ZN(n629) );
  AOI22_X1 U594 ( .A1(data_in[6]), .A2(n820), .B1(n918), .B2(\mem[31][6] ), 
        .ZN(n912) );
  INV_X1 U595 ( .A(n911), .ZN(n628) );
  AOI22_X1 U596 ( .A1(data_in[7]), .A2(n820), .B1(n918), .B2(\mem[31][7] ), 
        .ZN(n911) );
  MUX2_X1 U597 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n611), .Z(n1) );
  MUX2_X1 U598 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n611), .Z(n2) );
  MUX2_X1 U599 ( .A(n2), .B(n1), .S(n608), .Z(n3) );
  MUX2_X1 U600 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n611), .Z(n4) );
  MUX2_X1 U601 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n611), .Z(n5) );
  MUX2_X1 U602 ( .A(n5), .B(n4), .S(n608), .Z(n6) );
  MUX2_X1 U603 ( .A(n6), .B(n3), .S(N12), .Z(n7) );
  MUX2_X1 U604 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n611), .Z(n8) );
  MUX2_X1 U605 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n611), .Z(n9) );
  MUX2_X1 U606 ( .A(n9), .B(n8), .S(n608), .Z(n10) );
  MUX2_X1 U607 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n611), .Z(n11) );
  MUX2_X1 U608 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n611), .Z(n12) );
  MUX2_X1 U609 ( .A(n12), .B(n11), .S(n608), .Z(n13) );
  MUX2_X1 U610 ( .A(n13), .B(n10), .S(n606), .Z(n14) );
  MUX2_X1 U611 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U612 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n617), .Z(n16) );
  MUX2_X1 U613 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n617), .Z(n17) );
  MUX2_X1 U614 ( .A(n17), .B(n16), .S(n609), .Z(n18) );
  MUX2_X1 U615 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n617), .Z(n19) );
  MUX2_X1 U616 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n614), .Z(n20) );
  MUX2_X1 U617 ( .A(n20), .B(n19), .S(n609), .Z(n21) );
  MUX2_X1 U618 ( .A(n21), .B(n18), .S(n607), .Z(n22) );
  MUX2_X1 U619 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n617), .Z(n23) );
  MUX2_X1 U620 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n616), .Z(n24) );
  MUX2_X1 U621 ( .A(n24), .B(n23), .S(n609), .Z(n25) );
  MUX2_X1 U622 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n617), .Z(n26) );
  MUX2_X1 U623 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n615), .Z(n27) );
  MUX2_X1 U624 ( .A(n27), .B(n26), .S(n609), .Z(n28) );
  MUX2_X1 U625 ( .A(n28), .B(n25), .S(n607), .Z(n29) );
  MUX2_X1 U626 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U627 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U628 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n615), .Z(n31) );
  MUX2_X1 U629 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n617), .Z(n32) );
  MUX2_X1 U630 ( .A(n32), .B(n31), .S(n609), .Z(n33) );
  MUX2_X1 U631 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n616), .Z(n34) );
  MUX2_X1 U632 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n617), .Z(n35) );
  MUX2_X1 U633 ( .A(n35), .B(n34), .S(n609), .Z(n36) );
  MUX2_X1 U634 ( .A(n36), .B(n33), .S(n607), .Z(n37) );
  MUX2_X1 U635 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n617), .Z(n38) );
  MUX2_X1 U636 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n617), .Z(n39) );
  MUX2_X1 U637 ( .A(n39), .B(n38), .S(n609), .Z(n40) );
  MUX2_X1 U638 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n617), .Z(n41) );
  MUX2_X1 U639 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n617), .Z(n42) );
  MUX2_X1 U640 ( .A(n42), .B(n41), .S(n609), .Z(n43) );
  MUX2_X1 U641 ( .A(n43), .B(n40), .S(N12), .Z(n44) );
  MUX2_X1 U642 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U643 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n614), .Z(n46) );
  MUX2_X1 U644 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(N10), .Z(n47) );
  MUX2_X1 U645 ( .A(n47), .B(n46), .S(n609), .Z(n48) );
  MUX2_X1 U646 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n617), .Z(n49) );
  MUX2_X1 U647 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n617), .Z(n50) );
  MUX2_X1 U648 ( .A(n50), .B(n49), .S(n609), .Z(n51) );
  MUX2_X1 U649 ( .A(n51), .B(n48), .S(n606), .Z(n52) );
  MUX2_X1 U650 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n617), .Z(n53) );
  MUX2_X1 U651 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n617), .Z(n54) );
  MUX2_X1 U652 ( .A(n54), .B(n53), .S(n609), .Z(n55) );
  MUX2_X1 U653 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n617), .Z(n56) );
  MUX2_X1 U654 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n617), .Z(n57) );
  MUX2_X1 U655 ( .A(n57), .B(n56), .S(n609), .Z(n58) );
  MUX2_X1 U656 ( .A(n58), .B(n55), .S(N12), .Z(n59) );
  MUX2_X1 U657 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U658 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U659 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n613), .Z(n61) );
  MUX2_X1 U660 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n613), .Z(n62) );
  MUX2_X1 U661 ( .A(n62), .B(n61), .S(n610), .Z(n63) );
  MUX2_X1 U662 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n612), .Z(n64) );
  MUX2_X1 U663 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n613), .Z(n65) );
  MUX2_X1 U664 ( .A(n65), .B(n64), .S(n610), .Z(n66) );
  MUX2_X1 U665 ( .A(n66), .B(n63), .S(n606), .Z(n67) );
  MUX2_X1 U666 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n612), .Z(n68) );
  MUX2_X1 U667 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n614), .Z(n69) );
  MUX2_X1 U668 ( .A(n69), .B(n68), .S(n610), .Z(n70) );
  MUX2_X1 U669 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n612), .Z(n71) );
  MUX2_X1 U670 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n615), .Z(n72) );
  MUX2_X1 U671 ( .A(n72), .B(n71), .S(n610), .Z(n73) );
  MUX2_X1 U672 ( .A(n73), .B(n70), .S(n606), .Z(n74) );
  MUX2_X1 U673 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U674 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n613), .Z(n76) );
  MUX2_X1 U675 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n612), .Z(n77) );
  MUX2_X1 U676 ( .A(n77), .B(n76), .S(n610), .Z(n78) );
  MUX2_X1 U677 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n613), .Z(n79) );
  MUX2_X1 U678 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n616), .Z(n80) );
  MUX2_X1 U679 ( .A(n80), .B(n79), .S(n610), .Z(n81) );
  MUX2_X1 U680 ( .A(n81), .B(n78), .S(n606), .Z(n82) );
  MUX2_X1 U681 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n613), .Z(n83) );
  MUX2_X1 U682 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n613), .Z(n84) );
  MUX2_X1 U683 ( .A(n84), .B(n83), .S(n610), .Z(n85) );
  MUX2_X1 U684 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n612), .Z(n86) );
  MUX2_X1 U685 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n612), .Z(n87) );
  MUX2_X1 U686 ( .A(n87), .B(n86), .S(n610), .Z(n88) );
  MUX2_X1 U687 ( .A(n88), .B(n85), .S(n606), .Z(n89) );
  MUX2_X1 U688 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U689 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U690 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n613), .Z(n91) );
  MUX2_X1 U691 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n612), .Z(n92) );
  MUX2_X1 U692 ( .A(n92), .B(n91), .S(n610), .Z(n93) );
  MUX2_X1 U693 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n612), .Z(n94) );
  MUX2_X1 U694 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n612), .Z(n95) );
  MUX2_X1 U695 ( .A(n95), .B(n94), .S(n610), .Z(n96) );
  MUX2_X1 U696 ( .A(n96), .B(n93), .S(n606), .Z(n97) );
  MUX2_X1 U697 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n613), .Z(n98) );
  MUX2_X1 U698 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n613), .Z(n99) );
  MUX2_X1 U699 ( .A(n99), .B(n98), .S(n610), .Z(n100) );
  MUX2_X1 U700 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n613), .Z(n101) );
  MUX2_X1 U701 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n612), .Z(n102) );
  MUX2_X1 U702 ( .A(n102), .B(n101), .S(n610), .Z(n103) );
  MUX2_X1 U703 ( .A(n103), .B(n100), .S(n606), .Z(n104) );
  MUX2_X1 U704 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U705 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n612), .Z(n106) );
  MUX2_X1 U706 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n612), .Z(n107) );
  MUX2_X1 U707 ( .A(n107), .B(n106), .S(n610), .Z(n108) );
  MUX2_X1 U708 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n612), .Z(n109) );
  MUX2_X1 U709 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n612), .Z(n110) );
  MUX2_X1 U710 ( .A(n110), .B(n109), .S(n610), .Z(n111) );
  MUX2_X1 U711 ( .A(n111), .B(n108), .S(n606), .Z(n112) );
  MUX2_X1 U712 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n612), .Z(n113) );
  MUX2_X1 U713 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n612), .Z(n114) );
  MUX2_X1 U714 ( .A(n114), .B(n113), .S(n608), .Z(n115) );
  MUX2_X1 U715 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n612), .Z(n116) );
  MUX2_X1 U716 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n612), .Z(n117) );
  MUX2_X1 U717 ( .A(n117), .B(n116), .S(n609), .Z(n118) );
  MUX2_X1 U718 ( .A(n118), .B(n115), .S(n606), .Z(n119) );
  MUX2_X1 U719 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U720 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U721 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n612), .Z(n121) );
  MUX2_X1 U722 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n612), .Z(n122) );
  MUX2_X1 U723 ( .A(n122), .B(n121), .S(n608), .Z(n123) );
  MUX2_X1 U724 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n612), .Z(n124) );
  MUX2_X1 U725 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n612), .Z(n125) );
  MUX2_X1 U726 ( .A(n125), .B(n124), .S(n608), .Z(n126) );
  MUX2_X1 U727 ( .A(n126), .B(n123), .S(n606), .Z(n127) );
  MUX2_X1 U728 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n613), .Z(n128) );
  MUX2_X1 U729 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n613), .Z(n129) );
  MUX2_X1 U730 ( .A(n129), .B(n128), .S(n609), .Z(n130) );
  MUX2_X1 U731 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n613), .Z(n131) );
  MUX2_X1 U732 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n613), .Z(n132) );
  MUX2_X1 U733 ( .A(n132), .B(n131), .S(n609), .Z(n133) );
  MUX2_X1 U734 ( .A(n133), .B(n130), .S(n606), .Z(n134) );
  MUX2_X1 U735 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U736 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n613), .Z(n136) );
  MUX2_X1 U737 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n613), .Z(n137) );
  MUX2_X1 U738 ( .A(n137), .B(n136), .S(n610), .Z(n138) );
  MUX2_X1 U739 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n613), .Z(n139) );
  MUX2_X1 U740 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n613), .Z(n140) );
  MUX2_X1 U741 ( .A(n140), .B(n139), .S(n608), .Z(n141) );
  MUX2_X1 U742 ( .A(n141), .B(n138), .S(n606), .Z(n142) );
  MUX2_X1 U743 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n613), .Z(n143) );
  MUX2_X1 U744 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n613), .Z(n144) );
  MUX2_X1 U745 ( .A(n144), .B(n143), .S(n609), .Z(n145) );
  MUX2_X1 U746 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n613), .Z(n146) );
  MUX2_X1 U747 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n613), .Z(n147) );
  MUX2_X1 U748 ( .A(n147), .B(n146), .S(n610), .Z(n148) );
  MUX2_X1 U749 ( .A(n148), .B(n145), .S(n606), .Z(n149) );
  MUX2_X1 U750 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U751 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U752 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n614), .Z(n151) );
  MUX2_X1 U753 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n614), .Z(n152) );
  MUX2_X1 U754 ( .A(n152), .B(n151), .S(n609), .Z(n153) );
  MUX2_X1 U755 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n614), .Z(n154) );
  MUX2_X1 U756 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n614), .Z(n155) );
  MUX2_X1 U757 ( .A(n155), .B(n154), .S(n610), .Z(n156) );
  MUX2_X1 U758 ( .A(n156), .B(n153), .S(n607), .Z(n157) );
  MUX2_X1 U759 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n614), .Z(n158) );
  MUX2_X1 U760 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n614), .Z(n159) );
  MUX2_X1 U761 ( .A(n159), .B(n158), .S(N11), .Z(n160) );
  MUX2_X1 U762 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n614), .Z(n161) );
  MUX2_X1 U763 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n614), .Z(n162) );
  MUX2_X1 U764 ( .A(n162), .B(n161), .S(n608), .Z(n163) );
  MUX2_X1 U765 ( .A(n163), .B(n160), .S(n607), .Z(n164) );
  MUX2_X1 U766 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U767 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n614), .Z(n166) );
  MUX2_X1 U768 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n614), .Z(n167) );
  MUX2_X1 U769 ( .A(n167), .B(n166), .S(n608), .Z(n168) );
  MUX2_X1 U770 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n614), .Z(n169) );
  MUX2_X1 U771 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n614), .Z(n170) );
  MUX2_X1 U772 ( .A(n170), .B(n169), .S(N11), .Z(n171) );
  MUX2_X1 U773 ( .A(n171), .B(n168), .S(n607), .Z(n172) );
  MUX2_X1 U774 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n617), .Z(n173) );
  MUX2_X1 U775 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(N10), .Z(n174) );
  MUX2_X1 U776 ( .A(n174), .B(n173), .S(n609), .Z(n175) );
  MUX2_X1 U777 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n176) );
  MUX2_X1 U778 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n177) );
  MUX2_X1 U779 ( .A(n177), .B(n176), .S(n609), .Z(n178) );
  MUX2_X1 U780 ( .A(n178), .B(n175), .S(n607), .Z(n179) );
  MUX2_X1 U781 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U782 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U783 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n611), .Z(n181) );
  MUX2_X1 U784 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n611), .Z(n182) );
  MUX2_X1 U785 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U786 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n611), .Z(n184) );
  MUX2_X1 U787 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n612), .Z(n185) );
  MUX2_X1 U788 ( .A(n185), .B(n184), .S(N11), .Z(n186) );
  MUX2_X1 U789 ( .A(n186), .B(n183), .S(n607), .Z(n187) );
  MUX2_X1 U790 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n611), .Z(n188) );
  MUX2_X1 U791 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n617), .Z(n189) );
  MUX2_X1 U792 ( .A(n189), .B(n188), .S(n610), .Z(n190) );
  MUX2_X1 U793 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n617), .Z(n191) );
  MUX2_X1 U794 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(N10), .Z(n192) );
  MUX2_X1 U795 ( .A(n192), .B(n191), .S(N11), .Z(n193) );
  MUX2_X1 U796 ( .A(n193), .B(n190), .S(n607), .Z(n194) );
  MUX2_X1 U797 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U798 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n615), .Z(n196) );
  MUX2_X1 U799 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n615), .Z(n197) );
  MUX2_X1 U800 ( .A(n197), .B(n196), .S(n608), .Z(n198) );
  MUX2_X1 U801 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n615), .Z(n199) );
  MUX2_X1 U802 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n615), .Z(n200) );
  MUX2_X1 U803 ( .A(n200), .B(n199), .S(n610), .Z(n201) );
  MUX2_X1 U804 ( .A(n201), .B(n198), .S(n607), .Z(n202) );
  MUX2_X1 U805 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n615), .Z(n203) );
  MUX2_X1 U806 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n615), .Z(n204) );
  MUX2_X1 U807 ( .A(n204), .B(n203), .S(n608), .Z(n205) );
  MUX2_X1 U808 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n615), .Z(n206) );
  MUX2_X1 U809 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n615), .Z(n207) );
  MUX2_X1 U810 ( .A(n207), .B(n206), .S(n610), .Z(n208) );
  MUX2_X1 U811 ( .A(n208), .B(n205), .S(n607), .Z(n209) );
  MUX2_X1 U812 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U813 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U814 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n615), .Z(n211) );
  MUX2_X1 U815 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n615), .Z(n212) );
  MUX2_X1 U816 ( .A(n212), .B(n211), .S(n608), .Z(n213) );
  MUX2_X1 U817 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n615), .Z(n214) );
  MUX2_X1 U818 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n615), .Z(n215) );
  MUX2_X1 U819 ( .A(n215), .B(n214), .S(n608), .Z(n216) );
  MUX2_X1 U820 ( .A(n216), .B(n213), .S(n607), .Z(n217) );
  MUX2_X1 U821 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n616), .Z(n218) );
  MUX2_X1 U822 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n616), .Z(n219) );
  MUX2_X1 U823 ( .A(n219), .B(n218), .S(n608), .Z(n220) );
  MUX2_X1 U824 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n616), .Z(n221) );
  MUX2_X1 U825 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n616), .Z(n222) );
  MUX2_X1 U826 ( .A(n222), .B(n221), .S(n609), .Z(n223) );
  MUX2_X1 U827 ( .A(n223), .B(n220), .S(n607), .Z(n224) );
  MUX2_X1 U828 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U829 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n616), .Z(n226) );
  MUX2_X1 U830 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n616), .Z(n227) );
  MUX2_X1 U831 ( .A(n227), .B(n226), .S(n608), .Z(n228) );
  MUX2_X1 U832 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n616), .Z(n229) );
  MUX2_X1 U833 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n616), .Z(n595) );
  MUX2_X1 U834 ( .A(n595), .B(n229), .S(n610), .Z(n596) );
  MUX2_X1 U835 ( .A(n596), .B(n228), .S(n607), .Z(n597) );
  MUX2_X1 U836 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n616), .Z(n598) );
  MUX2_X1 U837 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n616), .Z(n599) );
  MUX2_X1 U838 ( .A(n599), .B(n598), .S(n608), .Z(n600) );
  MUX2_X1 U839 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n616), .Z(n601) );
  MUX2_X1 U840 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n616), .Z(n602) );
  MUX2_X1 U841 ( .A(n602), .B(n601), .S(n608), .Z(n603) );
  MUX2_X1 U842 ( .A(n603), .B(n600), .S(n607), .Z(n604) );
  MUX2_X1 U843 ( .A(n604), .B(n597), .S(N13), .Z(n605) );
  MUX2_X1 U844 ( .A(n605), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U845 ( .A(N11), .Z(n608) );
  CLKBUF_X1 U846 ( .A(n617), .Z(n611) );
  INV_X1 U847 ( .A(N10), .ZN(n618) );
  INV_X1 U848 ( .A(N11), .ZN(n619) );
  INV_X1 U849 ( .A(data_in[0]), .ZN(n620) );
  INV_X1 U850 ( .A(data_in[1]), .ZN(n621) );
  INV_X1 U851 ( .A(data_in[2]), .ZN(n622) );
  INV_X1 U852 ( .A(data_in[3]), .ZN(n623) );
  INV_X1 U853 ( .A(data_in[4]), .ZN(n624) );
  INV_X1 U854 ( .A(data_in[5]), .ZN(n625) );
  INV_X1 U855 ( .A(data_in[6]), .ZN(n626) );
  INV_X1 U856 ( .A(data_in[7]), .ZN(n627) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_27 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n627), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n628), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n629), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n630), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n631), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n632), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n633), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n634), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n635), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n636), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n637), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n638), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n639), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n640), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n641), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n642), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n643), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n644), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n645), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n646), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n647), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n648), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n649), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n650), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n651), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n652), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n653), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n654), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n655), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n656), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n657), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n658), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n659), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n660), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n661), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n662), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n663), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n664), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n665), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n666), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n667), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n668), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n669), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n670), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n671), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n672), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n673), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n674), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n675), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n676), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n677), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n678), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n679), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n680), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n681), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n682), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n683), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n684), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n685), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n686), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n687), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n688), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n689), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n690), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n691), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n692), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n693), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n694), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n695), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n696), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n697), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n698), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n699), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n700), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n701), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n702), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n703), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n704), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n705), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n706), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n707), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n708), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n709), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n710), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n711), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n712), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n713), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n714), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n715), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n716), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n717), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n718), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n719), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n720), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n721), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n722), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n723), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n724), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n725), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n726), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n727), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n728), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n729), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n730), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n731), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n732), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n733), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n734), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n735), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n736), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n737), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n738), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n739), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n740), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n741), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n742), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n743), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n744), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n745), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n746), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n747), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n748), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n749), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n750), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n751), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n752), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n753), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n754), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n755), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n756), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n757), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n758), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n759), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n760), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n761), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n762), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n763), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n764), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n765), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n766), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n767), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n768), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n769), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n770), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n771), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n772), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n773), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n774), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n775), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n776), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n777), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n778), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n779), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n780), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n781), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n782), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n783), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n784), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n785), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n786), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n787), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n788), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n789), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n790), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n791), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n792), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n793), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n794), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n795), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n796), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n797), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n798), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n799), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n800), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n801), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n802), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n803), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n804), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n805), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n806), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n807), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n808), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n809), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n810), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n811), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n812), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n813), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n814), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n815), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n816), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n817), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n818), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n846), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n847), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n848), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n849), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n850), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n851), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n852), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n853), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n854), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n855), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n856), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n857), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n858), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n859), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n860), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n861), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n862), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n863), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n864), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n865), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n866), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n867), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n868), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n869), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n870), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n871), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n872), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n873), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n874), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n875), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n876), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n877), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n878), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n879), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n880), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n881), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n882), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n883), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n884), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n885), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n886), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n887), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n888), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n889), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n890), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n891), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n892), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n893), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n894), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n895), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n896), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n897), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n898), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n899), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n900), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n901), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n902), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n903), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n904), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n905), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n906), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n907), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n908), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n909), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n616), .Z(n611) );
  BUF_X1 U4 ( .A(n616), .Z(n614) );
  BUF_X1 U5 ( .A(n616), .Z(n615) );
  BUF_X1 U6 ( .A(N10), .Z(n612) );
  BUF_X1 U7 ( .A(n616), .Z(n613) );
  BUF_X1 U8 ( .A(N11), .Z(n609) );
  BUF_X1 U9 ( .A(N11), .Z(n610) );
  BUF_X1 U10 ( .A(N10), .Z(n616) );
  NOR3_X1 U11 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1201) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(n617), .ZN(n1190) );
  NOR3_X1 U13 ( .A1(N10), .A2(N12), .A3(n618), .ZN(n1180) );
  NOR3_X1 U14 ( .A1(n617), .A2(N12), .A3(n618), .ZN(n1170) );
  INV_X1 U15 ( .A(n1127), .ZN(n842) );
  INV_X1 U16 ( .A(n1117), .ZN(n841) );
  INV_X1 U17 ( .A(n1108), .ZN(n840) );
  INV_X1 U18 ( .A(n1099), .ZN(n839) );
  INV_X1 U19 ( .A(n1054), .ZN(n834) );
  INV_X1 U20 ( .A(n1044), .ZN(n833) );
  INV_X1 U21 ( .A(n1035), .ZN(n832) );
  INV_X1 U22 ( .A(n1026), .ZN(n831) );
  INV_X1 U23 ( .A(n981), .ZN(n826) );
  INV_X1 U24 ( .A(n971), .ZN(n825) );
  INV_X1 U25 ( .A(n962), .ZN(n824) );
  INV_X1 U26 ( .A(n953), .ZN(n823) );
  INV_X1 U27 ( .A(n1090), .ZN(n838) );
  INV_X1 U28 ( .A(n1081), .ZN(n837) );
  INV_X1 U29 ( .A(n1072), .ZN(n836) );
  INV_X1 U30 ( .A(n1063), .ZN(n835) );
  INV_X1 U31 ( .A(n944), .ZN(n822) );
  INV_X1 U32 ( .A(n935), .ZN(n821) );
  INV_X1 U33 ( .A(n926), .ZN(n820) );
  INV_X1 U34 ( .A(n917), .ZN(n819) );
  INV_X1 U35 ( .A(n1017), .ZN(n830) );
  INV_X1 U36 ( .A(n1008), .ZN(n829) );
  INV_X1 U37 ( .A(n999), .ZN(n828) );
  INV_X1 U38 ( .A(n990), .ZN(n827) );
  BUF_X1 U39 ( .A(N12), .Z(n606) );
  BUF_X1 U40 ( .A(N12), .Z(n607) );
  INV_X1 U41 ( .A(N13), .ZN(n844) );
  AND3_X1 U42 ( .A1(n617), .A2(n618), .A3(N12), .ZN(n1160) );
  AND3_X1 U43 ( .A1(N10), .A2(n618), .A3(N12), .ZN(n1150) );
  AND3_X1 U44 ( .A1(N11), .A2(n617), .A3(N12), .ZN(n1140) );
  AND3_X1 U45 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1130) );
  INV_X1 U46 ( .A(N14), .ZN(n845) );
  NAND2_X1 U47 ( .A1(n1190), .A2(n1200), .ZN(n1199) );
  NAND2_X1 U48 ( .A1(n1180), .A2(n1200), .ZN(n1189) );
  NAND2_X1 U49 ( .A1(n1170), .A2(n1200), .ZN(n1179) );
  NAND2_X1 U50 ( .A1(n1160), .A2(n1200), .ZN(n1169) );
  NAND2_X1 U51 ( .A1(n1150), .A2(n1200), .ZN(n1159) );
  NAND2_X1 U52 ( .A1(n1140), .A2(n1200), .ZN(n1149) );
  NAND2_X1 U53 ( .A1(n1130), .A2(n1200), .ZN(n1139) );
  NAND2_X1 U54 ( .A1(n1201), .A2(n1200), .ZN(n1210) );
  NAND2_X1 U55 ( .A1(n1119), .A2(n1201), .ZN(n1127) );
  NAND2_X1 U56 ( .A1(n1119), .A2(n1190), .ZN(n1117) );
  NAND2_X1 U57 ( .A1(n1119), .A2(n1180), .ZN(n1108) );
  NAND2_X1 U58 ( .A1(n1119), .A2(n1170), .ZN(n1099) );
  NAND2_X1 U59 ( .A1(n1046), .A2(n1201), .ZN(n1054) );
  NAND2_X1 U60 ( .A1(n1046), .A2(n1190), .ZN(n1044) );
  NAND2_X1 U61 ( .A1(n1046), .A2(n1180), .ZN(n1035) );
  NAND2_X1 U62 ( .A1(n1046), .A2(n1170), .ZN(n1026) );
  NAND2_X1 U63 ( .A1(n973), .A2(n1201), .ZN(n981) );
  NAND2_X1 U64 ( .A1(n973), .A2(n1190), .ZN(n971) );
  NAND2_X1 U65 ( .A1(n973), .A2(n1180), .ZN(n962) );
  NAND2_X1 U66 ( .A1(n973), .A2(n1170), .ZN(n953) );
  NAND2_X1 U67 ( .A1(n1119), .A2(n1160), .ZN(n1090) );
  NAND2_X1 U68 ( .A1(n1119), .A2(n1150), .ZN(n1081) );
  NAND2_X1 U69 ( .A1(n1119), .A2(n1140), .ZN(n1072) );
  NAND2_X1 U70 ( .A1(n1119), .A2(n1130), .ZN(n1063) );
  NAND2_X1 U71 ( .A1(n1046), .A2(n1160), .ZN(n1017) );
  NAND2_X1 U72 ( .A1(n1046), .A2(n1150), .ZN(n1008) );
  NAND2_X1 U73 ( .A1(n1046), .A2(n1140), .ZN(n999) );
  NAND2_X1 U74 ( .A1(n1046), .A2(n1130), .ZN(n990) );
  NAND2_X1 U75 ( .A1(n973), .A2(n1160), .ZN(n944) );
  NAND2_X1 U76 ( .A1(n973), .A2(n1150), .ZN(n935) );
  NAND2_X1 U77 ( .A1(n973), .A2(n1140), .ZN(n926) );
  NAND2_X1 U78 ( .A1(n973), .A2(n1130), .ZN(n917) );
  AND3_X1 U79 ( .A1(n844), .A2(n845), .A3(n1129), .ZN(n1200) );
  AND3_X1 U80 ( .A1(N13), .A2(n1129), .A3(N14), .ZN(n973) );
  AND3_X1 U81 ( .A1(n1129), .A2(n845), .A3(N13), .ZN(n1119) );
  AND3_X1 U82 ( .A1(n1129), .A2(n844), .A3(N14), .ZN(n1046) );
  NOR2_X1 U83 ( .A1(n843), .A2(addr[5]), .ZN(n1129) );
  INV_X1 U84 ( .A(wr_en), .ZN(n843) );
  OAI21_X1 U85 ( .B1(n619), .B2(n1169), .A(n1168), .ZN(n877) );
  NAND2_X1 U86 ( .A1(\mem[4][0] ), .A2(n1169), .ZN(n1168) );
  OAI21_X1 U87 ( .B1(n620), .B2(n1169), .A(n1167), .ZN(n876) );
  NAND2_X1 U88 ( .A1(\mem[4][1] ), .A2(n1169), .ZN(n1167) );
  OAI21_X1 U89 ( .B1(n621), .B2(n1169), .A(n1166), .ZN(n875) );
  NAND2_X1 U90 ( .A1(\mem[4][2] ), .A2(n1169), .ZN(n1166) );
  OAI21_X1 U91 ( .B1(n622), .B2(n1169), .A(n1165), .ZN(n874) );
  NAND2_X1 U92 ( .A1(\mem[4][3] ), .A2(n1169), .ZN(n1165) );
  OAI21_X1 U93 ( .B1(n623), .B2(n1169), .A(n1164), .ZN(n873) );
  NAND2_X1 U94 ( .A1(\mem[4][4] ), .A2(n1169), .ZN(n1164) );
  OAI21_X1 U95 ( .B1(n624), .B2(n1169), .A(n1163), .ZN(n872) );
  NAND2_X1 U96 ( .A1(\mem[4][5] ), .A2(n1169), .ZN(n1163) );
  OAI21_X1 U97 ( .B1(n625), .B2(n1169), .A(n1162), .ZN(n871) );
  NAND2_X1 U98 ( .A1(\mem[4][6] ), .A2(n1169), .ZN(n1162) );
  OAI21_X1 U99 ( .B1(n626), .B2(n1169), .A(n1161), .ZN(n870) );
  NAND2_X1 U100 ( .A1(\mem[4][7] ), .A2(n1169), .ZN(n1161) );
  OAI21_X1 U101 ( .B1(n619), .B2(n1149), .A(n1148), .ZN(n861) );
  NAND2_X1 U102 ( .A1(\mem[6][0] ), .A2(n1149), .ZN(n1148) );
  OAI21_X1 U103 ( .B1(n620), .B2(n1149), .A(n1147), .ZN(n860) );
  NAND2_X1 U104 ( .A1(\mem[6][1] ), .A2(n1149), .ZN(n1147) );
  OAI21_X1 U105 ( .B1(n621), .B2(n1149), .A(n1146), .ZN(n859) );
  NAND2_X1 U106 ( .A1(\mem[6][2] ), .A2(n1149), .ZN(n1146) );
  OAI21_X1 U107 ( .B1(n622), .B2(n1149), .A(n1145), .ZN(n858) );
  NAND2_X1 U108 ( .A1(\mem[6][3] ), .A2(n1149), .ZN(n1145) );
  OAI21_X1 U109 ( .B1(n623), .B2(n1149), .A(n1144), .ZN(n857) );
  NAND2_X1 U110 ( .A1(\mem[6][4] ), .A2(n1149), .ZN(n1144) );
  OAI21_X1 U111 ( .B1(n624), .B2(n1149), .A(n1143), .ZN(n856) );
  NAND2_X1 U112 ( .A1(\mem[6][5] ), .A2(n1149), .ZN(n1143) );
  OAI21_X1 U113 ( .B1(n625), .B2(n1149), .A(n1142), .ZN(n855) );
  NAND2_X1 U114 ( .A1(\mem[6][6] ), .A2(n1149), .ZN(n1142) );
  OAI21_X1 U115 ( .B1(n626), .B2(n1149), .A(n1141), .ZN(n854) );
  NAND2_X1 U116 ( .A1(\mem[6][7] ), .A2(n1149), .ZN(n1141) );
  OAI21_X1 U117 ( .B1(n619), .B2(n1139), .A(n1138), .ZN(n853) );
  NAND2_X1 U118 ( .A1(\mem[7][0] ), .A2(n1139), .ZN(n1138) );
  OAI21_X1 U119 ( .B1(n620), .B2(n1139), .A(n1137), .ZN(n852) );
  NAND2_X1 U120 ( .A1(\mem[7][1] ), .A2(n1139), .ZN(n1137) );
  OAI21_X1 U121 ( .B1(n621), .B2(n1139), .A(n1136), .ZN(n851) );
  NAND2_X1 U122 ( .A1(\mem[7][2] ), .A2(n1139), .ZN(n1136) );
  OAI21_X1 U123 ( .B1(n622), .B2(n1139), .A(n1135), .ZN(n850) );
  NAND2_X1 U124 ( .A1(\mem[7][3] ), .A2(n1139), .ZN(n1135) );
  OAI21_X1 U125 ( .B1(n623), .B2(n1139), .A(n1134), .ZN(n849) );
  NAND2_X1 U126 ( .A1(\mem[7][4] ), .A2(n1139), .ZN(n1134) );
  OAI21_X1 U127 ( .B1(n624), .B2(n1139), .A(n1133), .ZN(n848) );
  NAND2_X1 U128 ( .A1(\mem[7][5] ), .A2(n1139), .ZN(n1133) );
  OAI21_X1 U129 ( .B1(n625), .B2(n1139), .A(n1132), .ZN(n847) );
  NAND2_X1 U130 ( .A1(\mem[7][6] ), .A2(n1139), .ZN(n1132) );
  OAI21_X1 U131 ( .B1(n626), .B2(n1139), .A(n1131), .ZN(n846) );
  NAND2_X1 U132 ( .A1(\mem[7][7] ), .A2(n1139), .ZN(n1131) );
  OAI21_X1 U133 ( .B1(n619), .B2(n1199), .A(n1198), .ZN(n901) );
  NAND2_X1 U134 ( .A1(\mem[1][0] ), .A2(n1199), .ZN(n1198) );
  OAI21_X1 U135 ( .B1(n620), .B2(n1199), .A(n1197), .ZN(n900) );
  NAND2_X1 U136 ( .A1(\mem[1][1] ), .A2(n1199), .ZN(n1197) );
  OAI21_X1 U137 ( .B1(n621), .B2(n1199), .A(n1196), .ZN(n899) );
  NAND2_X1 U138 ( .A1(\mem[1][2] ), .A2(n1199), .ZN(n1196) );
  OAI21_X1 U139 ( .B1(n622), .B2(n1199), .A(n1195), .ZN(n898) );
  NAND2_X1 U140 ( .A1(\mem[1][3] ), .A2(n1199), .ZN(n1195) );
  OAI21_X1 U141 ( .B1(n623), .B2(n1199), .A(n1194), .ZN(n897) );
  NAND2_X1 U142 ( .A1(\mem[1][4] ), .A2(n1199), .ZN(n1194) );
  OAI21_X1 U143 ( .B1(n624), .B2(n1199), .A(n1193), .ZN(n896) );
  NAND2_X1 U144 ( .A1(\mem[1][5] ), .A2(n1199), .ZN(n1193) );
  OAI21_X1 U145 ( .B1(n625), .B2(n1199), .A(n1192), .ZN(n895) );
  NAND2_X1 U146 ( .A1(\mem[1][6] ), .A2(n1199), .ZN(n1192) );
  OAI21_X1 U147 ( .B1(n626), .B2(n1199), .A(n1191), .ZN(n894) );
  NAND2_X1 U148 ( .A1(\mem[1][7] ), .A2(n1199), .ZN(n1191) );
  OAI21_X1 U149 ( .B1(n619), .B2(n1189), .A(n1188), .ZN(n893) );
  NAND2_X1 U150 ( .A1(\mem[2][0] ), .A2(n1189), .ZN(n1188) );
  OAI21_X1 U151 ( .B1(n620), .B2(n1189), .A(n1187), .ZN(n892) );
  NAND2_X1 U152 ( .A1(\mem[2][1] ), .A2(n1189), .ZN(n1187) );
  OAI21_X1 U153 ( .B1(n621), .B2(n1189), .A(n1186), .ZN(n891) );
  NAND2_X1 U154 ( .A1(\mem[2][2] ), .A2(n1189), .ZN(n1186) );
  OAI21_X1 U155 ( .B1(n622), .B2(n1189), .A(n1185), .ZN(n890) );
  NAND2_X1 U156 ( .A1(\mem[2][3] ), .A2(n1189), .ZN(n1185) );
  OAI21_X1 U157 ( .B1(n623), .B2(n1189), .A(n1184), .ZN(n889) );
  NAND2_X1 U158 ( .A1(\mem[2][4] ), .A2(n1189), .ZN(n1184) );
  OAI21_X1 U159 ( .B1(n624), .B2(n1189), .A(n1183), .ZN(n888) );
  NAND2_X1 U160 ( .A1(\mem[2][5] ), .A2(n1189), .ZN(n1183) );
  OAI21_X1 U161 ( .B1(n625), .B2(n1189), .A(n1182), .ZN(n887) );
  NAND2_X1 U162 ( .A1(\mem[2][6] ), .A2(n1189), .ZN(n1182) );
  OAI21_X1 U163 ( .B1(n626), .B2(n1189), .A(n1181), .ZN(n886) );
  NAND2_X1 U164 ( .A1(\mem[2][7] ), .A2(n1189), .ZN(n1181) );
  OAI21_X1 U165 ( .B1(n619), .B2(n1179), .A(n1178), .ZN(n885) );
  NAND2_X1 U166 ( .A1(\mem[3][0] ), .A2(n1179), .ZN(n1178) );
  OAI21_X1 U167 ( .B1(n620), .B2(n1179), .A(n1177), .ZN(n884) );
  NAND2_X1 U168 ( .A1(\mem[3][1] ), .A2(n1179), .ZN(n1177) );
  OAI21_X1 U169 ( .B1(n621), .B2(n1179), .A(n1176), .ZN(n883) );
  NAND2_X1 U170 ( .A1(\mem[3][2] ), .A2(n1179), .ZN(n1176) );
  OAI21_X1 U171 ( .B1(n622), .B2(n1179), .A(n1175), .ZN(n882) );
  NAND2_X1 U172 ( .A1(\mem[3][3] ), .A2(n1179), .ZN(n1175) );
  OAI21_X1 U173 ( .B1(n623), .B2(n1179), .A(n1174), .ZN(n881) );
  NAND2_X1 U174 ( .A1(\mem[3][4] ), .A2(n1179), .ZN(n1174) );
  OAI21_X1 U175 ( .B1(n624), .B2(n1179), .A(n1173), .ZN(n880) );
  NAND2_X1 U176 ( .A1(\mem[3][5] ), .A2(n1179), .ZN(n1173) );
  OAI21_X1 U177 ( .B1(n625), .B2(n1179), .A(n1172), .ZN(n879) );
  NAND2_X1 U178 ( .A1(\mem[3][6] ), .A2(n1179), .ZN(n1172) );
  OAI21_X1 U179 ( .B1(n626), .B2(n1179), .A(n1171), .ZN(n878) );
  NAND2_X1 U180 ( .A1(\mem[3][7] ), .A2(n1179), .ZN(n1171) );
  OAI21_X1 U181 ( .B1(n619), .B2(n1159), .A(n1158), .ZN(n869) );
  NAND2_X1 U182 ( .A1(\mem[5][0] ), .A2(n1159), .ZN(n1158) );
  OAI21_X1 U183 ( .B1(n620), .B2(n1159), .A(n1157), .ZN(n868) );
  NAND2_X1 U184 ( .A1(\mem[5][1] ), .A2(n1159), .ZN(n1157) );
  OAI21_X1 U185 ( .B1(n621), .B2(n1159), .A(n1156), .ZN(n867) );
  NAND2_X1 U186 ( .A1(\mem[5][2] ), .A2(n1159), .ZN(n1156) );
  OAI21_X1 U187 ( .B1(n622), .B2(n1159), .A(n1155), .ZN(n866) );
  NAND2_X1 U188 ( .A1(\mem[5][3] ), .A2(n1159), .ZN(n1155) );
  OAI21_X1 U189 ( .B1(n623), .B2(n1159), .A(n1154), .ZN(n865) );
  NAND2_X1 U190 ( .A1(\mem[5][4] ), .A2(n1159), .ZN(n1154) );
  OAI21_X1 U191 ( .B1(n624), .B2(n1159), .A(n1153), .ZN(n864) );
  NAND2_X1 U192 ( .A1(\mem[5][5] ), .A2(n1159), .ZN(n1153) );
  OAI21_X1 U193 ( .B1(n625), .B2(n1159), .A(n1152), .ZN(n863) );
  NAND2_X1 U194 ( .A1(\mem[5][6] ), .A2(n1159), .ZN(n1152) );
  OAI21_X1 U195 ( .B1(n626), .B2(n1159), .A(n1151), .ZN(n862) );
  NAND2_X1 U196 ( .A1(\mem[5][7] ), .A2(n1159), .ZN(n1151) );
  OAI21_X1 U197 ( .B1(n1210), .B2(n619), .A(n1209), .ZN(n909) );
  NAND2_X1 U198 ( .A1(\mem[0][0] ), .A2(n1210), .ZN(n1209) );
  OAI21_X1 U199 ( .B1(n1210), .B2(n620), .A(n1208), .ZN(n908) );
  NAND2_X1 U200 ( .A1(\mem[0][1] ), .A2(n1210), .ZN(n1208) );
  OAI21_X1 U201 ( .B1(n1210), .B2(n621), .A(n1207), .ZN(n907) );
  NAND2_X1 U202 ( .A1(\mem[0][2] ), .A2(n1210), .ZN(n1207) );
  OAI21_X1 U203 ( .B1(n1210), .B2(n622), .A(n1206), .ZN(n906) );
  NAND2_X1 U204 ( .A1(\mem[0][3] ), .A2(n1210), .ZN(n1206) );
  OAI21_X1 U205 ( .B1(n1210), .B2(n623), .A(n1205), .ZN(n905) );
  NAND2_X1 U206 ( .A1(\mem[0][4] ), .A2(n1210), .ZN(n1205) );
  OAI21_X1 U207 ( .B1(n1210), .B2(n624), .A(n1204), .ZN(n904) );
  NAND2_X1 U208 ( .A1(\mem[0][5] ), .A2(n1210), .ZN(n1204) );
  OAI21_X1 U209 ( .B1(n1210), .B2(n625), .A(n1203), .ZN(n903) );
  NAND2_X1 U210 ( .A1(\mem[0][6] ), .A2(n1210), .ZN(n1203) );
  OAI21_X1 U211 ( .B1(n1210), .B2(n626), .A(n1202), .ZN(n902) );
  NAND2_X1 U212 ( .A1(\mem[0][7] ), .A2(n1210), .ZN(n1202) );
  INV_X1 U213 ( .A(n1128), .ZN(n818) );
  AOI22_X1 U214 ( .A1(data_in[0]), .A2(n842), .B1(n1127), .B2(\mem[8][0] ), 
        .ZN(n1128) );
  INV_X1 U215 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U216 ( .A1(data_in[1]), .A2(n842), .B1(n1127), .B2(\mem[8][1] ), 
        .ZN(n1126) );
  INV_X1 U217 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U218 ( .A1(data_in[2]), .A2(n842), .B1(n1127), .B2(\mem[8][2] ), 
        .ZN(n1125) );
  INV_X1 U219 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U220 ( .A1(data_in[3]), .A2(n842), .B1(n1127), .B2(\mem[8][3] ), 
        .ZN(n1124) );
  INV_X1 U221 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U222 ( .A1(data_in[4]), .A2(n842), .B1(n1127), .B2(\mem[8][4] ), 
        .ZN(n1123) );
  INV_X1 U223 ( .A(n1122), .ZN(n813) );
  AOI22_X1 U224 ( .A1(data_in[5]), .A2(n842), .B1(n1127), .B2(\mem[8][5] ), 
        .ZN(n1122) );
  INV_X1 U225 ( .A(n1121), .ZN(n812) );
  AOI22_X1 U226 ( .A1(data_in[6]), .A2(n842), .B1(n1127), .B2(\mem[8][6] ), 
        .ZN(n1121) );
  INV_X1 U227 ( .A(n1120), .ZN(n811) );
  AOI22_X1 U228 ( .A1(data_in[7]), .A2(n842), .B1(n1127), .B2(\mem[8][7] ), 
        .ZN(n1120) );
  INV_X1 U229 ( .A(n1118), .ZN(n810) );
  AOI22_X1 U230 ( .A1(data_in[0]), .A2(n841), .B1(n1117), .B2(\mem[9][0] ), 
        .ZN(n1118) );
  INV_X1 U231 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U232 ( .A1(data_in[1]), .A2(n841), .B1(n1117), .B2(\mem[9][1] ), 
        .ZN(n1116) );
  INV_X1 U233 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U234 ( .A1(data_in[2]), .A2(n841), .B1(n1117), .B2(\mem[9][2] ), 
        .ZN(n1115) );
  INV_X1 U235 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U236 ( .A1(data_in[3]), .A2(n841), .B1(n1117), .B2(\mem[9][3] ), 
        .ZN(n1114) );
  INV_X1 U237 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U238 ( .A1(data_in[4]), .A2(n841), .B1(n1117), .B2(\mem[9][4] ), 
        .ZN(n1113) );
  INV_X1 U239 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U240 ( .A1(data_in[5]), .A2(n841), .B1(n1117), .B2(\mem[9][5] ), 
        .ZN(n1112) );
  INV_X1 U241 ( .A(n1111), .ZN(n804) );
  AOI22_X1 U242 ( .A1(data_in[6]), .A2(n841), .B1(n1117), .B2(\mem[9][6] ), 
        .ZN(n1111) );
  INV_X1 U243 ( .A(n1110), .ZN(n803) );
  AOI22_X1 U244 ( .A1(data_in[7]), .A2(n841), .B1(n1117), .B2(\mem[9][7] ), 
        .ZN(n1110) );
  INV_X1 U245 ( .A(n1109), .ZN(n802) );
  AOI22_X1 U246 ( .A1(data_in[0]), .A2(n840), .B1(n1108), .B2(\mem[10][0] ), 
        .ZN(n1109) );
  INV_X1 U247 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U248 ( .A1(data_in[1]), .A2(n840), .B1(n1108), .B2(\mem[10][1] ), 
        .ZN(n1107) );
  INV_X1 U249 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U250 ( .A1(data_in[2]), .A2(n840), .B1(n1108), .B2(\mem[10][2] ), 
        .ZN(n1106) );
  INV_X1 U251 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U252 ( .A1(data_in[3]), .A2(n840), .B1(n1108), .B2(\mem[10][3] ), 
        .ZN(n1105) );
  INV_X1 U253 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U254 ( .A1(data_in[4]), .A2(n840), .B1(n1108), .B2(\mem[10][4] ), 
        .ZN(n1104) );
  INV_X1 U255 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U256 ( .A1(data_in[5]), .A2(n840), .B1(n1108), .B2(\mem[10][5] ), 
        .ZN(n1103) );
  INV_X1 U257 ( .A(n1102), .ZN(n796) );
  AOI22_X1 U258 ( .A1(data_in[6]), .A2(n840), .B1(n1108), .B2(\mem[10][6] ), 
        .ZN(n1102) );
  INV_X1 U259 ( .A(n1101), .ZN(n795) );
  AOI22_X1 U260 ( .A1(data_in[7]), .A2(n840), .B1(n1108), .B2(\mem[10][7] ), 
        .ZN(n1101) );
  INV_X1 U261 ( .A(n1100), .ZN(n794) );
  AOI22_X1 U262 ( .A1(data_in[0]), .A2(n839), .B1(n1099), .B2(\mem[11][0] ), 
        .ZN(n1100) );
  INV_X1 U263 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U264 ( .A1(data_in[1]), .A2(n839), .B1(n1099), .B2(\mem[11][1] ), 
        .ZN(n1098) );
  INV_X1 U265 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U266 ( .A1(data_in[2]), .A2(n839), .B1(n1099), .B2(\mem[11][2] ), 
        .ZN(n1097) );
  INV_X1 U267 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U268 ( .A1(data_in[3]), .A2(n839), .B1(n1099), .B2(\mem[11][3] ), 
        .ZN(n1096) );
  INV_X1 U269 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U270 ( .A1(data_in[4]), .A2(n839), .B1(n1099), .B2(\mem[11][4] ), 
        .ZN(n1095) );
  INV_X1 U271 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U272 ( .A1(data_in[5]), .A2(n839), .B1(n1099), .B2(\mem[11][5] ), 
        .ZN(n1094) );
  INV_X1 U273 ( .A(n1093), .ZN(n788) );
  AOI22_X1 U274 ( .A1(data_in[6]), .A2(n839), .B1(n1099), .B2(\mem[11][6] ), 
        .ZN(n1093) );
  INV_X1 U275 ( .A(n1092), .ZN(n787) );
  AOI22_X1 U276 ( .A1(data_in[7]), .A2(n839), .B1(n1099), .B2(\mem[11][7] ), 
        .ZN(n1092) );
  INV_X1 U277 ( .A(n1091), .ZN(n786) );
  AOI22_X1 U278 ( .A1(data_in[0]), .A2(n838), .B1(n1090), .B2(\mem[12][0] ), 
        .ZN(n1091) );
  INV_X1 U279 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U280 ( .A1(data_in[1]), .A2(n838), .B1(n1090), .B2(\mem[12][1] ), 
        .ZN(n1089) );
  INV_X1 U281 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U282 ( .A1(data_in[2]), .A2(n838), .B1(n1090), .B2(\mem[12][2] ), 
        .ZN(n1088) );
  INV_X1 U283 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U284 ( .A1(data_in[3]), .A2(n838), .B1(n1090), .B2(\mem[12][3] ), 
        .ZN(n1087) );
  INV_X1 U285 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U286 ( .A1(data_in[4]), .A2(n838), .B1(n1090), .B2(\mem[12][4] ), 
        .ZN(n1086) );
  INV_X1 U287 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U288 ( .A1(data_in[5]), .A2(n838), .B1(n1090), .B2(\mem[12][5] ), 
        .ZN(n1085) );
  INV_X1 U289 ( .A(n1084), .ZN(n780) );
  AOI22_X1 U290 ( .A1(data_in[6]), .A2(n838), .B1(n1090), .B2(\mem[12][6] ), 
        .ZN(n1084) );
  INV_X1 U291 ( .A(n1083), .ZN(n779) );
  AOI22_X1 U292 ( .A1(data_in[7]), .A2(n838), .B1(n1090), .B2(\mem[12][7] ), 
        .ZN(n1083) );
  INV_X1 U293 ( .A(n1082), .ZN(n778) );
  AOI22_X1 U294 ( .A1(data_in[0]), .A2(n837), .B1(n1081), .B2(\mem[13][0] ), 
        .ZN(n1082) );
  INV_X1 U295 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U296 ( .A1(data_in[1]), .A2(n837), .B1(n1081), .B2(\mem[13][1] ), 
        .ZN(n1080) );
  INV_X1 U297 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U298 ( .A1(data_in[2]), .A2(n837), .B1(n1081), .B2(\mem[13][2] ), 
        .ZN(n1079) );
  INV_X1 U299 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U300 ( .A1(data_in[3]), .A2(n837), .B1(n1081), .B2(\mem[13][3] ), 
        .ZN(n1078) );
  INV_X1 U301 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U302 ( .A1(data_in[4]), .A2(n837), .B1(n1081), .B2(\mem[13][4] ), 
        .ZN(n1077) );
  INV_X1 U303 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U304 ( .A1(data_in[5]), .A2(n837), .B1(n1081), .B2(\mem[13][5] ), 
        .ZN(n1076) );
  INV_X1 U305 ( .A(n1075), .ZN(n772) );
  AOI22_X1 U306 ( .A1(data_in[6]), .A2(n837), .B1(n1081), .B2(\mem[13][6] ), 
        .ZN(n1075) );
  INV_X1 U307 ( .A(n1074), .ZN(n771) );
  AOI22_X1 U308 ( .A1(data_in[7]), .A2(n837), .B1(n1081), .B2(\mem[13][7] ), 
        .ZN(n1074) );
  INV_X1 U309 ( .A(n1073), .ZN(n770) );
  AOI22_X1 U310 ( .A1(data_in[0]), .A2(n836), .B1(n1072), .B2(\mem[14][0] ), 
        .ZN(n1073) );
  INV_X1 U311 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U312 ( .A1(data_in[1]), .A2(n836), .B1(n1072), .B2(\mem[14][1] ), 
        .ZN(n1071) );
  INV_X1 U313 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U314 ( .A1(data_in[2]), .A2(n836), .B1(n1072), .B2(\mem[14][2] ), 
        .ZN(n1070) );
  INV_X1 U315 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U316 ( .A1(data_in[3]), .A2(n836), .B1(n1072), .B2(\mem[14][3] ), 
        .ZN(n1069) );
  INV_X1 U317 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U318 ( .A1(data_in[4]), .A2(n836), .B1(n1072), .B2(\mem[14][4] ), 
        .ZN(n1068) );
  INV_X1 U319 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U320 ( .A1(data_in[5]), .A2(n836), .B1(n1072), .B2(\mem[14][5] ), 
        .ZN(n1067) );
  INV_X1 U321 ( .A(n1066), .ZN(n764) );
  AOI22_X1 U322 ( .A1(data_in[6]), .A2(n836), .B1(n1072), .B2(\mem[14][6] ), 
        .ZN(n1066) );
  INV_X1 U323 ( .A(n1065), .ZN(n763) );
  AOI22_X1 U324 ( .A1(data_in[7]), .A2(n836), .B1(n1072), .B2(\mem[14][7] ), 
        .ZN(n1065) );
  INV_X1 U325 ( .A(n1064), .ZN(n762) );
  AOI22_X1 U326 ( .A1(data_in[0]), .A2(n835), .B1(n1063), .B2(\mem[15][0] ), 
        .ZN(n1064) );
  INV_X1 U327 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U328 ( .A1(data_in[1]), .A2(n835), .B1(n1063), .B2(\mem[15][1] ), 
        .ZN(n1062) );
  INV_X1 U329 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U330 ( .A1(data_in[2]), .A2(n835), .B1(n1063), .B2(\mem[15][2] ), 
        .ZN(n1061) );
  INV_X1 U331 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U332 ( .A1(data_in[3]), .A2(n835), .B1(n1063), .B2(\mem[15][3] ), 
        .ZN(n1060) );
  INV_X1 U333 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U334 ( .A1(data_in[4]), .A2(n835), .B1(n1063), .B2(\mem[15][4] ), 
        .ZN(n1059) );
  INV_X1 U335 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U336 ( .A1(data_in[5]), .A2(n835), .B1(n1063), .B2(\mem[15][5] ), 
        .ZN(n1058) );
  INV_X1 U337 ( .A(n1057), .ZN(n756) );
  AOI22_X1 U338 ( .A1(data_in[6]), .A2(n835), .B1(n1063), .B2(\mem[15][6] ), 
        .ZN(n1057) );
  INV_X1 U339 ( .A(n1056), .ZN(n755) );
  AOI22_X1 U340 ( .A1(data_in[7]), .A2(n835), .B1(n1063), .B2(\mem[15][7] ), 
        .ZN(n1056) );
  INV_X1 U341 ( .A(n1055), .ZN(n754) );
  AOI22_X1 U342 ( .A1(data_in[0]), .A2(n834), .B1(n1054), .B2(\mem[16][0] ), 
        .ZN(n1055) );
  INV_X1 U343 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U344 ( .A1(data_in[1]), .A2(n834), .B1(n1054), .B2(\mem[16][1] ), 
        .ZN(n1053) );
  INV_X1 U345 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U346 ( .A1(data_in[2]), .A2(n834), .B1(n1054), .B2(\mem[16][2] ), 
        .ZN(n1052) );
  INV_X1 U347 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U348 ( .A1(data_in[3]), .A2(n834), .B1(n1054), .B2(\mem[16][3] ), 
        .ZN(n1051) );
  INV_X1 U349 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U350 ( .A1(data_in[4]), .A2(n834), .B1(n1054), .B2(\mem[16][4] ), 
        .ZN(n1050) );
  INV_X1 U351 ( .A(n1049), .ZN(n749) );
  AOI22_X1 U352 ( .A1(data_in[5]), .A2(n834), .B1(n1054), .B2(\mem[16][5] ), 
        .ZN(n1049) );
  INV_X1 U353 ( .A(n1048), .ZN(n748) );
  AOI22_X1 U354 ( .A1(data_in[6]), .A2(n834), .B1(n1054), .B2(\mem[16][6] ), 
        .ZN(n1048) );
  INV_X1 U355 ( .A(n1047), .ZN(n747) );
  AOI22_X1 U356 ( .A1(data_in[7]), .A2(n834), .B1(n1054), .B2(\mem[16][7] ), 
        .ZN(n1047) );
  INV_X1 U357 ( .A(n1045), .ZN(n746) );
  AOI22_X1 U358 ( .A1(data_in[0]), .A2(n833), .B1(n1044), .B2(\mem[17][0] ), 
        .ZN(n1045) );
  INV_X1 U359 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U360 ( .A1(data_in[1]), .A2(n833), .B1(n1044), .B2(\mem[17][1] ), 
        .ZN(n1043) );
  INV_X1 U361 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U362 ( .A1(data_in[2]), .A2(n833), .B1(n1044), .B2(\mem[17][2] ), 
        .ZN(n1042) );
  INV_X1 U363 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U364 ( .A1(data_in[3]), .A2(n833), .B1(n1044), .B2(\mem[17][3] ), 
        .ZN(n1041) );
  INV_X1 U365 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U366 ( .A1(data_in[4]), .A2(n833), .B1(n1044), .B2(\mem[17][4] ), 
        .ZN(n1040) );
  INV_X1 U367 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U368 ( .A1(data_in[5]), .A2(n833), .B1(n1044), .B2(\mem[17][5] ), 
        .ZN(n1039) );
  INV_X1 U369 ( .A(n1038), .ZN(n740) );
  AOI22_X1 U370 ( .A1(data_in[6]), .A2(n833), .B1(n1044), .B2(\mem[17][6] ), 
        .ZN(n1038) );
  INV_X1 U371 ( .A(n1037), .ZN(n739) );
  AOI22_X1 U372 ( .A1(data_in[7]), .A2(n833), .B1(n1044), .B2(\mem[17][7] ), 
        .ZN(n1037) );
  INV_X1 U373 ( .A(n1036), .ZN(n738) );
  AOI22_X1 U374 ( .A1(data_in[0]), .A2(n832), .B1(n1035), .B2(\mem[18][0] ), 
        .ZN(n1036) );
  INV_X1 U375 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U376 ( .A1(data_in[1]), .A2(n832), .B1(n1035), .B2(\mem[18][1] ), 
        .ZN(n1034) );
  INV_X1 U377 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U378 ( .A1(data_in[2]), .A2(n832), .B1(n1035), .B2(\mem[18][2] ), 
        .ZN(n1033) );
  INV_X1 U379 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U380 ( .A1(data_in[3]), .A2(n832), .B1(n1035), .B2(\mem[18][3] ), 
        .ZN(n1032) );
  INV_X1 U381 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U382 ( .A1(data_in[4]), .A2(n832), .B1(n1035), .B2(\mem[18][4] ), 
        .ZN(n1031) );
  INV_X1 U383 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U384 ( .A1(data_in[5]), .A2(n832), .B1(n1035), .B2(\mem[18][5] ), 
        .ZN(n1030) );
  INV_X1 U385 ( .A(n1029), .ZN(n732) );
  AOI22_X1 U386 ( .A1(data_in[6]), .A2(n832), .B1(n1035), .B2(\mem[18][6] ), 
        .ZN(n1029) );
  INV_X1 U387 ( .A(n1028), .ZN(n731) );
  AOI22_X1 U388 ( .A1(data_in[7]), .A2(n832), .B1(n1035), .B2(\mem[18][7] ), 
        .ZN(n1028) );
  INV_X1 U389 ( .A(n1027), .ZN(n730) );
  AOI22_X1 U390 ( .A1(data_in[0]), .A2(n831), .B1(n1026), .B2(\mem[19][0] ), 
        .ZN(n1027) );
  INV_X1 U391 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U392 ( .A1(data_in[1]), .A2(n831), .B1(n1026), .B2(\mem[19][1] ), 
        .ZN(n1025) );
  INV_X1 U393 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U394 ( .A1(data_in[2]), .A2(n831), .B1(n1026), .B2(\mem[19][2] ), 
        .ZN(n1024) );
  INV_X1 U395 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U396 ( .A1(data_in[3]), .A2(n831), .B1(n1026), .B2(\mem[19][3] ), 
        .ZN(n1023) );
  INV_X1 U397 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U398 ( .A1(data_in[4]), .A2(n831), .B1(n1026), .B2(\mem[19][4] ), 
        .ZN(n1022) );
  INV_X1 U399 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U400 ( .A1(data_in[5]), .A2(n831), .B1(n1026), .B2(\mem[19][5] ), 
        .ZN(n1021) );
  INV_X1 U401 ( .A(n1020), .ZN(n724) );
  AOI22_X1 U402 ( .A1(data_in[6]), .A2(n831), .B1(n1026), .B2(\mem[19][6] ), 
        .ZN(n1020) );
  INV_X1 U403 ( .A(n1019), .ZN(n723) );
  AOI22_X1 U404 ( .A1(data_in[7]), .A2(n831), .B1(n1026), .B2(\mem[19][7] ), 
        .ZN(n1019) );
  INV_X1 U405 ( .A(n1018), .ZN(n722) );
  AOI22_X1 U406 ( .A1(data_in[0]), .A2(n830), .B1(n1017), .B2(\mem[20][0] ), 
        .ZN(n1018) );
  INV_X1 U407 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U408 ( .A1(data_in[1]), .A2(n830), .B1(n1017), .B2(\mem[20][1] ), 
        .ZN(n1016) );
  INV_X1 U409 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U410 ( .A1(data_in[2]), .A2(n830), .B1(n1017), .B2(\mem[20][2] ), 
        .ZN(n1015) );
  INV_X1 U411 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U412 ( .A1(data_in[3]), .A2(n830), .B1(n1017), .B2(\mem[20][3] ), 
        .ZN(n1014) );
  INV_X1 U413 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U414 ( .A1(data_in[4]), .A2(n830), .B1(n1017), .B2(\mem[20][4] ), 
        .ZN(n1013) );
  INV_X1 U415 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U416 ( .A1(data_in[5]), .A2(n830), .B1(n1017), .B2(\mem[20][5] ), 
        .ZN(n1012) );
  INV_X1 U417 ( .A(n1011), .ZN(n716) );
  AOI22_X1 U418 ( .A1(data_in[6]), .A2(n830), .B1(n1017), .B2(\mem[20][6] ), 
        .ZN(n1011) );
  INV_X1 U419 ( .A(n1010), .ZN(n715) );
  AOI22_X1 U420 ( .A1(data_in[7]), .A2(n830), .B1(n1017), .B2(\mem[20][7] ), 
        .ZN(n1010) );
  INV_X1 U421 ( .A(n1009), .ZN(n714) );
  AOI22_X1 U422 ( .A1(data_in[0]), .A2(n829), .B1(n1008), .B2(\mem[21][0] ), 
        .ZN(n1009) );
  INV_X1 U423 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U424 ( .A1(data_in[1]), .A2(n829), .B1(n1008), .B2(\mem[21][1] ), 
        .ZN(n1007) );
  INV_X1 U425 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U426 ( .A1(data_in[2]), .A2(n829), .B1(n1008), .B2(\mem[21][2] ), 
        .ZN(n1006) );
  INV_X1 U427 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U428 ( .A1(data_in[3]), .A2(n829), .B1(n1008), .B2(\mem[21][3] ), 
        .ZN(n1005) );
  INV_X1 U429 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U430 ( .A1(data_in[4]), .A2(n829), .B1(n1008), .B2(\mem[21][4] ), 
        .ZN(n1004) );
  INV_X1 U431 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U432 ( .A1(data_in[5]), .A2(n829), .B1(n1008), .B2(\mem[21][5] ), 
        .ZN(n1003) );
  INV_X1 U433 ( .A(n1002), .ZN(n708) );
  AOI22_X1 U434 ( .A1(data_in[6]), .A2(n829), .B1(n1008), .B2(\mem[21][6] ), 
        .ZN(n1002) );
  INV_X1 U435 ( .A(n1001), .ZN(n707) );
  AOI22_X1 U436 ( .A1(data_in[7]), .A2(n829), .B1(n1008), .B2(\mem[21][7] ), 
        .ZN(n1001) );
  INV_X1 U437 ( .A(n1000), .ZN(n706) );
  AOI22_X1 U438 ( .A1(data_in[0]), .A2(n828), .B1(n999), .B2(\mem[22][0] ), 
        .ZN(n1000) );
  INV_X1 U439 ( .A(n998), .ZN(n705) );
  AOI22_X1 U440 ( .A1(data_in[1]), .A2(n828), .B1(n999), .B2(\mem[22][1] ), 
        .ZN(n998) );
  INV_X1 U441 ( .A(n997), .ZN(n704) );
  AOI22_X1 U442 ( .A1(data_in[2]), .A2(n828), .B1(n999), .B2(\mem[22][2] ), 
        .ZN(n997) );
  INV_X1 U443 ( .A(n996), .ZN(n703) );
  AOI22_X1 U444 ( .A1(data_in[3]), .A2(n828), .B1(n999), .B2(\mem[22][3] ), 
        .ZN(n996) );
  INV_X1 U445 ( .A(n995), .ZN(n702) );
  AOI22_X1 U446 ( .A1(data_in[4]), .A2(n828), .B1(n999), .B2(\mem[22][4] ), 
        .ZN(n995) );
  INV_X1 U447 ( .A(n994), .ZN(n701) );
  AOI22_X1 U448 ( .A1(data_in[5]), .A2(n828), .B1(n999), .B2(\mem[22][5] ), 
        .ZN(n994) );
  INV_X1 U449 ( .A(n993), .ZN(n700) );
  AOI22_X1 U450 ( .A1(data_in[6]), .A2(n828), .B1(n999), .B2(\mem[22][6] ), 
        .ZN(n993) );
  INV_X1 U451 ( .A(n992), .ZN(n699) );
  AOI22_X1 U452 ( .A1(data_in[7]), .A2(n828), .B1(n999), .B2(\mem[22][7] ), 
        .ZN(n992) );
  INV_X1 U453 ( .A(n991), .ZN(n698) );
  AOI22_X1 U454 ( .A1(data_in[0]), .A2(n827), .B1(n990), .B2(\mem[23][0] ), 
        .ZN(n991) );
  INV_X1 U455 ( .A(n989), .ZN(n697) );
  AOI22_X1 U456 ( .A1(data_in[1]), .A2(n827), .B1(n990), .B2(\mem[23][1] ), 
        .ZN(n989) );
  INV_X1 U457 ( .A(n988), .ZN(n696) );
  AOI22_X1 U458 ( .A1(data_in[2]), .A2(n827), .B1(n990), .B2(\mem[23][2] ), 
        .ZN(n988) );
  INV_X1 U459 ( .A(n987), .ZN(n695) );
  AOI22_X1 U460 ( .A1(data_in[3]), .A2(n827), .B1(n990), .B2(\mem[23][3] ), 
        .ZN(n987) );
  INV_X1 U461 ( .A(n986), .ZN(n694) );
  AOI22_X1 U462 ( .A1(data_in[4]), .A2(n827), .B1(n990), .B2(\mem[23][4] ), 
        .ZN(n986) );
  INV_X1 U463 ( .A(n985), .ZN(n693) );
  AOI22_X1 U464 ( .A1(data_in[5]), .A2(n827), .B1(n990), .B2(\mem[23][5] ), 
        .ZN(n985) );
  INV_X1 U465 ( .A(n984), .ZN(n692) );
  AOI22_X1 U466 ( .A1(data_in[6]), .A2(n827), .B1(n990), .B2(\mem[23][6] ), 
        .ZN(n984) );
  INV_X1 U467 ( .A(n983), .ZN(n691) );
  AOI22_X1 U468 ( .A1(data_in[7]), .A2(n827), .B1(n990), .B2(\mem[23][7] ), 
        .ZN(n983) );
  INV_X1 U469 ( .A(n982), .ZN(n690) );
  AOI22_X1 U470 ( .A1(data_in[0]), .A2(n826), .B1(n981), .B2(\mem[24][0] ), 
        .ZN(n982) );
  INV_X1 U471 ( .A(n980), .ZN(n689) );
  AOI22_X1 U472 ( .A1(data_in[1]), .A2(n826), .B1(n981), .B2(\mem[24][1] ), 
        .ZN(n980) );
  INV_X1 U473 ( .A(n979), .ZN(n688) );
  AOI22_X1 U474 ( .A1(data_in[2]), .A2(n826), .B1(n981), .B2(\mem[24][2] ), 
        .ZN(n979) );
  INV_X1 U475 ( .A(n978), .ZN(n687) );
  AOI22_X1 U476 ( .A1(data_in[3]), .A2(n826), .B1(n981), .B2(\mem[24][3] ), 
        .ZN(n978) );
  INV_X1 U477 ( .A(n977), .ZN(n686) );
  AOI22_X1 U478 ( .A1(data_in[4]), .A2(n826), .B1(n981), .B2(\mem[24][4] ), 
        .ZN(n977) );
  INV_X1 U479 ( .A(n976), .ZN(n685) );
  AOI22_X1 U480 ( .A1(data_in[5]), .A2(n826), .B1(n981), .B2(\mem[24][5] ), 
        .ZN(n976) );
  INV_X1 U481 ( .A(n975), .ZN(n684) );
  AOI22_X1 U482 ( .A1(data_in[6]), .A2(n826), .B1(n981), .B2(\mem[24][6] ), 
        .ZN(n975) );
  INV_X1 U483 ( .A(n974), .ZN(n683) );
  AOI22_X1 U484 ( .A1(data_in[7]), .A2(n826), .B1(n981), .B2(\mem[24][7] ), 
        .ZN(n974) );
  INV_X1 U485 ( .A(n972), .ZN(n682) );
  AOI22_X1 U486 ( .A1(data_in[0]), .A2(n825), .B1(n971), .B2(\mem[25][0] ), 
        .ZN(n972) );
  INV_X1 U487 ( .A(n970), .ZN(n681) );
  AOI22_X1 U488 ( .A1(data_in[1]), .A2(n825), .B1(n971), .B2(\mem[25][1] ), 
        .ZN(n970) );
  INV_X1 U489 ( .A(n969), .ZN(n680) );
  AOI22_X1 U490 ( .A1(data_in[2]), .A2(n825), .B1(n971), .B2(\mem[25][2] ), 
        .ZN(n969) );
  INV_X1 U491 ( .A(n968), .ZN(n679) );
  AOI22_X1 U492 ( .A1(data_in[3]), .A2(n825), .B1(n971), .B2(\mem[25][3] ), 
        .ZN(n968) );
  INV_X1 U493 ( .A(n967), .ZN(n678) );
  AOI22_X1 U494 ( .A1(data_in[4]), .A2(n825), .B1(n971), .B2(\mem[25][4] ), 
        .ZN(n967) );
  INV_X1 U495 ( .A(n966), .ZN(n677) );
  AOI22_X1 U496 ( .A1(data_in[5]), .A2(n825), .B1(n971), .B2(\mem[25][5] ), 
        .ZN(n966) );
  INV_X1 U497 ( .A(n965), .ZN(n676) );
  AOI22_X1 U498 ( .A1(data_in[6]), .A2(n825), .B1(n971), .B2(\mem[25][6] ), 
        .ZN(n965) );
  INV_X1 U499 ( .A(n964), .ZN(n675) );
  AOI22_X1 U500 ( .A1(data_in[7]), .A2(n825), .B1(n971), .B2(\mem[25][7] ), 
        .ZN(n964) );
  INV_X1 U501 ( .A(n963), .ZN(n674) );
  AOI22_X1 U502 ( .A1(data_in[0]), .A2(n824), .B1(n962), .B2(\mem[26][0] ), 
        .ZN(n963) );
  INV_X1 U503 ( .A(n961), .ZN(n673) );
  AOI22_X1 U504 ( .A1(data_in[1]), .A2(n824), .B1(n962), .B2(\mem[26][1] ), 
        .ZN(n961) );
  INV_X1 U505 ( .A(n960), .ZN(n672) );
  AOI22_X1 U506 ( .A1(data_in[2]), .A2(n824), .B1(n962), .B2(\mem[26][2] ), 
        .ZN(n960) );
  INV_X1 U507 ( .A(n959), .ZN(n671) );
  AOI22_X1 U508 ( .A1(data_in[3]), .A2(n824), .B1(n962), .B2(\mem[26][3] ), 
        .ZN(n959) );
  INV_X1 U509 ( .A(n958), .ZN(n670) );
  AOI22_X1 U510 ( .A1(data_in[4]), .A2(n824), .B1(n962), .B2(\mem[26][4] ), 
        .ZN(n958) );
  INV_X1 U511 ( .A(n957), .ZN(n669) );
  AOI22_X1 U512 ( .A1(data_in[5]), .A2(n824), .B1(n962), .B2(\mem[26][5] ), 
        .ZN(n957) );
  INV_X1 U513 ( .A(n956), .ZN(n668) );
  AOI22_X1 U514 ( .A1(data_in[6]), .A2(n824), .B1(n962), .B2(\mem[26][6] ), 
        .ZN(n956) );
  INV_X1 U515 ( .A(n955), .ZN(n667) );
  AOI22_X1 U516 ( .A1(data_in[7]), .A2(n824), .B1(n962), .B2(\mem[26][7] ), 
        .ZN(n955) );
  INV_X1 U517 ( .A(n954), .ZN(n666) );
  AOI22_X1 U518 ( .A1(data_in[0]), .A2(n823), .B1(n953), .B2(\mem[27][0] ), 
        .ZN(n954) );
  INV_X1 U519 ( .A(n952), .ZN(n665) );
  AOI22_X1 U520 ( .A1(data_in[1]), .A2(n823), .B1(n953), .B2(\mem[27][1] ), 
        .ZN(n952) );
  INV_X1 U521 ( .A(n951), .ZN(n664) );
  AOI22_X1 U522 ( .A1(data_in[2]), .A2(n823), .B1(n953), .B2(\mem[27][2] ), 
        .ZN(n951) );
  INV_X1 U523 ( .A(n950), .ZN(n663) );
  AOI22_X1 U524 ( .A1(data_in[3]), .A2(n823), .B1(n953), .B2(\mem[27][3] ), 
        .ZN(n950) );
  INV_X1 U525 ( .A(n949), .ZN(n662) );
  AOI22_X1 U526 ( .A1(data_in[4]), .A2(n823), .B1(n953), .B2(\mem[27][4] ), 
        .ZN(n949) );
  INV_X1 U527 ( .A(n948), .ZN(n661) );
  AOI22_X1 U528 ( .A1(data_in[5]), .A2(n823), .B1(n953), .B2(\mem[27][5] ), 
        .ZN(n948) );
  INV_X1 U529 ( .A(n947), .ZN(n660) );
  AOI22_X1 U530 ( .A1(data_in[6]), .A2(n823), .B1(n953), .B2(\mem[27][6] ), 
        .ZN(n947) );
  INV_X1 U531 ( .A(n946), .ZN(n659) );
  AOI22_X1 U532 ( .A1(data_in[7]), .A2(n823), .B1(n953), .B2(\mem[27][7] ), 
        .ZN(n946) );
  INV_X1 U533 ( .A(n945), .ZN(n658) );
  AOI22_X1 U534 ( .A1(data_in[0]), .A2(n822), .B1(n944), .B2(\mem[28][0] ), 
        .ZN(n945) );
  INV_X1 U535 ( .A(n943), .ZN(n657) );
  AOI22_X1 U536 ( .A1(data_in[1]), .A2(n822), .B1(n944), .B2(\mem[28][1] ), 
        .ZN(n943) );
  INV_X1 U537 ( .A(n942), .ZN(n656) );
  AOI22_X1 U538 ( .A1(data_in[2]), .A2(n822), .B1(n944), .B2(\mem[28][2] ), 
        .ZN(n942) );
  INV_X1 U539 ( .A(n941), .ZN(n655) );
  AOI22_X1 U540 ( .A1(data_in[3]), .A2(n822), .B1(n944), .B2(\mem[28][3] ), 
        .ZN(n941) );
  INV_X1 U541 ( .A(n940), .ZN(n654) );
  AOI22_X1 U542 ( .A1(data_in[4]), .A2(n822), .B1(n944), .B2(\mem[28][4] ), 
        .ZN(n940) );
  INV_X1 U543 ( .A(n939), .ZN(n653) );
  AOI22_X1 U544 ( .A1(data_in[5]), .A2(n822), .B1(n944), .B2(\mem[28][5] ), 
        .ZN(n939) );
  INV_X1 U545 ( .A(n938), .ZN(n652) );
  AOI22_X1 U546 ( .A1(data_in[6]), .A2(n822), .B1(n944), .B2(\mem[28][6] ), 
        .ZN(n938) );
  INV_X1 U547 ( .A(n937), .ZN(n651) );
  AOI22_X1 U548 ( .A1(data_in[7]), .A2(n822), .B1(n944), .B2(\mem[28][7] ), 
        .ZN(n937) );
  INV_X1 U549 ( .A(n936), .ZN(n650) );
  AOI22_X1 U550 ( .A1(data_in[0]), .A2(n821), .B1(n935), .B2(\mem[29][0] ), 
        .ZN(n936) );
  INV_X1 U551 ( .A(n934), .ZN(n649) );
  AOI22_X1 U552 ( .A1(data_in[1]), .A2(n821), .B1(n935), .B2(\mem[29][1] ), 
        .ZN(n934) );
  INV_X1 U553 ( .A(n933), .ZN(n648) );
  AOI22_X1 U554 ( .A1(data_in[2]), .A2(n821), .B1(n935), .B2(\mem[29][2] ), 
        .ZN(n933) );
  INV_X1 U555 ( .A(n932), .ZN(n647) );
  AOI22_X1 U556 ( .A1(data_in[3]), .A2(n821), .B1(n935), .B2(\mem[29][3] ), 
        .ZN(n932) );
  INV_X1 U557 ( .A(n931), .ZN(n646) );
  AOI22_X1 U558 ( .A1(data_in[4]), .A2(n821), .B1(n935), .B2(\mem[29][4] ), 
        .ZN(n931) );
  INV_X1 U559 ( .A(n930), .ZN(n645) );
  AOI22_X1 U560 ( .A1(data_in[5]), .A2(n821), .B1(n935), .B2(\mem[29][5] ), 
        .ZN(n930) );
  INV_X1 U561 ( .A(n929), .ZN(n644) );
  AOI22_X1 U562 ( .A1(data_in[6]), .A2(n821), .B1(n935), .B2(\mem[29][6] ), 
        .ZN(n929) );
  INV_X1 U563 ( .A(n928), .ZN(n643) );
  AOI22_X1 U564 ( .A1(data_in[7]), .A2(n821), .B1(n935), .B2(\mem[29][7] ), 
        .ZN(n928) );
  INV_X1 U565 ( .A(n927), .ZN(n642) );
  AOI22_X1 U566 ( .A1(data_in[0]), .A2(n820), .B1(n926), .B2(\mem[30][0] ), 
        .ZN(n927) );
  INV_X1 U567 ( .A(n925), .ZN(n641) );
  AOI22_X1 U568 ( .A1(data_in[1]), .A2(n820), .B1(n926), .B2(\mem[30][1] ), 
        .ZN(n925) );
  INV_X1 U569 ( .A(n924), .ZN(n640) );
  AOI22_X1 U570 ( .A1(data_in[2]), .A2(n820), .B1(n926), .B2(\mem[30][2] ), 
        .ZN(n924) );
  INV_X1 U571 ( .A(n923), .ZN(n639) );
  AOI22_X1 U572 ( .A1(data_in[3]), .A2(n820), .B1(n926), .B2(\mem[30][3] ), 
        .ZN(n923) );
  INV_X1 U573 ( .A(n922), .ZN(n638) );
  AOI22_X1 U574 ( .A1(data_in[4]), .A2(n820), .B1(n926), .B2(\mem[30][4] ), 
        .ZN(n922) );
  INV_X1 U575 ( .A(n921), .ZN(n637) );
  AOI22_X1 U576 ( .A1(data_in[5]), .A2(n820), .B1(n926), .B2(\mem[30][5] ), 
        .ZN(n921) );
  INV_X1 U577 ( .A(n920), .ZN(n636) );
  AOI22_X1 U578 ( .A1(data_in[6]), .A2(n820), .B1(n926), .B2(\mem[30][6] ), 
        .ZN(n920) );
  INV_X1 U579 ( .A(n919), .ZN(n635) );
  AOI22_X1 U580 ( .A1(data_in[7]), .A2(n820), .B1(n926), .B2(\mem[30][7] ), 
        .ZN(n919) );
  INV_X1 U581 ( .A(n918), .ZN(n634) );
  AOI22_X1 U582 ( .A1(data_in[0]), .A2(n819), .B1(n917), .B2(\mem[31][0] ), 
        .ZN(n918) );
  INV_X1 U583 ( .A(n916), .ZN(n633) );
  AOI22_X1 U584 ( .A1(data_in[1]), .A2(n819), .B1(n917), .B2(\mem[31][1] ), 
        .ZN(n916) );
  INV_X1 U585 ( .A(n915), .ZN(n632) );
  AOI22_X1 U586 ( .A1(data_in[2]), .A2(n819), .B1(n917), .B2(\mem[31][2] ), 
        .ZN(n915) );
  INV_X1 U587 ( .A(n914), .ZN(n631) );
  AOI22_X1 U588 ( .A1(data_in[3]), .A2(n819), .B1(n917), .B2(\mem[31][3] ), 
        .ZN(n914) );
  INV_X1 U589 ( .A(n913), .ZN(n630) );
  AOI22_X1 U590 ( .A1(data_in[4]), .A2(n819), .B1(n917), .B2(\mem[31][4] ), 
        .ZN(n913) );
  INV_X1 U591 ( .A(n912), .ZN(n629) );
  AOI22_X1 U592 ( .A1(data_in[5]), .A2(n819), .B1(n917), .B2(\mem[31][5] ), 
        .ZN(n912) );
  INV_X1 U593 ( .A(n911), .ZN(n628) );
  AOI22_X1 U594 ( .A1(data_in[6]), .A2(n819), .B1(n917), .B2(\mem[31][6] ), 
        .ZN(n911) );
  INV_X1 U595 ( .A(n910), .ZN(n627) );
  AOI22_X1 U596 ( .A1(data_in[7]), .A2(n819), .B1(n917), .B2(\mem[31][7] ), 
        .ZN(n910) );
  MUX2_X1 U597 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n611), .Z(n1) );
  MUX2_X1 U598 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n611), .Z(n2) );
  MUX2_X1 U599 ( .A(n2), .B(n1), .S(n608), .Z(n3) );
  MUX2_X1 U600 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n611), .Z(n4) );
  MUX2_X1 U601 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n611), .Z(n5) );
  MUX2_X1 U602 ( .A(n5), .B(n4), .S(n608), .Z(n6) );
  MUX2_X1 U603 ( .A(n6), .B(n3), .S(n607), .Z(n7) );
  MUX2_X1 U604 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n611), .Z(n8) );
  MUX2_X1 U605 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n611), .Z(n9) );
  MUX2_X1 U606 ( .A(n9), .B(n8), .S(n608), .Z(n10) );
  MUX2_X1 U607 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n611), .Z(n11) );
  MUX2_X1 U608 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n611), .Z(n12) );
  MUX2_X1 U609 ( .A(n12), .B(n11), .S(n608), .Z(n13) );
  MUX2_X1 U610 ( .A(n13), .B(n10), .S(N12), .Z(n14) );
  MUX2_X1 U611 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U612 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n611), .Z(n16) );
  MUX2_X1 U613 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n614), .Z(n17) );
  MUX2_X1 U614 ( .A(n17), .B(n16), .S(n609), .Z(n18) );
  MUX2_X1 U615 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n613), .Z(n19) );
  MUX2_X1 U616 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n611), .Z(n20) );
  MUX2_X1 U617 ( .A(n20), .B(n19), .S(n609), .Z(n21) );
  MUX2_X1 U618 ( .A(n21), .B(n18), .S(N12), .Z(n22) );
  MUX2_X1 U619 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n612), .Z(n23) );
  MUX2_X1 U620 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n615), .Z(n24) );
  MUX2_X1 U621 ( .A(n24), .B(n23), .S(n609), .Z(n25) );
  MUX2_X1 U622 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n616), .Z(n26) );
  MUX2_X1 U623 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n616), .Z(n27) );
  MUX2_X1 U624 ( .A(n27), .B(n26), .S(n609), .Z(n28) );
  MUX2_X1 U625 ( .A(n28), .B(n25), .S(n606), .Z(n29) );
  MUX2_X1 U626 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U627 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U628 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n611), .Z(n31) );
  MUX2_X1 U629 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n611), .Z(n32) );
  MUX2_X1 U630 ( .A(n32), .B(n31), .S(n609), .Z(n33) );
  MUX2_X1 U631 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n611), .Z(n34) );
  MUX2_X1 U632 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n616), .Z(n35) );
  MUX2_X1 U633 ( .A(n35), .B(n34), .S(n609), .Z(n36) );
  MUX2_X1 U634 ( .A(n36), .B(n33), .S(n606), .Z(n37) );
  MUX2_X1 U635 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n613), .Z(n38) );
  MUX2_X1 U636 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n616), .Z(n39) );
  MUX2_X1 U637 ( .A(n39), .B(n38), .S(n609), .Z(n40) );
  MUX2_X1 U638 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n613), .Z(n41) );
  MUX2_X1 U639 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(N10), .Z(n42) );
  MUX2_X1 U640 ( .A(n42), .B(n41), .S(n609), .Z(n43) );
  MUX2_X1 U641 ( .A(n43), .B(n40), .S(N12), .Z(n44) );
  MUX2_X1 U642 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U643 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n612), .Z(n46) );
  MUX2_X1 U644 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n614), .Z(n47) );
  MUX2_X1 U645 ( .A(n47), .B(n46), .S(n609), .Z(n48) );
  MUX2_X1 U646 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n613), .Z(n49) );
  MUX2_X1 U647 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n616), .Z(n50) );
  MUX2_X1 U648 ( .A(n50), .B(n49), .S(n609), .Z(n51) );
  MUX2_X1 U649 ( .A(n51), .B(n48), .S(n607), .Z(n52) );
  MUX2_X1 U650 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n615), .Z(n53) );
  MUX2_X1 U651 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n54) );
  MUX2_X1 U652 ( .A(n54), .B(n53), .S(n609), .Z(n55) );
  MUX2_X1 U653 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n615), .Z(n56) );
  MUX2_X1 U654 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(N10), .Z(n57) );
  MUX2_X1 U655 ( .A(n57), .B(n56), .S(n609), .Z(n58) );
  MUX2_X1 U656 ( .A(n58), .B(n55), .S(n607), .Z(n59) );
  MUX2_X1 U657 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U658 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U659 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n612), .Z(n61) );
  MUX2_X1 U660 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n612), .Z(n62) );
  MUX2_X1 U661 ( .A(n62), .B(n61), .S(n610), .Z(n63) );
  MUX2_X1 U662 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n612), .Z(n64) );
  MUX2_X1 U663 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n612), .Z(n65) );
  MUX2_X1 U664 ( .A(n65), .B(n64), .S(n610), .Z(n66) );
  MUX2_X1 U665 ( .A(n66), .B(n63), .S(n606), .Z(n67) );
  MUX2_X1 U666 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n612), .Z(n68) );
  MUX2_X1 U667 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n612), .Z(n69) );
  MUX2_X1 U668 ( .A(n69), .B(n68), .S(n610), .Z(n70) );
  MUX2_X1 U669 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n612), .Z(n71) );
  MUX2_X1 U670 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n612), .Z(n72) );
  MUX2_X1 U671 ( .A(n72), .B(n71), .S(n610), .Z(n73) );
  MUX2_X1 U672 ( .A(n73), .B(n70), .S(n606), .Z(n74) );
  MUX2_X1 U673 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U674 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n612), .Z(n76) );
  MUX2_X1 U675 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n612), .Z(n77) );
  MUX2_X1 U676 ( .A(n77), .B(n76), .S(n610), .Z(n78) );
  MUX2_X1 U677 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n612), .Z(n79) );
  MUX2_X1 U678 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n612), .Z(n80) );
  MUX2_X1 U679 ( .A(n80), .B(n79), .S(n610), .Z(n81) );
  MUX2_X1 U680 ( .A(n81), .B(n78), .S(n606), .Z(n82) );
  MUX2_X1 U681 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n613), .Z(n83) );
  MUX2_X1 U682 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n613), .Z(n84) );
  MUX2_X1 U683 ( .A(n84), .B(n83), .S(n610), .Z(n85) );
  MUX2_X1 U684 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n613), .Z(n86) );
  MUX2_X1 U685 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n613), .Z(n87) );
  MUX2_X1 U686 ( .A(n87), .B(n86), .S(n610), .Z(n88) );
  MUX2_X1 U687 ( .A(n88), .B(n85), .S(n606), .Z(n89) );
  MUX2_X1 U688 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U689 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U690 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n613), .Z(n91) );
  MUX2_X1 U691 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n613), .Z(n92) );
  MUX2_X1 U692 ( .A(n92), .B(n91), .S(n610), .Z(n93) );
  MUX2_X1 U693 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n613), .Z(n94) );
  MUX2_X1 U694 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n613), .Z(n95) );
  MUX2_X1 U695 ( .A(n95), .B(n94), .S(n610), .Z(n96) );
  MUX2_X1 U696 ( .A(n96), .B(n93), .S(n606), .Z(n97) );
  MUX2_X1 U697 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n613), .Z(n98) );
  MUX2_X1 U698 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n613), .Z(n99) );
  MUX2_X1 U699 ( .A(n99), .B(n98), .S(n610), .Z(n100) );
  MUX2_X1 U700 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n613), .Z(n101) );
  MUX2_X1 U701 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n613), .Z(n102) );
  MUX2_X1 U702 ( .A(n102), .B(n101), .S(n610), .Z(n103) );
  MUX2_X1 U703 ( .A(n103), .B(n100), .S(n606), .Z(n104) );
  MUX2_X1 U704 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U705 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n616), .Z(n106) );
  MUX2_X1 U706 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n616), .Z(n107) );
  MUX2_X1 U707 ( .A(n107), .B(n106), .S(n610), .Z(n108) );
  MUX2_X1 U708 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n616), .Z(n109) );
  MUX2_X1 U709 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n616), .Z(n110) );
  MUX2_X1 U710 ( .A(n110), .B(n109), .S(n609), .Z(n111) );
  MUX2_X1 U711 ( .A(n111), .B(n108), .S(n606), .Z(n112) );
  MUX2_X1 U712 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n616), .Z(n113) );
  MUX2_X1 U713 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n616), .Z(n114) );
  MUX2_X1 U714 ( .A(n114), .B(n113), .S(n608), .Z(n115) );
  MUX2_X1 U715 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n616), .Z(n116) );
  MUX2_X1 U716 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n616), .Z(n117) );
  MUX2_X1 U717 ( .A(n117), .B(n116), .S(n610), .Z(n118) );
  MUX2_X1 U718 ( .A(n118), .B(n115), .S(n606), .Z(n119) );
  MUX2_X1 U719 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U720 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U721 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n616), .Z(n121) );
  MUX2_X1 U722 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n614), .Z(n122) );
  MUX2_X1 U723 ( .A(n122), .B(n121), .S(n608), .Z(n123) );
  MUX2_X1 U724 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n611), .Z(n124) );
  MUX2_X1 U725 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n615), .Z(n125) );
  MUX2_X1 U726 ( .A(n125), .B(n124), .S(n608), .Z(n126) );
  MUX2_X1 U727 ( .A(n126), .B(n123), .S(n606), .Z(n127) );
  MUX2_X1 U728 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n615), .Z(n128) );
  MUX2_X1 U729 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n616), .Z(n129) );
  MUX2_X1 U730 ( .A(n129), .B(n128), .S(n610), .Z(n130) );
  MUX2_X1 U731 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n616), .Z(n131) );
  MUX2_X1 U732 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n616), .Z(n132) );
  MUX2_X1 U733 ( .A(n132), .B(n131), .S(n609), .Z(n133) );
  MUX2_X1 U734 ( .A(n133), .B(n130), .S(n606), .Z(n134) );
  MUX2_X1 U735 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U736 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n611), .Z(n136) );
  MUX2_X1 U737 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n616), .Z(n137) );
  MUX2_X1 U738 ( .A(n137), .B(n136), .S(n609), .Z(n138) );
  MUX2_X1 U739 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n611), .Z(n139) );
  MUX2_X1 U740 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n614), .Z(n140) );
  MUX2_X1 U741 ( .A(n140), .B(n139), .S(n608), .Z(n141) );
  MUX2_X1 U742 ( .A(n141), .B(n138), .S(n606), .Z(n142) );
  MUX2_X1 U743 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(N10), .Z(n143) );
  MUX2_X1 U744 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n616), .Z(n144) );
  MUX2_X1 U745 ( .A(n144), .B(n143), .S(n609), .Z(n145) );
  MUX2_X1 U746 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n616), .Z(n146) );
  MUX2_X1 U747 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n611), .Z(n147) );
  MUX2_X1 U748 ( .A(n147), .B(n146), .S(n608), .Z(n148) );
  MUX2_X1 U749 ( .A(n148), .B(n145), .S(n606), .Z(n149) );
  MUX2_X1 U750 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U751 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U752 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n612), .Z(n151) );
  MUX2_X1 U753 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n612), .Z(n152) );
  MUX2_X1 U754 ( .A(n152), .B(n151), .S(N11), .Z(n153) );
  MUX2_X1 U755 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n612), .Z(n154) );
  MUX2_X1 U756 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n613), .Z(n155) );
  MUX2_X1 U757 ( .A(n155), .B(n154), .S(n609), .Z(n156) );
  MUX2_X1 U758 ( .A(n156), .B(n153), .S(n607), .Z(n157) );
  MUX2_X1 U759 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n612), .Z(n158) );
  MUX2_X1 U760 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n612), .Z(n159) );
  MUX2_X1 U761 ( .A(n159), .B(n158), .S(N11), .Z(n160) );
  MUX2_X1 U762 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n612), .Z(n161) );
  MUX2_X1 U763 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(N10), .Z(n162) );
  MUX2_X1 U764 ( .A(n162), .B(n161), .S(n609), .Z(n163) );
  MUX2_X1 U765 ( .A(n163), .B(n160), .S(n607), .Z(n164) );
  MUX2_X1 U766 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U767 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n612), .Z(n166) );
  MUX2_X1 U768 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n612), .Z(n167) );
  MUX2_X1 U769 ( .A(n167), .B(n166), .S(n608), .Z(n168) );
  MUX2_X1 U770 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n612), .Z(n169) );
  MUX2_X1 U771 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n611), .Z(n170) );
  MUX2_X1 U772 ( .A(n170), .B(n169), .S(N11), .Z(n171) );
  MUX2_X1 U773 ( .A(n171), .B(n168), .S(n607), .Z(n172) );
  MUX2_X1 U774 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n614), .Z(n173) );
  MUX2_X1 U775 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n614), .Z(n174) );
  MUX2_X1 U776 ( .A(n174), .B(n173), .S(n610), .Z(n175) );
  MUX2_X1 U777 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n614), .Z(n176) );
  MUX2_X1 U778 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n614), .Z(n177) );
  MUX2_X1 U779 ( .A(n177), .B(n176), .S(n609), .Z(n178) );
  MUX2_X1 U780 ( .A(n178), .B(n175), .S(n607), .Z(n179) );
  MUX2_X1 U781 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U782 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U783 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n614), .Z(n181) );
  MUX2_X1 U784 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n614), .Z(n182) );
  MUX2_X1 U785 ( .A(n182), .B(n181), .S(n609), .Z(n183) );
  MUX2_X1 U786 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n614), .Z(n184) );
  MUX2_X1 U787 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n614), .Z(n185) );
  MUX2_X1 U788 ( .A(n185), .B(n184), .S(N11), .Z(n186) );
  MUX2_X1 U789 ( .A(n186), .B(n183), .S(n607), .Z(n187) );
  MUX2_X1 U790 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n614), .Z(n188) );
  MUX2_X1 U791 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n614), .Z(n189) );
  MUX2_X1 U792 ( .A(n189), .B(n188), .S(n610), .Z(n190) );
  MUX2_X1 U793 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n614), .Z(n191) );
  MUX2_X1 U794 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n614), .Z(n192) );
  MUX2_X1 U795 ( .A(n192), .B(n191), .S(N11), .Z(n193) );
  MUX2_X1 U796 ( .A(n193), .B(n190), .S(n607), .Z(n194) );
  MUX2_X1 U797 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U798 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n615), .Z(n196) );
  MUX2_X1 U799 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n615), .Z(n197) );
  MUX2_X1 U800 ( .A(n197), .B(n196), .S(n608), .Z(n198) );
  MUX2_X1 U801 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n615), .Z(n199) );
  MUX2_X1 U802 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n615), .Z(n200) );
  MUX2_X1 U803 ( .A(n200), .B(n199), .S(n609), .Z(n201) );
  MUX2_X1 U804 ( .A(n201), .B(n198), .S(n607), .Z(n202) );
  MUX2_X1 U805 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n615), .Z(n203) );
  MUX2_X1 U806 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n615), .Z(n204) );
  MUX2_X1 U807 ( .A(n204), .B(n203), .S(n608), .Z(n205) );
  MUX2_X1 U808 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n615), .Z(n206) );
  MUX2_X1 U809 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n615), .Z(n207) );
  MUX2_X1 U810 ( .A(n207), .B(n206), .S(n610), .Z(n208) );
  MUX2_X1 U811 ( .A(n208), .B(n205), .S(n607), .Z(n209) );
  MUX2_X1 U812 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U813 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U814 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n615), .Z(n211) );
  MUX2_X1 U815 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n615), .Z(n212) );
  MUX2_X1 U816 ( .A(n212), .B(n211), .S(n608), .Z(n213) );
  MUX2_X1 U817 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n615), .Z(n214) );
  MUX2_X1 U818 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n615), .Z(n215) );
  MUX2_X1 U819 ( .A(n215), .B(n214), .S(n608), .Z(n216) );
  MUX2_X1 U820 ( .A(n216), .B(n213), .S(n607), .Z(n217) );
  MUX2_X1 U821 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n611), .Z(n218) );
  MUX2_X1 U822 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n611), .Z(n219) );
  MUX2_X1 U823 ( .A(n219), .B(n218), .S(n608), .Z(n220) );
  MUX2_X1 U824 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n614), .Z(n221) );
  MUX2_X1 U825 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n615), .Z(n222) );
  MUX2_X1 U826 ( .A(n222), .B(n221), .S(n610), .Z(n223) );
  MUX2_X1 U827 ( .A(n223), .B(n220), .S(n607), .Z(n224) );
  MUX2_X1 U828 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U829 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n614), .Z(n226) );
  MUX2_X1 U830 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n614), .Z(n227) );
  MUX2_X1 U831 ( .A(n227), .B(n226), .S(n608), .Z(n228) );
  MUX2_X1 U832 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n615), .Z(n229) );
  MUX2_X1 U833 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n613), .Z(n595) );
  MUX2_X1 U834 ( .A(n595), .B(n229), .S(n610), .Z(n596) );
  MUX2_X1 U835 ( .A(n596), .B(n228), .S(n607), .Z(n597) );
  MUX2_X1 U836 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n613), .Z(n598) );
  MUX2_X1 U837 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n615), .Z(n599) );
  MUX2_X1 U838 ( .A(n599), .B(n598), .S(n608), .Z(n600) );
  MUX2_X1 U839 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n613), .Z(n601) );
  MUX2_X1 U840 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n614), .Z(n602) );
  MUX2_X1 U841 ( .A(n602), .B(n601), .S(n608), .Z(n603) );
  MUX2_X1 U842 ( .A(n603), .B(n600), .S(n607), .Z(n604) );
  MUX2_X1 U843 ( .A(n604), .B(n597), .S(N13), .Z(n605) );
  MUX2_X1 U844 ( .A(n605), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U845 ( .A(N11), .Z(n608) );
  INV_X1 U846 ( .A(N10), .ZN(n617) );
  INV_X1 U847 ( .A(N11), .ZN(n618) );
  INV_X1 U848 ( .A(data_in[0]), .ZN(n619) );
  INV_X1 U849 ( .A(data_in[1]), .ZN(n620) );
  INV_X1 U850 ( .A(data_in[2]), .ZN(n621) );
  INV_X1 U851 ( .A(data_in[3]), .ZN(n622) );
  INV_X1 U852 ( .A(data_in[4]), .ZN(n623) );
  INV_X1 U853 ( .A(data_in[5]), .ZN(n624) );
  INV_X1 U854 ( .A(data_in[6]), .ZN(n625) );
  INV_X1 U855 ( .A(data_in[7]), .ZN(n626) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_26 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n627), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n628), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n629), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n630), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n631), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n632), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n633), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n634), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n635), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n636), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n637), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n638), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n639), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n640), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n641), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n642), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n643), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n644), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n645), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n646), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n647), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n648), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n649), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n650), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n651), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n652), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n653), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n654), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n655), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n656), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n657), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n658), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n659), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n660), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n661), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n662), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n663), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n664), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n665), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n666), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n667), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n668), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n669), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n670), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n671), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n672), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n673), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n674), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n675), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n676), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n677), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n678), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n679), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n680), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n681), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n682), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n683), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n684), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n685), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n686), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n687), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n688), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n689), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n690), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n691), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n692), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n693), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n694), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n695), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n696), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n697), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n698), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n699), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n700), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n701), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n702), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n703), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n704), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n705), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n706), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n707), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n708), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n709), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n710), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n711), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n712), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n713), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n714), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n715), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n716), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n717), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n718), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n719), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n720), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n721), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n722), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n723), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n724), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n725), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n726), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n727), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n728), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n729), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n730), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n731), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n732), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n733), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n734), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n735), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n736), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n737), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n738), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n739), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n740), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n741), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n742), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n743), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n744), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n745), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n746), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n747), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n748), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n749), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n750), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n751), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n752), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n753), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n754), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n755), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n756), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n757), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n758), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n759), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n760), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n761), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n762), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n763), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n764), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n765), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n766), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n767), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n768), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n769), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n770), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n771), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n772), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n773), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n774), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n775), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n776), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n777), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n778), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n779), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n780), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n781), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n782), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n783), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n784), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n785), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n786), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n787), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n788), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n789), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n790), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n791), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n792), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n793), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n794), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n795), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n796), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n797), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n798), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n799), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n800), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n801), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n802), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n803), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n804), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n805), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n806), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n807), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n808), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n809), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n810), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n811), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n812), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n813), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n814), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n815), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n816), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n817), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n818), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n846), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n847), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n848), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n849), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n850), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n851), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n852), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n853), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n854), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n855), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n856), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n857), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n858), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n859), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n860), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n861), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n862), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n863), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n864), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n865), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n866), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n867), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n868), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n869), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n870), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n871), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n872), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n873), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n874), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n875), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n876), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n877), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n878), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n879), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n880), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n881), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n882), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n883), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n884), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n885), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n886), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n887), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n888), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n889), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n890), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n891), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n892), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n893), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n894), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n895), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n896), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n897), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n898), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n899), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n900), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n901), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n902), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n903), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n904), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n905), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n906), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n907), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n908), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n909), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  BUF_X1 U3 ( .A(N10), .Z(n613) );
  BUF_X1 U4 ( .A(n616), .Z(n614) );
  BUF_X1 U5 ( .A(n616), .Z(n615) );
  BUF_X1 U6 ( .A(n616), .Z(n612) );
  BUF_X1 U7 ( .A(n616), .Z(n611) );
  BUF_X1 U8 ( .A(N11), .Z(n609) );
  BUF_X1 U9 ( .A(N11), .Z(n610) );
  BUF_X1 U10 ( .A(N10), .Z(n616) );
  NOR3_X1 U11 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1201) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(n617), .ZN(n1190) );
  NOR3_X1 U13 ( .A1(N10), .A2(N12), .A3(n618), .ZN(n1180) );
  NOR3_X1 U14 ( .A1(n617), .A2(N12), .A3(n618), .ZN(n1170) );
  INV_X1 U15 ( .A(n1127), .ZN(n842) );
  INV_X1 U16 ( .A(n1117), .ZN(n841) );
  INV_X1 U17 ( .A(n1108), .ZN(n840) );
  INV_X1 U18 ( .A(n1099), .ZN(n839) );
  INV_X1 U19 ( .A(n1054), .ZN(n834) );
  INV_X1 U20 ( .A(n1044), .ZN(n833) );
  INV_X1 U21 ( .A(n1035), .ZN(n832) );
  INV_X1 U22 ( .A(n1026), .ZN(n831) );
  INV_X1 U23 ( .A(n981), .ZN(n826) );
  INV_X1 U24 ( .A(n971), .ZN(n825) );
  INV_X1 U25 ( .A(n962), .ZN(n824) );
  INV_X1 U26 ( .A(n953), .ZN(n823) );
  INV_X1 U27 ( .A(n1090), .ZN(n838) );
  INV_X1 U28 ( .A(n1081), .ZN(n837) );
  INV_X1 U29 ( .A(n1072), .ZN(n836) );
  INV_X1 U30 ( .A(n1063), .ZN(n835) );
  INV_X1 U31 ( .A(n944), .ZN(n822) );
  INV_X1 U32 ( .A(n935), .ZN(n821) );
  INV_X1 U33 ( .A(n926), .ZN(n820) );
  INV_X1 U34 ( .A(n917), .ZN(n819) );
  INV_X1 U35 ( .A(n1017), .ZN(n830) );
  INV_X1 U36 ( .A(n1008), .ZN(n829) );
  INV_X1 U37 ( .A(n999), .ZN(n828) );
  INV_X1 U38 ( .A(n990), .ZN(n827) );
  BUF_X1 U39 ( .A(N12), .Z(n607) );
  INV_X1 U40 ( .A(N13), .ZN(n844) );
  AND3_X1 U41 ( .A1(n617), .A2(n618), .A3(N12), .ZN(n1160) );
  AND3_X1 U42 ( .A1(N10), .A2(n618), .A3(N12), .ZN(n1150) );
  AND3_X1 U43 ( .A1(N11), .A2(n617), .A3(N12), .ZN(n1140) );
  AND3_X1 U44 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1130) );
  BUF_X1 U45 ( .A(N12), .Z(n606) );
  INV_X1 U46 ( .A(N14), .ZN(n845) );
  NAND2_X1 U47 ( .A1(n1190), .A2(n1200), .ZN(n1199) );
  NAND2_X1 U48 ( .A1(n1180), .A2(n1200), .ZN(n1189) );
  NAND2_X1 U49 ( .A1(n1170), .A2(n1200), .ZN(n1179) );
  NAND2_X1 U50 ( .A1(n1160), .A2(n1200), .ZN(n1169) );
  NAND2_X1 U51 ( .A1(n1150), .A2(n1200), .ZN(n1159) );
  NAND2_X1 U52 ( .A1(n1140), .A2(n1200), .ZN(n1149) );
  NAND2_X1 U53 ( .A1(n1130), .A2(n1200), .ZN(n1139) );
  NAND2_X1 U54 ( .A1(n1201), .A2(n1200), .ZN(n1210) );
  NAND2_X1 U55 ( .A1(n1119), .A2(n1201), .ZN(n1127) );
  NAND2_X1 U56 ( .A1(n1119), .A2(n1190), .ZN(n1117) );
  NAND2_X1 U57 ( .A1(n1119), .A2(n1180), .ZN(n1108) );
  NAND2_X1 U58 ( .A1(n1119), .A2(n1170), .ZN(n1099) );
  NAND2_X1 U59 ( .A1(n1046), .A2(n1201), .ZN(n1054) );
  NAND2_X1 U60 ( .A1(n1046), .A2(n1190), .ZN(n1044) );
  NAND2_X1 U61 ( .A1(n1046), .A2(n1180), .ZN(n1035) );
  NAND2_X1 U62 ( .A1(n1046), .A2(n1170), .ZN(n1026) );
  NAND2_X1 U63 ( .A1(n973), .A2(n1201), .ZN(n981) );
  NAND2_X1 U64 ( .A1(n973), .A2(n1190), .ZN(n971) );
  NAND2_X1 U65 ( .A1(n973), .A2(n1180), .ZN(n962) );
  NAND2_X1 U66 ( .A1(n973), .A2(n1170), .ZN(n953) );
  NAND2_X1 U67 ( .A1(n1119), .A2(n1160), .ZN(n1090) );
  NAND2_X1 U68 ( .A1(n1119), .A2(n1150), .ZN(n1081) );
  NAND2_X1 U69 ( .A1(n1119), .A2(n1140), .ZN(n1072) );
  NAND2_X1 U70 ( .A1(n1119), .A2(n1130), .ZN(n1063) );
  NAND2_X1 U71 ( .A1(n1046), .A2(n1160), .ZN(n1017) );
  NAND2_X1 U72 ( .A1(n1046), .A2(n1150), .ZN(n1008) );
  NAND2_X1 U73 ( .A1(n1046), .A2(n1140), .ZN(n999) );
  NAND2_X1 U74 ( .A1(n1046), .A2(n1130), .ZN(n990) );
  NAND2_X1 U75 ( .A1(n973), .A2(n1160), .ZN(n944) );
  NAND2_X1 U76 ( .A1(n973), .A2(n1150), .ZN(n935) );
  NAND2_X1 U77 ( .A1(n973), .A2(n1140), .ZN(n926) );
  NAND2_X1 U78 ( .A1(n973), .A2(n1130), .ZN(n917) );
  AND3_X1 U79 ( .A1(n844), .A2(n845), .A3(n1129), .ZN(n1200) );
  AND3_X1 U80 ( .A1(N13), .A2(n1129), .A3(N14), .ZN(n973) );
  AND3_X1 U81 ( .A1(n1129), .A2(n845), .A3(N13), .ZN(n1119) );
  AND3_X1 U82 ( .A1(n1129), .A2(n844), .A3(N14), .ZN(n1046) );
  NOR2_X1 U83 ( .A1(n843), .A2(addr[5]), .ZN(n1129) );
  INV_X1 U84 ( .A(wr_en), .ZN(n843) );
  OAI21_X1 U85 ( .B1(n619), .B2(n1169), .A(n1168), .ZN(n877) );
  NAND2_X1 U86 ( .A1(\mem[4][0] ), .A2(n1169), .ZN(n1168) );
  OAI21_X1 U87 ( .B1(n620), .B2(n1169), .A(n1167), .ZN(n876) );
  NAND2_X1 U88 ( .A1(\mem[4][1] ), .A2(n1169), .ZN(n1167) );
  OAI21_X1 U89 ( .B1(n621), .B2(n1169), .A(n1166), .ZN(n875) );
  NAND2_X1 U90 ( .A1(\mem[4][2] ), .A2(n1169), .ZN(n1166) );
  OAI21_X1 U91 ( .B1(n622), .B2(n1169), .A(n1165), .ZN(n874) );
  NAND2_X1 U92 ( .A1(\mem[4][3] ), .A2(n1169), .ZN(n1165) );
  OAI21_X1 U93 ( .B1(n623), .B2(n1169), .A(n1164), .ZN(n873) );
  NAND2_X1 U94 ( .A1(\mem[4][4] ), .A2(n1169), .ZN(n1164) );
  OAI21_X1 U95 ( .B1(n624), .B2(n1169), .A(n1163), .ZN(n872) );
  NAND2_X1 U96 ( .A1(\mem[4][5] ), .A2(n1169), .ZN(n1163) );
  OAI21_X1 U97 ( .B1(n625), .B2(n1169), .A(n1162), .ZN(n871) );
  NAND2_X1 U98 ( .A1(\mem[4][6] ), .A2(n1169), .ZN(n1162) );
  OAI21_X1 U99 ( .B1(n626), .B2(n1169), .A(n1161), .ZN(n870) );
  NAND2_X1 U100 ( .A1(\mem[4][7] ), .A2(n1169), .ZN(n1161) );
  OAI21_X1 U101 ( .B1(n619), .B2(n1149), .A(n1148), .ZN(n861) );
  NAND2_X1 U102 ( .A1(\mem[6][0] ), .A2(n1149), .ZN(n1148) );
  OAI21_X1 U103 ( .B1(n620), .B2(n1149), .A(n1147), .ZN(n860) );
  NAND2_X1 U104 ( .A1(\mem[6][1] ), .A2(n1149), .ZN(n1147) );
  OAI21_X1 U105 ( .B1(n621), .B2(n1149), .A(n1146), .ZN(n859) );
  NAND2_X1 U106 ( .A1(\mem[6][2] ), .A2(n1149), .ZN(n1146) );
  OAI21_X1 U107 ( .B1(n622), .B2(n1149), .A(n1145), .ZN(n858) );
  NAND2_X1 U108 ( .A1(\mem[6][3] ), .A2(n1149), .ZN(n1145) );
  OAI21_X1 U109 ( .B1(n623), .B2(n1149), .A(n1144), .ZN(n857) );
  NAND2_X1 U110 ( .A1(\mem[6][4] ), .A2(n1149), .ZN(n1144) );
  OAI21_X1 U111 ( .B1(n624), .B2(n1149), .A(n1143), .ZN(n856) );
  NAND2_X1 U112 ( .A1(\mem[6][5] ), .A2(n1149), .ZN(n1143) );
  OAI21_X1 U113 ( .B1(n625), .B2(n1149), .A(n1142), .ZN(n855) );
  NAND2_X1 U114 ( .A1(\mem[6][6] ), .A2(n1149), .ZN(n1142) );
  OAI21_X1 U115 ( .B1(n626), .B2(n1149), .A(n1141), .ZN(n854) );
  NAND2_X1 U116 ( .A1(\mem[6][7] ), .A2(n1149), .ZN(n1141) );
  OAI21_X1 U117 ( .B1(n619), .B2(n1139), .A(n1138), .ZN(n853) );
  NAND2_X1 U118 ( .A1(\mem[7][0] ), .A2(n1139), .ZN(n1138) );
  OAI21_X1 U119 ( .B1(n620), .B2(n1139), .A(n1137), .ZN(n852) );
  NAND2_X1 U120 ( .A1(\mem[7][1] ), .A2(n1139), .ZN(n1137) );
  OAI21_X1 U121 ( .B1(n621), .B2(n1139), .A(n1136), .ZN(n851) );
  NAND2_X1 U122 ( .A1(\mem[7][2] ), .A2(n1139), .ZN(n1136) );
  OAI21_X1 U123 ( .B1(n622), .B2(n1139), .A(n1135), .ZN(n850) );
  NAND2_X1 U124 ( .A1(\mem[7][3] ), .A2(n1139), .ZN(n1135) );
  OAI21_X1 U125 ( .B1(n623), .B2(n1139), .A(n1134), .ZN(n849) );
  NAND2_X1 U126 ( .A1(\mem[7][4] ), .A2(n1139), .ZN(n1134) );
  OAI21_X1 U127 ( .B1(n624), .B2(n1139), .A(n1133), .ZN(n848) );
  NAND2_X1 U128 ( .A1(\mem[7][5] ), .A2(n1139), .ZN(n1133) );
  OAI21_X1 U129 ( .B1(n625), .B2(n1139), .A(n1132), .ZN(n847) );
  NAND2_X1 U130 ( .A1(\mem[7][6] ), .A2(n1139), .ZN(n1132) );
  OAI21_X1 U131 ( .B1(n626), .B2(n1139), .A(n1131), .ZN(n846) );
  NAND2_X1 U132 ( .A1(\mem[7][7] ), .A2(n1139), .ZN(n1131) );
  OAI21_X1 U133 ( .B1(n619), .B2(n1199), .A(n1198), .ZN(n901) );
  NAND2_X1 U134 ( .A1(\mem[1][0] ), .A2(n1199), .ZN(n1198) );
  OAI21_X1 U135 ( .B1(n620), .B2(n1199), .A(n1197), .ZN(n900) );
  NAND2_X1 U136 ( .A1(\mem[1][1] ), .A2(n1199), .ZN(n1197) );
  OAI21_X1 U137 ( .B1(n621), .B2(n1199), .A(n1196), .ZN(n899) );
  NAND2_X1 U138 ( .A1(\mem[1][2] ), .A2(n1199), .ZN(n1196) );
  OAI21_X1 U139 ( .B1(n622), .B2(n1199), .A(n1195), .ZN(n898) );
  NAND2_X1 U140 ( .A1(\mem[1][3] ), .A2(n1199), .ZN(n1195) );
  OAI21_X1 U141 ( .B1(n623), .B2(n1199), .A(n1194), .ZN(n897) );
  NAND2_X1 U142 ( .A1(\mem[1][4] ), .A2(n1199), .ZN(n1194) );
  OAI21_X1 U143 ( .B1(n624), .B2(n1199), .A(n1193), .ZN(n896) );
  NAND2_X1 U144 ( .A1(\mem[1][5] ), .A2(n1199), .ZN(n1193) );
  OAI21_X1 U145 ( .B1(n625), .B2(n1199), .A(n1192), .ZN(n895) );
  NAND2_X1 U146 ( .A1(\mem[1][6] ), .A2(n1199), .ZN(n1192) );
  OAI21_X1 U147 ( .B1(n626), .B2(n1199), .A(n1191), .ZN(n894) );
  NAND2_X1 U148 ( .A1(\mem[1][7] ), .A2(n1199), .ZN(n1191) );
  OAI21_X1 U149 ( .B1(n619), .B2(n1189), .A(n1188), .ZN(n893) );
  NAND2_X1 U150 ( .A1(\mem[2][0] ), .A2(n1189), .ZN(n1188) );
  OAI21_X1 U151 ( .B1(n620), .B2(n1189), .A(n1187), .ZN(n892) );
  NAND2_X1 U152 ( .A1(\mem[2][1] ), .A2(n1189), .ZN(n1187) );
  OAI21_X1 U153 ( .B1(n621), .B2(n1189), .A(n1186), .ZN(n891) );
  NAND2_X1 U154 ( .A1(\mem[2][2] ), .A2(n1189), .ZN(n1186) );
  OAI21_X1 U155 ( .B1(n622), .B2(n1189), .A(n1185), .ZN(n890) );
  NAND2_X1 U156 ( .A1(\mem[2][3] ), .A2(n1189), .ZN(n1185) );
  OAI21_X1 U157 ( .B1(n623), .B2(n1189), .A(n1184), .ZN(n889) );
  NAND2_X1 U158 ( .A1(\mem[2][4] ), .A2(n1189), .ZN(n1184) );
  OAI21_X1 U159 ( .B1(n624), .B2(n1189), .A(n1183), .ZN(n888) );
  NAND2_X1 U160 ( .A1(\mem[2][5] ), .A2(n1189), .ZN(n1183) );
  OAI21_X1 U161 ( .B1(n625), .B2(n1189), .A(n1182), .ZN(n887) );
  NAND2_X1 U162 ( .A1(\mem[2][6] ), .A2(n1189), .ZN(n1182) );
  OAI21_X1 U163 ( .B1(n626), .B2(n1189), .A(n1181), .ZN(n886) );
  NAND2_X1 U164 ( .A1(\mem[2][7] ), .A2(n1189), .ZN(n1181) );
  OAI21_X1 U165 ( .B1(n619), .B2(n1179), .A(n1178), .ZN(n885) );
  NAND2_X1 U166 ( .A1(\mem[3][0] ), .A2(n1179), .ZN(n1178) );
  OAI21_X1 U167 ( .B1(n620), .B2(n1179), .A(n1177), .ZN(n884) );
  NAND2_X1 U168 ( .A1(\mem[3][1] ), .A2(n1179), .ZN(n1177) );
  OAI21_X1 U169 ( .B1(n621), .B2(n1179), .A(n1176), .ZN(n883) );
  NAND2_X1 U170 ( .A1(\mem[3][2] ), .A2(n1179), .ZN(n1176) );
  OAI21_X1 U171 ( .B1(n622), .B2(n1179), .A(n1175), .ZN(n882) );
  NAND2_X1 U172 ( .A1(\mem[3][3] ), .A2(n1179), .ZN(n1175) );
  OAI21_X1 U173 ( .B1(n623), .B2(n1179), .A(n1174), .ZN(n881) );
  NAND2_X1 U174 ( .A1(\mem[3][4] ), .A2(n1179), .ZN(n1174) );
  OAI21_X1 U175 ( .B1(n624), .B2(n1179), .A(n1173), .ZN(n880) );
  NAND2_X1 U176 ( .A1(\mem[3][5] ), .A2(n1179), .ZN(n1173) );
  OAI21_X1 U177 ( .B1(n625), .B2(n1179), .A(n1172), .ZN(n879) );
  NAND2_X1 U178 ( .A1(\mem[3][6] ), .A2(n1179), .ZN(n1172) );
  OAI21_X1 U179 ( .B1(n626), .B2(n1179), .A(n1171), .ZN(n878) );
  NAND2_X1 U180 ( .A1(\mem[3][7] ), .A2(n1179), .ZN(n1171) );
  OAI21_X1 U181 ( .B1(n619), .B2(n1159), .A(n1158), .ZN(n869) );
  NAND2_X1 U182 ( .A1(\mem[5][0] ), .A2(n1159), .ZN(n1158) );
  OAI21_X1 U183 ( .B1(n620), .B2(n1159), .A(n1157), .ZN(n868) );
  NAND2_X1 U184 ( .A1(\mem[5][1] ), .A2(n1159), .ZN(n1157) );
  OAI21_X1 U185 ( .B1(n621), .B2(n1159), .A(n1156), .ZN(n867) );
  NAND2_X1 U186 ( .A1(\mem[5][2] ), .A2(n1159), .ZN(n1156) );
  OAI21_X1 U187 ( .B1(n622), .B2(n1159), .A(n1155), .ZN(n866) );
  NAND2_X1 U188 ( .A1(\mem[5][3] ), .A2(n1159), .ZN(n1155) );
  OAI21_X1 U189 ( .B1(n623), .B2(n1159), .A(n1154), .ZN(n865) );
  NAND2_X1 U190 ( .A1(\mem[5][4] ), .A2(n1159), .ZN(n1154) );
  OAI21_X1 U191 ( .B1(n624), .B2(n1159), .A(n1153), .ZN(n864) );
  NAND2_X1 U192 ( .A1(\mem[5][5] ), .A2(n1159), .ZN(n1153) );
  OAI21_X1 U193 ( .B1(n625), .B2(n1159), .A(n1152), .ZN(n863) );
  NAND2_X1 U194 ( .A1(\mem[5][6] ), .A2(n1159), .ZN(n1152) );
  OAI21_X1 U195 ( .B1(n626), .B2(n1159), .A(n1151), .ZN(n862) );
  NAND2_X1 U196 ( .A1(\mem[5][7] ), .A2(n1159), .ZN(n1151) );
  OAI21_X1 U197 ( .B1(n1210), .B2(n619), .A(n1209), .ZN(n909) );
  NAND2_X1 U198 ( .A1(\mem[0][0] ), .A2(n1210), .ZN(n1209) );
  OAI21_X1 U199 ( .B1(n1210), .B2(n620), .A(n1208), .ZN(n908) );
  NAND2_X1 U200 ( .A1(\mem[0][1] ), .A2(n1210), .ZN(n1208) );
  OAI21_X1 U201 ( .B1(n1210), .B2(n621), .A(n1207), .ZN(n907) );
  NAND2_X1 U202 ( .A1(\mem[0][2] ), .A2(n1210), .ZN(n1207) );
  OAI21_X1 U203 ( .B1(n1210), .B2(n622), .A(n1206), .ZN(n906) );
  NAND2_X1 U204 ( .A1(\mem[0][3] ), .A2(n1210), .ZN(n1206) );
  OAI21_X1 U205 ( .B1(n1210), .B2(n623), .A(n1205), .ZN(n905) );
  NAND2_X1 U206 ( .A1(\mem[0][4] ), .A2(n1210), .ZN(n1205) );
  OAI21_X1 U207 ( .B1(n1210), .B2(n624), .A(n1204), .ZN(n904) );
  NAND2_X1 U208 ( .A1(\mem[0][5] ), .A2(n1210), .ZN(n1204) );
  OAI21_X1 U209 ( .B1(n1210), .B2(n625), .A(n1203), .ZN(n903) );
  NAND2_X1 U210 ( .A1(\mem[0][6] ), .A2(n1210), .ZN(n1203) );
  OAI21_X1 U211 ( .B1(n1210), .B2(n626), .A(n1202), .ZN(n902) );
  NAND2_X1 U212 ( .A1(\mem[0][7] ), .A2(n1210), .ZN(n1202) );
  INV_X1 U213 ( .A(n1128), .ZN(n818) );
  AOI22_X1 U214 ( .A1(data_in[0]), .A2(n842), .B1(n1127), .B2(\mem[8][0] ), 
        .ZN(n1128) );
  INV_X1 U215 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U216 ( .A1(data_in[1]), .A2(n842), .B1(n1127), .B2(\mem[8][1] ), 
        .ZN(n1126) );
  INV_X1 U217 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U218 ( .A1(data_in[2]), .A2(n842), .B1(n1127), .B2(\mem[8][2] ), 
        .ZN(n1125) );
  INV_X1 U219 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U220 ( .A1(data_in[3]), .A2(n842), .B1(n1127), .B2(\mem[8][3] ), 
        .ZN(n1124) );
  INV_X1 U221 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U222 ( .A1(data_in[4]), .A2(n842), .B1(n1127), .B2(\mem[8][4] ), 
        .ZN(n1123) );
  INV_X1 U223 ( .A(n1122), .ZN(n813) );
  AOI22_X1 U224 ( .A1(data_in[5]), .A2(n842), .B1(n1127), .B2(\mem[8][5] ), 
        .ZN(n1122) );
  INV_X1 U225 ( .A(n1121), .ZN(n812) );
  AOI22_X1 U226 ( .A1(data_in[6]), .A2(n842), .B1(n1127), .B2(\mem[8][6] ), 
        .ZN(n1121) );
  INV_X1 U227 ( .A(n1120), .ZN(n811) );
  AOI22_X1 U228 ( .A1(data_in[7]), .A2(n842), .B1(n1127), .B2(\mem[8][7] ), 
        .ZN(n1120) );
  INV_X1 U229 ( .A(n1118), .ZN(n810) );
  AOI22_X1 U230 ( .A1(data_in[0]), .A2(n841), .B1(n1117), .B2(\mem[9][0] ), 
        .ZN(n1118) );
  INV_X1 U231 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U232 ( .A1(data_in[1]), .A2(n841), .B1(n1117), .B2(\mem[9][1] ), 
        .ZN(n1116) );
  INV_X1 U233 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U234 ( .A1(data_in[2]), .A2(n841), .B1(n1117), .B2(\mem[9][2] ), 
        .ZN(n1115) );
  INV_X1 U235 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U236 ( .A1(data_in[3]), .A2(n841), .B1(n1117), .B2(\mem[9][3] ), 
        .ZN(n1114) );
  INV_X1 U237 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U238 ( .A1(data_in[4]), .A2(n841), .B1(n1117), .B2(\mem[9][4] ), 
        .ZN(n1113) );
  INV_X1 U239 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U240 ( .A1(data_in[5]), .A2(n841), .B1(n1117), .B2(\mem[9][5] ), 
        .ZN(n1112) );
  INV_X1 U241 ( .A(n1111), .ZN(n804) );
  AOI22_X1 U242 ( .A1(data_in[6]), .A2(n841), .B1(n1117), .B2(\mem[9][6] ), 
        .ZN(n1111) );
  INV_X1 U243 ( .A(n1110), .ZN(n803) );
  AOI22_X1 U244 ( .A1(data_in[7]), .A2(n841), .B1(n1117), .B2(\mem[9][7] ), 
        .ZN(n1110) );
  INV_X1 U245 ( .A(n1109), .ZN(n802) );
  AOI22_X1 U246 ( .A1(data_in[0]), .A2(n840), .B1(n1108), .B2(\mem[10][0] ), 
        .ZN(n1109) );
  INV_X1 U247 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U248 ( .A1(data_in[1]), .A2(n840), .B1(n1108), .B2(\mem[10][1] ), 
        .ZN(n1107) );
  INV_X1 U249 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U250 ( .A1(data_in[2]), .A2(n840), .B1(n1108), .B2(\mem[10][2] ), 
        .ZN(n1106) );
  INV_X1 U251 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U252 ( .A1(data_in[3]), .A2(n840), .B1(n1108), .B2(\mem[10][3] ), 
        .ZN(n1105) );
  INV_X1 U253 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U254 ( .A1(data_in[4]), .A2(n840), .B1(n1108), .B2(\mem[10][4] ), 
        .ZN(n1104) );
  INV_X1 U255 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U256 ( .A1(data_in[5]), .A2(n840), .B1(n1108), .B2(\mem[10][5] ), 
        .ZN(n1103) );
  INV_X1 U257 ( .A(n1102), .ZN(n796) );
  AOI22_X1 U258 ( .A1(data_in[6]), .A2(n840), .B1(n1108), .B2(\mem[10][6] ), 
        .ZN(n1102) );
  INV_X1 U259 ( .A(n1101), .ZN(n795) );
  AOI22_X1 U260 ( .A1(data_in[7]), .A2(n840), .B1(n1108), .B2(\mem[10][7] ), 
        .ZN(n1101) );
  INV_X1 U261 ( .A(n1100), .ZN(n794) );
  AOI22_X1 U262 ( .A1(data_in[0]), .A2(n839), .B1(n1099), .B2(\mem[11][0] ), 
        .ZN(n1100) );
  INV_X1 U263 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U264 ( .A1(data_in[1]), .A2(n839), .B1(n1099), .B2(\mem[11][1] ), 
        .ZN(n1098) );
  INV_X1 U265 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U266 ( .A1(data_in[2]), .A2(n839), .B1(n1099), .B2(\mem[11][2] ), 
        .ZN(n1097) );
  INV_X1 U267 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U268 ( .A1(data_in[3]), .A2(n839), .B1(n1099), .B2(\mem[11][3] ), 
        .ZN(n1096) );
  INV_X1 U269 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U270 ( .A1(data_in[4]), .A2(n839), .B1(n1099), .B2(\mem[11][4] ), 
        .ZN(n1095) );
  INV_X1 U271 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U272 ( .A1(data_in[5]), .A2(n839), .B1(n1099), .B2(\mem[11][5] ), 
        .ZN(n1094) );
  INV_X1 U273 ( .A(n1093), .ZN(n788) );
  AOI22_X1 U274 ( .A1(data_in[6]), .A2(n839), .B1(n1099), .B2(\mem[11][6] ), 
        .ZN(n1093) );
  INV_X1 U275 ( .A(n1092), .ZN(n787) );
  AOI22_X1 U276 ( .A1(data_in[7]), .A2(n839), .B1(n1099), .B2(\mem[11][7] ), 
        .ZN(n1092) );
  INV_X1 U277 ( .A(n1091), .ZN(n786) );
  AOI22_X1 U278 ( .A1(data_in[0]), .A2(n838), .B1(n1090), .B2(\mem[12][0] ), 
        .ZN(n1091) );
  INV_X1 U279 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U280 ( .A1(data_in[1]), .A2(n838), .B1(n1090), .B2(\mem[12][1] ), 
        .ZN(n1089) );
  INV_X1 U281 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U282 ( .A1(data_in[2]), .A2(n838), .B1(n1090), .B2(\mem[12][2] ), 
        .ZN(n1088) );
  INV_X1 U283 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U284 ( .A1(data_in[3]), .A2(n838), .B1(n1090), .B2(\mem[12][3] ), 
        .ZN(n1087) );
  INV_X1 U285 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U286 ( .A1(data_in[4]), .A2(n838), .B1(n1090), .B2(\mem[12][4] ), 
        .ZN(n1086) );
  INV_X1 U287 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U288 ( .A1(data_in[5]), .A2(n838), .B1(n1090), .B2(\mem[12][5] ), 
        .ZN(n1085) );
  INV_X1 U289 ( .A(n1084), .ZN(n780) );
  AOI22_X1 U290 ( .A1(data_in[6]), .A2(n838), .B1(n1090), .B2(\mem[12][6] ), 
        .ZN(n1084) );
  INV_X1 U291 ( .A(n1083), .ZN(n779) );
  AOI22_X1 U292 ( .A1(data_in[7]), .A2(n838), .B1(n1090), .B2(\mem[12][7] ), 
        .ZN(n1083) );
  INV_X1 U293 ( .A(n1082), .ZN(n778) );
  AOI22_X1 U294 ( .A1(data_in[0]), .A2(n837), .B1(n1081), .B2(\mem[13][0] ), 
        .ZN(n1082) );
  INV_X1 U295 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U296 ( .A1(data_in[1]), .A2(n837), .B1(n1081), .B2(\mem[13][1] ), 
        .ZN(n1080) );
  INV_X1 U297 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U298 ( .A1(data_in[2]), .A2(n837), .B1(n1081), .B2(\mem[13][2] ), 
        .ZN(n1079) );
  INV_X1 U299 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U300 ( .A1(data_in[3]), .A2(n837), .B1(n1081), .B2(\mem[13][3] ), 
        .ZN(n1078) );
  INV_X1 U301 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U302 ( .A1(data_in[4]), .A2(n837), .B1(n1081), .B2(\mem[13][4] ), 
        .ZN(n1077) );
  INV_X1 U303 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U304 ( .A1(data_in[5]), .A2(n837), .B1(n1081), .B2(\mem[13][5] ), 
        .ZN(n1076) );
  INV_X1 U305 ( .A(n1075), .ZN(n772) );
  AOI22_X1 U306 ( .A1(data_in[6]), .A2(n837), .B1(n1081), .B2(\mem[13][6] ), 
        .ZN(n1075) );
  INV_X1 U307 ( .A(n1074), .ZN(n771) );
  AOI22_X1 U308 ( .A1(data_in[7]), .A2(n837), .B1(n1081), .B2(\mem[13][7] ), 
        .ZN(n1074) );
  INV_X1 U309 ( .A(n1073), .ZN(n770) );
  AOI22_X1 U310 ( .A1(data_in[0]), .A2(n836), .B1(n1072), .B2(\mem[14][0] ), 
        .ZN(n1073) );
  INV_X1 U311 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U312 ( .A1(data_in[1]), .A2(n836), .B1(n1072), .B2(\mem[14][1] ), 
        .ZN(n1071) );
  INV_X1 U313 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U314 ( .A1(data_in[2]), .A2(n836), .B1(n1072), .B2(\mem[14][2] ), 
        .ZN(n1070) );
  INV_X1 U315 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U316 ( .A1(data_in[3]), .A2(n836), .B1(n1072), .B2(\mem[14][3] ), 
        .ZN(n1069) );
  INV_X1 U317 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U318 ( .A1(data_in[4]), .A2(n836), .B1(n1072), .B2(\mem[14][4] ), 
        .ZN(n1068) );
  INV_X1 U319 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U320 ( .A1(data_in[5]), .A2(n836), .B1(n1072), .B2(\mem[14][5] ), 
        .ZN(n1067) );
  INV_X1 U321 ( .A(n1066), .ZN(n764) );
  AOI22_X1 U322 ( .A1(data_in[6]), .A2(n836), .B1(n1072), .B2(\mem[14][6] ), 
        .ZN(n1066) );
  INV_X1 U323 ( .A(n1065), .ZN(n763) );
  AOI22_X1 U324 ( .A1(data_in[7]), .A2(n836), .B1(n1072), .B2(\mem[14][7] ), 
        .ZN(n1065) );
  INV_X1 U325 ( .A(n1064), .ZN(n762) );
  AOI22_X1 U326 ( .A1(data_in[0]), .A2(n835), .B1(n1063), .B2(\mem[15][0] ), 
        .ZN(n1064) );
  INV_X1 U327 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U328 ( .A1(data_in[1]), .A2(n835), .B1(n1063), .B2(\mem[15][1] ), 
        .ZN(n1062) );
  INV_X1 U329 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U330 ( .A1(data_in[2]), .A2(n835), .B1(n1063), .B2(\mem[15][2] ), 
        .ZN(n1061) );
  INV_X1 U331 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U332 ( .A1(data_in[3]), .A2(n835), .B1(n1063), .B2(\mem[15][3] ), 
        .ZN(n1060) );
  INV_X1 U333 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U334 ( .A1(data_in[4]), .A2(n835), .B1(n1063), .B2(\mem[15][4] ), 
        .ZN(n1059) );
  INV_X1 U335 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U336 ( .A1(data_in[5]), .A2(n835), .B1(n1063), .B2(\mem[15][5] ), 
        .ZN(n1058) );
  INV_X1 U337 ( .A(n1057), .ZN(n756) );
  AOI22_X1 U338 ( .A1(data_in[6]), .A2(n835), .B1(n1063), .B2(\mem[15][6] ), 
        .ZN(n1057) );
  INV_X1 U339 ( .A(n1056), .ZN(n755) );
  AOI22_X1 U340 ( .A1(data_in[7]), .A2(n835), .B1(n1063), .B2(\mem[15][7] ), 
        .ZN(n1056) );
  INV_X1 U341 ( .A(n1055), .ZN(n754) );
  AOI22_X1 U342 ( .A1(data_in[0]), .A2(n834), .B1(n1054), .B2(\mem[16][0] ), 
        .ZN(n1055) );
  INV_X1 U343 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U344 ( .A1(data_in[1]), .A2(n834), .B1(n1054), .B2(\mem[16][1] ), 
        .ZN(n1053) );
  INV_X1 U345 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U346 ( .A1(data_in[2]), .A2(n834), .B1(n1054), .B2(\mem[16][2] ), 
        .ZN(n1052) );
  INV_X1 U347 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U348 ( .A1(data_in[3]), .A2(n834), .B1(n1054), .B2(\mem[16][3] ), 
        .ZN(n1051) );
  INV_X1 U349 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U350 ( .A1(data_in[4]), .A2(n834), .B1(n1054), .B2(\mem[16][4] ), 
        .ZN(n1050) );
  INV_X1 U351 ( .A(n1049), .ZN(n749) );
  AOI22_X1 U352 ( .A1(data_in[5]), .A2(n834), .B1(n1054), .B2(\mem[16][5] ), 
        .ZN(n1049) );
  INV_X1 U353 ( .A(n1048), .ZN(n748) );
  AOI22_X1 U354 ( .A1(data_in[6]), .A2(n834), .B1(n1054), .B2(\mem[16][6] ), 
        .ZN(n1048) );
  INV_X1 U355 ( .A(n1047), .ZN(n747) );
  AOI22_X1 U356 ( .A1(data_in[7]), .A2(n834), .B1(n1054), .B2(\mem[16][7] ), 
        .ZN(n1047) );
  INV_X1 U357 ( .A(n1045), .ZN(n746) );
  AOI22_X1 U358 ( .A1(data_in[0]), .A2(n833), .B1(n1044), .B2(\mem[17][0] ), 
        .ZN(n1045) );
  INV_X1 U359 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U360 ( .A1(data_in[1]), .A2(n833), .B1(n1044), .B2(\mem[17][1] ), 
        .ZN(n1043) );
  INV_X1 U361 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U362 ( .A1(data_in[2]), .A2(n833), .B1(n1044), .B2(\mem[17][2] ), 
        .ZN(n1042) );
  INV_X1 U363 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U364 ( .A1(data_in[3]), .A2(n833), .B1(n1044), .B2(\mem[17][3] ), 
        .ZN(n1041) );
  INV_X1 U365 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U366 ( .A1(data_in[4]), .A2(n833), .B1(n1044), .B2(\mem[17][4] ), 
        .ZN(n1040) );
  INV_X1 U367 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U368 ( .A1(data_in[5]), .A2(n833), .B1(n1044), .B2(\mem[17][5] ), 
        .ZN(n1039) );
  INV_X1 U369 ( .A(n1038), .ZN(n740) );
  AOI22_X1 U370 ( .A1(data_in[6]), .A2(n833), .B1(n1044), .B2(\mem[17][6] ), 
        .ZN(n1038) );
  INV_X1 U371 ( .A(n1037), .ZN(n739) );
  AOI22_X1 U372 ( .A1(data_in[7]), .A2(n833), .B1(n1044), .B2(\mem[17][7] ), 
        .ZN(n1037) );
  INV_X1 U373 ( .A(n1036), .ZN(n738) );
  AOI22_X1 U374 ( .A1(data_in[0]), .A2(n832), .B1(n1035), .B2(\mem[18][0] ), 
        .ZN(n1036) );
  INV_X1 U375 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U376 ( .A1(data_in[1]), .A2(n832), .B1(n1035), .B2(\mem[18][1] ), 
        .ZN(n1034) );
  INV_X1 U377 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U378 ( .A1(data_in[2]), .A2(n832), .B1(n1035), .B2(\mem[18][2] ), 
        .ZN(n1033) );
  INV_X1 U379 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U380 ( .A1(data_in[3]), .A2(n832), .B1(n1035), .B2(\mem[18][3] ), 
        .ZN(n1032) );
  INV_X1 U381 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U382 ( .A1(data_in[4]), .A2(n832), .B1(n1035), .B2(\mem[18][4] ), 
        .ZN(n1031) );
  INV_X1 U383 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U384 ( .A1(data_in[5]), .A2(n832), .B1(n1035), .B2(\mem[18][5] ), 
        .ZN(n1030) );
  INV_X1 U385 ( .A(n1029), .ZN(n732) );
  AOI22_X1 U386 ( .A1(data_in[6]), .A2(n832), .B1(n1035), .B2(\mem[18][6] ), 
        .ZN(n1029) );
  INV_X1 U387 ( .A(n1028), .ZN(n731) );
  AOI22_X1 U388 ( .A1(data_in[7]), .A2(n832), .B1(n1035), .B2(\mem[18][7] ), 
        .ZN(n1028) );
  INV_X1 U389 ( .A(n1027), .ZN(n730) );
  AOI22_X1 U390 ( .A1(data_in[0]), .A2(n831), .B1(n1026), .B2(\mem[19][0] ), 
        .ZN(n1027) );
  INV_X1 U391 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U392 ( .A1(data_in[1]), .A2(n831), .B1(n1026), .B2(\mem[19][1] ), 
        .ZN(n1025) );
  INV_X1 U393 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U394 ( .A1(data_in[2]), .A2(n831), .B1(n1026), .B2(\mem[19][2] ), 
        .ZN(n1024) );
  INV_X1 U395 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U396 ( .A1(data_in[3]), .A2(n831), .B1(n1026), .B2(\mem[19][3] ), 
        .ZN(n1023) );
  INV_X1 U397 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U398 ( .A1(data_in[4]), .A2(n831), .B1(n1026), .B2(\mem[19][4] ), 
        .ZN(n1022) );
  INV_X1 U399 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U400 ( .A1(data_in[5]), .A2(n831), .B1(n1026), .B2(\mem[19][5] ), 
        .ZN(n1021) );
  INV_X1 U401 ( .A(n1020), .ZN(n724) );
  AOI22_X1 U402 ( .A1(data_in[6]), .A2(n831), .B1(n1026), .B2(\mem[19][6] ), 
        .ZN(n1020) );
  INV_X1 U403 ( .A(n1019), .ZN(n723) );
  AOI22_X1 U404 ( .A1(data_in[7]), .A2(n831), .B1(n1026), .B2(\mem[19][7] ), 
        .ZN(n1019) );
  INV_X1 U405 ( .A(n1018), .ZN(n722) );
  AOI22_X1 U406 ( .A1(data_in[0]), .A2(n830), .B1(n1017), .B2(\mem[20][0] ), 
        .ZN(n1018) );
  INV_X1 U407 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U408 ( .A1(data_in[1]), .A2(n830), .B1(n1017), .B2(\mem[20][1] ), 
        .ZN(n1016) );
  INV_X1 U409 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U410 ( .A1(data_in[2]), .A2(n830), .B1(n1017), .B2(\mem[20][2] ), 
        .ZN(n1015) );
  INV_X1 U411 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U412 ( .A1(data_in[3]), .A2(n830), .B1(n1017), .B2(\mem[20][3] ), 
        .ZN(n1014) );
  INV_X1 U413 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U414 ( .A1(data_in[4]), .A2(n830), .B1(n1017), .B2(\mem[20][4] ), 
        .ZN(n1013) );
  INV_X1 U415 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U416 ( .A1(data_in[5]), .A2(n830), .B1(n1017), .B2(\mem[20][5] ), 
        .ZN(n1012) );
  INV_X1 U417 ( .A(n1011), .ZN(n716) );
  AOI22_X1 U418 ( .A1(data_in[6]), .A2(n830), .B1(n1017), .B2(\mem[20][6] ), 
        .ZN(n1011) );
  INV_X1 U419 ( .A(n1010), .ZN(n715) );
  AOI22_X1 U420 ( .A1(data_in[7]), .A2(n830), .B1(n1017), .B2(\mem[20][7] ), 
        .ZN(n1010) );
  INV_X1 U421 ( .A(n1009), .ZN(n714) );
  AOI22_X1 U422 ( .A1(data_in[0]), .A2(n829), .B1(n1008), .B2(\mem[21][0] ), 
        .ZN(n1009) );
  INV_X1 U423 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U424 ( .A1(data_in[1]), .A2(n829), .B1(n1008), .B2(\mem[21][1] ), 
        .ZN(n1007) );
  INV_X1 U425 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U426 ( .A1(data_in[2]), .A2(n829), .B1(n1008), .B2(\mem[21][2] ), 
        .ZN(n1006) );
  INV_X1 U427 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U428 ( .A1(data_in[3]), .A2(n829), .B1(n1008), .B2(\mem[21][3] ), 
        .ZN(n1005) );
  INV_X1 U429 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U430 ( .A1(data_in[4]), .A2(n829), .B1(n1008), .B2(\mem[21][4] ), 
        .ZN(n1004) );
  INV_X1 U431 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U432 ( .A1(data_in[5]), .A2(n829), .B1(n1008), .B2(\mem[21][5] ), 
        .ZN(n1003) );
  INV_X1 U433 ( .A(n1002), .ZN(n708) );
  AOI22_X1 U434 ( .A1(data_in[6]), .A2(n829), .B1(n1008), .B2(\mem[21][6] ), 
        .ZN(n1002) );
  INV_X1 U435 ( .A(n1001), .ZN(n707) );
  AOI22_X1 U436 ( .A1(data_in[7]), .A2(n829), .B1(n1008), .B2(\mem[21][7] ), 
        .ZN(n1001) );
  INV_X1 U437 ( .A(n1000), .ZN(n706) );
  AOI22_X1 U438 ( .A1(data_in[0]), .A2(n828), .B1(n999), .B2(\mem[22][0] ), 
        .ZN(n1000) );
  INV_X1 U439 ( .A(n998), .ZN(n705) );
  AOI22_X1 U440 ( .A1(data_in[1]), .A2(n828), .B1(n999), .B2(\mem[22][1] ), 
        .ZN(n998) );
  INV_X1 U441 ( .A(n997), .ZN(n704) );
  AOI22_X1 U442 ( .A1(data_in[2]), .A2(n828), .B1(n999), .B2(\mem[22][2] ), 
        .ZN(n997) );
  INV_X1 U443 ( .A(n996), .ZN(n703) );
  AOI22_X1 U444 ( .A1(data_in[3]), .A2(n828), .B1(n999), .B2(\mem[22][3] ), 
        .ZN(n996) );
  INV_X1 U445 ( .A(n995), .ZN(n702) );
  AOI22_X1 U446 ( .A1(data_in[4]), .A2(n828), .B1(n999), .B2(\mem[22][4] ), 
        .ZN(n995) );
  INV_X1 U447 ( .A(n994), .ZN(n701) );
  AOI22_X1 U448 ( .A1(data_in[5]), .A2(n828), .B1(n999), .B2(\mem[22][5] ), 
        .ZN(n994) );
  INV_X1 U449 ( .A(n993), .ZN(n700) );
  AOI22_X1 U450 ( .A1(data_in[6]), .A2(n828), .B1(n999), .B2(\mem[22][6] ), 
        .ZN(n993) );
  INV_X1 U451 ( .A(n992), .ZN(n699) );
  AOI22_X1 U452 ( .A1(data_in[7]), .A2(n828), .B1(n999), .B2(\mem[22][7] ), 
        .ZN(n992) );
  INV_X1 U453 ( .A(n991), .ZN(n698) );
  AOI22_X1 U454 ( .A1(data_in[0]), .A2(n827), .B1(n990), .B2(\mem[23][0] ), 
        .ZN(n991) );
  INV_X1 U455 ( .A(n989), .ZN(n697) );
  AOI22_X1 U456 ( .A1(data_in[1]), .A2(n827), .B1(n990), .B2(\mem[23][1] ), 
        .ZN(n989) );
  INV_X1 U457 ( .A(n988), .ZN(n696) );
  AOI22_X1 U458 ( .A1(data_in[2]), .A2(n827), .B1(n990), .B2(\mem[23][2] ), 
        .ZN(n988) );
  INV_X1 U459 ( .A(n987), .ZN(n695) );
  AOI22_X1 U460 ( .A1(data_in[3]), .A2(n827), .B1(n990), .B2(\mem[23][3] ), 
        .ZN(n987) );
  INV_X1 U461 ( .A(n986), .ZN(n694) );
  AOI22_X1 U462 ( .A1(data_in[4]), .A2(n827), .B1(n990), .B2(\mem[23][4] ), 
        .ZN(n986) );
  INV_X1 U463 ( .A(n985), .ZN(n693) );
  AOI22_X1 U464 ( .A1(data_in[5]), .A2(n827), .B1(n990), .B2(\mem[23][5] ), 
        .ZN(n985) );
  INV_X1 U465 ( .A(n984), .ZN(n692) );
  AOI22_X1 U466 ( .A1(data_in[6]), .A2(n827), .B1(n990), .B2(\mem[23][6] ), 
        .ZN(n984) );
  INV_X1 U467 ( .A(n983), .ZN(n691) );
  AOI22_X1 U468 ( .A1(data_in[7]), .A2(n827), .B1(n990), .B2(\mem[23][7] ), 
        .ZN(n983) );
  INV_X1 U469 ( .A(n982), .ZN(n690) );
  AOI22_X1 U470 ( .A1(data_in[0]), .A2(n826), .B1(n981), .B2(\mem[24][0] ), 
        .ZN(n982) );
  INV_X1 U471 ( .A(n980), .ZN(n689) );
  AOI22_X1 U472 ( .A1(data_in[1]), .A2(n826), .B1(n981), .B2(\mem[24][1] ), 
        .ZN(n980) );
  INV_X1 U473 ( .A(n979), .ZN(n688) );
  AOI22_X1 U474 ( .A1(data_in[2]), .A2(n826), .B1(n981), .B2(\mem[24][2] ), 
        .ZN(n979) );
  INV_X1 U475 ( .A(n978), .ZN(n687) );
  AOI22_X1 U476 ( .A1(data_in[3]), .A2(n826), .B1(n981), .B2(\mem[24][3] ), 
        .ZN(n978) );
  INV_X1 U477 ( .A(n977), .ZN(n686) );
  AOI22_X1 U478 ( .A1(data_in[4]), .A2(n826), .B1(n981), .B2(\mem[24][4] ), 
        .ZN(n977) );
  INV_X1 U479 ( .A(n976), .ZN(n685) );
  AOI22_X1 U480 ( .A1(data_in[5]), .A2(n826), .B1(n981), .B2(\mem[24][5] ), 
        .ZN(n976) );
  INV_X1 U481 ( .A(n975), .ZN(n684) );
  AOI22_X1 U482 ( .A1(data_in[6]), .A2(n826), .B1(n981), .B2(\mem[24][6] ), 
        .ZN(n975) );
  INV_X1 U483 ( .A(n974), .ZN(n683) );
  AOI22_X1 U484 ( .A1(data_in[7]), .A2(n826), .B1(n981), .B2(\mem[24][7] ), 
        .ZN(n974) );
  INV_X1 U485 ( .A(n972), .ZN(n682) );
  AOI22_X1 U486 ( .A1(data_in[0]), .A2(n825), .B1(n971), .B2(\mem[25][0] ), 
        .ZN(n972) );
  INV_X1 U487 ( .A(n970), .ZN(n681) );
  AOI22_X1 U488 ( .A1(data_in[1]), .A2(n825), .B1(n971), .B2(\mem[25][1] ), 
        .ZN(n970) );
  INV_X1 U489 ( .A(n969), .ZN(n680) );
  AOI22_X1 U490 ( .A1(data_in[2]), .A2(n825), .B1(n971), .B2(\mem[25][2] ), 
        .ZN(n969) );
  INV_X1 U491 ( .A(n968), .ZN(n679) );
  AOI22_X1 U492 ( .A1(data_in[3]), .A2(n825), .B1(n971), .B2(\mem[25][3] ), 
        .ZN(n968) );
  INV_X1 U493 ( .A(n967), .ZN(n678) );
  AOI22_X1 U494 ( .A1(data_in[4]), .A2(n825), .B1(n971), .B2(\mem[25][4] ), 
        .ZN(n967) );
  INV_X1 U495 ( .A(n966), .ZN(n677) );
  AOI22_X1 U496 ( .A1(data_in[5]), .A2(n825), .B1(n971), .B2(\mem[25][5] ), 
        .ZN(n966) );
  INV_X1 U497 ( .A(n965), .ZN(n676) );
  AOI22_X1 U498 ( .A1(data_in[6]), .A2(n825), .B1(n971), .B2(\mem[25][6] ), 
        .ZN(n965) );
  INV_X1 U499 ( .A(n964), .ZN(n675) );
  AOI22_X1 U500 ( .A1(data_in[7]), .A2(n825), .B1(n971), .B2(\mem[25][7] ), 
        .ZN(n964) );
  INV_X1 U501 ( .A(n963), .ZN(n674) );
  AOI22_X1 U502 ( .A1(data_in[0]), .A2(n824), .B1(n962), .B2(\mem[26][0] ), 
        .ZN(n963) );
  INV_X1 U503 ( .A(n961), .ZN(n673) );
  AOI22_X1 U504 ( .A1(data_in[1]), .A2(n824), .B1(n962), .B2(\mem[26][1] ), 
        .ZN(n961) );
  INV_X1 U505 ( .A(n960), .ZN(n672) );
  AOI22_X1 U506 ( .A1(data_in[2]), .A2(n824), .B1(n962), .B2(\mem[26][2] ), 
        .ZN(n960) );
  INV_X1 U507 ( .A(n959), .ZN(n671) );
  AOI22_X1 U508 ( .A1(data_in[3]), .A2(n824), .B1(n962), .B2(\mem[26][3] ), 
        .ZN(n959) );
  INV_X1 U509 ( .A(n958), .ZN(n670) );
  AOI22_X1 U510 ( .A1(data_in[4]), .A2(n824), .B1(n962), .B2(\mem[26][4] ), 
        .ZN(n958) );
  INV_X1 U511 ( .A(n957), .ZN(n669) );
  AOI22_X1 U512 ( .A1(data_in[5]), .A2(n824), .B1(n962), .B2(\mem[26][5] ), 
        .ZN(n957) );
  INV_X1 U513 ( .A(n956), .ZN(n668) );
  AOI22_X1 U514 ( .A1(data_in[6]), .A2(n824), .B1(n962), .B2(\mem[26][6] ), 
        .ZN(n956) );
  INV_X1 U515 ( .A(n955), .ZN(n667) );
  AOI22_X1 U516 ( .A1(data_in[7]), .A2(n824), .B1(n962), .B2(\mem[26][7] ), 
        .ZN(n955) );
  INV_X1 U517 ( .A(n954), .ZN(n666) );
  AOI22_X1 U518 ( .A1(data_in[0]), .A2(n823), .B1(n953), .B2(\mem[27][0] ), 
        .ZN(n954) );
  INV_X1 U519 ( .A(n952), .ZN(n665) );
  AOI22_X1 U520 ( .A1(data_in[1]), .A2(n823), .B1(n953), .B2(\mem[27][1] ), 
        .ZN(n952) );
  INV_X1 U521 ( .A(n951), .ZN(n664) );
  AOI22_X1 U522 ( .A1(data_in[2]), .A2(n823), .B1(n953), .B2(\mem[27][2] ), 
        .ZN(n951) );
  INV_X1 U523 ( .A(n950), .ZN(n663) );
  AOI22_X1 U524 ( .A1(data_in[3]), .A2(n823), .B1(n953), .B2(\mem[27][3] ), 
        .ZN(n950) );
  INV_X1 U525 ( .A(n949), .ZN(n662) );
  AOI22_X1 U526 ( .A1(data_in[4]), .A2(n823), .B1(n953), .B2(\mem[27][4] ), 
        .ZN(n949) );
  INV_X1 U527 ( .A(n948), .ZN(n661) );
  AOI22_X1 U528 ( .A1(data_in[5]), .A2(n823), .B1(n953), .B2(\mem[27][5] ), 
        .ZN(n948) );
  INV_X1 U529 ( .A(n947), .ZN(n660) );
  AOI22_X1 U530 ( .A1(data_in[6]), .A2(n823), .B1(n953), .B2(\mem[27][6] ), 
        .ZN(n947) );
  INV_X1 U531 ( .A(n946), .ZN(n659) );
  AOI22_X1 U532 ( .A1(data_in[7]), .A2(n823), .B1(n953), .B2(\mem[27][7] ), 
        .ZN(n946) );
  INV_X1 U533 ( .A(n945), .ZN(n658) );
  AOI22_X1 U534 ( .A1(data_in[0]), .A2(n822), .B1(n944), .B2(\mem[28][0] ), 
        .ZN(n945) );
  INV_X1 U535 ( .A(n943), .ZN(n657) );
  AOI22_X1 U536 ( .A1(data_in[1]), .A2(n822), .B1(n944), .B2(\mem[28][1] ), 
        .ZN(n943) );
  INV_X1 U537 ( .A(n942), .ZN(n656) );
  AOI22_X1 U538 ( .A1(data_in[2]), .A2(n822), .B1(n944), .B2(\mem[28][2] ), 
        .ZN(n942) );
  INV_X1 U539 ( .A(n941), .ZN(n655) );
  AOI22_X1 U540 ( .A1(data_in[3]), .A2(n822), .B1(n944), .B2(\mem[28][3] ), 
        .ZN(n941) );
  INV_X1 U541 ( .A(n940), .ZN(n654) );
  AOI22_X1 U542 ( .A1(data_in[4]), .A2(n822), .B1(n944), .B2(\mem[28][4] ), 
        .ZN(n940) );
  INV_X1 U543 ( .A(n939), .ZN(n653) );
  AOI22_X1 U544 ( .A1(data_in[5]), .A2(n822), .B1(n944), .B2(\mem[28][5] ), 
        .ZN(n939) );
  INV_X1 U545 ( .A(n938), .ZN(n652) );
  AOI22_X1 U546 ( .A1(data_in[6]), .A2(n822), .B1(n944), .B2(\mem[28][6] ), 
        .ZN(n938) );
  INV_X1 U547 ( .A(n937), .ZN(n651) );
  AOI22_X1 U548 ( .A1(data_in[7]), .A2(n822), .B1(n944), .B2(\mem[28][7] ), 
        .ZN(n937) );
  INV_X1 U549 ( .A(n936), .ZN(n650) );
  AOI22_X1 U550 ( .A1(data_in[0]), .A2(n821), .B1(n935), .B2(\mem[29][0] ), 
        .ZN(n936) );
  INV_X1 U551 ( .A(n934), .ZN(n649) );
  AOI22_X1 U552 ( .A1(data_in[1]), .A2(n821), .B1(n935), .B2(\mem[29][1] ), 
        .ZN(n934) );
  INV_X1 U553 ( .A(n933), .ZN(n648) );
  AOI22_X1 U554 ( .A1(data_in[2]), .A2(n821), .B1(n935), .B2(\mem[29][2] ), 
        .ZN(n933) );
  INV_X1 U555 ( .A(n932), .ZN(n647) );
  AOI22_X1 U556 ( .A1(data_in[3]), .A2(n821), .B1(n935), .B2(\mem[29][3] ), 
        .ZN(n932) );
  INV_X1 U557 ( .A(n931), .ZN(n646) );
  AOI22_X1 U558 ( .A1(data_in[4]), .A2(n821), .B1(n935), .B2(\mem[29][4] ), 
        .ZN(n931) );
  INV_X1 U559 ( .A(n930), .ZN(n645) );
  AOI22_X1 U560 ( .A1(data_in[5]), .A2(n821), .B1(n935), .B2(\mem[29][5] ), 
        .ZN(n930) );
  INV_X1 U561 ( .A(n929), .ZN(n644) );
  AOI22_X1 U562 ( .A1(data_in[6]), .A2(n821), .B1(n935), .B2(\mem[29][6] ), 
        .ZN(n929) );
  INV_X1 U563 ( .A(n928), .ZN(n643) );
  AOI22_X1 U564 ( .A1(data_in[7]), .A2(n821), .B1(n935), .B2(\mem[29][7] ), 
        .ZN(n928) );
  INV_X1 U565 ( .A(n927), .ZN(n642) );
  AOI22_X1 U566 ( .A1(data_in[0]), .A2(n820), .B1(n926), .B2(\mem[30][0] ), 
        .ZN(n927) );
  INV_X1 U567 ( .A(n925), .ZN(n641) );
  AOI22_X1 U568 ( .A1(data_in[1]), .A2(n820), .B1(n926), .B2(\mem[30][1] ), 
        .ZN(n925) );
  INV_X1 U569 ( .A(n924), .ZN(n640) );
  AOI22_X1 U570 ( .A1(data_in[2]), .A2(n820), .B1(n926), .B2(\mem[30][2] ), 
        .ZN(n924) );
  INV_X1 U571 ( .A(n923), .ZN(n639) );
  AOI22_X1 U572 ( .A1(data_in[3]), .A2(n820), .B1(n926), .B2(\mem[30][3] ), 
        .ZN(n923) );
  INV_X1 U573 ( .A(n922), .ZN(n638) );
  AOI22_X1 U574 ( .A1(data_in[4]), .A2(n820), .B1(n926), .B2(\mem[30][4] ), 
        .ZN(n922) );
  INV_X1 U575 ( .A(n921), .ZN(n637) );
  AOI22_X1 U576 ( .A1(data_in[5]), .A2(n820), .B1(n926), .B2(\mem[30][5] ), 
        .ZN(n921) );
  INV_X1 U577 ( .A(n920), .ZN(n636) );
  AOI22_X1 U578 ( .A1(data_in[6]), .A2(n820), .B1(n926), .B2(\mem[30][6] ), 
        .ZN(n920) );
  INV_X1 U579 ( .A(n919), .ZN(n635) );
  AOI22_X1 U580 ( .A1(data_in[7]), .A2(n820), .B1(n926), .B2(\mem[30][7] ), 
        .ZN(n919) );
  INV_X1 U581 ( .A(n918), .ZN(n634) );
  AOI22_X1 U582 ( .A1(data_in[0]), .A2(n819), .B1(n917), .B2(\mem[31][0] ), 
        .ZN(n918) );
  INV_X1 U583 ( .A(n916), .ZN(n633) );
  AOI22_X1 U584 ( .A1(data_in[1]), .A2(n819), .B1(n917), .B2(\mem[31][1] ), 
        .ZN(n916) );
  INV_X1 U585 ( .A(n915), .ZN(n632) );
  AOI22_X1 U586 ( .A1(data_in[2]), .A2(n819), .B1(n917), .B2(\mem[31][2] ), 
        .ZN(n915) );
  INV_X1 U587 ( .A(n914), .ZN(n631) );
  AOI22_X1 U588 ( .A1(data_in[3]), .A2(n819), .B1(n917), .B2(\mem[31][3] ), 
        .ZN(n914) );
  INV_X1 U589 ( .A(n913), .ZN(n630) );
  AOI22_X1 U590 ( .A1(data_in[4]), .A2(n819), .B1(n917), .B2(\mem[31][4] ), 
        .ZN(n913) );
  INV_X1 U591 ( .A(n912), .ZN(n629) );
  AOI22_X1 U592 ( .A1(data_in[5]), .A2(n819), .B1(n917), .B2(\mem[31][5] ), 
        .ZN(n912) );
  INV_X1 U593 ( .A(n911), .ZN(n628) );
  AOI22_X1 U594 ( .A1(data_in[6]), .A2(n819), .B1(n917), .B2(\mem[31][6] ), 
        .ZN(n911) );
  INV_X1 U595 ( .A(n910), .ZN(n627) );
  AOI22_X1 U596 ( .A1(data_in[7]), .A2(n819), .B1(n917), .B2(\mem[31][7] ), 
        .ZN(n910) );
  MUX2_X1 U597 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n613), .Z(n1) );
  MUX2_X1 U598 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n613), .Z(n2) );
  MUX2_X1 U599 ( .A(n2), .B(n1), .S(n608), .Z(n3) );
  MUX2_X1 U600 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n613), .Z(n4) );
  MUX2_X1 U601 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n613), .Z(n5) );
  MUX2_X1 U602 ( .A(n5), .B(n4), .S(n608), .Z(n6) );
  MUX2_X1 U603 ( .A(n6), .B(n3), .S(n606), .Z(n7) );
  MUX2_X1 U604 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n613), .Z(n8) );
  MUX2_X1 U605 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n615), .Z(n9) );
  MUX2_X1 U606 ( .A(n9), .B(n8), .S(n608), .Z(n10) );
  MUX2_X1 U607 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n613), .Z(n11) );
  MUX2_X1 U608 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n614), .Z(n12) );
  MUX2_X1 U609 ( .A(n12), .B(n11), .S(n608), .Z(n13) );
  MUX2_X1 U610 ( .A(n13), .B(n10), .S(n606), .Z(n14) );
  MUX2_X1 U611 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U612 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n611), .Z(n16) );
  MUX2_X1 U613 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n611), .Z(n17) );
  MUX2_X1 U614 ( .A(n17), .B(n16), .S(n609), .Z(n18) );
  MUX2_X1 U615 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n611), .Z(n19) );
  MUX2_X1 U616 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n611), .Z(n20) );
  MUX2_X1 U617 ( .A(n20), .B(n19), .S(n609), .Z(n21) );
  MUX2_X1 U618 ( .A(n21), .B(n18), .S(n606), .Z(n22) );
  MUX2_X1 U619 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n611), .Z(n23) );
  MUX2_X1 U620 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n611), .Z(n24) );
  MUX2_X1 U621 ( .A(n24), .B(n23), .S(n609), .Z(n25) );
  MUX2_X1 U622 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n611), .Z(n26) );
  MUX2_X1 U623 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n611), .Z(n27) );
  MUX2_X1 U624 ( .A(n27), .B(n26), .S(n609), .Z(n28) );
  MUX2_X1 U625 ( .A(n28), .B(n25), .S(n606), .Z(n29) );
  MUX2_X1 U626 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U627 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U628 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n611), .Z(n31) );
  MUX2_X1 U629 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n611), .Z(n32) );
  MUX2_X1 U630 ( .A(n32), .B(n31), .S(n609), .Z(n33) );
  MUX2_X1 U631 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n611), .Z(n34) );
  MUX2_X1 U632 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n611), .Z(n35) );
  MUX2_X1 U633 ( .A(n35), .B(n34), .S(n609), .Z(n36) );
  MUX2_X1 U634 ( .A(n36), .B(n33), .S(n606), .Z(n37) );
  MUX2_X1 U635 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n612), .Z(n38) );
  MUX2_X1 U636 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n612), .Z(n39) );
  MUX2_X1 U637 ( .A(n39), .B(n38), .S(n609), .Z(n40) );
  MUX2_X1 U638 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n612), .Z(n41) );
  MUX2_X1 U639 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n612), .Z(n42) );
  MUX2_X1 U640 ( .A(n42), .B(n41), .S(n609), .Z(n43) );
  MUX2_X1 U641 ( .A(n43), .B(n40), .S(n606), .Z(n44) );
  MUX2_X1 U642 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U643 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n612), .Z(n46) );
  MUX2_X1 U644 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n612), .Z(n47) );
  MUX2_X1 U645 ( .A(n47), .B(n46), .S(n609), .Z(n48) );
  MUX2_X1 U646 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n612), .Z(n49) );
  MUX2_X1 U647 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n612), .Z(n50) );
  MUX2_X1 U648 ( .A(n50), .B(n49), .S(n609), .Z(n51) );
  MUX2_X1 U649 ( .A(n51), .B(n48), .S(n606), .Z(n52) );
  MUX2_X1 U650 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n612), .Z(n53) );
  MUX2_X1 U651 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n612), .Z(n54) );
  MUX2_X1 U652 ( .A(n54), .B(n53), .S(n609), .Z(n55) );
  MUX2_X1 U653 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n612), .Z(n56) );
  MUX2_X1 U654 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n612), .Z(n57) );
  MUX2_X1 U655 ( .A(n57), .B(n56), .S(n609), .Z(n58) );
  MUX2_X1 U656 ( .A(n58), .B(n55), .S(n606), .Z(n59) );
  MUX2_X1 U657 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U658 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U659 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n614), .Z(n61) );
  MUX2_X1 U660 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n615), .Z(n62) );
  MUX2_X1 U661 ( .A(n62), .B(n61), .S(n610), .Z(n63) );
  MUX2_X1 U662 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n612), .Z(n64) );
  MUX2_X1 U663 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n615), .Z(n65) );
  MUX2_X1 U664 ( .A(n65), .B(n64), .S(n610), .Z(n66) );
  MUX2_X1 U665 ( .A(n66), .B(n63), .S(n607), .Z(n67) );
  MUX2_X1 U666 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n614), .Z(n68) );
  MUX2_X1 U667 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n611), .Z(n69) );
  MUX2_X1 U668 ( .A(n69), .B(n68), .S(n610), .Z(n70) );
  MUX2_X1 U669 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n611), .Z(n71) );
  MUX2_X1 U670 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n615), .Z(n72) );
  MUX2_X1 U671 ( .A(n72), .B(n71), .S(n610), .Z(n73) );
  MUX2_X1 U672 ( .A(n73), .B(n70), .S(n607), .Z(n74) );
  MUX2_X1 U673 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U674 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n611), .Z(n76) );
  MUX2_X1 U675 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n612), .Z(n77) );
  MUX2_X1 U676 ( .A(n77), .B(n76), .S(n610), .Z(n78) );
  MUX2_X1 U677 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n612), .Z(n79) );
  MUX2_X1 U678 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n614), .Z(n80) );
  MUX2_X1 U679 ( .A(n80), .B(n79), .S(n610), .Z(n81) );
  MUX2_X1 U680 ( .A(n81), .B(n78), .S(n607), .Z(n82) );
  MUX2_X1 U681 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n614), .Z(n83) );
  MUX2_X1 U682 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n614), .Z(n84) );
  MUX2_X1 U683 ( .A(n84), .B(n83), .S(n610), .Z(n85) );
  MUX2_X1 U684 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n611), .Z(n86) );
  MUX2_X1 U685 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n615), .Z(n87) );
  MUX2_X1 U686 ( .A(n87), .B(n86), .S(n610), .Z(n88) );
  MUX2_X1 U687 ( .A(n88), .B(n85), .S(n607), .Z(n89) );
  MUX2_X1 U688 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U689 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U690 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n616), .Z(n91) );
  MUX2_X1 U691 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n616), .Z(n92) );
  MUX2_X1 U692 ( .A(n92), .B(n91), .S(n610), .Z(n93) );
  MUX2_X1 U693 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n616), .Z(n94) );
  MUX2_X1 U694 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n614), .Z(n95) );
  MUX2_X1 U695 ( .A(n95), .B(n94), .S(n610), .Z(n96) );
  MUX2_X1 U696 ( .A(n96), .B(n93), .S(n607), .Z(n97) );
  MUX2_X1 U697 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n616), .Z(n98) );
  MUX2_X1 U698 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n611), .Z(n99) );
  MUX2_X1 U699 ( .A(n99), .B(n98), .S(n610), .Z(n100) );
  MUX2_X1 U700 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n615), .Z(n101) );
  MUX2_X1 U701 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n612), .Z(n102) );
  MUX2_X1 U702 ( .A(n102), .B(n101), .S(n610), .Z(n103) );
  MUX2_X1 U703 ( .A(n103), .B(n100), .S(n607), .Z(n104) );
  MUX2_X1 U704 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U705 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n613), .Z(n106) );
  MUX2_X1 U706 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n613), .Z(n107) );
  MUX2_X1 U707 ( .A(n107), .B(n106), .S(n610), .Z(n108) );
  MUX2_X1 U708 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n613), .Z(n109) );
  MUX2_X1 U709 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n613), .Z(n110) );
  MUX2_X1 U710 ( .A(n110), .B(n109), .S(n609), .Z(n111) );
  MUX2_X1 U711 ( .A(n111), .B(n108), .S(n607), .Z(n112) );
  MUX2_X1 U712 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n613), .Z(n113) );
  MUX2_X1 U713 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n613), .Z(n114) );
  MUX2_X1 U714 ( .A(n114), .B(n113), .S(n608), .Z(n115) );
  MUX2_X1 U715 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n613), .Z(n116) );
  MUX2_X1 U716 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n613), .Z(n117) );
  MUX2_X1 U717 ( .A(n117), .B(n116), .S(n610), .Z(n118) );
  MUX2_X1 U718 ( .A(n118), .B(n115), .S(n607), .Z(n119) );
  MUX2_X1 U719 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U720 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U721 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n613), .Z(n121) );
  MUX2_X1 U722 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n613), .Z(n122) );
  MUX2_X1 U723 ( .A(n122), .B(n121), .S(n608), .Z(n123) );
  MUX2_X1 U724 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n613), .Z(n124) );
  MUX2_X1 U725 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n613), .Z(n125) );
  MUX2_X1 U726 ( .A(n125), .B(n124), .S(n608), .Z(n126) );
  MUX2_X1 U727 ( .A(n126), .B(n123), .S(n607), .Z(n127) );
  MUX2_X1 U728 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n614), .Z(n128) );
  MUX2_X1 U729 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n614), .Z(n129) );
  MUX2_X1 U730 ( .A(n129), .B(n128), .S(n610), .Z(n130) );
  MUX2_X1 U731 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n614), .Z(n131) );
  MUX2_X1 U732 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n614), .Z(n132) );
  MUX2_X1 U733 ( .A(n132), .B(n131), .S(n609), .Z(n133) );
  MUX2_X1 U734 ( .A(n133), .B(n130), .S(n607), .Z(n134) );
  MUX2_X1 U735 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U736 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n614), .Z(n136) );
  MUX2_X1 U737 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n614), .Z(n137) );
  MUX2_X1 U738 ( .A(n137), .B(n136), .S(n609), .Z(n138) );
  MUX2_X1 U739 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n614), .Z(n139) );
  MUX2_X1 U740 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n614), .Z(n140) );
  MUX2_X1 U741 ( .A(n140), .B(n139), .S(n608), .Z(n141) );
  MUX2_X1 U742 ( .A(n141), .B(n138), .S(n607), .Z(n142) );
  MUX2_X1 U743 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n614), .Z(n143) );
  MUX2_X1 U744 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n614), .Z(n144) );
  MUX2_X1 U745 ( .A(n144), .B(n143), .S(n609), .Z(n145) );
  MUX2_X1 U746 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n614), .Z(n146) );
  MUX2_X1 U747 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n614), .Z(n147) );
  MUX2_X1 U748 ( .A(n147), .B(n146), .S(n608), .Z(n148) );
  MUX2_X1 U749 ( .A(n148), .B(n145), .S(n607), .Z(n149) );
  MUX2_X1 U750 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U751 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U752 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n615), .Z(n151) );
  MUX2_X1 U753 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n615), .Z(n152) );
  MUX2_X1 U754 ( .A(n152), .B(n151), .S(n609), .Z(n153) );
  MUX2_X1 U755 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n615), .Z(n154) );
  MUX2_X1 U756 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n615), .Z(n155) );
  MUX2_X1 U757 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U758 ( .A(n156), .B(n153), .S(n606), .Z(n157) );
  MUX2_X1 U759 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n615), .Z(n158) );
  MUX2_X1 U760 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n615), .Z(n159) );
  MUX2_X1 U761 ( .A(n159), .B(n158), .S(n608), .Z(n160) );
  MUX2_X1 U762 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n615), .Z(n161) );
  MUX2_X1 U763 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n615), .Z(n162) );
  MUX2_X1 U764 ( .A(n162), .B(n161), .S(N11), .Z(n163) );
  MUX2_X1 U765 ( .A(n163), .B(n160), .S(n606), .Z(n164) );
  MUX2_X1 U766 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U767 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n615), .Z(n166) );
  MUX2_X1 U768 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n615), .Z(n167) );
  MUX2_X1 U769 ( .A(n167), .B(n166), .S(n610), .Z(n168) );
  MUX2_X1 U770 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n615), .Z(n169) );
  MUX2_X1 U771 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n615), .Z(n170) );
  MUX2_X1 U772 ( .A(n170), .B(n169), .S(n610), .Z(n171) );
  MUX2_X1 U773 ( .A(n171), .B(n168), .S(n606), .Z(n172) );
  MUX2_X1 U774 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n616), .Z(n173) );
  MUX2_X1 U775 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n615), .Z(n174) );
  MUX2_X1 U776 ( .A(n174), .B(n173), .S(n610), .Z(n175) );
  MUX2_X1 U777 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n616), .Z(n176) );
  MUX2_X1 U778 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n616), .Z(n177) );
  MUX2_X1 U779 ( .A(n177), .B(n176), .S(n609), .Z(n178) );
  MUX2_X1 U780 ( .A(n178), .B(n175), .S(n607), .Z(n179) );
  MUX2_X1 U781 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U782 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U783 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n616), .Z(n181) );
  MUX2_X1 U784 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n612), .Z(n182) );
  MUX2_X1 U785 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U786 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n615), .Z(n184) );
  MUX2_X1 U787 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n616), .Z(n185) );
  MUX2_X1 U788 ( .A(n185), .B(n184), .S(n609), .Z(n186) );
  MUX2_X1 U789 ( .A(n186), .B(n183), .S(n606), .Z(n187) );
  MUX2_X1 U790 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n616), .Z(n188) );
  MUX2_X1 U791 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n611), .Z(n189) );
  MUX2_X1 U792 ( .A(n189), .B(n188), .S(N11), .Z(n190) );
  MUX2_X1 U793 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n616), .Z(n191) );
  MUX2_X1 U794 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n614), .Z(n192) );
  MUX2_X1 U795 ( .A(n192), .B(n191), .S(n609), .Z(n193) );
  MUX2_X1 U796 ( .A(n193), .B(n190), .S(n607), .Z(n194) );
  MUX2_X1 U797 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U798 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n611), .Z(n196) );
  MUX2_X1 U799 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n616), .Z(n197) );
  MUX2_X1 U800 ( .A(n197), .B(n196), .S(n608), .Z(n198) );
  MUX2_X1 U801 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n616), .Z(n199) );
  MUX2_X1 U802 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n616), .Z(n200) );
  MUX2_X1 U803 ( .A(n200), .B(n199), .S(n609), .Z(n201) );
  MUX2_X1 U804 ( .A(n201), .B(n198), .S(n606), .Z(n202) );
  MUX2_X1 U805 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n612), .Z(n203) );
  MUX2_X1 U806 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n616), .Z(n204) );
  MUX2_X1 U807 ( .A(n204), .B(n203), .S(n608), .Z(n205) );
  MUX2_X1 U808 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n616), .Z(n206) );
  MUX2_X1 U809 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n207) );
  MUX2_X1 U810 ( .A(n207), .B(n206), .S(n610), .Z(n208) );
  MUX2_X1 U811 ( .A(n208), .B(n205), .S(n606), .Z(n209) );
  MUX2_X1 U812 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U813 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U814 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n612), .Z(n211) );
  MUX2_X1 U815 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n612), .Z(n212) );
  MUX2_X1 U816 ( .A(n212), .B(n211), .S(n608), .Z(n213) );
  MUX2_X1 U817 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n611), .Z(n214) );
  MUX2_X1 U818 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n613), .Z(n215) );
  MUX2_X1 U819 ( .A(n215), .B(n214), .S(n608), .Z(n216) );
  MUX2_X1 U820 ( .A(n216), .B(n213), .S(n606), .Z(n217) );
  MUX2_X1 U821 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n613), .Z(n218) );
  MUX2_X1 U822 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n616), .Z(n219) );
  MUX2_X1 U823 ( .A(n219), .B(n218), .S(n608), .Z(n220) );
  MUX2_X1 U824 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(N10), .Z(n221) );
  MUX2_X1 U825 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n222) );
  MUX2_X1 U826 ( .A(n222), .B(n221), .S(n610), .Z(n223) );
  MUX2_X1 U827 ( .A(n223), .B(n220), .S(n606), .Z(n224) );
  MUX2_X1 U828 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U829 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n613), .Z(n226) );
  MUX2_X1 U830 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n613), .Z(n227) );
  MUX2_X1 U831 ( .A(n227), .B(n226), .S(n608), .Z(n228) );
  MUX2_X1 U832 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(N10), .Z(n229) );
  MUX2_X1 U833 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n595) );
  MUX2_X1 U834 ( .A(n595), .B(n229), .S(N11), .Z(n596) );
  MUX2_X1 U835 ( .A(n596), .B(n228), .S(n607), .Z(n597) );
  MUX2_X1 U836 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n613), .Z(n598) );
  MUX2_X1 U837 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n616), .Z(n599) );
  MUX2_X1 U838 ( .A(n599), .B(n598), .S(n608), .Z(n600) );
  MUX2_X1 U839 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n616), .Z(n601) );
  MUX2_X1 U840 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n616), .Z(n602) );
  MUX2_X1 U841 ( .A(n602), .B(n601), .S(n608), .Z(n603) );
  MUX2_X1 U842 ( .A(n603), .B(n600), .S(n607), .Z(n604) );
  MUX2_X1 U843 ( .A(n604), .B(n597), .S(N13), .Z(n605) );
  MUX2_X1 U844 ( .A(n605), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U845 ( .A(N11), .Z(n608) );
  INV_X1 U846 ( .A(N10), .ZN(n617) );
  INV_X1 U847 ( .A(N11), .ZN(n618) );
  INV_X1 U848 ( .A(data_in[0]), .ZN(n619) );
  INV_X1 U849 ( .A(data_in[1]), .ZN(n620) );
  INV_X1 U850 ( .A(data_in[2]), .ZN(n621) );
  INV_X1 U851 ( .A(data_in[3]), .ZN(n622) );
  INV_X1 U852 ( .A(data_in[4]), .ZN(n623) );
  INV_X1 U853 ( .A(data_in[5]), .ZN(n624) );
  INV_X1 U854 ( .A(data_in[6]), .ZN(n625) );
  INV_X1 U855 ( .A(data_in[7]), .ZN(n626) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_25 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n630), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n631), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n632), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n633), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n634), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n635), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n636), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n637), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n638), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n639), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n640), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n641), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n642), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n643), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n644), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n645), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n646), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n647), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n648), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n649), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n650), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n651), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n652), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n653), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n654), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n655), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n656), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n657), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n658), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n659), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n660), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n661), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n662), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n663), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n664), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n665), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n666), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n667), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n668), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n669), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n670), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n671), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n672), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n673), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n674), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n675), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n676), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n677), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n678), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n679), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n680), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n681), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n682), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n683), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n684), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n685), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n686), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n687), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n688), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n689), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n690), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n691), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n692), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n693), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n694), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n695), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n696), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n697), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n698), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n699), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n700), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n701), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n702), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n703), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n704), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n705), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n706), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n707), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n708), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n709), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n710), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n711), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n712), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n713), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n714), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n715), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n716), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n717), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n718), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n719), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n720), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n721), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n722), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n723), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n724), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n725), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n726), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n727), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n728), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n729), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n730), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n731), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n732), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n733), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n734), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n735), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n736), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n737), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n738), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n739), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n740), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n741), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n742), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n743), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n744), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n745), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n746), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n747), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n748), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n749), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n750), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n751), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n752), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n753), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n754), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n755), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n756), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n757), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n758), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n759), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n760), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n761), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n762), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n763), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n764), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n765), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n766), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n767), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n768), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n769), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n770), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n771), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n772), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n773), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n774), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n775), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n776), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n777), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n778), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n779), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n780), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n781), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n782), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n783), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n784), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n785), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n786), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n787), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n788), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n789), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n790), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n791), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n792), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n793), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n794), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n795), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n796), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n797), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n798), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n799), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n800), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n801), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n802), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n803), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n804), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n805), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n806), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n807), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n808), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n809), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n810), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n811), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n812), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n813), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n814), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n815), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n816), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n817), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n818), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n819), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n820), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n821), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n849), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n850), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n851), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n852), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n853), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n854), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n855), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n856), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n857), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n858), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n859), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n860), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n861), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n862), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n863), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n864), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n865), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n866), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n867), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n868), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n869), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n870), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n871), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n872), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n873), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n874), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n875), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n876), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n877), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n878), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n879), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n880), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n881), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n882), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n883), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n884), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n885), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n886), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n887), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n888), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n889), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n890), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n891), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n892), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n893), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n894), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n895), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n896), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n897), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n898), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n899), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n900), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n901), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n902), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n903), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n904), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n905), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n906), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n907), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n908), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n909), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n910), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n911), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n912), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X2 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  BUF_X1 U3 ( .A(n619), .Z(n612) );
  BUF_X1 U4 ( .A(N10), .Z(n617) );
  BUF_X1 U5 ( .A(n619), .Z(n618) );
  BUF_X1 U6 ( .A(N10), .Z(n614) );
  BUF_X1 U7 ( .A(n619), .Z(n615) );
  BUF_X1 U8 ( .A(n619), .Z(n616) );
  BUF_X1 U9 ( .A(n619), .Z(n613) );
  BUF_X1 U10 ( .A(N11), .Z(n610) );
  BUF_X1 U11 ( .A(N11), .Z(n611) );
  BUF_X1 U12 ( .A(N10), .Z(n619) );
  NOR3_X1 U13 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1204) );
  NOR3_X1 U14 ( .A1(N11), .A2(N12), .A3(n620), .ZN(n1193) );
  NOR3_X1 U15 ( .A1(N10), .A2(N12), .A3(n621), .ZN(n1183) );
  NOR3_X1 U16 ( .A1(n620), .A2(N12), .A3(n621), .ZN(n1173) );
  INV_X1 U17 ( .A(n1130), .ZN(n845) );
  INV_X1 U18 ( .A(n1120), .ZN(n844) );
  INV_X1 U19 ( .A(n1111), .ZN(n843) );
  INV_X1 U20 ( .A(n1102), .ZN(n842) );
  INV_X1 U21 ( .A(n1057), .ZN(n837) );
  INV_X1 U22 ( .A(n1047), .ZN(n836) );
  INV_X1 U23 ( .A(n1038), .ZN(n835) );
  INV_X1 U24 ( .A(n1029), .ZN(n834) );
  INV_X1 U25 ( .A(n984), .ZN(n829) );
  INV_X1 U26 ( .A(n974), .ZN(n828) );
  INV_X1 U27 ( .A(n965), .ZN(n827) );
  INV_X1 U28 ( .A(n956), .ZN(n826) );
  INV_X1 U29 ( .A(n920), .ZN(n822) );
  INV_X1 U30 ( .A(n1093), .ZN(n841) );
  INV_X1 U31 ( .A(n1084), .ZN(n840) );
  INV_X1 U32 ( .A(n1075), .ZN(n839) );
  INV_X1 U33 ( .A(n1066), .ZN(n838) );
  INV_X1 U34 ( .A(n947), .ZN(n825) );
  INV_X1 U35 ( .A(n938), .ZN(n824) );
  INV_X1 U36 ( .A(n929), .ZN(n823) );
  INV_X1 U37 ( .A(n1020), .ZN(n833) );
  INV_X1 U38 ( .A(n1011), .ZN(n832) );
  INV_X1 U39 ( .A(n1002), .ZN(n831) );
  INV_X1 U40 ( .A(n993), .ZN(n830) );
  BUF_X1 U41 ( .A(N12), .Z(n607) );
  BUF_X1 U42 ( .A(N12), .Z(n608) );
  INV_X1 U43 ( .A(N13), .ZN(n847) );
  AND3_X1 U44 ( .A1(n620), .A2(n621), .A3(N12), .ZN(n1163) );
  AND3_X1 U45 ( .A1(N10), .A2(n621), .A3(N12), .ZN(n1153) );
  AND3_X1 U46 ( .A1(N11), .A2(n620), .A3(N12), .ZN(n1143) );
  AND3_X1 U47 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1133) );
  INV_X1 U48 ( .A(N14), .ZN(n848) );
  NAND2_X1 U49 ( .A1(n1193), .A2(n1203), .ZN(n1202) );
  NAND2_X1 U50 ( .A1(n1183), .A2(n1203), .ZN(n1192) );
  NAND2_X1 U51 ( .A1(n1173), .A2(n1203), .ZN(n1182) );
  NAND2_X1 U52 ( .A1(n1163), .A2(n1203), .ZN(n1172) );
  NAND2_X1 U53 ( .A1(n1153), .A2(n1203), .ZN(n1162) );
  NAND2_X1 U54 ( .A1(n1143), .A2(n1203), .ZN(n1152) );
  NAND2_X1 U55 ( .A1(n1133), .A2(n1203), .ZN(n1142) );
  NAND2_X1 U56 ( .A1(n1204), .A2(n1203), .ZN(n1213) );
  NAND2_X1 U57 ( .A1(n1122), .A2(n1204), .ZN(n1130) );
  NAND2_X1 U58 ( .A1(n1122), .A2(n1193), .ZN(n1120) );
  NAND2_X1 U59 ( .A1(n1122), .A2(n1183), .ZN(n1111) );
  NAND2_X1 U60 ( .A1(n1122), .A2(n1173), .ZN(n1102) );
  NAND2_X1 U61 ( .A1(n1049), .A2(n1204), .ZN(n1057) );
  NAND2_X1 U62 ( .A1(n1049), .A2(n1193), .ZN(n1047) );
  NAND2_X1 U63 ( .A1(n1049), .A2(n1183), .ZN(n1038) );
  NAND2_X1 U64 ( .A1(n1049), .A2(n1173), .ZN(n1029) );
  NAND2_X1 U65 ( .A1(n976), .A2(n1204), .ZN(n984) );
  NAND2_X1 U66 ( .A1(n976), .A2(n1193), .ZN(n974) );
  NAND2_X1 U67 ( .A1(n976), .A2(n1183), .ZN(n965) );
  NAND2_X1 U68 ( .A1(n976), .A2(n1173), .ZN(n956) );
  NAND2_X1 U69 ( .A1(n1122), .A2(n1163), .ZN(n1093) );
  NAND2_X1 U70 ( .A1(n1122), .A2(n1153), .ZN(n1084) );
  NAND2_X1 U71 ( .A1(n1122), .A2(n1143), .ZN(n1075) );
  NAND2_X1 U72 ( .A1(n1122), .A2(n1133), .ZN(n1066) );
  NAND2_X1 U73 ( .A1(n1049), .A2(n1163), .ZN(n1020) );
  NAND2_X1 U74 ( .A1(n1049), .A2(n1153), .ZN(n1011) );
  NAND2_X1 U75 ( .A1(n1049), .A2(n1143), .ZN(n1002) );
  NAND2_X1 U76 ( .A1(n1049), .A2(n1133), .ZN(n993) );
  NAND2_X1 U77 ( .A1(n976), .A2(n1163), .ZN(n947) );
  NAND2_X1 U78 ( .A1(n976), .A2(n1153), .ZN(n938) );
  NAND2_X1 U79 ( .A1(n976), .A2(n1143), .ZN(n929) );
  NAND2_X1 U80 ( .A1(n976), .A2(n1133), .ZN(n920) );
  AND3_X1 U81 ( .A1(n847), .A2(n848), .A3(n1132), .ZN(n1203) );
  AND3_X1 U82 ( .A1(N13), .A2(n1132), .A3(N14), .ZN(n976) );
  AND3_X1 U83 ( .A1(n1132), .A2(n848), .A3(N13), .ZN(n1122) );
  AND3_X1 U84 ( .A1(n1132), .A2(n847), .A3(N14), .ZN(n1049) );
  NOR2_X1 U85 ( .A1(n846), .A2(addr[5]), .ZN(n1132) );
  INV_X1 U86 ( .A(wr_en), .ZN(n846) );
  OAI21_X1 U87 ( .B1(n622), .B2(n1172), .A(n1171), .ZN(n880) );
  NAND2_X1 U88 ( .A1(\mem[4][0] ), .A2(n1172), .ZN(n1171) );
  OAI21_X1 U89 ( .B1(n623), .B2(n1172), .A(n1170), .ZN(n879) );
  NAND2_X1 U90 ( .A1(\mem[4][1] ), .A2(n1172), .ZN(n1170) );
  OAI21_X1 U91 ( .B1(n624), .B2(n1172), .A(n1169), .ZN(n878) );
  NAND2_X1 U92 ( .A1(\mem[4][2] ), .A2(n1172), .ZN(n1169) );
  OAI21_X1 U93 ( .B1(n625), .B2(n1172), .A(n1168), .ZN(n877) );
  NAND2_X1 U94 ( .A1(\mem[4][3] ), .A2(n1172), .ZN(n1168) );
  OAI21_X1 U95 ( .B1(n626), .B2(n1172), .A(n1167), .ZN(n876) );
  NAND2_X1 U96 ( .A1(\mem[4][4] ), .A2(n1172), .ZN(n1167) );
  OAI21_X1 U97 ( .B1(n627), .B2(n1172), .A(n1166), .ZN(n875) );
  NAND2_X1 U98 ( .A1(\mem[4][5] ), .A2(n1172), .ZN(n1166) );
  OAI21_X1 U99 ( .B1(n628), .B2(n1172), .A(n1165), .ZN(n874) );
  NAND2_X1 U100 ( .A1(\mem[4][6] ), .A2(n1172), .ZN(n1165) );
  OAI21_X1 U101 ( .B1(n629), .B2(n1172), .A(n1164), .ZN(n873) );
  NAND2_X1 U102 ( .A1(\mem[4][7] ), .A2(n1172), .ZN(n1164) );
  OAI21_X1 U103 ( .B1(n622), .B2(n1152), .A(n1151), .ZN(n864) );
  NAND2_X1 U104 ( .A1(\mem[6][0] ), .A2(n1152), .ZN(n1151) );
  OAI21_X1 U105 ( .B1(n623), .B2(n1152), .A(n1150), .ZN(n863) );
  NAND2_X1 U106 ( .A1(\mem[6][1] ), .A2(n1152), .ZN(n1150) );
  OAI21_X1 U107 ( .B1(n624), .B2(n1152), .A(n1149), .ZN(n862) );
  NAND2_X1 U108 ( .A1(\mem[6][2] ), .A2(n1152), .ZN(n1149) );
  OAI21_X1 U109 ( .B1(n625), .B2(n1152), .A(n1148), .ZN(n861) );
  NAND2_X1 U110 ( .A1(\mem[6][3] ), .A2(n1152), .ZN(n1148) );
  OAI21_X1 U111 ( .B1(n626), .B2(n1152), .A(n1147), .ZN(n860) );
  NAND2_X1 U112 ( .A1(\mem[6][4] ), .A2(n1152), .ZN(n1147) );
  OAI21_X1 U113 ( .B1(n627), .B2(n1152), .A(n1146), .ZN(n859) );
  NAND2_X1 U114 ( .A1(\mem[6][5] ), .A2(n1152), .ZN(n1146) );
  OAI21_X1 U115 ( .B1(n628), .B2(n1152), .A(n1145), .ZN(n858) );
  NAND2_X1 U116 ( .A1(\mem[6][6] ), .A2(n1152), .ZN(n1145) );
  OAI21_X1 U117 ( .B1(n629), .B2(n1152), .A(n1144), .ZN(n857) );
  NAND2_X1 U118 ( .A1(\mem[6][7] ), .A2(n1152), .ZN(n1144) );
  OAI21_X1 U119 ( .B1(n622), .B2(n1142), .A(n1141), .ZN(n856) );
  NAND2_X1 U120 ( .A1(\mem[7][0] ), .A2(n1142), .ZN(n1141) );
  OAI21_X1 U121 ( .B1(n623), .B2(n1142), .A(n1140), .ZN(n855) );
  NAND2_X1 U122 ( .A1(\mem[7][1] ), .A2(n1142), .ZN(n1140) );
  OAI21_X1 U123 ( .B1(n624), .B2(n1142), .A(n1139), .ZN(n854) );
  NAND2_X1 U124 ( .A1(\mem[7][2] ), .A2(n1142), .ZN(n1139) );
  OAI21_X1 U125 ( .B1(n625), .B2(n1142), .A(n1138), .ZN(n853) );
  NAND2_X1 U126 ( .A1(\mem[7][3] ), .A2(n1142), .ZN(n1138) );
  OAI21_X1 U127 ( .B1(n626), .B2(n1142), .A(n1137), .ZN(n852) );
  NAND2_X1 U128 ( .A1(\mem[7][4] ), .A2(n1142), .ZN(n1137) );
  OAI21_X1 U129 ( .B1(n627), .B2(n1142), .A(n1136), .ZN(n851) );
  NAND2_X1 U130 ( .A1(\mem[7][5] ), .A2(n1142), .ZN(n1136) );
  OAI21_X1 U131 ( .B1(n628), .B2(n1142), .A(n1135), .ZN(n850) );
  NAND2_X1 U132 ( .A1(\mem[7][6] ), .A2(n1142), .ZN(n1135) );
  OAI21_X1 U133 ( .B1(n629), .B2(n1142), .A(n1134), .ZN(n849) );
  NAND2_X1 U134 ( .A1(\mem[7][7] ), .A2(n1142), .ZN(n1134) );
  OAI21_X1 U135 ( .B1(n622), .B2(n1202), .A(n1201), .ZN(n904) );
  NAND2_X1 U136 ( .A1(\mem[1][0] ), .A2(n1202), .ZN(n1201) );
  OAI21_X1 U137 ( .B1(n623), .B2(n1202), .A(n1200), .ZN(n903) );
  NAND2_X1 U138 ( .A1(\mem[1][1] ), .A2(n1202), .ZN(n1200) );
  OAI21_X1 U139 ( .B1(n624), .B2(n1202), .A(n1199), .ZN(n902) );
  NAND2_X1 U140 ( .A1(\mem[1][2] ), .A2(n1202), .ZN(n1199) );
  OAI21_X1 U141 ( .B1(n625), .B2(n1202), .A(n1198), .ZN(n901) );
  NAND2_X1 U142 ( .A1(\mem[1][3] ), .A2(n1202), .ZN(n1198) );
  OAI21_X1 U143 ( .B1(n626), .B2(n1202), .A(n1197), .ZN(n900) );
  NAND2_X1 U144 ( .A1(\mem[1][4] ), .A2(n1202), .ZN(n1197) );
  OAI21_X1 U145 ( .B1(n627), .B2(n1202), .A(n1196), .ZN(n899) );
  NAND2_X1 U146 ( .A1(\mem[1][5] ), .A2(n1202), .ZN(n1196) );
  OAI21_X1 U147 ( .B1(n628), .B2(n1202), .A(n1195), .ZN(n898) );
  NAND2_X1 U148 ( .A1(\mem[1][6] ), .A2(n1202), .ZN(n1195) );
  OAI21_X1 U149 ( .B1(n629), .B2(n1202), .A(n1194), .ZN(n897) );
  NAND2_X1 U150 ( .A1(\mem[1][7] ), .A2(n1202), .ZN(n1194) );
  OAI21_X1 U151 ( .B1(n622), .B2(n1192), .A(n1191), .ZN(n896) );
  NAND2_X1 U152 ( .A1(\mem[2][0] ), .A2(n1192), .ZN(n1191) );
  OAI21_X1 U153 ( .B1(n623), .B2(n1192), .A(n1190), .ZN(n895) );
  NAND2_X1 U154 ( .A1(\mem[2][1] ), .A2(n1192), .ZN(n1190) );
  OAI21_X1 U155 ( .B1(n624), .B2(n1192), .A(n1189), .ZN(n894) );
  NAND2_X1 U156 ( .A1(\mem[2][2] ), .A2(n1192), .ZN(n1189) );
  OAI21_X1 U157 ( .B1(n625), .B2(n1192), .A(n1188), .ZN(n893) );
  NAND2_X1 U158 ( .A1(\mem[2][3] ), .A2(n1192), .ZN(n1188) );
  OAI21_X1 U159 ( .B1(n626), .B2(n1192), .A(n1187), .ZN(n892) );
  NAND2_X1 U160 ( .A1(\mem[2][4] ), .A2(n1192), .ZN(n1187) );
  OAI21_X1 U161 ( .B1(n627), .B2(n1192), .A(n1186), .ZN(n891) );
  NAND2_X1 U162 ( .A1(\mem[2][5] ), .A2(n1192), .ZN(n1186) );
  OAI21_X1 U163 ( .B1(n628), .B2(n1192), .A(n1185), .ZN(n890) );
  NAND2_X1 U164 ( .A1(\mem[2][6] ), .A2(n1192), .ZN(n1185) );
  OAI21_X1 U165 ( .B1(n629), .B2(n1192), .A(n1184), .ZN(n889) );
  NAND2_X1 U166 ( .A1(\mem[2][7] ), .A2(n1192), .ZN(n1184) );
  OAI21_X1 U167 ( .B1(n622), .B2(n1182), .A(n1181), .ZN(n888) );
  NAND2_X1 U168 ( .A1(\mem[3][0] ), .A2(n1182), .ZN(n1181) );
  OAI21_X1 U169 ( .B1(n623), .B2(n1182), .A(n1180), .ZN(n887) );
  NAND2_X1 U170 ( .A1(\mem[3][1] ), .A2(n1182), .ZN(n1180) );
  OAI21_X1 U171 ( .B1(n624), .B2(n1182), .A(n1179), .ZN(n886) );
  NAND2_X1 U172 ( .A1(\mem[3][2] ), .A2(n1182), .ZN(n1179) );
  OAI21_X1 U173 ( .B1(n625), .B2(n1182), .A(n1178), .ZN(n885) );
  NAND2_X1 U174 ( .A1(\mem[3][3] ), .A2(n1182), .ZN(n1178) );
  OAI21_X1 U175 ( .B1(n626), .B2(n1182), .A(n1177), .ZN(n884) );
  NAND2_X1 U176 ( .A1(\mem[3][4] ), .A2(n1182), .ZN(n1177) );
  OAI21_X1 U177 ( .B1(n627), .B2(n1182), .A(n1176), .ZN(n883) );
  NAND2_X1 U178 ( .A1(\mem[3][5] ), .A2(n1182), .ZN(n1176) );
  OAI21_X1 U179 ( .B1(n628), .B2(n1182), .A(n1175), .ZN(n882) );
  NAND2_X1 U180 ( .A1(\mem[3][6] ), .A2(n1182), .ZN(n1175) );
  OAI21_X1 U181 ( .B1(n629), .B2(n1182), .A(n1174), .ZN(n881) );
  NAND2_X1 U182 ( .A1(\mem[3][7] ), .A2(n1182), .ZN(n1174) );
  OAI21_X1 U183 ( .B1(n622), .B2(n1162), .A(n1161), .ZN(n872) );
  NAND2_X1 U184 ( .A1(\mem[5][0] ), .A2(n1162), .ZN(n1161) );
  OAI21_X1 U185 ( .B1(n623), .B2(n1162), .A(n1160), .ZN(n871) );
  NAND2_X1 U186 ( .A1(\mem[5][1] ), .A2(n1162), .ZN(n1160) );
  OAI21_X1 U187 ( .B1(n624), .B2(n1162), .A(n1159), .ZN(n870) );
  NAND2_X1 U188 ( .A1(\mem[5][2] ), .A2(n1162), .ZN(n1159) );
  OAI21_X1 U189 ( .B1(n625), .B2(n1162), .A(n1158), .ZN(n869) );
  NAND2_X1 U190 ( .A1(\mem[5][3] ), .A2(n1162), .ZN(n1158) );
  OAI21_X1 U191 ( .B1(n626), .B2(n1162), .A(n1157), .ZN(n868) );
  NAND2_X1 U192 ( .A1(\mem[5][4] ), .A2(n1162), .ZN(n1157) );
  OAI21_X1 U193 ( .B1(n627), .B2(n1162), .A(n1156), .ZN(n867) );
  NAND2_X1 U194 ( .A1(\mem[5][5] ), .A2(n1162), .ZN(n1156) );
  OAI21_X1 U195 ( .B1(n628), .B2(n1162), .A(n1155), .ZN(n866) );
  NAND2_X1 U196 ( .A1(\mem[5][6] ), .A2(n1162), .ZN(n1155) );
  OAI21_X1 U197 ( .B1(n629), .B2(n1162), .A(n1154), .ZN(n865) );
  NAND2_X1 U198 ( .A1(\mem[5][7] ), .A2(n1162), .ZN(n1154) );
  OAI21_X1 U199 ( .B1(n1213), .B2(n622), .A(n1212), .ZN(n912) );
  NAND2_X1 U200 ( .A1(\mem[0][0] ), .A2(n1213), .ZN(n1212) );
  OAI21_X1 U201 ( .B1(n1213), .B2(n623), .A(n1211), .ZN(n911) );
  NAND2_X1 U202 ( .A1(\mem[0][1] ), .A2(n1213), .ZN(n1211) );
  OAI21_X1 U203 ( .B1(n1213), .B2(n624), .A(n1210), .ZN(n910) );
  NAND2_X1 U204 ( .A1(\mem[0][2] ), .A2(n1213), .ZN(n1210) );
  OAI21_X1 U205 ( .B1(n1213), .B2(n625), .A(n1209), .ZN(n909) );
  NAND2_X1 U206 ( .A1(\mem[0][3] ), .A2(n1213), .ZN(n1209) );
  OAI21_X1 U207 ( .B1(n1213), .B2(n626), .A(n1208), .ZN(n908) );
  NAND2_X1 U208 ( .A1(\mem[0][4] ), .A2(n1213), .ZN(n1208) );
  OAI21_X1 U209 ( .B1(n1213), .B2(n627), .A(n1207), .ZN(n907) );
  NAND2_X1 U210 ( .A1(\mem[0][5] ), .A2(n1213), .ZN(n1207) );
  OAI21_X1 U211 ( .B1(n1213), .B2(n628), .A(n1206), .ZN(n906) );
  NAND2_X1 U212 ( .A1(\mem[0][6] ), .A2(n1213), .ZN(n1206) );
  OAI21_X1 U213 ( .B1(n1213), .B2(n629), .A(n1205), .ZN(n905) );
  NAND2_X1 U214 ( .A1(\mem[0][7] ), .A2(n1213), .ZN(n1205) );
  INV_X1 U215 ( .A(n1131), .ZN(n821) );
  AOI22_X1 U216 ( .A1(data_in[0]), .A2(n845), .B1(n1130), .B2(\mem[8][0] ), 
        .ZN(n1131) );
  INV_X1 U217 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U218 ( .A1(data_in[1]), .A2(n845), .B1(n1130), .B2(\mem[8][1] ), 
        .ZN(n1129) );
  INV_X1 U219 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U220 ( .A1(data_in[2]), .A2(n845), .B1(n1130), .B2(\mem[8][2] ), 
        .ZN(n1128) );
  INV_X1 U221 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U222 ( .A1(data_in[3]), .A2(n845), .B1(n1130), .B2(\mem[8][3] ), 
        .ZN(n1127) );
  INV_X1 U223 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U224 ( .A1(data_in[4]), .A2(n845), .B1(n1130), .B2(\mem[8][4] ), 
        .ZN(n1126) );
  INV_X1 U225 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U226 ( .A1(data_in[5]), .A2(n845), .B1(n1130), .B2(\mem[8][5] ), 
        .ZN(n1125) );
  INV_X1 U227 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U228 ( .A1(data_in[6]), .A2(n845), .B1(n1130), .B2(\mem[8][6] ), 
        .ZN(n1124) );
  INV_X1 U229 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U230 ( .A1(data_in[7]), .A2(n845), .B1(n1130), .B2(\mem[8][7] ), 
        .ZN(n1123) );
  INV_X1 U231 ( .A(n1121), .ZN(n813) );
  AOI22_X1 U232 ( .A1(data_in[0]), .A2(n844), .B1(n1120), .B2(\mem[9][0] ), 
        .ZN(n1121) );
  INV_X1 U233 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U234 ( .A1(data_in[1]), .A2(n844), .B1(n1120), .B2(\mem[9][1] ), 
        .ZN(n1119) );
  INV_X1 U235 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U236 ( .A1(data_in[2]), .A2(n844), .B1(n1120), .B2(\mem[9][2] ), 
        .ZN(n1118) );
  INV_X1 U237 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U238 ( .A1(data_in[3]), .A2(n844), .B1(n1120), .B2(\mem[9][3] ), 
        .ZN(n1117) );
  INV_X1 U239 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U240 ( .A1(data_in[4]), .A2(n844), .B1(n1120), .B2(\mem[9][4] ), 
        .ZN(n1116) );
  INV_X1 U241 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U242 ( .A1(data_in[5]), .A2(n844), .B1(n1120), .B2(\mem[9][5] ), 
        .ZN(n1115) );
  INV_X1 U243 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U244 ( .A1(data_in[6]), .A2(n844), .B1(n1120), .B2(\mem[9][6] ), 
        .ZN(n1114) );
  INV_X1 U245 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U246 ( .A1(data_in[7]), .A2(n844), .B1(n1120), .B2(\mem[9][7] ), 
        .ZN(n1113) );
  INV_X1 U247 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U248 ( .A1(data_in[0]), .A2(n843), .B1(n1111), .B2(\mem[10][0] ), 
        .ZN(n1112) );
  INV_X1 U249 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U250 ( .A1(data_in[1]), .A2(n843), .B1(n1111), .B2(\mem[10][1] ), 
        .ZN(n1110) );
  INV_X1 U251 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U252 ( .A1(data_in[2]), .A2(n843), .B1(n1111), .B2(\mem[10][2] ), 
        .ZN(n1109) );
  INV_X1 U253 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U254 ( .A1(data_in[3]), .A2(n843), .B1(n1111), .B2(\mem[10][3] ), 
        .ZN(n1108) );
  INV_X1 U255 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U256 ( .A1(data_in[4]), .A2(n843), .B1(n1111), .B2(\mem[10][4] ), 
        .ZN(n1107) );
  INV_X1 U257 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U258 ( .A1(data_in[5]), .A2(n843), .B1(n1111), .B2(\mem[10][5] ), 
        .ZN(n1106) );
  INV_X1 U259 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U260 ( .A1(data_in[6]), .A2(n843), .B1(n1111), .B2(\mem[10][6] ), 
        .ZN(n1105) );
  INV_X1 U261 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U262 ( .A1(data_in[7]), .A2(n843), .B1(n1111), .B2(\mem[10][7] ), 
        .ZN(n1104) );
  INV_X1 U263 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U264 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[11][0] ), 
        .ZN(n1103) );
  INV_X1 U265 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U266 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[11][1] ), 
        .ZN(n1101) );
  INV_X1 U267 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U268 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[11][2] ), 
        .ZN(n1100) );
  INV_X1 U269 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U270 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[11][3] ), 
        .ZN(n1099) );
  INV_X1 U271 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U272 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[11][4] ), 
        .ZN(n1098) );
  INV_X1 U273 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U274 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[11][5] ), 
        .ZN(n1097) );
  INV_X1 U275 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U276 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[11][6] ), 
        .ZN(n1096) );
  INV_X1 U277 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U278 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[11][7] ), 
        .ZN(n1095) );
  INV_X1 U279 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U280 ( .A1(data_in[0]), .A2(n841), .B1(n1093), .B2(\mem[12][0] ), 
        .ZN(n1094) );
  INV_X1 U281 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U282 ( .A1(data_in[1]), .A2(n841), .B1(n1093), .B2(\mem[12][1] ), 
        .ZN(n1092) );
  INV_X1 U283 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U284 ( .A1(data_in[2]), .A2(n841), .B1(n1093), .B2(\mem[12][2] ), 
        .ZN(n1091) );
  INV_X1 U285 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U286 ( .A1(data_in[3]), .A2(n841), .B1(n1093), .B2(\mem[12][3] ), 
        .ZN(n1090) );
  INV_X1 U287 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U288 ( .A1(data_in[4]), .A2(n841), .B1(n1093), .B2(\mem[12][4] ), 
        .ZN(n1089) );
  INV_X1 U289 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U290 ( .A1(data_in[5]), .A2(n841), .B1(n1093), .B2(\mem[12][5] ), 
        .ZN(n1088) );
  INV_X1 U291 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U292 ( .A1(data_in[6]), .A2(n841), .B1(n1093), .B2(\mem[12][6] ), 
        .ZN(n1087) );
  INV_X1 U293 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U294 ( .A1(data_in[7]), .A2(n841), .B1(n1093), .B2(\mem[12][7] ), 
        .ZN(n1086) );
  INV_X1 U295 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U296 ( .A1(data_in[0]), .A2(n840), .B1(n1084), .B2(\mem[13][0] ), 
        .ZN(n1085) );
  INV_X1 U297 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U298 ( .A1(data_in[1]), .A2(n840), .B1(n1084), .B2(\mem[13][1] ), 
        .ZN(n1083) );
  INV_X1 U299 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U300 ( .A1(data_in[2]), .A2(n840), .B1(n1084), .B2(\mem[13][2] ), 
        .ZN(n1082) );
  INV_X1 U301 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U302 ( .A1(data_in[3]), .A2(n840), .B1(n1084), .B2(\mem[13][3] ), 
        .ZN(n1081) );
  INV_X1 U303 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U304 ( .A1(data_in[4]), .A2(n840), .B1(n1084), .B2(\mem[13][4] ), 
        .ZN(n1080) );
  INV_X1 U305 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U306 ( .A1(data_in[5]), .A2(n840), .B1(n1084), .B2(\mem[13][5] ), 
        .ZN(n1079) );
  INV_X1 U307 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U308 ( .A1(data_in[6]), .A2(n840), .B1(n1084), .B2(\mem[13][6] ), 
        .ZN(n1078) );
  INV_X1 U309 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U310 ( .A1(data_in[7]), .A2(n840), .B1(n1084), .B2(\mem[13][7] ), 
        .ZN(n1077) );
  INV_X1 U311 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U312 ( .A1(data_in[0]), .A2(n839), .B1(n1075), .B2(\mem[14][0] ), 
        .ZN(n1076) );
  INV_X1 U313 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U314 ( .A1(data_in[1]), .A2(n839), .B1(n1075), .B2(\mem[14][1] ), 
        .ZN(n1074) );
  INV_X1 U315 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U316 ( .A1(data_in[2]), .A2(n839), .B1(n1075), .B2(\mem[14][2] ), 
        .ZN(n1073) );
  INV_X1 U317 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U318 ( .A1(data_in[3]), .A2(n839), .B1(n1075), .B2(\mem[14][3] ), 
        .ZN(n1072) );
  INV_X1 U319 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U320 ( .A1(data_in[4]), .A2(n839), .B1(n1075), .B2(\mem[14][4] ), 
        .ZN(n1071) );
  INV_X1 U321 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U322 ( .A1(data_in[5]), .A2(n839), .B1(n1075), .B2(\mem[14][5] ), 
        .ZN(n1070) );
  INV_X1 U323 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U324 ( .A1(data_in[6]), .A2(n839), .B1(n1075), .B2(\mem[14][6] ), 
        .ZN(n1069) );
  INV_X1 U325 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U326 ( .A1(data_in[7]), .A2(n839), .B1(n1075), .B2(\mem[14][7] ), 
        .ZN(n1068) );
  INV_X1 U327 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U328 ( .A1(data_in[0]), .A2(n838), .B1(n1066), .B2(\mem[15][0] ), 
        .ZN(n1067) );
  INV_X1 U329 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U330 ( .A1(data_in[1]), .A2(n838), .B1(n1066), .B2(\mem[15][1] ), 
        .ZN(n1065) );
  INV_X1 U331 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U332 ( .A1(data_in[2]), .A2(n838), .B1(n1066), .B2(\mem[15][2] ), 
        .ZN(n1064) );
  INV_X1 U333 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U334 ( .A1(data_in[3]), .A2(n838), .B1(n1066), .B2(\mem[15][3] ), 
        .ZN(n1063) );
  INV_X1 U335 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U336 ( .A1(data_in[4]), .A2(n838), .B1(n1066), .B2(\mem[15][4] ), 
        .ZN(n1062) );
  INV_X1 U337 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U338 ( .A1(data_in[5]), .A2(n838), .B1(n1066), .B2(\mem[15][5] ), 
        .ZN(n1061) );
  INV_X1 U339 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U340 ( .A1(data_in[6]), .A2(n838), .B1(n1066), .B2(\mem[15][6] ), 
        .ZN(n1060) );
  INV_X1 U341 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U342 ( .A1(data_in[7]), .A2(n838), .B1(n1066), .B2(\mem[15][7] ), 
        .ZN(n1059) );
  INV_X1 U343 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U344 ( .A1(data_in[0]), .A2(n837), .B1(n1057), .B2(\mem[16][0] ), 
        .ZN(n1058) );
  INV_X1 U345 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U346 ( .A1(data_in[1]), .A2(n837), .B1(n1057), .B2(\mem[16][1] ), 
        .ZN(n1056) );
  INV_X1 U347 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U348 ( .A1(data_in[2]), .A2(n837), .B1(n1057), .B2(\mem[16][2] ), 
        .ZN(n1055) );
  INV_X1 U349 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U350 ( .A1(data_in[3]), .A2(n837), .B1(n1057), .B2(\mem[16][3] ), 
        .ZN(n1054) );
  INV_X1 U351 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U352 ( .A1(data_in[4]), .A2(n837), .B1(n1057), .B2(\mem[16][4] ), 
        .ZN(n1053) );
  INV_X1 U353 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U354 ( .A1(data_in[5]), .A2(n837), .B1(n1057), .B2(\mem[16][5] ), 
        .ZN(n1052) );
  INV_X1 U355 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U356 ( .A1(data_in[6]), .A2(n837), .B1(n1057), .B2(\mem[16][6] ), 
        .ZN(n1051) );
  INV_X1 U357 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U358 ( .A1(data_in[7]), .A2(n837), .B1(n1057), .B2(\mem[16][7] ), 
        .ZN(n1050) );
  INV_X1 U359 ( .A(n1048), .ZN(n749) );
  AOI22_X1 U360 ( .A1(data_in[0]), .A2(n836), .B1(n1047), .B2(\mem[17][0] ), 
        .ZN(n1048) );
  INV_X1 U361 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U362 ( .A1(data_in[1]), .A2(n836), .B1(n1047), .B2(\mem[17][1] ), 
        .ZN(n1046) );
  INV_X1 U363 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U364 ( .A1(data_in[2]), .A2(n836), .B1(n1047), .B2(\mem[17][2] ), 
        .ZN(n1045) );
  INV_X1 U365 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U366 ( .A1(data_in[3]), .A2(n836), .B1(n1047), .B2(\mem[17][3] ), 
        .ZN(n1044) );
  INV_X1 U367 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U368 ( .A1(data_in[4]), .A2(n836), .B1(n1047), .B2(\mem[17][4] ), 
        .ZN(n1043) );
  INV_X1 U369 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U370 ( .A1(data_in[5]), .A2(n836), .B1(n1047), .B2(\mem[17][5] ), 
        .ZN(n1042) );
  INV_X1 U371 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U372 ( .A1(data_in[6]), .A2(n836), .B1(n1047), .B2(\mem[17][6] ), 
        .ZN(n1041) );
  INV_X1 U373 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U374 ( .A1(data_in[7]), .A2(n836), .B1(n1047), .B2(\mem[17][7] ), 
        .ZN(n1040) );
  INV_X1 U375 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U376 ( .A1(data_in[0]), .A2(n835), .B1(n1038), .B2(\mem[18][0] ), 
        .ZN(n1039) );
  INV_X1 U377 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U378 ( .A1(data_in[1]), .A2(n835), .B1(n1038), .B2(\mem[18][1] ), 
        .ZN(n1037) );
  INV_X1 U379 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U380 ( .A1(data_in[2]), .A2(n835), .B1(n1038), .B2(\mem[18][2] ), 
        .ZN(n1036) );
  INV_X1 U381 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U382 ( .A1(data_in[3]), .A2(n835), .B1(n1038), .B2(\mem[18][3] ), 
        .ZN(n1035) );
  INV_X1 U383 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U384 ( .A1(data_in[4]), .A2(n835), .B1(n1038), .B2(\mem[18][4] ), 
        .ZN(n1034) );
  INV_X1 U385 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U386 ( .A1(data_in[5]), .A2(n835), .B1(n1038), .B2(\mem[18][5] ), 
        .ZN(n1033) );
  INV_X1 U387 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U388 ( .A1(data_in[6]), .A2(n835), .B1(n1038), .B2(\mem[18][6] ), 
        .ZN(n1032) );
  INV_X1 U389 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U390 ( .A1(data_in[7]), .A2(n835), .B1(n1038), .B2(\mem[18][7] ), 
        .ZN(n1031) );
  INV_X1 U391 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U392 ( .A1(data_in[0]), .A2(n834), .B1(n1029), .B2(\mem[19][0] ), 
        .ZN(n1030) );
  INV_X1 U393 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U394 ( .A1(data_in[1]), .A2(n834), .B1(n1029), .B2(\mem[19][1] ), 
        .ZN(n1028) );
  INV_X1 U395 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U396 ( .A1(data_in[2]), .A2(n834), .B1(n1029), .B2(\mem[19][2] ), 
        .ZN(n1027) );
  INV_X1 U397 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U398 ( .A1(data_in[3]), .A2(n834), .B1(n1029), .B2(\mem[19][3] ), 
        .ZN(n1026) );
  INV_X1 U399 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U400 ( .A1(data_in[4]), .A2(n834), .B1(n1029), .B2(\mem[19][4] ), 
        .ZN(n1025) );
  INV_X1 U401 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U402 ( .A1(data_in[5]), .A2(n834), .B1(n1029), .B2(\mem[19][5] ), 
        .ZN(n1024) );
  INV_X1 U403 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U404 ( .A1(data_in[6]), .A2(n834), .B1(n1029), .B2(\mem[19][6] ), 
        .ZN(n1023) );
  INV_X1 U405 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U406 ( .A1(data_in[7]), .A2(n834), .B1(n1029), .B2(\mem[19][7] ), 
        .ZN(n1022) );
  INV_X1 U407 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U408 ( .A1(data_in[0]), .A2(n833), .B1(n1020), .B2(\mem[20][0] ), 
        .ZN(n1021) );
  INV_X1 U409 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U410 ( .A1(data_in[1]), .A2(n833), .B1(n1020), .B2(\mem[20][1] ), 
        .ZN(n1019) );
  INV_X1 U411 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U412 ( .A1(data_in[2]), .A2(n833), .B1(n1020), .B2(\mem[20][2] ), 
        .ZN(n1018) );
  INV_X1 U413 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U414 ( .A1(data_in[3]), .A2(n833), .B1(n1020), .B2(\mem[20][3] ), 
        .ZN(n1017) );
  INV_X1 U415 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U416 ( .A1(data_in[4]), .A2(n833), .B1(n1020), .B2(\mem[20][4] ), 
        .ZN(n1016) );
  INV_X1 U417 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U418 ( .A1(data_in[5]), .A2(n833), .B1(n1020), .B2(\mem[20][5] ), 
        .ZN(n1015) );
  INV_X1 U419 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U420 ( .A1(data_in[6]), .A2(n833), .B1(n1020), .B2(\mem[20][6] ), 
        .ZN(n1014) );
  INV_X1 U421 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U422 ( .A1(data_in[7]), .A2(n833), .B1(n1020), .B2(\mem[20][7] ), 
        .ZN(n1013) );
  INV_X1 U423 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U424 ( .A1(data_in[0]), .A2(n832), .B1(n1011), .B2(\mem[21][0] ), 
        .ZN(n1012) );
  INV_X1 U425 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U426 ( .A1(data_in[1]), .A2(n832), .B1(n1011), .B2(\mem[21][1] ), 
        .ZN(n1010) );
  INV_X1 U427 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U428 ( .A1(data_in[2]), .A2(n832), .B1(n1011), .B2(\mem[21][2] ), 
        .ZN(n1009) );
  INV_X1 U429 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U430 ( .A1(data_in[3]), .A2(n832), .B1(n1011), .B2(\mem[21][3] ), 
        .ZN(n1008) );
  INV_X1 U431 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U432 ( .A1(data_in[4]), .A2(n832), .B1(n1011), .B2(\mem[21][4] ), 
        .ZN(n1007) );
  INV_X1 U433 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U434 ( .A1(data_in[5]), .A2(n832), .B1(n1011), .B2(\mem[21][5] ), 
        .ZN(n1006) );
  INV_X1 U435 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U436 ( .A1(data_in[6]), .A2(n832), .B1(n1011), .B2(\mem[21][6] ), 
        .ZN(n1005) );
  INV_X1 U437 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U438 ( .A1(data_in[7]), .A2(n832), .B1(n1011), .B2(\mem[21][7] ), 
        .ZN(n1004) );
  INV_X1 U439 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U440 ( .A1(data_in[0]), .A2(n831), .B1(n1002), .B2(\mem[22][0] ), 
        .ZN(n1003) );
  INV_X1 U441 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U442 ( .A1(data_in[1]), .A2(n831), .B1(n1002), .B2(\mem[22][1] ), 
        .ZN(n1001) );
  INV_X1 U443 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U444 ( .A1(data_in[2]), .A2(n831), .B1(n1002), .B2(\mem[22][2] ), 
        .ZN(n1000) );
  INV_X1 U445 ( .A(n999), .ZN(n706) );
  AOI22_X1 U446 ( .A1(data_in[3]), .A2(n831), .B1(n1002), .B2(\mem[22][3] ), 
        .ZN(n999) );
  INV_X1 U447 ( .A(n998), .ZN(n705) );
  AOI22_X1 U448 ( .A1(data_in[4]), .A2(n831), .B1(n1002), .B2(\mem[22][4] ), 
        .ZN(n998) );
  INV_X1 U449 ( .A(n997), .ZN(n704) );
  AOI22_X1 U450 ( .A1(data_in[5]), .A2(n831), .B1(n1002), .B2(\mem[22][5] ), 
        .ZN(n997) );
  INV_X1 U451 ( .A(n996), .ZN(n703) );
  AOI22_X1 U452 ( .A1(data_in[6]), .A2(n831), .B1(n1002), .B2(\mem[22][6] ), 
        .ZN(n996) );
  INV_X1 U453 ( .A(n995), .ZN(n702) );
  AOI22_X1 U454 ( .A1(data_in[7]), .A2(n831), .B1(n1002), .B2(\mem[22][7] ), 
        .ZN(n995) );
  INV_X1 U455 ( .A(n994), .ZN(n701) );
  AOI22_X1 U456 ( .A1(data_in[0]), .A2(n830), .B1(n993), .B2(\mem[23][0] ), 
        .ZN(n994) );
  INV_X1 U457 ( .A(n992), .ZN(n700) );
  AOI22_X1 U458 ( .A1(data_in[1]), .A2(n830), .B1(n993), .B2(\mem[23][1] ), 
        .ZN(n992) );
  INV_X1 U459 ( .A(n991), .ZN(n699) );
  AOI22_X1 U460 ( .A1(data_in[2]), .A2(n830), .B1(n993), .B2(\mem[23][2] ), 
        .ZN(n991) );
  INV_X1 U461 ( .A(n990), .ZN(n698) );
  AOI22_X1 U462 ( .A1(data_in[3]), .A2(n830), .B1(n993), .B2(\mem[23][3] ), 
        .ZN(n990) );
  INV_X1 U463 ( .A(n989), .ZN(n697) );
  AOI22_X1 U464 ( .A1(data_in[4]), .A2(n830), .B1(n993), .B2(\mem[23][4] ), 
        .ZN(n989) );
  INV_X1 U465 ( .A(n988), .ZN(n696) );
  AOI22_X1 U466 ( .A1(data_in[5]), .A2(n830), .B1(n993), .B2(\mem[23][5] ), 
        .ZN(n988) );
  INV_X1 U467 ( .A(n987), .ZN(n695) );
  AOI22_X1 U468 ( .A1(data_in[6]), .A2(n830), .B1(n993), .B2(\mem[23][6] ), 
        .ZN(n987) );
  INV_X1 U469 ( .A(n986), .ZN(n694) );
  AOI22_X1 U470 ( .A1(data_in[7]), .A2(n830), .B1(n993), .B2(\mem[23][7] ), 
        .ZN(n986) );
  INV_X1 U471 ( .A(n985), .ZN(n693) );
  AOI22_X1 U472 ( .A1(data_in[0]), .A2(n829), .B1(n984), .B2(\mem[24][0] ), 
        .ZN(n985) );
  INV_X1 U473 ( .A(n983), .ZN(n692) );
  AOI22_X1 U474 ( .A1(data_in[1]), .A2(n829), .B1(n984), .B2(\mem[24][1] ), 
        .ZN(n983) );
  INV_X1 U475 ( .A(n982), .ZN(n691) );
  AOI22_X1 U476 ( .A1(data_in[2]), .A2(n829), .B1(n984), .B2(\mem[24][2] ), 
        .ZN(n982) );
  INV_X1 U477 ( .A(n981), .ZN(n690) );
  AOI22_X1 U478 ( .A1(data_in[3]), .A2(n829), .B1(n984), .B2(\mem[24][3] ), 
        .ZN(n981) );
  INV_X1 U479 ( .A(n980), .ZN(n689) );
  AOI22_X1 U480 ( .A1(data_in[4]), .A2(n829), .B1(n984), .B2(\mem[24][4] ), 
        .ZN(n980) );
  INV_X1 U481 ( .A(n979), .ZN(n688) );
  AOI22_X1 U482 ( .A1(data_in[5]), .A2(n829), .B1(n984), .B2(\mem[24][5] ), 
        .ZN(n979) );
  INV_X1 U483 ( .A(n978), .ZN(n687) );
  AOI22_X1 U484 ( .A1(data_in[6]), .A2(n829), .B1(n984), .B2(\mem[24][6] ), 
        .ZN(n978) );
  INV_X1 U485 ( .A(n977), .ZN(n686) );
  AOI22_X1 U486 ( .A1(data_in[7]), .A2(n829), .B1(n984), .B2(\mem[24][7] ), 
        .ZN(n977) );
  INV_X1 U487 ( .A(n975), .ZN(n685) );
  AOI22_X1 U488 ( .A1(data_in[0]), .A2(n828), .B1(n974), .B2(\mem[25][0] ), 
        .ZN(n975) );
  INV_X1 U489 ( .A(n973), .ZN(n684) );
  AOI22_X1 U490 ( .A1(data_in[1]), .A2(n828), .B1(n974), .B2(\mem[25][1] ), 
        .ZN(n973) );
  INV_X1 U491 ( .A(n972), .ZN(n683) );
  AOI22_X1 U492 ( .A1(data_in[2]), .A2(n828), .B1(n974), .B2(\mem[25][2] ), 
        .ZN(n972) );
  INV_X1 U493 ( .A(n971), .ZN(n682) );
  AOI22_X1 U494 ( .A1(data_in[3]), .A2(n828), .B1(n974), .B2(\mem[25][3] ), 
        .ZN(n971) );
  INV_X1 U495 ( .A(n970), .ZN(n681) );
  AOI22_X1 U496 ( .A1(data_in[4]), .A2(n828), .B1(n974), .B2(\mem[25][4] ), 
        .ZN(n970) );
  INV_X1 U497 ( .A(n969), .ZN(n680) );
  AOI22_X1 U498 ( .A1(data_in[5]), .A2(n828), .B1(n974), .B2(\mem[25][5] ), 
        .ZN(n969) );
  INV_X1 U499 ( .A(n968), .ZN(n679) );
  AOI22_X1 U500 ( .A1(data_in[6]), .A2(n828), .B1(n974), .B2(\mem[25][6] ), 
        .ZN(n968) );
  INV_X1 U501 ( .A(n967), .ZN(n678) );
  AOI22_X1 U502 ( .A1(data_in[7]), .A2(n828), .B1(n974), .B2(\mem[25][7] ), 
        .ZN(n967) );
  INV_X1 U503 ( .A(n966), .ZN(n677) );
  AOI22_X1 U504 ( .A1(data_in[0]), .A2(n827), .B1(n965), .B2(\mem[26][0] ), 
        .ZN(n966) );
  INV_X1 U505 ( .A(n964), .ZN(n676) );
  AOI22_X1 U506 ( .A1(data_in[1]), .A2(n827), .B1(n965), .B2(\mem[26][1] ), 
        .ZN(n964) );
  INV_X1 U507 ( .A(n963), .ZN(n675) );
  AOI22_X1 U508 ( .A1(data_in[2]), .A2(n827), .B1(n965), .B2(\mem[26][2] ), 
        .ZN(n963) );
  INV_X1 U509 ( .A(n962), .ZN(n674) );
  AOI22_X1 U510 ( .A1(data_in[3]), .A2(n827), .B1(n965), .B2(\mem[26][3] ), 
        .ZN(n962) );
  INV_X1 U511 ( .A(n961), .ZN(n673) );
  AOI22_X1 U512 ( .A1(data_in[4]), .A2(n827), .B1(n965), .B2(\mem[26][4] ), 
        .ZN(n961) );
  INV_X1 U513 ( .A(n960), .ZN(n672) );
  AOI22_X1 U514 ( .A1(data_in[5]), .A2(n827), .B1(n965), .B2(\mem[26][5] ), 
        .ZN(n960) );
  INV_X1 U515 ( .A(n959), .ZN(n671) );
  AOI22_X1 U516 ( .A1(data_in[6]), .A2(n827), .B1(n965), .B2(\mem[26][6] ), 
        .ZN(n959) );
  INV_X1 U517 ( .A(n958), .ZN(n670) );
  AOI22_X1 U518 ( .A1(data_in[7]), .A2(n827), .B1(n965), .B2(\mem[26][7] ), 
        .ZN(n958) );
  INV_X1 U519 ( .A(n957), .ZN(n669) );
  AOI22_X1 U520 ( .A1(data_in[0]), .A2(n826), .B1(n956), .B2(\mem[27][0] ), 
        .ZN(n957) );
  INV_X1 U521 ( .A(n955), .ZN(n668) );
  AOI22_X1 U522 ( .A1(data_in[1]), .A2(n826), .B1(n956), .B2(\mem[27][1] ), 
        .ZN(n955) );
  INV_X1 U523 ( .A(n954), .ZN(n667) );
  AOI22_X1 U524 ( .A1(data_in[2]), .A2(n826), .B1(n956), .B2(\mem[27][2] ), 
        .ZN(n954) );
  INV_X1 U525 ( .A(n953), .ZN(n666) );
  AOI22_X1 U526 ( .A1(data_in[3]), .A2(n826), .B1(n956), .B2(\mem[27][3] ), 
        .ZN(n953) );
  INV_X1 U527 ( .A(n952), .ZN(n665) );
  AOI22_X1 U528 ( .A1(data_in[4]), .A2(n826), .B1(n956), .B2(\mem[27][4] ), 
        .ZN(n952) );
  INV_X1 U529 ( .A(n951), .ZN(n664) );
  AOI22_X1 U530 ( .A1(data_in[5]), .A2(n826), .B1(n956), .B2(\mem[27][5] ), 
        .ZN(n951) );
  INV_X1 U531 ( .A(n950), .ZN(n663) );
  AOI22_X1 U532 ( .A1(data_in[6]), .A2(n826), .B1(n956), .B2(\mem[27][6] ), 
        .ZN(n950) );
  INV_X1 U533 ( .A(n949), .ZN(n662) );
  AOI22_X1 U534 ( .A1(data_in[7]), .A2(n826), .B1(n956), .B2(\mem[27][7] ), 
        .ZN(n949) );
  INV_X1 U535 ( .A(n948), .ZN(n661) );
  AOI22_X1 U536 ( .A1(data_in[0]), .A2(n825), .B1(n947), .B2(\mem[28][0] ), 
        .ZN(n948) );
  INV_X1 U537 ( .A(n946), .ZN(n660) );
  AOI22_X1 U538 ( .A1(data_in[1]), .A2(n825), .B1(n947), .B2(\mem[28][1] ), 
        .ZN(n946) );
  INV_X1 U539 ( .A(n945), .ZN(n659) );
  AOI22_X1 U540 ( .A1(data_in[2]), .A2(n825), .B1(n947), .B2(\mem[28][2] ), 
        .ZN(n945) );
  INV_X1 U541 ( .A(n944), .ZN(n658) );
  AOI22_X1 U542 ( .A1(data_in[3]), .A2(n825), .B1(n947), .B2(\mem[28][3] ), 
        .ZN(n944) );
  INV_X1 U543 ( .A(n943), .ZN(n657) );
  AOI22_X1 U544 ( .A1(data_in[4]), .A2(n825), .B1(n947), .B2(\mem[28][4] ), 
        .ZN(n943) );
  INV_X1 U545 ( .A(n942), .ZN(n656) );
  AOI22_X1 U546 ( .A1(data_in[5]), .A2(n825), .B1(n947), .B2(\mem[28][5] ), 
        .ZN(n942) );
  INV_X1 U547 ( .A(n941), .ZN(n655) );
  AOI22_X1 U548 ( .A1(data_in[6]), .A2(n825), .B1(n947), .B2(\mem[28][6] ), 
        .ZN(n941) );
  INV_X1 U549 ( .A(n940), .ZN(n654) );
  AOI22_X1 U550 ( .A1(data_in[7]), .A2(n825), .B1(n947), .B2(\mem[28][7] ), 
        .ZN(n940) );
  INV_X1 U551 ( .A(n939), .ZN(n653) );
  AOI22_X1 U552 ( .A1(data_in[0]), .A2(n824), .B1(n938), .B2(\mem[29][0] ), 
        .ZN(n939) );
  INV_X1 U553 ( .A(n937), .ZN(n652) );
  AOI22_X1 U554 ( .A1(data_in[1]), .A2(n824), .B1(n938), .B2(\mem[29][1] ), 
        .ZN(n937) );
  INV_X1 U555 ( .A(n936), .ZN(n651) );
  AOI22_X1 U556 ( .A1(data_in[2]), .A2(n824), .B1(n938), .B2(\mem[29][2] ), 
        .ZN(n936) );
  INV_X1 U557 ( .A(n935), .ZN(n650) );
  AOI22_X1 U558 ( .A1(data_in[3]), .A2(n824), .B1(n938), .B2(\mem[29][3] ), 
        .ZN(n935) );
  INV_X1 U559 ( .A(n934), .ZN(n649) );
  AOI22_X1 U560 ( .A1(data_in[4]), .A2(n824), .B1(n938), .B2(\mem[29][4] ), 
        .ZN(n934) );
  INV_X1 U561 ( .A(n933), .ZN(n648) );
  AOI22_X1 U562 ( .A1(data_in[5]), .A2(n824), .B1(n938), .B2(\mem[29][5] ), 
        .ZN(n933) );
  INV_X1 U563 ( .A(n932), .ZN(n647) );
  AOI22_X1 U564 ( .A1(data_in[6]), .A2(n824), .B1(n938), .B2(\mem[29][6] ), 
        .ZN(n932) );
  INV_X1 U565 ( .A(n931), .ZN(n646) );
  AOI22_X1 U566 ( .A1(data_in[7]), .A2(n824), .B1(n938), .B2(\mem[29][7] ), 
        .ZN(n931) );
  INV_X1 U567 ( .A(n930), .ZN(n645) );
  AOI22_X1 U568 ( .A1(data_in[0]), .A2(n823), .B1(n929), .B2(\mem[30][0] ), 
        .ZN(n930) );
  INV_X1 U569 ( .A(n928), .ZN(n644) );
  AOI22_X1 U570 ( .A1(data_in[1]), .A2(n823), .B1(n929), .B2(\mem[30][1] ), 
        .ZN(n928) );
  INV_X1 U571 ( .A(n927), .ZN(n643) );
  AOI22_X1 U572 ( .A1(data_in[2]), .A2(n823), .B1(n929), .B2(\mem[30][2] ), 
        .ZN(n927) );
  INV_X1 U573 ( .A(n926), .ZN(n642) );
  AOI22_X1 U574 ( .A1(data_in[3]), .A2(n823), .B1(n929), .B2(\mem[30][3] ), 
        .ZN(n926) );
  INV_X1 U575 ( .A(n925), .ZN(n641) );
  AOI22_X1 U576 ( .A1(data_in[4]), .A2(n823), .B1(n929), .B2(\mem[30][4] ), 
        .ZN(n925) );
  INV_X1 U577 ( .A(n924), .ZN(n640) );
  AOI22_X1 U578 ( .A1(data_in[5]), .A2(n823), .B1(n929), .B2(\mem[30][5] ), 
        .ZN(n924) );
  INV_X1 U579 ( .A(n923), .ZN(n639) );
  AOI22_X1 U580 ( .A1(data_in[6]), .A2(n823), .B1(n929), .B2(\mem[30][6] ), 
        .ZN(n923) );
  INV_X1 U581 ( .A(n922), .ZN(n638) );
  AOI22_X1 U582 ( .A1(data_in[7]), .A2(n823), .B1(n929), .B2(\mem[30][7] ), 
        .ZN(n922) );
  INV_X1 U583 ( .A(n921), .ZN(n637) );
  AOI22_X1 U584 ( .A1(data_in[0]), .A2(n822), .B1(n920), .B2(\mem[31][0] ), 
        .ZN(n921) );
  INV_X1 U585 ( .A(n919), .ZN(n636) );
  AOI22_X1 U586 ( .A1(data_in[1]), .A2(n822), .B1(n920), .B2(\mem[31][1] ), 
        .ZN(n919) );
  INV_X1 U587 ( .A(n918), .ZN(n635) );
  AOI22_X1 U588 ( .A1(data_in[2]), .A2(n822), .B1(n920), .B2(\mem[31][2] ), 
        .ZN(n918) );
  INV_X1 U589 ( .A(n917), .ZN(n634) );
  AOI22_X1 U590 ( .A1(data_in[3]), .A2(n822), .B1(n920), .B2(\mem[31][3] ), 
        .ZN(n917) );
  INV_X1 U591 ( .A(n916), .ZN(n633) );
  AOI22_X1 U592 ( .A1(data_in[4]), .A2(n822), .B1(n920), .B2(\mem[31][4] ), 
        .ZN(n916) );
  INV_X1 U593 ( .A(n915), .ZN(n632) );
  AOI22_X1 U594 ( .A1(data_in[5]), .A2(n822), .B1(n920), .B2(\mem[31][5] ), 
        .ZN(n915) );
  INV_X1 U595 ( .A(n914), .ZN(n631) );
  AOI22_X1 U596 ( .A1(data_in[6]), .A2(n822), .B1(n920), .B2(\mem[31][6] ), 
        .ZN(n914) );
  INV_X1 U597 ( .A(n913), .ZN(n630) );
  AOI22_X1 U598 ( .A1(data_in[7]), .A2(n822), .B1(n920), .B2(\mem[31][7] ), 
        .ZN(n913) );
  MUX2_X1 U599 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n612), .Z(n2) );
  MUX2_X1 U600 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n612), .Z(n3) );
  MUX2_X1 U601 ( .A(n3), .B(n2), .S(n609), .Z(n4) );
  MUX2_X1 U602 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n612), .Z(n5) );
  MUX2_X1 U603 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n612), .Z(n6) );
  MUX2_X1 U604 ( .A(n6), .B(n5), .S(n609), .Z(n7) );
  MUX2_X1 U605 ( .A(n7), .B(n4), .S(n607), .Z(n8) );
  MUX2_X1 U606 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n612), .Z(n9) );
  MUX2_X1 U607 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n612), .Z(n10) );
  MUX2_X1 U608 ( .A(n10), .B(n9), .S(n609), .Z(n11) );
  MUX2_X1 U609 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n612), .Z(n12) );
  MUX2_X1 U610 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n612), .Z(n13) );
  MUX2_X1 U611 ( .A(n13), .B(n12), .S(n609), .Z(n14) );
  MUX2_X1 U612 ( .A(n14), .B(n11), .S(N12), .Z(n15) );
  MUX2_X1 U613 ( .A(n15), .B(n8), .S(N13), .Z(n16) );
  MUX2_X1 U614 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n613), .Z(n17) );
  MUX2_X1 U615 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n619), .Z(n18) );
  MUX2_X1 U616 ( .A(n18), .B(n17), .S(n609), .Z(n19) );
  MUX2_X1 U617 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n619), .Z(n20) );
  MUX2_X1 U618 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n619), .Z(n21) );
  MUX2_X1 U619 ( .A(n21), .B(n20), .S(n610), .Z(n22) );
  MUX2_X1 U620 ( .A(n22), .B(n19), .S(N12), .Z(n23) );
  MUX2_X1 U621 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n612), .Z(n24) );
  MUX2_X1 U622 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n619), .Z(n25) );
  MUX2_X1 U623 ( .A(n25), .B(n24), .S(n609), .Z(n26) );
  MUX2_X1 U624 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n619), .Z(n27) );
  MUX2_X1 U625 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n619), .Z(n28) );
  MUX2_X1 U626 ( .A(n28), .B(n27), .S(n611), .Z(n29) );
  MUX2_X1 U627 ( .A(n29), .B(n26), .S(n608), .Z(n30) );
  MUX2_X1 U628 ( .A(n30), .B(n23), .S(N13), .Z(n31) );
  MUX2_X1 U629 ( .A(n31), .B(n16), .S(N14), .Z(N22) );
  MUX2_X1 U630 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n619), .Z(n32) );
  MUX2_X1 U631 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n615), .Z(n33) );
  MUX2_X1 U632 ( .A(n33), .B(n32), .S(n609), .Z(n34) );
  MUX2_X1 U633 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n618), .Z(n35) );
  MUX2_X1 U634 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n619), .Z(n36) );
  MUX2_X1 U635 ( .A(n36), .B(n35), .S(n609), .Z(n37) );
  MUX2_X1 U636 ( .A(n37), .B(n34), .S(n608), .Z(n38) );
  MUX2_X1 U637 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n613), .Z(n39) );
  MUX2_X1 U638 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n613), .Z(n40) );
  MUX2_X1 U639 ( .A(n40), .B(n39), .S(n609), .Z(n41) );
  MUX2_X1 U640 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n613), .Z(n42) );
  MUX2_X1 U641 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n613), .Z(n43) );
  MUX2_X1 U642 ( .A(n43), .B(n42), .S(N11), .Z(n44) );
  MUX2_X1 U643 ( .A(n44), .B(n41), .S(N12), .Z(n45) );
  MUX2_X1 U644 ( .A(n45), .B(n38), .S(N13), .Z(n46) );
  MUX2_X1 U645 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n613), .Z(n47) );
  MUX2_X1 U646 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n613), .Z(n48) );
  MUX2_X1 U647 ( .A(n48), .B(n47), .S(n609), .Z(n49) );
  MUX2_X1 U648 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n613), .Z(n50) );
  MUX2_X1 U649 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n613), .Z(n51) );
  MUX2_X1 U650 ( .A(n51), .B(n50), .S(n611), .Z(n52) );
  MUX2_X1 U651 ( .A(n52), .B(n49), .S(n607), .Z(n53) );
  MUX2_X1 U652 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n613), .Z(n54) );
  MUX2_X1 U653 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n613), .Z(n55) );
  MUX2_X1 U654 ( .A(n55), .B(n54), .S(n609), .Z(n56) );
  MUX2_X1 U655 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n613), .Z(n57) );
  MUX2_X1 U656 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n613), .Z(n58) );
  MUX2_X1 U657 ( .A(n58), .B(n57), .S(n609), .Z(n59) );
  MUX2_X1 U658 ( .A(n59), .B(n56), .S(n607), .Z(n60) );
  MUX2_X1 U659 ( .A(n60), .B(n53), .S(N13), .Z(n61) );
  MUX2_X1 U660 ( .A(n61), .B(n46), .S(N14), .Z(N21) );
  MUX2_X1 U661 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n617), .Z(n62) );
  MUX2_X1 U662 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n617), .Z(n63) );
  MUX2_X1 U663 ( .A(n63), .B(n62), .S(n610), .Z(n64) );
  MUX2_X1 U664 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n614), .Z(n65) );
  MUX2_X1 U665 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n614), .Z(n66) );
  MUX2_X1 U666 ( .A(n66), .B(n65), .S(n610), .Z(n67) );
  MUX2_X1 U667 ( .A(n67), .B(n64), .S(n607), .Z(n68) );
  MUX2_X1 U668 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n614), .Z(n69) );
  MUX2_X1 U669 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n617), .Z(n70) );
  MUX2_X1 U670 ( .A(n70), .B(n69), .S(n610), .Z(n71) );
  MUX2_X1 U671 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n617), .Z(n72) );
  MUX2_X1 U672 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n619), .Z(n73) );
  MUX2_X1 U673 ( .A(n73), .B(n72), .S(n610), .Z(n74) );
  MUX2_X1 U674 ( .A(n74), .B(n71), .S(n607), .Z(n75) );
  MUX2_X1 U675 ( .A(n75), .B(n68), .S(N13), .Z(n76) );
  MUX2_X1 U676 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n617), .Z(n77) );
  MUX2_X1 U677 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n619), .Z(n78) );
  MUX2_X1 U678 ( .A(n78), .B(n77), .S(n610), .Z(n79) );
  MUX2_X1 U679 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n614), .Z(n80) );
  MUX2_X1 U680 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n614), .Z(n81) );
  MUX2_X1 U681 ( .A(n81), .B(n80), .S(n610), .Z(n82) );
  MUX2_X1 U682 ( .A(n82), .B(n79), .S(n607), .Z(n83) );
  MUX2_X1 U683 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n614), .Z(n84) );
  MUX2_X1 U684 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n617), .Z(n85) );
  MUX2_X1 U685 ( .A(n85), .B(n84), .S(n610), .Z(n86) );
  MUX2_X1 U686 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n617), .Z(n87) );
  MUX2_X1 U687 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n614), .Z(n88) );
  MUX2_X1 U688 ( .A(n88), .B(n87), .S(n610), .Z(n89) );
  MUX2_X1 U689 ( .A(n89), .B(n86), .S(n607), .Z(n90) );
  MUX2_X1 U690 ( .A(n90), .B(n83), .S(N13), .Z(n91) );
  MUX2_X1 U691 ( .A(n91), .B(n76), .S(N14), .Z(N20) );
  MUX2_X1 U692 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n617), .Z(n92) );
  MUX2_X1 U693 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n614), .Z(n93) );
  MUX2_X1 U694 ( .A(n93), .B(n92), .S(n610), .Z(n94) );
  MUX2_X1 U695 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n614), .Z(n95) );
  MUX2_X1 U696 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n617), .Z(n96) );
  MUX2_X1 U697 ( .A(n96), .B(n95), .S(n610), .Z(n97) );
  MUX2_X1 U698 ( .A(n97), .B(n94), .S(n607), .Z(n98) );
  MUX2_X1 U699 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n617), .Z(n99) );
  MUX2_X1 U700 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n614), .Z(n100) );
  MUX2_X1 U701 ( .A(n100), .B(n99), .S(n610), .Z(n101) );
  MUX2_X1 U702 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n617), .Z(n102) );
  MUX2_X1 U703 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n614), .Z(n103) );
  MUX2_X1 U704 ( .A(n103), .B(n102), .S(n610), .Z(n104) );
  MUX2_X1 U705 ( .A(n104), .B(n101), .S(n607), .Z(n105) );
  MUX2_X1 U706 ( .A(n105), .B(n98), .S(N13), .Z(n106) );
  MUX2_X1 U707 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n614), .Z(n107) );
  MUX2_X1 U708 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n614), .Z(n108) );
  MUX2_X1 U709 ( .A(n108), .B(n107), .S(n611), .Z(n109) );
  MUX2_X1 U710 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n614), .Z(n110) );
  MUX2_X1 U711 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n614), .Z(n111) );
  MUX2_X1 U712 ( .A(n111), .B(n110), .S(n611), .Z(n112) );
  MUX2_X1 U713 ( .A(n112), .B(n109), .S(n607), .Z(n113) );
  MUX2_X1 U714 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n614), .Z(n114) );
  MUX2_X1 U715 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n614), .Z(n115) );
  MUX2_X1 U716 ( .A(n115), .B(n114), .S(n611), .Z(n116) );
  MUX2_X1 U717 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n614), .Z(n117) );
  MUX2_X1 U718 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n614), .Z(n118) );
  MUX2_X1 U719 ( .A(n118), .B(n117), .S(n611), .Z(n119) );
  MUX2_X1 U720 ( .A(n119), .B(n116), .S(n607), .Z(n120) );
  MUX2_X1 U721 ( .A(n120), .B(n113), .S(N13), .Z(n121) );
  MUX2_X1 U722 ( .A(n121), .B(n106), .S(N14), .Z(N19) );
  MUX2_X1 U723 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n614), .Z(n122) );
  MUX2_X1 U724 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n614), .Z(n123) );
  MUX2_X1 U725 ( .A(n123), .B(n122), .S(n611), .Z(n124) );
  MUX2_X1 U726 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n614), .Z(n125) );
  MUX2_X1 U727 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n614), .Z(n126) );
  MUX2_X1 U728 ( .A(n126), .B(n125), .S(n611), .Z(n127) );
  MUX2_X1 U729 ( .A(n127), .B(n124), .S(n607), .Z(n128) );
  MUX2_X1 U730 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n615), .Z(n129) );
  MUX2_X1 U731 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n615), .Z(n130) );
  MUX2_X1 U732 ( .A(n130), .B(n129), .S(n611), .Z(n131) );
  MUX2_X1 U733 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n615), .Z(n132) );
  MUX2_X1 U734 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n615), .Z(n133) );
  MUX2_X1 U735 ( .A(n133), .B(n132), .S(n611), .Z(n134) );
  MUX2_X1 U736 ( .A(n134), .B(n131), .S(n607), .Z(n135) );
  MUX2_X1 U737 ( .A(n135), .B(n128), .S(N13), .Z(n136) );
  MUX2_X1 U738 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n615), .Z(n137) );
  MUX2_X1 U739 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n615), .Z(n138) );
  MUX2_X1 U740 ( .A(n138), .B(n137), .S(n611), .Z(n139) );
  MUX2_X1 U741 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n615), .Z(n140) );
  MUX2_X1 U742 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n615), .Z(n141) );
  MUX2_X1 U743 ( .A(n141), .B(n140), .S(n611), .Z(n142) );
  MUX2_X1 U744 ( .A(n142), .B(n139), .S(n607), .Z(n143) );
  MUX2_X1 U745 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n615), .Z(n144) );
  MUX2_X1 U746 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n615), .Z(n145) );
  MUX2_X1 U747 ( .A(n145), .B(n144), .S(n611), .Z(n146) );
  MUX2_X1 U748 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n615), .Z(n147) );
  MUX2_X1 U749 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n615), .Z(n148) );
  MUX2_X1 U750 ( .A(n148), .B(n147), .S(n611), .Z(n149) );
  MUX2_X1 U751 ( .A(n149), .B(n146), .S(n607), .Z(n150) );
  MUX2_X1 U752 ( .A(n150), .B(n143), .S(N13), .Z(n151) );
  MUX2_X1 U753 ( .A(n151), .B(n136), .S(N14), .Z(N18) );
  MUX2_X1 U754 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n616), .Z(n152) );
  MUX2_X1 U755 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n616), .Z(n153) );
  MUX2_X1 U756 ( .A(n153), .B(n152), .S(n609), .Z(n154) );
  MUX2_X1 U757 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n616), .Z(n155) );
  MUX2_X1 U758 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n616), .Z(n156) );
  MUX2_X1 U759 ( .A(n156), .B(n155), .S(n609), .Z(n157) );
  MUX2_X1 U760 ( .A(n157), .B(n154), .S(n608), .Z(n158) );
  MUX2_X1 U761 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n616), .Z(n159) );
  MUX2_X1 U762 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n616), .Z(n160) );
  MUX2_X1 U763 ( .A(n160), .B(n159), .S(n611), .Z(n161) );
  MUX2_X1 U764 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n616), .Z(n162) );
  MUX2_X1 U765 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n616), .Z(n163) );
  MUX2_X1 U766 ( .A(n163), .B(n162), .S(n610), .Z(n164) );
  MUX2_X1 U767 ( .A(n164), .B(n161), .S(n608), .Z(n165) );
  MUX2_X1 U768 ( .A(n165), .B(n158), .S(N13), .Z(n166) );
  MUX2_X1 U769 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n616), .Z(n167) );
  MUX2_X1 U770 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n616), .Z(n168) );
  MUX2_X1 U771 ( .A(n168), .B(n167), .S(n610), .Z(n169) );
  MUX2_X1 U772 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n616), .Z(n170) );
  MUX2_X1 U773 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n616), .Z(n171) );
  MUX2_X1 U774 ( .A(n171), .B(n170), .S(n611), .Z(n172) );
  MUX2_X1 U775 ( .A(n172), .B(n169), .S(n608), .Z(n173) );
  MUX2_X1 U776 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n612), .Z(n174) );
  MUX2_X1 U777 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n619), .Z(n175) );
  MUX2_X1 U778 ( .A(n175), .B(n174), .S(N11), .Z(n176) );
  MUX2_X1 U779 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n612), .Z(n177) );
  MUX2_X1 U780 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n612), .Z(n178) );
  MUX2_X1 U781 ( .A(n178), .B(n177), .S(n609), .Z(n179) );
  MUX2_X1 U782 ( .A(n179), .B(n176), .S(n608), .Z(n180) );
  MUX2_X1 U783 ( .A(n180), .B(n173), .S(N13), .Z(n181) );
  MUX2_X1 U784 ( .A(n181), .B(n166), .S(N14), .Z(N17) );
  MUX2_X1 U785 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(N10), .Z(n182) );
  MUX2_X1 U786 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(N10), .Z(n183) );
  MUX2_X1 U787 ( .A(n183), .B(n182), .S(n611), .Z(n184) );
  MUX2_X1 U788 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(N10), .Z(n185) );
  MUX2_X1 U789 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(N10), .Z(n186) );
  MUX2_X1 U790 ( .A(n186), .B(n185), .S(n611), .Z(n187) );
  MUX2_X1 U791 ( .A(n187), .B(n184), .S(n608), .Z(n188) );
  MUX2_X1 U792 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n612), .Z(n189) );
  MUX2_X1 U793 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n619), .Z(n190) );
  MUX2_X1 U794 ( .A(n190), .B(n189), .S(n609), .Z(n191) );
  MUX2_X1 U795 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n619), .Z(n192) );
  MUX2_X1 U796 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(N10), .Z(n193) );
  MUX2_X1 U797 ( .A(n193), .B(n192), .S(n609), .Z(n194) );
  MUX2_X1 U798 ( .A(n194), .B(n191), .S(n608), .Z(n195) );
  MUX2_X1 U799 ( .A(n195), .B(n188), .S(N13), .Z(n196) );
  MUX2_X1 U800 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n617), .Z(n197) );
  MUX2_X1 U801 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n617), .Z(n198) );
  MUX2_X1 U802 ( .A(n198), .B(n197), .S(n611), .Z(n199) );
  MUX2_X1 U803 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n617), .Z(n200) );
  MUX2_X1 U804 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n617), .Z(n201) );
  MUX2_X1 U805 ( .A(n201), .B(n200), .S(n611), .Z(n202) );
  MUX2_X1 U806 ( .A(n202), .B(n199), .S(n608), .Z(n203) );
  MUX2_X1 U807 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n617), .Z(n204) );
  MUX2_X1 U808 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n617), .Z(n205) );
  MUX2_X1 U809 ( .A(n205), .B(n204), .S(N11), .Z(n206) );
  MUX2_X1 U810 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n617), .Z(n207) );
  MUX2_X1 U811 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n617), .Z(n208) );
  MUX2_X1 U812 ( .A(n208), .B(n207), .S(n610), .Z(n209) );
  MUX2_X1 U813 ( .A(n209), .B(n206), .S(n608), .Z(n210) );
  MUX2_X1 U814 ( .A(n210), .B(n203), .S(N13), .Z(n211) );
  MUX2_X1 U815 ( .A(n211), .B(n196), .S(N14), .Z(N16) );
  MUX2_X1 U816 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n617), .Z(n212) );
  MUX2_X1 U817 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n617), .Z(n213) );
  MUX2_X1 U818 ( .A(n213), .B(n212), .S(n610), .Z(n214) );
  MUX2_X1 U819 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n617), .Z(n215) );
  MUX2_X1 U820 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n617), .Z(n216) );
  MUX2_X1 U821 ( .A(n216), .B(n215), .S(N11), .Z(n217) );
  MUX2_X1 U822 ( .A(n217), .B(n214), .S(n608), .Z(n218) );
  MUX2_X1 U823 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n618), .Z(n219) );
  MUX2_X1 U824 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n618), .Z(n220) );
  MUX2_X1 U825 ( .A(n220), .B(n219), .S(n609), .Z(n221) );
  MUX2_X1 U826 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n618), .Z(n222) );
  MUX2_X1 U827 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n618), .Z(n223) );
  MUX2_X1 U828 ( .A(n223), .B(n222), .S(N11), .Z(n224) );
  MUX2_X1 U829 ( .A(n224), .B(n221), .S(n608), .Z(n225) );
  MUX2_X1 U830 ( .A(n225), .B(n218), .S(N13), .Z(n226) );
  MUX2_X1 U831 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n618), .Z(n227) );
  MUX2_X1 U832 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n618), .Z(n228) );
  MUX2_X1 U833 ( .A(n228), .B(n227), .S(n610), .Z(n229) );
  MUX2_X1 U834 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n618), .Z(n595) );
  MUX2_X1 U835 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n618), .Z(n596) );
  MUX2_X1 U836 ( .A(n596), .B(n595), .S(n610), .Z(n597) );
  MUX2_X1 U837 ( .A(n597), .B(n229), .S(n608), .Z(n598) );
  MUX2_X1 U838 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n618), .Z(n599) );
  MUX2_X1 U839 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n618), .Z(n600) );
  MUX2_X1 U840 ( .A(n600), .B(n599), .S(n610), .Z(n601) );
  MUX2_X1 U841 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n618), .Z(n602) );
  MUX2_X1 U842 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n618), .Z(n603) );
  MUX2_X1 U843 ( .A(n603), .B(n602), .S(n611), .Z(n604) );
  MUX2_X1 U844 ( .A(n604), .B(n601), .S(n608), .Z(n605) );
  MUX2_X1 U845 ( .A(n605), .B(n598), .S(N13), .Z(n606) );
  MUX2_X1 U846 ( .A(n606), .B(n226), .S(N14), .Z(N15) );
  CLKBUF_X1 U847 ( .A(N11), .Z(n609) );
  INV_X1 U848 ( .A(N10), .ZN(n620) );
  INV_X1 U849 ( .A(N11), .ZN(n621) );
  INV_X1 U850 ( .A(data_in[0]), .ZN(n622) );
  INV_X1 U851 ( .A(data_in[1]), .ZN(n623) );
  INV_X1 U852 ( .A(data_in[2]), .ZN(n624) );
  INV_X1 U853 ( .A(data_in[3]), .ZN(n625) );
  INV_X1 U854 ( .A(data_in[4]), .ZN(n626) );
  INV_X1 U855 ( .A(data_in[5]), .ZN(n627) );
  INV_X1 U856 ( .A(data_in[6]), .ZN(n628) );
  INV_X1 U857 ( .A(data_in[7]), .ZN(n629) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_24 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n628), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n629), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n630), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n631), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n632), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n633), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n634), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n635), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n636), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n637), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n638), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n639), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n640), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n641), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n642), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n643), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n644), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n645), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n646), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n647), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n648), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n649), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n650), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n651), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n652), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n653), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n654), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n655), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n656), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n657), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n658), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n659), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n660), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n661), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n662), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n663), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n664), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n665), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n666), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n667), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n668), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n669), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n670), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n671), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n672), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n673), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n674), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n675), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n676), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n677), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n678), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n679), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n680), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n681), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n682), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n683), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n684), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n685), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n686), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n687), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n688), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n689), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n690), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n691), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n692), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n693), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n694), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n695), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n696), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n697), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n698), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n699), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n700), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n701), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n702), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n703), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n704), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n705), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n706), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n707), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n708), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n709), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n710), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n711), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n712), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n713), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n714), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n715), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n716), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n717), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n718), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n719), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n720), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n721), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n722), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n723), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n724), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n725), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n726), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n727), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n728), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n729), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n730), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n731), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n732), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n733), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n734), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n735), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n736), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n737), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n738), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n739), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n740), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n741), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n742), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n743), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n744), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n745), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n746), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n747), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n748), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n749), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n750), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n751), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n752), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n753), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n754), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n755), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n756), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n757), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n758), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n759), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n760), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n761), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n762), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n763), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n764), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n765), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n766), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n767), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n768), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n769), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n770), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n771), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n772), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n773), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n774), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n775), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n776), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n777), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n778), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n779), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n780), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n781), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n782), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n783), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n784), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n785), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n786), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n787), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n788), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n789), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n790), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n791), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n792), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n793), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n794), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n795), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n796), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n797), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n798), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n799), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n800), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n801), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n802), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n803), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n804), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n805), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n806), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n807), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n808), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n809), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n810), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n811), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n812), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n813), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n814), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n815), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n816), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n817), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n818), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n819), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n847), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n848), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n849), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n850), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n851), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n852), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n853), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n854), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n855), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n856), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n857), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n858), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n859), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n860), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n861), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n862), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n863), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n864), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n865), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n866), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n867), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n868), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n869), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n870), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n871), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n872), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n873), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n874), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n875), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n876), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n877), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n878), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n879), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n880), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n881), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n882), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n883), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n884), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n885), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n886), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n887), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n888), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n889), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n890), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n891), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n892), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n893), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n894), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n895), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n896), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n897), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n898), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n899), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n900), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n901), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n902), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n903), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n904), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n905), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n906), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n907), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n908), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n909), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n910), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n617), .Z(n616) );
  BUF_X1 U4 ( .A(n617), .Z(n613) );
  BUF_X1 U5 ( .A(N10), .Z(n614) );
  BUF_X1 U6 ( .A(n617), .Z(n615) );
  BUF_X1 U7 ( .A(n617), .Z(n612) );
  BUF_X1 U8 ( .A(N11), .Z(n610) );
  BUF_X1 U9 ( .A(N11), .Z(n611) );
  BUF_X1 U10 ( .A(N10), .Z(n617) );
  NOR3_X1 U11 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1202) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(n618), .ZN(n1191) );
  NOR3_X1 U13 ( .A1(N10), .A2(N12), .A3(n619), .ZN(n1181) );
  NOR3_X1 U14 ( .A1(n618), .A2(N12), .A3(n619), .ZN(n1171) );
  INV_X1 U15 ( .A(n1128), .ZN(n843) );
  INV_X1 U16 ( .A(n1118), .ZN(n842) );
  INV_X1 U17 ( .A(n1109), .ZN(n841) );
  INV_X1 U18 ( .A(n1100), .ZN(n840) );
  INV_X1 U19 ( .A(n1055), .ZN(n835) );
  INV_X1 U20 ( .A(n1045), .ZN(n834) );
  INV_X1 U21 ( .A(n1036), .ZN(n833) );
  INV_X1 U22 ( .A(n1027), .ZN(n832) );
  INV_X1 U23 ( .A(n982), .ZN(n827) );
  INV_X1 U24 ( .A(n972), .ZN(n826) );
  INV_X1 U25 ( .A(n963), .ZN(n825) );
  INV_X1 U26 ( .A(n954), .ZN(n824) );
  INV_X1 U27 ( .A(n1091), .ZN(n839) );
  INV_X1 U28 ( .A(n1082), .ZN(n838) );
  INV_X1 U29 ( .A(n1073), .ZN(n837) );
  INV_X1 U30 ( .A(n1064), .ZN(n836) );
  INV_X1 U31 ( .A(n945), .ZN(n823) );
  INV_X1 U32 ( .A(n936), .ZN(n822) );
  INV_X1 U33 ( .A(n927), .ZN(n821) );
  INV_X1 U34 ( .A(n918), .ZN(n820) );
  INV_X1 U35 ( .A(n1018), .ZN(n831) );
  INV_X1 U36 ( .A(n1009), .ZN(n830) );
  INV_X1 U37 ( .A(n1000), .ZN(n829) );
  INV_X1 U38 ( .A(n991), .ZN(n828) );
  BUF_X1 U39 ( .A(N12), .Z(n608) );
  INV_X1 U40 ( .A(N13), .ZN(n845) );
  AND3_X1 U41 ( .A1(n618), .A2(n619), .A3(N12), .ZN(n1161) );
  AND3_X1 U42 ( .A1(N10), .A2(n619), .A3(N12), .ZN(n1151) );
  AND3_X1 U43 ( .A1(N11), .A2(n618), .A3(N12), .ZN(n1141) );
  AND3_X1 U44 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1131) );
  BUF_X1 U45 ( .A(N12), .Z(n607) );
  INV_X1 U46 ( .A(N14), .ZN(n846) );
  NAND2_X1 U47 ( .A1(n1191), .A2(n1201), .ZN(n1200) );
  NAND2_X1 U48 ( .A1(n1181), .A2(n1201), .ZN(n1190) );
  NAND2_X1 U49 ( .A1(n1171), .A2(n1201), .ZN(n1180) );
  NAND2_X1 U50 ( .A1(n1161), .A2(n1201), .ZN(n1170) );
  NAND2_X1 U51 ( .A1(n1151), .A2(n1201), .ZN(n1160) );
  NAND2_X1 U52 ( .A1(n1141), .A2(n1201), .ZN(n1150) );
  NAND2_X1 U53 ( .A1(n1131), .A2(n1201), .ZN(n1140) );
  NAND2_X1 U54 ( .A1(n1202), .A2(n1201), .ZN(n1211) );
  NAND2_X1 U55 ( .A1(n1120), .A2(n1202), .ZN(n1128) );
  NAND2_X1 U56 ( .A1(n1120), .A2(n1191), .ZN(n1118) );
  NAND2_X1 U57 ( .A1(n1120), .A2(n1181), .ZN(n1109) );
  NAND2_X1 U58 ( .A1(n1120), .A2(n1171), .ZN(n1100) );
  NAND2_X1 U59 ( .A1(n1047), .A2(n1202), .ZN(n1055) );
  NAND2_X1 U60 ( .A1(n1047), .A2(n1191), .ZN(n1045) );
  NAND2_X1 U61 ( .A1(n1047), .A2(n1181), .ZN(n1036) );
  NAND2_X1 U62 ( .A1(n1047), .A2(n1171), .ZN(n1027) );
  NAND2_X1 U63 ( .A1(n974), .A2(n1202), .ZN(n982) );
  NAND2_X1 U64 ( .A1(n974), .A2(n1191), .ZN(n972) );
  NAND2_X1 U65 ( .A1(n974), .A2(n1181), .ZN(n963) );
  NAND2_X1 U66 ( .A1(n974), .A2(n1171), .ZN(n954) );
  NAND2_X1 U67 ( .A1(n1120), .A2(n1161), .ZN(n1091) );
  NAND2_X1 U68 ( .A1(n1120), .A2(n1151), .ZN(n1082) );
  NAND2_X1 U69 ( .A1(n1120), .A2(n1141), .ZN(n1073) );
  NAND2_X1 U70 ( .A1(n1120), .A2(n1131), .ZN(n1064) );
  NAND2_X1 U71 ( .A1(n1047), .A2(n1161), .ZN(n1018) );
  NAND2_X1 U72 ( .A1(n1047), .A2(n1151), .ZN(n1009) );
  NAND2_X1 U73 ( .A1(n1047), .A2(n1141), .ZN(n1000) );
  NAND2_X1 U74 ( .A1(n1047), .A2(n1131), .ZN(n991) );
  NAND2_X1 U75 ( .A1(n974), .A2(n1161), .ZN(n945) );
  NAND2_X1 U76 ( .A1(n974), .A2(n1151), .ZN(n936) );
  NAND2_X1 U77 ( .A1(n974), .A2(n1141), .ZN(n927) );
  NAND2_X1 U78 ( .A1(n974), .A2(n1131), .ZN(n918) );
  AND3_X1 U79 ( .A1(n845), .A2(n846), .A3(n1130), .ZN(n1201) );
  AND3_X1 U80 ( .A1(N13), .A2(n1130), .A3(N14), .ZN(n974) );
  AND3_X1 U81 ( .A1(n1130), .A2(n846), .A3(N13), .ZN(n1120) );
  AND3_X1 U82 ( .A1(n1130), .A2(n845), .A3(N14), .ZN(n1047) );
  NOR2_X1 U83 ( .A1(n844), .A2(addr[5]), .ZN(n1130) );
  INV_X1 U84 ( .A(wr_en), .ZN(n844) );
  OAI21_X1 U85 ( .B1(n620), .B2(n1170), .A(n1169), .ZN(n878) );
  NAND2_X1 U86 ( .A1(\mem[4][0] ), .A2(n1170), .ZN(n1169) );
  OAI21_X1 U87 ( .B1(n621), .B2(n1170), .A(n1168), .ZN(n877) );
  NAND2_X1 U88 ( .A1(\mem[4][1] ), .A2(n1170), .ZN(n1168) );
  OAI21_X1 U89 ( .B1(n622), .B2(n1170), .A(n1167), .ZN(n876) );
  NAND2_X1 U90 ( .A1(\mem[4][2] ), .A2(n1170), .ZN(n1167) );
  OAI21_X1 U91 ( .B1(n623), .B2(n1170), .A(n1166), .ZN(n875) );
  NAND2_X1 U92 ( .A1(\mem[4][3] ), .A2(n1170), .ZN(n1166) );
  OAI21_X1 U93 ( .B1(n624), .B2(n1170), .A(n1165), .ZN(n874) );
  NAND2_X1 U94 ( .A1(\mem[4][4] ), .A2(n1170), .ZN(n1165) );
  OAI21_X1 U95 ( .B1(n625), .B2(n1170), .A(n1164), .ZN(n873) );
  NAND2_X1 U96 ( .A1(\mem[4][5] ), .A2(n1170), .ZN(n1164) );
  OAI21_X1 U97 ( .B1(n626), .B2(n1170), .A(n1163), .ZN(n872) );
  NAND2_X1 U98 ( .A1(\mem[4][6] ), .A2(n1170), .ZN(n1163) );
  OAI21_X1 U99 ( .B1(n627), .B2(n1170), .A(n1162), .ZN(n871) );
  NAND2_X1 U100 ( .A1(\mem[4][7] ), .A2(n1170), .ZN(n1162) );
  OAI21_X1 U101 ( .B1(n620), .B2(n1150), .A(n1149), .ZN(n862) );
  NAND2_X1 U102 ( .A1(\mem[6][0] ), .A2(n1150), .ZN(n1149) );
  OAI21_X1 U103 ( .B1(n621), .B2(n1150), .A(n1148), .ZN(n861) );
  NAND2_X1 U104 ( .A1(\mem[6][1] ), .A2(n1150), .ZN(n1148) );
  OAI21_X1 U105 ( .B1(n622), .B2(n1150), .A(n1147), .ZN(n860) );
  NAND2_X1 U106 ( .A1(\mem[6][2] ), .A2(n1150), .ZN(n1147) );
  OAI21_X1 U107 ( .B1(n623), .B2(n1150), .A(n1146), .ZN(n859) );
  NAND2_X1 U108 ( .A1(\mem[6][3] ), .A2(n1150), .ZN(n1146) );
  OAI21_X1 U109 ( .B1(n624), .B2(n1150), .A(n1145), .ZN(n858) );
  NAND2_X1 U110 ( .A1(\mem[6][4] ), .A2(n1150), .ZN(n1145) );
  OAI21_X1 U111 ( .B1(n625), .B2(n1150), .A(n1144), .ZN(n857) );
  NAND2_X1 U112 ( .A1(\mem[6][5] ), .A2(n1150), .ZN(n1144) );
  OAI21_X1 U113 ( .B1(n626), .B2(n1150), .A(n1143), .ZN(n856) );
  NAND2_X1 U114 ( .A1(\mem[6][6] ), .A2(n1150), .ZN(n1143) );
  OAI21_X1 U115 ( .B1(n627), .B2(n1150), .A(n1142), .ZN(n855) );
  NAND2_X1 U116 ( .A1(\mem[6][7] ), .A2(n1150), .ZN(n1142) );
  OAI21_X1 U117 ( .B1(n620), .B2(n1140), .A(n1139), .ZN(n854) );
  NAND2_X1 U118 ( .A1(\mem[7][0] ), .A2(n1140), .ZN(n1139) );
  OAI21_X1 U119 ( .B1(n621), .B2(n1140), .A(n1138), .ZN(n853) );
  NAND2_X1 U120 ( .A1(\mem[7][1] ), .A2(n1140), .ZN(n1138) );
  OAI21_X1 U121 ( .B1(n622), .B2(n1140), .A(n1137), .ZN(n852) );
  NAND2_X1 U122 ( .A1(\mem[7][2] ), .A2(n1140), .ZN(n1137) );
  OAI21_X1 U123 ( .B1(n623), .B2(n1140), .A(n1136), .ZN(n851) );
  NAND2_X1 U124 ( .A1(\mem[7][3] ), .A2(n1140), .ZN(n1136) );
  OAI21_X1 U125 ( .B1(n624), .B2(n1140), .A(n1135), .ZN(n850) );
  NAND2_X1 U126 ( .A1(\mem[7][4] ), .A2(n1140), .ZN(n1135) );
  OAI21_X1 U127 ( .B1(n625), .B2(n1140), .A(n1134), .ZN(n849) );
  NAND2_X1 U128 ( .A1(\mem[7][5] ), .A2(n1140), .ZN(n1134) );
  OAI21_X1 U129 ( .B1(n626), .B2(n1140), .A(n1133), .ZN(n848) );
  NAND2_X1 U130 ( .A1(\mem[7][6] ), .A2(n1140), .ZN(n1133) );
  OAI21_X1 U131 ( .B1(n627), .B2(n1140), .A(n1132), .ZN(n847) );
  NAND2_X1 U132 ( .A1(\mem[7][7] ), .A2(n1140), .ZN(n1132) );
  OAI21_X1 U133 ( .B1(n620), .B2(n1200), .A(n1199), .ZN(n902) );
  NAND2_X1 U134 ( .A1(\mem[1][0] ), .A2(n1200), .ZN(n1199) );
  OAI21_X1 U135 ( .B1(n621), .B2(n1200), .A(n1198), .ZN(n901) );
  NAND2_X1 U136 ( .A1(\mem[1][1] ), .A2(n1200), .ZN(n1198) );
  OAI21_X1 U137 ( .B1(n622), .B2(n1200), .A(n1197), .ZN(n900) );
  NAND2_X1 U138 ( .A1(\mem[1][2] ), .A2(n1200), .ZN(n1197) );
  OAI21_X1 U139 ( .B1(n623), .B2(n1200), .A(n1196), .ZN(n899) );
  NAND2_X1 U140 ( .A1(\mem[1][3] ), .A2(n1200), .ZN(n1196) );
  OAI21_X1 U141 ( .B1(n624), .B2(n1200), .A(n1195), .ZN(n898) );
  NAND2_X1 U142 ( .A1(\mem[1][4] ), .A2(n1200), .ZN(n1195) );
  OAI21_X1 U143 ( .B1(n625), .B2(n1200), .A(n1194), .ZN(n897) );
  NAND2_X1 U144 ( .A1(\mem[1][5] ), .A2(n1200), .ZN(n1194) );
  OAI21_X1 U145 ( .B1(n626), .B2(n1200), .A(n1193), .ZN(n896) );
  NAND2_X1 U146 ( .A1(\mem[1][6] ), .A2(n1200), .ZN(n1193) );
  OAI21_X1 U147 ( .B1(n627), .B2(n1200), .A(n1192), .ZN(n895) );
  NAND2_X1 U148 ( .A1(\mem[1][7] ), .A2(n1200), .ZN(n1192) );
  OAI21_X1 U149 ( .B1(n620), .B2(n1190), .A(n1189), .ZN(n894) );
  NAND2_X1 U150 ( .A1(\mem[2][0] ), .A2(n1190), .ZN(n1189) );
  OAI21_X1 U151 ( .B1(n621), .B2(n1190), .A(n1188), .ZN(n893) );
  NAND2_X1 U152 ( .A1(\mem[2][1] ), .A2(n1190), .ZN(n1188) );
  OAI21_X1 U153 ( .B1(n622), .B2(n1190), .A(n1187), .ZN(n892) );
  NAND2_X1 U154 ( .A1(\mem[2][2] ), .A2(n1190), .ZN(n1187) );
  OAI21_X1 U155 ( .B1(n623), .B2(n1190), .A(n1186), .ZN(n891) );
  NAND2_X1 U156 ( .A1(\mem[2][3] ), .A2(n1190), .ZN(n1186) );
  OAI21_X1 U157 ( .B1(n624), .B2(n1190), .A(n1185), .ZN(n890) );
  NAND2_X1 U158 ( .A1(\mem[2][4] ), .A2(n1190), .ZN(n1185) );
  OAI21_X1 U159 ( .B1(n625), .B2(n1190), .A(n1184), .ZN(n889) );
  NAND2_X1 U160 ( .A1(\mem[2][5] ), .A2(n1190), .ZN(n1184) );
  OAI21_X1 U161 ( .B1(n626), .B2(n1190), .A(n1183), .ZN(n888) );
  NAND2_X1 U162 ( .A1(\mem[2][6] ), .A2(n1190), .ZN(n1183) );
  OAI21_X1 U163 ( .B1(n627), .B2(n1190), .A(n1182), .ZN(n887) );
  NAND2_X1 U164 ( .A1(\mem[2][7] ), .A2(n1190), .ZN(n1182) );
  OAI21_X1 U165 ( .B1(n620), .B2(n1180), .A(n1179), .ZN(n886) );
  NAND2_X1 U166 ( .A1(\mem[3][0] ), .A2(n1180), .ZN(n1179) );
  OAI21_X1 U167 ( .B1(n621), .B2(n1180), .A(n1178), .ZN(n885) );
  NAND2_X1 U168 ( .A1(\mem[3][1] ), .A2(n1180), .ZN(n1178) );
  OAI21_X1 U169 ( .B1(n622), .B2(n1180), .A(n1177), .ZN(n884) );
  NAND2_X1 U170 ( .A1(\mem[3][2] ), .A2(n1180), .ZN(n1177) );
  OAI21_X1 U171 ( .B1(n623), .B2(n1180), .A(n1176), .ZN(n883) );
  NAND2_X1 U172 ( .A1(\mem[3][3] ), .A2(n1180), .ZN(n1176) );
  OAI21_X1 U173 ( .B1(n624), .B2(n1180), .A(n1175), .ZN(n882) );
  NAND2_X1 U174 ( .A1(\mem[3][4] ), .A2(n1180), .ZN(n1175) );
  OAI21_X1 U175 ( .B1(n625), .B2(n1180), .A(n1174), .ZN(n881) );
  NAND2_X1 U176 ( .A1(\mem[3][5] ), .A2(n1180), .ZN(n1174) );
  OAI21_X1 U177 ( .B1(n626), .B2(n1180), .A(n1173), .ZN(n880) );
  NAND2_X1 U178 ( .A1(\mem[3][6] ), .A2(n1180), .ZN(n1173) );
  OAI21_X1 U179 ( .B1(n627), .B2(n1180), .A(n1172), .ZN(n879) );
  NAND2_X1 U180 ( .A1(\mem[3][7] ), .A2(n1180), .ZN(n1172) );
  OAI21_X1 U181 ( .B1(n620), .B2(n1160), .A(n1159), .ZN(n870) );
  NAND2_X1 U182 ( .A1(\mem[5][0] ), .A2(n1160), .ZN(n1159) );
  OAI21_X1 U183 ( .B1(n621), .B2(n1160), .A(n1158), .ZN(n869) );
  NAND2_X1 U184 ( .A1(\mem[5][1] ), .A2(n1160), .ZN(n1158) );
  OAI21_X1 U185 ( .B1(n622), .B2(n1160), .A(n1157), .ZN(n868) );
  NAND2_X1 U186 ( .A1(\mem[5][2] ), .A2(n1160), .ZN(n1157) );
  OAI21_X1 U187 ( .B1(n623), .B2(n1160), .A(n1156), .ZN(n867) );
  NAND2_X1 U188 ( .A1(\mem[5][3] ), .A2(n1160), .ZN(n1156) );
  OAI21_X1 U189 ( .B1(n624), .B2(n1160), .A(n1155), .ZN(n866) );
  NAND2_X1 U190 ( .A1(\mem[5][4] ), .A2(n1160), .ZN(n1155) );
  OAI21_X1 U191 ( .B1(n625), .B2(n1160), .A(n1154), .ZN(n865) );
  NAND2_X1 U192 ( .A1(\mem[5][5] ), .A2(n1160), .ZN(n1154) );
  OAI21_X1 U193 ( .B1(n626), .B2(n1160), .A(n1153), .ZN(n864) );
  NAND2_X1 U194 ( .A1(\mem[5][6] ), .A2(n1160), .ZN(n1153) );
  OAI21_X1 U195 ( .B1(n627), .B2(n1160), .A(n1152), .ZN(n863) );
  NAND2_X1 U196 ( .A1(\mem[5][7] ), .A2(n1160), .ZN(n1152) );
  OAI21_X1 U197 ( .B1(n1211), .B2(n620), .A(n1210), .ZN(n910) );
  NAND2_X1 U198 ( .A1(\mem[0][0] ), .A2(n1211), .ZN(n1210) );
  OAI21_X1 U199 ( .B1(n1211), .B2(n621), .A(n1209), .ZN(n909) );
  NAND2_X1 U200 ( .A1(\mem[0][1] ), .A2(n1211), .ZN(n1209) );
  OAI21_X1 U201 ( .B1(n1211), .B2(n622), .A(n1208), .ZN(n908) );
  NAND2_X1 U202 ( .A1(\mem[0][2] ), .A2(n1211), .ZN(n1208) );
  OAI21_X1 U203 ( .B1(n1211), .B2(n623), .A(n1207), .ZN(n907) );
  NAND2_X1 U204 ( .A1(\mem[0][3] ), .A2(n1211), .ZN(n1207) );
  OAI21_X1 U205 ( .B1(n1211), .B2(n624), .A(n1206), .ZN(n906) );
  NAND2_X1 U206 ( .A1(\mem[0][4] ), .A2(n1211), .ZN(n1206) );
  OAI21_X1 U207 ( .B1(n1211), .B2(n625), .A(n1205), .ZN(n905) );
  NAND2_X1 U208 ( .A1(\mem[0][5] ), .A2(n1211), .ZN(n1205) );
  OAI21_X1 U209 ( .B1(n1211), .B2(n626), .A(n1204), .ZN(n904) );
  NAND2_X1 U210 ( .A1(\mem[0][6] ), .A2(n1211), .ZN(n1204) );
  OAI21_X1 U211 ( .B1(n1211), .B2(n627), .A(n1203), .ZN(n903) );
  NAND2_X1 U212 ( .A1(\mem[0][7] ), .A2(n1211), .ZN(n1203) );
  INV_X1 U213 ( .A(n1129), .ZN(n819) );
  AOI22_X1 U214 ( .A1(data_in[0]), .A2(n843), .B1(n1128), .B2(\mem[8][0] ), 
        .ZN(n1129) );
  INV_X1 U215 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U216 ( .A1(data_in[1]), .A2(n843), .B1(n1128), .B2(\mem[8][1] ), 
        .ZN(n1127) );
  INV_X1 U217 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U218 ( .A1(data_in[2]), .A2(n843), .B1(n1128), .B2(\mem[8][2] ), 
        .ZN(n1126) );
  INV_X1 U219 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U220 ( .A1(data_in[3]), .A2(n843), .B1(n1128), .B2(\mem[8][3] ), 
        .ZN(n1125) );
  INV_X1 U221 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U222 ( .A1(data_in[4]), .A2(n843), .B1(n1128), .B2(\mem[8][4] ), 
        .ZN(n1124) );
  INV_X1 U223 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U224 ( .A1(data_in[5]), .A2(n843), .B1(n1128), .B2(\mem[8][5] ), 
        .ZN(n1123) );
  INV_X1 U225 ( .A(n1122), .ZN(n813) );
  AOI22_X1 U226 ( .A1(data_in[6]), .A2(n843), .B1(n1128), .B2(\mem[8][6] ), 
        .ZN(n1122) );
  INV_X1 U227 ( .A(n1121), .ZN(n812) );
  AOI22_X1 U228 ( .A1(data_in[7]), .A2(n843), .B1(n1128), .B2(\mem[8][7] ), 
        .ZN(n1121) );
  INV_X1 U229 ( .A(n1119), .ZN(n811) );
  AOI22_X1 U230 ( .A1(data_in[0]), .A2(n842), .B1(n1118), .B2(\mem[9][0] ), 
        .ZN(n1119) );
  INV_X1 U231 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U232 ( .A1(data_in[1]), .A2(n842), .B1(n1118), .B2(\mem[9][1] ), 
        .ZN(n1117) );
  INV_X1 U233 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U234 ( .A1(data_in[2]), .A2(n842), .B1(n1118), .B2(\mem[9][2] ), 
        .ZN(n1116) );
  INV_X1 U235 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U236 ( .A1(data_in[3]), .A2(n842), .B1(n1118), .B2(\mem[9][3] ), 
        .ZN(n1115) );
  INV_X1 U237 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U238 ( .A1(data_in[4]), .A2(n842), .B1(n1118), .B2(\mem[9][4] ), 
        .ZN(n1114) );
  INV_X1 U239 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U240 ( .A1(data_in[5]), .A2(n842), .B1(n1118), .B2(\mem[9][5] ), 
        .ZN(n1113) );
  INV_X1 U241 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U242 ( .A1(data_in[6]), .A2(n842), .B1(n1118), .B2(\mem[9][6] ), 
        .ZN(n1112) );
  INV_X1 U243 ( .A(n1111), .ZN(n804) );
  AOI22_X1 U244 ( .A1(data_in[7]), .A2(n842), .B1(n1118), .B2(\mem[9][7] ), 
        .ZN(n1111) );
  INV_X1 U245 ( .A(n1110), .ZN(n803) );
  AOI22_X1 U246 ( .A1(data_in[0]), .A2(n841), .B1(n1109), .B2(\mem[10][0] ), 
        .ZN(n1110) );
  INV_X1 U247 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U248 ( .A1(data_in[1]), .A2(n841), .B1(n1109), .B2(\mem[10][1] ), 
        .ZN(n1108) );
  INV_X1 U249 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U250 ( .A1(data_in[2]), .A2(n841), .B1(n1109), .B2(\mem[10][2] ), 
        .ZN(n1107) );
  INV_X1 U251 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U252 ( .A1(data_in[3]), .A2(n841), .B1(n1109), .B2(\mem[10][3] ), 
        .ZN(n1106) );
  INV_X1 U253 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U254 ( .A1(data_in[4]), .A2(n841), .B1(n1109), .B2(\mem[10][4] ), 
        .ZN(n1105) );
  INV_X1 U255 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U256 ( .A1(data_in[5]), .A2(n841), .B1(n1109), .B2(\mem[10][5] ), 
        .ZN(n1104) );
  INV_X1 U257 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U258 ( .A1(data_in[6]), .A2(n841), .B1(n1109), .B2(\mem[10][6] ), 
        .ZN(n1103) );
  INV_X1 U259 ( .A(n1102), .ZN(n796) );
  AOI22_X1 U260 ( .A1(data_in[7]), .A2(n841), .B1(n1109), .B2(\mem[10][7] ), 
        .ZN(n1102) );
  INV_X1 U261 ( .A(n1101), .ZN(n795) );
  AOI22_X1 U262 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[11][0] ), 
        .ZN(n1101) );
  INV_X1 U263 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U264 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[11][1] ), 
        .ZN(n1099) );
  INV_X1 U265 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U266 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[11][2] ), 
        .ZN(n1098) );
  INV_X1 U267 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U268 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[11][3] ), 
        .ZN(n1097) );
  INV_X1 U269 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U270 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[11][4] ), 
        .ZN(n1096) );
  INV_X1 U271 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U272 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[11][5] ), 
        .ZN(n1095) );
  INV_X1 U273 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U274 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[11][6] ), 
        .ZN(n1094) );
  INV_X1 U275 ( .A(n1093), .ZN(n788) );
  AOI22_X1 U276 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[11][7] ), 
        .ZN(n1093) );
  INV_X1 U277 ( .A(n1092), .ZN(n787) );
  AOI22_X1 U278 ( .A1(data_in[0]), .A2(n839), .B1(n1091), .B2(\mem[12][0] ), 
        .ZN(n1092) );
  INV_X1 U279 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U280 ( .A1(data_in[1]), .A2(n839), .B1(n1091), .B2(\mem[12][1] ), 
        .ZN(n1090) );
  INV_X1 U281 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U282 ( .A1(data_in[2]), .A2(n839), .B1(n1091), .B2(\mem[12][2] ), 
        .ZN(n1089) );
  INV_X1 U283 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U284 ( .A1(data_in[3]), .A2(n839), .B1(n1091), .B2(\mem[12][3] ), 
        .ZN(n1088) );
  INV_X1 U285 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U286 ( .A1(data_in[4]), .A2(n839), .B1(n1091), .B2(\mem[12][4] ), 
        .ZN(n1087) );
  INV_X1 U287 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U288 ( .A1(data_in[5]), .A2(n839), .B1(n1091), .B2(\mem[12][5] ), 
        .ZN(n1086) );
  INV_X1 U289 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U290 ( .A1(data_in[6]), .A2(n839), .B1(n1091), .B2(\mem[12][6] ), 
        .ZN(n1085) );
  INV_X1 U291 ( .A(n1084), .ZN(n780) );
  AOI22_X1 U292 ( .A1(data_in[7]), .A2(n839), .B1(n1091), .B2(\mem[12][7] ), 
        .ZN(n1084) );
  INV_X1 U293 ( .A(n1083), .ZN(n779) );
  AOI22_X1 U294 ( .A1(data_in[0]), .A2(n838), .B1(n1082), .B2(\mem[13][0] ), 
        .ZN(n1083) );
  INV_X1 U295 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U296 ( .A1(data_in[1]), .A2(n838), .B1(n1082), .B2(\mem[13][1] ), 
        .ZN(n1081) );
  INV_X1 U297 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U298 ( .A1(data_in[2]), .A2(n838), .B1(n1082), .B2(\mem[13][2] ), 
        .ZN(n1080) );
  INV_X1 U299 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U300 ( .A1(data_in[3]), .A2(n838), .B1(n1082), .B2(\mem[13][3] ), 
        .ZN(n1079) );
  INV_X1 U301 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U302 ( .A1(data_in[4]), .A2(n838), .B1(n1082), .B2(\mem[13][4] ), 
        .ZN(n1078) );
  INV_X1 U303 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U304 ( .A1(data_in[5]), .A2(n838), .B1(n1082), .B2(\mem[13][5] ), 
        .ZN(n1077) );
  INV_X1 U305 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U306 ( .A1(data_in[6]), .A2(n838), .B1(n1082), .B2(\mem[13][6] ), 
        .ZN(n1076) );
  INV_X1 U307 ( .A(n1075), .ZN(n772) );
  AOI22_X1 U308 ( .A1(data_in[7]), .A2(n838), .B1(n1082), .B2(\mem[13][7] ), 
        .ZN(n1075) );
  INV_X1 U309 ( .A(n1074), .ZN(n771) );
  AOI22_X1 U310 ( .A1(data_in[0]), .A2(n837), .B1(n1073), .B2(\mem[14][0] ), 
        .ZN(n1074) );
  INV_X1 U311 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U312 ( .A1(data_in[1]), .A2(n837), .B1(n1073), .B2(\mem[14][1] ), 
        .ZN(n1072) );
  INV_X1 U313 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U314 ( .A1(data_in[2]), .A2(n837), .B1(n1073), .B2(\mem[14][2] ), 
        .ZN(n1071) );
  INV_X1 U315 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U316 ( .A1(data_in[3]), .A2(n837), .B1(n1073), .B2(\mem[14][3] ), 
        .ZN(n1070) );
  INV_X1 U317 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U318 ( .A1(data_in[4]), .A2(n837), .B1(n1073), .B2(\mem[14][4] ), 
        .ZN(n1069) );
  INV_X1 U319 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U320 ( .A1(data_in[5]), .A2(n837), .B1(n1073), .B2(\mem[14][5] ), 
        .ZN(n1068) );
  INV_X1 U321 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U322 ( .A1(data_in[6]), .A2(n837), .B1(n1073), .B2(\mem[14][6] ), 
        .ZN(n1067) );
  INV_X1 U323 ( .A(n1066), .ZN(n764) );
  AOI22_X1 U324 ( .A1(data_in[7]), .A2(n837), .B1(n1073), .B2(\mem[14][7] ), 
        .ZN(n1066) );
  INV_X1 U325 ( .A(n1065), .ZN(n763) );
  AOI22_X1 U326 ( .A1(data_in[0]), .A2(n836), .B1(n1064), .B2(\mem[15][0] ), 
        .ZN(n1065) );
  INV_X1 U327 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U328 ( .A1(data_in[1]), .A2(n836), .B1(n1064), .B2(\mem[15][1] ), 
        .ZN(n1063) );
  INV_X1 U329 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U330 ( .A1(data_in[2]), .A2(n836), .B1(n1064), .B2(\mem[15][2] ), 
        .ZN(n1062) );
  INV_X1 U331 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U332 ( .A1(data_in[3]), .A2(n836), .B1(n1064), .B2(\mem[15][3] ), 
        .ZN(n1061) );
  INV_X1 U333 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U334 ( .A1(data_in[4]), .A2(n836), .B1(n1064), .B2(\mem[15][4] ), 
        .ZN(n1060) );
  INV_X1 U335 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U336 ( .A1(data_in[5]), .A2(n836), .B1(n1064), .B2(\mem[15][5] ), 
        .ZN(n1059) );
  INV_X1 U337 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U338 ( .A1(data_in[6]), .A2(n836), .B1(n1064), .B2(\mem[15][6] ), 
        .ZN(n1058) );
  INV_X1 U339 ( .A(n1057), .ZN(n756) );
  AOI22_X1 U340 ( .A1(data_in[7]), .A2(n836), .B1(n1064), .B2(\mem[15][7] ), 
        .ZN(n1057) );
  INV_X1 U341 ( .A(n1056), .ZN(n755) );
  AOI22_X1 U342 ( .A1(data_in[0]), .A2(n835), .B1(n1055), .B2(\mem[16][0] ), 
        .ZN(n1056) );
  INV_X1 U343 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U344 ( .A1(data_in[1]), .A2(n835), .B1(n1055), .B2(\mem[16][1] ), 
        .ZN(n1054) );
  INV_X1 U345 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U346 ( .A1(data_in[2]), .A2(n835), .B1(n1055), .B2(\mem[16][2] ), 
        .ZN(n1053) );
  INV_X1 U347 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U348 ( .A1(data_in[3]), .A2(n835), .B1(n1055), .B2(\mem[16][3] ), 
        .ZN(n1052) );
  INV_X1 U349 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U350 ( .A1(data_in[4]), .A2(n835), .B1(n1055), .B2(\mem[16][4] ), 
        .ZN(n1051) );
  INV_X1 U351 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U352 ( .A1(data_in[5]), .A2(n835), .B1(n1055), .B2(\mem[16][5] ), 
        .ZN(n1050) );
  INV_X1 U353 ( .A(n1049), .ZN(n749) );
  AOI22_X1 U354 ( .A1(data_in[6]), .A2(n835), .B1(n1055), .B2(\mem[16][6] ), 
        .ZN(n1049) );
  INV_X1 U355 ( .A(n1048), .ZN(n748) );
  AOI22_X1 U356 ( .A1(data_in[7]), .A2(n835), .B1(n1055), .B2(\mem[16][7] ), 
        .ZN(n1048) );
  INV_X1 U357 ( .A(n1046), .ZN(n747) );
  AOI22_X1 U358 ( .A1(data_in[0]), .A2(n834), .B1(n1045), .B2(\mem[17][0] ), 
        .ZN(n1046) );
  INV_X1 U359 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U360 ( .A1(data_in[1]), .A2(n834), .B1(n1045), .B2(\mem[17][1] ), 
        .ZN(n1044) );
  INV_X1 U361 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U362 ( .A1(data_in[2]), .A2(n834), .B1(n1045), .B2(\mem[17][2] ), 
        .ZN(n1043) );
  INV_X1 U363 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U364 ( .A1(data_in[3]), .A2(n834), .B1(n1045), .B2(\mem[17][3] ), 
        .ZN(n1042) );
  INV_X1 U365 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U366 ( .A1(data_in[4]), .A2(n834), .B1(n1045), .B2(\mem[17][4] ), 
        .ZN(n1041) );
  INV_X1 U367 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U368 ( .A1(data_in[5]), .A2(n834), .B1(n1045), .B2(\mem[17][5] ), 
        .ZN(n1040) );
  INV_X1 U369 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U370 ( .A1(data_in[6]), .A2(n834), .B1(n1045), .B2(\mem[17][6] ), 
        .ZN(n1039) );
  INV_X1 U371 ( .A(n1038), .ZN(n740) );
  AOI22_X1 U372 ( .A1(data_in[7]), .A2(n834), .B1(n1045), .B2(\mem[17][7] ), 
        .ZN(n1038) );
  INV_X1 U373 ( .A(n1037), .ZN(n739) );
  AOI22_X1 U374 ( .A1(data_in[0]), .A2(n833), .B1(n1036), .B2(\mem[18][0] ), 
        .ZN(n1037) );
  INV_X1 U375 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U376 ( .A1(data_in[1]), .A2(n833), .B1(n1036), .B2(\mem[18][1] ), 
        .ZN(n1035) );
  INV_X1 U377 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U378 ( .A1(data_in[2]), .A2(n833), .B1(n1036), .B2(\mem[18][2] ), 
        .ZN(n1034) );
  INV_X1 U379 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U380 ( .A1(data_in[3]), .A2(n833), .B1(n1036), .B2(\mem[18][3] ), 
        .ZN(n1033) );
  INV_X1 U381 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U382 ( .A1(data_in[4]), .A2(n833), .B1(n1036), .B2(\mem[18][4] ), 
        .ZN(n1032) );
  INV_X1 U383 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U384 ( .A1(data_in[5]), .A2(n833), .B1(n1036), .B2(\mem[18][5] ), 
        .ZN(n1031) );
  INV_X1 U385 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U386 ( .A1(data_in[6]), .A2(n833), .B1(n1036), .B2(\mem[18][6] ), 
        .ZN(n1030) );
  INV_X1 U387 ( .A(n1029), .ZN(n732) );
  AOI22_X1 U388 ( .A1(data_in[7]), .A2(n833), .B1(n1036), .B2(\mem[18][7] ), 
        .ZN(n1029) );
  INV_X1 U389 ( .A(n1028), .ZN(n731) );
  AOI22_X1 U390 ( .A1(data_in[0]), .A2(n832), .B1(n1027), .B2(\mem[19][0] ), 
        .ZN(n1028) );
  INV_X1 U391 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U392 ( .A1(data_in[1]), .A2(n832), .B1(n1027), .B2(\mem[19][1] ), 
        .ZN(n1026) );
  INV_X1 U393 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U394 ( .A1(data_in[2]), .A2(n832), .B1(n1027), .B2(\mem[19][2] ), 
        .ZN(n1025) );
  INV_X1 U395 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U396 ( .A1(data_in[3]), .A2(n832), .B1(n1027), .B2(\mem[19][3] ), 
        .ZN(n1024) );
  INV_X1 U397 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U398 ( .A1(data_in[4]), .A2(n832), .B1(n1027), .B2(\mem[19][4] ), 
        .ZN(n1023) );
  INV_X1 U399 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U400 ( .A1(data_in[5]), .A2(n832), .B1(n1027), .B2(\mem[19][5] ), 
        .ZN(n1022) );
  INV_X1 U401 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U402 ( .A1(data_in[6]), .A2(n832), .B1(n1027), .B2(\mem[19][6] ), 
        .ZN(n1021) );
  INV_X1 U403 ( .A(n1020), .ZN(n724) );
  AOI22_X1 U404 ( .A1(data_in[7]), .A2(n832), .B1(n1027), .B2(\mem[19][7] ), 
        .ZN(n1020) );
  INV_X1 U405 ( .A(n1019), .ZN(n723) );
  AOI22_X1 U406 ( .A1(data_in[0]), .A2(n831), .B1(n1018), .B2(\mem[20][0] ), 
        .ZN(n1019) );
  INV_X1 U407 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U408 ( .A1(data_in[1]), .A2(n831), .B1(n1018), .B2(\mem[20][1] ), 
        .ZN(n1017) );
  INV_X1 U409 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U410 ( .A1(data_in[2]), .A2(n831), .B1(n1018), .B2(\mem[20][2] ), 
        .ZN(n1016) );
  INV_X1 U411 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U412 ( .A1(data_in[3]), .A2(n831), .B1(n1018), .B2(\mem[20][3] ), 
        .ZN(n1015) );
  INV_X1 U413 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U414 ( .A1(data_in[4]), .A2(n831), .B1(n1018), .B2(\mem[20][4] ), 
        .ZN(n1014) );
  INV_X1 U415 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U416 ( .A1(data_in[5]), .A2(n831), .B1(n1018), .B2(\mem[20][5] ), 
        .ZN(n1013) );
  INV_X1 U417 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U418 ( .A1(data_in[6]), .A2(n831), .B1(n1018), .B2(\mem[20][6] ), 
        .ZN(n1012) );
  INV_X1 U419 ( .A(n1011), .ZN(n716) );
  AOI22_X1 U420 ( .A1(data_in[7]), .A2(n831), .B1(n1018), .B2(\mem[20][7] ), 
        .ZN(n1011) );
  INV_X1 U421 ( .A(n1010), .ZN(n715) );
  AOI22_X1 U422 ( .A1(data_in[0]), .A2(n830), .B1(n1009), .B2(\mem[21][0] ), 
        .ZN(n1010) );
  INV_X1 U423 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U424 ( .A1(data_in[1]), .A2(n830), .B1(n1009), .B2(\mem[21][1] ), 
        .ZN(n1008) );
  INV_X1 U425 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U426 ( .A1(data_in[2]), .A2(n830), .B1(n1009), .B2(\mem[21][2] ), 
        .ZN(n1007) );
  INV_X1 U427 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U428 ( .A1(data_in[3]), .A2(n830), .B1(n1009), .B2(\mem[21][3] ), 
        .ZN(n1006) );
  INV_X1 U429 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U430 ( .A1(data_in[4]), .A2(n830), .B1(n1009), .B2(\mem[21][4] ), 
        .ZN(n1005) );
  INV_X1 U431 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U432 ( .A1(data_in[5]), .A2(n830), .B1(n1009), .B2(\mem[21][5] ), 
        .ZN(n1004) );
  INV_X1 U433 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U434 ( .A1(data_in[6]), .A2(n830), .B1(n1009), .B2(\mem[21][6] ), 
        .ZN(n1003) );
  INV_X1 U435 ( .A(n1002), .ZN(n708) );
  AOI22_X1 U436 ( .A1(data_in[7]), .A2(n830), .B1(n1009), .B2(\mem[21][7] ), 
        .ZN(n1002) );
  INV_X1 U437 ( .A(n1001), .ZN(n707) );
  AOI22_X1 U438 ( .A1(data_in[0]), .A2(n829), .B1(n1000), .B2(\mem[22][0] ), 
        .ZN(n1001) );
  INV_X1 U439 ( .A(n999), .ZN(n706) );
  AOI22_X1 U440 ( .A1(data_in[1]), .A2(n829), .B1(n1000), .B2(\mem[22][1] ), 
        .ZN(n999) );
  INV_X1 U441 ( .A(n998), .ZN(n705) );
  AOI22_X1 U442 ( .A1(data_in[2]), .A2(n829), .B1(n1000), .B2(\mem[22][2] ), 
        .ZN(n998) );
  INV_X1 U443 ( .A(n997), .ZN(n704) );
  AOI22_X1 U444 ( .A1(data_in[3]), .A2(n829), .B1(n1000), .B2(\mem[22][3] ), 
        .ZN(n997) );
  INV_X1 U445 ( .A(n996), .ZN(n703) );
  AOI22_X1 U446 ( .A1(data_in[4]), .A2(n829), .B1(n1000), .B2(\mem[22][4] ), 
        .ZN(n996) );
  INV_X1 U447 ( .A(n995), .ZN(n702) );
  AOI22_X1 U448 ( .A1(data_in[5]), .A2(n829), .B1(n1000), .B2(\mem[22][5] ), 
        .ZN(n995) );
  INV_X1 U449 ( .A(n994), .ZN(n701) );
  AOI22_X1 U450 ( .A1(data_in[6]), .A2(n829), .B1(n1000), .B2(\mem[22][6] ), 
        .ZN(n994) );
  INV_X1 U451 ( .A(n993), .ZN(n700) );
  AOI22_X1 U452 ( .A1(data_in[7]), .A2(n829), .B1(n1000), .B2(\mem[22][7] ), 
        .ZN(n993) );
  INV_X1 U453 ( .A(n992), .ZN(n699) );
  AOI22_X1 U454 ( .A1(data_in[0]), .A2(n828), .B1(n991), .B2(\mem[23][0] ), 
        .ZN(n992) );
  INV_X1 U455 ( .A(n990), .ZN(n698) );
  AOI22_X1 U456 ( .A1(data_in[1]), .A2(n828), .B1(n991), .B2(\mem[23][1] ), 
        .ZN(n990) );
  INV_X1 U457 ( .A(n989), .ZN(n697) );
  AOI22_X1 U458 ( .A1(data_in[2]), .A2(n828), .B1(n991), .B2(\mem[23][2] ), 
        .ZN(n989) );
  INV_X1 U459 ( .A(n988), .ZN(n696) );
  AOI22_X1 U460 ( .A1(data_in[3]), .A2(n828), .B1(n991), .B2(\mem[23][3] ), 
        .ZN(n988) );
  INV_X1 U461 ( .A(n987), .ZN(n695) );
  AOI22_X1 U462 ( .A1(data_in[4]), .A2(n828), .B1(n991), .B2(\mem[23][4] ), 
        .ZN(n987) );
  INV_X1 U463 ( .A(n986), .ZN(n694) );
  AOI22_X1 U464 ( .A1(data_in[5]), .A2(n828), .B1(n991), .B2(\mem[23][5] ), 
        .ZN(n986) );
  INV_X1 U465 ( .A(n985), .ZN(n693) );
  AOI22_X1 U466 ( .A1(data_in[6]), .A2(n828), .B1(n991), .B2(\mem[23][6] ), 
        .ZN(n985) );
  INV_X1 U467 ( .A(n984), .ZN(n692) );
  AOI22_X1 U468 ( .A1(data_in[7]), .A2(n828), .B1(n991), .B2(\mem[23][7] ), 
        .ZN(n984) );
  INV_X1 U469 ( .A(n983), .ZN(n691) );
  AOI22_X1 U470 ( .A1(data_in[0]), .A2(n827), .B1(n982), .B2(\mem[24][0] ), 
        .ZN(n983) );
  INV_X1 U471 ( .A(n981), .ZN(n690) );
  AOI22_X1 U472 ( .A1(data_in[1]), .A2(n827), .B1(n982), .B2(\mem[24][1] ), 
        .ZN(n981) );
  INV_X1 U473 ( .A(n980), .ZN(n689) );
  AOI22_X1 U474 ( .A1(data_in[2]), .A2(n827), .B1(n982), .B2(\mem[24][2] ), 
        .ZN(n980) );
  INV_X1 U475 ( .A(n979), .ZN(n688) );
  AOI22_X1 U476 ( .A1(data_in[3]), .A2(n827), .B1(n982), .B2(\mem[24][3] ), 
        .ZN(n979) );
  INV_X1 U477 ( .A(n978), .ZN(n687) );
  AOI22_X1 U478 ( .A1(data_in[4]), .A2(n827), .B1(n982), .B2(\mem[24][4] ), 
        .ZN(n978) );
  INV_X1 U479 ( .A(n977), .ZN(n686) );
  AOI22_X1 U480 ( .A1(data_in[5]), .A2(n827), .B1(n982), .B2(\mem[24][5] ), 
        .ZN(n977) );
  INV_X1 U481 ( .A(n976), .ZN(n685) );
  AOI22_X1 U482 ( .A1(data_in[6]), .A2(n827), .B1(n982), .B2(\mem[24][6] ), 
        .ZN(n976) );
  INV_X1 U483 ( .A(n975), .ZN(n684) );
  AOI22_X1 U484 ( .A1(data_in[7]), .A2(n827), .B1(n982), .B2(\mem[24][7] ), 
        .ZN(n975) );
  INV_X1 U485 ( .A(n973), .ZN(n683) );
  AOI22_X1 U486 ( .A1(data_in[0]), .A2(n826), .B1(n972), .B2(\mem[25][0] ), 
        .ZN(n973) );
  INV_X1 U487 ( .A(n971), .ZN(n682) );
  AOI22_X1 U488 ( .A1(data_in[1]), .A2(n826), .B1(n972), .B2(\mem[25][1] ), 
        .ZN(n971) );
  INV_X1 U489 ( .A(n970), .ZN(n681) );
  AOI22_X1 U490 ( .A1(data_in[2]), .A2(n826), .B1(n972), .B2(\mem[25][2] ), 
        .ZN(n970) );
  INV_X1 U491 ( .A(n969), .ZN(n680) );
  AOI22_X1 U492 ( .A1(data_in[3]), .A2(n826), .B1(n972), .B2(\mem[25][3] ), 
        .ZN(n969) );
  INV_X1 U493 ( .A(n968), .ZN(n679) );
  AOI22_X1 U494 ( .A1(data_in[4]), .A2(n826), .B1(n972), .B2(\mem[25][4] ), 
        .ZN(n968) );
  INV_X1 U495 ( .A(n967), .ZN(n678) );
  AOI22_X1 U496 ( .A1(data_in[5]), .A2(n826), .B1(n972), .B2(\mem[25][5] ), 
        .ZN(n967) );
  INV_X1 U497 ( .A(n966), .ZN(n677) );
  AOI22_X1 U498 ( .A1(data_in[6]), .A2(n826), .B1(n972), .B2(\mem[25][6] ), 
        .ZN(n966) );
  INV_X1 U499 ( .A(n965), .ZN(n676) );
  AOI22_X1 U500 ( .A1(data_in[7]), .A2(n826), .B1(n972), .B2(\mem[25][7] ), 
        .ZN(n965) );
  INV_X1 U501 ( .A(n964), .ZN(n675) );
  AOI22_X1 U502 ( .A1(data_in[0]), .A2(n825), .B1(n963), .B2(\mem[26][0] ), 
        .ZN(n964) );
  INV_X1 U503 ( .A(n962), .ZN(n674) );
  AOI22_X1 U504 ( .A1(data_in[1]), .A2(n825), .B1(n963), .B2(\mem[26][1] ), 
        .ZN(n962) );
  INV_X1 U505 ( .A(n961), .ZN(n673) );
  AOI22_X1 U506 ( .A1(data_in[2]), .A2(n825), .B1(n963), .B2(\mem[26][2] ), 
        .ZN(n961) );
  INV_X1 U507 ( .A(n960), .ZN(n672) );
  AOI22_X1 U508 ( .A1(data_in[3]), .A2(n825), .B1(n963), .B2(\mem[26][3] ), 
        .ZN(n960) );
  INV_X1 U509 ( .A(n959), .ZN(n671) );
  AOI22_X1 U510 ( .A1(data_in[4]), .A2(n825), .B1(n963), .B2(\mem[26][4] ), 
        .ZN(n959) );
  INV_X1 U511 ( .A(n958), .ZN(n670) );
  AOI22_X1 U512 ( .A1(data_in[5]), .A2(n825), .B1(n963), .B2(\mem[26][5] ), 
        .ZN(n958) );
  INV_X1 U513 ( .A(n957), .ZN(n669) );
  AOI22_X1 U514 ( .A1(data_in[6]), .A2(n825), .B1(n963), .B2(\mem[26][6] ), 
        .ZN(n957) );
  INV_X1 U515 ( .A(n956), .ZN(n668) );
  AOI22_X1 U516 ( .A1(data_in[7]), .A2(n825), .B1(n963), .B2(\mem[26][7] ), 
        .ZN(n956) );
  INV_X1 U517 ( .A(n955), .ZN(n667) );
  AOI22_X1 U518 ( .A1(data_in[0]), .A2(n824), .B1(n954), .B2(\mem[27][0] ), 
        .ZN(n955) );
  INV_X1 U519 ( .A(n953), .ZN(n666) );
  AOI22_X1 U520 ( .A1(data_in[1]), .A2(n824), .B1(n954), .B2(\mem[27][1] ), 
        .ZN(n953) );
  INV_X1 U521 ( .A(n952), .ZN(n665) );
  AOI22_X1 U522 ( .A1(data_in[2]), .A2(n824), .B1(n954), .B2(\mem[27][2] ), 
        .ZN(n952) );
  INV_X1 U523 ( .A(n951), .ZN(n664) );
  AOI22_X1 U524 ( .A1(data_in[3]), .A2(n824), .B1(n954), .B2(\mem[27][3] ), 
        .ZN(n951) );
  INV_X1 U525 ( .A(n950), .ZN(n663) );
  AOI22_X1 U526 ( .A1(data_in[4]), .A2(n824), .B1(n954), .B2(\mem[27][4] ), 
        .ZN(n950) );
  INV_X1 U527 ( .A(n949), .ZN(n662) );
  AOI22_X1 U528 ( .A1(data_in[5]), .A2(n824), .B1(n954), .B2(\mem[27][5] ), 
        .ZN(n949) );
  INV_X1 U529 ( .A(n948), .ZN(n661) );
  AOI22_X1 U530 ( .A1(data_in[6]), .A2(n824), .B1(n954), .B2(\mem[27][6] ), 
        .ZN(n948) );
  INV_X1 U531 ( .A(n947), .ZN(n660) );
  AOI22_X1 U532 ( .A1(data_in[7]), .A2(n824), .B1(n954), .B2(\mem[27][7] ), 
        .ZN(n947) );
  INV_X1 U533 ( .A(n946), .ZN(n659) );
  AOI22_X1 U534 ( .A1(data_in[0]), .A2(n823), .B1(n945), .B2(\mem[28][0] ), 
        .ZN(n946) );
  INV_X1 U535 ( .A(n944), .ZN(n658) );
  AOI22_X1 U536 ( .A1(data_in[1]), .A2(n823), .B1(n945), .B2(\mem[28][1] ), 
        .ZN(n944) );
  INV_X1 U537 ( .A(n943), .ZN(n657) );
  AOI22_X1 U538 ( .A1(data_in[2]), .A2(n823), .B1(n945), .B2(\mem[28][2] ), 
        .ZN(n943) );
  INV_X1 U539 ( .A(n942), .ZN(n656) );
  AOI22_X1 U540 ( .A1(data_in[3]), .A2(n823), .B1(n945), .B2(\mem[28][3] ), 
        .ZN(n942) );
  INV_X1 U541 ( .A(n941), .ZN(n655) );
  AOI22_X1 U542 ( .A1(data_in[4]), .A2(n823), .B1(n945), .B2(\mem[28][4] ), 
        .ZN(n941) );
  INV_X1 U543 ( .A(n940), .ZN(n654) );
  AOI22_X1 U544 ( .A1(data_in[5]), .A2(n823), .B1(n945), .B2(\mem[28][5] ), 
        .ZN(n940) );
  INV_X1 U545 ( .A(n939), .ZN(n653) );
  AOI22_X1 U546 ( .A1(data_in[6]), .A2(n823), .B1(n945), .B2(\mem[28][6] ), 
        .ZN(n939) );
  INV_X1 U547 ( .A(n938), .ZN(n652) );
  AOI22_X1 U548 ( .A1(data_in[7]), .A2(n823), .B1(n945), .B2(\mem[28][7] ), 
        .ZN(n938) );
  INV_X1 U549 ( .A(n937), .ZN(n651) );
  AOI22_X1 U550 ( .A1(data_in[0]), .A2(n822), .B1(n936), .B2(\mem[29][0] ), 
        .ZN(n937) );
  INV_X1 U551 ( .A(n935), .ZN(n650) );
  AOI22_X1 U552 ( .A1(data_in[1]), .A2(n822), .B1(n936), .B2(\mem[29][1] ), 
        .ZN(n935) );
  INV_X1 U553 ( .A(n934), .ZN(n649) );
  AOI22_X1 U554 ( .A1(data_in[2]), .A2(n822), .B1(n936), .B2(\mem[29][2] ), 
        .ZN(n934) );
  INV_X1 U555 ( .A(n933), .ZN(n648) );
  AOI22_X1 U556 ( .A1(data_in[3]), .A2(n822), .B1(n936), .B2(\mem[29][3] ), 
        .ZN(n933) );
  INV_X1 U557 ( .A(n932), .ZN(n647) );
  AOI22_X1 U558 ( .A1(data_in[4]), .A2(n822), .B1(n936), .B2(\mem[29][4] ), 
        .ZN(n932) );
  INV_X1 U559 ( .A(n931), .ZN(n646) );
  AOI22_X1 U560 ( .A1(data_in[5]), .A2(n822), .B1(n936), .B2(\mem[29][5] ), 
        .ZN(n931) );
  INV_X1 U561 ( .A(n930), .ZN(n645) );
  AOI22_X1 U562 ( .A1(data_in[6]), .A2(n822), .B1(n936), .B2(\mem[29][6] ), 
        .ZN(n930) );
  INV_X1 U563 ( .A(n929), .ZN(n644) );
  AOI22_X1 U564 ( .A1(data_in[7]), .A2(n822), .B1(n936), .B2(\mem[29][7] ), 
        .ZN(n929) );
  INV_X1 U565 ( .A(n928), .ZN(n643) );
  AOI22_X1 U566 ( .A1(data_in[0]), .A2(n821), .B1(n927), .B2(\mem[30][0] ), 
        .ZN(n928) );
  INV_X1 U567 ( .A(n926), .ZN(n642) );
  AOI22_X1 U568 ( .A1(data_in[1]), .A2(n821), .B1(n927), .B2(\mem[30][1] ), 
        .ZN(n926) );
  INV_X1 U569 ( .A(n925), .ZN(n641) );
  AOI22_X1 U570 ( .A1(data_in[2]), .A2(n821), .B1(n927), .B2(\mem[30][2] ), 
        .ZN(n925) );
  INV_X1 U571 ( .A(n924), .ZN(n640) );
  AOI22_X1 U572 ( .A1(data_in[3]), .A2(n821), .B1(n927), .B2(\mem[30][3] ), 
        .ZN(n924) );
  INV_X1 U573 ( .A(n923), .ZN(n639) );
  AOI22_X1 U574 ( .A1(data_in[4]), .A2(n821), .B1(n927), .B2(\mem[30][4] ), 
        .ZN(n923) );
  INV_X1 U575 ( .A(n922), .ZN(n638) );
  AOI22_X1 U576 ( .A1(data_in[5]), .A2(n821), .B1(n927), .B2(\mem[30][5] ), 
        .ZN(n922) );
  INV_X1 U577 ( .A(n921), .ZN(n637) );
  AOI22_X1 U578 ( .A1(data_in[6]), .A2(n821), .B1(n927), .B2(\mem[30][6] ), 
        .ZN(n921) );
  INV_X1 U579 ( .A(n920), .ZN(n636) );
  AOI22_X1 U580 ( .A1(data_in[7]), .A2(n821), .B1(n927), .B2(\mem[30][7] ), 
        .ZN(n920) );
  INV_X1 U581 ( .A(n919), .ZN(n635) );
  AOI22_X1 U582 ( .A1(data_in[0]), .A2(n820), .B1(n918), .B2(\mem[31][0] ), 
        .ZN(n919) );
  INV_X1 U583 ( .A(n917), .ZN(n634) );
  AOI22_X1 U584 ( .A1(data_in[1]), .A2(n820), .B1(n918), .B2(\mem[31][1] ), 
        .ZN(n917) );
  INV_X1 U585 ( .A(n916), .ZN(n633) );
  AOI22_X1 U586 ( .A1(data_in[2]), .A2(n820), .B1(n918), .B2(\mem[31][2] ), 
        .ZN(n916) );
  INV_X1 U587 ( .A(n915), .ZN(n632) );
  AOI22_X1 U588 ( .A1(data_in[3]), .A2(n820), .B1(n918), .B2(\mem[31][3] ), 
        .ZN(n915) );
  INV_X1 U589 ( .A(n914), .ZN(n631) );
  AOI22_X1 U590 ( .A1(data_in[4]), .A2(n820), .B1(n918), .B2(\mem[31][4] ), 
        .ZN(n914) );
  INV_X1 U591 ( .A(n913), .ZN(n630) );
  AOI22_X1 U592 ( .A1(data_in[5]), .A2(n820), .B1(n918), .B2(\mem[31][5] ), 
        .ZN(n913) );
  INV_X1 U593 ( .A(n912), .ZN(n629) );
  AOI22_X1 U594 ( .A1(data_in[6]), .A2(n820), .B1(n918), .B2(\mem[31][6] ), 
        .ZN(n912) );
  INV_X1 U595 ( .A(n911), .ZN(n628) );
  AOI22_X1 U596 ( .A1(data_in[7]), .A2(n820), .B1(n918), .B2(\mem[31][7] ), 
        .ZN(n911) );
  MUX2_X1 U597 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n614), .Z(n2) );
  MUX2_X1 U598 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n614), .Z(n3) );
  MUX2_X1 U599 ( .A(n3), .B(n2), .S(n609), .Z(n4) );
  MUX2_X1 U600 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n614), .Z(n5) );
  MUX2_X1 U601 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n614), .Z(n6) );
  MUX2_X1 U602 ( .A(n6), .B(n5), .S(n609), .Z(n7) );
  MUX2_X1 U603 ( .A(n7), .B(n4), .S(n607), .Z(n8) );
  MUX2_X1 U604 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n614), .Z(n9) );
  MUX2_X1 U605 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n614), .Z(n10) );
  MUX2_X1 U606 ( .A(n10), .B(n9), .S(n609), .Z(n11) );
  MUX2_X1 U607 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n614), .Z(n12) );
  MUX2_X1 U608 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n614), .Z(n13) );
  MUX2_X1 U609 ( .A(n13), .B(n12), .S(n609), .Z(n14) );
  MUX2_X1 U610 ( .A(n14), .B(n11), .S(n607), .Z(n15) );
  MUX2_X1 U611 ( .A(n15), .B(n8), .S(N13), .Z(n16) );
  MUX2_X1 U612 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n612), .Z(n17) );
  MUX2_X1 U613 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n612), .Z(n18) );
  MUX2_X1 U614 ( .A(n18), .B(n17), .S(n609), .Z(n19) );
  MUX2_X1 U615 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n612), .Z(n20) );
  MUX2_X1 U616 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n612), .Z(n21) );
  MUX2_X1 U617 ( .A(n21), .B(n20), .S(n610), .Z(n22) );
  MUX2_X1 U618 ( .A(n22), .B(n19), .S(n607), .Z(n23) );
  MUX2_X1 U619 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n612), .Z(n24) );
  MUX2_X1 U620 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n612), .Z(n25) );
  MUX2_X1 U621 ( .A(n25), .B(n24), .S(n609), .Z(n26) );
  MUX2_X1 U622 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n612), .Z(n27) );
  MUX2_X1 U623 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n612), .Z(n28) );
  MUX2_X1 U624 ( .A(n28), .B(n27), .S(N11), .Z(n29) );
  MUX2_X1 U625 ( .A(n29), .B(n26), .S(n607), .Z(n30) );
  MUX2_X1 U626 ( .A(n30), .B(n23), .S(N13), .Z(n31) );
  MUX2_X1 U627 ( .A(n31), .B(n16), .S(N14), .Z(N22) );
  MUX2_X1 U628 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n612), .Z(n32) );
  MUX2_X1 U629 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n612), .Z(n33) );
  MUX2_X1 U630 ( .A(n33), .B(n32), .S(n609), .Z(n34) );
  MUX2_X1 U631 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n612), .Z(n35) );
  MUX2_X1 U632 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n612), .Z(n36) );
  MUX2_X1 U633 ( .A(n36), .B(n35), .S(n609), .Z(n37) );
  MUX2_X1 U634 ( .A(n37), .B(n34), .S(n607), .Z(n38) );
  MUX2_X1 U635 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n613), .Z(n39) );
  MUX2_X1 U636 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n615), .Z(n40) );
  MUX2_X1 U637 ( .A(n40), .B(n39), .S(n609), .Z(n41) );
  MUX2_X1 U638 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n612), .Z(n42) );
  MUX2_X1 U639 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n616), .Z(n43) );
  MUX2_X1 U640 ( .A(n43), .B(n42), .S(n609), .Z(n44) );
  MUX2_X1 U641 ( .A(n44), .B(n41), .S(n607), .Z(n45) );
  MUX2_X1 U642 ( .A(n45), .B(n38), .S(N13), .Z(n46) );
  MUX2_X1 U643 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n616), .Z(n47) );
  MUX2_X1 U644 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n616), .Z(n48) );
  MUX2_X1 U645 ( .A(n48), .B(n47), .S(n609), .Z(n49) );
  MUX2_X1 U646 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n615), .Z(n50) );
  MUX2_X1 U647 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n612), .Z(n51) );
  MUX2_X1 U648 ( .A(n51), .B(n50), .S(n611), .Z(n52) );
  MUX2_X1 U649 ( .A(n52), .B(n49), .S(n607), .Z(n53) );
  MUX2_X1 U650 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n613), .Z(n54) );
  MUX2_X1 U651 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n615), .Z(n55) );
  MUX2_X1 U652 ( .A(n55), .B(n54), .S(n609), .Z(n56) );
  MUX2_X1 U653 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n613), .Z(n57) );
  MUX2_X1 U654 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n612), .Z(n58) );
  MUX2_X1 U655 ( .A(n58), .B(n57), .S(n609), .Z(n59) );
  MUX2_X1 U656 ( .A(n59), .B(n56), .S(n607), .Z(n60) );
  MUX2_X1 U657 ( .A(n60), .B(n53), .S(N13), .Z(n61) );
  MUX2_X1 U658 ( .A(n61), .B(n46), .S(N14), .Z(N21) );
  MUX2_X1 U659 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n615), .Z(n62) );
  MUX2_X1 U660 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n613), .Z(n63) );
  MUX2_X1 U661 ( .A(n63), .B(n62), .S(n610), .Z(n64) );
  MUX2_X1 U662 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n617), .Z(n65) );
  MUX2_X1 U663 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n613), .Z(n66) );
  MUX2_X1 U664 ( .A(n66), .B(n65), .S(n610), .Z(n67) );
  MUX2_X1 U665 ( .A(n67), .B(n64), .S(n607), .Z(n68) );
  MUX2_X1 U666 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n613), .Z(n69) );
  MUX2_X1 U667 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n616), .Z(n70) );
  MUX2_X1 U668 ( .A(n70), .B(n69), .S(n610), .Z(n71) );
  MUX2_X1 U669 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n616), .Z(n72) );
  MUX2_X1 U670 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n616), .Z(n73) );
  MUX2_X1 U671 ( .A(n73), .B(n72), .S(n610), .Z(n74) );
  MUX2_X1 U672 ( .A(n74), .B(n71), .S(N12), .Z(n75) );
  MUX2_X1 U673 ( .A(n75), .B(n68), .S(N13), .Z(n76) );
  MUX2_X1 U674 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n612), .Z(n77) );
  MUX2_X1 U675 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n612), .Z(n78) );
  MUX2_X1 U676 ( .A(n78), .B(n77), .S(n610), .Z(n79) );
  MUX2_X1 U677 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n615), .Z(n80) );
  MUX2_X1 U678 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n615), .Z(n81) );
  MUX2_X1 U679 ( .A(n81), .B(n80), .S(n610), .Z(n82) );
  MUX2_X1 U680 ( .A(n82), .B(n79), .S(n607), .Z(n83) );
  MUX2_X1 U681 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n617), .Z(n84) );
  MUX2_X1 U682 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n613), .Z(n85) );
  MUX2_X1 U683 ( .A(n85), .B(n84), .S(n610), .Z(n86) );
  MUX2_X1 U684 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n617), .Z(n87) );
  MUX2_X1 U685 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n616), .Z(n88) );
  MUX2_X1 U686 ( .A(n88), .B(n87), .S(n610), .Z(n89) );
  MUX2_X1 U687 ( .A(n89), .B(n86), .S(n608), .Z(n90) );
  MUX2_X1 U688 ( .A(n90), .B(n83), .S(N13), .Z(n91) );
  MUX2_X1 U689 ( .A(n91), .B(n76), .S(N14), .Z(N20) );
  MUX2_X1 U690 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n616), .Z(n92) );
  MUX2_X1 U691 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n617), .Z(n93) );
  MUX2_X1 U692 ( .A(n93), .B(n92), .S(n610), .Z(n94) );
  MUX2_X1 U693 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n615), .Z(n95) );
  MUX2_X1 U694 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n617), .Z(n96) );
  MUX2_X1 U695 ( .A(n96), .B(n95), .S(n610), .Z(n97) );
  MUX2_X1 U696 ( .A(n97), .B(n94), .S(n607), .Z(n98) );
  MUX2_X1 U697 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n617), .Z(n99) );
  MUX2_X1 U698 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n617), .Z(n100) );
  MUX2_X1 U699 ( .A(n100), .B(n99), .S(n610), .Z(n101) );
  MUX2_X1 U700 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n617), .Z(n102) );
  MUX2_X1 U701 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n612), .Z(n103) );
  MUX2_X1 U702 ( .A(n103), .B(n102), .S(n610), .Z(n104) );
  MUX2_X1 U703 ( .A(n104), .B(n101), .S(N12), .Z(n105) );
  MUX2_X1 U704 ( .A(n105), .B(n98), .S(N13), .Z(n106) );
  MUX2_X1 U705 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n613), .Z(n107) );
  MUX2_X1 U706 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n613), .Z(n108) );
  MUX2_X1 U707 ( .A(n108), .B(n107), .S(n611), .Z(n109) );
  MUX2_X1 U708 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n613), .Z(n110) );
  MUX2_X1 U709 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n613), .Z(n111) );
  MUX2_X1 U710 ( .A(n111), .B(n110), .S(n611), .Z(n112) );
  MUX2_X1 U711 ( .A(n112), .B(n109), .S(n608), .Z(n113) );
  MUX2_X1 U712 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n613), .Z(n114) );
  MUX2_X1 U713 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n613), .Z(n115) );
  MUX2_X1 U714 ( .A(n115), .B(n114), .S(n611), .Z(n116) );
  MUX2_X1 U715 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n613), .Z(n117) );
  MUX2_X1 U716 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n613), .Z(n118) );
  MUX2_X1 U717 ( .A(n118), .B(n117), .S(n611), .Z(n119) );
  MUX2_X1 U718 ( .A(n119), .B(n116), .S(n607), .Z(n120) );
  MUX2_X1 U719 ( .A(n120), .B(n113), .S(N13), .Z(n121) );
  MUX2_X1 U720 ( .A(n121), .B(n106), .S(N14), .Z(N19) );
  MUX2_X1 U721 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n613), .Z(n122) );
  MUX2_X1 U722 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n613), .Z(n123) );
  MUX2_X1 U723 ( .A(n123), .B(n122), .S(n611), .Z(n124) );
  MUX2_X1 U724 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n613), .Z(n125) );
  MUX2_X1 U725 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n613), .Z(n126) );
  MUX2_X1 U726 ( .A(n126), .B(n125), .S(n611), .Z(n127) );
  MUX2_X1 U727 ( .A(n127), .B(n124), .S(n607), .Z(n128) );
  MUX2_X1 U728 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n614), .Z(n129) );
  MUX2_X1 U729 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n614), .Z(n130) );
  MUX2_X1 U730 ( .A(n130), .B(n129), .S(n611), .Z(n131) );
  MUX2_X1 U731 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n614), .Z(n132) );
  MUX2_X1 U732 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n614), .Z(n133) );
  MUX2_X1 U733 ( .A(n133), .B(n132), .S(n611), .Z(n134) );
  MUX2_X1 U734 ( .A(n134), .B(n131), .S(N12), .Z(n135) );
  MUX2_X1 U735 ( .A(n135), .B(n128), .S(N13), .Z(n136) );
  MUX2_X1 U736 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n614), .Z(n137) );
  MUX2_X1 U737 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n614), .Z(n138) );
  MUX2_X1 U738 ( .A(n138), .B(n137), .S(n611), .Z(n139) );
  MUX2_X1 U739 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n614), .Z(n140) );
  MUX2_X1 U740 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n614), .Z(n141) );
  MUX2_X1 U741 ( .A(n141), .B(n140), .S(n611), .Z(n142) );
  MUX2_X1 U742 ( .A(n142), .B(n139), .S(n607), .Z(n143) );
  MUX2_X1 U743 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n614), .Z(n144) );
  MUX2_X1 U744 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n614), .Z(n145) );
  MUX2_X1 U745 ( .A(n145), .B(n144), .S(n611), .Z(n146) );
  MUX2_X1 U746 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n614), .Z(n147) );
  MUX2_X1 U747 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n614), .Z(n148) );
  MUX2_X1 U748 ( .A(n148), .B(n147), .S(n611), .Z(n149) );
  MUX2_X1 U749 ( .A(n149), .B(n146), .S(n608), .Z(n150) );
  MUX2_X1 U750 ( .A(n150), .B(n143), .S(N13), .Z(n151) );
  MUX2_X1 U751 ( .A(n151), .B(n136), .S(N14), .Z(N18) );
  MUX2_X1 U752 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n615), .Z(n152) );
  MUX2_X1 U753 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n615), .Z(n153) );
  MUX2_X1 U754 ( .A(n153), .B(n152), .S(n610), .Z(n154) );
  MUX2_X1 U755 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n615), .Z(n155) );
  MUX2_X1 U756 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n615), .Z(n156) );
  MUX2_X1 U757 ( .A(n156), .B(n155), .S(n609), .Z(n157) );
  MUX2_X1 U758 ( .A(n157), .B(n154), .S(n608), .Z(n158) );
  MUX2_X1 U759 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n615), .Z(n159) );
  MUX2_X1 U760 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n615), .Z(n160) );
  MUX2_X1 U761 ( .A(n160), .B(n159), .S(n610), .Z(n161) );
  MUX2_X1 U762 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n615), .Z(n162) );
  MUX2_X1 U763 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n615), .Z(n163) );
  MUX2_X1 U764 ( .A(n163), .B(n162), .S(n609), .Z(n164) );
  MUX2_X1 U765 ( .A(n164), .B(n161), .S(n608), .Z(n165) );
  MUX2_X1 U766 ( .A(n165), .B(n158), .S(N13), .Z(n166) );
  MUX2_X1 U767 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n615), .Z(n167) );
  MUX2_X1 U768 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n615), .Z(n168) );
  MUX2_X1 U769 ( .A(n168), .B(n167), .S(N11), .Z(n169) );
  MUX2_X1 U770 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n615), .Z(n170) );
  MUX2_X1 U771 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n615), .Z(n171) );
  MUX2_X1 U772 ( .A(n171), .B(n170), .S(n611), .Z(n172) );
  MUX2_X1 U773 ( .A(n172), .B(n169), .S(n608), .Z(n173) );
  MUX2_X1 U774 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n617), .Z(n174) );
  MUX2_X1 U775 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n617), .Z(n175) );
  MUX2_X1 U776 ( .A(n175), .B(n174), .S(n610), .Z(n176) );
  MUX2_X1 U777 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n617), .Z(n177) );
  MUX2_X1 U778 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n178) );
  MUX2_X1 U779 ( .A(n178), .B(n177), .S(n610), .Z(n179) );
  MUX2_X1 U780 ( .A(n179), .B(n176), .S(n608), .Z(n180) );
  MUX2_X1 U781 ( .A(n180), .B(n173), .S(N13), .Z(n181) );
  MUX2_X1 U782 ( .A(n181), .B(n166), .S(N14), .Z(N17) );
  MUX2_X1 U783 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n617), .Z(n182) );
  MUX2_X1 U784 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n615), .Z(n183) );
  MUX2_X1 U785 ( .A(n183), .B(n182), .S(n609), .Z(n184) );
  MUX2_X1 U786 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n617), .Z(n185) );
  MUX2_X1 U787 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n617), .Z(n186) );
  MUX2_X1 U788 ( .A(n186), .B(n185), .S(n611), .Z(n187) );
  MUX2_X1 U789 ( .A(n187), .B(n184), .S(n608), .Z(n188) );
  MUX2_X1 U790 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n612), .Z(n189) );
  MUX2_X1 U791 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n612), .Z(n190) );
  MUX2_X1 U792 ( .A(n190), .B(n189), .S(n609), .Z(n191) );
  MUX2_X1 U793 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n617), .Z(n192) );
  MUX2_X1 U794 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n617), .Z(n193) );
  MUX2_X1 U795 ( .A(n193), .B(n192), .S(n610), .Z(n194) );
  MUX2_X1 U796 ( .A(n194), .B(n191), .S(n608), .Z(n195) );
  MUX2_X1 U797 ( .A(n195), .B(n188), .S(N13), .Z(n196) );
  MUX2_X1 U798 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n614), .Z(n197) );
  MUX2_X1 U799 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n617), .Z(n198) );
  MUX2_X1 U800 ( .A(n198), .B(n197), .S(n611), .Z(n199) );
  MUX2_X1 U801 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n617), .Z(n200) );
  MUX2_X1 U802 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n201) );
  MUX2_X1 U803 ( .A(n201), .B(n200), .S(n611), .Z(n202) );
  MUX2_X1 U804 ( .A(n202), .B(n199), .S(n608), .Z(n203) );
  MUX2_X1 U805 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n617), .Z(n204) );
  MUX2_X1 U806 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n205) );
  MUX2_X1 U807 ( .A(n205), .B(n204), .S(N11), .Z(n206) );
  MUX2_X1 U808 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n207) );
  MUX2_X1 U809 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n208) );
  MUX2_X1 U810 ( .A(n208), .B(n207), .S(n610), .Z(n209) );
  MUX2_X1 U811 ( .A(n209), .B(n206), .S(n608), .Z(n210) );
  MUX2_X1 U812 ( .A(n210), .B(n203), .S(N13), .Z(n211) );
  MUX2_X1 U813 ( .A(n211), .B(n196), .S(N14), .Z(N16) );
  MUX2_X1 U814 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n614), .Z(n212) );
  MUX2_X1 U815 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n614), .Z(n213) );
  MUX2_X1 U816 ( .A(n213), .B(n212), .S(n610), .Z(n214) );
  MUX2_X1 U817 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n613), .Z(n215) );
  MUX2_X1 U818 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n617), .Z(n216) );
  MUX2_X1 U819 ( .A(n216), .B(n215), .S(N11), .Z(n217) );
  MUX2_X1 U820 ( .A(n217), .B(n214), .S(n608), .Z(n218) );
  MUX2_X1 U821 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n616), .Z(n219) );
  MUX2_X1 U822 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n616), .Z(n220) );
  MUX2_X1 U823 ( .A(n220), .B(n219), .S(n609), .Z(n221) );
  MUX2_X1 U824 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n616), .Z(n222) );
  MUX2_X1 U825 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n616), .Z(n223) );
  MUX2_X1 U826 ( .A(n223), .B(n222), .S(N11), .Z(n224) );
  MUX2_X1 U827 ( .A(n224), .B(n221), .S(n608), .Z(n225) );
  MUX2_X1 U828 ( .A(n225), .B(n218), .S(N13), .Z(n226) );
  MUX2_X1 U829 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n616), .Z(n227) );
  MUX2_X1 U830 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n616), .Z(n228) );
  MUX2_X1 U831 ( .A(n228), .B(n227), .S(n611), .Z(n229) );
  MUX2_X1 U832 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n616), .Z(n595) );
  MUX2_X1 U833 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n616), .Z(n596) );
  MUX2_X1 U834 ( .A(n596), .B(n595), .S(n611), .Z(n597) );
  MUX2_X1 U835 ( .A(n597), .B(n229), .S(n608), .Z(n598) );
  MUX2_X1 U836 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n616), .Z(n599) );
  MUX2_X1 U837 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n616), .Z(n600) );
  MUX2_X1 U838 ( .A(n600), .B(n599), .S(n610), .Z(n601) );
  MUX2_X1 U839 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n616), .Z(n602) );
  MUX2_X1 U840 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n616), .Z(n603) );
  MUX2_X1 U841 ( .A(n603), .B(n602), .S(n611), .Z(n604) );
  MUX2_X1 U842 ( .A(n604), .B(n601), .S(n608), .Z(n605) );
  MUX2_X1 U843 ( .A(n605), .B(n598), .S(N13), .Z(n606) );
  MUX2_X1 U844 ( .A(n606), .B(n226), .S(N14), .Z(N15) );
  CLKBUF_X1 U845 ( .A(N11), .Z(n609) );
  INV_X1 U846 ( .A(N10), .ZN(n618) );
  INV_X1 U847 ( .A(N11), .ZN(n619) );
  INV_X1 U848 ( .A(data_in[0]), .ZN(n620) );
  INV_X1 U849 ( .A(data_in[1]), .ZN(n621) );
  INV_X1 U850 ( .A(data_in[2]), .ZN(n622) );
  INV_X1 U851 ( .A(data_in[3]), .ZN(n623) );
  INV_X1 U852 ( .A(data_in[4]), .ZN(n624) );
  INV_X1 U853 ( .A(data_in[5]), .ZN(n625) );
  INV_X1 U854 ( .A(data_in[6]), .ZN(n626) );
  INV_X1 U855 ( .A(data_in[7]), .ZN(n627) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_23 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n631), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n632), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n633), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n634), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n635), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n636), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n637), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n638), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n639), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n640), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n641), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n642), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n643), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n644), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n645), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n646), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n647), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n648), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n649), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n650), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n651), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n652), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n653), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n654), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n655), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n656), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n657), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n658), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n659), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n660), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n661), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n662), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n663), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n664), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n665), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n666), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n667), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n668), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n669), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n670), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n671), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n672), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n673), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n674), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n675), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n676), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n677), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n678), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n679), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n680), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n681), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n682), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n683), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n684), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n685), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n686), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n687), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n688), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n689), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n690), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n691), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n692), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n693), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n694), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n695), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n696), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n697), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n698), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n699), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n700), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n701), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n702), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n703), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n704), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n705), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n706), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n707), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n708), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n709), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n710), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n711), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n712), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n713), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n714), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n715), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n716), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n717), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n718), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n719), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n720), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n721), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n722), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n723), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n724), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n725), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n726), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n727), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n728), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n729), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n730), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n731), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n732), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n733), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n734), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n735), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n736), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n737), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n738), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n739), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n740), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n741), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n742), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n743), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n744), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n745), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n746), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n747), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n748), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n749), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n750), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n751), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n752), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n753), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n754), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n755), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n756), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n757), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n758), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n759), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n760), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n761), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n762), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n763), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n764), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n765), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n766), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n767), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n768), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n769), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n770), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n771), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n772), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n773), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n774), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n775), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n776), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n777), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n778), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n779), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n780), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n781), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n782), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n783), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n784), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n785), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n786), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n787), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n788), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n789), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n790), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n791), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n792), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n793), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n794), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n795), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n796), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n797), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n798), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n799), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n800), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n801), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n802), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n803), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n804), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n805), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n806), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n807), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n808), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n809), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n810), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n811), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n812), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n813), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n814), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n815), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n816), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n817), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n818), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n819), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n820), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n821), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n822), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n850), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n851), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n852), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n853), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n854), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n855), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n856), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n857), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n858), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n859), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n860), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n861), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n862), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n863), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n864), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n865), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n866), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n867), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n868), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n869), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n870), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n871), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n872), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n873), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n874), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n875), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n876), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n877), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n878), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n879), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n880), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n881), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n882), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n883), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n884), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n885), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n886), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n887), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n888), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n889), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n890), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n891), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n892), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n893), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n894), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n895), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n896), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n897), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n898), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n899), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n900), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n901), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n902), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n903), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n904), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n905), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n906), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n907), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n908), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n909), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n910), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n911), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n912), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n913), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n3) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n619), .Z(n615) );
  INV_X2 U4 ( .A(n3), .ZN(data_out[3]) );
  BUF_X1 U5 ( .A(n619), .Z(n617) );
  BUF_X1 U6 ( .A(n619), .Z(n616) );
  BUF_X1 U7 ( .A(n619), .Z(n618) );
  BUF_X1 U8 ( .A(N11), .Z(n613) );
  BUF_X1 U9 ( .A(N11), .Z(n614) );
  BUF_X1 U10 ( .A(N10), .Z(n620) );
  BUF_X1 U11 ( .A(N10), .Z(n619) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1205) );
  NOR3_X1 U13 ( .A1(N11), .A2(N12), .A3(n621), .ZN(n1194) );
  NOR3_X1 U14 ( .A1(N10), .A2(N12), .A3(n622), .ZN(n1184) );
  NOR3_X1 U15 ( .A1(n621), .A2(N12), .A3(n622), .ZN(n1174) );
  INV_X1 U16 ( .A(n1131), .ZN(n846) );
  INV_X1 U17 ( .A(n1121), .ZN(n845) );
  INV_X1 U18 ( .A(n1112), .ZN(n844) );
  INV_X1 U19 ( .A(n1103), .ZN(n843) );
  INV_X1 U20 ( .A(n1058), .ZN(n838) );
  INV_X1 U21 ( .A(n1048), .ZN(n837) );
  INV_X1 U22 ( .A(n1039), .ZN(n836) );
  INV_X1 U23 ( .A(n1030), .ZN(n835) );
  INV_X1 U24 ( .A(n985), .ZN(n830) );
  INV_X1 U25 ( .A(n975), .ZN(n829) );
  INV_X1 U26 ( .A(n966), .ZN(n828) );
  INV_X1 U27 ( .A(n957), .ZN(n827) );
  INV_X1 U28 ( .A(n921), .ZN(n823) );
  INV_X1 U29 ( .A(n1094), .ZN(n842) );
  INV_X1 U30 ( .A(n1085), .ZN(n841) );
  INV_X1 U31 ( .A(n1076), .ZN(n840) );
  INV_X1 U32 ( .A(n1067), .ZN(n839) );
  INV_X1 U33 ( .A(n948), .ZN(n826) );
  INV_X1 U34 ( .A(n939), .ZN(n825) );
  INV_X1 U35 ( .A(n930), .ZN(n824) );
  INV_X1 U36 ( .A(n1021), .ZN(n834) );
  INV_X1 U37 ( .A(n1012), .ZN(n833) );
  INV_X1 U38 ( .A(n1003), .ZN(n832) );
  INV_X1 U39 ( .A(n994), .ZN(n831) );
  BUF_X1 U40 ( .A(N12), .Z(n611) );
  INV_X1 U41 ( .A(N13), .ZN(n848) );
  AND3_X1 U42 ( .A1(n621), .A2(n622), .A3(N12), .ZN(n1164) );
  AND3_X1 U43 ( .A1(N10), .A2(n622), .A3(N12), .ZN(n1154) );
  AND3_X1 U44 ( .A1(N11), .A2(n621), .A3(N12), .ZN(n1144) );
  AND3_X1 U45 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1134) );
  BUF_X1 U46 ( .A(N12), .Z(n610) );
  INV_X1 U47 ( .A(N14), .ZN(n849) );
  NAND2_X1 U48 ( .A1(n1194), .A2(n1204), .ZN(n1203) );
  NAND2_X1 U49 ( .A1(n1184), .A2(n1204), .ZN(n1193) );
  NAND2_X1 U50 ( .A1(n1174), .A2(n1204), .ZN(n1183) );
  NAND2_X1 U51 ( .A1(n1164), .A2(n1204), .ZN(n1173) );
  NAND2_X1 U52 ( .A1(n1154), .A2(n1204), .ZN(n1163) );
  NAND2_X1 U53 ( .A1(n1144), .A2(n1204), .ZN(n1153) );
  NAND2_X1 U54 ( .A1(n1134), .A2(n1204), .ZN(n1143) );
  NAND2_X1 U55 ( .A1(n1205), .A2(n1204), .ZN(n1214) );
  NAND2_X1 U56 ( .A1(n1123), .A2(n1205), .ZN(n1131) );
  NAND2_X1 U57 ( .A1(n1123), .A2(n1194), .ZN(n1121) );
  NAND2_X1 U58 ( .A1(n1123), .A2(n1184), .ZN(n1112) );
  NAND2_X1 U59 ( .A1(n1123), .A2(n1174), .ZN(n1103) );
  NAND2_X1 U60 ( .A1(n1050), .A2(n1205), .ZN(n1058) );
  NAND2_X1 U61 ( .A1(n1050), .A2(n1194), .ZN(n1048) );
  NAND2_X1 U62 ( .A1(n1050), .A2(n1184), .ZN(n1039) );
  NAND2_X1 U63 ( .A1(n1050), .A2(n1174), .ZN(n1030) );
  NAND2_X1 U64 ( .A1(n977), .A2(n1205), .ZN(n985) );
  NAND2_X1 U65 ( .A1(n977), .A2(n1194), .ZN(n975) );
  NAND2_X1 U66 ( .A1(n977), .A2(n1184), .ZN(n966) );
  NAND2_X1 U67 ( .A1(n977), .A2(n1174), .ZN(n957) );
  NAND2_X1 U68 ( .A1(n1123), .A2(n1164), .ZN(n1094) );
  NAND2_X1 U69 ( .A1(n1123), .A2(n1154), .ZN(n1085) );
  NAND2_X1 U70 ( .A1(n1123), .A2(n1144), .ZN(n1076) );
  NAND2_X1 U71 ( .A1(n1123), .A2(n1134), .ZN(n1067) );
  NAND2_X1 U72 ( .A1(n1050), .A2(n1164), .ZN(n1021) );
  NAND2_X1 U73 ( .A1(n1050), .A2(n1154), .ZN(n1012) );
  NAND2_X1 U74 ( .A1(n1050), .A2(n1144), .ZN(n1003) );
  NAND2_X1 U75 ( .A1(n1050), .A2(n1134), .ZN(n994) );
  NAND2_X1 U76 ( .A1(n977), .A2(n1164), .ZN(n948) );
  NAND2_X1 U77 ( .A1(n977), .A2(n1154), .ZN(n939) );
  NAND2_X1 U78 ( .A1(n977), .A2(n1144), .ZN(n930) );
  NAND2_X1 U79 ( .A1(n977), .A2(n1134), .ZN(n921) );
  AND3_X1 U80 ( .A1(n848), .A2(n849), .A3(n1133), .ZN(n1204) );
  AND3_X1 U81 ( .A1(N13), .A2(n1133), .A3(N14), .ZN(n977) );
  AND3_X1 U82 ( .A1(n1133), .A2(n849), .A3(N13), .ZN(n1123) );
  AND3_X1 U83 ( .A1(n1133), .A2(n848), .A3(N14), .ZN(n1050) );
  NOR2_X1 U84 ( .A1(n847), .A2(addr[5]), .ZN(n1133) );
  INV_X1 U85 ( .A(wr_en), .ZN(n847) );
  OAI21_X1 U86 ( .B1(n623), .B2(n1173), .A(n1172), .ZN(n881) );
  NAND2_X1 U87 ( .A1(\mem[4][0] ), .A2(n1173), .ZN(n1172) );
  OAI21_X1 U88 ( .B1(n624), .B2(n1173), .A(n1171), .ZN(n880) );
  NAND2_X1 U89 ( .A1(\mem[4][1] ), .A2(n1173), .ZN(n1171) );
  OAI21_X1 U90 ( .B1(n625), .B2(n1173), .A(n1170), .ZN(n879) );
  NAND2_X1 U91 ( .A1(\mem[4][2] ), .A2(n1173), .ZN(n1170) );
  OAI21_X1 U92 ( .B1(n626), .B2(n1173), .A(n1169), .ZN(n878) );
  NAND2_X1 U93 ( .A1(\mem[4][3] ), .A2(n1173), .ZN(n1169) );
  OAI21_X1 U94 ( .B1(n627), .B2(n1173), .A(n1168), .ZN(n877) );
  NAND2_X1 U95 ( .A1(\mem[4][4] ), .A2(n1173), .ZN(n1168) );
  OAI21_X1 U96 ( .B1(n628), .B2(n1173), .A(n1167), .ZN(n876) );
  NAND2_X1 U97 ( .A1(\mem[4][5] ), .A2(n1173), .ZN(n1167) );
  OAI21_X1 U98 ( .B1(n629), .B2(n1173), .A(n1166), .ZN(n875) );
  NAND2_X1 U99 ( .A1(\mem[4][6] ), .A2(n1173), .ZN(n1166) );
  OAI21_X1 U100 ( .B1(n630), .B2(n1173), .A(n1165), .ZN(n874) );
  NAND2_X1 U101 ( .A1(\mem[4][7] ), .A2(n1173), .ZN(n1165) );
  OAI21_X1 U102 ( .B1(n623), .B2(n1153), .A(n1152), .ZN(n865) );
  NAND2_X1 U103 ( .A1(\mem[6][0] ), .A2(n1153), .ZN(n1152) );
  OAI21_X1 U104 ( .B1(n624), .B2(n1153), .A(n1151), .ZN(n864) );
  NAND2_X1 U105 ( .A1(\mem[6][1] ), .A2(n1153), .ZN(n1151) );
  OAI21_X1 U106 ( .B1(n625), .B2(n1153), .A(n1150), .ZN(n863) );
  NAND2_X1 U107 ( .A1(\mem[6][2] ), .A2(n1153), .ZN(n1150) );
  OAI21_X1 U108 ( .B1(n626), .B2(n1153), .A(n1149), .ZN(n862) );
  NAND2_X1 U109 ( .A1(\mem[6][3] ), .A2(n1153), .ZN(n1149) );
  OAI21_X1 U110 ( .B1(n627), .B2(n1153), .A(n1148), .ZN(n861) );
  NAND2_X1 U111 ( .A1(\mem[6][4] ), .A2(n1153), .ZN(n1148) );
  OAI21_X1 U112 ( .B1(n628), .B2(n1153), .A(n1147), .ZN(n860) );
  NAND2_X1 U113 ( .A1(\mem[6][5] ), .A2(n1153), .ZN(n1147) );
  OAI21_X1 U114 ( .B1(n629), .B2(n1153), .A(n1146), .ZN(n859) );
  NAND2_X1 U115 ( .A1(\mem[6][6] ), .A2(n1153), .ZN(n1146) );
  OAI21_X1 U116 ( .B1(n630), .B2(n1153), .A(n1145), .ZN(n858) );
  NAND2_X1 U117 ( .A1(\mem[6][7] ), .A2(n1153), .ZN(n1145) );
  OAI21_X1 U118 ( .B1(n623), .B2(n1143), .A(n1142), .ZN(n857) );
  NAND2_X1 U119 ( .A1(\mem[7][0] ), .A2(n1143), .ZN(n1142) );
  OAI21_X1 U120 ( .B1(n624), .B2(n1143), .A(n1141), .ZN(n856) );
  NAND2_X1 U121 ( .A1(\mem[7][1] ), .A2(n1143), .ZN(n1141) );
  OAI21_X1 U122 ( .B1(n625), .B2(n1143), .A(n1140), .ZN(n855) );
  NAND2_X1 U123 ( .A1(\mem[7][2] ), .A2(n1143), .ZN(n1140) );
  OAI21_X1 U124 ( .B1(n626), .B2(n1143), .A(n1139), .ZN(n854) );
  NAND2_X1 U125 ( .A1(\mem[7][3] ), .A2(n1143), .ZN(n1139) );
  OAI21_X1 U126 ( .B1(n627), .B2(n1143), .A(n1138), .ZN(n853) );
  NAND2_X1 U127 ( .A1(\mem[7][4] ), .A2(n1143), .ZN(n1138) );
  OAI21_X1 U128 ( .B1(n628), .B2(n1143), .A(n1137), .ZN(n852) );
  NAND2_X1 U129 ( .A1(\mem[7][5] ), .A2(n1143), .ZN(n1137) );
  OAI21_X1 U130 ( .B1(n629), .B2(n1143), .A(n1136), .ZN(n851) );
  NAND2_X1 U131 ( .A1(\mem[7][6] ), .A2(n1143), .ZN(n1136) );
  OAI21_X1 U132 ( .B1(n630), .B2(n1143), .A(n1135), .ZN(n850) );
  NAND2_X1 U133 ( .A1(\mem[7][7] ), .A2(n1143), .ZN(n1135) );
  OAI21_X1 U134 ( .B1(n623), .B2(n1203), .A(n1202), .ZN(n905) );
  NAND2_X1 U135 ( .A1(\mem[1][0] ), .A2(n1203), .ZN(n1202) );
  OAI21_X1 U136 ( .B1(n624), .B2(n1203), .A(n1201), .ZN(n904) );
  NAND2_X1 U137 ( .A1(\mem[1][1] ), .A2(n1203), .ZN(n1201) );
  OAI21_X1 U138 ( .B1(n625), .B2(n1203), .A(n1200), .ZN(n903) );
  NAND2_X1 U139 ( .A1(\mem[1][2] ), .A2(n1203), .ZN(n1200) );
  OAI21_X1 U140 ( .B1(n626), .B2(n1203), .A(n1199), .ZN(n902) );
  NAND2_X1 U141 ( .A1(\mem[1][3] ), .A2(n1203), .ZN(n1199) );
  OAI21_X1 U142 ( .B1(n627), .B2(n1203), .A(n1198), .ZN(n901) );
  NAND2_X1 U143 ( .A1(\mem[1][4] ), .A2(n1203), .ZN(n1198) );
  OAI21_X1 U144 ( .B1(n628), .B2(n1203), .A(n1197), .ZN(n900) );
  NAND2_X1 U145 ( .A1(\mem[1][5] ), .A2(n1203), .ZN(n1197) );
  OAI21_X1 U146 ( .B1(n629), .B2(n1203), .A(n1196), .ZN(n899) );
  NAND2_X1 U147 ( .A1(\mem[1][6] ), .A2(n1203), .ZN(n1196) );
  OAI21_X1 U148 ( .B1(n630), .B2(n1203), .A(n1195), .ZN(n898) );
  NAND2_X1 U149 ( .A1(\mem[1][7] ), .A2(n1203), .ZN(n1195) );
  OAI21_X1 U150 ( .B1(n623), .B2(n1193), .A(n1192), .ZN(n897) );
  NAND2_X1 U151 ( .A1(\mem[2][0] ), .A2(n1193), .ZN(n1192) );
  OAI21_X1 U152 ( .B1(n624), .B2(n1193), .A(n1191), .ZN(n896) );
  NAND2_X1 U153 ( .A1(\mem[2][1] ), .A2(n1193), .ZN(n1191) );
  OAI21_X1 U154 ( .B1(n625), .B2(n1193), .A(n1190), .ZN(n895) );
  NAND2_X1 U155 ( .A1(\mem[2][2] ), .A2(n1193), .ZN(n1190) );
  OAI21_X1 U156 ( .B1(n626), .B2(n1193), .A(n1189), .ZN(n894) );
  NAND2_X1 U157 ( .A1(\mem[2][3] ), .A2(n1193), .ZN(n1189) );
  OAI21_X1 U158 ( .B1(n627), .B2(n1193), .A(n1188), .ZN(n893) );
  NAND2_X1 U159 ( .A1(\mem[2][4] ), .A2(n1193), .ZN(n1188) );
  OAI21_X1 U160 ( .B1(n628), .B2(n1193), .A(n1187), .ZN(n892) );
  NAND2_X1 U161 ( .A1(\mem[2][5] ), .A2(n1193), .ZN(n1187) );
  OAI21_X1 U162 ( .B1(n629), .B2(n1193), .A(n1186), .ZN(n891) );
  NAND2_X1 U163 ( .A1(\mem[2][6] ), .A2(n1193), .ZN(n1186) );
  OAI21_X1 U164 ( .B1(n630), .B2(n1193), .A(n1185), .ZN(n890) );
  NAND2_X1 U165 ( .A1(\mem[2][7] ), .A2(n1193), .ZN(n1185) );
  OAI21_X1 U166 ( .B1(n623), .B2(n1183), .A(n1182), .ZN(n889) );
  NAND2_X1 U167 ( .A1(\mem[3][0] ), .A2(n1183), .ZN(n1182) );
  OAI21_X1 U168 ( .B1(n624), .B2(n1183), .A(n1181), .ZN(n888) );
  NAND2_X1 U169 ( .A1(\mem[3][1] ), .A2(n1183), .ZN(n1181) );
  OAI21_X1 U170 ( .B1(n625), .B2(n1183), .A(n1180), .ZN(n887) );
  NAND2_X1 U171 ( .A1(\mem[3][2] ), .A2(n1183), .ZN(n1180) );
  OAI21_X1 U172 ( .B1(n626), .B2(n1183), .A(n1179), .ZN(n886) );
  NAND2_X1 U173 ( .A1(\mem[3][3] ), .A2(n1183), .ZN(n1179) );
  OAI21_X1 U174 ( .B1(n627), .B2(n1183), .A(n1178), .ZN(n885) );
  NAND2_X1 U175 ( .A1(\mem[3][4] ), .A2(n1183), .ZN(n1178) );
  OAI21_X1 U176 ( .B1(n628), .B2(n1183), .A(n1177), .ZN(n884) );
  NAND2_X1 U177 ( .A1(\mem[3][5] ), .A2(n1183), .ZN(n1177) );
  OAI21_X1 U178 ( .B1(n629), .B2(n1183), .A(n1176), .ZN(n883) );
  NAND2_X1 U179 ( .A1(\mem[3][6] ), .A2(n1183), .ZN(n1176) );
  OAI21_X1 U180 ( .B1(n630), .B2(n1183), .A(n1175), .ZN(n882) );
  NAND2_X1 U181 ( .A1(\mem[3][7] ), .A2(n1183), .ZN(n1175) );
  OAI21_X1 U182 ( .B1(n623), .B2(n1163), .A(n1162), .ZN(n873) );
  NAND2_X1 U183 ( .A1(\mem[5][0] ), .A2(n1163), .ZN(n1162) );
  OAI21_X1 U184 ( .B1(n624), .B2(n1163), .A(n1161), .ZN(n872) );
  NAND2_X1 U185 ( .A1(\mem[5][1] ), .A2(n1163), .ZN(n1161) );
  OAI21_X1 U186 ( .B1(n625), .B2(n1163), .A(n1160), .ZN(n871) );
  NAND2_X1 U187 ( .A1(\mem[5][2] ), .A2(n1163), .ZN(n1160) );
  OAI21_X1 U188 ( .B1(n626), .B2(n1163), .A(n1159), .ZN(n870) );
  NAND2_X1 U189 ( .A1(\mem[5][3] ), .A2(n1163), .ZN(n1159) );
  OAI21_X1 U190 ( .B1(n627), .B2(n1163), .A(n1158), .ZN(n869) );
  NAND2_X1 U191 ( .A1(\mem[5][4] ), .A2(n1163), .ZN(n1158) );
  OAI21_X1 U192 ( .B1(n628), .B2(n1163), .A(n1157), .ZN(n868) );
  NAND2_X1 U193 ( .A1(\mem[5][5] ), .A2(n1163), .ZN(n1157) );
  OAI21_X1 U194 ( .B1(n629), .B2(n1163), .A(n1156), .ZN(n867) );
  NAND2_X1 U195 ( .A1(\mem[5][6] ), .A2(n1163), .ZN(n1156) );
  OAI21_X1 U196 ( .B1(n630), .B2(n1163), .A(n1155), .ZN(n866) );
  NAND2_X1 U197 ( .A1(\mem[5][7] ), .A2(n1163), .ZN(n1155) );
  OAI21_X1 U198 ( .B1(n1214), .B2(n623), .A(n1213), .ZN(n913) );
  NAND2_X1 U199 ( .A1(\mem[0][0] ), .A2(n1214), .ZN(n1213) );
  OAI21_X1 U200 ( .B1(n1214), .B2(n624), .A(n1212), .ZN(n912) );
  NAND2_X1 U201 ( .A1(\mem[0][1] ), .A2(n1214), .ZN(n1212) );
  OAI21_X1 U202 ( .B1(n1214), .B2(n625), .A(n1211), .ZN(n911) );
  NAND2_X1 U203 ( .A1(\mem[0][2] ), .A2(n1214), .ZN(n1211) );
  OAI21_X1 U204 ( .B1(n1214), .B2(n626), .A(n1210), .ZN(n910) );
  NAND2_X1 U205 ( .A1(\mem[0][3] ), .A2(n1214), .ZN(n1210) );
  OAI21_X1 U206 ( .B1(n1214), .B2(n627), .A(n1209), .ZN(n909) );
  NAND2_X1 U207 ( .A1(\mem[0][4] ), .A2(n1214), .ZN(n1209) );
  OAI21_X1 U208 ( .B1(n1214), .B2(n628), .A(n1208), .ZN(n908) );
  NAND2_X1 U209 ( .A1(\mem[0][5] ), .A2(n1214), .ZN(n1208) );
  OAI21_X1 U210 ( .B1(n1214), .B2(n629), .A(n1207), .ZN(n907) );
  NAND2_X1 U211 ( .A1(\mem[0][6] ), .A2(n1214), .ZN(n1207) );
  OAI21_X1 U212 ( .B1(n1214), .B2(n630), .A(n1206), .ZN(n906) );
  NAND2_X1 U213 ( .A1(\mem[0][7] ), .A2(n1214), .ZN(n1206) );
  INV_X1 U214 ( .A(n1132), .ZN(n822) );
  AOI22_X1 U215 ( .A1(data_in[0]), .A2(n846), .B1(n1131), .B2(\mem[8][0] ), 
        .ZN(n1132) );
  INV_X1 U216 ( .A(n1130), .ZN(n821) );
  AOI22_X1 U217 ( .A1(data_in[1]), .A2(n846), .B1(n1131), .B2(\mem[8][1] ), 
        .ZN(n1130) );
  INV_X1 U218 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U219 ( .A1(data_in[2]), .A2(n846), .B1(n1131), .B2(\mem[8][2] ), 
        .ZN(n1129) );
  INV_X1 U220 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U221 ( .A1(data_in[3]), .A2(n846), .B1(n1131), .B2(\mem[8][3] ), 
        .ZN(n1128) );
  INV_X1 U222 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U223 ( .A1(data_in[4]), .A2(n846), .B1(n1131), .B2(\mem[8][4] ), 
        .ZN(n1127) );
  INV_X1 U224 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U225 ( .A1(data_in[5]), .A2(n846), .B1(n1131), .B2(\mem[8][5] ), 
        .ZN(n1126) );
  INV_X1 U226 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U227 ( .A1(data_in[6]), .A2(n846), .B1(n1131), .B2(\mem[8][6] ), 
        .ZN(n1125) );
  INV_X1 U228 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U229 ( .A1(data_in[7]), .A2(n846), .B1(n1131), .B2(\mem[8][7] ), 
        .ZN(n1124) );
  INV_X1 U230 ( .A(n1122), .ZN(n814) );
  AOI22_X1 U231 ( .A1(data_in[0]), .A2(n845), .B1(n1121), .B2(\mem[9][0] ), 
        .ZN(n1122) );
  INV_X1 U232 ( .A(n1120), .ZN(n813) );
  AOI22_X1 U233 ( .A1(data_in[1]), .A2(n845), .B1(n1121), .B2(\mem[9][1] ), 
        .ZN(n1120) );
  INV_X1 U234 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U235 ( .A1(data_in[2]), .A2(n845), .B1(n1121), .B2(\mem[9][2] ), 
        .ZN(n1119) );
  INV_X1 U236 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U237 ( .A1(data_in[3]), .A2(n845), .B1(n1121), .B2(\mem[9][3] ), 
        .ZN(n1118) );
  INV_X1 U238 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U239 ( .A1(data_in[4]), .A2(n845), .B1(n1121), .B2(\mem[9][4] ), 
        .ZN(n1117) );
  INV_X1 U240 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U241 ( .A1(data_in[5]), .A2(n845), .B1(n1121), .B2(\mem[9][5] ), 
        .ZN(n1116) );
  INV_X1 U242 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U243 ( .A1(data_in[6]), .A2(n845), .B1(n1121), .B2(\mem[9][6] ), 
        .ZN(n1115) );
  INV_X1 U244 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U245 ( .A1(data_in[7]), .A2(n845), .B1(n1121), .B2(\mem[9][7] ), 
        .ZN(n1114) );
  INV_X1 U246 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U247 ( .A1(data_in[0]), .A2(n844), .B1(n1112), .B2(\mem[10][0] ), 
        .ZN(n1113) );
  INV_X1 U248 ( .A(n1111), .ZN(n805) );
  AOI22_X1 U249 ( .A1(data_in[1]), .A2(n844), .B1(n1112), .B2(\mem[10][1] ), 
        .ZN(n1111) );
  INV_X1 U250 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U251 ( .A1(data_in[2]), .A2(n844), .B1(n1112), .B2(\mem[10][2] ), 
        .ZN(n1110) );
  INV_X1 U252 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U253 ( .A1(data_in[3]), .A2(n844), .B1(n1112), .B2(\mem[10][3] ), 
        .ZN(n1109) );
  INV_X1 U254 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U255 ( .A1(data_in[4]), .A2(n844), .B1(n1112), .B2(\mem[10][4] ), 
        .ZN(n1108) );
  INV_X1 U256 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U257 ( .A1(data_in[5]), .A2(n844), .B1(n1112), .B2(\mem[10][5] ), 
        .ZN(n1107) );
  INV_X1 U258 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U259 ( .A1(data_in[6]), .A2(n844), .B1(n1112), .B2(\mem[10][6] ), 
        .ZN(n1106) );
  INV_X1 U260 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U261 ( .A1(data_in[7]), .A2(n844), .B1(n1112), .B2(\mem[10][7] ), 
        .ZN(n1105) );
  INV_X1 U262 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U263 ( .A1(data_in[0]), .A2(n843), .B1(n1103), .B2(\mem[11][0] ), 
        .ZN(n1104) );
  INV_X1 U264 ( .A(n1102), .ZN(n797) );
  AOI22_X1 U265 ( .A1(data_in[1]), .A2(n843), .B1(n1103), .B2(\mem[11][1] ), 
        .ZN(n1102) );
  INV_X1 U266 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U267 ( .A1(data_in[2]), .A2(n843), .B1(n1103), .B2(\mem[11][2] ), 
        .ZN(n1101) );
  INV_X1 U268 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U269 ( .A1(data_in[3]), .A2(n843), .B1(n1103), .B2(\mem[11][3] ), 
        .ZN(n1100) );
  INV_X1 U270 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U271 ( .A1(data_in[4]), .A2(n843), .B1(n1103), .B2(\mem[11][4] ), 
        .ZN(n1099) );
  INV_X1 U272 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U273 ( .A1(data_in[5]), .A2(n843), .B1(n1103), .B2(\mem[11][5] ), 
        .ZN(n1098) );
  INV_X1 U274 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U275 ( .A1(data_in[6]), .A2(n843), .B1(n1103), .B2(\mem[11][6] ), 
        .ZN(n1097) );
  INV_X1 U276 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U277 ( .A1(data_in[7]), .A2(n843), .B1(n1103), .B2(\mem[11][7] ), 
        .ZN(n1096) );
  INV_X1 U278 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U279 ( .A1(data_in[0]), .A2(n842), .B1(n1094), .B2(\mem[12][0] ), 
        .ZN(n1095) );
  INV_X1 U280 ( .A(n1093), .ZN(n789) );
  AOI22_X1 U281 ( .A1(data_in[1]), .A2(n842), .B1(n1094), .B2(\mem[12][1] ), 
        .ZN(n1093) );
  INV_X1 U282 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U283 ( .A1(data_in[2]), .A2(n842), .B1(n1094), .B2(\mem[12][2] ), 
        .ZN(n1092) );
  INV_X1 U284 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U285 ( .A1(data_in[3]), .A2(n842), .B1(n1094), .B2(\mem[12][3] ), 
        .ZN(n1091) );
  INV_X1 U286 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U287 ( .A1(data_in[4]), .A2(n842), .B1(n1094), .B2(\mem[12][4] ), 
        .ZN(n1090) );
  INV_X1 U288 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U289 ( .A1(data_in[5]), .A2(n842), .B1(n1094), .B2(\mem[12][5] ), 
        .ZN(n1089) );
  INV_X1 U290 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U291 ( .A1(data_in[6]), .A2(n842), .B1(n1094), .B2(\mem[12][6] ), 
        .ZN(n1088) );
  INV_X1 U292 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U293 ( .A1(data_in[7]), .A2(n842), .B1(n1094), .B2(\mem[12][7] ), 
        .ZN(n1087) );
  INV_X1 U294 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U295 ( .A1(data_in[0]), .A2(n841), .B1(n1085), .B2(\mem[13][0] ), 
        .ZN(n1086) );
  INV_X1 U296 ( .A(n1084), .ZN(n781) );
  AOI22_X1 U297 ( .A1(data_in[1]), .A2(n841), .B1(n1085), .B2(\mem[13][1] ), 
        .ZN(n1084) );
  INV_X1 U298 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U299 ( .A1(data_in[2]), .A2(n841), .B1(n1085), .B2(\mem[13][2] ), 
        .ZN(n1083) );
  INV_X1 U300 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U301 ( .A1(data_in[3]), .A2(n841), .B1(n1085), .B2(\mem[13][3] ), 
        .ZN(n1082) );
  INV_X1 U302 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U303 ( .A1(data_in[4]), .A2(n841), .B1(n1085), .B2(\mem[13][4] ), 
        .ZN(n1081) );
  INV_X1 U304 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U305 ( .A1(data_in[5]), .A2(n841), .B1(n1085), .B2(\mem[13][5] ), 
        .ZN(n1080) );
  INV_X1 U306 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U307 ( .A1(data_in[6]), .A2(n841), .B1(n1085), .B2(\mem[13][6] ), 
        .ZN(n1079) );
  INV_X1 U308 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U309 ( .A1(data_in[7]), .A2(n841), .B1(n1085), .B2(\mem[13][7] ), 
        .ZN(n1078) );
  INV_X1 U310 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U311 ( .A1(data_in[0]), .A2(n840), .B1(n1076), .B2(\mem[14][0] ), 
        .ZN(n1077) );
  INV_X1 U312 ( .A(n1075), .ZN(n773) );
  AOI22_X1 U313 ( .A1(data_in[1]), .A2(n840), .B1(n1076), .B2(\mem[14][1] ), 
        .ZN(n1075) );
  INV_X1 U314 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U315 ( .A1(data_in[2]), .A2(n840), .B1(n1076), .B2(\mem[14][2] ), 
        .ZN(n1074) );
  INV_X1 U316 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U317 ( .A1(data_in[3]), .A2(n840), .B1(n1076), .B2(\mem[14][3] ), 
        .ZN(n1073) );
  INV_X1 U318 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U319 ( .A1(data_in[4]), .A2(n840), .B1(n1076), .B2(\mem[14][4] ), 
        .ZN(n1072) );
  INV_X1 U320 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U321 ( .A1(data_in[5]), .A2(n840), .B1(n1076), .B2(\mem[14][5] ), 
        .ZN(n1071) );
  INV_X1 U322 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U323 ( .A1(data_in[6]), .A2(n840), .B1(n1076), .B2(\mem[14][6] ), 
        .ZN(n1070) );
  INV_X1 U324 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U325 ( .A1(data_in[7]), .A2(n840), .B1(n1076), .B2(\mem[14][7] ), 
        .ZN(n1069) );
  INV_X1 U326 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U327 ( .A1(data_in[0]), .A2(n839), .B1(n1067), .B2(\mem[15][0] ), 
        .ZN(n1068) );
  INV_X1 U328 ( .A(n1066), .ZN(n765) );
  AOI22_X1 U329 ( .A1(data_in[1]), .A2(n839), .B1(n1067), .B2(\mem[15][1] ), 
        .ZN(n1066) );
  INV_X1 U330 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U331 ( .A1(data_in[2]), .A2(n839), .B1(n1067), .B2(\mem[15][2] ), 
        .ZN(n1065) );
  INV_X1 U332 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U333 ( .A1(data_in[3]), .A2(n839), .B1(n1067), .B2(\mem[15][3] ), 
        .ZN(n1064) );
  INV_X1 U334 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U335 ( .A1(data_in[4]), .A2(n839), .B1(n1067), .B2(\mem[15][4] ), 
        .ZN(n1063) );
  INV_X1 U336 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U337 ( .A1(data_in[5]), .A2(n839), .B1(n1067), .B2(\mem[15][5] ), 
        .ZN(n1062) );
  INV_X1 U338 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U339 ( .A1(data_in[6]), .A2(n839), .B1(n1067), .B2(\mem[15][6] ), 
        .ZN(n1061) );
  INV_X1 U340 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U341 ( .A1(data_in[7]), .A2(n839), .B1(n1067), .B2(\mem[15][7] ), 
        .ZN(n1060) );
  INV_X1 U342 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U343 ( .A1(data_in[0]), .A2(n838), .B1(n1058), .B2(\mem[16][0] ), 
        .ZN(n1059) );
  INV_X1 U344 ( .A(n1057), .ZN(n757) );
  AOI22_X1 U345 ( .A1(data_in[1]), .A2(n838), .B1(n1058), .B2(\mem[16][1] ), 
        .ZN(n1057) );
  INV_X1 U346 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U347 ( .A1(data_in[2]), .A2(n838), .B1(n1058), .B2(\mem[16][2] ), 
        .ZN(n1056) );
  INV_X1 U348 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U349 ( .A1(data_in[3]), .A2(n838), .B1(n1058), .B2(\mem[16][3] ), 
        .ZN(n1055) );
  INV_X1 U350 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U351 ( .A1(data_in[4]), .A2(n838), .B1(n1058), .B2(\mem[16][4] ), 
        .ZN(n1054) );
  INV_X1 U352 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U353 ( .A1(data_in[5]), .A2(n838), .B1(n1058), .B2(\mem[16][5] ), 
        .ZN(n1053) );
  INV_X1 U354 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U355 ( .A1(data_in[6]), .A2(n838), .B1(n1058), .B2(\mem[16][6] ), 
        .ZN(n1052) );
  INV_X1 U356 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U357 ( .A1(data_in[7]), .A2(n838), .B1(n1058), .B2(\mem[16][7] ), 
        .ZN(n1051) );
  INV_X1 U358 ( .A(n1049), .ZN(n750) );
  AOI22_X1 U359 ( .A1(data_in[0]), .A2(n837), .B1(n1048), .B2(\mem[17][0] ), 
        .ZN(n1049) );
  INV_X1 U360 ( .A(n1047), .ZN(n749) );
  AOI22_X1 U361 ( .A1(data_in[1]), .A2(n837), .B1(n1048), .B2(\mem[17][1] ), 
        .ZN(n1047) );
  INV_X1 U362 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U363 ( .A1(data_in[2]), .A2(n837), .B1(n1048), .B2(\mem[17][2] ), 
        .ZN(n1046) );
  INV_X1 U364 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U365 ( .A1(data_in[3]), .A2(n837), .B1(n1048), .B2(\mem[17][3] ), 
        .ZN(n1045) );
  INV_X1 U366 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U367 ( .A1(data_in[4]), .A2(n837), .B1(n1048), .B2(\mem[17][4] ), 
        .ZN(n1044) );
  INV_X1 U368 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U369 ( .A1(data_in[5]), .A2(n837), .B1(n1048), .B2(\mem[17][5] ), 
        .ZN(n1043) );
  INV_X1 U370 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U371 ( .A1(data_in[6]), .A2(n837), .B1(n1048), .B2(\mem[17][6] ), 
        .ZN(n1042) );
  INV_X1 U372 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U373 ( .A1(data_in[7]), .A2(n837), .B1(n1048), .B2(\mem[17][7] ), 
        .ZN(n1041) );
  INV_X1 U374 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U375 ( .A1(data_in[0]), .A2(n836), .B1(n1039), .B2(\mem[18][0] ), 
        .ZN(n1040) );
  INV_X1 U376 ( .A(n1038), .ZN(n741) );
  AOI22_X1 U377 ( .A1(data_in[1]), .A2(n836), .B1(n1039), .B2(\mem[18][1] ), 
        .ZN(n1038) );
  INV_X1 U378 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U379 ( .A1(data_in[2]), .A2(n836), .B1(n1039), .B2(\mem[18][2] ), 
        .ZN(n1037) );
  INV_X1 U380 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U381 ( .A1(data_in[3]), .A2(n836), .B1(n1039), .B2(\mem[18][3] ), 
        .ZN(n1036) );
  INV_X1 U382 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U383 ( .A1(data_in[4]), .A2(n836), .B1(n1039), .B2(\mem[18][4] ), 
        .ZN(n1035) );
  INV_X1 U384 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U385 ( .A1(data_in[5]), .A2(n836), .B1(n1039), .B2(\mem[18][5] ), 
        .ZN(n1034) );
  INV_X1 U386 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U387 ( .A1(data_in[6]), .A2(n836), .B1(n1039), .B2(\mem[18][6] ), 
        .ZN(n1033) );
  INV_X1 U388 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U389 ( .A1(data_in[7]), .A2(n836), .B1(n1039), .B2(\mem[18][7] ), 
        .ZN(n1032) );
  INV_X1 U390 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U391 ( .A1(data_in[0]), .A2(n835), .B1(n1030), .B2(\mem[19][0] ), 
        .ZN(n1031) );
  INV_X1 U392 ( .A(n1029), .ZN(n733) );
  AOI22_X1 U393 ( .A1(data_in[1]), .A2(n835), .B1(n1030), .B2(\mem[19][1] ), 
        .ZN(n1029) );
  INV_X1 U394 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U395 ( .A1(data_in[2]), .A2(n835), .B1(n1030), .B2(\mem[19][2] ), 
        .ZN(n1028) );
  INV_X1 U396 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U397 ( .A1(data_in[3]), .A2(n835), .B1(n1030), .B2(\mem[19][3] ), 
        .ZN(n1027) );
  INV_X1 U398 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U399 ( .A1(data_in[4]), .A2(n835), .B1(n1030), .B2(\mem[19][4] ), 
        .ZN(n1026) );
  INV_X1 U400 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U401 ( .A1(data_in[5]), .A2(n835), .B1(n1030), .B2(\mem[19][5] ), 
        .ZN(n1025) );
  INV_X1 U402 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U403 ( .A1(data_in[6]), .A2(n835), .B1(n1030), .B2(\mem[19][6] ), 
        .ZN(n1024) );
  INV_X1 U404 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U405 ( .A1(data_in[7]), .A2(n835), .B1(n1030), .B2(\mem[19][7] ), 
        .ZN(n1023) );
  INV_X1 U406 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U407 ( .A1(data_in[0]), .A2(n834), .B1(n1021), .B2(\mem[20][0] ), 
        .ZN(n1022) );
  INV_X1 U408 ( .A(n1020), .ZN(n725) );
  AOI22_X1 U409 ( .A1(data_in[1]), .A2(n834), .B1(n1021), .B2(\mem[20][1] ), 
        .ZN(n1020) );
  INV_X1 U410 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U411 ( .A1(data_in[2]), .A2(n834), .B1(n1021), .B2(\mem[20][2] ), 
        .ZN(n1019) );
  INV_X1 U412 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U413 ( .A1(data_in[3]), .A2(n834), .B1(n1021), .B2(\mem[20][3] ), 
        .ZN(n1018) );
  INV_X1 U414 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U415 ( .A1(data_in[4]), .A2(n834), .B1(n1021), .B2(\mem[20][4] ), 
        .ZN(n1017) );
  INV_X1 U416 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U417 ( .A1(data_in[5]), .A2(n834), .B1(n1021), .B2(\mem[20][5] ), 
        .ZN(n1016) );
  INV_X1 U418 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U419 ( .A1(data_in[6]), .A2(n834), .B1(n1021), .B2(\mem[20][6] ), 
        .ZN(n1015) );
  INV_X1 U420 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U421 ( .A1(data_in[7]), .A2(n834), .B1(n1021), .B2(\mem[20][7] ), 
        .ZN(n1014) );
  INV_X1 U422 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U423 ( .A1(data_in[0]), .A2(n833), .B1(n1012), .B2(\mem[21][0] ), 
        .ZN(n1013) );
  INV_X1 U424 ( .A(n1011), .ZN(n717) );
  AOI22_X1 U425 ( .A1(data_in[1]), .A2(n833), .B1(n1012), .B2(\mem[21][1] ), 
        .ZN(n1011) );
  INV_X1 U426 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U427 ( .A1(data_in[2]), .A2(n833), .B1(n1012), .B2(\mem[21][2] ), 
        .ZN(n1010) );
  INV_X1 U428 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U429 ( .A1(data_in[3]), .A2(n833), .B1(n1012), .B2(\mem[21][3] ), 
        .ZN(n1009) );
  INV_X1 U430 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U431 ( .A1(data_in[4]), .A2(n833), .B1(n1012), .B2(\mem[21][4] ), 
        .ZN(n1008) );
  INV_X1 U432 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U433 ( .A1(data_in[5]), .A2(n833), .B1(n1012), .B2(\mem[21][5] ), 
        .ZN(n1007) );
  INV_X1 U434 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U435 ( .A1(data_in[6]), .A2(n833), .B1(n1012), .B2(\mem[21][6] ), 
        .ZN(n1006) );
  INV_X1 U436 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U437 ( .A1(data_in[7]), .A2(n833), .B1(n1012), .B2(\mem[21][7] ), 
        .ZN(n1005) );
  INV_X1 U438 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U439 ( .A1(data_in[0]), .A2(n832), .B1(n1003), .B2(\mem[22][0] ), 
        .ZN(n1004) );
  INV_X1 U440 ( .A(n1002), .ZN(n709) );
  AOI22_X1 U441 ( .A1(data_in[1]), .A2(n832), .B1(n1003), .B2(\mem[22][1] ), 
        .ZN(n1002) );
  INV_X1 U442 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U443 ( .A1(data_in[2]), .A2(n832), .B1(n1003), .B2(\mem[22][2] ), 
        .ZN(n1001) );
  INV_X1 U444 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U445 ( .A1(data_in[3]), .A2(n832), .B1(n1003), .B2(\mem[22][3] ), 
        .ZN(n1000) );
  INV_X1 U446 ( .A(n999), .ZN(n706) );
  AOI22_X1 U447 ( .A1(data_in[4]), .A2(n832), .B1(n1003), .B2(\mem[22][4] ), 
        .ZN(n999) );
  INV_X1 U448 ( .A(n998), .ZN(n705) );
  AOI22_X1 U449 ( .A1(data_in[5]), .A2(n832), .B1(n1003), .B2(\mem[22][5] ), 
        .ZN(n998) );
  INV_X1 U450 ( .A(n997), .ZN(n704) );
  AOI22_X1 U451 ( .A1(data_in[6]), .A2(n832), .B1(n1003), .B2(\mem[22][6] ), 
        .ZN(n997) );
  INV_X1 U452 ( .A(n996), .ZN(n703) );
  AOI22_X1 U453 ( .A1(data_in[7]), .A2(n832), .B1(n1003), .B2(\mem[22][7] ), 
        .ZN(n996) );
  INV_X1 U454 ( .A(n995), .ZN(n702) );
  AOI22_X1 U455 ( .A1(data_in[0]), .A2(n831), .B1(n994), .B2(\mem[23][0] ), 
        .ZN(n995) );
  INV_X1 U456 ( .A(n993), .ZN(n701) );
  AOI22_X1 U457 ( .A1(data_in[1]), .A2(n831), .B1(n994), .B2(\mem[23][1] ), 
        .ZN(n993) );
  INV_X1 U458 ( .A(n992), .ZN(n700) );
  AOI22_X1 U459 ( .A1(data_in[2]), .A2(n831), .B1(n994), .B2(\mem[23][2] ), 
        .ZN(n992) );
  INV_X1 U460 ( .A(n991), .ZN(n699) );
  AOI22_X1 U461 ( .A1(data_in[3]), .A2(n831), .B1(n994), .B2(\mem[23][3] ), 
        .ZN(n991) );
  INV_X1 U462 ( .A(n990), .ZN(n698) );
  AOI22_X1 U463 ( .A1(data_in[4]), .A2(n831), .B1(n994), .B2(\mem[23][4] ), 
        .ZN(n990) );
  INV_X1 U464 ( .A(n989), .ZN(n697) );
  AOI22_X1 U465 ( .A1(data_in[5]), .A2(n831), .B1(n994), .B2(\mem[23][5] ), 
        .ZN(n989) );
  INV_X1 U466 ( .A(n988), .ZN(n696) );
  AOI22_X1 U467 ( .A1(data_in[6]), .A2(n831), .B1(n994), .B2(\mem[23][6] ), 
        .ZN(n988) );
  INV_X1 U468 ( .A(n987), .ZN(n695) );
  AOI22_X1 U469 ( .A1(data_in[7]), .A2(n831), .B1(n994), .B2(\mem[23][7] ), 
        .ZN(n987) );
  INV_X1 U470 ( .A(n986), .ZN(n694) );
  AOI22_X1 U471 ( .A1(data_in[0]), .A2(n830), .B1(n985), .B2(\mem[24][0] ), 
        .ZN(n986) );
  INV_X1 U472 ( .A(n984), .ZN(n693) );
  AOI22_X1 U473 ( .A1(data_in[1]), .A2(n830), .B1(n985), .B2(\mem[24][1] ), 
        .ZN(n984) );
  INV_X1 U474 ( .A(n983), .ZN(n692) );
  AOI22_X1 U475 ( .A1(data_in[2]), .A2(n830), .B1(n985), .B2(\mem[24][2] ), 
        .ZN(n983) );
  INV_X1 U476 ( .A(n982), .ZN(n691) );
  AOI22_X1 U477 ( .A1(data_in[3]), .A2(n830), .B1(n985), .B2(\mem[24][3] ), 
        .ZN(n982) );
  INV_X1 U478 ( .A(n981), .ZN(n690) );
  AOI22_X1 U479 ( .A1(data_in[4]), .A2(n830), .B1(n985), .B2(\mem[24][4] ), 
        .ZN(n981) );
  INV_X1 U480 ( .A(n980), .ZN(n689) );
  AOI22_X1 U481 ( .A1(data_in[5]), .A2(n830), .B1(n985), .B2(\mem[24][5] ), 
        .ZN(n980) );
  INV_X1 U482 ( .A(n979), .ZN(n688) );
  AOI22_X1 U483 ( .A1(data_in[6]), .A2(n830), .B1(n985), .B2(\mem[24][6] ), 
        .ZN(n979) );
  INV_X1 U484 ( .A(n978), .ZN(n687) );
  AOI22_X1 U485 ( .A1(data_in[7]), .A2(n830), .B1(n985), .B2(\mem[24][7] ), 
        .ZN(n978) );
  INV_X1 U486 ( .A(n976), .ZN(n686) );
  AOI22_X1 U487 ( .A1(data_in[0]), .A2(n829), .B1(n975), .B2(\mem[25][0] ), 
        .ZN(n976) );
  INV_X1 U488 ( .A(n974), .ZN(n685) );
  AOI22_X1 U489 ( .A1(data_in[1]), .A2(n829), .B1(n975), .B2(\mem[25][1] ), 
        .ZN(n974) );
  INV_X1 U490 ( .A(n973), .ZN(n684) );
  AOI22_X1 U491 ( .A1(data_in[2]), .A2(n829), .B1(n975), .B2(\mem[25][2] ), 
        .ZN(n973) );
  INV_X1 U492 ( .A(n972), .ZN(n683) );
  AOI22_X1 U493 ( .A1(data_in[3]), .A2(n829), .B1(n975), .B2(\mem[25][3] ), 
        .ZN(n972) );
  INV_X1 U494 ( .A(n971), .ZN(n682) );
  AOI22_X1 U495 ( .A1(data_in[4]), .A2(n829), .B1(n975), .B2(\mem[25][4] ), 
        .ZN(n971) );
  INV_X1 U496 ( .A(n970), .ZN(n681) );
  AOI22_X1 U497 ( .A1(data_in[5]), .A2(n829), .B1(n975), .B2(\mem[25][5] ), 
        .ZN(n970) );
  INV_X1 U498 ( .A(n969), .ZN(n680) );
  AOI22_X1 U499 ( .A1(data_in[6]), .A2(n829), .B1(n975), .B2(\mem[25][6] ), 
        .ZN(n969) );
  INV_X1 U500 ( .A(n968), .ZN(n679) );
  AOI22_X1 U501 ( .A1(data_in[7]), .A2(n829), .B1(n975), .B2(\mem[25][7] ), 
        .ZN(n968) );
  INV_X1 U502 ( .A(n967), .ZN(n678) );
  AOI22_X1 U503 ( .A1(data_in[0]), .A2(n828), .B1(n966), .B2(\mem[26][0] ), 
        .ZN(n967) );
  INV_X1 U504 ( .A(n965), .ZN(n677) );
  AOI22_X1 U505 ( .A1(data_in[1]), .A2(n828), .B1(n966), .B2(\mem[26][1] ), 
        .ZN(n965) );
  INV_X1 U506 ( .A(n964), .ZN(n676) );
  AOI22_X1 U507 ( .A1(data_in[2]), .A2(n828), .B1(n966), .B2(\mem[26][2] ), 
        .ZN(n964) );
  INV_X1 U508 ( .A(n963), .ZN(n675) );
  AOI22_X1 U509 ( .A1(data_in[3]), .A2(n828), .B1(n966), .B2(\mem[26][3] ), 
        .ZN(n963) );
  INV_X1 U510 ( .A(n962), .ZN(n674) );
  AOI22_X1 U511 ( .A1(data_in[4]), .A2(n828), .B1(n966), .B2(\mem[26][4] ), 
        .ZN(n962) );
  INV_X1 U512 ( .A(n961), .ZN(n673) );
  AOI22_X1 U513 ( .A1(data_in[5]), .A2(n828), .B1(n966), .B2(\mem[26][5] ), 
        .ZN(n961) );
  INV_X1 U514 ( .A(n960), .ZN(n672) );
  AOI22_X1 U515 ( .A1(data_in[6]), .A2(n828), .B1(n966), .B2(\mem[26][6] ), 
        .ZN(n960) );
  INV_X1 U516 ( .A(n959), .ZN(n671) );
  AOI22_X1 U517 ( .A1(data_in[7]), .A2(n828), .B1(n966), .B2(\mem[26][7] ), 
        .ZN(n959) );
  INV_X1 U518 ( .A(n958), .ZN(n670) );
  AOI22_X1 U519 ( .A1(data_in[0]), .A2(n827), .B1(n957), .B2(\mem[27][0] ), 
        .ZN(n958) );
  INV_X1 U520 ( .A(n956), .ZN(n669) );
  AOI22_X1 U521 ( .A1(data_in[1]), .A2(n827), .B1(n957), .B2(\mem[27][1] ), 
        .ZN(n956) );
  INV_X1 U522 ( .A(n955), .ZN(n668) );
  AOI22_X1 U523 ( .A1(data_in[2]), .A2(n827), .B1(n957), .B2(\mem[27][2] ), 
        .ZN(n955) );
  INV_X1 U524 ( .A(n954), .ZN(n667) );
  AOI22_X1 U525 ( .A1(data_in[3]), .A2(n827), .B1(n957), .B2(\mem[27][3] ), 
        .ZN(n954) );
  INV_X1 U526 ( .A(n953), .ZN(n666) );
  AOI22_X1 U527 ( .A1(data_in[4]), .A2(n827), .B1(n957), .B2(\mem[27][4] ), 
        .ZN(n953) );
  INV_X1 U528 ( .A(n952), .ZN(n665) );
  AOI22_X1 U529 ( .A1(data_in[5]), .A2(n827), .B1(n957), .B2(\mem[27][5] ), 
        .ZN(n952) );
  INV_X1 U530 ( .A(n951), .ZN(n664) );
  AOI22_X1 U531 ( .A1(data_in[6]), .A2(n827), .B1(n957), .B2(\mem[27][6] ), 
        .ZN(n951) );
  INV_X1 U532 ( .A(n950), .ZN(n663) );
  AOI22_X1 U533 ( .A1(data_in[7]), .A2(n827), .B1(n957), .B2(\mem[27][7] ), 
        .ZN(n950) );
  INV_X1 U534 ( .A(n949), .ZN(n662) );
  AOI22_X1 U535 ( .A1(data_in[0]), .A2(n826), .B1(n948), .B2(\mem[28][0] ), 
        .ZN(n949) );
  INV_X1 U536 ( .A(n947), .ZN(n661) );
  AOI22_X1 U537 ( .A1(data_in[1]), .A2(n826), .B1(n948), .B2(\mem[28][1] ), 
        .ZN(n947) );
  INV_X1 U538 ( .A(n946), .ZN(n660) );
  AOI22_X1 U539 ( .A1(data_in[2]), .A2(n826), .B1(n948), .B2(\mem[28][2] ), 
        .ZN(n946) );
  INV_X1 U540 ( .A(n945), .ZN(n659) );
  AOI22_X1 U541 ( .A1(data_in[3]), .A2(n826), .B1(n948), .B2(\mem[28][3] ), 
        .ZN(n945) );
  INV_X1 U542 ( .A(n944), .ZN(n658) );
  AOI22_X1 U543 ( .A1(data_in[4]), .A2(n826), .B1(n948), .B2(\mem[28][4] ), 
        .ZN(n944) );
  INV_X1 U544 ( .A(n943), .ZN(n657) );
  AOI22_X1 U545 ( .A1(data_in[5]), .A2(n826), .B1(n948), .B2(\mem[28][5] ), 
        .ZN(n943) );
  INV_X1 U546 ( .A(n942), .ZN(n656) );
  AOI22_X1 U547 ( .A1(data_in[6]), .A2(n826), .B1(n948), .B2(\mem[28][6] ), 
        .ZN(n942) );
  INV_X1 U548 ( .A(n941), .ZN(n655) );
  AOI22_X1 U549 ( .A1(data_in[7]), .A2(n826), .B1(n948), .B2(\mem[28][7] ), 
        .ZN(n941) );
  INV_X1 U550 ( .A(n940), .ZN(n654) );
  AOI22_X1 U551 ( .A1(data_in[0]), .A2(n825), .B1(n939), .B2(\mem[29][0] ), 
        .ZN(n940) );
  INV_X1 U552 ( .A(n938), .ZN(n653) );
  AOI22_X1 U553 ( .A1(data_in[1]), .A2(n825), .B1(n939), .B2(\mem[29][1] ), 
        .ZN(n938) );
  INV_X1 U554 ( .A(n937), .ZN(n652) );
  AOI22_X1 U555 ( .A1(data_in[2]), .A2(n825), .B1(n939), .B2(\mem[29][2] ), 
        .ZN(n937) );
  INV_X1 U556 ( .A(n936), .ZN(n651) );
  AOI22_X1 U557 ( .A1(data_in[3]), .A2(n825), .B1(n939), .B2(\mem[29][3] ), 
        .ZN(n936) );
  INV_X1 U558 ( .A(n935), .ZN(n650) );
  AOI22_X1 U559 ( .A1(data_in[4]), .A2(n825), .B1(n939), .B2(\mem[29][4] ), 
        .ZN(n935) );
  INV_X1 U560 ( .A(n934), .ZN(n649) );
  AOI22_X1 U561 ( .A1(data_in[5]), .A2(n825), .B1(n939), .B2(\mem[29][5] ), 
        .ZN(n934) );
  INV_X1 U562 ( .A(n933), .ZN(n648) );
  AOI22_X1 U563 ( .A1(data_in[6]), .A2(n825), .B1(n939), .B2(\mem[29][6] ), 
        .ZN(n933) );
  INV_X1 U564 ( .A(n932), .ZN(n647) );
  AOI22_X1 U565 ( .A1(data_in[7]), .A2(n825), .B1(n939), .B2(\mem[29][7] ), 
        .ZN(n932) );
  INV_X1 U566 ( .A(n931), .ZN(n646) );
  AOI22_X1 U567 ( .A1(data_in[0]), .A2(n824), .B1(n930), .B2(\mem[30][0] ), 
        .ZN(n931) );
  INV_X1 U568 ( .A(n929), .ZN(n645) );
  AOI22_X1 U569 ( .A1(data_in[1]), .A2(n824), .B1(n930), .B2(\mem[30][1] ), 
        .ZN(n929) );
  INV_X1 U570 ( .A(n928), .ZN(n644) );
  AOI22_X1 U571 ( .A1(data_in[2]), .A2(n824), .B1(n930), .B2(\mem[30][2] ), 
        .ZN(n928) );
  INV_X1 U572 ( .A(n927), .ZN(n643) );
  AOI22_X1 U573 ( .A1(data_in[3]), .A2(n824), .B1(n930), .B2(\mem[30][3] ), 
        .ZN(n927) );
  INV_X1 U574 ( .A(n926), .ZN(n642) );
  AOI22_X1 U575 ( .A1(data_in[4]), .A2(n824), .B1(n930), .B2(\mem[30][4] ), 
        .ZN(n926) );
  INV_X1 U576 ( .A(n925), .ZN(n641) );
  AOI22_X1 U577 ( .A1(data_in[5]), .A2(n824), .B1(n930), .B2(\mem[30][5] ), 
        .ZN(n925) );
  INV_X1 U578 ( .A(n924), .ZN(n640) );
  AOI22_X1 U579 ( .A1(data_in[6]), .A2(n824), .B1(n930), .B2(\mem[30][6] ), 
        .ZN(n924) );
  INV_X1 U580 ( .A(n923), .ZN(n639) );
  AOI22_X1 U581 ( .A1(data_in[7]), .A2(n824), .B1(n930), .B2(\mem[30][7] ), 
        .ZN(n923) );
  INV_X1 U582 ( .A(n922), .ZN(n638) );
  AOI22_X1 U583 ( .A1(data_in[0]), .A2(n823), .B1(n921), .B2(\mem[31][0] ), 
        .ZN(n922) );
  INV_X1 U584 ( .A(n920), .ZN(n637) );
  AOI22_X1 U585 ( .A1(data_in[1]), .A2(n823), .B1(n921), .B2(\mem[31][1] ), 
        .ZN(n920) );
  INV_X1 U586 ( .A(n919), .ZN(n636) );
  AOI22_X1 U587 ( .A1(data_in[2]), .A2(n823), .B1(n921), .B2(\mem[31][2] ), 
        .ZN(n919) );
  INV_X1 U588 ( .A(n918), .ZN(n635) );
  AOI22_X1 U589 ( .A1(data_in[3]), .A2(n823), .B1(n921), .B2(\mem[31][3] ), 
        .ZN(n918) );
  INV_X1 U590 ( .A(n917), .ZN(n634) );
  AOI22_X1 U591 ( .A1(data_in[4]), .A2(n823), .B1(n921), .B2(\mem[31][4] ), 
        .ZN(n917) );
  INV_X1 U592 ( .A(n916), .ZN(n633) );
  AOI22_X1 U593 ( .A1(data_in[5]), .A2(n823), .B1(n921), .B2(\mem[31][5] ), 
        .ZN(n916) );
  INV_X1 U594 ( .A(n915), .ZN(n632) );
  AOI22_X1 U595 ( .A1(data_in[6]), .A2(n823), .B1(n921), .B2(\mem[31][6] ), 
        .ZN(n915) );
  INV_X1 U596 ( .A(n914), .ZN(n631) );
  AOI22_X1 U597 ( .A1(data_in[7]), .A2(n823), .B1(n921), .B2(\mem[31][7] ), 
        .ZN(n914) );
  MUX2_X1 U598 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n615), .Z(n5) );
  MUX2_X1 U599 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n615), .Z(n6) );
  MUX2_X1 U600 ( .A(n6), .B(n5), .S(n612), .Z(n7) );
  MUX2_X1 U601 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n615), .Z(n8) );
  MUX2_X1 U602 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n615), .Z(n9) );
  MUX2_X1 U603 ( .A(n9), .B(n8), .S(n612), .Z(n10) );
  MUX2_X1 U604 ( .A(n10), .B(n7), .S(n610), .Z(n11) );
  MUX2_X1 U605 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n615), .Z(n12) );
  MUX2_X1 U606 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n615), .Z(n13) );
  MUX2_X1 U607 ( .A(n13), .B(n12), .S(n612), .Z(n14) );
  MUX2_X1 U608 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n615), .Z(n15) );
  MUX2_X1 U609 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n615), .Z(n16) );
  MUX2_X1 U610 ( .A(n16), .B(n15), .S(n612), .Z(n17) );
  MUX2_X1 U611 ( .A(n17), .B(n14), .S(n610), .Z(n18) );
  MUX2_X1 U612 ( .A(n18), .B(n11), .S(N13), .Z(n19) );
  MUX2_X1 U613 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n616), .Z(n20) );
  MUX2_X1 U614 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n616), .Z(n21) );
  MUX2_X1 U615 ( .A(n21), .B(n20), .S(n613), .Z(n22) );
  MUX2_X1 U616 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n616), .Z(n23) );
  MUX2_X1 U617 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n616), .Z(n24) );
  MUX2_X1 U618 ( .A(n24), .B(n23), .S(n613), .Z(n25) );
  MUX2_X1 U619 ( .A(n25), .B(n22), .S(n610), .Z(n26) );
  MUX2_X1 U620 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n616), .Z(n27) );
  MUX2_X1 U621 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n616), .Z(n28) );
  MUX2_X1 U622 ( .A(n28), .B(n27), .S(n613), .Z(n29) );
  MUX2_X1 U623 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n616), .Z(n30) );
  MUX2_X1 U624 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n616), .Z(n31) );
  MUX2_X1 U625 ( .A(n31), .B(n30), .S(n613), .Z(n32) );
  MUX2_X1 U626 ( .A(n32), .B(n29), .S(n610), .Z(n33) );
  MUX2_X1 U627 ( .A(n33), .B(n26), .S(N13), .Z(n34) );
  MUX2_X1 U628 ( .A(n34), .B(n19), .S(N14), .Z(N22) );
  MUX2_X1 U629 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n616), .Z(n35) );
  MUX2_X1 U630 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n616), .Z(n36) );
  MUX2_X1 U631 ( .A(n36), .B(n35), .S(n613), .Z(n37) );
  MUX2_X1 U632 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n616), .Z(n38) );
  MUX2_X1 U633 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n616), .Z(n39) );
  MUX2_X1 U634 ( .A(n39), .B(n38), .S(n613), .Z(n40) );
  MUX2_X1 U635 ( .A(n40), .B(n37), .S(n610), .Z(n41) );
  MUX2_X1 U636 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n617), .Z(n42) );
  MUX2_X1 U637 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n617), .Z(n43) );
  MUX2_X1 U638 ( .A(n43), .B(n42), .S(n613), .Z(n44) );
  MUX2_X1 U639 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n617), .Z(n45) );
  MUX2_X1 U640 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n617), .Z(n46) );
  MUX2_X1 U641 ( .A(n46), .B(n45), .S(n613), .Z(n47) );
  MUX2_X1 U642 ( .A(n47), .B(n44), .S(n610), .Z(n48) );
  MUX2_X1 U643 ( .A(n48), .B(n41), .S(N13), .Z(n49) );
  MUX2_X1 U644 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n617), .Z(n50) );
  MUX2_X1 U645 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n617), .Z(n51) );
  MUX2_X1 U646 ( .A(n51), .B(n50), .S(n613), .Z(n52) );
  MUX2_X1 U647 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n617), .Z(n53) );
  MUX2_X1 U648 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n617), .Z(n54) );
  MUX2_X1 U649 ( .A(n54), .B(n53), .S(n613), .Z(n55) );
  MUX2_X1 U650 ( .A(n55), .B(n52), .S(n610), .Z(n56) );
  MUX2_X1 U651 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n617), .Z(n57) );
  MUX2_X1 U652 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n617), .Z(n58) );
  MUX2_X1 U653 ( .A(n58), .B(n57), .S(n613), .Z(n59) );
  MUX2_X1 U654 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n617), .Z(n60) );
  MUX2_X1 U655 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n617), .Z(n61) );
  MUX2_X1 U656 ( .A(n61), .B(n60), .S(n613), .Z(n62) );
  MUX2_X1 U657 ( .A(n62), .B(n59), .S(n610), .Z(n63) );
  MUX2_X1 U658 ( .A(n63), .B(n56), .S(N13), .Z(n64) );
  MUX2_X1 U659 ( .A(n64), .B(n49), .S(N14), .Z(N21) );
  MUX2_X1 U660 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n618), .Z(n65) );
  MUX2_X1 U661 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n618), .Z(n66) );
  MUX2_X1 U662 ( .A(n66), .B(n65), .S(n614), .Z(n67) );
  MUX2_X1 U663 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n618), .Z(n68) );
  MUX2_X1 U664 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n618), .Z(n69) );
  MUX2_X1 U665 ( .A(n69), .B(n68), .S(n614), .Z(n70) );
  MUX2_X1 U666 ( .A(n70), .B(n67), .S(n610), .Z(n71) );
  MUX2_X1 U667 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n618), .Z(n72) );
  MUX2_X1 U668 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n618), .Z(n73) );
  MUX2_X1 U669 ( .A(n73), .B(n72), .S(n614), .Z(n74) );
  MUX2_X1 U670 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n618), .Z(n75) );
  MUX2_X1 U671 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n618), .Z(n76) );
  MUX2_X1 U672 ( .A(n76), .B(n75), .S(n614), .Z(n77) );
  MUX2_X1 U673 ( .A(n77), .B(n74), .S(N12), .Z(n78) );
  MUX2_X1 U674 ( .A(n78), .B(n71), .S(N13), .Z(n79) );
  MUX2_X1 U675 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n618), .Z(n80) );
  MUX2_X1 U676 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n618), .Z(n81) );
  MUX2_X1 U677 ( .A(n81), .B(n80), .S(n614), .Z(n82) );
  MUX2_X1 U678 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n618), .Z(n83) );
  MUX2_X1 U679 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n618), .Z(n84) );
  MUX2_X1 U680 ( .A(n84), .B(n83), .S(n614), .Z(n85) );
  MUX2_X1 U681 ( .A(n85), .B(n82), .S(n610), .Z(n86) );
  MUX2_X1 U682 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n616), .Z(n87) );
  MUX2_X1 U683 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n617), .Z(n88) );
  MUX2_X1 U684 ( .A(n88), .B(n87), .S(n614), .Z(n89) );
  MUX2_X1 U685 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n615), .Z(n90) );
  MUX2_X1 U686 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n615), .Z(n91) );
  MUX2_X1 U687 ( .A(n91), .B(n90), .S(n614), .Z(n92) );
  MUX2_X1 U688 ( .A(n92), .B(n89), .S(n611), .Z(n93) );
  MUX2_X1 U689 ( .A(n93), .B(n86), .S(N13), .Z(n94) );
  MUX2_X1 U690 ( .A(n94), .B(n79), .S(N14), .Z(N20) );
  MUX2_X1 U691 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n618), .Z(n95) );
  MUX2_X1 U692 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n617), .Z(n96) );
  MUX2_X1 U693 ( .A(n96), .B(n95), .S(n614), .Z(n97) );
  MUX2_X1 U694 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n616), .Z(n98) );
  MUX2_X1 U695 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n617), .Z(n99) );
  MUX2_X1 U696 ( .A(n99), .B(n98), .S(n614), .Z(n100) );
  MUX2_X1 U697 ( .A(n100), .B(n97), .S(n610), .Z(n101) );
  MUX2_X1 U698 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n615), .Z(n102) );
  MUX2_X1 U699 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n618), .Z(n103) );
  MUX2_X1 U700 ( .A(n103), .B(n102), .S(n614), .Z(n104) );
  MUX2_X1 U701 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n615), .Z(n105) );
  MUX2_X1 U702 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n618), .Z(n106) );
  MUX2_X1 U703 ( .A(n106), .B(n105), .S(n614), .Z(n107) );
  MUX2_X1 U704 ( .A(n107), .B(n104), .S(N12), .Z(n108) );
  MUX2_X1 U705 ( .A(n108), .B(n101), .S(N13), .Z(n109) );
  MUX2_X1 U706 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n617), .Z(n110) );
  MUX2_X1 U707 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n620), .Z(n111) );
  MUX2_X1 U708 ( .A(n111), .B(n110), .S(n613), .Z(n112) );
  MUX2_X1 U709 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n619), .Z(n113) );
  MUX2_X1 U710 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n619), .Z(n114) );
  MUX2_X1 U711 ( .A(n114), .B(n113), .S(n613), .Z(n115) );
  MUX2_X1 U712 ( .A(n115), .B(n112), .S(n611), .Z(n116) );
  MUX2_X1 U713 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n620), .Z(n117) );
  MUX2_X1 U714 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n620), .Z(n118) );
  MUX2_X1 U715 ( .A(n118), .B(n117), .S(n614), .Z(n119) );
  MUX2_X1 U716 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n616), .Z(n120) );
  MUX2_X1 U717 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n618), .Z(n121) );
  MUX2_X1 U718 ( .A(n121), .B(n120), .S(n612), .Z(n122) );
  MUX2_X1 U719 ( .A(n122), .B(n119), .S(n610), .Z(n123) );
  MUX2_X1 U720 ( .A(n123), .B(n116), .S(N13), .Z(n124) );
  MUX2_X1 U721 ( .A(n124), .B(n109), .S(N14), .Z(N19) );
  MUX2_X1 U722 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n620), .Z(n125) );
  MUX2_X1 U723 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n620), .Z(n126) );
  MUX2_X1 U724 ( .A(n126), .B(n125), .S(n612), .Z(n127) );
  MUX2_X1 U725 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n617), .Z(n128) );
  MUX2_X1 U726 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n619), .Z(n129) );
  MUX2_X1 U727 ( .A(n129), .B(n128), .S(n613), .Z(n130) );
  MUX2_X1 U728 ( .A(n130), .B(n127), .S(n610), .Z(n131) );
  MUX2_X1 U729 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n620), .Z(n132) );
  MUX2_X1 U730 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n620), .Z(n133) );
  MUX2_X1 U731 ( .A(n133), .B(n132), .S(N11), .Z(n134) );
  MUX2_X1 U732 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n619), .Z(n135) );
  MUX2_X1 U733 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n619), .Z(n136) );
  MUX2_X1 U734 ( .A(n136), .B(n135), .S(n613), .Z(n137) );
  MUX2_X1 U735 ( .A(n137), .B(n134), .S(N12), .Z(n138) );
  MUX2_X1 U736 ( .A(n138), .B(n131), .S(N13), .Z(n139) );
  MUX2_X1 U737 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n619), .Z(n140) );
  MUX2_X1 U738 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n619), .Z(n141) );
  MUX2_X1 U739 ( .A(n141), .B(n140), .S(n614), .Z(n142) );
  MUX2_X1 U740 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n620), .Z(n143) );
  MUX2_X1 U741 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n620), .Z(n144) );
  MUX2_X1 U742 ( .A(n144), .B(n143), .S(n614), .Z(n145) );
  MUX2_X1 U743 ( .A(n145), .B(n142), .S(n610), .Z(n146) );
  MUX2_X1 U744 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n620), .Z(n147) );
  MUX2_X1 U745 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n619), .Z(n148) );
  MUX2_X1 U746 ( .A(n148), .B(n147), .S(n612), .Z(n149) );
  MUX2_X1 U747 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n620), .Z(n150) );
  MUX2_X1 U748 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n619), .Z(n151) );
  MUX2_X1 U749 ( .A(n151), .B(n150), .S(n613), .Z(n152) );
  MUX2_X1 U750 ( .A(n152), .B(n149), .S(n611), .Z(n153) );
  MUX2_X1 U751 ( .A(n153), .B(n146), .S(N13), .Z(n154) );
  MUX2_X1 U752 ( .A(n154), .B(n139), .S(N14), .Z(N18) );
  MUX2_X1 U753 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n620), .Z(n155) );
  MUX2_X1 U754 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(N10), .Z(n156) );
  MUX2_X1 U755 ( .A(n156), .B(n155), .S(n613), .Z(n157) );
  MUX2_X1 U756 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(N10), .Z(n158) );
  MUX2_X1 U757 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(N10), .Z(n159) );
  MUX2_X1 U758 ( .A(n159), .B(n158), .S(N11), .Z(n160) );
  MUX2_X1 U759 ( .A(n160), .B(n157), .S(n611), .Z(n161) );
  MUX2_X1 U760 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n615), .Z(n162) );
  MUX2_X1 U761 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n620), .Z(n163) );
  MUX2_X1 U762 ( .A(n163), .B(n162), .S(n612), .Z(n164) );
  MUX2_X1 U763 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(N10), .Z(n165) );
  MUX2_X1 U764 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(N10), .Z(n166) );
  MUX2_X1 U765 ( .A(n166), .B(n165), .S(N11), .Z(n167) );
  MUX2_X1 U766 ( .A(n167), .B(n164), .S(n611), .Z(n168) );
  MUX2_X1 U767 ( .A(n168), .B(n161), .S(N13), .Z(n169) );
  MUX2_X1 U768 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n615), .Z(n170) );
  MUX2_X1 U769 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n619), .Z(n171) );
  MUX2_X1 U770 ( .A(n171), .B(n170), .S(n612), .Z(n172) );
  MUX2_X1 U771 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n615), .Z(n173) );
  MUX2_X1 U772 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n619), .Z(n174) );
  MUX2_X1 U773 ( .A(n174), .B(n173), .S(n612), .Z(n175) );
  MUX2_X1 U774 ( .A(n175), .B(n172), .S(n611), .Z(n176) );
  MUX2_X1 U775 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n615), .Z(n177) );
  MUX2_X1 U776 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n616), .Z(n178) );
  MUX2_X1 U777 ( .A(n178), .B(n177), .S(n614), .Z(n179) );
  MUX2_X1 U778 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n616), .Z(n180) );
  MUX2_X1 U779 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n615), .Z(n181) );
  MUX2_X1 U780 ( .A(n181), .B(n180), .S(n613), .Z(n182) );
  MUX2_X1 U781 ( .A(n182), .B(n179), .S(n611), .Z(n183) );
  MUX2_X1 U782 ( .A(n183), .B(n176), .S(N13), .Z(n184) );
  MUX2_X1 U783 ( .A(n184), .B(n169), .S(N14), .Z(N17) );
  MUX2_X1 U784 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n618), .Z(n185) );
  MUX2_X1 U785 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n617), .Z(n186) );
  MUX2_X1 U786 ( .A(n186), .B(n185), .S(n614), .Z(n187) );
  MUX2_X1 U787 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n615), .Z(n188) );
  MUX2_X1 U788 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n616), .Z(n189) );
  MUX2_X1 U789 ( .A(n189), .B(n188), .S(n613), .Z(n190) );
  MUX2_X1 U790 ( .A(n190), .B(n187), .S(n611), .Z(n191) );
  MUX2_X1 U791 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n616), .Z(n192) );
  MUX2_X1 U792 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n618), .Z(n193) );
  MUX2_X1 U793 ( .A(n193), .B(n192), .S(N11), .Z(n194) );
  MUX2_X1 U794 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n618), .Z(n195) );
  MUX2_X1 U795 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n617), .Z(n196) );
  MUX2_X1 U796 ( .A(n196), .B(n195), .S(N11), .Z(n197) );
  MUX2_X1 U797 ( .A(n197), .B(n194), .S(n611), .Z(n198) );
  MUX2_X1 U798 ( .A(n198), .B(n191), .S(N13), .Z(n199) );
  MUX2_X1 U799 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n619), .Z(n200) );
  MUX2_X1 U800 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n619), .Z(n201) );
  MUX2_X1 U801 ( .A(n201), .B(n200), .S(n612), .Z(n202) );
  MUX2_X1 U802 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n619), .Z(n203) );
  MUX2_X1 U803 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n618), .Z(n204) );
  MUX2_X1 U804 ( .A(n204), .B(n203), .S(n613), .Z(n205) );
  MUX2_X1 U805 ( .A(n205), .B(n202), .S(n611), .Z(n206) );
  MUX2_X1 U806 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n619), .Z(n207) );
  MUX2_X1 U807 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n620), .Z(n208) );
  MUX2_X1 U808 ( .A(n208), .B(n207), .S(n612), .Z(n209) );
  MUX2_X1 U809 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n617), .Z(n210) );
  MUX2_X1 U810 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n616), .Z(n211) );
  MUX2_X1 U811 ( .A(n211), .B(n210), .S(n614), .Z(n212) );
  MUX2_X1 U812 ( .A(n212), .B(n209), .S(n611), .Z(n213) );
  MUX2_X1 U813 ( .A(n213), .B(n206), .S(N13), .Z(n214) );
  MUX2_X1 U814 ( .A(n214), .B(n199), .S(N14), .Z(N16) );
  MUX2_X1 U815 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n620), .Z(n215) );
  MUX2_X1 U816 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n620), .Z(n216) );
  MUX2_X1 U817 ( .A(n216), .B(n215), .S(n612), .Z(n217) );
  MUX2_X1 U818 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n615), .Z(n218) );
  MUX2_X1 U819 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n620), .Z(n219) );
  MUX2_X1 U820 ( .A(n219), .B(n218), .S(n612), .Z(n220) );
  MUX2_X1 U821 ( .A(n220), .B(n217), .S(n611), .Z(n221) );
  MUX2_X1 U822 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n620), .Z(n222) );
  MUX2_X1 U823 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n620), .Z(n223) );
  MUX2_X1 U824 ( .A(n223), .B(n222), .S(n612), .Z(n224) );
  MUX2_X1 U825 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n619), .Z(n225) );
  MUX2_X1 U826 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n619), .Z(n226) );
  MUX2_X1 U827 ( .A(n226), .B(n225), .S(n614), .Z(n227) );
  MUX2_X1 U828 ( .A(n227), .B(n224), .S(n611), .Z(n228) );
  MUX2_X1 U829 ( .A(n228), .B(n221), .S(N13), .Z(n229) );
  MUX2_X1 U830 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n620), .Z(n595) );
  MUX2_X1 U831 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n619), .Z(n596) );
  MUX2_X1 U832 ( .A(n596), .B(n595), .S(n612), .Z(n597) );
  MUX2_X1 U833 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n620), .Z(n598) );
  MUX2_X1 U834 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n620), .Z(n599) );
  MUX2_X1 U835 ( .A(n599), .B(n598), .S(n614), .Z(n600) );
  MUX2_X1 U836 ( .A(n600), .B(n597), .S(n611), .Z(n601) );
  MUX2_X1 U837 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n615), .Z(n602) );
  MUX2_X1 U838 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n620), .Z(n603) );
  MUX2_X1 U839 ( .A(n603), .B(n602), .S(n612), .Z(n604) );
  MUX2_X1 U840 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n619), .Z(n605) );
  MUX2_X1 U841 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n619), .Z(n606) );
  MUX2_X1 U842 ( .A(n606), .B(n605), .S(n612), .Z(n607) );
  MUX2_X1 U843 ( .A(n607), .B(n604), .S(n611), .Z(n608) );
  MUX2_X1 U844 ( .A(n608), .B(n601), .S(N13), .Z(n609) );
  MUX2_X1 U845 ( .A(n609), .B(n229), .S(N14), .Z(N15) );
  CLKBUF_X1 U846 ( .A(N11), .Z(n612) );
  INV_X1 U847 ( .A(N10), .ZN(n621) );
  INV_X1 U848 ( .A(N11), .ZN(n622) );
  INV_X1 U849 ( .A(data_in[0]), .ZN(n623) );
  INV_X1 U850 ( .A(data_in[1]), .ZN(n624) );
  INV_X1 U851 ( .A(data_in[2]), .ZN(n625) );
  INV_X1 U852 ( .A(data_in[3]), .ZN(n626) );
  INV_X1 U853 ( .A(data_in[4]), .ZN(n627) );
  INV_X1 U854 ( .A(data_in[5]), .ZN(n628) );
  INV_X1 U855 ( .A(data_in[6]), .ZN(n629) );
  INV_X1 U856 ( .A(data_in[7]), .ZN(n630) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_22 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n2) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n631), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n632), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n633), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n634), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n635), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n636), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n637), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n638), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n639), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n640), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n641), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n642), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n643), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n644), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n645), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n646), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n647), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n648), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n649), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n650), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n651), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n652), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n653), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n654), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n655), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n656), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n657), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n658), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n659), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n660), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n661), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n662), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n663), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n664), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n665), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n666), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n667), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n668), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n669), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n670), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n671), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n672), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n673), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n674), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n675), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n676), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n677), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n678), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n679), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n680), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n681), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n682), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n683), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n684), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n685), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n686), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n687), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n688), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n689), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n690), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n691), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n692), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n693), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n694), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n695), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n696), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n697), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n698), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n699), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n700), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n701), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n702), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n703), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n704), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n705), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n706), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n707), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n708), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n709), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n710), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n711), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n712), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n713), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n714), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n715), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n716), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n717), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n718), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n719), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n720), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n721), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n722), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n723), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n724), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n725), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n726), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n727), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n728), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n729), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n730), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n731), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n732), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n733), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n734), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n735), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n736), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n737), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n738), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n739), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n740), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n741), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n742), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n743), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n744), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n745), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n746), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n747), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n748), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n749), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n750), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n751), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n752), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n753), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n754), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n755), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n756), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n757), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n758), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n759), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n760), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n761), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n762), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n763), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n764), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n765), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n766), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n767), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n768), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n769), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n770), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n771), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n772), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n773), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n774), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n775), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n776), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n777), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n778), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n779), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n780), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n781), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n782), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n783), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n784), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n785), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n786), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n787), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n788), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n789), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n790), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n791), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n792), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n793), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n794), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n795), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n796), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n797), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n798), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n799), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n800), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n801), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n802), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n803), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n804), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n805), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n806), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n807), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n808), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n809), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n810), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n811), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n812), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n813), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n814), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n815), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n816), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n817), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n818), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n819), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n820), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n821), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n822), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n850), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n851), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n852), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n853), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n854), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n855), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n856), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n857), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n858), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n859), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n860), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n861), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n862), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n863), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n864), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n865), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n866), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n867), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n868), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n869), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n870), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n871), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n872), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n873), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n874), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n875), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n876), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n877), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n878), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n879), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n880), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n881), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n882), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n883), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n884), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n885), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n886), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n887), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n888), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n889), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n890), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n891), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n892), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n893), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n894), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n895), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n896), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n897), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n898), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n899), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n900), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n901), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n902), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n903), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n904), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n905), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n906), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n907), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n908), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n909), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n910), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n911), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n912), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n913), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  CLKBUF_X1 U3 ( .A(n620), .Z(n618) );
  CLKBUF_X1 U4 ( .A(n620), .Z(n615) );
  CLKBUF_X1 U5 ( .A(n620), .Z(n616) );
  INV_X2 U6 ( .A(n2), .ZN(data_out[3]) );
  BUF_X1 U7 ( .A(N10), .Z(n619) );
  BUF_X1 U8 ( .A(N10), .Z(n617) );
  BUF_X1 U9 ( .A(N11), .Z(n612) );
  BUF_X1 U10 ( .A(N11), .Z(n613) );
  BUF_X1 U11 ( .A(N10), .Z(n620) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1205) );
  NOR3_X1 U13 ( .A1(N11), .A2(N12), .A3(n621), .ZN(n1194) );
  NOR3_X1 U14 ( .A1(N10), .A2(N12), .A3(n622), .ZN(n1184) );
  NOR3_X1 U15 ( .A1(n621), .A2(N12), .A3(n622), .ZN(n1174) );
  INV_X1 U16 ( .A(n1131), .ZN(n846) );
  INV_X1 U17 ( .A(n1121), .ZN(n845) );
  INV_X1 U18 ( .A(n1112), .ZN(n844) );
  INV_X1 U19 ( .A(n1103), .ZN(n843) );
  INV_X1 U20 ( .A(n1058), .ZN(n838) );
  INV_X1 U21 ( .A(n1048), .ZN(n837) );
  INV_X1 U22 ( .A(n1039), .ZN(n836) );
  INV_X1 U23 ( .A(n1030), .ZN(n835) );
  INV_X1 U24 ( .A(n985), .ZN(n830) );
  INV_X1 U25 ( .A(n975), .ZN(n829) );
  INV_X1 U26 ( .A(n966), .ZN(n828) );
  INV_X1 U27 ( .A(n957), .ZN(n827) );
  INV_X1 U28 ( .A(n1094), .ZN(n842) );
  INV_X1 U29 ( .A(n1085), .ZN(n841) );
  INV_X1 U30 ( .A(n1076), .ZN(n840) );
  INV_X1 U31 ( .A(n1067), .ZN(n839) );
  INV_X1 U32 ( .A(n948), .ZN(n826) );
  INV_X1 U33 ( .A(n939), .ZN(n825) );
  INV_X1 U34 ( .A(n930), .ZN(n824) );
  INV_X1 U35 ( .A(n921), .ZN(n823) );
  INV_X1 U36 ( .A(n1021), .ZN(n834) );
  INV_X1 U37 ( .A(n1012), .ZN(n833) );
  INV_X1 U38 ( .A(n1003), .ZN(n832) );
  INV_X1 U39 ( .A(n994), .ZN(n831) );
  BUF_X1 U40 ( .A(N12), .Z(n609) );
  BUF_X1 U41 ( .A(N12), .Z(n610) );
  INV_X1 U42 ( .A(N13), .ZN(n848) );
  AND3_X1 U43 ( .A1(n621), .A2(n622), .A3(N12), .ZN(n1164) );
  AND3_X1 U44 ( .A1(N10), .A2(n622), .A3(N12), .ZN(n1154) );
  AND3_X1 U45 ( .A1(N11), .A2(n621), .A3(N12), .ZN(n1144) );
  AND3_X1 U46 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1134) );
  INV_X1 U47 ( .A(N14), .ZN(n849) );
  NAND2_X1 U48 ( .A1(n1194), .A2(n1204), .ZN(n1203) );
  NAND2_X1 U49 ( .A1(n1184), .A2(n1204), .ZN(n1193) );
  NAND2_X1 U50 ( .A1(n1174), .A2(n1204), .ZN(n1183) );
  NAND2_X1 U51 ( .A1(n1164), .A2(n1204), .ZN(n1173) );
  NAND2_X1 U52 ( .A1(n1154), .A2(n1204), .ZN(n1163) );
  NAND2_X1 U53 ( .A1(n1144), .A2(n1204), .ZN(n1153) );
  NAND2_X1 U54 ( .A1(n1134), .A2(n1204), .ZN(n1143) );
  NAND2_X1 U55 ( .A1(n1205), .A2(n1204), .ZN(n1214) );
  NAND2_X1 U56 ( .A1(n1123), .A2(n1205), .ZN(n1131) );
  NAND2_X1 U57 ( .A1(n1123), .A2(n1194), .ZN(n1121) );
  NAND2_X1 U58 ( .A1(n1123), .A2(n1184), .ZN(n1112) );
  NAND2_X1 U59 ( .A1(n1123), .A2(n1174), .ZN(n1103) );
  NAND2_X1 U60 ( .A1(n1050), .A2(n1205), .ZN(n1058) );
  NAND2_X1 U61 ( .A1(n1050), .A2(n1194), .ZN(n1048) );
  NAND2_X1 U62 ( .A1(n1050), .A2(n1184), .ZN(n1039) );
  NAND2_X1 U63 ( .A1(n1050), .A2(n1174), .ZN(n1030) );
  NAND2_X1 U64 ( .A1(n977), .A2(n1205), .ZN(n985) );
  NAND2_X1 U65 ( .A1(n977), .A2(n1194), .ZN(n975) );
  NAND2_X1 U66 ( .A1(n977), .A2(n1184), .ZN(n966) );
  NAND2_X1 U67 ( .A1(n977), .A2(n1174), .ZN(n957) );
  NAND2_X1 U68 ( .A1(n1123), .A2(n1164), .ZN(n1094) );
  NAND2_X1 U69 ( .A1(n1123), .A2(n1154), .ZN(n1085) );
  NAND2_X1 U70 ( .A1(n1123), .A2(n1144), .ZN(n1076) );
  NAND2_X1 U71 ( .A1(n1123), .A2(n1134), .ZN(n1067) );
  NAND2_X1 U72 ( .A1(n1050), .A2(n1164), .ZN(n1021) );
  NAND2_X1 U73 ( .A1(n1050), .A2(n1154), .ZN(n1012) );
  NAND2_X1 U74 ( .A1(n1050), .A2(n1144), .ZN(n1003) );
  NAND2_X1 U75 ( .A1(n1050), .A2(n1134), .ZN(n994) );
  NAND2_X1 U76 ( .A1(n977), .A2(n1164), .ZN(n948) );
  NAND2_X1 U77 ( .A1(n977), .A2(n1154), .ZN(n939) );
  NAND2_X1 U78 ( .A1(n977), .A2(n1144), .ZN(n930) );
  NAND2_X1 U79 ( .A1(n977), .A2(n1134), .ZN(n921) );
  AND3_X1 U80 ( .A1(n848), .A2(n849), .A3(n1133), .ZN(n1204) );
  AND3_X1 U81 ( .A1(N13), .A2(n1133), .A3(N14), .ZN(n977) );
  AND3_X1 U82 ( .A1(n1133), .A2(n849), .A3(N13), .ZN(n1123) );
  AND3_X1 U83 ( .A1(n1133), .A2(n848), .A3(N14), .ZN(n1050) );
  NOR2_X1 U84 ( .A1(n847), .A2(addr[5]), .ZN(n1133) );
  INV_X1 U85 ( .A(wr_en), .ZN(n847) );
  OAI21_X1 U86 ( .B1(n623), .B2(n1173), .A(n1172), .ZN(n881) );
  NAND2_X1 U87 ( .A1(\mem[4][0] ), .A2(n1173), .ZN(n1172) );
  OAI21_X1 U88 ( .B1(n624), .B2(n1173), .A(n1171), .ZN(n880) );
  NAND2_X1 U89 ( .A1(\mem[4][1] ), .A2(n1173), .ZN(n1171) );
  OAI21_X1 U90 ( .B1(n625), .B2(n1173), .A(n1170), .ZN(n879) );
  NAND2_X1 U91 ( .A1(\mem[4][2] ), .A2(n1173), .ZN(n1170) );
  OAI21_X1 U92 ( .B1(n626), .B2(n1173), .A(n1169), .ZN(n878) );
  NAND2_X1 U93 ( .A1(\mem[4][3] ), .A2(n1173), .ZN(n1169) );
  OAI21_X1 U94 ( .B1(n627), .B2(n1173), .A(n1168), .ZN(n877) );
  NAND2_X1 U95 ( .A1(\mem[4][4] ), .A2(n1173), .ZN(n1168) );
  OAI21_X1 U96 ( .B1(n628), .B2(n1173), .A(n1167), .ZN(n876) );
  NAND2_X1 U97 ( .A1(\mem[4][5] ), .A2(n1173), .ZN(n1167) );
  OAI21_X1 U98 ( .B1(n629), .B2(n1173), .A(n1166), .ZN(n875) );
  NAND2_X1 U99 ( .A1(\mem[4][6] ), .A2(n1173), .ZN(n1166) );
  OAI21_X1 U100 ( .B1(n630), .B2(n1173), .A(n1165), .ZN(n874) );
  NAND2_X1 U101 ( .A1(\mem[4][7] ), .A2(n1173), .ZN(n1165) );
  OAI21_X1 U102 ( .B1(n623), .B2(n1153), .A(n1152), .ZN(n865) );
  NAND2_X1 U103 ( .A1(\mem[6][0] ), .A2(n1153), .ZN(n1152) );
  OAI21_X1 U104 ( .B1(n624), .B2(n1153), .A(n1151), .ZN(n864) );
  NAND2_X1 U105 ( .A1(\mem[6][1] ), .A2(n1153), .ZN(n1151) );
  OAI21_X1 U106 ( .B1(n625), .B2(n1153), .A(n1150), .ZN(n863) );
  NAND2_X1 U107 ( .A1(\mem[6][2] ), .A2(n1153), .ZN(n1150) );
  OAI21_X1 U108 ( .B1(n626), .B2(n1153), .A(n1149), .ZN(n862) );
  NAND2_X1 U109 ( .A1(\mem[6][3] ), .A2(n1153), .ZN(n1149) );
  OAI21_X1 U110 ( .B1(n627), .B2(n1153), .A(n1148), .ZN(n861) );
  NAND2_X1 U111 ( .A1(\mem[6][4] ), .A2(n1153), .ZN(n1148) );
  OAI21_X1 U112 ( .B1(n628), .B2(n1153), .A(n1147), .ZN(n860) );
  NAND2_X1 U113 ( .A1(\mem[6][5] ), .A2(n1153), .ZN(n1147) );
  OAI21_X1 U114 ( .B1(n629), .B2(n1153), .A(n1146), .ZN(n859) );
  NAND2_X1 U115 ( .A1(\mem[6][6] ), .A2(n1153), .ZN(n1146) );
  OAI21_X1 U116 ( .B1(n630), .B2(n1153), .A(n1145), .ZN(n858) );
  NAND2_X1 U117 ( .A1(\mem[6][7] ), .A2(n1153), .ZN(n1145) );
  OAI21_X1 U118 ( .B1(n623), .B2(n1143), .A(n1142), .ZN(n857) );
  NAND2_X1 U119 ( .A1(\mem[7][0] ), .A2(n1143), .ZN(n1142) );
  OAI21_X1 U120 ( .B1(n624), .B2(n1143), .A(n1141), .ZN(n856) );
  NAND2_X1 U121 ( .A1(\mem[7][1] ), .A2(n1143), .ZN(n1141) );
  OAI21_X1 U122 ( .B1(n625), .B2(n1143), .A(n1140), .ZN(n855) );
  NAND2_X1 U123 ( .A1(\mem[7][2] ), .A2(n1143), .ZN(n1140) );
  OAI21_X1 U124 ( .B1(n626), .B2(n1143), .A(n1139), .ZN(n854) );
  NAND2_X1 U125 ( .A1(\mem[7][3] ), .A2(n1143), .ZN(n1139) );
  OAI21_X1 U126 ( .B1(n627), .B2(n1143), .A(n1138), .ZN(n853) );
  NAND2_X1 U127 ( .A1(\mem[7][4] ), .A2(n1143), .ZN(n1138) );
  OAI21_X1 U128 ( .B1(n628), .B2(n1143), .A(n1137), .ZN(n852) );
  NAND2_X1 U129 ( .A1(\mem[7][5] ), .A2(n1143), .ZN(n1137) );
  OAI21_X1 U130 ( .B1(n629), .B2(n1143), .A(n1136), .ZN(n851) );
  NAND2_X1 U131 ( .A1(\mem[7][6] ), .A2(n1143), .ZN(n1136) );
  OAI21_X1 U132 ( .B1(n630), .B2(n1143), .A(n1135), .ZN(n850) );
  NAND2_X1 U133 ( .A1(\mem[7][7] ), .A2(n1143), .ZN(n1135) );
  OAI21_X1 U134 ( .B1(n623), .B2(n1203), .A(n1202), .ZN(n905) );
  NAND2_X1 U135 ( .A1(\mem[1][0] ), .A2(n1203), .ZN(n1202) );
  OAI21_X1 U136 ( .B1(n624), .B2(n1203), .A(n1201), .ZN(n904) );
  NAND2_X1 U137 ( .A1(\mem[1][1] ), .A2(n1203), .ZN(n1201) );
  OAI21_X1 U138 ( .B1(n625), .B2(n1203), .A(n1200), .ZN(n903) );
  NAND2_X1 U139 ( .A1(\mem[1][2] ), .A2(n1203), .ZN(n1200) );
  OAI21_X1 U140 ( .B1(n626), .B2(n1203), .A(n1199), .ZN(n902) );
  NAND2_X1 U141 ( .A1(\mem[1][3] ), .A2(n1203), .ZN(n1199) );
  OAI21_X1 U142 ( .B1(n627), .B2(n1203), .A(n1198), .ZN(n901) );
  NAND2_X1 U143 ( .A1(\mem[1][4] ), .A2(n1203), .ZN(n1198) );
  OAI21_X1 U144 ( .B1(n628), .B2(n1203), .A(n1197), .ZN(n900) );
  NAND2_X1 U145 ( .A1(\mem[1][5] ), .A2(n1203), .ZN(n1197) );
  OAI21_X1 U146 ( .B1(n629), .B2(n1203), .A(n1196), .ZN(n899) );
  NAND2_X1 U147 ( .A1(\mem[1][6] ), .A2(n1203), .ZN(n1196) );
  OAI21_X1 U148 ( .B1(n630), .B2(n1203), .A(n1195), .ZN(n898) );
  NAND2_X1 U149 ( .A1(\mem[1][7] ), .A2(n1203), .ZN(n1195) );
  OAI21_X1 U150 ( .B1(n623), .B2(n1193), .A(n1192), .ZN(n897) );
  NAND2_X1 U151 ( .A1(\mem[2][0] ), .A2(n1193), .ZN(n1192) );
  OAI21_X1 U152 ( .B1(n624), .B2(n1193), .A(n1191), .ZN(n896) );
  NAND2_X1 U153 ( .A1(\mem[2][1] ), .A2(n1193), .ZN(n1191) );
  OAI21_X1 U154 ( .B1(n625), .B2(n1193), .A(n1190), .ZN(n895) );
  NAND2_X1 U155 ( .A1(\mem[2][2] ), .A2(n1193), .ZN(n1190) );
  OAI21_X1 U156 ( .B1(n626), .B2(n1193), .A(n1189), .ZN(n894) );
  NAND2_X1 U157 ( .A1(\mem[2][3] ), .A2(n1193), .ZN(n1189) );
  OAI21_X1 U158 ( .B1(n627), .B2(n1193), .A(n1188), .ZN(n893) );
  NAND2_X1 U159 ( .A1(\mem[2][4] ), .A2(n1193), .ZN(n1188) );
  OAI21_X1 U160 ( .B1(n628), .B2(n1193), .A(n1187), .ZN(n892) );
  NAND2_X1 U161 ( .A1(\mem[2][5] ), .A2(n1193), .ZN(n1187) );
  OAI21_X1 U162 ( .B1(n629), .B2(n1193), .A(n1186), .ZN(n891) );
  NAND2_X1 U163 ( .A1(\mem[2][6] ), .A2(n1193), .ZN(n1186) );
  OAI21_X1 U164 ( .B1(n630), .B2(n1193), .A(n1185), .ZN(n890) );
  NAND2_X1 U165 ( .A1(\mem[2][7] ), .A2(n1193), .ZN(n1185) );
  OAI21_X1 U166 ( .B1(n623), .B2(n1183), .A(n1182), .ZN(n889) );
  NAND2_X1 U167 ( .A1(\mem[3][0] ), .A2(n1183), .ZN(n1182) );
  OAI21_X1 U168 ( .B1(n624), .B2(n1183), .A(n1181), .ZN(n888) );
  NAND2_X1 U169 ( .A1(\mem[3][1] ), .A2(n1183), .ZN(n1181) );
  OAI21_X1 U170 ( .B1(n625), .B2(n1183), .A(n1180), .ZN(n887) );
  NAND2_X1 U171 ( .A1(\mem[3][2] ), .A2(n1183), .ZN(n1180) );
  OAI21_X1 U172 ( .B1(n626), .B2(n1183), .A(n1179), .ZN(n886) );
  NAND2_X1 U173 ( .A1(\mem[3][3] ), .A2(n1183), .ZN(n1179) );
  OAI21_X1 U174 ( .B1(n627), .B2(n1183), .A(n1178), .ZN(n885) );
  NAND2_X1 U175 ( .A1(\mem[3][4] ), .A2(n1183), .ZN(n1178) );
  OAI21_X1 U176 ( .B1(n628), .B2(n1183), .A(n1177), .ZN(n884) );
  NAND2_X1 U177 ( .A1(\mem[3][5] ), .A2(n1183), .ZN(n1177) );
  OAI21_X1 U178 ( .B1(n629), .B2(n1183), .A(n1176), .ZN(n883) );
  NAND2_X1 U179 ( .A1(\mem[3][6] ), .A2(n1183), .ZN(n1176) );
  OAI21_X1 U180 ( .B1(n630), .B2(n1183), .A(n1175), .ZN(n882) );
  NAND2_X1 U181 ( .A1(\mem[3][7] ), .A2(n1183), .ZN(n1175) );
  OAI21_X1 U182 ( .B1(n623), .B2(n1163), .A(n1162), .ZN(n873) );
  NAND2_X1 U183 ( .A1(\mem[5][0] ), .A2(n1163), .ZN(n1162) );
  OAI21_X1 U184 ( .B1(n624), .B2(n1163), .A(n1161), .ZN(n872) );
  NAND2_X1 U185 ( .A1(\mem[5][1] ), .A2(n1163), .ZN(n1161) );
  OAI21_X1 U186 ( .B1(n625), .B2(n1163), .A(n1160), .ZN(n871) );
  NAND2_X1 U187 ( .A1(\mem[5][2] ), .A2(n1163), .ZN(n1160) );
  OAI21_X1 U188 ( .B1(n626), .B2(n1163), .A(n1159), .ZN(n870) );
  NAND2_X1 U189 ( .A1(\mem[5][3] ), .A2(n1163), .ZN(n1159) );
  OAI21_X1 U190 ( .B1(n627), .B2(n1163), .A(n1158), .ZN(n869) );
  NAND2_X1 U191 ( .A1(\mem[5][4] ), .A2(n1163), .ZN(n1158) );
  OAI21_X1 U192 ( .B1(n628), .B2(n1163), .A(n1157), .ZN(n868) );
  NAND2_X1 U193 ( .A1(\mem[5][5] ), .A2(n1163), .ZN(n1157) );
  OAI21_X1 U194 ( .B1(n629), .B2(n1163), .A(n1156), .ZN(n867) );
  NAND2_X1 U195 ( .A1(\mem[5][6] ), .A2(n1163), .ZN(n1156) );
  OAI21_X1 U196 ( .B1(n630), .B2(n1163), .A(n1155), .ZN(n866) );
  NAND2_X1 U197 ( .A1(\mem[5][7] ), .A2(n1163), .ZN(n1155) );
  OAI21_X1 U198 ( .B1(n1214), .B2(n623), .A(n1213), .ZN(n913) );
  NAND2_X1 U199 ( .A1(\mem[0][0] ), .A2(n1214), .ZN(n1213) );
  OAI21_X1 U200 ( .B1(n1214), .B2(n624), .A(n1212), .ZN(n912) );
  NAND2_X1 U201 ( .A1(\mem[0][1] ), .A2(n1214), .ZN(n1212) );
  OAI21_X1 U202 ( .B1(n1214), .B2(n625), .A(n1211), .ZN(n911) );
  NAND2_X1 U203 ( .A1(\mem[0][2] ), .A2(n1214), .ZN(n1211) );
  OAI21_X1 U204 ( .B1(n1214), .B2(n626), .A(n1210), .ZN(n910) );
  NAND2_X1 U205 ( .A1(\mem[0][3] ), .A2(n1214), .ZN(n1210) );
  OAI21_X1 U206 ( .B1(n1214), .B2(n627), .A(n1209), .ZN(n909) );
  NAND2_X1 U207 ( .A1(\mem[0][4] ), .A2(n1214), .ZN(n1209) );
  OAI21_X1 U208 ( .B1(n1214), .B2(n628), .A(n1208), .ZN(n908) );
  NAND2_X1 U209 ( .A1(\mem[0][5] ), .A2(n1214), .ZN(n1208) );
  OAI21_X1 U210 ( .B1(n1214), .B2(n629), .A(n1207), .ZN(n907) );
  NAND2_X1 U211 ( .A1(\mem[0][6] ), .A2(n1214), .ZN(n1207) );
  OAI21_X1 U212 ( .B1(n1214), .B2(n630), .A(n1206), .ZN(n906) );
  NAND2_X1 U213 ( .A1(\mem[0][7] ), .A2(n1214), .ZN(n1206) );
  INV_X1 U214 ( .A(n1132), .ZN(n822) );
  AOI22_X1 U215 ( .A1(data_in[0]), .A2(n846), .B1(n1131), .B2(\mem[8][0] ), 
        .ZN(n1132) );
  INV_X1 U216 ( .A(n1130), .ZN(n821) );
  AOI22_X1 U217 ( .A1(data_in[1]), .A2(n846), .B1(n1131), .B2(\mem[8][1] ), 
        .ZN(n1130) );
  INV_X1 U218 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U219 ( .A1(data_in[2]), .A2(n846), .B1(n1131), .B2(\mem[8][2] ), 
        .ZN(n1129) );
  INV_X1 U220 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U221 ( .A1(data_in[3]), .A2(n846), .B1(n1131), .B2(\mem[8][3] ), 
        .ZN(n1128) );
  INV_X1 U222 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U223 ( .A1(data_in[4]), .A2(n846), .B1(n1131), .B2(\mem[8][4] ), 
        .ZN(n1127) );
  INV_X1 U224 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U225 ( .A1(data_in[5]), .A2(n846), .B1(n1131), .B2(\mem[8][5] ), 
        .ZN(n1126) );
  INV_X1 U226 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U227 ( .A1(data_in[6]), .A2(n846), .B1(n1131), .B2(\mem[8][6] ), 
        .ZN(n1125) );
  INV_X1 U228 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U229 ( .A1(data_in[7]), .A2(n846), .B1(n1131), .B2(\mem[8][7] ), 
        .ZN(n1124) );
  INV_X1 U230 ( .A(n1122), .ZN(n814) );
  AOI22_X1 U231 ( .A1(data_in[0]), .A2(n845), .B1(n1121), .B2(\mem[9][0] ), 
        .ZN(n1122) );
  INV_X1 U232 ( .A(n1120), .ZN(n813) );
  AOI22_X1 U233 ( .A1(data_in[1]), .A2(n845), .B1(n1121), .B2(\mem[9][1] ), 
        .ZN(n1120) );
  INV_X1 U234 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U235 ( .A1(data_in[2]), .A2(n845), .B1(n1121), .B2(\mem[9][2] ), 
        .ZN(n1119) );
  INV_X1 U236 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U237 ( .A1(data_in[3]), .A2(n845), .B1(n1121), .B2(\mem[9][3] ), 
        .ZN(n1118) );
  INV_X1 U238 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U239 ( .A1(data_in[4]), .A2(n845), .B1(n1121), .B2(\mem[9][4] ), 
        .ZN(n1117) );
  INV_X1 U240 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U241 ( .A1(data_in[5]), .A2(n845), .B1(n1121), .B2(\mem[9][5] ), 
        .ZN(n1116) );
  INV_X1 U242 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U243 ( .A1(data_in[6]), .A2(n845), .B1(n1121), .B2(\mem[9][6] ), 
        .ZN(n1115) );
  INV_X1 U244 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U245 ( .A1(data_in[7]), .A2(n845), .B1(n1121), .B2(\mem[9][7] ), 
        .ZN(n1114) );
  INV_X1 U246 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U247 ( .A1(data_in[0]), .A2(n844), .B1(n1112), .B2(\mem[10][0] ), 
        .ZN(n1113) );
  INV_X1 U248 ( .A(n1111), .ZN(n805) );
  AOI22_X1 U249 ( .A1(data_in[1]), .A2(n844), .B1(n1112), .B2(\mem[10][1] ), 
        .ZN(n1111) );
  INV_X1 U250 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U251 ( .A1(data_in[2]), .A2(n844), .B1(n1112), .B2(\mem[10][2] ), 
        .ZN(n1110) );
  INV_X1 U252 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U253 ( .A1(data_in[3]), .A2(n844), .B1(n1112), .B2(\mem[10][3] ), 
        .ZN(n1109) );
  INV_X1 U254 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U255 ( .A1(data_in[4]), .A2(n844), .B1(n1112), .B2(\mem[10][4] ), 
        .ZN(n1108) );
  INV_X1 U256 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U257 ( .A1(data_in[5]), .A2(n844), .B1(n1112), .B2(\mem[10][5] ), 
        .ZN(n1107) );
  INV_X1 U258 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U259 ( .A1(data_in[6]), .A2(n844), .B1(n1112), .B2(\mem[10][6] ), 
        .ZN(n1106) );
  INV_X1 U260 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U261 ( .A1(data_in[7]), .A2(n844), .B1(n1112), .B2(\mem[10][7] ), 
        .ZN(n1105) );
  INV_X1 U262 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U263 ( .A1(data_in[0]), .A2(n843), .B1(n1103), .B2(\mem[11][0] ), 
        .ZN(n1104) );
  INV_X1 U264 ( .A(n1102), .ZN(n797) );
  AOI22_X1 U265 ( .A1(data_in[1]), .A2(n843), .B1(n1103), .B2(\mem[11][1] ), 
        .ZN(n1102) );
  INV_X1 U266 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U267 ( .A1(data_in[2]), .A2(n843), .B1(n1103), .B2(\mem[11][2] ), 
        .ZN(n1101) );
  INV_X1 U268 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U269 ( .A1(data_in[3]), .A2(n843), .B1(n1103), .B2(\mem[11][3] ), 
        .ZN(n1100) );
  INV_X1 U270 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U271 ( .A1(data_in[4]), .A2(n843), .B1(n1103), .B2(\mem[11][4] ), 
        .ZN(n1099) );
  INV_X1 U272 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U273 ( .A1(data_in[5]), .A2(n843), .B1(n1103), .B2(\mem[11][5] ), 
        .ZN(n1098) );
  INV_X1 U274 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U275 ( .A1(data_in[6]), .A2(n843), .B1(n1103), .B2(\mem[11][6] ), 
        .ZN(n1097) );
  INV_X1 U276 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U277 ( .A1(data_in[7]), .A2(n843), .B1(n1103), .B2(\mem[11][7] ), 
        .ZN(n1096) );
  INV_X1 U278 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U279 ( .A1(data_in[0]), .A2(n842), .B1(n1094), .B2(\mem[12][0] ), 
        .ZN(n1095) );
  INV_X1 U280 ( .A(n1093), .ZN(n789) );
  AOI22_X1 U281 ( .A1(data_in[1]), .A2(n842), .B1(n1094), .B2(\mem[12][1] ), 
        .ZN(n1093) );
  INV_X1 U282 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U283 ( .A1(data_in[2]), .A2(n842), .B1(n1094), .B2(\mem[12][2] ), 
        .ZN(n1092) );
  INV_X1 U284 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U285 ( .A1(data_in[3]), .A2(n842), .B1(n1094), .B2(\mem[12][3] ), 
        .ZN(n1091) );
  INV_X1 U286 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U287 ( .A1(data_in[4]), .A2(n842), .B1(n1094), .B2(\mem[12][4] ), 
        .ZN(n1090) );
  INV_X1 U288 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U289 ( .A1(data_in[5]), .A2(n842), .B1(n1094), .B2(\mem[12][5] ), 
        .ZN(n1089) );
  INV_X1 U290 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U291 ( .A1(data_in[6]), .A2(n842), .B1(n1094), .B2(\mem[12][6] ), 
        .ZN(n1088) );
  INV_X1 U292 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U293 ( .A1(data_in[7]), .A2(n842), .B1(n1094), .B2(\mem[12][7] ), 
        .ZN(n1087) );
  INV_X1 U294 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U295 ( .A1(data_in[0]), .A2(n841), .B1(n1085), .B2(\mem[13][0] ), 
        .ZN(n1086) );
  INV_X1 U296 ( .A(n1084), .ZN(n781) );
  AOI22_X1 U297 ( .A1(data_in[1]), .A2(n841), .B1(n1085), .B2(\mem[13][1] ), 
        .ZN(n1084) );
  INV_X1 U298 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U299 ( .A1(data_in[2]), .A2(n841), .B1(n1085), .B2(\mem[13][2] ), 
        .ZN(n1083) );
  INV_X1 U300 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U301 ( .A1(data_in[3]), .A2(n841), .B1(n1085), .B2(\mem[13][3] ), 
        .ZN(n1082) );
  INV_X1 U302 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U303 ( .A1(data_in[4]), .A2(n841), .B1(n1085), .B2(\mem[13][4] ), 
        .ZN(n1081) );
  INV_X1 U304 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U305 ( .A1(data_in[5]), .A2(n841), .B1(n1085), .B2(\mem[13][5] ), 
        .ZN(n1080) );
  INV_X1 U306 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U307 ( .A1(data_in[6]), .A2(n841), .B1(n1085), .B2(\mem[13][6] ), 
        .ZN(n1079) );
  INV_X1 U308 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U309 ( .A1(data_in[7]), .A2(n841), .B1(n1085), .B2(\mem[13][7] ), 
        .ZN(n1078) );
  INV_X1 U310 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U311 ( .A1(data_in[0]), .A2(n840), .B1(n1076), .B2(\mem[14][0] ), 
        .ZN(n1077) );
  INV_X1 U312 ( .A(n1075), .ZN(n773) );
  AOI22_X1 U313 ( .A1(data_in[1]), .A2(n840), .B1(n1076), .B2(\mem[14][1] ), 
        .ZN(n1075) );
  INV_X1 U314 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U315 ( .A1(data_in[2]), .A2(n840), .B1(n1076), .B2(\mem[14][2] ), 
        .ZN(n1074) );
  INV_X1 U316 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U317 ( .A1(data_in[3]), .A2(n840), .B1(n1076), .B2(\mem[14][3] ), 
        .ZN(n1073) );
  INV_X1 U318 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U319 ( .A1(data_in[4]), .A2(n840), .B1(n1076), .B2(\mem[14][4] ), 
        .ZN(n1072) );
  INV_X1 U320 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U321 ( .A1(data_in[5]), .A2(n840), .B1(n1076), .B2(\mem[14][5] ), 
        .ZN(n1071) );
  INV_X1 U322 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U323 ( .A1(data_in[6]), .A2(n840), .B1(n1076), .B2(\mem[14][6] ), 
        .ZN(n1070) );
  INV_X1 U324 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U325 ( .A1(data_in[7]), .A2(n840), .B1(n1076), .B2(\mem[14][7] ), 
        .ZN(n1069) );
  INV_X1 U326 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U327 ( .A1(data_in[0]), .A2(n839), .B1(n1067), .B2(\mem[15][0] ), 
        .ZN(n1068) );
  INV_X1 U328 ( .A(n1066), .ZN(n765) );
  AOI22_X1 U329 ( .A1(data_in[1]), .A2(n839), .B1(n1067), .B2(\mem[15][1] ), 
        .ZN(n1066) );
  INV_X1 U330 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U331 ( .A1(data_in[2]), .A2(n839), .B1(n1067), .B2(\mem[15][2] ), 
        .ZN(n1065) );
  INV_X1 U332 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U333 ( .A1(data_in[3]), .A2(n839), .B1(n1067), .B2(\mem[15][3] ), 
        .ZN(n1064) );
  INV_X1 U334 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U335 ( .A1(data_in[4]), .A2(n839), .B1(n1067), .B2(\mem[15][4] ), 
        .ZN(n1063) );
  INV_X1 U336 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U337 ( .A1(data_in[5]), .A2(n839), .B1(n1067), .B2(\mem[15][5] ), 
        .ZN(n1062) );
  INV_X1 U338 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U339 ( .A1(data_in[6]), .A2(n839), .B1(n1067), .B2(\mem[15][6] ), 
        .ZN(n1061) );
  INV_X1 U340 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U341 ( .A1(data_in[7]), .A2(n839), .B1(n1067), .B2(\mem[15][7] ), 
        .ZN(n1060) );
  INV_X1 U342 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U343 ( .A1(data_in[0]), .A2(n838), .B1(n1058), .B2(\mem[16][0] ), 
        .ZN(n1059) );
  INV_X1 U344 ( .A(n1057), .ZN(n757) );
  AOI22_X1 U345 ( .A1(data_in[1]), .A2(n838), .B1(n1058), .B2(\mem[16][1] ), 
        .ZN(n1057) );
  INV_X1 U346 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U347 ( .A1(data_in[2]), .A2(n838), .B1(n1058), .B2(\mem[16][2] ), 
        .ZN(n1056) );
  INV_X1 U348 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U349 ( .A1(data_in[3]), .A2(n838), .B1(n1058), .B2(\mem[16][3] ), 
        .ZN(n1055) );
  INV_X1 U350 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U351 ( .A1(data_in[4]), .A2(n838), .B1(n1058), .B2(\mem[16][4] ), 
        .ZN(n1054) );
  INV_X1 U352 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U353 ( .A1(data_in[5]), .A2(n838), .B1(n1058), .B2(\mem[16][5] ), 
        .ZN(n1053) );
  INV_X1 U354 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U355 ( .A1(data_in[6]), .A2(n838), .B1(n1058), .B2(\mem[16][6] ), 
        .ZN(n1052) );
  INV_X1 U356 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U357 ( .A1(data_in[7]), .A2(n838), .B1(n1058), .B2(\mem[16][7] ), 
        .ZN(n1051) );
  INV_X1 U358 ( .A(n1049), .ZN(n750) );
  AOI22_X1 U359 ( .A1(data_in[0]), .A2(n837), .B1(n1048), .B2(\mem[17][0] ), 
        .ZN(n1049) );
  INV_X1 U360 ( .A(n1047), .ZN(n749) );
  AOI22_X1 U361 ( .A1(data_in[1]), .A2(n837), .B1(n1048), .B2(\mem[17][1] ), 
        .ZN(n1047) );
  INV_X1 U362 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U363 ( .A1(data_in[2]), .A2(n837), .B1(n1048), .B2(\mem[17][2] ), 
        .ZN(n1046) );
  INV_X1 U364 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U365 ( .A1(data_in[3]), .A2(n837), .B1(n1048), .B2(\mem[17][3] ), 
        .ZN(n1045) );
  INV_X1 U366 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U367 ( .A1(data_in[4]), .A2(n837), .B1(n1048), .B2(\mem[17][4] ), 
        .ZN(n1044) );
  INV_X1 U368 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U369 ( .A1(data_in[5]), .A2(n837), .B1(n1048), .B2(\mem[17][5] ), 
        .ZN(n1043) );
  INV_X1 U370 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U371 ( .A1(data_in[6]), .A2(n837), .B1(n1048), .B2(\mem[17][6] ), 
        .ZN(n1042) );
  INV_X1 U372 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U373 ( .A1(data_in[7]), .A2(n837), .B1(n1048), .B2(\mem[17][7] ), 
        .ZN(n1041) );
  INV_X1 U374 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U375 ( .A1(data_in[0]), .A2(n836), .B1(n1039), .B2(\mem[18][0] ), 
        .ZN(n1040) );
  INV_X1 U376 ( .A(n1038), .ZN(n741) );
  AOI22_X1 U377 ( .A1(data_in[1]), .A2(n836), .B1(n1039), .B2(\mem[18][1] ), 
        .ZN(n1038) );
  INV_X1 U378 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U379 ( .A1(data_in[2]), .A2(n836), .B1(n1039), .B2(\mem[18][2] ), 
        .ZN(n1037) );
  INV_X1 U380 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U381 ( .A1(data_in[3]), .A2(n836), .B1(n1039), .B2(\mem[18][3] ), 
        .ZN(n1036) );
  INV_X1 U382 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U383 ( .A1(data_in[4]), .A2(n836), .B1(n1039), .B2(\mem[18][4] ), 
        .ZN(n1035) );
  INV_X1 U384 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U385 ( .A1(data_in[5]), .A2(n836), .B1(n1039), .B2(\mem[18][5] ), 
        .ZN(n1034) );
  INV_X1 U386 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U387 ( .A1(data_in[6]), .A2(n836), .B1(n1039), .B2(\mem[18][6] ), 
        .ZN(n1033) );
  INV_X1 U388 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U389 ( .A1(data_in[7]), .A2(n836), .B1(n1039), .B2(\mem[18][7] ), 
        .ZN(n1032) );
  INV_X1 U390 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U391 ( .A1(data_in[0]), .A2(n835), .B1(n1030), .B2(\mem[19][0] ), 
        .ZN(n1031) );
  INV_X1 U392 ( .A(n1029), .ZN(n733) );
  AOI22_X1 U393 ( .A1(data_in[1]), .A2(n835), .B1(n1030), .B2(\mem[19][1] ), 
        .ZN(n1029) );
  INV_X1 U394 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U395 ( .A1(data_in[2]), .A2(n835), .B1(n1030), .B2(\mem[19][2] ), 
        .ZN(n1028) );
  INV_X1 U396 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U397 ( .A1(data_in[3]), .A2(n835), .B1(n1030), .B2(\mem[19][3] ), 
        .ZN(n1027) );
  INV_X1 U398 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U399 ( .A1(data_in[4]), .A2(n835), .B1(n1030), .B2(\mem[19][4] ), 
        .ZN(n1026) );
  INV_X1 U400 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U401 ( .A1(data_in[5]), .A2(n835), .B1(n1030), .B2(\mem[19][5] ), 
        .ZN(n1025) );
  INV_X1 U402 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U403 ( .A1(data_in[6]), .A2(n835), .B1(n1030), .B2(\mem[19][6] ), 
        .ZN(n1024) );
  INV_X1 U404 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U405 ( .A1(data_in[7]), .A2(n835), .B1(n1030), .B2(\mem[19][7] ), 
        .ZN(n1023) );
  INV_X1 U406 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U407 ( .A1(data_in[0]), .A2(n834), .B1(n1021), .B2(\mem[20][0] ), 
        .ZN(n1022) );
  INV_X1 U408 ( .A(n1020), .ZN(n725) );
  AOI22_X1 U409 ( .A1(data_in[1]), .A2(n834), .B1(n1021), .B2(\mem[20][1] ), 
        .ZN(n1020) );
  INV_X1 U410 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U411 ( .A1(data_in[2]), .A2(n834), .B1(n1021), .B2(\mem[20][2] ), 
        .ZN(n1019) );
  INV_X1 U412 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U413 ( .A1(data_in[3]), .A2(n834), .B1(n1021), .B2(\mem[20][3] ), 
        .ZN(n1018) );
  INV_X1 U414 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U415 ( .A1(data_in[4]), .A2(n834), .B1(n1021), .B2(\mem[20][4] ), 
        .ZN(n1017) );
  INV_X1 U416 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U417 ( .A1(data_in[5]), .A2(n834), .B1(n1021), .B2(\mem[20][5] ), 
        .ZN(n1016) );
  INV_X1 U418 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U419 ( .A1(data_in[6]), .A2(n834), .B1(n1021), .B2(\mem[20][6] ), 
        .ZN(n1015) );
  INV_X1 U420 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U421 ( .A1(data_in[7]), .A2(n834), .B1(n1021), .B2(\mem[20][7] ), 
        .ZN(n1014) );
  INV_X1 U422 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U423 ( .A1(data_in[0]), .A2(n833), .B1(n1012), .B2(\mem[21][0] ), 
        .ZN(n1013) );
  INV_X1 U424 ( .A(n1011), .ZN(n717) );
  AOI22_X1 U425 ( .A1(data_in[1]), .A2(n833), .B1(n1012), .B2(\mem[21][1] ), 
        .ZN(n1011) );
  INV_X1 U426 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U427 ( .A1(data_in[2]), .A2(n833), .B1(n1012), .B2(\mem[21][2] ), 
        .ZN(n1010) );
  INV_X1 U428 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U429 ( .A1(data_in[3]), .A2(n833), .B1(n1012), .B2(\mem[21][3] ), 
        .ZN(n1009) );
  INV_X1 U430 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U431 ( .A1(data_in[4]), .A2(n833), .B1(n1012), .B2(\mem[21][4] ), 
        .ZN(n1008) );
  INV_X1 U432 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U433 ( .A1(data_in[5]), .A2(n833), .B1(n1012), .B2(\mem[21][5] ), 
        .ZN(n1007) );
  INV_X1 U434 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U435 ( .A1(data_in[6]), .A2(n833), .B1(n1012), .B2(\mem[21][6] ), 
        .ZN(n1006) );
  INV_X1 U436 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U437 ( .A1(data_in[7]), .A2(n833), .B1(n1012), .B2(\mem[21][7] ), 
        .ZN(n1005) );
  INV_X1 U438 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U439 ( .A1(data_in[0]), .A2(n832), .B1(n1003), .B2(\mem[22][0] ), 
        .ZN(n1004) );
  INV_X1 U440 ( .A(n1002), .ZN(n709) );
  AOI22_X1 U441 ( .A1(data_in[1]), .A2(n832), .B1(n1003), .B2(\mem[22][1] ), 
        .ZN(n1002) );
  INV_X1 U442 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U443 ( .A1(data_in[2]), .A2(n832), .B1(n1003), .B2(\mem[22][2] ), 
        .ZN(n1001) );
  INV_X1 U444 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U445 ( .A1(data_in[3]), .A2(n832), .B1(n1003), .B2(\mem[22][3] ), 
        .ZN(n1000) );
  INV_X1 U446 ( .A(n999), .ZN(n706) );
  AOI22_X1 U447 ( .A1(data_in[4]), .A2(n832), .B1(n1003), .B2(\mem[22][4] ), 
        .ZN(n999) );
  INV_X1 U448 ( .A(n998), .ZN(n705) );
  AOI22_X1 U449 ( .A1(data_in[5]), .A2(n832), .B1(n1003), .B2(\mem[22][5] ), 
        .ZN(n998) );
  INV_X1 U450 ( .A(n997), .ZN(n704) );
  AOI22_X1 U451 ( .A1(data_in[6]), .A2(n832), .B1(n1003), .B2(\mem[22][6] ), 
        .ZN(n997) );
  INV_X1 U452 ( .A(n996), .ZN(n703) );
  AOI22_X1 U453 ( .A1(data_in[7]), .A2(n832), .B1(n1003), .B2(\mem[22][7] ), 
        .ZN(n996) );
  INV_X1 U454 ( .A(n995), .ZN(n702) );
  AOI22_X1 U455 ( .A1(data_in[0]), .A2(n831), .B1(n994), .B2(\mem[23][0] ), 
        .ZN(n995) );
  INV_X1 U456 ( .A(n993), .ZN(n701) );
  AOI22_X1 U457 ( .A1(data_in[1]), .A2(n831), .B1(n994), .B2(\mem[23][1] ), 
        .ZN(n993) );
  INV_X1 U458 ( .A(n992), .ZN(n700) );
  AOI22_X1 U459 ( .A1(data_in[2]), .A2(n831), .B1(n994), .B2(\mem[23][2] ), 
        .ZN(n992) );
  INV_X1 U460 ( .A(n991), .ZN(n699) );
  AOI22_X1 U461 ( .A1(data_in[3]), .A2(n831), .B1(n994), .B2(\mem[23][3] ), 
        .ZN(n991) );
  INV_X1 U462 ( .A(n990), .ZN(n698) );
  AOI22_X1 U463 ( .A1(data_in[4]), .A2(n831), .B1(n994), .B2(\mem[23][4] ), 
        .ZN(n990) );
  INV_X1 U464 ( .A(n989), .ZN(n697) );
  AOI22_X1 U465 ( .A1(data_in[5]), .A2(n831), .B1(n994), .B2(\mem[23][5] ), 
        .ZN(n989) );
  INV_X1 U466 ( .A(n988), .ZN(n696) );
  AOI22_X1 U467 ( .A1(data_in[6]), .A2(n831), .B1(n994), .B2(\mem[23][6] ), 
        .ZN(n988) );
  INV_X1 U468 ( .A(n987), .ZN(n695) );
  AOI22_X1 U469 ( .A1(data_in[7]), .A2(n831), .B1(n994), .B2(\mem[23][7] ), 
        .ZN(n987) );
  INV_X1 U470 ( .A(n986), .ZN(n694) );
  AOI22_X1 U471 ( .A1(data_in[0]), .A2(n830), .B1(n985), .B2(\mem[24][0] ), 
        .ZN(n986) );
  INV_X1 U472 ( .A(n984), .ZN(n693) );
  AOI22_X1 U473 ( .A1(data_in[1]), .A2(n830), .B1(n985), .B2(\mem[24][1] ), 
        .ZN(n984) );
  INV_X1 U474 ( .A(n983), .ZN(n692) );
  AOI22_X1 U475 ( .A1(data_in[2]), .A2(n830), .B1(n985), .B2(\mem[24][2] ), 
        .ZN(n983) );
  INV_X1 U476 ( .A(n982), .ZN(n691) );
  AOI22_X1 U477 ( .A1(data_in[3]), .A2(n830), .B1(n985), .B2(\mem[24][3] ), 
        .ZN(n982) );
  INV_X1 U478 ( .A(n981), .ZN(n690) );
  AOI22_X1 U479 ( .A1(data_in[4]), .A2(n830), .B1(n985), .B2(\mem[24][4] ), 
        .ZN(n981) );
  INV_X1 U480 ( .A(n980), .ZN(n689) );
  AOI22_X1 U481 ( .A1(data_in[5]), .A2(n830), .B1(n985), .B2(\mem[24][5] ), 
        .ZN(n980) );
  INV_X1 U482 ( .A(n979), .ZN(n688) );
  AOI22_X1 U483 ( .A1(data_in[6]), .A2(n830), .B1(n985), .B2(\mem[24][6] ), 
        .ZN(n979) );
  INV_X1 U484 ( .A(n978), .ZN(n687) );
  AOI22_X1 U485 ( .A1(data_in[7]), .A2(n830), .B1(n985), .B2(\mem[24][7] ), 
        .ZN(n978) );
  INV_X1 U486 ( .A(n976), .ZN(n686) );
  AOI22_X1 U487 ( .A1(data_in[0]), .A2(n829), .B1(n975), .B2(\mem[25][0] ), 
        .ZN(n976) );
  INV_X1 U488 ( .A(n974), .ZN(n685) );
  AOI22_X1 U489 ( .A1(data_in[1]), .A2(n829), .B1(n975), .B2(\mem[25][1] ), 
        .ZN(n974) );
  INV_X1 U490 ( .A(n973), .ZN(n684) );
  AOI22_X1 U491 ( .A1(data_in[2]), .A2(n829), .B1(n975), .B2(\mem[25][2] ), 
        .ZN(n973) );
  INV_X1 U492 ( .A(n972), .ZN(n683) );
  AOI22_X1 U493 ( .A1(data_in[3]), .A2(n829), .B1(n975), .B2(\mem[25][3] ), 
        .ZN(n972) );
  INV_X1 U494 ( .A(n971), .ZN(n682) );
  AOI22_X1 U495 ( .A1(data_in[4]), .A2(n829), .B1(n975), .B2(\mem[25][4] ), 
        .ZN(n971) );
  INV_X1 U496 ( .A(n970), .ZN(n681) );
  AOI22_X1 U497 ( .A1(data_in[5]), .A2(n829), .B1(n975), .B2(\mem[25][5] ), 
        .ZN(n970) );
  INV_X1 U498 ( .A(n969), .ZN(n680) );
  AOI22_X1 U499 ( .A1(data_in[6]), .A2(n829), .B1(n975), .B2(\mem[25][6] ), 
        .ZN(n969) );
  INV_X1 U500 ( .A(n968), .ZN(n679) );
  AOI22_X1 U501 ( .A1(data_in[7]), .A2(n829), .B1(n975), .B2(\mem[25][7] ), 
        .ZN(n968) );
  INV_X1 U502 ( .A(n967), .ZN(n678) );
  AOI22_X1 U503 ( .A1(data_in[0]), .A2(n828), .B1(n966), .B2(\mem[26][0] ), 
        .ZN(n967) );
  INV_X1 U504 ( .A(n965), .ZN(n677) );
  AOI22_X1 U505 ( .A1(data_in[1]), .A2(n828), .B1(n966), .B2(\mem[26][1] ), 
        .ZN(n965) );
  INV_X1 U506 ( .A(n964), .ZN(n676) );
  AOI22_X1 U507 ( .A1(data_in[2]), .A2(n828), .B1(n966), .B2(\mem[26][2] ), 
        .ZN(n964) );
  INV_X1 U508 ( .A(n963), .ZN(n675) );
  AOI22_X1 U509 ( .A1(data_in[3]), .A2(n828), .B1(n966), .B2(\mem[26][3] ), 
        .ZN(n963) );
  INV_X1 U510 ( .A(n962), .ZN(n674) );
  AOI22_X1 U511 ( .A1(data_in[4]), .A2(n828), .B1(n966), .B2(\mem[26][4] ), 
        .ZN(n962) );
  INV_X1 U512 ( .A(n961), .ZN(n673) );
  AOI22_X1 U513 ( .A1(data_in[5]), .A2(n828), .B1(n966), .B2(\mem[26][5] ), 
        .ZN(n961) );
  INV_X1 U514 ( .A(n960), .ZN(n672) );
  AOI22_X1 U515 ( .A1(data_in[6]), .A2(n828), .B1(n966), .B2(\mem[26][6] ), 
        .ZN(n960) );
  INV_X1 U516 ( .A(n959), .ZN(n671) );
  AOI22_X1 U517 ( .A1(data_in[7]), .A2(n828), .B1(n966), .B2(\mem[26][7] ), 
        .ZN(n959) );
  INV_X1 U518 ( .A(n958), .ZN(n670) );
  AOI22_X1 U519 ( .A1(data_in[0]), .A2(n827), .B1(n957), .B2(\mem[27][0] ), 
        .ZN(n958) );
  INV_X1 U520 ( .A(n956), .ZN(n669) );
  AOI22_X1 U521 ( .A1(data_in[1]), .A2(n827), .B1(n957), .B2(\mem[27][1] ), 
        .ZN(n956) );
  INV_X1 U522 ( .A(n955), .ZN(n668) );
  AOI22_X1 U523 ( .A1(data_in[2]), .A2(n827), .B1(n957), .B2(\mem[27][2] ), 
        .ZN(n955) );
  INV_X1 U524 ( .A(n954), .ZN(n667) );
  AOI22_X1 U525 ( .A1(data_in[3]), .A2(n827), .B1(n957), .B2(\mem[27][3] ), 
        .ZN(n954) );
  INV_X1 U526 ( .A(n953), .ZN(n666) );
  AOI22_X1 U527 ( .A1(data_in[4]), .A2(n827), .B1(n957), .B2(\mem[27][4] ), 
        .ZN(n953) );
  INV_X1 U528 ( .A(n952), .ZN(n665) );
  AOI22_X1 U529 ( .A1(data_in[5]), .A2(n827), .B1(n957), .B2(\mem[27][5] ), 
        .ZN(n952) );
  INV_X1 U530 ( .A(n951), .ZN(n664) );
  AOI22_X1 U531 ( .A1(data_in[6]), .A2(n827), .B1(n957), .B2(\mem[27][6] ), 
        .ZN(n951) );
  INV_X1 U532 ( .A(n950), .ZN(n663) );
  AOI22_X1 U533 ( .A1(data_in[7]), .A2(n827), .B1(n957), .B2(\mem[27][7] ), 
        .ZN(n950) );
  INV_X1 U534 ( .A(n949), .ZN(n662) );
  AOI22_X1 U535 ( .A1(data_in[0]), .A2(n826), .B1(n948), .B2(\mem[28][0] ), 
        .ZN(n949) );
  INV_X1 U536 ( .A(n947), .ZN(n661) );
  AOI22_X1 U537 ( .A1(data_in[1]), .A2(n826), .B1(n948), .B2(\mem[28][1] ), 
        .ZN(n947) );
  INV_X1 U538 ( .A(n946), .ZN(n660) );
  AOI22_X1 U539 ( .A1(data_in[2]), .A2(n826), .B1(n948), .B2(\mem[28][2] ), 
        .ZN(n946) );
  INV_X1 U540 ( .A(n945), .ZN(n659) );
  AOI22_X1 U541 ( .A1(data_in[3]), .A2(n826), .B1(n948), .B2(\mem[28][3] ), 
        .ZN(n945) );
  INV_X1 U542 ( .A(n944), .ZN(n658) );
  AOI22_X1 U543 ( .A1(data_in[4]), .A2(n826), .B1(n948), .B2(\mem[28][4] ), 
        .ZN(n944) );
  INV_X1 U544 ( .A(n943), .ZN(n657) );
  AOI22_X1 U545 ( .A1(data_in[5]), .A2(n826), .B1(n948), .B2(\mem[28][5] ), 
        .ZN(n943) );
  INV_X1 U546 ( .A(n942), .ZN(n656) );
  AOI22_X1 U547 ( .A1(data_in[6]), .A2(n826), .B1(n948), .B2(\mem[28][6] ), 
        .ZN(n942) );
  INV_X1 U548 ( .A(n941), .ZN(n655) );
  AOI22_X1 U549 ( .A1(data_in[7]), .A2(n826), .B1(n948), .B2(\mem[28][7] ), 
        .ZN(n941) );
  INV_X1 U550 ( .A(n940), .ZN(n654) );
  AOI22_X1 U551 ( .A1(data_in[0]), .A2(n825), .B1(n939), .B2(\mem[29][0] ), 
        .ZN(n940) );
  INV_X1 U552 ( .A(n938), .ZN(n653) );
  AOI22_X1 U553 ( .A1(data_in[1]), .A2(n825), .B1(n939), .B2(\mem[29][1] ), 
        .ZN(n938) );
  INV_X1 U554 ( .A(n937), .ZN(n652) );
  AOI22_X1 U555 ( .A1(data_in[2]), .A2(n825), .B1(n939), .B2(\mem[29][2] ), 
        .ZN(n937) );
  INV_X1 U556 ( .A(n936), .ZN(n651) );
  AOI22_X1 U557 ( .A1(data_in[3]), .A2(n825), .B1(n939), .B2(\mem[29][3] ), 
        .ZN(n936) );
  INV_X1 U558 ( .A(n935), .ZN(n650) );
  AOI22_X1 U559 ( .A1(data_in[4]), .A2(n825), .B1(n939), .B2(\mem[29][4] ), 
        .ZN(n935) );
  INV_X1 U560 ( .A(n934), .ZN(n649) );
  AOI22_X1 U561 ( .A1(data_in[5]), .A2(n825), .B1(n939), .B2(\mem[29][5] ), 
        .ZN(n934) );
  INV_X1 U562 ( .A(n933), .ZN(n648) );
  AOI22_X1 U563 ( .A1(data_in[6]), .A2(n825), .B1(n939), .B2(\mem[29][6] ), 
        .ZN(n933) );
  INV_X1 U564 ( .A(n932), .ZN(n647) );
  AOI22_X1 U565 ( .A1(data_in[7]), .A2(n825), .B1(n939), .B2(\mem[29][7] ), 
        .ZN(n932) );
  INV_X1 U566 ( .A(n931), .ZN(n646) );
  AOI22_X1 U567 ( .A1(data_in[0]), .A2(n824), .B1(n930), .B2(\mem[30][0] ), 
        .ZN(n931) );
  INV_X1 U568 ( .A(n929), .ZN(n645) );
  AOI22_X1 U569 ( .A1(data_in[1]), .A2(n824), .B1(n930), .B2(\mem[30][1] ), 
        .ZN(n929) );
  INV_X1 U570 ( .A(n928), .ZN(n644) );
  AOI22_X1 U571 ( .A1(data_in[2]), .A2(n824), .B1(n930), .B2(\mem[30][2] ), 
        .ZN(n928) );
  INV_X1 U572 ( .A(n927), .ZN(n643) );
  AOI22_X1 U573 ( .A1(data_in[3]), .A2(n824), .B1(n930), .B2(\mem[30][3] ), 
        .ZN(n927) );
  INV_X1 U574 ( .A(n926), .ZN(n642) );
  AOI22_X1 U575 ( .A1(data_in[4]), .A2(n824), .B1(n930), .B2(\mem[30][4] ), 
        .ZN(n926) );
  INV_X1 U576 ( .A(n925), .ZN(n641) );
  AOI22_X1 U577 ( .A1(data_in[5]), .A2(n824), .B1(n930), .B2(\mem[30][5] ), 
        .ZN(n925) );
  INV_X1 U578 ( .A(n924), .ZN(n640) );
  AOI22_X1 U579 ( .A1(data_in[6]), .A2(n824), .B1(n930), .B2(\mem[30][6] ), 
        .ZN(n924) );
  INV_X1 U580 ( .A(n923), .ZN(n639) );
  AOI22_X1 U581 ( .A1(data_in[7]), .A2(n824), .B1(n930), .B2(\mem[30][7] ), 
        .ZN(n923) );
  INV_X1 U582 ( .A(n922), .ZN(n638) );
  AOI22_X1 U583 ( .A1(data_in[0]), .A2(n823), .B1(n921), .B2(\mem[31][0] ), 
        .ZN(n922) );
  INV_X1 U584 ( .A(n920), .ZN(n637) );
  AOI22_X1 U585 ( .A1(data_in[1]), .A2(n823), .B1(n921), .B2(\mem[31][1] ), 
        .ZN(n920) );
  INV_X1 U586 ( .A(n919), .ZN(n636) );
  AOI22_X1 U587 ( .A1(data_in[2]), .A2(n823), .B1(n921), .B2(\mem[31][2] ), 
        .ZN(n919) );
  INV_X1 U588 ( .A(n918), .ZN(n635) );
  AOI22_X1 U589 ( .A1(data_in[3]), .A2(n823), .B1(n921), .B2(\mem[31][3] ), 
        .ZN(n918) );
  INV_X1 U590 ( .A(n917), .ZN(n634) );
  AOI22_X1 U591 ( .A1(data_in[4]), .A2(n823), .B1(n921), .B2(\mem[31][4] ), 
        .ZN(n917) );
  INV_X1 U592 ( .A(n916), .ZN(n633) );
  AOI22_X1 U593 ( .A1(data_in[5]), .A2(n823), .B1(n921), .B2(\mem[31][5] ), 
        .ZN(n916) );
  INV_X1 U594 ( .A(n915), .ZN(n632) );
  AOI22_X1 U595 ( .A1(data_in[6]), .A2(n823), .B1(n921), .B2(\mem[31][6] ), 
        .ZN(n915) );
  INV_X1 U596 ( .A(n914), .ZN(n631) );
  AOI22_X1 U597 ( .A1(data_in[7]), .A2(n823), .B1(n921), .B2(\mem[31][7] ), 
        .ZN(n914) );
  MUX2_X1 U598 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n614), .Z(n4) );
  MUX2_X1 U599 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n614), .Z(n5) );
  MUX2_X1 U600 ( .A(n5), .B(n4), .S(n611), .Z(n6) );
  MUX2_X1 U601 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n614), .Z(n7) );
  MUX2_X1 U602 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n614), .Z(n8) );
  MUX2_X1 U603 ( .A(n8), .B(n7), .S(n611), .Z(n9) );
  MUX2_X1 U604 ( .A(n9), .B(n6), .S(n609), .Z(n10) );
  MUX2_X1 U605 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n614), .Z(n11) );
  MUX2_X1 U606 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n614), .Z(n12) );
  MUX2_X1 U607 ( .A(n12), .B(n11), .S(n611), .Z(n13) );
  MUX2_X1 U608 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n614), .Z(n14) );
  MUX2_X1 U609 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n614), .Z(n15) );
  MUX2_X1 U610 ( .A(n15), .B(n14), .S(n611), .Z(n16) );
  MUX2_X1 U611 ( .A(n16), .B(n13), .S(N12), .Z(n17) );
  MUX2_X1 U612 ( .A(n17), .B(n10), .S(N13), .Z(n18) );
  MUX2_X1 U613 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n614), .Z(n19) );
  MUX2_X1 U614 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n620), .Z(n20) );
  MUX2_X1 U615 ( .A(n20), .B(n19), .S(n612), .Z(n21) );
  MUX2_X1 U616 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n620), .Z(n22) );
  MUX2_X1 U617 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n616), .Z(n23) );
  MUX2_X1 U618 ( .A(n23), .B(n22), .S(n612), .Z(n24) );
  MUX2_X1 U619 ( .A(n24), .B(n21), .S(N12), .Z(n25) );
  MUX2_X1 U620 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n620), .Z(n26) );
  MUX2_X1 U621 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n618), .Z(n27) );
  MUX2_X1 U622 ( .A(n27), .B(n26), .S(n612), .Z(n28) );
  MUX2_X1 U623 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n614), .Z(n29) );
  MUX2_X1 U624 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n615), .Z(n30) );
  MUX2_X1 U625 ( .A(n30), .B(n29), .S(n612), .Z(n31) );
  MUX2_X1 U626 ( .A(n31), .B(n28), .S(n610), .Z(n32) );
  MUX2_X1 U627 ( .A(n32), .B(n25), .S(N13), .Z(n33) );
  MUX2_X1 U628 ( .A(n33), .B(n18), .S(N14), .Z(N22) );
  MUX2_X1 U629 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n614), .Z(n34) );
  MUX2_X1 U630 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n620), .Z(n35) );
  MUX2_X1 U631 ( .A(n35), .B(n34), .S(n612), .Z(n36) );
  MUX2_X1 U632 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n620), .Z(n37) );
  MUX2_X1 U633 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n620), .Z(n38) );
  MUX2_X1 U634 ( .A(n38), .B(n37), .S(n612), .Z(n39) );
  MUX2_X1 U635 ( .A(n39), .B(n36), .S(n610), .Z(n40) );
  MUX2_X1 U636 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n620), .Z(n41) );
  MUX2_X1 U637 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n620), .Z(n42) );
  MUX2_X1 U638 ( .A(n42), .B(n41), .S(n612), .Z(n43) );
  MUX2_X1 U639 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n615), .Z(n44) );
  MUX2_X1 U640 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n620), .Z(n45) );
  MUX2_X1 U641 ( .A(n45), .B(n44), .S(n612), .Z(n46) );
  MUX2_X1 U642 ( .A(n46), .B(n43), .S(n609), .Z(n47) );
  MUX2_X1 U643 ( .A(n47), .B(n40), .S(N13), .Z(n48) );
  MUX2_X1 U644 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n620), .Z(n49) );
  MUX2_X1 U645 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n620), .Z(n50) );
  MUX2_X1 U646 ( .A(n50), .B(n49), .S(n612), .Z(n51) );
  MUX2_X1 U647 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n616), .Z(n52) );
  MUX2_X1 U648 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n620), .Z(n53) );
  MUX2_X1 U649 ( .A(n53), .B(n52), .S(n612), .Z(n54) );
  MUX2_X1 U650 ( .A(n54), .B(n51), .S(N12), .Z(n55) );
  MUX2_X1 U651 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n618), .Z(n56) );
  MUX2_X1 U652 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n620), .Z(n57) );
  MUX2_X1 U653 ( .A(n57), .B(n56), .S(n612), .Z(n58) );
  MUX2_X1 U654 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n620), .Z(n59) );
  MUX2_X1 U655 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n620), .Z(n60) );
  MUX2_X1 U656 ( .A(n60), .B(n59), .S(n612), .Z(n61) );
  MUX2_X1 U657 ( .A(n61), .B(n58), .S(n609), .Z(n62) );
  MUX2_X1 U658 ( .A(n62), .B(n55), .S(N13), .Z(n63) );
  MUX2_X1 U659 ( .A(n63), .B(n48), .S(N14), .Z(N21) );
  MUX2_X1 U660 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n617), .Z(n64) );
  MUX2_X1 U661 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n617), .Z(n65) );
  MUX2_X1 U662 ( .A(n65), .B(n64), .S(n613), .Z(n66) );
  MUX2_X1 U663 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n617), .Z(n67) );
  MUX2_X1 U664 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n617), .Z(n68) );
  MUX2_X1 U665 ( .A(n68), .B(n67), .S(n613), .Z(n69) );
  MUX2_X1 U666 ( .A(n69), .B(n66), .S(n609), .Z(n70) );
  MUX2_X1 U667 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n619), .Z(n71) );
  MUX2_X1 U668 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n619), .Z(n72) );
  MUX2_X1 U669 ( .A(n72), .B(n71), .S(n613), .Z(n73) );
  MUX2_X1 U670 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n617), .Z(n74) );
  MUX2_X1 U671 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n620), .Z(n75) );
  MUX2_X1 U672 ( .A(n75), .B(n74), .S(n613), .Z(n76) );
  MUX2_X1 U673 ( .A(n76), .B(n73), .S(n609), .Z(n77) );
  MUX2_X1 U674 ( .A(n77), .B(n70), .S(N13), .Z(n78) );
  MUX2_X1 U675 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n619), .Z(n79) );
  MUX2_X1 U676 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n619), .Z(n80) );
  MUX2_X1 U677 ( .A(n80), .B(n79), .S(n613), .Z(n81) );
  MUX2_X1 U678 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n619), .Z(n82) );
  MUX2_X1 U679 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n620), .Z(n83) );
  MUX2_X1 U680 ( .A(n83), .B(n82), .S(n613), .Z(n84) );
  MUX2_X1 U681 ( .A(n84), .B(n81), .S(n609), .Z(n85) );
  MUX2_X1 U682 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n617), .Z(n86) );
  MUX2_X1 U683 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n619), .Z(n87) );
  MUX2_X1 U684 ( .A(n87), .B(n86), .S(n613), .Z(n88) );
  MUX2_X1 U685 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n617), .Z(n89) );
  MUX2_X1 U686 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n619), .Z(n90) );
  MUX2_X1 U687 ( .A(n90), .B(n89), .S(n613), .Z(n91) );
  MUX2_X1 U688 ( .A(n91), .B(n88), .S(n609), .Z(n92) );
  MUX2_X1 U689 ( .A(n92), .B(n85), .S(N13), .Z(n93) );
  MUX2_X1 U690 ( .A(n93), .B(n78), .S(N14), .Z(N20) );
  MUX2_X1 U691 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n617), .Z(n94) );
  MUX2_X1 U692 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n619), .Z(n95) );
  MUX2_X1 U693 ( .A(n95), .B(n94), .S(n613), .Z(n96) );
  MUX2_X1 U694 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n619), .Z(n97) );
  MUX2_X1 U695 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n617), .Z(n98) );
  MUX2_X1 U696 ( .A(n98), .B(n97), .S(n613), .Z(n99) );
  MUX2_X1 U697 ( .A(n99), .B(n96), .S(n609), .Z(n100) );
  MUX2_X1 U698 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n617), .Z(n101) );
  MUX2_X1 U699 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n619), .Z(n102) );
  MUX2_X1 U700 ( .A(n102), .B(n101), .S(n613), .Z(n103) );
  MUX2_X1 U701 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n619), .Z(n104) );
  MUX2_X1 U702 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n617), .Z(n105) );
  MUX2_X1 U703 ( .A(n105), .B(n104), .S(n613), .Z(n106) );
  MUX2_X1 U704 ( .A(n106), .B(n103), .S(n609), .Z(n107) );
  MUX2_X1 U705 ( .A(n107), .B(n100), .S(N13), .Z(n108) );
  MUX2_X1 U706 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n615), .Z(n109) );
  MUX2_X1 U707 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n615), .Z(n110) );
  MUX2_X1 U708 ( .A(n110), .B(n109), .S(n612), .Z(n111) );
  MUX2_X1 U709 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n615), .Z(n112) );
  MUX2_X1 U710 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n615), .Z(n113) );
  MUX2_X1 U711 ( .A(n113), .B(n112), .S(n613), .Z(n114) );
  MUX2_X1 U712 ( .A(n114), .B(n111), .S(n609), .Z(n115) );
  MUX2_X1 U713 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n615), .Z(n116) );
  MUX2_X1 U714 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n615), .Z(n117) );
  MUX2_X1 U715 ( .A(n117), .B(n116), .S(n611), .Z(n118) );
  MUX2_X1 U716 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n615), .Z(n119) );
  MUX2_X1 U717 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n615), .Z(n120) );
  MUX2_X1 U718 ( .A(n120), .B(n119), .S(n611), .Z(n121) );
  MUX2_X1 U719 ( .A(n121), .B(n118), .S(n609), .Z(n122) );
  MUX2_X1 U720 ( .A(n122), .B(n115), .S(N13), .Z(n123) );
  MUX2_X1 U721 ( .A(n123), .B(n108), .S(N14), .Z(N19) );
  MUX2_X1 U722 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n615), .Z(n124) );
  MUX2_X1 U723 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n615), .Z(n125) );
  MUX2_X1 U724 ( .A(n125), .B(n124), .S(n611), .Z(n126) );
  MUX2_X1 U725 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n615), .Z(n127) );
  MUX2_X1 U726 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n615), .Z(n128) );
  MUX2_X1 U727 ( .A(n128), .B(n127), .S(n612), .Z(n129) );
  MUX2_X1 U728 ( .A(n129), .B(n126), .S(n609), .Z(n130) );
  MUX2_X1 U729 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n616), .Z(n131) );
  MUX2_X1 U730 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n616), .Z(n132) );
  MUX2_X1 U731 ( .A(n132), .B(n131), .S(N11), .Z(n133) );
  MUX2_X1 U732 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n616), .Z(n134) );
  MUX2_X1 U733 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n616), .Z(n135) );
  MUX2_X1 U734 ( .A(n135), .B(n134), .S(n612), .Z(n136) );
  MUX2_X1 U735 ( .A(n136), .B(n133), .S(n609), .Z(n137) );
  MUX2_X1 U736 ( .A(n137), .B(n130), .S(N13), .Z(n138) );
  MUX2_X1 U737 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n616), .Z(n139) );
  MUX2_X1 U738 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n616), .Z(n140) );
  MUX2_X1 U739 ( .A(n140), .B(n139), .S(n613), .Z(n141) );
  MUX2_X1 U740 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n616), .Z(n142) );
  MUX2_X1 U741 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n616), .Z(n143) );
  MUX2_X1 U742 ( .A(n143), .B(n142), .S(n611), .Z(n144) );
  MUX2_X1 U743 ( .A(n144), .B(n141), .S(n609), .Z(n145) );
  MUX2_X1 U744 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n616), .Z(n146) );
  MUX2_X1 U745 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n616), .Z(n147) );
  MUX2_X1 U746 ( .A(n147), .B(n146), .S(n612), .Z(n148) );
  MUX2_X1 U747 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n616), .Z(n149) );
  MUX2_X1 U748 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n616), .Z(n150) );
  MUX2_X1 U749 ( .A(n150), .B(n149), .S(n612), .Z(n151) );
  MUX2_X1 U750 ( .A(n151), .B(n148), .S(n609), .Z(n152) );
  MUX2_X1 U751 ( .A(n152), .B(n145), .S(N13), .Z(n153) );
  MUX2_X1 U752 ( .A(n153), .B(n138), .S(N14), .Z(N18) );
  MUX2_X1 U753 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n617), .Z(n154) );
  MUX2_X1 U754 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n617), .Z(n155) );
  MUX2_X1 U755 ( .A(n155), .B(n154), .S(n612), .Z(n156) );
  MUX2_X1 U756 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n617), .Z(n157) );
  MUX2_X1 U757 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n617), .Z(n158) );
  MUX2_X1 U758 ( .A(n158), .B(n157), .S(n613), .Z(n159) );
  MUX2_X1 U759 ( .A(n159), .B(n156), .S(n610), .Z(n160) );
  MUX2_X1 U760 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n617), .Z(n161) );
  MUX2_X1 U761 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n617), .Z(n162) );
  MUX2_X1 U762 ( .A(n162), .B(n161), .S(n611), .Z(n163) );
  MUX2_X1 U763 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n617), .Z(n164) );
  MUX2_X1 U764 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n617), .Z(n165) );
  MUX2_X1 U765 ( .A(n165), .B(n164), .S(N11), .Z(n166) );
  MUX2_X1 U766 ( .A(n166), .B(n163), .S(n610), .Z(n167) );
  MUX2_X1 U767 ( .A(n167), .B(n160), .S(N13), .Z(n168) );
  MUX2_X1 U768 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n617), .Z(n169) );
  MUX2_X1 U769 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n617), .Z(n170) );
  MUX2_X1 U770 ( .A(n170), .B(n169), .S(n611), .Z(n171) );
  MUX2_X1 U771 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n617), .Z(n172) );
  MUX2_X1 U772 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n617), .Z(n173) );
  MUX2_X1 U773 ( .A(n173), .B(n172), .S(N11), .Z(n174) );
  MUX2_X1 U774 ( .A(n174), .B(n171), .S(n610), .Z(n175) );
  MUX2_X1 U775 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n620), .Z(n176) );
  MUX2_X1 U776 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(N10), .Z(n177) );
  MUX2_X1 U777 ( .A(n177), .B(n176), .S(N11), .Z(n178) );
  MUX2_X1 U778 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n179) );
  MUX2_X1 U779 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n180) );
  MUX2_X1 U780 ( .A(n180), .B(n179), .S(n612), .Z(n181) );
  MUX2_X1 U781 ( .A(n181), .B(n178), .S(n610), .Z(n182) );
  MUX2_X1 U782 ( .A(n182), .B(n175), .S(N13), .Z(n183) );
  MUX2_X1 U783 ( .A(n183), .B(n168), .S(N14), .Z(N17) );
  MUX2_X1 U784 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n614), .Z(n184) );
  MUX2_X1 U785 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n620), .Z(n185) );
  MUX2_X1 U786 ( .A(n185), .B(n184), .S(n613), .Z(n186) );
  MUX2_X1 U787 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n614), .Z(n187) );
  MUX2_X1 U788 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(N10), .Z(n188) );
  MUX2_X1 U789 ( .A(n188), .B(n187), .S(n613), .Z(n189) );
  MUX2_X1 U790 ( .A(n189), .B(n186), .S(n610), .Z(n190) );
  MUX2_X1 U791 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n614), .Z(n191) );
  MUX2_X1 U792 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n620), .Z(n192) );
  MUX2_X1 U793 ( .A(n192), .B(n191), .S(n612), .Z(n193) );
  MUX2_X1 U794 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n620), .Z(n194) );
  MUX2_X1 U795 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(N10), .Z(n195) );
  MUX2_X1 U796 ( .A(n195), .B(n194), .S(N11), .Z(n196) );
  MUX2_X1 U797 ( .A(n196), .B(n193), .S(n610), .Z(n197) );
  MUX2_X1 U798 ( .A(n197), .B(n190), .S(N13), .Z(n198) );
  MUX2_X1 U799 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n618), .Z(n199) );
  MUX2_X1 U800 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n618), .Z(n200) );
  MUX2_X1 U801 ( .A(n200), .B(n199), .S(n611), .Z(n201) );
  MUX2_X1 U802 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n618), .Z(n202) );
  MUX2_X1 U803 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n618), .Z(n203) );
  MUX2_X1 U804 ( .A(n203), .B(n202), .S(n612), .Z(n204) );
  MUX2_X1 U805 ( .A(n204), .B(n201), .S(n610), .Z(n205) );
  MUX2_X1 U806 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n618), .Z(n206) );
  MUX2_X1 U807 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n618), .Z(n207) );
  MUX2_X1 U808 ( .A(n207), .B(n206), .S(n611), .Z(n208) );
  MUX2_X1 U809 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n618), .Z(n209) );
  MUX2_X1 U810 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n618), .Z(n210) );
  MUX2_X1 U811 ( .A(n210), .B(n209), .S(n613), .Z(n211) );
  MUX2_X1 U812 ( .A(n211), .B(n208), .S(n610), .Z(n212) );
  MUX2_X1 U813 ( .A(n212), .B(n205), .S(N13), .Z(n213) );
  MUX2_X1 U814 ( .A(n213), .B(n198), .S(N14), .Z(N16) );
  MUX2_X1 U815 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n618), .Z(n214) );
  MUX2_X1 U816 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n618), .Z(n215) );
  MUX2_X1 U817 ( .A(n215), .B(n214), .S(n611), .Z(n216) );
  MUX2_X1 U818 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n618), .Z(n217) );
  MUX2_X1 U819 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n618), .Z(n218) );
  MUX2_X1 U820 ( .A(n218), .B(n217), .S(n611), .Z(n219) );
  MUX2_X1 U821 ( .A(n219), .B(n216), .S(n610), .Z(n220) );
  MUX2_X1 U822 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n619), .Z(n221) );
  MUX2_X1 U823 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n619), .Z(n222) );
  MUX2_X1 U824 ( .A(n222), .B(n221), .S(n611), .Z(n223) );
  MUX2_X1 U825 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n619), .Z(n224) );
  MUX2_X1 U826 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n619), .Z(n225) );
  MUX2_X1 U827 ( .A(n225), .B(n224), .S(n613), .Z(n226) );
  MUX2_X1 U828 ( .A(n226), .B(n223), .S(n610), .Z(n227) );
  MUX2_X1 U829 ( .A(n227), .B(n220), .S(N13), .Z(n228) );
  MUX2_X1 U830 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n619), .Z(n229) );
  MUX2_X1 U831 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n619), .Z(n595) );
  MUX2_X1 U832 ( .A(n595), .B(n229), .S(n611), .Z(n596) );
  MUX2_X1 U833 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n619), .Z(n597) );
  MUX2_X1 U834 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n619), .Z(n598) );
  MUX2_X1 U835 ( .A(n598), .B(n597), .S(n613), .Z(n599) );
  MUX2_X1 U836 ( .A(n599), .B(n596), .S(n610), .Z(n600) );
  MUX2_X1 U837 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n619), .Z(n601) );
  MUX2_X1 U838 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n619), .Z(n602) );
  MUX2_X1 U839 ( .A(n602), .B(n601), .S(n611), .Z(n603) );
  MUX2_X1 U840 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n619), .Z(n604) );
  MUX2_X1 U841 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n619), .Z(n605) );
  MUX2_X1 U842 ( .A(n605), .B(n604), .S(n611), .Z(n606) );
  MUX2_X1 U843 ( .A(n606), .B(n603), .S(n610), .Z(n607) );
  MUX2_X1 U844 ( .A(n607), .B(n600), .S(N13), .Z(n608) );
  MUX2_X1 U845 ( .A(n608), .B(n228), .S(N14), .Z(N15) );
  CLKBUF_X1 U846 ( .A(N11), .Z(n611) );
  CLKBUF_X1 U847 ( .A(n620), .Z(n614) );
  INV_X1 U848 ( .A(N10), .ZN(n621) );
  INV_X1 U849 ( .A(N11), .ZN(n622) );
  INV_X1 U850 ( .A(data_in[0]), .ZN(n623) );
  INV_X1 U851 ( .A(data_in[1]), .ZN(n624) );
  INV_X1 U852 ( .A(data_in[2]), .ZN(n625) );
  INV_X1 U853 ( .A(data_in[3]), .ZN(n626) );
  INV_X1 U854 ( .A(data_in[4]), .ZN(n627) );
  INV_X1 U855 ( .A(data_in[5]), .ZN(n628) );
  INV_X1 U856 ( .A(data_in[6]), .ZN(n629) );
  INV_X1 U857 ( .A(data_in[7]), .ZN(n630) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_21 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n629), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n630), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n631), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n632), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n633), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n634), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n635), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n636), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n637), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n638), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n639), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n640), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n641), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n642), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n643), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n644), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n645), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n646), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n647), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n648), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n649), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n650), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n651), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n652), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n653), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n654), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n655), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n656), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n657), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n658), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n659), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n660), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n661), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n662), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n663), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n664), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n665), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n666), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n667), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n668), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n669), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n670), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n671), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n672), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n673), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n674), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n675), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n676), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n677), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n678), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n679), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n680), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n681), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n682), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n683), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n684), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n685), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n686), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n687), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n688), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n689), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n690), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n691), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n692), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n693), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n694), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n695), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n696), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n697), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n698), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n699), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n700), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n701), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n702), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n703), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n704), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n705), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n706), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n707), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n708), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n709), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n710), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n711), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n712), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n713), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n714), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n715), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n716), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n717), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n718), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n719), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n720), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n721), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n722), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n723), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n724), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n725), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n726), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n727), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n728), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n729), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n730), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n731), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n732), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n733), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n734), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n735), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n736), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n737), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n738), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n739), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n740), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n741), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n742), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n743), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n744), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n745), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n746), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n747), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n748), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n749), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n750), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n751), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n752), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n753), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n754), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n755), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n756), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n757), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n758), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n759), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n760), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n761), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n762), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n763), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n764), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n765), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n766), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n767), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n768), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n769), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n770), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n771), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n772), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n773), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n774), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n775), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n776), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n777), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n778), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n779), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n780), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n781), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n782), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n783), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n784), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n785), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n786), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n787), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n788), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n789), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n790), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n791), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n792), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n793), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n794), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n795), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n796), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n797), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n798), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n799), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n800), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n801), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n802), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n803), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n804), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n805), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n806), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n807), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n808), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n809), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n810), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n811), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n812), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n813), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n814), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n815), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n816), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n817), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n818), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n819), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n820), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n848), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n849), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n850), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n851), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n852), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n853), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n854), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n855), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n856), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n857), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n858), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n859), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n860), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n861), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n862), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n863), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n864), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n865), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n866), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n867), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n868), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n869), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n870), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n871), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n872), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n873), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n874), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n875), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n876), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n877), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n878), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n879), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n880), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n881), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n882), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n883), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n884), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n885), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n886), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n887), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n888), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n889), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n890), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n891), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n892), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n893), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n894), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n895), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n896), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n897), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n898), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n899), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n900), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n901), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n902), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n903), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n904), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n905), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n906), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n907), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n908), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n909), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n910), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n911), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[5]) );
  BUF_X1 U4 ( .A(n618), .Z(n617) );
  BUF_X1 U5 ( .A(n618), .Z(n614) );
  BUF_X1 U6 ( .A(N10), .Z(n615) );
  BUF_X1 U7 ( .A(n618), .Z(n616) );
  BUF_X1 U8 ( .A(n618), .Z(n613) );
  BUF_X1 U9 ( .A(N11), .Z(n611) );
  BUF_X1 U10 ( .A(N11), .Z(n612) );
  BUF_X1 U11 ( .A(N10), .Z(n618) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1203) );
  NOR3_X1 U13 ( .A1(N11), .A2(N12), .A3(n619), .ZN(n1192) );
  NOR3_X1 U14 ( .A1(N10), .A2(N12), .A3(n620), .ZN(n1182) );
  NOR3_X1 U15 ( .A1(n619), .A2(N12), .A3(n620), .ZN(n1172) );
  INV_X1 U16 ( .A(n1129), .ZN(n844) );
  INV_X1 U17 ( .A(n1119), .ZN(n843) );
  INV_X1 U18 ( .A(n1110), .ZN(n842) );
  INV_X1 U19 ( .A(n1101), .ZN(n841) );
  INV_X1 U20 ( .A(n1056), .ZN(n836) );
  INV_X1 U21 ( .A(n1046), .ZN(n835) );
  INV_X1 U22 ( .A(n1037), .ZN(n834) );
  INV_X1 U23 ( .A(n1028), .ZN(n833) );
  INV_X1 U24 ( .A(n983), .ZN(n828) );
  INV_X1 U25 ( .A(n973), .ZN(n827) );
  INV_X1 U26 ( .A(n964), .ZN(n826) );
  INV_X1 U27 ( .A(n955), .ZN(n825) );
  INV_X1 U28 ( .A(n946), .ZN(n824) );
  INV_X1 U29 ( .A(n937), .ZN(n823) );
  INV_X1 U30 ( .A(n928), .ZN(n822) );
  INV_X1 U31 ( .A(n919), .ZN(n821) );
  INV_X1 U32 ( .A(n1092), .ZN(n840) );
  INV_X1 U33 ( .A(n1083), .ZN(n839) );
  INV_X1 U34 ( .A(n1074), .ZN(n838) );
  INV_X1 U35 ( .A(n1065), .ZN(n837) );
  INV_X1 U36 ( .A(n1019), .ZN(n832) );
  INV_X1 U37 ( .A(n1010), .ZN(n831) );
  INV_X1 U38 ( .A(n1001), .ZN(n830) );
  INV_X1 U39 ( .A(n992), .ZN(n829) );
  BUF_X1 U40 ( .A(N12), .Z(n608) );
  BUF_X1 U41 ( .A(N12), .Z(n609) );
  INV_X1 U42 ( .A(N13), .ZN(n846) );
  AND3_X1 U43 ( .A1(n619), .A2(n620), .A3(N12), .ZN(n1162) );
  AND3_X1 U44 ( .A1(N10), .A2(n620), .A3(N12), .ZN(n1152) );
  AND3_X1 U45 ( .A1(N11), .A2(n619), .A3(N12), .ZN(n1142) );
  AND3_X1 U46 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1132) );
  INV_X1 U47 ( .A(N14), .ZN(n847) );
  NAND2_X1 U48 ( .A1(n1192), .A2(n1202), .ZN(n1201) );
  NAND2_X1 U49 ( .A1(n1182), .A2(n1202), .ZN(n1191) );
  NAND2_X1 U50 ( .A1(n1172), .A2(n1202), .ZN(n1181) );
  NAND2_X1 U51 ( .A1(n1162), .A2(n1202), .ZN(n1171) );
  NAND2_X1 U52 ( .A1(n1152), .A2(n1202), .ZN(n1161) );
  NAND2_X1 U53 ( .A1(n1142), .A2(n1202), .ZN(n1151) );
  NAND2_X1 U54 ( .A1(n1132), .A2(n1202), .ZN(n1141) );
  NAND2_X1 U55 ( .A1(n1203), .A2(n1202), .ZN(n1212) );
  NAND2_X1 U56 ( .A1(n1121), .A2(n1203), .ZN(n1129) );
  NAND2_X1 U57 ( .A1(n1121), .A2(n1192), .ZN(n1119) );
  NAND2_X1 U58 ( .A1(n1121), .A2(n1182), .ZN(n1110) );
  NAND2_X1 U59 ( .A1(n1121), .A2(n1172), .ZN(n1101) );
  NAND2_X1 U60 ( .A1(n1048), .A2(n1203), .ZN(n1056) );
  NAND2_X1 U61 ( .A1(n1048), .A2(n1192), .ZN(n1046) );
  NAND2_X1 U62 ( .A1(n1048), .A2(n1182), .ZN(n1037) );
  NAND2_X1 U63 ( .A1(n1048), .A2(n1172), .ZN(n1028) );
  NAND2_X1 U64 ( .A1(n975), .A2(n1203), .ZN(n983) );
  NAND2_X1 U65 ( .A1(n975), .A2(n1192), .ZN(n973) );
  NAND2_X1 U66 ( .A1(n975), .A2(n1182), .ZN(n964) );
  NAND2_X1 U67 ( .A1(n975), .A2(n1172), .ZN(n955) );
  NAND2_X1 U68 ( .A1(n1121), .A2(n1162), .ZN(n1092) );
  NAND2_X1 U69 ( .A1(n1121), .A2(n1152), .ZN(n1083) );
  NAND2_X1 U70 ( .A1(n1121), .A2(n1142), .ZN(n1074) );
  NAND2_X1 U71 ( .A1(n1121), .A2(n1132), .ZN(n1065) );
  NAND2_X1 U72 ( .A1(n1048), .A2(n1162), .ZN(n1019) );
  NAND2_X1 U73 ( .A1(n1048), .A2(n1152), .ZN(n1010) );
  NAND2_X1 U74 ( .A1(n1048), .A2(n1142), .ZN(n1001) );
  NAND2_X1 U75 ( .A1(n1048), .A2(n1132), .ZN(n992) );
  NAND2_X1 U76 ( .A1(n975), .A2(n1162), .ZN(n946) );
  NAND2_X1 U77 ( .A1(n975), .A2(n1152), .ZN(n937) );
  NAND2_X1 U78 ( .A1(n975), .A2(n1142), .ZN(n928) );
  NAND2_X1 U79 ( .A1(n975), .A2(n1132), .ZN(n919) );
  AND3_X1 U80 ( .A1(n846), .A2(n847), .A3(n1131), .ZN(n1202) );
  AND3_X1 U81 ( .A1(N13), .A2(n1131), .A3(N14), .ZN(n975) );
  AND3_X1 U82 ( .A1(n1131), .A2(n847), .A3(N13), .ZN(n1121) );
  AND3_X1 U83 ( .A1(n1131), .A2(n846), .A3(N14), .ZN(n1048) );
  NOR2_X1 U84 ( .A1(n845), .A2(addr[5]), .ZN(n1131) );
  INV_X1 U85 ( .A(wr_en), .ZN(n845) );
  OAI21_X1 U86 ( .B1(n621), .B2(n1171), .A(n1170), .ZN(n879) );
  NAND2_X1 U87 ( .A1(\mem[4][0] ), .A2(n1171), .ZN(n1170) );
  OAI21_X1 U88 ( .B1(n622), .B2(n1171), .A(n1169), .ZN(n878) );
  NAND2_X1 U89 ( .A1(\mem[4][1] ), .A2(n1171), .ZN(n1169) );
  OAI21_X1 U90 ( .B1(n623), .B2(n1171), .A(n1168), .ZN(n877) );
  NAND2_X1 U91 ( .A1(\mem[4][2] ), .A2(n1171), .ZN(n1168) );
  OAI21_X1 U92 ( .B1(n624), .B2(n1171), .A(n1167), .ZN(n876) );
  NAND2_X1 U93 ( .A1(\mem[4][3] ), .A2(n1171), .ZN(n1167) );
  OAI21_X1 U94 ( .B1(n625), .B2(n1171), .A(n1166), .ZN(n875) );
  NAND2_X1 U95 ( .A1(\mem[4][4] ), .A2(n1171), .ZN(n1166) );
  OAI21_X1 U96 ( .B1(n626), .B2(n1171), .A(n1165), .ZN(n874) );
  NAND2_X1 U97 ( .A1(\mem[4][5] ), .A2(n1171), .ZN(n1165) );
  OAI21_X1 U98 ( .B1(n627), .B2(n1171), .A(n1164), .ZN(n873) );
  NAND2_X1 U99 ( .A1(\mem[4][6] ), .A2(n1171), .ZN(n1164) );
  OAI21_X1 U100 ( .B1(n628), .B2(n1171), .A(n1163), .ZN(n872) );
  NAND2_X1 U101 ( .A1(\mem[4][7] ), .A2(n1171), .ZN(n1163) );
  OAI21_X1 U102 ( .B1(n621), .B2(n1151), .A(n1150), .ZN(n863) );
  NAND2_X1 U103 ( .A1(\mem[6][0] ), .A2(n1151), .ZN(n1150) );
  OAI21_X1 U104 ( .B1(n622), .B2(n1151), .A(n1149), .ZN(n862) );
  NAND2_X1 U105 ( .A1(\mem[6][1] ), .A2(n1151), .ZN(n1149) );
  OAI21_X1 U106 ( .B1(n623), .B2(n1151), .A(n1148), .ZN(n861) );
  NAND2_X1 U107 ( .A1(\mem[6][2] ), .A2(n1151), .ZN(n1148) );
  OAI21_X1 U108 ( .B1(n624), .B2(n1151), .A(n1147), .ZN(n860) );
  NAND2_X1 U109 ( .A1(\mem[6][3] ), .A2(n1151), .ZN(n1147) );
  OAI21_X1 U110 ( .B1(n625), .B2(n1151), .A(n1146), .ZN(n859) );
  NAND2_X1 U111 ( .A1(\mem[6][4] ), .A2(n1151), .ZN(n1146) );
  OAI21_X1 U112 ( .B1(n626), .B2(n1151), .A(n1145), .ZN(n858) );
  NAND2_X1 U113 ( .A1(\mem[6][5] ), .A2(n1151), .ZN(n1145) );
  OAI21_X1 U114 ( .B1(n627), .B2(n1151), .A(n1144), .ZN(n857) );
  NAND2_X1 U115 ( .A1(\mem[6][6] ), .A2(n1151), .ZN(n1144) );
  OAI21_X1 U116 ( .B1(n628), .B2(n1151), .A(n1143), .ZN(n856) );
  NAND2_X1 U117 ( .A1(\mem[6][7] ), .A2(n1151), .ZN(n1143) );
  OAI21_X1 U118 ( .B1(n621), .B2(n1141), .A(n1140), .ZN(n855) );
  NAND2_X1 U119 ( .A1(\mem[7][0] ), .A2(n1141), .ZN(n1140) );
  OAI21_X1 U120 ( .B1(n622), .B2(n1141), .A(n1139), .ZN(n854) );
  NAND2_X1 U121 ( .A1(\mem[7][1] ), .A2(n1141), .ZN(n1139) );
  OAI21_X1 U122 ( .B1(n623), .B2(n1141), .A(n1138), .ZN(n853) );
  NAND2_X1 U123 ( .A1(\mem[7][2] ), .A2(n1141), .ZN(n1138) );
  OAI21_X1 U124 ( .B1(n624), .B2(n1141), .A(n1137), .ZN(n852) );
  NAND2_X1 U125 ( .A1(\mem[7][3] ), .A2(n1141), .ZN(n1137) );
  OAI21_X1 U126 ( .B1(n625), .B2(n1141), .A(n1136), .ZN(n851) );
  NAND2_X1 U127 ( .A1(\mem[7][4] ), .A2(n1141), .ZN(n1136) );
  OAI21_X1 U128 ( .B1(n626), .B2(n1141), .A(n1135), .ZN(n850) );
  NAND2_X1 U129 ( .A1(\mem[7][5] ), .A2(n1141), .ZN(n1135) );
  OAI21_X1 U130 ( .B1(n627), .B2(n1141), .A(n1134), .ZN(n849) );
  NAND2_X1 U131 ( .A1(\mem[7][6] ), .A2(n1141), .ZN(n1134) );
  OAI21_X1 U132 ( .B1(n628), .B2(n1141), .A(n1133), .ZN(n848) );
  NAND2_X1 U133 ( .A1(\mem[7][7] ), .A2(n1141), .ZN(n1133) );
  OAI21_X1 U134 ( .B1(n621), .B2(n1201), .A(n1200), .ZN(n903) );
  NAND2_X1 U135 ( .A1(\mem[1][0] ), .A2(n1201), .ZN(n1200) );
  OAI21_X1 U136 ( .B1(n622), .B2(n1201), .A(n1199), .ZN(n902) );
  NAND2_X1 U137 ( .A1(\mem[1][1] ), .A2(n1201), .ZN(n1199) );
  OAI21_X1 U138 ( .B1(n623), .B2(n1201), .A(n1198), .ZN(n901) );
  NAND2_X1 U139 ( .A1(\mem[1][2] ), .A2(n1201), .ZN(n1198) );
  OAI21_X1 U140 ( .B1(n624), .B2(n1201), .A(n1197), .ZN(n900) );
  NAND2_X1 U141 ( .A1(\mem[1][3] ), .A2(n1201), .ZN(n1197) );
  OAI21_X1 U142 ( .B1(n625), .B2(n1201), .A(n1196), .ZN(n899) );
  NAND2_X1 U143 ( .A1(\mem[1][4] ), .A2(n1201), .ZN(n1196) );
  OAI21_X1 U144 ( .B1(n626), .B2(n1201), .A(n1195), .ZN(n898) );
  NAND2_X1 U145 ( .A1(\mem[1][5] ), .A2(n1201), .ZN(n1195) );
  OAI21_X1 U146 ( .B1(n627), .B2(n1201), .A(n1194), .ZN(n897) );
  NAND2_X1 U147 ( .A1(\mem[1][6] ), .A2(n1201), .ZN(n1194) );
  OAI21_X1 U148 ( .B1(n628), .B2(n1201), .A(n1193), .ZN(n896) );
  NAND2_X1 U149 ( .A1(\mem[1][7] ), .A2(n1201), .ZN(n1193) );
  OAI21_X1 U150 ( .B1(n621), .B2(n1191), .A(n1190), .ZN(n895) );
  NAND2_X1 U151 ( .A1(\mem[2][0] ), .A2(n1191), .ZN(n1190) );
  OAI21_X1 U152 ( .B1(n622), .B2(n1191), .A(n1189), .ZN(n894) );
  NAND2_X1 U153 ( .A1(\mem[2][1] ), .A2(n1191), .ZN(n1189) );
  OAI21_X1 U154 ( .B1(n623), .B2(n1191), .A(n1188), .ZN(n893) );
  NAND2_X1 U155 ( .A1(\mem[2][2] ), .A2(n1191), .ZN(n1188) );
  OAI21_X1 U156 ( .B1(n624), .B2(n1191), .A(n1187), .ZN(n892) );
  NAND2_X1 U157 ( .A1(\mem[2][3] ), .A2(n1191), .ZN(n1187) );
  OAI21_X1 U158 ( .B1(n625), .B2(n1191), .A(n1186), .ZN(n891) );
  NAND2_X1 U159 ( .A1(\mem[2][4] ), .A2(n1191), .ZN(n1186) );
  OAI21_X1 U160 ( .B1(n626), .B2(n1191), .A(n1185), .ZN(n890) );
  NAND2_X1 U161 ( .A1(\mem[2][5] ), .A2(n1191), .ZN(n1185) );
  OAI21_X1 U162 ( .B1(n627), .B2(n1191), .A(n1184), .ZN(n889) );
  NAND2_X1 U163 ( .A1(\mem[2][6] ), .A2(n1191), .ZN(n1184) );
  OAI21_X1 U164 ( .B1(n628), .B2(n1191), .A(n1183), .ZN(n888) );
  NAND2_X1 U165 ( .A1(\mem[2][7] ), .A2(n1191), .ZN(n1183) );
  OAI21_X1 U166 ( .B1(n621), .B2(n1181), .A(n1180), .ZN(n887) );
  NAND2_X1 U167 ( .A1(\mem[3][0] ), .A2(n1181), .ZN(n1180) );
  OAI21_X1 U168 ( .B1(n622), .B2(n1181), .A(n1179), .ZN(n886) );
  NAND2_X1 U169 ( .A1(\mem[3][1] ), .A2(n1181), .ZN(n1179) );
  OAI21_X1 U170 ( .B1(n623), .B2(n1181), .A(n1178), .ZN(n885) );
  NAND2_X1 U171 ( .A1(\mem[3][2] ), .A2(n1181), .ZN(n1178) );
  OAI21_X1 U172 ( .B1(n624), .B2(n1181), .A(n1177), .ZN(n884) );
  NAND2_X1 U173 ( .A1(\mem[3][3] ), .A2(n1181), .ZN(n1177) );
  OAI21_X1 U174 ( .B1(n625), .B2(n1181), .A(n1176), .ZN(n883) );
  NAND2_X1 U175 ( .A1(\mem[3][4] ), .A2(n1181), .ZN(n1176) );
  OAI21_X1 U176 ( .B1(n626), .B2(n1181), .A(n1175), .ZN(n882) );
  NAND2_X1 U177 ( .A1(\mem[3][5] ), .A2(n1181), .ZN(n1175) );
  OAI21_X1 U178 ( .B1(n627), .B2(n1181), .A(n1174), .ZN(n881) );
  NAND2_X1 U179 ( .A1(\mem[3][6] ), .A2(n1181), .ZN(n1174) );
  OAI21_X1 U180 ( .B1(n628), .B2(n1181), .A(n1173), .ZN(n880) );
  NAND2_X1 U181 ( .A1(\mem[3][7] ), .A2(n1181), .ZN(n1173) );
  OAI21_X1 U182 ( .B1(n621), .B2(n1161), .A(n1160), .ZN(n871) );
  NAND2_X1 U183 ( .A1(\mem[5][0] ), .A2(n1161), .ZN(n1160) );
  OAI21_X1 U184 ( .B1(n622), .B2(n1161), .A(n1159), .ZN(n870) );
  NAND2_X1 U185 ( .A1(\mem[5][1] ), .A2(n1161), .ZN(n1159) );
  OAI21_X1 U186 ( .B1(n623), .B2(n1161), .A(n1158), .ZN(n869) );
  NAND2_X1 U187 ( .A1(\mem[5][2] ), .A2(n1161), .ZN(n1158) );
  OAI21_X1 U188 ( .B1(n624), .B2(n1161), .A(n1157), .ZN(n868) );
  NAND2_X1 U189 ( .A1(\mem[5][3] ), .A2(n1161), .ZN(n1157) );
  OAI21_X1 U190 ( .B1(n625), .B2(n1161), .A(n1156), .ZN(n867) );
  NAND2_X1 U191 ( .A1(\mem[5][4] ), .A2(n1161), .ZN(n1156) );
  OAI21_X1 U192 ( .B1(n626), .B2(n1161), .A(n1155), .ZN(n866) );
  NAND2_X1 U193 ( .A1(\mem[5][5] ), .A2(n1161), .ZN(n1155) );
  OAI21_X1 U194 ( .B1(n627), .B2(n1161), .A(n1154), .ZN(n865) );
  NAND2_X1 U195 ( .A1(\mem[5][6] ), .A2(n1161), .ZN(n1154) );
  OAI21_X1 U196 ( .B1(n628), .B2(n1161), .A(n1153), .ZN(n864) );
  NAND2_X1 U197 ( .A1(\mem[5][7] ), .A2(n1161), .ZN(n1153) );
  OAI21_X1 U198 ( .B1(n1212), .B2(n621), .A(n1211), .ZN(n911) );
  NAND2_X1 U199 ( .A1(\mem[0][0] ), .A2(n1212), .ZN(n1211) );
  OAI21_X1 U200 ( .B1(n1212), .B2(n622), .A(n1210), .ZN(n910) );
  NAND2_X1 U201 ( .A1(\mem[0][1] ), .A2(n1212), .ZN(n1210) );
  OAI21_X1 U202 ( .B1(n1212), .B2(n623), .A(n1209), .ZN(n909) );
  NAND2_X1 U203 ( .A1(\mem[0][2] ), .A2(n1212), .ZN(n1209) );
  OAI21_X1 U204 ( .B1(n1212), .B2(n624), .A(n1208), .ZN(n908) );
  NAND2_X1 U205 ( .A1(\mem[0][3] ), .A2(n1212), .ZN(n1208) );
  OAI21_X1 U206 ( .B1(n1212), .B2(n625), .A(n1207), .ZN(n907) );
  NAND2_X1 U207 ( .A1(\mem[0][4] ), .A2(n1212), .ZN(n1207) );
  OAI21_X1 U208 ( .B1(n1212), .B2(n626), .A(n1206), .ZN(n906) );
  NAND2_X1 U209 ( .A1(\mem[0][5] ), .A2(n1212), .ZN(n1206) );
  OAI21_X1 U210 ( .B1(n1212), .B2(n627), .A(n1205), .ZN(n905) );
  NAND2_X1 U211 ( .A1(\mem[0][6] ), .A2(n1212), .ZN(n1205) );
  OAI21_X1 U212 ( .B1(n1212), .B2(n628), .A(n1204), .ZN(n904) );
  NAND2_X1 U213 ( .A1(\mem[0][7] ), .A2(n1212), .ZN(n1204) );
  INV_X1 U214 ( .A(n1130), .ZN(n820) );
  AOI22_X1 U215 ( .A1(data_in[0]), .A2(n844), .B1(n1129), .B2(\mem[8][0] ), 
        .ZN(n1130) );
  INV_X1 U216 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U217 ( .A1(data_in[1]), .A2(n844), .B1(n1129), .B2(\mem[8][1] ), 
        .ZN(n1128) );
  INV_X1 U218 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U219 ( .A1(data_in[2]), .A2(n844), .B1(n1129), .B2(\mem[8][2] ), 
        .ZN(n1127) );
  INV_X1 U220 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U221 ( .A1(data_in[3]), .A2(n844), .B1(n1129), .B2(\mem[8][3] ), 
        .ZN(n1126) );
  INV_X1 U222 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U223 ( .A1(data_in[4]), .A2(n844), .B1(n1129), .B2(\mem[8][4] ), 
        .ZN(n1125) );
  INV_X1 U224 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U225 ( .A1(data_in[5]), .A2(n844), .B1(n1129), .B2(\mem[8][5] ), 
        .ZN(n1124) );
  INV_X1 U226 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U227 ( .A1(data_in[6]), .A2(n844), .B1(n1129), .B2(\mem[8][6] ), 
        .ZN(n1123) );
  INV_X1 U228 ( .A(n1122), .ZN(n813) );
  AOI22_X1 U229 ( .A1(data_in[7]), .A2(n844), .B1(n1129), .B2(\mem[8][7] ), 
        .ZN(n1122) );
  INV_X1 U230 ( .A(n1120), .ZN(n812) );
  AOI22_X1 U231 ( .A1(data_in[0]), .A2(n843), .B1(n1119), .B2(\mem[9][0] ), 
        .ZN(n1120) );
  INV_X1 U232 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U233 ( .A1(data_in[1]), .A2(n843), .B1(n1119), .B2(\mem[9][1] ), 
        .ZN(n1118) );
  INV_X1 U234 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U235 ( .A1(data_in[2]), .A2(n843), .B1(n1119), .B2(\mem[9][2] ), 
        .ZN(n1117) );
  INV_X1 U236 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U237 ( .A1(data_in[3]), .A2(n843), .B1(n1119), .B2(\mem[9][3] ), 
        .ZN(n1116) );
  INV_X1 U238 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U239 ( .A1(data_in[4]), .A2(n843), .B1(n1119), .B2(\mem[9][4] ), 
        .ZN(n1115) );
  INV_X1 U240 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U241 ( .A1(data_in[5]), .A2(n843), .B1(n1119), .B2(\mem[9][5] ), 
        .ZN(n1114) );
  INV_X1 U242 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U243 ( .A1(data_in[6]), .A2(n843), .B1(n1119), .B2(\mem[9][6] ), 
        .ZN(n1113) );
  INV_X1 U244 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U245 ( .A1(data_in[7]), .A2(n843), .B1(n1119), .B2(\mem[9][7] ), 
        .ZN(n1112) );
  INV_X1 U246 ( .A(n1111), .ZN(n804) );
  AOI22_X1 U247 ( .A1(data_in[0]), .A2(n842), .B1(n1110), .B2(\mem[10][0] ), 
        .ZN(n1111) );
  INV_X1 U248 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U249 ( .A1(data_in[1]), .A2(n842), .B1(n1110), .B2(\mem[10][1] ), 
        .ZN(n1109) );
  INV_X1 U250 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U251 ( .A1(data_in[2]), .A2(n842), .B1(n1110), .B2(\mem[10][2] ), 
        .ZN(n1108) );
  INV_X1 U252 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U253 ( .A1(data_in[3]), .A2(n842), .B1(n1110), .B2(\mem[10][3] ), 
        .ZN(n1107) );
  INV_X1 U254 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U255 ( .A1(data_in[4]), .A2(n842), .B1(n1110), .B2(\mem[10][4] ), 
        .ZN(n1106) );
  INV_X1 U256 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U257 ( .A1(data_in[5]), .A2(n842), .B1(n1110), .B2(\mem[10][5] ), 
        .ZN(n1105) );
  INV_X1 U258 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U259 ( .A1(data_in[6]), .A2(n842), .B1(n1110), .B2(\mem[10][6] ), 
        .ZN(n1104) );
  INV_X1 U260 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U261 ( .A1(data_in[7]), .A2(n842), .B1(n1110), .B2(\mem[10][7] ), 
        .ZN(n1103) );
  INV_X1 U262 ( .A(n1102), .ZN(n796) );
  AOI22_X1 U263 ( .A1(data_in[0]), .A2(n841), .B1(n1101), .B2(\mem[11][0] ), 
        .ZN(n1102) );
  INV_X1 U264 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U265 ( .A1(data_in[1]), .A2(n841), .B1(n1101), .B2(\mem[11][1] ), 
        .ZN(n1100) );
  INV_X1 U266 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U267 ( .A1(data_in[2]), .A2(n841), .B1(n1101), .B2(\mem[11][2] ), 
        .ZN(n1099) );
  INV_X1 U268 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U269 ( .A1(data_in[3]), .A2(n841), .B1(n1101), .B2(\mem[11][3] ), 
        .ZN(n1098) );
  INV_X1 U270 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U271 ( .A1(data_in[4]), .A2(n841), .B1(n1101), .B2(\mem[11][4] ), 
        .ZN(n1097) );
  INV_X1 U272 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U273 ( .A1(data_in[5]), .A2(n841), .B1(n1101), .B2(\mem[11][5] ), 
        .ZN(n1096) );
  INV_X1 U274 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U275 ( .A1(data_in[6]), .A2(n841), .B1(n1101), .B2(\mem[11][6] ), 
        .ZN(n1095) );
  INV_X1 U276 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U277 ( .A1(data_in[7]), .A2(n841), .B1(n1101), .B2(\mem[11][7] ), 
        .ZN(n1094) );
  INV_X1 U278 ( .A(n1093), .ZN(n788) );
  AOI22_X1 U279 ( .A1(data_in[0]), .A2(n840), .B1(n1092), .B2(\mem[12][0] ), 
        .ZN(n1093) );
  INV_X1 U280 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U281 ( .A1(data_in[1]), .A2(n840), .B1(n1092), .B2(\mem[12][1] ), 
        .ZN(n1091) );
  INV_X1 U282 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U283 ( .A1(data_in[2]), .A2(n840), .B1(n1092), .B2(\mem[12][2] ), 
        .ZN(n1090) );
  INV_X1 U284 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U285 ( .A1(data_in[3]), .A2(n840), .B1(n1092), .B2(\mem[12][3] ), 
        .ZN(n1089) );
  INV_X1 U286 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U287 ( .A1(data_in[4]), .A2(n840), .B1(n1092), .B2(\mem[12][4] ), 
        .ZN(n1088) );
  INV_X1 U288 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U289 ( .A1(data_in[5]), .A2(n840), .B1(n1092), .B2(\mem[12][5] ), 
        .ZN(n1087) );
  INV_X1 U290 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U291 ( .A1(data_in[6]), .A2(n840), .B1(n1092), .B2(\mem[12][6] ), 
        .ZN(n1086) );
  INV_X1 U292 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U293 ( .A1(data_in[7]), .A2(n840), .B1(n1092), .B2(\mem[12][7] ), 
        .ZN(n1085) );
  INV_X1 U294 ( .A(n1084), .ZN(n780) );
  AOI22_X1 U295 ( .A1(data_in[0]), .A2(n839), .B1(n1083), .B2(\mem[13][0] ), 
        .ZN(n1084) );
  INV_X1 U296 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U297 ( .A1(data_in[1]), .A2(n839), .B1(n1083), .B2(\mem[13][1] ), 
        .ZN(n1082) );
  INV_X1 U298 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U299 ( .A1(data_in[2]), .A2(n839), .B1(n1083), .B2(\mem[13][2] ), 
        .ZN(n1081) );
  INV_X1 U300 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U301 ( .A1(data_in[3]), .A2(n839), .B1(n1083), .B2(\mem[13][3] ), 
        .ZN(n1080) );
  INV_X1 U302 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U303 ( .A1(data_in[4]), .A2(n839), .B1(n1083), .B2(\mem[13][4] ), 
        .ZN(n1079) );
  INV_X1 U304 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U305 ( .A1(data_in[5]), .A2(n839), .B1(n1083), .B2(\mem[13][5] ), 
        .ZN(n1078) );
  INV_X1 U306 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U307 ( .A1(data_in[6]), .A2(n839), .B1(n1083), .B2(\mem[13][6] ), 
        .ZN(n1077) );
  INV_X1 U308 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U309 ( .A1(data_in[7]), .A2(n839), .B1(n1083), .B2(\mem[13][7] ), 
        .ZN(n1076) );
  INV_X1 U310 ( .A(n1075), .ZN(n772) );
  AOI22_X1 U311 ( .A1(data_in[0]), .A2(n838), .B1(n1074), .B2(\mem[14][0] ), 
        .ZN(n1075) );
  INV_X1 U312 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U313 ( .A1(data_in[1]), .A2(n838), .B1(n1074), .B2(\mem[14][1] ), 
        .ZN(n1073) );
  INV_X1 U314 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U315 ( .A1(data_in[2]), .A2(n838), .B1(n1074), .B2(\mem[14][2] ), 
        .ZN(n1072) );
  INV_X1 U316 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U317 ( .A1(data_in[3]), .A2(n838), .B1(n1074), .B2(\mem[14][3] ), 
        .ZN(n1071) );
  INV_X1 U318 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U319 ( .A1(data_in[4]), .A2(n838), .B1(n1074), .B2(\mem[14][4] ), 
        .ZN(n1070) );
  INV_X1 U320 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U321 ( .A1(data_in[5]), .A2(n838), .B1(n1074), .B2(\mem[14][5] ), 
        .ZN(n1069) );
  INV_X1 U322 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U323 ( .A1(data_in[6]), .A2(n838), .B1(n1074), .B2(\mem[14][6] ), 
        .ZN(n1068) );
  INV_X1 U324 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U325 ( .A1(data_in[7]), .A2(n838), .B1(n1074), .B2(\mem[14][7] ), 
        .ZN(n1067) );
  INV_X1 U326 ( .A(n1066), .ZN(n764) );
  AOI22_X1 U327 ( .A1(data_in[0]), .A2(n837), .B1(n1065), .B2(\mem[15][0] ), 
        .ZN(n1066) );
  INV_X1 U328 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U329 ( .A1(data_in[1]), .A2(n837), .B1(n1065), .B2(\mem[15][1] ), 
        .ZN(n1064) );
  INV_X1 U330 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U331 ( .A1(data_in[2]), .A2(n837), .B1(n1065), .B2(\mem[15][2] ), 
        .ZN(n1063) );
  INV_X1 U332 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U333 ( .A1(data_in[3]), .A2(n837), .B1(n1065), .B2(\mem[15][3] ), 
        .ZN(n1062) );
  INV_X1 U334 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U335 ( .A1(data_in[4]), .A2(n837), .B1(n1065), .B2(\mem[15][4] ), 
        .ZN(n1061) );
  INV_X1 U336 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U337 ( .A1(data_in[5]), .A2(n837), .B1(n1065), .B2(\mem[15][5] ), 
        .ZN(n1060) );
  INV_X1 U338 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U339 ( .A1(data_in[6]), .A2(n837), .B1(n1065), .B2(\mem[15][6] ), 
        .ZN(n1059) );
  INV_X1 U340 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U341 ( .A1(data_in[7]), .A2(n837), .B1(n1065), .B2(\mem[15][7] ), 
        .ZN(n1058) );
  INV_X1 U342 ( .A(n1057), .ZN(n756) );
  AOI22_X1 U343 ( .A1(data_in[0]), .A2(n836), .B1(n1056), .B2(\mem[16][0] ), 
        .ZN(n1057) );
  INV_X1 U344 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U345 ( .A1(data_in[1]), .A2(n836), .B1(n1056), .B2(\mem[16][1] ), 
        .ZN(n1055) );
  INV_X1 U346 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U347 ( .A1(data_in[2]), .A2(n836), .B1(n1056), .B2(\mem[16][2] ), 
        .ZN(n1054) );
  INV_X1 U348 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U349 ( .A1(data_in[3]), .A2(n836), .B1(n1056), .B2(\mem[16][3] ), 
        .ZN(n1053) );
  INV_X1 U350 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U351 ( .A1(data_in[4]), .A2(n836), .B1(n1056), .B2(\mem[16][4] ), 
        .ZN(n1052) );
  INV_X1 U352 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U353 ( .A1(data_in[5]), .A2(n836), .B1(n1056), .B2(\mem[16][5] ), 
        .ZN(n1051) );
  INV_X1 U354 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U355 ( .A1(data_in[6]), .A2(n836), .B1(n1056), .B2(\mem[16][6] ), 
        .ZN(n1050) );
  INV_X1 U356 ( .A(n1049), .ZN(n749) );
  AOI22_X1 U357 ( .A1(data_in[7]), .A2(n836), .B1(n1056), .B2(\mem[16][7] ), 
        .ZN(n1049) );
  INV_X1 U358 ( .A(n1047), .ZN(n748) );
  AOI22_X1 U359 ( .A1(data_in[0]), .A2(n835), .B1(n1046), .B2(\mem[17][0] ), 
        .ZN(n1047) );
  INV_X1 U360 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U361 ( .A1(data_in[1]), .A2(n835), .B1(n1046), .B2(\mem[17][1] ), 
        .ZN(n1045) );
  INV_X1 U362 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U363 ( .A1(data_in[2]), .A2(n835), .B1(n1046), .B2(\mem[17][2] ), 
        .ZN(n1044) );
  INV_X1 U364 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[3]), .A2(n835), .B1(n1046), .B2(\mem[17][3] ), 
        .ZN(n1043) );
  INV_X1 U366 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[4]), .A2(n835), .B1(n1046), .B2(\mem[17][4] ), 
        .ZN(n1042) );
  INV_X1 U368 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[5]), .A2(n835), .B1(n1046), .B2(\mem[17][5] ), 
        .ZN(n1041) );
  INV_X1 U370 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[6]), .A2(n835), .B1(n1046), .B2(\mem[17][6] ), 
        .ZN(n1040) );
  INV_X1 U372 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[7]), .A2(n835), .B1(n1046), .B2(\mem[17][7] ), 
        .ZN(n1039) );
  INV_X1 U374 ( .A(n1038), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[0]), .A2(n834), .B1(n1037), .B2(\mem[18][0] ), 
        .ZN(n1038) );
  INV_X1 U376 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[1]), .A2(n834), .B1(n1037), .B2(\mem[18][1] ), 
        .ZN(n1036) );
  INV_X1 U378 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[2]), .A2(n834), .B1(n1037), .B2(\mem[18][2] ), 
        .ZN(n1035) );
  INV_X1 U380 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U381 ( .A1(data_in[3]), .A2(n834), .B1(n1037), .B2(\mem[18][3] ), 
        .ZN(n1034) );
  INV_X1 U382 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U383 ( .A1(data_in[4]), .A2(n834), .B1(n1037), .B2(\mem[18][4] ), 
        .ZN(n1033) );
  INV_X1 U384 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U385 ( .A1(data_in[5]), .A2(n834), .B1(n1037), .B2(\mem[18][5] ), 
        .ZN(n1032) );
  INV_X1 U386 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U387 ( .A1(data_in[6]), .A2(n834), .B1(n1037), .B2(\mem[18][6] ), 
        .ZN(n1031) );
  INV_X1 U388 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U389 ( .A1(data_in[7]), .A2(n834), .B1(n1037), .B2(\mem[18][7] ), 
        .ZN(n1030) );
  INV_X1 U390 ( .A(n1029), .ZN(n732) );
  AOI22_X1 U391 ( .A1(data_in[0]), .A2(n833), .B1(n1028), .B2(\mem[19][0] ), 
        .ZN(n1029) );
  INV_X1 U392 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U393 ( .A1(data_in[1]), .A2(n833), .B1(n1028), .B2(\mem[19][1] ), 
        .ZN(n1027) );
  INV_X1 U394 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U395 ( .A1(data_in[2]), .A2(n833), .B1(n1028), .B2(\mem[19][2] ), 
        .ZN(n1026) );
  INV_X1 U396 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U397 ( .A1(data_in[3]), .A2(n833), .B1(n1028), .B2(\mem[19][3] ), 
        .ZN(n1025) );
  INV_X1 U398 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U399 ( .A1(data_in[4]), .A2(n833), .B1(n1028), .B2(\mem[19][4] ), 
        .ZN(n1024) );
  INV_X1 U400 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U401 ( .A1(data_in[5]), .A2(n833), .B1(n1028), .B2(\mem[19][5] ), 
        .ZN(n1023) );
  INV_X1 U402 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U403 ( .A1(data_in[6]), .A2(n833), .B1(n1028), .B2(\mem[19][6] ), 
        .ZN(n1022) );
  INV_X1 U404 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U405 ( .A1(data_in[7]), .A2(n833), .B1(n1028), .B2(\mem[19][7] ), 
        .ZN(n1021) );
  INV_X1 U406 ( .A(n1020), .ZN(n724) );
  AOI22_X1 U407 ( .A1(data_in[0]), .A2(n832), .B1(n1019), .B2(\mem[20][0] ), 
        .ZN(n1020) );
  INV_X1 U408 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U409 ( .A1(data_in[1]), .A2(n832), .B1(n1019), .B2(\mem[20][1] ), 
        .ZN(n1018) );
  INV_X1 U410 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U411 ( .A1(data_in[2]), .A2(n832), .B1(n1019), .B2(\mem[20][2] ), 
        .ZN(n1017) );
  INV_X1 U412 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U413 ( .A1(data_in[3]), .A2(n832), .B1(n1019), .B2(\mem[20][3] ), 
        .ZN(n1016) );
  INV_X1 U414 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U415 ( .A1(data_in[4]), .A2(n832), .B1(n1019), .B2(\mem[20][4] ), 
        .ZN(n1015) );
  INV_X1 U416 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U417 ( .A1(data_in[5]), .A2(n832), .B1(n1019), .B2(\mem[20][5] ), 
        .ZN(n1014) );
  INV_X1 U418 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U419 ( .A1(data_in[6]), .A2(n832), .B1(n1019), .B2(\mem[20][6] ), 
        .ZN(n1013) );
  INV_X1 U420 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U421 ( .A1(data_in[7]), .A2(n832), .B1(n1019), .B2(\mem[20][7] ), 
        .ZN(n1012) );
  INV_X1 U422 ( .A(n1011), .ZN(n716) );
  AOI22_X1 U423 ( .A1(data_in[0]), .A2(n831), .B1(n1010), .B2(\mem[21][0] ), 
        .ZN(n1011) );
  INV_X1 U424 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U425 ( .A1(data_in[1]), .A2(n831), .B1(n1010), .B2(\mem[21][1] ), 
        .ZN(n1009) );
  INV_X1 U426 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U427 ( .A1(data_in[2]), .A2(n831), .B1(n1010), .B2(\mem[21][2] ), 
        .ZN(n1008) );
  INV_X1 U428 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U429 ( .A1(data_in[3]), .A2(n831), .B1(n1010), .B2(\mem[21][3] ), 
        .ZN(n1007) );
  INV_X1 U430 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U431 ( .A1(data_in[4]), .A2(n831), .B1(n1010), .B2(\mem[21][4] ), 
        .ZN(n1006) );
  INV_X1 U432 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U433 ( .A1(data_in[5]), .A2(n831), .B1(n1010), .B2(\mem[21][5] ), 
        .ZN(n1005) );
  INV_X1 U434 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U435 ( .A1(data_in[6]), .A2(n831), .B1(n1010), .B2(\mem[21][6] ), 
        .ZN(n1004) );
  INV_X1 U436 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U437 ( .A1(data_in[7]), .A2(n831), .B1(n1010), .B2(\mem[21][7] ), 
        .ZN(n1003) );
  INV_X1 U438 ( .A(n1002), .ZN(n708) );
  AOI22_X1 U439 ( .A1(data_in[0]), .A2(n830), .B1(n1001), .B2(\mem[22][0] ), 
        .ZN(n1002) );
  INV_X1 U440 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U441 ( .A1(data_in[1]), .A2(n830), .B1(n1001), .B2(\mem[22][1] ), 
        .ZN(n1000) );
  INV_X1 U442 ( .A(n999), .ZN(n706) );
  AOI22_X1 U443 ( .A1(data_in[2]), .A2(n830), .B1(n1001), .B2(\mem[22][2] ), 
        .ZN(n999) );
  INV_X1 U444 ( .A(n998), .ZN(n705) );
  AOI22_X1 U445 ( .A1(data_in[3]), .A2(n830), .B1(n1001), .B2(\mem[22][3] ), 
        .ZN(n998) );
  INV_X1 U446 ( .A(n997), .ZN(n704) );
  AOI22_X1 U447 ( .A1(data_in[4]), .A2(n830), .B1(n1001), .B2(\mem[22][4] ), 
        .ZN(n997) );
  INV_X1 U448 ( .A(n996), .ZN(n703) );
  AOI22_X1 U449 ( .A1(data_in[5]), .A2(n830), .B1(n1001), .B2(\mem[22][5] ), 
        .ZN(n996) );
  INV_X1 U450 ( .A(n995), .ZN(n702) );
  AOI22_X1 U451 ( .A1(data_in[6]), .A2(n830), .B1(n1001), .B2(\mem[22][6] ), 
        .ZN(n995) );
  INV_X1 U452 ( .A(n994), .ZN(n701) );
  AOI22_X1 U453 ( .A1(data_in[7]), .A2(n830), .B1(n1001), .B2(\mem[22][7] ), 
        .ZN(n994) );
  INV_X1 U454 ( .A(n993), .ZN(n700) );
  AOI22_X1 U455 ( .A1(data_in[0]), .A2(n829), .B1(n992), .B2(\mem[23][0] ), 
        .ZN(n993) );
  INV_X1 U456 ( .A(n991), .ZN(n699) );
  AOI22_X1 U457 ( .A1(data_in[1]), .A2(n829), .B1(n992), .B2(\mem[23][1] ), 
        .ZN(n991) );
  INV_X1 U458 ( .A(n990), .ZN(n698) );
  AOI22_X1 U459 ( .A1(data_in[2]), .A2(n829), .B1(n992), .B2(\mem[23][2] ), 
        .ZN(n990) );
  INV_X1 U460 ( .A(n989), .ZN(n697) );
  AOI22_X1 U461 ( .A1(data_in[3]), .A2(n829), .B1(n992), .B2(\mem[23][3] ), 
        .ZN(n989) );
  INV_X1 U462 ( .A(n988), .ZN(n696) );
  AOI22_X1 U463 ( .A1(data_in[4]), .A2(n829), .B1(n992), .B2(\mem[23][4] ), 
        .ZN(n988) );
  INV_X1 U464 ( .A(n987), .ZN(n695) );
  AOI22_X1 U465 ( .A1(data_in[5]), .A2(n829), .B1(n992), .B2(\mem[23][5] ), 
        .ZN(n987) );
  INV_X1 U466 ( .A(n986), .ZN(n694) );
  AOI22_X1 U467 ( .A1(data_in[6]), .A2(n829), .B1(n992), .B2(\mem[23][6] ), 
        .ZN(n986) );
  INV_X1 U468 ( .A(n985), .ZN(n693) );
  AOI22_X1 U469 ( .A1(data_in[7]), .A2(n829), .B1(n992), .B2(\mem[23][7] ), 
        .ZN(n985) );
  INV_X1 U470 ( .A(n984), .ZN(n692) );
  AOI22_X1 U471 ( .A1(data_in[0]), .A2(n828), .B1(n983), .B2(\mem[24][0] ), 
        .ZN(n984) );
  INV_X1 U472 ( .A(n982), .ZN(n691) );
  AOI22_X1 U473 ( .A1(data_in[1]), .A2(n828), .B1(n983), .B2(\mem[24][1] ), 
        .ZN(n982) );
  INV_X1 U474 ( .A(n981), .ZN(n690) );
  AOI22_X1 U475 ( .A1(data_in[2]), .A2(n828), .B1(n983), .B2(\mem[24][2] ), 
        .ZN(n981) );
  INV_X1 U476 ( .A(n980), .ZN(n689) );
  AOI22_X1 U477 ( .A1(data_in[3]), .A2(n828), .B1(n983), .B2(\mem[24][3] ), 
        .ZN(n980) );
  INV_X1 U478 ( .A(n979), .ZN(n688) );
  AOI22_X1 U479 ( .A1(data_in[4]), .A2(n828), .B1(n983), .B2(\mem[24][4] ), 
        .ZN(n979) );
  INV_X1 U480 ( .A(n978), .ZN(n687) );
  AOI22_X1 U481 ( .A1(data_in[5]), .A2(n828), .B1(n983), .B2(\mem[24][5] ), 
        .ZN(n978) );
  INV_X1 U482 ( .A(n977), .ZN(n686) );
  AOI22_X1 U483 ( .A1(data_in[6]), .A2(n828), .B1(n983), .B2(\mem[24][6] ), 
        .ZN(n977) );
  INV_X1 U484 ( .A(n976), .ZN(n685) );
  AOI22_X1 U485 ( .A1(data_in[7]), .A2(n828), .B1(n983), .B2(\mem[24][7] ), 
        .ZN(n976) );
  INV_X1 U486 ( .A(n974), .ZN(n684) );
  AOI22_X1 U487 ( .A1(data_in[0]), .A2(n827), .B1(n973), .B2(\mem[25][0] ), 
        .ZN(n974) );
  INV_X1 U488 ( .A(n972), .ZN(n683) );
  AOI22_X1 U489 ( .A1(data_in[1]), .A2(n827), .B1(n973), .B2(\mem[25][1] ), 
        .ZN(n972) );
  INV_X1 U490 ( .A(n971), .ZN(n682) );
  AOI22_X1 U491 ( .A1(data_in[2]), .A2(n827), .B1(n973), .B2(\mem[25][2] ), 
        .ZN(n971) );
  INV_X1 U492 ( .A(n970), .ZN(n681) );
  AOI22_X1 U493 ( .A1(data_in[3]), .A2(n827), .B1(n973), .B2(\mem[25][3] ), 
        .ZN(n970) );
  INV_X1 U494 ( .A(n969), .ZN(n680) );
  AOI22_X1 U495 ( .A1(data_in[4]), .A2(n827), .B1(n973), .B2(\mem[25][4] ), 
        .ZN(n969) );
  INV_X1 U496 ( .A(n968), .ZN(n679) );
  AOI22_X1 U497 ( .A1(data_in[5]), .A2(n827), .B1(n973), .B2(\mem[25][5] ), 
        .ZN(n968) );
  INV_X1 U498 ( .A(n967), .ZN(n678) );
  AOI22_X1 U499 ( .A1(data_in[6]), .A2(n827), .B1(n973), .B2(\mem[25][6] ), 
        .ZN(n967) );
  INV_X1 U500 ( .A(n966), .ZN(n677) );
  AOI22_X1 U501 ( .A1(data_in[7]), .A2(n827), .B1(n973), .B2(\mem[25][7] ), 
        .ZN(n966) );
  INV_X1 U502 ( .A(n965), .ZN(n676) );
  AOI22_X1 U503 ( .A1(data_in[0]), .A2(n826), .B1(n964), .B2(\mem[26][0] ), 
        .ZN(n965) );
  INV_X1 U504 ( .A(n963), .ZN(n675) );
  AOI22_X1 U505 ( .A1(data_in[1]), .A2(n826), .B1(n964), .B2(\mem[26][1] ), 
        .ZN(n963) );
  INV_X1 U506 ( .A(n962), .ZN(n674) );
  AOI22_X1 U507 ( .A1(data_in[2]), .A2(n826), .B1(n964), .B2(\mem[26][2] ), 
        .ZN(n962) );
  INV_X1 U508 ( .A(n961), .ZN(n673) );
  AOI22_X1 U509 ( .A1(data_in[3]), .A2(n826), .B1(n964), .B2(\mem[26][3] ), 
        .ZN(n961) );
  INV_X1 U510 ( .A(n960), .ZN(n672) );
  AOI22_X1 U511 ( .A1(data_in[4]), .A2(n826), .B1(n964), .B2(\mem[26][4] ), 
        .ZN(n960) );
  INV_X1 U512 ( .A(n959), .ZN(n671) );
  AOI22_X1 U513 ( .A1(data_in[5]), .A2(n826), .B1(n964), .B2(\mem[26][5] ), 
        .ZN(n959) );
  INV_X1 U514 ( .A(n958), .ZN(n670) );
  AOI22_X1 U515 ( .A1(data_in[6]), .A2(n826), .B1(n964), .B2(\mem[26][6] ), 
        .ZN(n958) );
  INV_X1 U516 ( .A(n957), .ZN(n669) );
  AOI22_X1 U517 ( .A1(data_in[7]), .A2(n826), .B1(n964), .B2(\mem[26][7] ), 
        .ZN(n957) );
  INV_X1 U518 ( .A(n956), .ZN(n668) );
  AOI22_X1 U519 ( .A1(data_in[0]), .A2(n825), .B1(n955), .B2(\mem[27][0] ), 
        .ZN(n956) );
  INV_X1 U520 ( .A(n954), .ZN(n667) );
  AOI22_X1 U521 ( .A1(data_in[1]), .A2(n825), .B1(n955), .B2(\mem[27][1] ), 
        .ZN(n954) );
  INV_X1 U522 ( .A(n953), .ZN(n666) );
  AOI22_X1 U523 ( .A1(data_in[2]), .A2(n825), .B1(n955), .B2(\mem[27][2] ), 
        .ZN(n953) );
  INV_X1 U524 ( .A(n952), .ZN(n665) );
  AOI22_X1 U525 ( .A1(data_in[3]), .A2(n825), .B1(n955), .B2(\mem[27][3] ), 
        .ZN(n952) );
  INV_X1 U526 ( .A(n951), .ZN(n664) );
  AOI22_X1 U527 ( .A1(data_in[4]), .A2(n825), .B1(n955), .B2(\mem[27][4] ), 
        .ZN(n951) );
  INV_X1 U528 ( .A(n950), .ZN(n663) );
  AOI22_X1 U529 ( .A1(data_in[5]), .A2(n825), .B1(n955), .B2(\mem[27][5] ), 
        .ZN(n950) );
  INV_X1 U530 ( .A(n949), .ZN(n662) );
  AOI22_X1 U531 ( .A1(data_in[6]), .A2(n825), .B1(n955), .B2(\mem[27][6] ), 
        .ZN(n949) );
  INV_X1 U532 ( .A(n948), .ZN(n661) );
  AOI22_X1 U533 ( .A1(data_in[7]), .A2(n825), .B1(n955), .B2(\mem[27][7] ), 
        .ZN(n948) );
  INV_X1 U534 ( .A(n947), .ZN(n660) );
  AOI22_X1 U535 ( .A1(data_in[0]), .A2(n824), .B1(n946), .B2(\mem[28][0] ), 
        .ZN(n947) );
  INV_X1 U536 ( .A(n945), .ZN(n659) );
  AOI22_X1 U537 ( .A1(data_in[1]), .A2(n824), .B1(n946), .B2(\mem[28][1] ), 
        .ZN(n945) );
  INV_X1 U538 ( .A(n944), .ZN(n658) );
  AOI22_X1 U539 ( .A1(data_in[2]), .A2(n824), .B1(n946), .B2(\mem[28][2] ), 
        .ZN(n944) );
  INV_X1 U540 ( .A(n943), .ZN(n657) );
  AOI22_X1 U541 ( .A1(data_in[3]), .A2(n824), .B1(n946), .B2(\mem[28][3] ), 
        .ZN(n943) );
  INV_X1 U542 ( .A(n942), .ZN(n656) );
  AOI22_X1 U543 ( .A1(data_in[4]), .A2(n824), .B1(n946), .B2(\mem[28][4] ), 
        .ZN(n942) );
  INV_X1 U544 ( .A(n941), .ZN(n655) );
  AOI22_X1 U545 ( .A1(data_in[5]), .A2(n824), .B1(n946), .B2(\mem[28][5] ), 
        .ZN(n941) );
  INV_X1 U546 ( .A(n940), .ZN(n654) );
  AOI22_X1 U547 ( .A1(data_in[6]), .A2(n824), .B1(n946), .B2(\mem[28][6] ), 
        .ZN(n940) );
  INV_X1 U548 ( .A(n939), .ZN(n653) );
  AOI22_X1 U549 ( .A1(data_in[7]), .A2(n824), .B1(n946), .B2(\mem[28][7] ), 
        .ZN(n939) );
  INV_X1 U550 ( .A(n938), .ZN(n652) );
  AOI22_X1 U551 ( .A1(data_in[0]), .A2(n823), .B1(n937), .B2(\mem[29][0] ), 
        .ZN(n938) );
  INV_X1 U552 ( .A(n936), .ZN(n651) );
  AOI22_X1 U553 ( .A1(data_in[1]), .A2(n823), .B1(n937), .B2(\mem[29][1] ), 
        .ZN(n936) );
  INV_X1 U554 ( .A(n935), .ZN(n650) );
  AOI22_X1 U555 ( .A1(data_in[2]), .A2(n823), .B1(n937), .B2(\mem[29][2] ), 
        .ZN(n935) );
  INV_X1 U556 ( .A(n934), .ZN(n649) );
  AOI22_X1 U557 ( .A1(data_in[3]), .A2(n823), .B1(n937), .B2(\mem[29][3] ), 
        .ZN(n934) );
  INV_X1 U558 ( .A(n933), .ZN(n648) );
  AOI22_X1 U559 ( .A1(data_in[4]), .A2(n823), .B1(n937), .B2(\mem[29][4] ), 
        .ZN(n933) );
  INV_X1 U560 ( .A(n932), .ZN(n647) );
  AOI22_X1 U561 ( .A1(data_in[5]), .A2(n823), .B1(n937), .B2(\mem[29][5] ), 
        .ZN(n932) );
  INV_X1 U562 ( .A(n931), .ZN(n646) );
  AOI22_X1 U563 ( .A1(data_in[6]), .A2(n823), .B1(n937), .B2(\mem[29][6] ), 
        .ZN(n931) );
  INV_X1 U564 ( .A(n930), .ZN(n645) );
  AOI22_X1 U565 ( .A1(data_in[7]), .A2(n823), .B1(n937), .B2(\mem[29][7] ), 
        .ZN(n930) );
  INV_X1 U566 ( .A(n929), .ZN(n644) );
  AOI22_X1 U567 ( .A1(data_in[0]), .A2(n822), .B1(n928), .B2(\mem[30][0] ), 
        .ZN(n929) );
  INV_X1 U568 ( .A(n927), .ZN(n643) );
  AOI22_X1 U569 ( .A1(data_in[1]), .A2(n822), .B1(n928), .B2(\mem[30][1] ), 
        .ZN(n927) );
  INV_X1 U570 ( .A(n926), .ZN(n642) );
  AOI22_X1 U571 ( .A1(data_in[2]), .A2(n822), .B1(n928), .B2(\mem[30][2] ), 
        .ZN(n926) );
  INV_X1 U572 ( .A(n925), .ZN(n641) );
  AOI22_X1 U573 ( .A1(data_in[3]), .A2(n822), .B1(n928), .B2(\mem[30][3] ), 
        .ZN(n925) );
  INV_X1 U574 ( .A(n924), .ZN(n640) );
  AOI22_X1 U575 ( .A1(data_in[4]), .A2(n822), .B1(n928), .B2(\mem[30][4] ), 
        .ZN(n924) );
  INV_X1 U576 ( .A(n923), .ZN(n639) );
  AOI22_X1 U577 ( .A1(data_in[5]), .A2(n822), .B1(n928), .B2(\mem[30][5] ), 
        .ZN(n923) );
  INV_X1 U578 ( .A(n922), .ZN(n638) );
  AOI22_X1 U579 ( .A1(data_in[6]), .A2(n822), .B1(n928), .B2(\mem[30][6] ), 
        .ZN(n922) );
  INV_X1 U580 ( .A(n921), .ZN(n637) );
  AOI22_X1 U581 ( .A1(data_in[7]), .A2(n822), .B1(n928), .B2(\mem[30][7] ), 
        .ZN(n921) );
  INV_X1 U582 ( .A(n920), .ZN(n636) );
  AOI22_X1 U583 ( .A1(data_in[0]), .A2(n821), .B1(n919), .B2(\mem[31][0] ), 
        .ZN(n920) );
  INV_X1 U584 ( .A(n918), .ZN(n635) );
  AOI22_X1 U585 ( .A1(data_in[1]), .A2(n821), .B1(n919), .B2(\mem[31][1] ), 
        .ZN(n918) );
  INV_X1 U586 ( .A(n917), .ZN(n634) );
  AOI22_X1 U587 ( .A1(data_in[2]), .A2(n821), .B1(n919), .B2(\mem[31][2] ), 
        .ZN(n917) );
  INV_X1 U588 ( .A(n916), .ZN(n633) );
  AOI22_X1 U589 ( .A1(data_in[3]), .A2(n821), .B1(n919), .B2(\mem[31][3] ), 
        .ZN(n916) );
  INV_X1 U590 ( .A(n915), .ZN(n632) );
  AOI22_X1 U591 ( .A1(data_in[4]), .A2(n821), .B1(n919), .B2(\mem[31][4] ), 
        .ZN(n915) );
  INV_X1 U592 ( .A(n914), .ZN(n631) );
  AOI22_X1 U593 ( .A1(data_in[5]), .A2(n821), .B1(n919), .B2(\mem[31][5] ), 
        .ZN(n914) );
  INV_X1 U594 ( .A(n913), .ZN(n630) );
  AOI22_X1 U595 ( .A1(data_in[6]), .A2(n821), .B1(n919), .B2(\mem[31][6] ), 
        .ZN(n913) );
  INV_X1 U596 ( .A(n912), .ZN(n629) );
  AOI22_X1 U597 ( .A1(data_in[7]), .A2(n821), .B1(n919), .B2(\mem[31][7] ), 
        .ZN(n912) );
  MUX2_X1 U598 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n615), .Z(n3) );
  MUX2_X1 U599 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n615), .Z(n4) );
  MUX2_X1 U600 ( .A(n4), .B(n3), .S(n610), .Z(n5) );
  MUX2_X1 U601 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n615), .Z(n6) );
  MUX2_X1 U602 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n615), .Z(n7) );
  MUX2_X1 U603 ( .A(n7), .B(n6), .S(n610), .Z(n8) );
  MUX2_X1 U604 ( .A(n8), .B(n5), .S(n608), .Z(n9) );
  MUX2_X1 U605 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n615), .Z(n10) );
  MUX2_X1 U606 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n615), .Z(n11) );
  MUX2_X1 U607 ( .A(n11), .B(n10), .S(n610), .Z(n12) );
  MUX2_X1 U608 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n615), .Z(n13) );
  MUX2_X1 U609 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n615), .Z(n14) );
  MUX2_X1 U610 ( .A(n14), .B(n13), .S(n610), .Z(n15) );
  MUX2_X1 U611 ( .A(n15), .B(n12), .S(N12), .Z(n16) );
  MUX2_X1 U612 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U613 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n613), .Z(n18) );
  MUX2_X1 U614 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n617), .Z(n19) );
  MUX2_X1 U615 ( .A(n19), .B(n18), .S(n610), .Z(n20) );
  MUX2_X1 U616 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n617), .Z(n21) );
  MUX2_X1 U617 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n613), .Z(n22) );
  MUX2_X1 U618 ( .A(n22), .B(n21), .S(n611), .Z(n23) );
  MUX2_X1 U619 ( .A(n23), .B(n20), .S(N12), .Z(n24) );
  MUX2_X1 U620 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n614), .Z(n25) );
  MUX2_X1 U621 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n616), .Z(n26) );
  MUX2_X1 U622 ( .A(n26), .B(n25), .S(n610), .Z(n27) );
  MUX2_X1 U623 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n614), .Z(n28) );
  MUX2_X1 U624 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n616), .Z(n29) );
  MUX2_X1 U625 ( .A(n29), .B(n28), .S(N11), .Z(n30) );
  MUX2_X1 U626 ( .A(n30), .B(n27), .S(n609), .Z(n31) );
  MUX2_X1 U627 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U628 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U629 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n616), .Z(n33) );
  MUX2_X1 U630 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n614), .Z(n34) );
  MUX2_X1 U631 ( .A(n34), .B(n33), .S(n610), .Z(n35) );
  MUX2_X1 U632 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n617), .Z(n36) );
  MUX2_X1 U633 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n613), .Z(n37) );
  MUX2_X1 U634 ( .A(n37), .B(n36), .S(n610), .Z(n38) );
  MUX2_X1 U635 ( .A(n38), .B(n35), .S(n609), .Z(n39) );
  MUX2_X1 U636 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n613), .Z(n40) );
  MUX2_X1 U637 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n613), .Z(n41) );
  MUX2_X1 U638 ( .A(n41), .B(n40), .S(n610), .Z(n42) );
  MUX2_X1 U639 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n613), .Z(n43) );
  MUX2_X1 U640 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n613), .Z(n44) );
  MUX2_X1 U641 ( .A(n44), .B(n43), .S(n611), .Z(n45) );
  MUX2_X1 U642 ( .A(n45), .B(n42), .S(n608), .Z(n46) );
  MUX2_X1 U643 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U644 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n613), .Z(n48) );
  MUX2_X1 U645 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n613), .Z(n49) );
  MUX2_X1 U646 ( .A(n49), .B(n48), .S(n610), .Z(n50) );
  MUX2_X1 U647 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n613), .Z(n51) );
  MUX2_X1 U648 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n613), .Z(n52) );
  MUX2_X1 U649 ( .A(n52), .B(n51), .S(n612), .Z(n53) );
  MUX2_X1 U650 ( .A(n53), .B(n50), .S(N12), .Z(n54) );
  MUX2_X1 U651 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n613), .Z(n55) );
  MUX2_X1 U652 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n613), .Z(n56) );
  MUX2_X1 U653 ( .A(n56), .B(n55), .S(n610), .Z(n57) );
  MUX2_X1 U654 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n613), .Z(n58) );
  MUX2_X1 U655 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n613), .Z(n59) );
  MUX2_X1 U656 ( .A(n59), .B(n58), .S(n610), .Z(n60) );
  MUX2_X1 U657 ( .A(n60), .B(n57), .S(n608), .Z(n61) );
  MUX2_X1 U658 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U659 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U660 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n616), .Z(n63) );
  MUX2_X1 U661 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n613), .Z(n64) );
  MUX2_X1 U662 ( .A(n64), .B(n63), .S(n611), .Z(n65) );
  MUX2_X1 U663 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n618), .Z(n66) );
  MUX2_X1 U664 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n614), .Z(n67) );
  MUX2_X1 U665 ( .A(n67), .B(n66), .S(n611), .Z(n68) );
  MUX2_X1 U666 ( .A(n68), .B(n65), .S(n608), .Z(n69) );
  MUX2_X1 U667 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n614), .Z(n70) );
  MUX2_X1 U668 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n613), .Z(n71) );
  MUX2_X1 U669 ( .A(n71), .B(n70), .S(n611), .Z(n72) );
  MUX2_X1 U670 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n616), .Z(n73) );
  MUX2_X1 U671 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n616), .Z(n74) );
  MUX2_X1 U672 ( .A(n74), .B(n73), .S(n611), .Z(n75) );
  MUX2_X1 U673 ( .A(n75), .B(n72), .S(n608), .Z(n76) );
  MUX2_X1 U674 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U675 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n613), .Z(n78) );
  MUX2_X1 U676 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n616), .Z(n79) );
  MUX2_X1 U677 ( .A(n79), .B(n78), .S(n611), .Z(n80) );
  MUX2_X1 U678 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n617), .Z(n81) );
  MUX2_X1 U679 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n617), .Z(n82) );
  MUX2_X1 U680 ( .A(n82), .B(n81), .S(n611), .Z(n83) );
  MUX2_X1 U681 ( .A(n83), .B(n80), .S(n608), .Z(n84) );
  MUX2_X1 U682 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n618), .Z(n85) );
  MUX2_X1 U683 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n614), .Z(n86) );
  MUX2_X1 U684 ( .A(n86), .B(n85), .S(n611), .Z(n87) );
  MUX2_X1 U685 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n618), .Z(n88) );
  MUX2_X1 U686 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n617), .Z(n89) );
  MUX2_X1 U687 ( .A(n89), .B(n88), .S(n611), .Z(n90) );
  MUX2_X1 U688 ( .A(n90), .B(n87), .S(n608), .Z(n91) );
  MUX2_X1 U689 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U690 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U691 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n616), .Z(n93) );
  MUX2_X1 U692 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n618), .Z(n94) );
  MUX2_X1 U693 ( .A(n94), .B(n93), .S(n611), .Z(n95) );
  MUX2_X1 U694 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n618), .Z(n96) );
  MUX2_X1 U695 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n618), .Z(n97) );
  MUX2_X1 U696 ( .A(n97), .B(n96), .S(n611), .Z(n98) );
  MUX2_X1 U697 ( .A(n98), .B(n95), .S(n608), .Z(n99) );
  MUX2_X1 U698 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n618), .Z(n100) );
  MUX2_X1 U699 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n618), .Z(n101) );
  MUX2_X1 U700 ( .A(n101), .B(n100), .S(n611), .Z(n102) );
  MUX2_X1 U701 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n618), .Z(n103) );
  MUX2_X1 U702 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n617), .Z(n104) );
  MUX2_X1 U703 ( .A(n104), .B(n103), .S(n611), .Z(n105) );
  MUX2_X1 U704 ( .A(n105), .B(n102), .S(n608), .Z(n106) );
  MUX2_X1 U705 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U706 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n614), .Z(n108) );
  MUX2_X1 U707 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n614), .Z(n109) );
  MUX2_X1 U708 ( .A(n109), .B(n108), .S(n612), .Z(n110) );
  MUX2_X1 U709 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n614), .Z(n111) );
  MUX2_X1 U710 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n614), .Z(n112) );
  MUX2_X1 U711 ( .A(n112), .B(n111), .S(n612), .Z(n113) );
  MUX2_X1 U712 ( .A(n113), .B(n110), .S(n608), .Z(n114) );
  MUX2_X1 U713 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n614), .Z(n115) );
  MUX2_X1 U714 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n614), .Z(n116) );
  MUX2_X1 U715 ( .A(n116), .B(n115), .S(n612), .Z(n117) );
  MUX2_X1 U716 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n614), .Z(n118) );
  MUX2_X1 U717 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n614), .Z(n119) );
  MUX2_X1 U718 ( .A(n119), .B(n118), .S(n612), .Z(n120) );
  MUX2_X1 U719 ( .A(n120), .B(n117), .S(n608), .Z(n121) );
  MUX2_X1 U720 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U721 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U722 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n614), .Z(n123) );
  MUX2_X1 U723 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n614), .Z(n124) );
  MUX2_X1 U724 ( .A(n124), .B(n123), .S(n612), .Z(n125) );
  MUX2_X1 U725 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n614), .Z(n126) );
  MUX2_X1 U726 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n614), .Z(n127) );
  MUX2_X1 U727 ( .A(n127), .B(n126), .S(n612), .Z(n128) );
  MUX2_X1 U728 ( .A(n128), .B(n125), .S(n608), .Z(n129) );
  MUX2_X1 U729 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n615), .Z(n130) );
  MUX2_X1 U730 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n615), .Z(n131) );
  MUX2_X1 U731 ( .A(n131), .B(n130), .S(n612), .Z(n132) );
  MUX2_X1 U732 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n615), .Z(n133) );
  MUX2_X1 U733 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n615), .Z(n134) );
  MUX2_X1 U734 ( .A(n134), .B(n133), .S(n612), .Z(n135) );
  MUX2_X1 U735 ( .A(n135), .B(n132), .S(n608), .Z(n136) );
  MUX2_X1 U736 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U737 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n615), .Z(n138) );
  MUX2_X1 U738 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n615), .Z(n139) );
  MUX2_X1 U739 ( .A(n139), .B(n138), .S(n612), .Z(n140) );
  MUX2_X1 U740 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n615), .Z(n141) );
  MUX2_X1 U741 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n615), .Z(n142) );
  MUX2_X1 U742 ( .A(n142), .B(n141), .S(n612), .Z(n143) );
  MUX2_X1 U743 ( .A(n143), .B(n140), .S(n608), .Z(n144) );
  MUX2_X1 U744 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n615), .Z(n145) );
  MUX2_X1 U745 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n615), .Z(n146) );
  MUX2_X1 U746 ( .A(n146), .B(n145), .S(n612), .Z(n147) );
  MUX2_X1 U747 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n615), .Z(n148) );
  MUX2_X1 U748 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n615), .Z(n149) );
  MUX2_X1 U749 ( .A(n149), .B(n148), .S(n612), .Z(n150) );
  MUX2_X1 U750 ( .A(n150), .B(n147), .S(n608), .Z(n151) );
  MUX2_X1 U751 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U752 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U753 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n616), .Z(n153) );
  MUX2_X1 U754 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n616), .Z(n154) );
  MUX2_X1 U755 ( .A(n154), .B(n153), .S(n610), .Z(n155) );
  MUX2_X1 U756 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n616), .Z(n156) );
  MUX2_X1 U757 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n616), .Z(n157) );
  MUX2_X1 U758 ( .A(n157), .B(n156), .S(n612), .Z(n158) );
  MUX2_X1 U759 ( .A(n158), .B(n155), .S(n609), .Z(n159) );
  MUX2_X1 U760 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n616), .Z(n160) );
  MUX2_X1 U761 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n616), .Z(n161) );
  MUX2_X1 U762 ( .A(n161), .B(n160), .S(N11), .Z(n162) );
  MUX2_X1 U763 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n616), .Z(n163) );
  MUX2_X1 U764 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n616), .Z(n164) );
  MUX2_X1 U765 ( .A(n164), .B(n163), .S(n612), .Z(n165) );
  MUX2_X1 U766 ( .A(n165), .B(n162), .S(n609), .Z(n166) );
  MUX2_X1 U767 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U768 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n616), .Z(n168) );
  MUX2_X1 U769 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n616), .Z(n169) );
  MUX2_X1 U770 ( .A(n169), .B(n168), .S(n612), .Z(n170) );
  MUX2_X1 U771 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n616), .Z(n171) );
  MUX2_X1 U772 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n616), .Z(n172) );
  MUX2_X1 U773 ( .A(n172), .B(n171), .S(n610), .Z(n173) );
  MUX2_X1 U774 ( .A(n173), .B(n170), .S(n609), .Z(n174) );
  MUX2_X1 U775 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n618), .Z(n175) );
  MUX2_X1 U776 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n618), .Z(n176) );
  MUX2_X1 U777 ( .A(n176), .B(n175), .S(n611), .Z(n177) );
  MUX2_X1 U778 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n618), .Z(n178) );
  MUX2_X1 U779 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n179) );
  MUX2_X1 U780 ( .A(n179), .B(n178), .S(n611), .Z(n180) );
  MUX2_X1 U781 ( .A(n180), .B(n177), .S(n609), .Z(n181) );
  MUX2_X1 U782 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U783 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U784 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n614), .Z(n183) );
  MUX2_X1 U785 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n618), .Z(n184) );
  MUX2_X1 U786 ( .A(n184), .B(n183), .S(n611), .Z(n185) );
  MUX2_X1 U787 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n618), .Z(n186) );
  MUX2_X1 U788 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n613), .Z(n187) );
  MUX2_X1 U789 ( .A(n187), .B(n186), .S(n610), .Z(n188) );
  MUX2_X1 U790 ( .A(n188), .B(n185), .S(n609), .Z(n189) );
  MUX2_X1 U791 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n618), .Z(n190) );
  MUX2_X1 U792 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n618), .Z(n191) );
  MUX2_X1 U793 ( .A(n191), .B(n190), .S(n611), .Z(n192) );
  MUX2_X1 U794 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n613), .Z(n193) );
  MUX2_X1 U795 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n617), .Z(n194) );
  MUX2_X1 U796 ( .A(n194), .B(n193), .S(n610), .Z(n195) );
  MUX2_X1 U797 ( .A(n195), .B(n192), .S(n609), .Z(n196) );
  MUX2_X1 U798 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U799 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n614), .Z(n198) );
  MUX2_X1 U800 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n618), .Z(n199) );
  MUX2_X1 U801 ( .A(n199), .B(n198), .S(n612), .Z(n200) );
  MUX2_X1 U802 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n618), .Z(n201) );
  MUX2_X1 U803 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n202) );
  MUX2_X1 U804 ( .A(n202), .B(n201), .S(N11), .Z(n203) );
  MUX2_X1 U805 ( .A(n203), .B(n200), .S(n609), .Z(n204) );
  MUX2_X1 U806 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n618), .Z(n205) );
  MUX2_X1 U807 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n206) );
  MUX2_X1 U808 ( .A(n206), .B(n205), .S(n612), .Z(n207) );
  MUX2_X1 U809 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n208) );
  MUX2_X1 U810 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n209) );
  MUX2_X1 U811 ( .A(n209), .B(n208), .S(n611), .Z(n210) );
  MUX2_X1 U812 ( .A(n210), .B(n207), .S(n609), .Z(n211) );
  MUX2_X1 U813 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U814 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U815 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n615), .Z(n213) );
  MUX2_X1 U816 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n615), .Z(n214) );
  MUX2_X1 U817 ( .A(n214), .B(n213), .S(n611), .Z(n215) );
  MUX2_X1 U818 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n615), .Z(n216) );
  MUX2_X1 U819 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n618), .Z(n217) );
  MUX2_X1 U820 ( .A(n217), .B(n216), .S(n611), .Z(n218) );
  MUX2_X1 U821 ( .A(n218), .B(n215), .S(n609), .Z(n219) );
  MUX2_X1 U822 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n617), .Z(n220) );
  MUX2_X1 U823 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n617), .Z(n221) );
  MUX2_X1 U824 ( .A(n221), .B(n220), .S(n610), .Z(n222) );
  MUX2_X1 U825 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n617), .Z(n223) );
  MUX2_X1 U826 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n617), .Z(n224) );
  MUX2_X1 U827 ( .A(n224), .B(n223), .S(N11), .Z(n225) );
  MUX2_X1 U828 ( .A(n225), .B(n222), .S(n609), .Z(n226) );
  MUX2_X1 U829 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U830 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n617), .Z(n228) );
  MUX2_X1 U831 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n617), .Z(n229) );
  MUX2_X1 U832 ( .A(n229), .B(n228), .S(n610), .Z(n595) );
  MUX2_X1 U833 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n617), .Z(n596) );
  MUX2_X1 U834 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n617), .Z(n597) );
  MUX2_X1 U835 ( .A(n597), .B(n596), .S(N11), .Z(n598) );
  MUX2_X1 U836 ( .A(n598), .B(n595), .S(n609), .Z(n599) );
  MUX2_X1 U837 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n617), .Z(n600) );
  MUX2_X1 U838 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n617), .Z(n601) );
  MUX2_X1 U839 ( .A(n601), .B(n600), .S(n612), .Z(n602) );
  MUX2_X1 U840 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n617), .Z(n603) );
  MUX2_X1 U841 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n617), .Z(n604) );
  MUX2_X1 U842 ( .A(n604), .B(n603), .S(n612), .Z(n605) );
  MUX2_X1 U843 ( .A(n605), .B(n602), .S(n609), .Z(n606) );
  MUX2_X1 U844 ( .A(n606), .B(n599), .S(N13), .Z(n607) );
  MUX2_X1 U845 ( .A(n607), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U846 ( .A(N11), .Z(n610) );
  INV_X1 U847 ( .A(N10), .ZN(n619) );
  INV_X1 U848 ( .A(N11), .ZN(n620) );
  INV_X1 U849 ( .A(data_in[0]), .ZN(n621) );
  INV_X1 U850 ( .A(data_in[1]), .ZN(n622) );
  INV_X1 U851 ( .A(data_in[2]), .ZN(n623) );
  INV_X1 U852 ( .A(data_in[3]), .ZN(n624) );
  INV_X1 U853 ( .A(data_in[4]), .ZN(n625) );
  INV_X1 U854 ( .A(data_in[5]), .ZN(n626) );
  INV_X1 U855 ( .A(data_in[6]), .ZN(n627) );
  INV_X1 U856 ( .A(data_in[7]), .ZN(n628) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_20 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n629), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n630), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n631), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n632), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n633), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n634), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n635), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n636), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n637), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n638), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n639), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n640), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n641), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n642), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n643), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n644), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n645), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n646), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n647), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n648), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n649), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n650), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n651), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n652), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n653), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n654), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n655), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n656), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n657), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n658), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n659), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n660), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n661), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n662), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n663), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n664), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n665), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n666), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n667), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n668), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n669), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n670), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n671), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n672), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n673), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n674), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n675), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n676), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n677), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n678), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n679), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n680), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n681), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n682), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n683), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n684), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n685), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n686), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n687), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n688), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n689), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n690), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n691), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n692), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n693), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n694), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n695), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n696), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n697), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n698), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n699), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n700), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n701), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n702), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n703), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n704), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n705), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n706), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n707), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n708), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n709), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n710), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n711), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n712), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n713), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n714), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n715), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n716), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n717), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n718), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n719), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n720), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n721), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n722), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n723), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n724), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n725), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n726), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n727), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n728), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n729), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n730), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n731), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n732), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n733), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n734), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n735), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n736), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n737), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n738), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n739), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n740), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n741), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n742), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n743), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n744), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n745), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n746), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n747), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n748), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n749), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n750), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n751), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n752), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n753), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n754), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n755), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n756), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n757), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n758), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n759), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n760), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n761), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n762), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n763), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n764), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n765), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n766), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n767), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n768), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n769), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n770), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n771), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n772), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n773), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n774), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n775), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n776), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n777), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n778), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n779), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n780), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n781), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n782), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n783), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n784), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n785), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n786), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n787), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n788), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n789), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n790), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n791), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n792), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n793), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n794), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n795), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n796), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n797), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n798), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n799), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n800), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n801), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n802), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n803), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n804), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n805), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n806), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n807), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n808), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n809), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n810), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n811), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n812), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n813), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n814), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n815), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n816), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n817), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n818), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n819), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n820), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n848), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n849), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n850), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n851), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n852), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n853), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n854), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n855), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n856), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n857), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n858), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n859), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n860), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n861), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n862), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n863), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n864), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n865), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n866), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n867), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n868), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n869), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n870), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n871), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n872), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n873), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n874), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n875), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n876), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n877), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n878), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n879), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n880), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n881), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n882), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n883), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n884), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n885), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n886), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n887), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n888), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n889), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n890), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n891), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n892), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n893), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n894), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n895), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n896), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n897), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n898), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n899), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n900), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n901), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n902), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n903), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n904), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n905), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n906), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n907), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n908), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n909), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n910), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n911), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[5]) );
  BUF_X1 U4 ( .A(n618), .Z(n616) );
  BUF_X1 U5 ( .A(n618), .Z(n617) );
  BUF_X1 U6 ( .A(N10), .Z(n613) );
  BUF_X1 U7 ( .A(n618), .Z(n614) );
  BUF_X1 U8 ( .A(n618), .Z(n615) );
  BUF_X1 U9 ( .A(N11), .Z(n611) );
  BUF_X1 U10 ( .A(N11), .Z(n612) );
  BUF_X1 U11 ( .A(N10), .Z(n618) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1203) );
  NOR3_X1 U13 ( .A1(N11), .A2(N12), .A3(n619), .ZN(n1192) );
  NOR3_X1 U14 ( .A1(N10), .A2(N12), .A3(n620), .ZN(n1182) );
  NOR3_X1 U15 ( .A1(n619), .A2(N12), .A3(n620), .ZN(n1172) );
  INV_X1 U16 ( .A(n1129), .ZN(n844) );
  INV_X1 U17 ( .A(n1119), .ZN(n843) );
  INV_X1 U18 ( .A(n1110), .ZN(n842) );
  INV_X1 U19 ( .A(n1101), .ZN(n841) );
  INV_X1 U20 ( .A(n1056), .ZN(n836) );
  INV_X1 U21 ( .A(n1046), .ZN(n835) );
  INV_X1 U22 ( .A(n1037), .ZN(n834) );
  INV_X1 U23 ( .A(n1028), .ZN(n833) );
  INV_X1 U24 ( .A(n983), .ZN(n828) );
  INV_X1 U25 ( .A(n973), .ZN(n827) );
  INV_X1 U26 ( .A(n964), .ZN(n826) );
  INV_X1 U27 ( .A(n955), .ZN(n825) );
  INV_X1 U28 ( .A(n1092), .ZN(n840) );
  INV_X1 U29 ( .A(n1083), .ZN(n839) );
  INV_X1 U30 ( .A(n1074), .ZN(n838) );
  INV_X1 U31 ( .A(n1065), .ZN(n837) );
  INV_X1 U32 ( .A(n946), .ZN(n824) );
  INV_X1 U33 ( .A(n937), .ZN(n823) );
  INV_X1 U34 ( .A(n928), .ZN(n822) );
  INV_X1 U35 ( .A(n919), .ZN(n821) );
  INV_X1 U36 ( .A(n1019), .ZN(n832) );
  INV_X1 U37 ( .A(n1010), .ZN(n831) );
  INV_X1 U38 ( .A(n1001), .ZN(n830) );
  INV_X1 U39 ( .A(n992), .ZN(n829) );
  BUF_X1 U40 ( .A(N12), .Z(n609) );
  INV_X1 U41 ( .A(N13), .ZN(n846) );
  AND3_X1 U42 ( .A1(n619), .A2(n620), .A3(N12), .ZN(n1162) );
  AND3_X1 U43 ( .A1(N10), .A2(n620), .A3(N12), .ZN(n1152) );
  AND3_X1 U44 ( .A1(N11), .A2(n619), .A3(N12), .ZN(n1142) );
  AND3_X1 U45 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1132) );
  BUF_X1 U46 ( .A(N12), .Z(n608) );
  INV_X1 U47 ( .A(N14), .ZN(n847) );
  NAND2_X1 U48 ( .A1(n1192), .A2(n1202), .ZN(n1201) );
  NAND2_X1 U49 ( .A1(n1182), .A2(n1202), .ZN(n1191) );
  NAND2_X1 U50 ( .A1(n1172), .A2(n1202), .ZN(n1181) );
  NAND2_X1 U51 ( .A1(n1162), .A2(n1202), .ZN(n1171) );
  NAND2_X1 U52 ( .A1(n1152), .A2(n1202), .ZN(n1161) );
  NAND2_X1 U53 ( .A1(n1142), .A2(n1202), .ZN(n1151) );
  NAND2_X1 U54 ( .A1(n1132), .A2(n1202), .ZN(n1141) );
  NAND2_X1 U55 ( .A1(n1203), .A2(n1202), .ZN(n1212) );
  NAND2_X1 U56 ( .A1(n1121), .A2(n1203), .ZN(n1129) );
  NAND2_X1 U57 ( .A1(n1121), .A2(n1192), .ZN(n1119) );
  NAND2_X1 U58 ( .A1(n1121), .A2(n1182), .ZN(n1110) );
  NAND2_X1 U59 ( .A1(n1121), .A2(n1172), .ZN(n1101) );
  NAND2_X1 U60 ( .A1(n1048), .A2(n1203), .ZN(n1056) );
  NAND2_X1 U61 ( .A1(n1048), .A2(n1192), .ZN(n1046) );
  NAND2_X1 U62 ( .A1(n1048), .A2(n1182), .ZN(n1037) );
  NAND2_X1 U63 ( .A1(n1048), .A2(n1172), .ZN(n1028) );
  NAND2_X1 U64 ( .A1(n975), .A2(n1203), .ZN(n983) );
  NAND2_X1 U65 ( .A1(n975), .A2(n1192), .ZN(n973) );
  NAND2_X1 U66 ( .A1(n975), .A2(n1182), .ZN(n964) );
  NAND2_X1 U67 ( .A1(n975), .A2(n1172), .ZN(n955) );
  NAND2_X1 U68 ( .A1(n1121), .A2(n1162), .ZN(n1092) );
  NAND2_X1 U69 ( .A1(n1121), .A2(n1152), .ZN(n1083) );
  NAND2_X1 U70 ( .A1(n1121), .A2(n1142), .ZN(n1074) );
  NAND2_X1 U71 ( .A1(n1121), .A2(n1132), .ZN(n1065) );
  NAND2_X1 U72 ( .A1(n1048), .A2(n1162), .ZN(n1019) );
  NAND2_X1 U73 ( .A1(n1048), .A2(n1152), .ZN(n1010) );
  NAND2_X1 U74 ( .A1(n1048), .A2(n1142), .ZN(n1001) );
  NAND2_X1 U75 ( .A1(n1048), .A2(n1132), .ZN(n992) );
  NAND2_X1 U76 ( .A1(n975), .A2(n1162), .ZN(n946) );
  NAND2_X1 U77 ( .A1(n975), .A2(n1152), .ZN(n937) );
  NAND2_X1 U78 ( .A1(n975), .A2(n1142), .ZN(n928) );
  NAND2_X1 U79 ( .A1(n975), .A2(n1132), .ZN(n919) );
  AND3_X1 U80 ( .A1(n846), .A2(n847), .A3(n1131), .ZN(n1202) );
  AND3_X1 U81 ( .A1(N13), .A2(n1131), .A3(N14), .ZN(n975) );
  AND3_X1 U82 ( .A1(n1131), .A2(n847), .A3(N13), .ZN(n1121) );
  AND3_X1 U83 ( .A1(n1131), .A2(n846), .A3(N14), .ZN(n1048) );
  NOR2_X1 U84 ( .A1(n845), .A2(addr[5]), .ZN(n1131) );
  INV_X1 U85 ( .A(wr_en), .ZN(n845) );
  OAI21_X1 U86 ( .B1(n621), .B2(n1171), .A(n1170), .ZN(n879) );
  NAND2_X1 U87 ( .A1(\mem[4][0] ), .A2(n1171), .ZN(n1170) );
  OAI21_X1 U88 ( .B1(n622), .B2(n1171), .A(n1169), .ZN(n878) );
  NAND2_X1 U89 ( .A1(\mem[4][1] ), .A2(n1171), .ZN(n1169) );
  OAI21_X1 U90 ( .B1(n623), .B2(n1171), .A(n1168), .ZN(n877) );
  NAND2_X1 U91 ( .A1(\mem[4][2] ), .A2(n1171), .ZN(n1168) );
  OAI21_X1 U92 ( .B1(n624), .B2(n1171), .A(n1167), .ZN(n876) );
  NAND2_X1 U93 ( .A1(\mem[4][3] ), .A2(n1171), .ZN(n1167) );
  OAI21_X1 U94 ( .B1(n625), .B2(n1171), .A(n1166), .ZN(n875) );
  NAND2_X1 U95 ( .A1(\mem[4][4] ), .A2(n1171), .ZN(n1166) );
  OAI21_X1 U96 ( .B1(n626), .B2(n1171), .A(n1165), .ZN(n874) );
  NAND2_X1 U97 ( .A1(\mem[4][5] ), .A2(n1171), .ZN(n1165) );
  OAI21_X1 U98 ( .B1(n627), .B2(n1171), .A(n1164), .ZN(n873) );
  NAND2_X1 U99 ( .A1(\mem[4][6] ), .A2(n1171), .ZN(n1164) );
  OAI21_X1 U100 ( .B1(n628), .B2(n1171), .A(n1163), .ZN(n872) );
  NAND2_X1 U101 ( .A1(\mem[4][7] ), .A2(n1171), .ZN(n1163) );
  OAI21_X1 U102 ( .B1(n621), .B2(n1151), .A(n1150), .ZN(n863) );
  NAND2_X1 U103 ( .A1(\mem[6][0] ), .A2(n1151), .ZN(n1150) );
  OAI21_X1 U104 ( .B1(n622), .B2(n1151), .A(n1149), .ZN(n862) );
  NAND2_X1 U105 ( .A1(\mem[6][1] ), .A2(n1151), .ZN(n1149) );
  OAI21_X1 U106 ( .B1(n623), .B2(n1151), .A(n1148), .ZN(n861) );
  NAND2_X1 U107 ( .A1(\mem[6][2] ), .A2(n1151), .ZN(n1148) );
  OAI21_X1 U108 ( .B1(n624), .B2(n1151), .A(n1147), .ZN(n860) );
  NAND2_X1 U109 ( .A1(\mem[6][3] ), .A2(n1151), .ZN(n1147) );
  OAI21_X1 U110 ( .B1(n625), .B2(n1151), .A(n1146), .ZN(n859) );
  NAND2_X1 U111 ( .A1(\mem[6][4] ), .A2(n1151), .ZN(n1146) );
  OAI21_X1 U112 ( .B1(n626), .B2(n1151), .A(n1145), .ZN(n858) );
  NAND2_X1 U113 ( .A1(\mem[6][5] ), .A2(n1151), .ZN(n1145) );
  OAI21_X1 U114 ( .B1(n627), .B2(n1151), .A(n1144), .ZN(n857) );
  NAND2_X1 U115 ( .A1(\mem[6][6] ), .A2(n1151), .ZN(n1144) );
  OAI21_X1 U116 ( .B1(n628), .B2(n1151), .A(n1143), .ZN(n856) );
  NAND2_X1 U117 ( .A1(\mem[6][7] ), .A2(n1151), .ZN(n1143) );
  OAI21_X1 U118 ( .B1(n621), .B2(n1141), .A(n1140), .ZN(n855) );
  NAND2_X1 U119 ( .A1(\mem[7][0] ), .A2(n1141), .ZN(n1140) );
  OAI21_X1 U120 ( .B1(n622), .B2(n1141), .A(n1139), .ZN(n854) );
  NAND2_X1 U121 ( .A1(\mem[7][1] ), .A2(n1141), .ZN(n1139) );
  OAI21_X1 U122 ( .B1(n623), .B2(n1141), .A(n1138), .ZN(n853) );
  NAND2_X1 U123 ( .A1(\mem[7][2] ), .A2(n1141), .ZN(n1138) );
  OAI21_X1 U124 ( .B1(n624), .B2(n1141), .A(n1137), .ZN(n852) );
  NAND2_X1 U125 ( .A1(\mem[7][3] ), .A2(n1141), .ZN(n1137) );
  OAI21_X1 U126 ( .B1(n625), .B2(n1141), .A(n1136), .ZN(n851) );
  NAND2_X1 U127 ( .A1(\mem[7][4] ), .A2(n1141), .ZN(n1136) );
  OAI21_X1 U128 ( .B1(n626), .B2(n1141), .A(n1135), .ZN(n850) );
  NAND2_X1 U129 ( .A1(\mem[7][5] ), .A2(n1141), .ZN(n1135) );
  OAI21_X1 U130 ( .B1(n627), .B2(n1141), .A(n1134), .ZN(n849) );
  NAND2_X1 U131 ( .A1(\mem[7][6] ), .A2(n1141), .ZN(n1134) );
  OAI21_X1 U132 ( .B1(n628), .B2(n1141), .A(n1133), .ZN(n848) );
  NAND2_X1 U133 ( .A1(\mem[7][7] ), .A2(n1141), .ZN(n1133) );
  OAI21_X1 U134 ( .B1(n621), .B2(n1201), .A(n1200), .ZN(n903) );
  NAND2_X1 U135 ( .A1(\mem[1][0] ), .A2(n1201), .ZN(n1200) );
  OAI21_X1 U136 ( .B1(n622), .B2(n1201), .A(n1199), .ZN(n902) );
  NAND2_X1 U137 ( .A1(\mem[1][1] ), .A2(n1201), .ZN(n1199) );
  OAI21_X1 U138 ( .B1(n623), .B2(n1201), .A(n1198), .ZN(n901) );
  NAND2_X1 U139 ( .A1(\mem[1][2] ), .A2(n1201), .ZN(n1198) );
  OAI21_X1 U140 ( .B1(n624), .B2(n1201), .A(n1197), .ZN(n900) );
  NAND2_X1 U141 ( .A1(\mem[1][3] ), .A2(n1201), .ZN(n1197) );
  OAI21_X1 U142 ( .B1(n625), .B2(n1201), .A(n1196), .ZN(n899) );
  NAND2_X1 U143 ( .A1(\mem[1][4] ), .A2(n1201), .ZN(n1196) );
  OAI21_X1 U144 ( .B1(n626), .B2(n1201), .A(n1195), .ZN(n898) );
  NAND2_X1 U145 ( .A1(\mem[1][5] ), .A2(n1201), .ZN(n1195) );
  OAI21_X1 U146 ( .B1(n627), .B2(n1201), .A(n1194), .ZN(n897) );
  NAND2_X1 U147 ( .A1(\mem[1][6] ), .A2(n1201), .ZN(n1194) );
  OAI21_X1 U148 ( .B1(n628), .B2(n1201), .A(n1193), .ZN(n896) );
  NAND2_X1 U149 ( .A1(\mem[1][7] ), .A2(n1201), .ZN(n1193) );
  OAI21_X1 U150 ( .B1(n621), .B2(n1191), .A(n1190), .ZN(n895) );
  NAND2_X1 U151 ( .A1(\mem[2][0] ), .A2(n1191), .ZN(n1190) );
  OAI21_X1 U152 ( .B1(n622), .B2(n1191), .A(n1189), .ZN(n894) );
  NAND2_X1 U153 ( .A1(\mem[2][1] ), .A2(n1191), .ZN(n1189) );
  OAI21_X1 U154 ( .B1(n623), .B2(n1191), .A(n1188), .ZN(n893) );
  NAND2_X1 U155 ( .A1(\mem[2][2] ), .A2(n1191), .ZN(n1188) );
  OAI21_X1 U156 ( .B1(n624), .B2(n1191), .A(n1187), .ZN(n892) );
  NAND2_X1 U157 ( .A1(\mem[2][3] ), .A2(n1191), .ZN(n1187) );
  OAI21_X1 U158 ( .B1(n625), .B2(n1191), .A(n1186), .ZN(n891) );
  NAND2_X1 U159 ( .A1(\mem[2][4] ), .A2(n1191), .ZN(n1186) );
  OAI21_X1 U160 ( .B1(n626), .B2(n1191), .A(n1185), .ZN(n890) );
  NAND2_X1 U161 ( .A1(\mem[2][5] ), .A2(n1191), .ZN(n1185) );
  OAI21_X1 U162 ( .B1(n627), .B2(n1191), .A(n1184), .ZN(n889) );
  NAND2_X1 U163 ( .A1(\mem[2][6] ), .A2(n1191), .ZN(n1184) );
  OAI21_X1 U164 ( .B1(n628), .B2(n1191), .A(n1183), .ZN(n888) );
  NAND2_X1 U165 ( .A1(\mem[2][7] ), .A2(n1191), .ZN(n1183) );
  OAI21_X1 U166 ( .B1(n621), .B2(n1181), .A(n1180), .ZN(n887) );
  NAND2_X1 U167 ( .A1(\mem[3][0] ), .A2(n1181), .ZN(n1180) );
  OAI21_X1 U168 ( .B1(n622), .B2(n1181), .A(n1179), .ZN(n886) );
  NAND2_X1 U169 ( .A1(\mem[3][1] ), .A2(n1181), .ZN(n1179) );
  OAI21_X1 U170 ( .B1(n623), .B2(n1181), .A(n1178), .ZN(n885) );
  NAND2_X1 U171 ( .A1(\mem[3][2] ), .A2(n1181), .ZN(n1178) );
  OAI21_X1 U172 ( .B1(n624), .B2(n1181), .A(n1177), .ZN(n884) );
  NAND2_X1 U173 ( .A1(\mem[3][3] ), .A2(n1181), .ZN(n1177) );
  OAI21_X1 U174 ( .B1(n625), .B2(n1181), .A(n1176), .ZN(n883) );
  NAND2_X1 U175 ( .A1(\mem[3][4] ), .A2(n1181), .ZN(n1176) );
  OAI21_X1 U176 ( .B1(n626), .B2(n1181), .A(n1175), .ZN(n882) );
  NAND2_X1 U177 ( .A1(\mem[3][5] ), .A2(n1181), .ZN(n1175) );
  OAI21_X1 U178 ( .B1(n627), .B2(n1181), .A(n1174), .ZN(n881) );
  NAND2_X1 U179 ( .A1(\mem[3][6] ), .A2(n1181), .ZN(n1174) );
  OAI21_X1 U180 ( .B1(n628), .B2(n1181), .A(n1173), .ZN(n880) );
  NAND2_X1 U181 ( .A1(\mem[3][7] ), .A2(n1181), .ZN(n1173) );
  OAI21_X1 U182 ( .B1(n621), .B2(n1161), .A(n1160), .ZN(n871) );
  NAND2_X1 U183 ( .A1(\mem[5][0] ), .A2(n1161), .ZN(n1160) );
  OAI21_X1 U184 ( .B1(n622), .B2(n1161), .A(n1159), .ZN(n870) );
  NAND2_X1 U185 ( .A1(\mem[5][1] ), .A2(n1161), .ZN(n1159) );
  OAI21_X1 U186 ( .B1(n623), .B2(n1161), .A(n1158), .ZN(n869) );
  NAND2_X1 U187 ( .A1(\mem[5][2] ), .A2(n1161), .ZN(n1158) );
  OAI21_X1 U188 ( .B1(n624), .B2(n1161), .A(n1157), .ZN(n868) );
  NAND2_X1 U189 ( .A1(\mem[5][3] ), .A2(n1161), .ZN(n1157) );
  OAI21_X1 U190 ( .B1(n625), .B2(n1161), .A(n1156), .ZN(n867) );
  NAND2_X1 U191 ( .A1(\mem[5][4] ), .A2(n1161), .ZN(n1156) );
  OAI21_X1 U192 ( .B1(n626), .B2(n1161), .A(n1155), .ZN(n866) );
  NAND2_X1 U193 ( .A1(\mem[5][5] ), .A2(n1161), .ZN(n1155) );
  OAI21_X1 U194 ( .B1(n627), .B2(n1161), .A(n1154), .ZN(n865) );
  NAND2_X1 U195 ( .A1(\mem[5][6] ), .A2(n1161), .ZN(n1154) );
  OAI21_X1 U196 ( .B1(n628), .B2(n1161), .A(n1153), .ZN(n864) );
  NAND2_X1 U197 ( .A1(\mem[5][7] ), .A2(n1161), .ZN(n1153) );
  OAI21_X1 U198 ( .B1(n1212), .B2(n621), .A(n1211), .ZN(n911) );
  NAND2_X1 U199 ( .A1(\mem[0][0] ), .A2(n1212), .ZN(n1211) );
  OAI21_X1 U200 ( .B1(n1212), .B2(n622), .A(n1210), .ZN(n910) );
  NAND2_X1 U201 ( .A1(\mem[0][1] ), .A2(n1212), .ZN(n1210) );
  OAI21_X1 U202 ( .B1(n1212), .B2(n623), .A(n1209), .ZN(n909) );
  NAND2_X1 U203 ( .A1(\mem[0][2] ), .A2(n1212), .ZN(n1209) );
  OAI21_X1 U204 ( .B1(n1212), .B2(n624), .A(n1208), .ZN(n908) );
  NAND2_X1 U205 ( .A1(\mem[0][3] ), .A2(n1212), .ZN(n1208) );
  OAI21_X1 U206 ( .B1(n1212), .B2(n625), .A(n1207), .ZN(n907) );
  NAND2_X1 U207 ( .A1(\mem[0][4] ), .A2(n1212), .ZN(n1207) );
  OAI21_X1 U208 ( .B1(n1212), .B2(n626), .A(n1206), .ZN(n906) );
  NAND2_X1 U209 ( .A1(\mem[0][5] ), .A2(n1212), .ZN(n1206) );
  OAI21_X1 U210 ( .B1(n1212), .B2(n627), .A(n1205), .ZN(n905) );
  NAND2_X1 U211 ( .A1(\mem[0][6] ), .A2(n1212), .ZN(n1205) );
  OAI21_X1 U212 ( .B1(n1212), .B2(n628), .A(n1204), .ZN(n904) );
  NAND2_X1 U213 ( .A1(\mem[0][7] ), .A2(n1212), .ZN(n1204) );
  INV_X1 U214 ( .A(n1130), .ZN(n820) );
  AOI22_X1 U215 ( .A1(data_in[0]), .A2(n844), .B1(n1129), .B2(\mem[8][0] ), 
        .ZN(n1130) );
  INV_X1 U216 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U217 ( .A1(data_in[1]), .A2(n844), .B1(n1129), .B2(\mem[8][1] ), 
        .ZN(n1128) );
  INV_X1 U218 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U219 ( .A1(data_in[2]), .A2(n844), .B1(n1129), .B2(\mem[8][2] ), 
        .ZN(n1127) );
  INV_X1 U220 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U221 ( .A1(data_in[3]), .A2(n844), .B1(n1129), .B2(\mem[8][3] ), 
        .ZN(n1126) );
  INV_X1 U222 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U223 ( .A1(data_in[4]), .A2(n844), .B1(n1129), .B2(\mem[8][4] ), 
        .ZN(n1125) );
  INV_X1 U224 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U225 ( .A1(data_in[5]), .A2(n844), .B1(n1129), .B2(\mem[8][5] ), 
        .ZN(n1124) );
  INV_X1 U226 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U227 ( .A1(data_in[6]), .A2(n844), .B1(n1129), .B2(\mem[8][6] ), 
        .ZN(n1123) );
  INV_X1 U228 ( .A(n1122), .ZN(n813) );
  AOI22_X1 U229 ( .A1(data_in[7]), .A2(n844), .B1(n1129), .B2(\mem[8][7] ), 
        .ZN(n1122) );
  INV_X1 U230 ( .A(n1120), .ZN(n812) );
  AOI22_X1 U231 ( .A1(data_in[0]), .A2(n843), .B1(n1119), .B2(\mem[9][0] ), 
        .ZN(n1120) );
  INV_X1 U232 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U233 ( .A1(data_in[1]), .A2(n843), .B1(n1119), .B2(\mem[9][1] ), 
        .ZN(n1118) );
  INV_X1 U234 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U235 ( .A1(data_in[2]), .A2(n843), .B1(n1119), .B2(\mem[9][2] ), 
        .ZN(n1117) );
  INV_X1 U236 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U237 ( .A1(data_in[3]), .A2(n843), .B1(n1119), .B2(\mem[9][3] ), 
        .ZN(n1116) );
  INV_X1 U238 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U239 ( .A1(data_in[4]), .A2(n843), .B1(n1119), .B2(\mem[9][4] ), 
        .ZN(n1115) );
  INV_X1 U240 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U241 ( .A1(data_in[5]), .A2(n843), .B1(n1119), .B2(\mem[9][5] ), 
        .ZN(n1114) );
  INV_X1 U242 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U243 ( .A1(data_in[6]), .A2(n843), .B1(n1119), .B2(\mem[9][6] ), 
        .ZN(n1113) );
  INV_X1 U244 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U245 ( .A1(data_in[7]), .A2(n843), .B1(n1119), .B2(\mem[9][7] ), 
        .ZN(n1112) );
  INV_X1 U246 ( .A(n1111), .ZN(n804) );
  AOI22_X1 U247 ( .A1(data_in[0]), .A2(n842), .B1(n1110), .B2(\mem[10][0] ), 
        .ZN(n1111) );
  INV_X1 U248 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U249 ( .A1(data_in[1]), .A2(n842), .B1(n1110), .B2(\mem[10][1] ), 
        .ZN(n1109) );
  INV_X1 U250 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U251 ( .A1(data_in[2]), .A2(n842), .B1(n1110), .B2(\mem[10][2] ), 
        .ZN(n1108) );
  INV_X1 U252 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U253 ( .A1(data_in[3]), .A2(n842), .B1(n1110), .B2(\mem[10][3] ), 
        .ZN(n1107) );
  INV_X1 U254 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U255 ( .A1(data_in[4]), .A2(n842), .B1(n1110), .B2(\mem[10][4] ), 
        .ZN(n1106) );
  INV_X1 U256 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U257 ( .A1(data_in[5]), .A2(n842), .B1(n1110), .B2(\mem[10][5] ), 
        .ZN(n1105) );
  INV_X1 U258 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U259 ( .A1(data_in[6]), .A2(n842), .B1(n1110), .B2(\mem[10][6] ), 
        .ZN(n1104) );
  INV_X1 U260 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U261 ( .A1(data_in[7]), .A2(n842), .B1(n1110), .B2(\mem[10][7] ), 
        .ZN(n1103) );
  INV_X1 U262 ( .A(n1102), .ZN(n796) );
  AOI22_X1 U263 ( .A1(data_in[0]), .A2(n841), .B1(n1101), .B2(\mem[11][0] ), 
        .ZN(n1102) );
  INV_X1 U264 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U265 ( .A1(data_in[1]), .A2(n841), .B1(n1101), .B2(\mem[11][1] ), 
        .ZN(n1100) );
  INV_X1 U266 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U267 ( .A1(data_in[2]), .A2(n841), .B1(n1101), .B2(\mem[11][2] ), 
        .ZN(n1099) );
  INV_X1 U268 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U269 ( .A1(data_in[3]), .A2(n841), .B1(n1101), .B2(\mem[11][3] ), 
        .ZN(n1098) );
  INV_X1 U270 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U271 ( .A1(data_in[4]), .A2(n841), .B1(n1101), .B2(\mem[11][4] ), 
        .ZN(n1097) );
  INV_X1 U272 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U273 ( .A1(data_in[5]), .A2(n841), .B1(n1101), .B2(\mem[11][5] ), 
        .ZN(n1096) );
  INV_X1 U274 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U275 ( .A1(data_in[6]), .A2(n841), .B1(n1101), .B2(\mem[11][6] ), 
        .ZN(n1095) );
  INV_X1 U276 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U277 ( .A1(data_in[7]), .A2(n841), .B1(n1101), .B2(\mem[11][7] ), 
        .ZN(n1094) );
  INV_X1 U278 ( .A(n1093), .ZN(n788) );
  AOI22_X1 U279 ( .A1(data_in[0]), .A2(n840), .B1(n1092), .B2(\mem[12][0] ), 
        .ZN(n1093) );
  INV_X1 U280 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U281 ( .A1(data_in[1]), .A2(n840), .B1(n1092), .B2(\mem[12][1] ), 
        .ZN(n1091) );
  INV_X1 U282 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U283 ( .A1(data_in[2]), .A2(n840), .B1(n1092), .B2(\mem[12][2] ), 
        .ZN(n1090) );
  INV_X1 U284 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U285 ( .A1(data_in[3]), .A2(n840), .B1(n1092), .B2(\mem[12][3] ), 
        .ZN(n1089) );
  INV_X1 U286 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U287 ( .A1(data_in[4]), .A2(n840), .B1(n1092), .B2(\mem[12][4] ), 
        .ZN(n1088) );
  INV_X1 U288 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U289 ( .A1(data_in[5]), .A2(n840), .B1(n1092), .B2(\mem[12][5] ), 
        .ZN(n1087) );
  INV_X1 U290 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U291 ( .A1(data_in[6]), .A2(n840), .B1(n1092), .B2(\mem[12][6] ), 
        .ZN(n1086) );
  INV_X1 U292 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U293 ( .A1(data_in[7]), .A2(n840), .B1(n1092), .B2(\mem[12][7] ), 
        .ZN(n1085) );
  INV_X1 U294 ( .A(n1084), .ZN(n780) );
  AOI22_X1 U295 ( .A1(data_in[0]), .A2(n839), .B1(n1083), .B2(\mem[13][0] ), 
        .ZN(n1084) );
  INV_X1 U296 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U297 ( .A1(data_in[1]), .A2(n839), .B1(n1083), .B2(\mem[13][1] ), 
        .ZN(n1082) );
  INV_X1 U298 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U299 ( .A1(data_in[2]), .A2(n839), .B1(n1083), .B2(\mem[13][2] ), 
        .ZN(n1081) );
  INV_X1 U300 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U301 ( .A1(data_in[3]), .A2(n839), .B1(n1083), .B2(\mem[13][3] ), 
        .ZN(n1080) );
  INV_X1 U302 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U303 ( .A1(data_in[4]), .A2(n839), .B1(n1083), .B2(\mem[13][4] ), 
        .ZN(n1079) );
  INV_X1 U304 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U305 ( .A1(data_in[5]), .A2(n839), .B1(n1083), .B2(\mem[13][5] ), 
        .ZN(n1078) );
  INV_X1 U306 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U307 ( .A1(data_in[6]), .A2(n839), .B1(n1083), .B2(\mem[13][6] ), 
        .ZN(n1077) );
  INV_X1 U308 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U309 ( .A1(data_in[7]), .A2(n839), .B1(n1083), .B2(\mem[13][7] ), 
        .ZN(n1076) );
  INV_X1 U310 ( .A(n1075), .ZN(n772) );
  AOI22_X1 U311 ( .A1(data_in[0]), .A2(n838), .B1(n1074), .B2(\mem[14][0] ), 
        .ZN(n1075) );
  INV_X1 U312 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U313 ( .A1(data_in[1]), .A2(n838), .B1(n1074), .B2(\mem[14][1] ), 
        .ZN(n1073) );
  INV_X1 U314 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U315 ( .A1(data_in[2]), .A2(n838), .B1(n1074), .B2(\mem[14][2] ), 
        .ZN(n1072) );
  INV_X1 U316 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U317 ( .A1(data_in[3]), .A2(n838), .B1(n1074), .B2(\mem[14][3] ), 
        .ZN(n1071) );
  INV_X1 U318 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U319 ( .A1(data_in[4]), .A2(n838), .B1(n1074), .B2(\mem[14][4] ), 
        .ZN(n1070) );
  INV_X1 U320 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U321 ( .A1(data_in[5]), .A2(n838), .B1(n1074), .B2(\mem[14][5] ), 
        .ZN(n1069) );
  INV_X1 U322 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U323 ( .A1(data_in[6]), .A2(n838), .B1(n1074), .B2(\mem[14][6] ), 
        .ZN(n1068) );
  INV_X1 U324 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U325 ( .A1(data_in[7]), .A2(n838), .B1(n1074), .B2(\mem[14][7] ), 
        .ZN(n1067) );
  INV_X1 U326 ( .A(n1066), .ZN(n764) );
  AOI22_X1 U327 ( .A1(data_in[0]), .A2(n837), .B1(n1065), .B2(\mem[15][0] ), 
        .ZN(n1066) );
  INV_X1 U328 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U329 ( .A1(data_in[1]), .A2(n837), .B1(n1065), .B2(\mem[15][1] ), 
        .ZN(n1064) );
  INV_X1 U330 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U331 ( .A1(data_in[2]), .A2(n837), .B1(n1065), .B2(\mem[15][2] ), 
        .ZN(n1063) );
  INV_X1 U332 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U333 ( .A1(data_in[3]), .A2(n837), .B1(n1065), .B2(\mem[15][3] ), 
        .ZN(n1062) );
  INV_X1 U334 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U335 ( .A1(data_in[4]), .A2(n837), .B1(n1065), .B2(\mem[15][4] ), 
        .ZN(n1061) );
  INV_X1 U336 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U337 ( .A1(data_in[5]), .A2(n837), .B1(n1065), .B2(\mem[15][5] ), 
        .ZN(n1060) );
  INV_X1 U338 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U339 ( .A1(data_in[6]), .A2(n837), .B1(n1065), .B2(\mem[15][6] ), 
        .ZN(n1059) );
  INV_X1 U340 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U341 ( .A1(data_in[7]), .A2(n837), .B1(n1065), .B2(\mem[15][7] ), 
        .ZN(n1058) );
  INV_X1 U342 ( .A(n1057), .ZN(n756) );
  AOI22_X1 U343 ( .A1(data_in[0]), .A2(n836), .B1(n1056), .B2(\mem[16][0] ), 
        .ZN(n1057) );
  INV_X1 U344 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U345 ( .A1(data_in[1]), .A2(n836), .B1(n1056), .B2(\mem[16][1] ), 
        .ZN(n1055) );
  INV_X1 U346 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U347 ( .A1(data_in[2]), .A2(n836), .B1(n1056), .B2(\mem[16][2] ), 
        .ZN(n1054) );
  INV_X1 U348 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U349 ( .A1(data_in[3]), .A2(n836), .B1(n1056), .B2(\mem[16][3] ), 
        .ZN(n1053) );
  INV_X1 U350 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U351 ( .A1(data_in[4]), .A2(n836), .B1(n1056), .B2(\mem[16][4] ), 
        .ZN(n1052) );
  INV_X1 U352 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U353 ( .A1(data_in[5]), .A2(n836), .B1(n1056), .B2(\mem[16][5] ), 
        .ZN(n1051) );
  INV_X1 U354 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U355 ( .A1(data_in[6]), .A2(n836), .B1(n1056), .B2(\mem[16][6] ), 
        .ZN(n1050) );
  INV_X1 U356 ( .A(n1049), .ZN(n749) );
  AOI22_X1 U357 ( .A1(data_in[7]), .A2(n836), .B1(n1056), .B2(\mem[16][7] ), 
        .ZN(n1049) );
  INV_X1 U358 ( .A(n1047), .ZN(n748) );
  AOI22_X1 U359 ( .A1(data_in[0]), .A2(n835), .B1(n1046), .B2(\mem[17][0] ), 
        .ZN(n1047) );
  INV_X1 U360 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U361 ( .A1(data_in[1]), .A2(n835), .B1(n1046), .B2(\mem[17][1] ), 
        .ZN(n1045) );
  INV_X1 U362 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U363 ( .A1(data_in[2]), .A2(n835), .B1(n1046), .B2(\mem[17][2] ), 
        .ZN(n1044) );
  INV_X1 U364 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[3]), .A2(n835), .B1(n1046), .B2(\mem[17][3] ), 
        .ZN(n1043) );
  INV_X1 U366 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[4]), .A2(n835), .B1(n1046), .B2(\mem[17][4] ), 
        .ZN(n1042) );
  INV_X1 U368 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[5]), .A2(n835), .B1(n1046), .B2(\mem[17][5] ), 
        .ZN(n1041) );
  INV_X1 U370 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[6]), .A2(n835), .B1(n1046), .B2(\mem[17][6] ), 
        .ZN(n1040) );
  INV_X1 U372 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[7]), .A2(n835), .B1(n1046), .B2(\mem[17][7] ), 
        .ZN(n1039) );
  INV_X1 U374 ( .A(n1038), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[0]), .A2(n834), .B1(n1037), .B2(\mem[18][0] ), 
        .ZN(n1038) );
  INV_X1 U376 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[1]), .A2(n834), .B1(n1037), .B2(\mem[18][1] ), 
        .ZN(n1036) );
  INV_X1 U378 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[2]), .A2(n834), .B1(n1037), .B2(\mem[18][2] ), 
        .ZN(n1035) );
  INV_X1 U380 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U381 ( .A1(data_in[3]), .A2(n834), .B1(n1037), .B2(\mem[18][3] ), 
        .ZN(n1034) );
  INV_X1 U382 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U383 ( .A1(data_in[4]), .A2(n834), .B1(n1037), .B2(\mem[18][4] ), 
        .ZN(n1033) );
  INV_X1 U384 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U385 ( .A1(data_in[5]), .A2(n834), .B1(n1037), .B2(\mem[18][5] ), 
        .ZN(n1032) );
  INV_X1 U386 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U387 ( .A1(data_in[6]), .A2(n834), .B1(n1037), .B2(\mem[18][6] ), 
        .ZN(n1031) );
  INV_X1 U388 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U389 ( .A1(data_in[7]), .A2(n834), .B1(n1037), .B2(\mem[18][7] ), 
        .ZN(n1030) );
  INV_X1 U390 ( .A(n1029), .ZN(n732) );
  AOI22_X1 U391 ( .A1(data_in[0]), .A2(n833), .B1(n1028), .B2(\mem[19][0] ), 
        .ZN(n1029) );
  INV_X1 U392 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U393 ( .A1(data_in[1]), .A2(n833), .B1(n1028), .B2(\mem[19][1] ), 
        .ZN(n1027) );
  INV_X1 U394 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U395 ( .A1(data_in[2]), .A2(n833), .B1(n1028), .B2(\mem[19][2] ), 
        .ZN(n1026) );
  INV_X1 U396 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U397 ( .A1(data_in[3]), .A2(n833), .B1(n1028), .B2(\mem[19][3] ), 
        .ZN(n1025) );
  INV_X1 U398 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U399 ( .A1(data_in[4]), .A2(n833), .B1(n1028), .B2(\mem[19][4] ), 
        .ZN(n1024) );
  INV_X1 U400 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U401 ( .A1(data_in[5]), .A2(n833), .B1(n1028), .B2(\mem[19][5] ), 
        .ZN(n1023) );
  INV_X1 U402 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U403 ( .A1(data_in[6]), .A2(n833), .B1(n1028), .B2(\mem[19][6] ), 
        .ZN(n1022) );
  INV_X1 U404 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U405 ( .A1(data_in[7]), .A2(n833), .B1(n1028), .B2(\mem[19][7] ), 
        .ZN(n1021) );
  INV_X1 U406 ( .A(n1020), .ZN(n724) );
  AOI22_X1 U407 ( .A1(data_in[0]), .A2(n832), .B1(n1019), .B2(\mem[20][0] ), 
        .ZN(n1020) );
  INV_X1 U408 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U409 ( .A1(data_in[1]), .A2(n832), .B1(n1019), .B2(\mem[20][1] ), 
        .ZN(n1018) );
  INV_X1 U410 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U411 ( .A1(data_in[2]), .A2(n832), .B1(n1019), .B2(\mem[20][2] ), 
        .ZN(n1017) );
  INV_X1 U412 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U413 ( .A1(data_in[3]), .A2(n832), .B1(n1019), .B2(\mem[20][3] ), 
        .ZN(n1016) );
  INV_X1 U414 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U415 ( .A1(data_in[4]), .A2(n832), .B1(n1019), .B2(\mem[20][4] ), 
        .ZN(n1015) );
  INV_X1 U416 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U417 ( .A1(data_in[5]), .A2(n832), .B1(n1019), .B2(\mem[20][5] ), 
        .ZN(n1014) );
  INV_X1 U418 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U419 ( .A1(data_in[6]), .A2(n832), .B1(n1019), .B2(\mem[20][6] ), 
        .ZN(n1013) );
  INV_X1 U420 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U421 ( .A1(data_in[7]), .A2(n832), .B1(n1019), .B2(\mem[20][7] ), 
        .ZN(n1012) );
  INV_X1 U422 ( .A(n1011), .ZN(n716) );
  AOI22_X1 U423 ( .A1(data_in[0]), .A2(n831), .B1(n1010), .B2(\mem[21][0] ), 
        .ZN(n1011) );
  INV_X1 U424 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U425 ( .A1(data_in[1]), .A2(n831), .B1(n1010), .B2(\mem[21][1] ), 
        .ZN(n1009) );
  INV_X1 U426 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U427 ( .A1(data_in[2]), .A2(n831), .B1(n1010), .B2(\mem[21][2] ), 
        .ZN(n1008) );
  INV_X1 U428 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U429 ( .A1(data_in[3]), .A2(n831), .B1(n1010), .B2(\mem[21][3] ), 
        .ZN(n1007) );
  INV_X1 U430 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U431 ( .A1(data_in[4]), .A2(n831), .B1(n1010), .B2(\mem[21][4] ), 
        .ZN(n1006) );
  INV_X1 U432 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U433 ( .A1(data_in[5]), .A2(n831), .B1(n1010), .B2(\mem[21][5] ), 
        .ZN(n1005) );
  INV_X1 U434 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U435 ( .A1(data_in[6]), .A2(n831), .B1(n1010), .B2(\mem[21][6] ), 
        .ZN(n1004) );
  INV_X1 U436 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U437 ( .A1(data_in[7]), .A2(n831), .B1(n1010), .B2(\mem[21][7] ), 
        .ZN(n1003) );
  INV_X1 U438 ( .A(n1002), .ZN(n708) );
  AOI22_X1 U439 ( .A1(data_in[0]), .A2(n830), .B1(n1001), .B2(\mem[22][0] ), 
        .ZN(n1002) );
  INV_X1 U440 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U441 ( .A1(data_in[1]), .A2(n830), .B1(n1001), .B2(\mem[22][1] ), 
        .ZN(n1000) );
  INV_X1 U442 ( .A(n999), .ZN(n706) );
  AOI22_X1 U443 ( .A1(data_in[2]), .A2(n830), .B1(n1001), .B2(\mem[22][2] ), 
        .ZN(n999) );
  INV_X1 U444 ( .A(n998), .ZN(n705) );
  AOI22_X1 U445 ( .A1(data_in[3]), .A2(n830), .B1(n1001), .B2(\mem[22][3] ), 
        .ZN(n998) );
  INV_X1 U446 ( .A(n997), .ZN(n704) );
  AOI22_X1 U447 ( .A1(data_in[4]), .A2(n830), .B1(n1001), .B2(\mem[22][4] ), 
        .ZN(n997) );
  INV_X1 U448 ( .A(n996), .ZN(n703) );
  AOI22_X1 U449 ( .A1(data_in[5]), .A2(n830), .B1(n1001), .B2(\mem[22][5] ), 
        .ZN(n996) );
  INV_X1 U450 ( .A(n995), .ZN(n702) );
  AOI22_X1 U451 ( .A1(data_in[6]), .A2(n830), .B1(n1001), .B2(\mem[22][6] ), 
        .ZN(n995) );
  INV_X1 U452 ( .A(n994), .ZN(n701) );
  AOI22_X1 U453 ( .A1(data_in[7]), .A2(n830), .B1(n1001), .B2(\mem[22][7] ), 
        .ZN(n994) );
  INV_X1 U454 ( .A(n993), .ZN(n700) );
  AOI22_X1 U455 ( .A1(data_in[0]), .A2(n829), .B1(n992), .B2(\mem[23][0] ), 
        .ZN(n993) );
  INV_X1 U456 ( .A(n991), .ZN(n699) );
  AOI22_X1 U457 ( .A1(data_in[1]), .A2(n829), .B1(n992), .B2(\mem[23][1] ), 
        .ZN(n991) );
  INV_X1 U458 ( .A(n990), .ZN(n698) );
  AOI22_X1 U459 ( .A1(data_in[2]), .A2(n829), .B1(n992), .B2(\mem[23][2] ), 
        .ZN(n990) );
  INV_X1 U460 ( .A(n989), .ZN(n697) );
  AOI22_X1 U461 ( .A1(data_in[3]), .A2(n829), .B1(n992), .B2(\mem[23][3] ), 
        .ZN(n989) );
  INV_X1 U462 ( .A(n988), .ZN(n696) );
  AOI22_X1 U463 ( .A1(data_in[4]), .A2(n829), .B1(n992), .B2(\mem[23][4] ), 
        .ZN(n988) );
  INV_X1 U464 ( .A(n987), .ZN(n695) );
  AOI22_X1 U465 ( .A1(data_in[5]), .A2(n829), .B1(n992), .B2(\mem[23][5] ), 
        .ZN(n987) );
  INV_X1 U466 ( .A(n986), .ZN(n694) );
  AOI22_X1 U467 ( .A1(data_in[6]), .A2(n829), .B1(n992), .B2(\mem[23][6] ), 
        .ZN(n986) );
  INV_X1 U468 ( .A(n985), .ZN(n693) );
  AOI22_X1 U469 ( .A1(data_in[7]), .A2(n829), .B1(n992), .B2(\mem[23][7] ), 
        .ZN(n985) );
  INV_X1 U470 ( .A(n984), .ZN(n692) );
  AOI22_X1 U471 ( .A1(data_in[0]), .A2(n828), .B1(n983), .B2(\mem[24][0] ), 
        .ZN(n984) );
  INV_X1 U472 ( .A(n982), .ZN(n691) );
  AOI22_X1 U473 ( .A1(data_in[1]), .A2(n828), .B1(n983), .B2(\mem[24][1] ), 
        .ZN(n982) );
  INV_X1 U474 ( .A(n981), .ZN(n690) );
  AOI22_X1 U475 ( .A1(data_in[2]), .A2(n828), .B1(n983), .B2(\mem[24][2] ), 
        .ZN(n981) );
  INV_X1 U476 ( .A(n980), .ZN(n689) );
  AOI22_X1 U477 ( .A1(data_in[3]), .A2(n828), .B1(n983), .B2(\mem[24][3] ), 
        .ZN(n980) );
  INV_X1 U478 ( .A(n979), .ZN(n688) );
  AOI22_X1 U479 ( .A1(data_in[4]), .A2(n828), .B1(n983), .B2(\mem[24][4] ), 
        .ZN(n979) );
  INV_X1 U480 ( .A(n978), .ZN(n687) );
  AOI22_X1 U481 ( .A1(data_in[5]), .A2(n828), .B1(n983), .B2(\mem[24][5] ), 
        .ZN(n978) );
  INV_X1 U482 ( .A(n977), .ZN(n686) );
  AOI22_X1 U483 ( .A1(data_in[6]), .A2(n828), .B1(n983), .B2(\mem[24][6] ), 
        .ZN(n977) );
  INV_X1 U484 ( .A(n976), .ZN(n685) );
  AOI22_X1 U485 ( .A1(data_in[7]), .A2(n828), .B1(n983), .B2(\mem[24][7] ), 
        .ZN(n976) );
  INV_X1 U486 ( .A(n974), .ZN(n684) );
  AOI22_X1 U487 ( .A1(data_in[0]), .A2(n827), .B1(n973), .B2(\mem[25][0] ), 
        .ZN(n974) );
  INV_X1 U488 ( .A(n972), .ZN(n683) );
  AOI22_X1 U489 ( .A1(data_in[1]), .A2(n827), .B1(n973), .B2(\mem[25][1] ), 
        .ZN(n972) );
  INV_X1 U490 ( .A(n971), .ZN(n682) );
  AOI22_X1 U491 ( .A1(data_in[2]), .A2(n827), .B1(n973), .B2(\mem[25][2] ), 
        .ZN(n971) );
  INV_X1 U492 ( .A(n970), .ZN(n681) );
  AOI22_X1 U493 ( .A1(data_in[3]), .A2(n827), .B1(n973), .B2(\mem[25][3] ), 
        .ZN(n970) );
  INV_X1 U494 ( .A(n969), .ZN(n680) );
  AOI22_X1 U495 ( .A1(data_in[4]), .A2(n827), .B1(n973), .B2(\mem[25][4] ), 
        .ZN(n969) );
  INV_X1 U496 ( .A(n968), .ZN(n679) );
  AOI22_X1 U497 ( .A1(data_in[5]), .A2(n827), .B1(n973), .B2(\mem[25][5] ), 
        .ZN(n968) );
  INV_X1 U498 ( .A(n967), .ZN(n678) );
  AOI22_X1 U499 ( .A1(data_in[6]), .A2(n827), .B1(n973), .B2(\mem[25][6] ), 
        .ZN(n967) );
  INV_X1 U500 ( .A(n966), .ZN(n677) );
  AOI22_X1 U501 ( .A1(data_in[7]), .A2(n827), .B1(n973), .B2(\mem[25][7] ), 
        .ZN(n966) );
  INV_X1 U502 ( .A(n965), .ZN(n676) );
  AOI22_X1 U503 ( .A1(data_in[0]), .A2(n826), .B1(n964), .B2(\mem[26][0] ), 
        .ZN(n965) );
  INV_X1 U504 ( .A(n963), .ZN(n675) );
  AOI22_X1 U505 ( .A1(data_in[1]), .A2(n826), .B1(n964), .B2(\mem[26][1] ), 
        .ZN(n963) );
  INV_X1 U506 ( .A(n962), .ZN(n674) );
  AOI22_X1 U507 ( .A1(data_in[2]), .A2(n826), .B1(n964), .B2(\mem[26][2] ), 
        .ZN(n962) );
  INV_X1 U508 ( .A(n961), .ZN(n673) );
  AOI22_X1 U509 ( .A1(data_in[3]), .A2(n826), .B1(n964), .B2(\mem[26][3] ), 
        .ZN(n961) );
  INV_X1 U510 ( .A(n960), .ZN(n672) );
  AOI22_X1 U511 ( .A1(data_in[4]), .A2(n826), .B1(n964), .B2(\mem[26][4] ), 
        .ZN(n960) );
  INV_X1 U512 ( .A(n959), .ZN(n671) );
  AOI22_X1 U513 ( .A1(data_in[5]), .A2(n826), .B1(n964), .B2(\mem[26][5] ), 
        .ZN(n959) );
  INV_X1 U514 ( .A(n958), .ZN(n670) );
  AOI22_X1 U515 ( .A1(data_in[6]), .A2(n826), .B1(n964), .B2(\mem[26][6] ), 
        .ZN(n958) );
  INV_X1 U516 ( .A(n957), .ZN(n669) );
  AOI22_X1 U517 ( .A1(data_in[7]), .A2(n826), .B1(n964), .B2(\mem[26][7] ), 
        .ZN(n957) );
  INV_X1 U518 ( .A(n956), .ZN(n668) );
  AOI22_X1 U519 ( .A1(data_in[0]), .A2(n825), .B1(n955), .B2(\mem[27][0] ), 
        .ZN(n956) );
  INV_X1 U520 ( .A(n954), .ZN(n667) );
  AOI22_X1 U521 ( .A1(data_in[1]), .A2(n825), .B1(n955), .B2(\mem[27][1] ), 
        .ZN(n954) );
  INV_X1 U522 ( .A(n953), .ZN(n666) );
  AOI22_X1 U523 ( .A1(data_in[2]), .A2(n825), .B1(n955), .B2(\mem[27][2] ), 
        .ZN(n953) );
  INV_X1 U524 ( .A(n952), .ZN(n665) );
  AOI22_X1 U525 ( .A1(data_in[3]), .A2(n825), .B1(n955), .B2(\mem[27][3] ), 
        .ZN(n952) );
  INV_X1 U526 ( .A(n951), .ZN(n664) );
  AOI22_X1 U527 ( .A1(data_in[4]), .A2(n825), .B1(n955), .B2(\mem[27][4] ), 
        .ZN(n951) );
  INV_X1 U528 ( .A(n950), .ZN(n663) );
  AOI22_X1 U529 ( .A1(data_in[5]), .A2(n825), .B1(n955), .B2(\mem[27][5] ), 
        .ZN(n950) );
  INV_X1 U530 ( .A(n949), .ZN(n662) );
  AOI22_X1 U531 ( .A1(data_in[6]), .A2(n825), .B1(n955), .B2(\mem[27][6] ), 
        .ZN(n949) );
  INV_X1 U532 ( .A(n948), .ZN(n661) );
  AOI22_X1 U533 ( .A1(data_in[7]), .A2(n825), .B1(n955), .B2(\mem[27][7] ), 
        .ZN(n948) );
  INV_X1 U534 ( .A(n947), .ZN(n660) );
  AOI22_X1 U535 ( .A1(data_in[0]), .A2(n824), .B1(n946), .B2(\mem[28][0] ), 
        .ZN(n947) );
  INV_X1 U536 ( .A(n945), .ZN(n659) );
  AOI22_X1 U537 ( .A1(data_in[1]), .A2(n824), .B1(n946), .B2(\mem[28][1] ), 
        .ZN(n945) );
  INV_X1 U538 ( .A(n944), .ZN(n658) );
  AOI22_X1 U539 ( .A1(data_in[2]), .A2(n824), .B1(n946), .B2(\mem[28][2] ), 
        .ZN(n944) );
  INV_X1 U540 ( .A(n943), .ZN(n657) );
  AOI22_X1 U541 ( .A1(data_in[3]), .A2(n824), .B1(n946), .B2(\mem[28][3] ), 
        .ZN(n943) );
  INV_X1 U542 ( .A(n942), .ZN(n656) );
  AOI22_X1 U543 ( .A1(data_in[4]), .A2(n824), .B1(n946), .B2(\mem[28][4] ), 
        .ZN(n942) );
  INV_X1 U544 ( .A(n941), .ZN(n655) );
  AOI22_X1 U545 ( .A1(data_in[5]), .A2(n824), .B1(n946), .B2(\mem[28][5] ), 
        .ZN(n941) );
  INV_X1 U546 ( .A(n940), .ZN(n654) );
  AOI22_X1 U547 ( .A1(data_in[6]), .A2(n824), .B1(n946), .B2(\mem[28][6] ), 
        .ZN(n940) );
  INV_X1 U548 ( .A(n939), .ZN(n653) );
  AOI22_X1 U549 ( .A1(data_in[7]), .A2(n824), .B1(n946), .B2(\mem[28][7] ), 
        .ZN(n939) );
  INV_X1 U550 ( .A(n938), .ZN(n652) );
  AOI22_X1 U551 ( .A1(data_in[0]), .A2(n823), .B1(n937), .B2(\mem[29][0] ), 
        .ZN(n938) );
  INV_X1 U552 ( .A(n936), .ZN(n651) );
  AOI22_X1 U553 ( .A1(data_in[1]), .A2(n823), .B1(n937), .B2(\mem[29][1] ), 
        .ZN(n936) );
  INV_X1 U554 ( .A(n935), .ZN(n650) );
  AOI22_X1 U555 ( .A1(data_in[2]), .A2(n823), .B1(n937), .B2(\mem[29][2] ), 
        .ZN(n935) );
  INV_X1 U556 ( .A(n934), .ZN(n649) );
  AOI22_X1 U557 ( .A1(data_in[3]), .A2(n823), .B1(n937), .B2(\mem[29][3] ), 
        .ZN(n934) );
  INV_X1 U558 ( .A(n933), .ZN(n648) );
  AOI22_X1 U559 ( .A1(data_in[4]), .A2(n823), .B1(n937), .B2(\mem[29][4] ), 
        .ZN(n933) );
  INV_X1 U560 ( .A(n932), .ZN(n647) );
  AOI22_X1 U561 ( .A1(data_in[5]), .A2(n823), .B1(n937), .B2(\mem[29][5] ), 
        .ZN(n932) );
  INV_X1 U562 ( .A(n931), .ZN(n646) );
  AOI22_X1 U563 ( .A1(data_in[6]), .A2(n823), .B1(n937), .B2(\mem[29][6] ), 
        .ZN(n931) );
  INV_X1 U564 ( .A(n930), .ZN(n645) );
  AOI22_X1 U565 ( .A1(data_in[7]), .A2(n823), .B1(n937), .B2(\mem[29][7] ), 
        .ZN(n930) );
  INV_X1 U566 ( .A(n929), .ZN(n644) );
  AOI22_X1 U567 ( .A1(data_in[0]), .A2(n822), .B1(n928), .B2(\mem[30][0] ), 
        .ZN(n929) );
  INV_X1 U568 ( .A(n927), .ZN(n643) );
  AOI22_X1 U569 ( .A1(data_in[1]), .A2(n822), .B1(n928), .B2(\mem[30][1] ), 
        .ZN(n927) );
  INV_X1 U570 ( .A(n926), .ZN(n642) );
  AOI22_X1 U571 ( .A1(data_in[2]), .A2(n822), .B1(n928), .B2(\mem[30][2] ), 
        .ZN(n926) );
  INV_X1 U572 ( .A(n925), .ZN(n641) );
  AOI22_X1 U573 ( .A1(data_in[3]), .A2(n822), .B1(n928), .B2(\mem[30][3] ), 
        .ZN(n925) );
  INV_X1 U574 ( .A(n924), .ZN(n640) );
  AOI22_X1 U575 ( .A1(data_in[4]), .A2(n822), .B1(n928), .B2(\mem[30][4] ), 
        .ZN(n924) );
  INV_X1 U576 ( .A(n923), .ZN(n639) );
  AOI22_X1 U577 ( .A1(data_in[5]), .A2(n822), .B1(n928), .B2(\mem[30][5] ), 
        .ZN(n923) );
  INV_X1 U578 ( .A(n922), .ZN(n638) );
  AOI22_X1 U579 ( .A1(data_in[6]), .A2(n822), .B1(n928), .B2(\mem[30][6] ), 
        .ZN(n922) );
  INV_X1 U580 ( .A(n921), .ZN(n637) );
  AOI22_X1 U581 ( .A1(data_in[7]), .A2(n822), .B1(n928), .B2(\mem[30][7] ), 
        .ZN(n921) );
  INV_X1 U582 ( .A(n920), .ZN(n636) );
  AOI22_X1 U583 ( .A1(data_in[0]), .A2(n821), .B1(n919), .B2(\mem[31][0] ), 
        .ZN(n920) );
  INV_X1 U584 ( .A(n918), .ZN(n635) );
  AOI22_X1 U585 ( .A1(data_in[1]), .A2(n821), .B1(n919), .B2(\mem[31][1] ), 
        .ZN(n918) );
  INV_X1 U586 ( .A(n917), .ZN(n634) );
  AOI22_X1 U587 ( .A1(data_in[2]), .A2(n821), .B1(n919), .B2(\mem[31][2] ), 
        .ZN(n917) );
  INV_X1 U588 ( .A(n916), .ZN(n633) );
  AOI22_X1 U589 ( .A1(data_in[3]), .A2(n821), .B1(n919), .B2(\mem[31][3] ), 
        .ZN(n916) );
  INV_X1 U590 ( .A(n915), .ZN(n632) );
  AOI22_X1 U591 ( .A1(data_in[4]), .A2(n821), .B1(n919), .B2(\mem[31][4] ), 
        .ZN(n915) );
  INV_X1 U592 ( .A(n914), .ZN(n631) );
  AOI22_X1 U593 ( .A1(data_in[5]), .A2(n821), .B1(n919), .B2(\mem[31][5] ), 
        .ZN(n914) );
  INV_X1 U594 ( .A(n913), .ZN(n630) );
  AOI22_X1 U595 ( .A1(data_in[6]), .A2(n821), .B1(n919), .B2(\mem[31][6] ), 
        .ZN(n913) );
  INV_X1 U596 ( .A(n912), .ZN(n629) );
  AOI22_X1 U597 ( .A1(data_in[7]), .A2(n821), .B1(n919), .B2(\mem[31][7] ), 
        .ZN(n912) );
  MUX2_X1 U598 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n616), .Z(n3) );
  MUX2_X1 U599 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n615), .Z(n4) );
  MUX2_X1 U600 ( .A(n4), .B(n3), .S(n610), .Z(n5) );
  MUX2_X1 U601 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n617), .Z(n6) );
  MUX2_X1 U602 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n616), .Z(n7) );
  MUX2_X1 U603 ( .A(n7), .B(n6), .S(n610), .Z(n8) );
  MUX2_X1 U604 ( .A(n8), .B(n5), .S(n608), .Z(n9) );
  MUX2_X1 U605 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n614), .Z(n10) );
  MUX2_X1 U606 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n615), .Z(n11) );
  MUX2_X1 U607 ( .A(n11), .B(n10), .S(n610), .Z(n12) );
  MUX2_X1 U608 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n617), .Z(n13) );
  MUX2_X1 U609 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n614), .Z(n14) );
  MUX2_X1 U610 ( .A(n14), .B(n13), .S(n610), .Z(n15) );
  MUX2_X1 U611 ( .A(n15), .B(n12), .S(n608), .Z(n16) );
  MUX2_X1 U612 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U613 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n615), .Z(n18) );
  MUX2_X1 U614 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n618), .Z(n19) );
  MUX2_X1 U615 ( .A(n19), .B(n18), .S(n611), .Z(n20) );
  MUX2_X1 U616 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n618), .Z(n21) );
  MUX2_X1 U617 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n22) );
  MUX2_X1 U618 ( .A(n22), .B(n21), .S(n611), .Z(n23) );
  MUX2_X1 U619 ( .A(n23), .B(n20), .S(n608), .Z(n24) );
  MUX2_X1 U620 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n618), .Z(n25) );
  MUX2_X1 U621 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n26) );
  MUX2_X1 U622 ( .A(n26), .B(n25), .S(n611), .Z(n27) );
  MUX2_X1 U623 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n28) );
  MUX2_X1 U624 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n29) );
  MUX2_X1 U625 ( .A(n29), .B(n28), .S(n611), .Z(n30) );
  MUX2_X1 U626 ( .A(n30), .B(n27), .S(n608), .Z(n31) );
  MUX2_X1 U627 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U628 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U629 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n616), .Z(n33) );
  MUX2_X1 U630 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n618), .Z(n34) );
  MUX2_X1 U631 ( .A(n34), .B(n33), .S(n611), .Z(n35) );
  MUX2_X1 U632 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n614), .Z(n36) );
  MUX2_X1 U633 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(N10), .Z(n37) );
  MUX2_X1 U634 ( .A(n37), .B(n36), .S(n611), .Z(n38) );
  MUX2_X1 U635 ( .A(n38), .B(n35), .S(n608), .Z(n39) );
  MUX2_X1 U636 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n613), .Z(n40) );
  MUX2_X1 U637 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n613), .Z(n41) );
  MUX2_X1 U638 ( .A(n41), .B(n40), .S(n611), .Z(n42) );
  MUX2_X1 U639 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n613), .Z(n43) );
  MUX2_X1 U640 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n613), .Z(n44) );
  MUX2_X1 U641 ( .A(n44), .B(n43), .S(n611), .Z(n45) );
  MUX2_X1 U642 ( .A(n45), .B(n42), .S(n608), .Z(n46) );
  MUX2_X1 U643 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U644 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n613), .Z(n48) );
  MUX2_X1 U645 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n613), .Z(n49) );
  MUX2_X1 U646 ( .A(n49), .B(n48), .S(n611), .Z(n50) );
  MUX2_X1 U647 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n613), .Z(n51) );
  MUX2_X1 U648 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n613), .Z(n52) );
  MUX2_X1 U649 ( .A(n52), .B(n51), .S(n611), .Z(n53) );
  MUX2_X1 U650 ( .A(n53), .B(n50), .S(n608), .Z(n54) );
  MUX2_X1 U651 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n613), .Z(n55) );
  MUX2_X1 U652 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n613), .Z(n56) );
  MUX2_X1 U653 ( .A(n56), .B(n55), .S(n611), .Z(n57) );
  MUX2_X1 U654 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n613), .Z(n58) );
  MUX2_X1 U655 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n613), .Z(n59) );
  MUX2_X1 U656 ( .A(n59), .B(n58), .S(n611), .Z(n60) );
  MUX2_X1 U657 ( .A(n60), .B(n57), .S(n608), .Z(n61) );
  MUX2_X1 U658 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U659 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U660 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n614), .Z(n63) );
  MUX2_X1 U661 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n614), .Z(n64) );
  MUX2_X1 U662 ( .A(n64), .B(n63), .S(n612), .Z(n65) );
  MUX2_X1 U663 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n614), .Z(n66) );
  MUX2_X1 U664 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n614), .Z(n67) );
  MUX2_X1 U665 ( .A(n67), .B(n66), .S(n612), .Z(n68) );
  MUX2_X1 U666 ( .A(n68), .B(n65), .S(n609), .Z(n69) );
  MUX2_X1 U667 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n614), .Z(n70) );
  MUX2_X1 U668 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n614), .Z(n71) );
  MUX2_X1 U669 ( .A(n71), .B(n70), .S(n612), .Z(n72) );
  MUX2_X1 U670 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n614), .Z(n73) );
  MUX2_X1 U671 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n614), .Z(n74) );
  MUX2_X1 U672 ( .A(n74), .B(n73), .S(n612), .Z(n75) );
  MUX2_X1 U673 ( .A(n75), .B(n72), .S(n609), .Z(n76) );
  MUX2_X1 U674 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U675 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n614), .Z(n78) );
  MUX2_X1 U676 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n614), .Z(n79) );
  MUX2_X1 U677 ( .A(n79), .B(n78), .S(n612), .Z(n80) );
  MUX2_X1 U678 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n614), .Z(n81) );
  MUX2_X1 U679 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n614), .Z(n82) );
  MUX2_X1 U680 ( .A(n82), .B(n81), .S(n612), .Z(n83) );
  MUX2_X1 U681 ( .A(n83), .B(n80), .S(n609), .Z(n84) );
  MUX2_X1 U682 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n615), .Z(n85) );
  MUX2_X1 U683 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n615), .Z(n86) );
  MUX2_X1 U684 ( .A(n86), .B(n85), .S(n612), .Z(n87) );
  MUX2_X1 U685 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n615), .Z(n88) );
  MUX2_X1 U686 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n615), .Z(n89) );
  MUX2_X1 U687 ( .A(n89), .B(n88), .S(n612), .Z(n90) );
  MUX2_X1 U688 ( .A(n90), .B(n87), .S(n609), .Z(n91) );
  MUX2_X1 U689 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U690 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U691 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n615), .Z(n93) );
  MUX2_X1 U692 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n615), .Z(n94) );
  MUX2_X1 U693 ( .A(n94), .B(n93), .S(n612), .Z(n95) );
  MUX2_X1 U694 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n615), .Z(n96) );
  MUX2_X1 U695 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n615), .Z(n97) );
  MUX2_X1 U696 ( .A(n97), .B(n96), .S(n612), .Z(n98) );
  MUX2_X1 U697 ( .A(n98), .B(n95), .S(n609), .Z(n99) );
  MUX2_X1 U698 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n615), .Z(n100) );
  MUX2_X1 U699 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n615), .Z(n101) );
  MUX2_X1 U700 ( .A(n101), .B(n100), .S(n612), .Z(n102) );
  MUX2_X1 U701 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n615), .Z(n103) );
  MUX2_X1 U702 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n615), .Z(n104) );
  MUX2_X1 U703 ( .A(n104), .B(n103), .S(n612), .Z(n105) );
  MUX2_X1 U704 ( .A(n105), .B(n102), .S(n609), .Z(n106) );
  MUX2_X1 U705 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U706 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n618), .Z(n108) );
  MUX2_X1 U707 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n618), .Z(n109) );
  MUX2_X1 U708 ( .A(n109), .B(n108), .S(n611), .Z(n110) );
  MUX2_X1 U709 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n618), .Z(n111) );
  MUX2_X1 U710 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n618), .Z(n112) );
  MUX2_X1 U711 ( .A(n112), .B(n111), .S(n612), .Z(n113) );
  MUX2_X1 U712 ( .A(n113), .B(n110), .S(n609), .Z(n114) );
  MUX2_X1 U713 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n615), .Z(n115) );
  MUX2_X1 U714 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n614), .Z(n116) );
  MUX2_X1 U715 ( .A(n116), .B(n115), .S(n610), .Z(n117) );
  MUX2_X1 U716 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n614), .Z(n118) );
  MUX2_X1 U717 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n618), .Z(n119) );
  MUX2_X1 U718 ( .A(n119), .B(n118), .S(n610), .Z(n120) );
  MUX2_X1 U719 ( .A(n120), .B(n117), .S(n609), .Z(n121) );
  MUX2_X1 U720 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U721 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U722 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n617), .Z(n123) );
  MUX2_X1 U723 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n616), .Z(n124) );
  MUX2_X1 U724 ( .A(n124), .B(n123), .S(n610), .Z(n125) );
  MUX2_X1 U725 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n618), .Z(n126) );
  MUX2_X1 U726 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n618), .Z(n127) );
  MUX2_X1 U727 ( .A(n127), .B(n126), .S(n611), .Z(n128) );
  MUX2_X1 U728 ( .A(n128), .B(n125), .S(n609), .Z(n129) );
  MUX2_X1 U729 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n616), .Z(n130) );
  MUX2_X1 U730 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n618), .Z(n131) );
  MUX2_X1 U731 ( .A(n131), .B(n130), .S(N11), .Z(n132) );
  MUX2_X1 U732 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n618), .Z(n133) );
  MUX2_X1 U733 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n618), .Z(n134) );
  MUX2_X1 U734 ( .A(n134), .B(n133), .S(n611), .Z(n135) );
  MUX2_X1 U735 ( .A(n135), .B(n132), .S(n609), .Z(n136) );
  MUX2_X1 U736 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U737 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n617), .Z(n138) );
  MUX2_X1 U738 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n618), .Z(n139) );
  MUX2_X1 U739 ( .A(n139), .B(n138), .S(n612), .Z(n140) );
  MUX2_X1 U740 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n616), .Z(n141) );
  MUX2_X1 U741 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n615), .Z(n142) );
  MUX2_X1 U742 ( .A(n142), .B(n141), .S(n610), .Z(n143) );
  MUX2_X1 U743 ( .A(n143), .B(n140), .S(n609), .Z(n144) );
  MUX2_X1 U744 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n617), .Z(n145) );
  MUX2_X1 U745 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n618), .Z(n146) );
  MUX2_X1 U746 ( .A(n146), .B(n145), .S(n611), .Z(n147) );
  MUX2_X1 U747 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n618), .Z(n148) );
  MUX2_X1 U748 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n618), .Z(n149) );
  MUX2_X1 U749 ( .A(n149), .B(n148), .S(n611), .Z(n150) );
  MUX2_X1 U750 ( .A(n150), .B(n147), .S(n609), .Z(n151) );
  MUX2_X1 U751 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U752 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U753 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n613), .Z(n153) );
  MUX2_X1 U754 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n613), .Z(n154) );
  MUX2_X1 U755 ( .A(n154), .B(n153), .S(n611), .Z(n155) );
  MUX2_X1 U756 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n613), .Z(n156) );
  MUX2_X1 U757 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n613), .Z(n157) );
  MUX2_X1 U758 ( .A(n157), .B(n156), .S(n612), .Z(n158) );
  MUX2_X1 U759 ( .A(n158), .B(n155), .S(n608), .Z(n159) );
  MUX2_X1 U760 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n613), .Z(n160) );
  MUX2_X1 U761 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n613), .Z(n161) );
  MUX2_X1 U762 ( .A(n161), .B(n160), .S(n610), .Z(n162) );
  MUX2_X1 U763 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n613), .Z(n163) );
  MUX2_X1 U764 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n614), .Z(n164) );
  MUX2_X1 U765 ( .A(n164), .B(n163), .S(N11), .Z(n165) );
  MUX2_X1 U766 ( .A(n165), .B(n162), .S(N12), .Z(n166) );
  MUX2_X1 U767 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U768 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n613), .Z(n168) );
  MUX2_X1 U769 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n613), .Z(n169) );
  MUX2_X1 U770 ( .A(n169), .B(n168), .S(n610), .Z(n170) );
  MUX2_X1 U771 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n613), .Z(n171) );
  MUX2_X1 U772 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n613), .Z(n172) );
  MUX2_X1 U773 ( .A(n172), .B(n171), .S(N11), .Z(n173) );
  MUX2_X1 U774 ( .A(n173), .B(n170), .S(n608), .Z(n174) );
  MUX2_X1 U775 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n616), .Z(n175) );
  MUX2_X1 U776 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n616), .Z(n176) );
  MUX2_X1 U777 ( .A(n176), .B(n175), .S(N11), .Z(n177) );
  MUX2_X1 U778 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n616), .Z(n178) );
  MUX2_X1 U779 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n616), .Z(n179) );
  MUX2_X1 U780 ( .A(n179), .B(n178), .S(n611), .Z(n180) );
  MUX2_X1 U781 ( .A(n180), .B(n177), .S(n609), .Z(n181) );
  MUX2_X1 U782 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U783 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U784 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n616), .Z(n183) );
  MUX2_X1 U785 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n616), .Z(n184) );
  MUX2_X1 U786 ( .A(n184), .B(n183), .S(n612), .Z(n185) );
  MUX2_X1 U787 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n616), .Z(n186) );
  MUX2_X1 U788 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n616), .Z(n187) );
  MUX2_X1 U789 ( .A(n187), .B(n186), .S(n612), .Z(n188) );
  MUX2_X1 U790 ( .A(n188), .B(n185), .S(n608), .Z(n189) );
  MUX2_X1 U791 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n616), .Z(n190) );
  MUX2_X1 U792 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n616), .Z(n191) );
  MUX2_X1 U793 ( .A(n191), .B(n190), .S(n611), .Z(n192) );
  MUX2_X1 U794 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n616), .Z(n193) );
  MUX2_X1 U795 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n616), .Z(n194) );
  MUX2_X1 U796 ( .A(n194), .B(n193), .S(N11), .Z(n195) );
  MUX2_X1 U797 ( .A(n195), .B(n192), .S(N12), .Z(n196) );
  MUX2_X1 U798 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U799 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n617), .Z(n198) );
  MUX2_X1 U800 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n617), .Z(n199) );
  MUX2_X1 U801 ( .A(n199), .B(n198), .S(n610), .Z(n200) );
  MUX2_X1 U802 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n617), .Z(n201) );
  MUX2_X1 U803 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n617), .Z(n202) );
  MUX2_X1 U804 ( .A(n202), .B(n201), .S(n611), .Z(n203) );
  MUX2_X1 U805 ( .A(n203), .B(n200), .S(n609), .Z(n204) );
  MUX2_X1 U806 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n617), .Z(n205) );
  MUX2_X1 U807 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n617), .Z(n206) );
  MUX2_X1 U808 ( .A(n206), .B(n205), .S(n610), .Z(n207) );
  MUX2_X1 U809 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n617), .Z(n208) );
  MUX2_X1 U810 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n617), .Z(n209) );
  MUX2_X1 U811 ( .A(n209), .B(n208), .S(n612), .Z(n210) );
  MUX2_X1 U812 ( .A(n210), .B(n207), .S(n608), .Z(n211) );
  MUX2_X1 U813 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U814 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U815 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n617), .Z(n213) );
  MUX2_X1 U816 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n617), .Z(n214) );
  MUX2_X1 U817 ( .A(n214), .B(n213), .S(n610), .Z(n215) );
  MUX2_X1 U818 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n617), .Z(n216) );
  MUX2_X1 U819 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n617), .Z(n217) );
  MUX2_X1 U820 ( .A(n217), .B(n216), .S(n610), .Z(n218) );
  MUX2_X1 U821 ( .A(n218), .B(n215), .S(n608), .Z(n219) );
  MUX2_X1 U822 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n615), .Z(n220) );
  MUX2_X1 U823 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n618), .Z(n221) );
  MUX2_X1 U824 ( .A(n221), .B(n220), .S(n610), .Z(n222) );
  MUX2_X1 U825 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n616), .Z(n223) );
  MUX2_X1 U826 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n615), .Z(n224) );
  MUX2_X1 U827 ( .A(n224), .B(n223), .S(n612), .Z(n225) );
  MUX2_X1 U828 ( .A(n225), .B(n222), .S(N12), .Z(n226) );
  MUX2_X1 U829 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U830 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n616), .Z(n228) );
  MUX2_X1 U831 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n617), .Z(n229) );
  MUX2_X1 U832 ( .A(n229), .B(n228), .S(n610), .Z(n595) );
  MUX2_X1 U833 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n617), .Z(n596) );
  MUX2_X1 U834 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n614), .Z(n597) );
  MUX2_X1 U835 ( .A(n597), .B(n596), .S(n612), .Z(n598) );
  MUX2_X1 U836 ( .A(n598), .B(n595), .S(n608), .Z(n599) );
  MUX2_X1 U837 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n614), .Z(n600) );
  MUX2_X1 U838 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n617), .Z(n601) );
  MUX2_X1 U839 ( .A(n601), .B(n600), .S(n610), .Z(n602) );
  MUX2_X1 U840 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n618), .Z(n603) );
  MUX2_X1 U841 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n615), .Z(n604) );
  MUX2_X1 U842 ( .A(n604), .B(n603), .S(n610), .Z(n605) );
  MUX2_X1 U843 ( .A(n605), .B(n602), .S(n609), .Z(n606) );
  MUX2_X1 U844 ( .A(n606), .B(n599), .S(N13), .Z(n607) );
  MUX2_X1 U845 ( .A(n607), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U846 ( .A(N11), .Z(n610) );
  INV_X1 U847 ( .A(N10), .ZN(n619) );
  INV_X1 U848 ( .A(N11), .ZN(n620) );
  INV_X1 U849 ( .A(data_in[0]), .ZN(n621) );
  INV_X1 U850 ( .A(data_in[1]), .ZN(n622) );
  INV_X1 U851 ( .A(data_in[2]), .ZN(n623) );
  INV_X1 U852 ( .A(data_in[3]), .ZN(n624) );
  INV_X1 U853 ( .A(data_in[4]), .ZN(n625) );
  INV_X1 U854 ( .A(data_in[5]), .ZN(n626) );
  INV_X1 U855 ( .A(data_in[6]), .ZN(n627) );
  INV_X1 U856 ( .A(data_in[7]), .ZN(n628) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_19 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n630), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n631), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n632), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n633), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n634), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n635), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n636), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n637), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n638), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n639), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n640), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n641), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n642), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n643), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n644), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n645), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n646), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n647), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n648), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n649), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n650), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n651), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n652), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n653), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n654), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n655), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n656), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n657), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n658), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n659), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n660), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n661), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n662), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n663), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n664), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n665), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n666), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n667), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n668), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n669), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n670), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n671), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n672), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n673), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n674), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n675), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n676), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n677), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n678), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n679), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n680), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n681), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n682), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n683), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n684), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n685), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n686), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n687), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n688), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n689), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n690), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n691), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n692), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n693), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n694), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n695), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n696), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n697), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n698), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n699), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n700), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n701), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n702), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n703), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n704), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n705), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n706), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n707), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n708), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n709), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n710), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n711), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n712), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n713), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n714), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n715), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n716), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n717), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n718), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n719), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n720), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n721), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n722), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n723), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n724), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n725), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n726), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n727), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n728), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n729), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n730), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n731), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n732), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n733), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n734), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n735), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n736), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n737), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n738), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n739), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n740), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n741), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n742), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n743), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n744), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n745), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n746), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n747), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n748), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n749), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n750), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n751), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n752), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n753), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n754), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n755), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n756), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n757), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n758), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n759), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n760), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n761), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n762), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n763), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n764), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n765), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n766), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n767), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n768), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n769), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n770), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n771), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n772), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n773), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n774), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n775), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n776), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n777), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n778), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n779), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n780), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n781), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n782), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n783), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n784), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n785), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n786), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n787), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n788), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n789), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n790), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n791), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n792), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n793), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n794), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n795), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n796), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n797), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n798), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n799), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n800), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n801), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n802), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n803), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n804), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n805), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n806), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n807), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n808), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n809), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n810), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n811), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n812), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n813), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n814), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n815), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n816), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n817), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n818), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n819), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n820), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n821), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n849), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n850), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n851), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n852), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n853), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n854), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n855), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n856), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n857), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n858), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n859), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n860), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n861), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n862), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n863), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n864), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n865), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n866), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n867), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n868), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n869), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n870), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n871), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n872), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n873), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n874), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n875), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n876), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n877), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n878), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n879), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n880), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n881), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n882), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n883), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n884), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n885), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n886), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n887), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n888), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n889), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n890), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n891), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n892), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n893), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n894), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n895), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n896), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n897), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n898), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n899), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n900), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n901), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n902), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n903), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n904), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n905), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n906), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n907), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n908), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n909), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n910), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n911), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n912), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n619), .Z(n613) );
  INV_X2 U4 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U5 ( .A(n619), .Z(n617) );
  BUF_X1 U6 ( .A(n619), .Z(n618) );
  BUF_X1 U7 ( .A(n619), .Z(n615) );
  BUF_X1 U8 ( .A(n619), .Z(n614) );
  BUF_X1 U9 ( .A(n619), .Z(n616) );
  BUF_X1 U10 ( .A(N11), .Z(n611) );
  BUF_X1 U11 ( .A(N11), .Z(n612) );
  BUF_X1 U12 ( .A(N10), .Z(n619) );
  NOR3_X1 U13 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1204) );
  NOR3_X1 U14 ( .A1(N11), .A2(N12), .A3(n620), .ZN(n1193) );
  NOR3_X1 U15 ( .A1(N10), .A2(N12), .A3(n621), .ZN(n1183) );
  NOR3_X1 U16 ( .A1(n620), .A2(N12), .A3(n621), .ZN(n1173) );
  INV_X1 U17 ( .A(n1130), .ZN(n845) );
  INV_X1 U18 ( .A(n1120), .ZN(n844) );
  INV_X1 U19 ( .A(n1111), .ZN(n843) );
  INV_X1 U20 ( .A(n1102), .ZN(n842) );
  INV_X1 U21 ( .A(n1057), .ZN(n837) );
  INV_X1 U22 ( .A(n1047), .ZN(n836) );
  INV_X1 U23 ( .A(n1038), .ZN(n835) );
  INV_X1 U24 ( .A(n1029), .ZN(n834) );
  INV_X1 U25 ( .A(n984), .ZN(n829) );
  INV_X1 U26 ( .A(n974), .ZN(n828) );
  INV_X1 U27 ( .A(n965), .ZN(n827) );
  INV_X1 U28 ( .A(n956), .ZN(n826) );
  INV_X1 U29 ( .A(n947), .ZN(n825) );
  INV_X1 U30 ( .A(n938), .ZN(n824) );
  INV_X1 U31 ( .A(n929), .ZN(n823) );
  INV_X1 U32 ( .A(n920), .ZN(n822) );
  INV_X1 U33 ( .A(n1093), .ZN(n841) );
  INV_X1 U34 ( .A(n1084), .ZN(n840) );
  INV_X1 U35 ( .A(n1075), .ZN(n839) );
  INV_X1 U36 ( .A(n1066), .ZN(n838) );
  INV_X1 U37 ( .A(n1020), .ZN(n833) );
  INV_X1 U38 ( .A(n1011), .ZN(n832) );
  INV_X1 U39 ( .A(n1002), .ZN(n831) );
  INV_X1 U40 ( .A(n993), .ZN(n830) );
  BUF_X1 U41 ( .A(N12), .Z(n608) );
  BUF_X1 U42 ( .A(N12), .Z(n609) );
  INV_X1 U43 ( .A(N13), .ZN(n847) );
  AND3_X1 U44 ( .A1(n620), .A2(n621), .A3(N12), .ZN(n1163) );
  AND3_X1 U45 ( .A1(N10), .A2(n621), .A3(N12), .ZN(n1153) );
  AND3_X1 U46 ( .A1(N11), .A2(n620), .A3(N12), .ZN(n1143) );
  AND3_X1 U47 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1133) );
  INV_X1 U48 ( .A(N14), .ZN(n848) );
  NAND2_X1 U49 ( .A1(n1193), .A2(n1203), .ZN(n1202) );
  NAND2_X1 U50 ( .A1(n1183), .A2(n1203), .ZN(n1192) );
  NAND2_X1 U51 ( .A1(n1173), .A2(n1203), .ZN(n1182) );
  NAND2_X1 U52 ( .A1(n1163), .A2(n1203), .ZN(n1172) );
  NAND2_X1 U53 ( .A1(n1153), .A2(n1203), .ZN(n1162) );
  NAND2_X1 U54 ( .A1(n1143), .A2(n1203), .ZN(n1152) );
  NAND2_X1 U55 ( .A1(n1133), .A2(n1203), .ZN(n1142) );
  NAND2_X1 U56 ( .A1(n1204), .A2(n1203), .ZN(n1213) );
  NAND2_X1 U57 ( .A1(n1122), .A2(n1204), .ZN(n1130) );
  NAND2_X1 U58 ( .A1(n1122), .A2(n1193), .ZN(n1120) );
  NAND2_X1 U59 ( .A1(n1122), .A2(n1183), .ZN(n1111) );
  NAND2_X1 U60 ( .A1(n1122), .A2(n1173), .ZN(n1102) );
  NAND2_X1 U61 ( .A1(n1049), .A2(n1204), .ZN(n1057) );
  NAND2_X1 U62 ( .A1(n1049), .A2(n1193), .ZN(n1047) );
  NAND2_X1 U63 ( .A1(n1049), .A2(n1183), .ZN(n1038) );
  NAND2_X1 U64 ( .A1(n1049), .A2(n1173), .ZN(n1029) );
  NAND2_X1 U65 ( .A1(n976), .A2(n1204), .ZN(n984) );
  NAND2_X1 U66 ( .A1(n976), .A2(n1193), .ZN(n974) );
  NAND2_X1 U67 ( .A1(n976), .A2(n1183), .ZN(n965) );
  NAND2_X1 U68 ( .A1(n976), .A2(n1173), .ZN(n956) );
  NAND2_X1 U69 ( .A1(n1122), .A2(n1163), .ZN(n1093) );
  NAND2_X1 U70 ( .A1(n1122), .A2(n1153), .ZN(n1084) );
  NAND2_X1 U71 ( .A1(n1122), .A2(n1143), .ZN(n1075) );
  NAND2_X1 U72 ( .A1(n1122), .A2(n1133), .ZN(n1066) );
  NAND2_X1 U73 ( .A1(n1049), .A2(n1163), .ZN(n1020) );
  NAND2_X1 U74 ( .A1(n1049), .A2(n1153), .ZN(n1011) );
  NAND2_X1 U75 ( .A1(n1049), .A2(n1143), .ZN(n1002) );
  NAND2_X1 U76 ( .A1(n1049), .A2(n1133), .ZN(n993) );
  NAND2_X1 U77 ( .A1(n976), .A2(n1163), .ZN(n947) );
  NAND2_X1 U78 ( .A1(n976), .A2(n1153), .ZN(n938) );
  NAND2_X1 U79 ( .A1(n976), .A2(n1143), .ZN(n929) );
  NAND2_X1 U80 ( .A1(n976), .A2(n1133), .ZN(n920) );
  AND3_X1 U81 ( .A1(n847), .A2(n848), .A3(n1132), .ZN(n1203) );
  AND3_X1 U82 ( .A1(N13), .A2(n1132), .A3(N14), .ZN(n976) );
  AND3_X1 U83 ( .A1(n1132), .A2(n848), .A3(N13), .ZN(n1122) );
  AND3_X1 U84 ( .A1(n1132), .A2(n847), .A3(N14), .ZN(n1049) );
  NOR2_X1 U85 ( .A1(n846), .A2(addr[5]), .ZN(n1132) );
  INV_X1 U86 ( .A(wr_en), .ZN(n846) );
  OAI21_X1 U87 ( .B1(n622), .B2(n1172), .A(n1171), .ZN(n880) );
  NAND2_X1 U88 ( .A1(\mem[4][0] ), .A2(n1172), .ZN(n1171) );
  OAI21_X1 U89 ( .B1(n623), .B2(n1172), .A(n1170), .ZN(n879) );
  NAND2_X1 U90 ( .A1(\mem[4][1] ), .A2(n1172), .ZN(n1170) );
  OAI21_X1 U91 ( .B1(n624), .B2(n1172), .A(n1169), .ZN(n878) );
  NAND2_X1 U92 ( .A1(\mem[4][2] ), .A2(n1172), .ZN(n1169) );
  OAI21_X1 U93 ( .B1(n625), .B2(n1172), .A(n1168), .ZN(n877) );
  NAND2_X1 U94 ( .A1(\mem[4][3] ), .A2(n1172), .ZN(n1168) );
  OAI21_X1 U95 ( .B1(n626), .B2(n1172), .A(n1167), .ZN(n876) );
  NAND2_X1 U96 ( .A1(\mem[4][4] ), .A2(n1172), .ZN(n1167) );
  OAI21_X1 U97 ( .B1(n627), .B2(n1172), .A(n1166), .ZN(n875) );
  NAND2_X1 U98 ( .A1(\mem[4][5] ), .A2(n1172), .ZN(n1166) );
  OAI21_X1 U99 ( .B1(n628), .B2(n1172), .A(n1165), .ZN(n874) );
  NAND2_X1 U100 ( .A1(\mem[4][6] ), .A2(n1172), .ZN(n1165) );
  OAI21_X1 U101 ( .B1(n629), .B2(n1172), .A(n1164), .ZN(n873) );
  NAND2_X1 U102 ( .A1(\mem[4][7] ), .A2(n1172), .ZN(n1164) );
  OAI21_X1 U103 ( .B1(n622), .B2(n1152), .A(n1151), .ZN(n864) );
  NAND2_X1 U104 ( .A1(\mem[6][0] ), .A2(n1152), .ZN(n1151) );
  OAI21_X1 U105 ( .B1(n623), .B2(n1152), .A(n1150), .ZN(n863) );
  NAND2_X1 U106 ( .A1(\mem[6][1] ), .A2(n1152), .ZN(n1150) );
  OAI21_X1 U107 ( .B1(n624), .B2(n1152), .A(n1149), .ZN(n862) );
  NAND2_X1 U108 ( .A1(\mem[6][2] ), .A2(n1152), .ZN(n1149) );
  OAI21_X1 U109 ( .B1(n625), .B2(n1152), .A(n1148), .ZN(n861) );
  NAND2_X1 U110 ( .A1(\mem[6][3] ), .A2(n1152), .ZN(n1148) );
  OAI21_X1 U111 ( .B1(n626), .B2(n1152), .A(n1147), .ZN(n860) );
  NAND2_X1 U112 ( .A1(\mem[6][4] ), .A2(n1152), .ZN(n1147) );
  OAI21_X1 U113 ( .B1(n627), .B2(n1152), .A(n1146), .ZN(n859) );
  NAND2_X1 U114 ( .A1(\mem[6][5] ), .A2(n1152), .ZN(n1146) );
  OAI21_X1 U115 ( .B1(n628), .B2(n1152), .A(n1145), .ZN(n858) );
  NAND2_X1 U116 ( .A1(\mem[6][6] ), .A2(n1152), .ZN(n1145) );
  OAI21_X1 U117 ( .B1(n629), .B2(n1152), .A(n1144), .ZN(n857) );
  NAND2_X1 U118 ( .A1(\mem[6][7] ), .A2(n1152), .ZN(n1144) );
  OAI21_X1 U119 ( .B1(n622), .B2(n1142), .A(n1141), .ZN(n856) );
  NAND2_X1 U120 ( .A1(\mem[7][0] ), .A2(n1142), .ZN(n1141) );
  OAI21_X1 U121 ( .B1(n623), .B2(n1142), .A(n1140), .ZN(n855) );
  NAND2_X1 U122 ( .A1(\mem[7][1] ), .A2(n1142), .ZN(n1140) );
  OAI21_X1 U123 ( .B1(n624), .B2(n1142), .A(n1139), .ZN(n854) );
  NAND2_X1 U124 ( .A1(\mem[7][2] ), .A2(n1142), .ZN(n1139) );
  OAI21_X1 U125 ( .B1(n625), .B2(n1142), .A(n1138), .ZN(n853) );
  NAND2_X1 U126 ( .A1(\mem[7][3] ), .A2(n1142), .ZN(n1138) );
  OAI21_X1 U127 ( .B1(n626), .B2(n1142), .A(n1137), .ZN(n852) );
  NAND2_X1 U128 ( .A1(\mem[7][4] ), .A2(n1142), .ZN(n1137) );
  OAI21_X1 U129 ( .B1(n627), .B2(n1142), .A(n1136), .ZN(n851) );
  NAND2_X1 U130 ( .A1(\mem[7][5] ), .A2(n1142), .ZN(n1136) );
  OAI21_X1 U131 ( .B1(n628), .B2(n1142), .A(n1135), .ZN(n850) );
  NAND2_X1 U132 ( .A1(\mem[7][6] ), .A2(n1142), .ZN(n1135) );
  OAI21_X1 U133 ( .B1(n629), .B2(n1142), .A(n1134), .ZN(n849) );
  NAND2_X1 U134 ( .A1(\mem[7][7] ), .A2(n1142), .ZN(n1134) );
  OAI21_X1 U135 ( .B1(n622), .B2(n1202), .A(n1201), .ZN(n904) );
  NAND2_X1 U136 ( .A1(\mem[1][0] ), .A2(n1202), .ZN(n1201) );
  OAI21_X1 U137 ( .B1(n623), .B2(n1202), .A(n1200), .ZN(n903) );
  NAND2_X1 U138 ( .A1(\mem[1][1] ), .A2(n1202), .ZN(n1200) );
  OAI21_X1 U139 ( .B1(n624), .B2(n1202), .A(n1199), .ZN(n902) );
  NAND2_X1 U140 ( .A1(\mem[1][2] ), .A2(n1202), .ZN(n1199) );
  OAI21_X1 U141 ( .B1(n625), .B2(n1202), .A(n1198), .ZN(n901) );
  NAND2_X1 U142 ( .A1(\mem[1][3] ), .A2(n1202), .ZN(n1198) );
  OAI21_X1 U143 ( .B1(n626), .B2(n1202), .A(n1197), .ZN(n900) );
  NAND2_X1 U144 ( .A1(\mem[1][4] ), .A2(n1202), .ZN(n1197) );
  OAI21_X1 U145 ( .B1(n627), .B2(n1202), .A(n1196), .ZN(n899) );
  NAND2_X1 U146 ( .A1(\mem[1][5] ), .A2(n1202), .ZN(n1196) );
  OAI21_X1 U147 ( .B1(n628), .B2(n1202), .A(n1195), .ZN(n898) );
  NAND2_X1 U148 ( .A1(\mem[1][6] ), .A2(n1202), .ZN(n1195) );
  OAI21_X1 U149 ( .B1(n629), .B2(n1202), .A(n1194), .ZN(n897) );
  NAND2_X1 U150 ( .A1(\mem[1][7] ), .A2(n1202), .ZN(n1194) );
  OAI21_X1 U151 ( .B1(n622), .B2(n1192), .A(n1191), .ZN(n896) );
  NAND2_X1 U152 ( .A1(\mem[2][0] ), .A2(n1192), .ZN(n1191) );
  OAI21_X1 U153 ( .B1(n623), .B2(n1192), .A(n1190), .ZN(n895) );
  NAND2_X1 U154 ( .A1(\mem[2][1] ), .A2(n1192), .ZN(n1190) );
  OAI21_X1 U155 ( .B1(n624), .B2(n1192), .A(n1189), .ZN(n894) );
  NAND2_X1 U156 ( .A1(\mem[2][2] ), .A2(n1192), .ZN(n1189) );
  OAI21_X1 U157 ( .B1(n625), .B2(n1192), .A(n1188), .ZN(n893) );
  NAND2_X1 U158 ( .A1(\mem[2][3] ), .A2(n1192), .ZN(n1188) );
  OAI21_X1 U159 ( .B1(n626), .B2(n1192), .A(n1187), .ZN(n892) );
  NAND2_X1 U160 ( .A1(\mem[2][4] ), .A2(n1192), .ZN(n1187) );
  OAI21_X1 U161 ( .B1(n627), .B2(n1192), .A(n1186), .ZN(n891) );
  NAND2_X1 U162 ( .A1(\mem[2][5] ), .A2(n1192), .ZN(n1186) );
  OAI21_X1 U163 ( .B1(n628), .B2(n1192), .A(n1185), .ZN(n890) );
  NAND2_X1 U164 ( .A1(\mem[2][6] ), .A2(n1192), .ZN(n1185) );
  OAI21_X1 U165 ( .B1(n629), .B2(n1192), .A(n1184), .ZN(n889) );
  NAND2_X1 U166 ( .A1(\mem[2][7] ), .A2(n1192), .ZN(n1184) );
  OAI21_X1 U167 ( .B1(n622), .B2(n1182), .A(n1181), .ZN(n888) );
  NAND2_X1 U168 ( .A1(\mem[3][0] ), .A2(n1182), .ZN(n1181) );
  OAI21_X1 U169 ( .B1(n623), .B2(n1182), .A(n1180), .ZN(n887) );
  NAND2_X1 U170 ( .A1(\mem[3][1] ), .A2(n1182), .ZN(n1180) );
  OAI21_X1 U171 ( .B1(n624), .B2(n1182), .A(n1179), .ZN(n886) );
  NAND2_X1 U172 ( .A1(\mem[3][2] ), .A2(n1182), .ZN(n1179) );
  OAI21_X1 U173 ( .B1(n625), .B2(n1182), .A(n1178), .ZN(n885) );
  NAND2_X1 U174 ( .A1(\mem[3][3] ), .A2(n1182), .ZN(n1178) );
  OAI21_X1 U175 ( .B1(n626), .B2(n1182), .A(n1177), .ZN(n884) );
  NAND2_X1 U176 ( .A1(\mem[3][4] ), .A2(n1182), .ZN(n1177) );
  OAI21_X1 U177 ( .B1(n627), .B2(n1182), .A(n1176), .ZN(n883) );
  NAND2_X1 U178 ( .A1(\mem[3][5] ), .A2(n1182), .ZN(n1176) );
  OAI21_X1 U179 ( .B1(n628), .B2(n1182), .A(n1175), .ZN(n882) );
  NAND2_X1 U180 ( .A1(\mem[3][6] ), .A2(n1182), .ZN(n1175) );
  OAI21_X1 U181 ( .B1(n629), .B2(n1182), .A(n1174), .ZN(n881) );
  NAND2_X1 U182 ( .A1(\mem[3][7] ), .A2(n1182), .ZN(n1174) );
  OAI21_X1 U183 ( .B1(n622), .B2(n1162), .A(n1161), .ZN(n872) );
  NAND2_X1 U184 ( .A1(\mem[5][0] ), .A2(n1162), .ZN(n1161) );
  OAI21_X1 U185 ( .B1(n623), .B2(n1162), .A(n1160), .ZN(n871) );
  NAND2_X1 U186 ( .A1(\mem[5][1] ), .A2(n1162), .ZN(n1160) );
  OAI21_X1 U187 ( .B1(n624), .B2(n1162), .A(n1159), .ZN(n870) );
  NAND2_X1 U188 ( .A1(\mem[5][2] ), .A2(n1162), .ZN(n1159) );
  OAI21_X1 U189 ( .B1(n625), .B2(n1162), .A(n1158), .ZN(n869) );
  NAND2_X1 U190 ( .A1(\mem[5][3] ), .A2(n1162), .ZN(n1158) );
  OAI21_X1 U191 ( .B1(n626), .B2(n1162), .A(n1157), .ZN(n868) );
  NAND2_X1 U192 ( .A1(\mem[5][4] ), .A2(n1162), .ZN(n1157) );
  OAI21_X1 U193 ( .B1(n627), .B2(n1162), .A(n1156), .ZN(n867) );
  NAND2_X1 U194 ( .A1(\mem[5][5] ), .A2(n1162), .ZN(n1156) );
  OAI21_X1 U195 ( .B1(n628), .B2(n1162), .A(n1155), .ZN(n866) );
  NAND2_X1 U196 ( .A1(\mem[5][6] ), .A2(n1162), .ZN(n1155) );
  OAI21_X1 U197 ( .B1(n629), .B2(n1162), .A(n1154), .ZN(n865) );
  NAND2_X1 U198 ( .A1(\mem[5][7] ), .A2(n1162), .ZN(n1154) );
  OAI21_X1 U199 ( .B1(n1213), .B2(n622), .A(n1212), .ZN(n912) );
  NAND2_X1 U200 ( .A1(\mem[0][0] ), .A2(n1213), .ZN(n1212) );
  OAI21_X1 U201 ( .B1(n1213), .B2(n623), .A(n1211), .ZN(n911) );
  NAND2_X1 U202 ( .A1(\mem[0][1] ), .A2(n1213), .ZN(n1211) );
  OAI21_X1 U203 ( .B1(n1213), .B2(n624), .A(n1210), .ZN(n910) );
  NAND2_X1 U204 ( .A1(\mem[0][2] ), .A2(n1213), .ZN(n1210) );
  OAI21_X1 U205 ( .B1(n1213), .B2(n625), .A(n1209), .ZN(n909) );
  NAND2_X1 U206 ( .A1(\mem[0][3] ), .A2(n1213), .ZN(n1209) );
  OAI21_X1 U207 ( .B1(n1213), .B2(n626), .A(n1208), .ZN(n908) );
  NAND2_X1 U208 ( .A1(\mem[0][4] ), .A2(n1213), .ZN(n1208) );
  OAI21_X1 U209 ( .B1(n1213), .B2(n627), .A(n1207), .ZN(n907) );
  NAND2_X1 U210 ( .A1(\mem[0][5] ), .A2(n1213), .ZN(n1207) );
  OAI21_X1 U211 ( .B1(n1213), .B2(n628), .A(n1206), .ZN(n906) );
  NAND2_X1 U212 ( .A1(\mem[0][6] ), .A2(n1213), .ZN(n1206) );
  OAI21_X1 U213 ( .B1(n1213), .B2(n629), .A(n1205), .ZN(n905) );
  NAND2_X1 U214 ( .A1(\mem[0][7] ), .A2(n1213), .ZN(n1205) );
  INV_X1 U215 ( .A(n1131), .ZN(n821) );
  AOI22_X1 U216 ( .A1(data_in[0]), .A2(n845), .B1(n1130), .B2(\mem[8][0] ), 
        .ZN(n1131) );
  INV_X1 U217 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U218 ( .A1(data_in[1]), .A2(n845), .B1(n1130), .B2(\mem[8][1] ), 
        .ZN(n1129) );
  INV_X1 U219 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U220 ( .A1(data_in[2]), .A2(n845), .B1(n1130), .B2(\mem[8][2] ), 
        .ZN(n1128) );
  INV_X1 U221 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U222 ( .A1(data_in[3]), .A2(n845), .B1(n1130), .B2(\mem[8][3] ), 
        .ZN(n1127) );
  INV_X1 U223 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U224 ( .A1(data_in[4]), .A2(n845), .B1(n1130), .B2(\mem[8][4] ), 
        .ZN(n1126) );
  INV_X1 U225 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U226 ( .A1(data_in[5]), .A2(n845), .B1(n1130), .B2(\mem[8][5] ), 
        .ZN(n1125) );
  INV_X1 U227 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U228 ( .A1(data_in[6]), .A2(n845), .B1(n1130), .B2(\mem[8][6] ), 
        .ZN(n1124) );
  INV_X1 U229 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U230 ( .A1(data_in[7]), .A2(n845), .B1(n1130), .B2(\mem[8][7] ), 
        .ZN(n1123) );
  INV_X1 U231 ( .A(n1121), .ZN(n813) );
  AOI22_X1 U232 ( .A1(data_in[0]), .A2(n844), .B1(n1120), .B2(\mem[9][0] ), 
        .ZN(n1121) );
  INV_X1 U233 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U234 ( .A1(data_in[1]), .A2(n844), .B1(n1120), .B2(\mem[9][1] ), 
        .ZN(n1119) );
  INV_X1 U235 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U236 ( .A1(data_in[2]), .A2(n844), .B1(n1120), .B2(\mem[9][2] ), 
        .ZN(n1118) );
  INV_X1 U237 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U238 ( .A1(data_in[3]), .A2(n844), .B1(n1120), .B2(\mem[9][3] ), 
        .ZN(n1117) );
  INV_X1 U239 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U240 ( .A1(data_in[4]), .A2(n844), .B1(n1120), .B2(\mem[9][4] ), 
        .ZN(n1116) );
  INV_X1 U241 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U242 ( .A1(data_in[5]), .A2(n844), .B1(n1120), .B2(\mem[9][5] ), 
        .ZN(n1115) );
  INV_X1 U243 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U244 ( .A1(data_in[6]), .A2(n844), .B1(n1120), .B2(\mem[9][6] ), 
        .ZN(n1114) );
  INV_X1 U245 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U246 ( .A1(data_in[7]), .A2(n844), .B1(n1120), .B2(\mem[9][7] ), 
        .ZN(n1113) );
  INV_X1 U247 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U248 ( .A1(data_in[0]), .A2(n843), .B1(n1111), .B2(\mem[10][0] ), 
        .ZN(n1112) );
  INV_X1 U249 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U250 ( .A1(data_in[1]), .A2(n843), .B1(n1111), .B2(\mem[10][1] ), 
        .ZN(n1110) );
  INV_X1 U251 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U252 ( .A1(data_in[2]), .A2(n843), .B1(n1111), .B2(\mem[10][2] ), 
        .ZN(n1109) );
  INV_X1 U253 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U254 ( .A1(data_in[3]), .A2(n843), .B1(n1111), .B2(\mem[10][3] ), 
        .ZN(n1108) );
  INV_X1 U255 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U256 ( .A1(data_in[4]), .A2(n843), .B1(n1111), .B2(\mem[10][4] ), 
        .ZN(n1107) );
  INV_X1 U257 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U258 ( .A1(data_in[5]), .A2(n843), .B1(n1111), .B2(\mem[10][5] ), 
        .ZN(n1106) );
  INV_X1 U259 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U260 ( .A1(data_in[6]), .A2(n843), .B1(n1111), .B2(\mem[10][6] ), 
        .ZN(n1105) );
  INV_X1 U261 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U262 ( .A1(data_in[7]), .A2(n843), .B1(n1111), .B2(\mem[10][7] ), 
        .ZN(n1104) );
  INV_X1 U263 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U264 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[11][0] ), 
        .ZN(n1103) );
  INV_X1 U265 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U266 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[11][1] ), 
        .ZN(n1101) );
  INV_X1 U267 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U268 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[11][2] ), 
        .ZN(n1100) );
  INV_X1 U269 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U270 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[11][3] ), 
        .ZN(n1099) );
  INV_X1 U271 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U272 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[11][4] ), 
        .ZN(n1098) );
  INV_X1 U273 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U274 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[11][5] ), 
        .ZN(n1097) );
  INV_X1 U275 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U276 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[11][6] ), 
        .ZN(n1096) );
  INV_X1 U277 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U278 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[11][7] ), 
        .ZN(n1095) );
  INV_X1 U279 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U280 ( .A1(data_in[0]), .A2(n841), .B1(n1093), .B2(\mem[12][0] ), 
        .ZN(n1094) );
  INV_X1 U281 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U282 ( .A1(data_in[1]), .A2(n841), .B1(n1093), .B2(\mem[12][1] ), 
        .ZN(n1092) );
  INV_X1 U283 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U284 ( .A1(data_in[2]), .A2(n841), .B1(n1093), .B2(\mem[12][2] ), 
        .ZN(n1091) );
  INV_X1 U285 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U286 ( .A1(data_in[3]), .A2(n841), .B1(n1093), .B2(\mem[12][3] ), 
        .ZN(n1090) );
  INV_X1 U287 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U288 ( .A1(data_in[4]), .A2(n841), .B1(n1093), .B2(\mem[12][4] ), 
        .ZN(n1089) );
  INV_X1 U289 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U290 ( .A1(data_in[5]), .A2(n841), .B1(n1093), .B2(\mem[12][5] ), 
        .ZN(n1088) );
  INV_X1 U291 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U292 ( .A1(data_in[6]), .A2(n841), .B1(n1093), .B2(\mem[12][6] ), 
        .ZN(n1087) );
  INV_X1 U293 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U294 ( .A1(data_in[7]), .A2(n841), .B1(n1093), .B2(\mem[12][7] ), 
        .ZN(n1086) );
  INV_X1 U295 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U296 ( .A1(data_in[0]), .A2(n840), .B1(n1084), .B2(\mem[13][0] ), 
        .ZN(n1085) );
  INV_X1 U297 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U298 ( .A1(data_in[1]), .A2(n840), .B1(n1084), .B2(\mem[13][1] ), 
        .ZN(n1083) );
  INV_X1 U299 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U300 ( .A1(data_in[2]), .A2(n840), .B1(n1084), .B2(\mem[13][2] ), 
        .ZN(n1082) );
  INV_X1 U301 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U302 ( .A1(data_in[3]), .A2(n840), .B1(n1084), .B2(\mem[13][3] ), 
        .ZN(n1081) );
  INV_X1 U303 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U304 ( .A1(data_in[4]), .A2(n840), .B1(n1084), .B2(\mem[13][4] ), 
        .ZN(n1080) );
  INV_X1 U305 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U306 ( .A1(data_in[5]), .A2(n840), .B1(n1084), .B2(\mem[13][5] ), 
        .ZN(n1079) );
  INV_X1 U307 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U308 ( .A1(data_in[6]), .A2(n840), .B1(n1084), .B2(\mem[13][6] ), 
        .ZN(n1078) );
  INV_X1 U309 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U310 ( .A1(data_in[7]), .A2(n840), .B1(n1084), .B2(\mem[13][7] ), 
        .ZN(n1077) );
  INV_X1 U311 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U312 ( .A1(data_in[0]), .A2(n839), .B1(n1075), .B2(\mem[14][0] ), 
        .ZN(n1076) );
  INV_X1 U313 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U314 ( .A1(data_in[1]), .A2(n839), .B1(n1075), .B2(\mem[14][1] ), 
        .ZN(n1074) );
  INV_X1 U315 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U316 ( .A1(data_in[2]), .A2(n839), .B1(n1075), .B2(\mem[14][2] ), 
        .ZN(n1073) );
  INV_X1 U317 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U318 ( .A1(data_in[3]), .A2(n839), .B1(n1075), .B2(\mem[14][3] ), 
        .ZN(n1072) );
  INV_X1 U319 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U320 ( .A1(data_in[4]), .A2(n839), .B1(n1075), .B2(\mem[14][4] ), 
        .ZN(n1071) );
  INV_X1 U321 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U322 ( .A1(data_in[5]), .A2(n839), .B1(n1075), .B2(\mem[14][5] ), 
        .ZN(n1070) );
  INV_X1 U323 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U324 ( .A1(data_in[6]), .A2(n839), .B1(n1075), .B2(\mem[14][6] ), 
        .ZN(n1069) );
  INV_X1 U325 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U326 ( .A1(data_in[7]), .A2(n839), .B1(n1075), .B2(\mem[14][7] ), 
        .ZN(n1068) );
  INV_X1 U327 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U328 ( .A1(data_in[0]), .A2(n838), .B1(n1066), .B2(\mem[15][0] ), 
        .ZN(n1067) );
  INV_X1 U329 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U330 ( .A1(data_in[1]), .A2(n838), .B1(n1066), .B2(\mem[15][1] ), 
        .ZN(n1065) );
  INV_X1 U331 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U332 ( .A1(data_in[2]), .A2(n838), .B1(n1066), .B2(\mem[15][2] ), 
        .ZN(n1064) );
  INV_X1 U333 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U334 ( .A1(data_in[3]), .A2(n838), .B1(n1066), .B2(\mem[15][3] ), 
        .ZN(n1063) );
  INV_X1 U335 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U336 ( .A1(data_in[4]), .A2(n838), .B1(n1066), .B2(\mem[15][4] ), 
        .ZN(n1062) );
  INV_X1 U337 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U338 ( .A1(data_in[5]), .A2(n838), .B1(n1066), .B2(\mem[15][5] ), 
        .ZN(n1061) );
  INV_X1 U339 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U340 ( .A1(data_in[6]), .A2(n838), .B1(n1066), .B2(\mem[15][6] ), 
        .ZN(n1060) );
  INV_X1 U341 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U342 ( .A1(data_in[7]), .A2(n838), .B1(n1066), .B2(\mem[15][7] ), 
        .ZN(n1059) );
  INV_X1 U343 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U344 ( .A1(data_in[0]), .A2(n837), .B1(n1057), .B2(\mem[16][0] ), 
        .ZN(n1058) );
  INV_X1 U345 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U346 ( .A1(data_in[1]), .A2(n837), .B1(n1057), .B2(\mem[16][1] ), 
        .ZN(n1056) );
  INV_X1 U347 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U348 ( .A1(data_in[2]), .A2(n837), .B1(n1057), .B2(\mem[16][2] ), 
        .ZN(n1055) );
  INV_X1 U349 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U350 ( .A1(data_in[3]), .A2(n837), .B1(n1057), .B2(\mem[16][3] ), 
        .ZN(n1054) );
  INV_X1 U351 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U352 ( .A1(data_in[4]), .A2(n837), .B1(n1057), .B2(\mem[16][4] ), 
        .ZN(n1053) );
  INV_X1 U353 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U354 ( .A1(data_in[5]), .A2(n837), .B1(n1057), .B2(\mem[16][5] ), 
        .ZN(n1052) );
  INV_X1 U355 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U356 ( .A1(data_in[6]), .A2(n837), .B1(n1057), .B2(\mem[16][6] ), 
        .ZN(n1051) );
  INV_X1 U357 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U358 ( .A1(data_in[7]), .A2(n837), .B1(n1057), .B2(\mem[16][7] ), 
        .ZN(n1050) );
  INV_X1 U359 ( .A(n1048), .ZN(n749) );
  AOI22_X1 U360 ( .A1(data_in[0]), .A2(n836), .B1(n1047), .B2(\mem[17][0] ), 
        .ZN(n1048) );
  INV_X1 U361 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U362 ( .A1(data_in[1]), .A2(n836), .B1(n1047), .B2(\mem[17][1] ), 
        .ZN(n1046) );
  INV_X1 U363 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U364 ( .A1(data_in[2]), .A2(n836), .B1(n1047), .B2(\mem[17][2] ), 
        .ZN(n1045) );
  INV_X1 U365 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U366 ( .A1(data_in[3]), .A2(n836), .B1(n1047), .B2(\mem[17][3] ), 
        .ZN(n1044) );
  INV_X1 U367 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U368 ( .A1(data_in[4]), .A2(n836), .B1(n1047), .B2(\mem[17][4] ), 
        .ZN(n1043) );
  INV_X1 U369 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U370 ( .A1(data_in[5]), .A2(n836), .B1(n1047), .B2(\mem[17][5] ), 
        .ZN(n1042) );
  INV_X1 U371 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U372 ( .A1(data_in[6]), .A2(n836), .B1(n1047), .B2(\mem[17][6] ), 
        .ZN(n1041) );
  INV_X1 U373 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U374 ( .A1(data_in[7]), .A2(n836), .B1(n1047), .B2(\mem[17][7] ), 
        .ZN(n1040) );
  INV_X1 U375 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U376 ( .A1(data_in[0]), .A2(n835), .B1(n1038), .B2(\mem[18][0] ), 
        .ZN(n1039) );
  INV_X1 U377 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U378 ( .A1(data_in[1]), .A2(n835), .B1(n1038), .B2(\mem[18][1] ), 
        .ZN(n1037) );
  INV_X1 U379 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U380 ( .A1(data_in[2]), .A2(n835), .B1(n1038), .B2(\mem[18][2] ), 
        .ZN(n1036) );
  INV_X1 U381 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U382 ( .A1(data_in[3]), .A2(n835), .B1(n1038), .B2(\mem[18][3] ), 
        .ZN(n1035) );
  INV_X1 U383 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U384 ( .A1(data_in[4]), .A2(n835), .B1(n1038), .B2(\mem[18][4] ), 
        .ZN(n1034) );
  INV_X1 U385 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U386 ( .A1(data_in[5]), .A2(n835), .B1(n1038), .B2(\mem[18][5] ), 
        .ZN(n1033) );
  INV_X1 U387 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U388 ( .A1(data_in[6]), .A2(n835), .B1(n1038), .B2(\mem[18][6] ), 
        .ZN(n1032) );
  INV_X1 U389 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U390 ( .A1(data_in[7]), .A2(n835), .B1(n1038), .B2(\mem[18][7] ), 
        .ZN(n1031) );
  INV_X1 U391 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U392 ( .A1(data_in[0]), .A2(n834), .B1(n1029), .B2(\mem[19][0] ), 
        .ZN(n1030) );
  INV_X1 U393 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U394 ( .A1(data_in[1]), .A2(n834), .B1(n1029), .B2(\mem[19][1] ), 
        .ZN(n1028) );
  INV_X1 U395 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U396 ( .A1(data_in[2]), .A2(n834), .B1(n1029), .B2(\mem[19][2] ), 
        .ZN(n1027) );
  INV_X1 U397 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U398 ( .A1(data_in[3]), .A2(n834), .B1(n1029), .B2(\mem[19][3] ), 
        .ZN(n1026) );
  INV_X1 U399 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U400 ( .A1(data_in[4]), .A2(n834), .B1(n1029), .B2(\mem[19][4] ), 
        .ZN(n1025) );
  INV_X1 U401 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U402 ( .A1(data_in[5]), .A2(n834), .B1(n1029), .B2(\mem[19][5] ), 
        .ZN(n1024) );
  INV_X1 U403 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U404 ( .A1(data_in[6]), .A2(n834), .B1(n1029), .B2(\mem[19][6] ), 
        .ZN(n1023) );
  INV_X1 U405 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U406 ( .A1(data_in[7]), .A2(n834), .B1(n1029), .B2(\mem[19][7] ), 
        .ZN(n1022) );
  INV_X1 U407 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U408 ( .A1(data_in[0]), .A2(n833), .B1(n1020), .B2(\mem[20][0] ), 
        .ZN(n1021) );
  INV_X1 U409 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U410 ( .A1(data_in[1]), .A2(n833), .B1(n1020), .B2(\mem[20][1] ), 
        .ZN(n1019) );
  INV_X1 U411 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U412 ( .A1(data_in[2]), .A2(n833), .B1(n1020), .B2(\mem[20][2] ), 
        .ZN(n1018) );
  INV_X1 U413 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U414 ( .A1(data_in[3]), .A2(n833), .B1(n1020), .B2(\mem[20][3] ), 
        .ZN(n1017) );
  INV_X1 U415 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U416 ( .A1(data_in[4]), .A2(n833), .B1(n1020), .B2(\mem[20][4] ), 
        .ZN(n1016) );
  INV_X1 U417 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U418 ( .A1(data_in[5]), .A2(n833), .B1(n1020), .B2(\mem[20][5] ), 
        .ZN(n1015) );
  INV_X1 U419 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U420 ( .A1(data_in[6]), .A2(n833), .B1(n1020), .B2(\mem[20][6] ), 
        .ZN(n1014) );
  INV_X1 U421 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U422 ( .A1(data_in[7]), .A2(n833), .B1(n1020), .B2(\mem[20][7] ), 
        .ZN(n1013) );
  INV_X1 U423 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U424 ( .A1(data_in[0]), .A2(n832), .B1(n1011), .B2(\mem[21][0] ), 
        .ZN(n1012) );
  INV_X1 U425 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U426 ( .A1(data_in[1]), .A2(n832), .B1(n1011), .B2(\mem[21][1] ), 
        .ZN(n1010) );
  INV_X1 U427 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U428 ( .A1(data_in[2]), .A2(n832), .B1(n1011), .B2(\mem[21][2] ), 
        .ZN(n1009) );
  INV_X1 U429 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U430 ( .A1(data_in[3]), .A2(n832), .B1(n1011), .B2(\mem[21][3] ), 
        .ZN(n1008) );
  INV_X1 U431 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U432 ( .A1(data_in[4]), .A2(n832), .B1(n1011), .B2(\mem[21][4] ), 
        .ZN(n1007) );
  INV_X1 U433 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U434 ( .A1(data_in[5]), .A2(n832), .B1(n1011), .B2(\mem[21][5] ), 
        .ZN(n1006) );
  INV_X1 U435 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U436 ( .A1(data_in[6]), .A2(n832), .B1(n1011), .B2(\mem[21][6] ), 
        .ZN(n1005) );
  INV_X1 U437 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U438 ( .A1(data_in[7]), .A2(n832), .B1(n1011), .B2(\mem[21][7] ), 
        .ZN(n1004) );
  INV_X1 U439 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U440 ( .A1(data_in[0]), .A2(n831), .B1(n1002), .B2(\mem[22][0] ), 
        .ZN(n1003) );
  INV_X1 U441 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U442 ( .A1(data_in[1]), .A2(n831), .B1(n1002), .B2(\mem[22][1] ), 
        .ZN(n1001) );
  INV_X1 U443 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U444 ( .A1(data_in[2]), .A2(n831), .B1(n1002), .B2(\mem[22][2] ), 
        .ZN(n1000) );
  INV_X1 U445 ( .A(n999), .ZN(n706) );
  AOI22_X1 U446 ( .A1(data_in[3]), .A2(n831), .B1(n1002), .B2(\mem[22][3] ), 
        .ZN(n999) );
  INV_X1 U447 ( .A(n998), .ZN(n705) );
  AOI22_X1 U448 ( .A1(data_in[4]), .A2(n831), .B1(n1002), .B2(\mem[22][4] ), 
        .ZN(n998) );
  INV_X1 U449 ( .A(n997), .ZN(n704) );
  AOI22_X1 U450 ( .A1(data_in[5]), .A2(n831), .B1(n1002), .B2(\mem[22][5] ), 
        .ZN(n997) );
  INV_X1 U451 ( .A(n996), .ZN(n703) );
  AOI22_X1 U452 ( .A1(data_in[6]), .A2(n831), .B1(n1002), .B2(\mem[22][6] ), 
        .ZN(n996) );
  INV_X1 U453 ( .A(n995), .ZN(n702) );
  AOI22_X1 U454 ( .A1(data_in[7]), .A2(n831), .B1(n1002), .B2(\mem[22][7] ), 
        .ZN(n995) );
  INV_X1 U455 ( .A(n994), .ZN(n701) );
  AOI22_X1 U456 ( .A1(data_in[0]), .A2(n830), .B1(n993), .B2(\mem[23][0] ), 
        .ZN(n994) );
  INV_X1 U457 ( .A(n992), .ZN(n700) );
  AOI22_X1 U458 ( .A1(data_in[1]), .A2(n830), .B1(n993), .B2(\mem[23][1] ), 
        .ZN(n992) );
  INV_X1 U459 ( .A(n991), .ZN(n699) );
  AOI22_X1 U460 ( .A1(data_in[2]), .A2(n830), .B1(n993), .B2(\mem[23][2] ), 
        .ZN(n991) );
  INV_X1 U461 ( .A(n990), .ZN(n698) );
  AOI22_X1 U462 ( .A1(data_in[3]), .A2(n830), .B1(n993), .B2(\mem[23][3] ), 
        .ZN(n990) );
  INV_X1 U463 ( .A(n989), .ZN(n697) );
  AOI22_X1 U464 ( .A1(data_in[4]), .A2(n830), .B1(n993), .B2(\mem[23][4] ), 
        .ZN(n989) );
  INV_X1 U465 ( .A(n988), .ZN(n696) );
  AOI22_X1 U466 ( .A1(data_in[5]), .A2(n830), .B1(n993), .B2(\mem[23][5] ), 
        .ZN(n988) );
  INV_X1 U467 ( .A(n987), .ZN(n695) );
  AOI22_X1 U468 ( .A1(data_in[6]), .A2(n830), .B1(n993), .B2(\mem[23][6] ), 
        .ZN(n987) );
  INV_X1 U469 ( .A(n986), .ZN(n694) );
  AOI22_X1 U470 ( .A1(data_in[7]), .A2(n830), .B1(n993), .B2(\mem[23][7] ), 
        .ZN(n986) );
  INV_X1 U471 ( .A(n985), .ZN(n693) );
  AOI22_X1 U472 ( .A1(data_in[0]), .A2(n829), .B1(n984), .B2(\mem[24][0] ), 
        .ZN(n985) );
  INV_X1 U473 ( .A(n983), .ZN(n692) );
  AOI22_X1 U474 ( .A1(data_in[1]), .A2(n829), .B1(n984), .B2(\mem[24][1] ), 
        .ZN(n983) );
  INV_X1 U475 ( .A(n982), .ZN(n691) );
  AOI22_X1 U476 ( .A1(data_in[2]), .A2(n829), .B1(n984), .B2(\mem[24][2] ), 
        .ZN(n982) );
  INV_X1 U477 ( .A(n981), .ZN(n690) );
  AOI22_X1 U478 ( .A1(data_in[3]), .A2(n829), .B1(n984), .B2(\mem[24][3] ), 
        .ZN(n981) );
  INV_X1 U479 ( .A(n980), .ZN(n689) );
  AOI22_X1 U480 ( .A1(data_in[4]), .A2(n829), .B1(n984), .B2(\mem[24][4] ), 
        .ZN(n980) );
  INV_X1 U481 ( .A(n979), .ZN(n688) );
  AOI22_X1 U482 ( .A1(data_in[5]), .A2(n829), .B1(n984), .B2(\mem[24][5] ), 
        .ZN(n979) );
  INV_X1 U483 ( .A(n978), .ZN(n687) );
  AOI22_X1 U484 ( .A1(data_in[6]), .A2(n829), .B1(n984), .B2(\mem[24][6] ), 
        .ZN(n978) );
  INV_X1 U485 ( .A(n977), .ZN(n686) );
  AOI22_X1 U486 ( .A1(data_in[7]), .A2(n829), .B1(n984), .B2(\mem[24][7] ), 
        .ZN(n977) );
  INV_X1 U487 ( .A(n975), .ZN(n685) );
  AOI22_X1 U488 ( .A1(data_in[0]), .A2(n828), .B1(n974), .B2(\mem[25][0] ), 
        .ZN(n975) );
  INV_X1 U489 ( .A(n973), .ZN(n684) );
  AOI22_X1 U490 ( .A1(data_in[1]), .A2(n828), .B1(n974), .B2(\mem[25][1] ), 
        .ZN(n973) );
  INV_X1 U491 ( .A(n972), .ZN(n683) );
  AOI22_X1 U492 ( .A1(data_in[2]), .A2(n828), .B1(n974), .B2(\mem[25][2] ), 
        .ZN(n972) );
  INV_X1 U493 ( .A(n971), .ZN(n682) );
  AOI22_X1 U494 ( .A1(data_in[3]), .A2(n828), .B1(n974), .B2(\mem[25][3] ), 
        .ZN(n971) );
  INV_X1 U495 ( .A(n970), .ZN(n681) );
  AOI22_X1 U496 ( .A1(data_in[4]), .A2(n828), .B1(n974), .B2(\mem[25][4] ), 
        .ZN(n970) );
  INV_X1 U497 ( .A(n969), .ZN(n680) );
  AOI22_X1 U498 ( .A1(data_in[5]), .A2(n828), .B1(n974), .B2(\mem[25][5] ), 
        .ZN(n969) );
  INV_X1 U499 ( .A(n968), .ZN(n679) );
  AOI22_X1 U500 ( .A1(data_in[6]), .A2(n828), .B1(n974), .B2(\mem[25][6] ), 
        .ZN(n968) );
  INV_X1 U501 ( .A(n967), .ZN(n678) );
  AOI22_X1 U502 ( .A1(data_in[7]), .A2(n828), .B1(n974), .B2(\mem[25][7] ), 
        .ZN(n967) );
  INV_X1 U503 ( .A(n966), .ZN(n677) );
  AOI22_X1 U504 ( .A1(data_in[0]), .A2(n827), .B1(n965), .B2(\mem[26][0] ), 
        .ZN(n966) );
  INV_X1 U505 ( .A(n964), .ZN(n676) );
  AOI22_X1 U506 ( .A1(data_in[1]), .A2(n827), .B1(n965), .B2(\mem[26][1] ), 
        .ZN(n964) );
  INV_X1 U507 ( .A(n963), .ZN(n675) );
  AOI22_X1 U508 ( .A1(data_in[2]), .A2(n827), .B1(n965), .B2(\mem[26][2] ), 
        .ZN(n963) );
  INV_X1 U509 ( .A(n962), .ZN(n674) );
  AOI22_X1 U510 ( .A1(data_in[3]), .A2(n827), .B1(n965), .B2(\mem[26][3] ), 
        .ZN(n962) );
  INV_X1 U511 ( .A(n961), .ZN(n673) );
  AOI22_X1 U512 ( .A1(data_in[4]), .A2(n827), .B1(n965), .B2(\mem[26][4] ), 
        .ZN(n961) );
  INV_X1 U513 ( .A(n960), .ZN(n672) );
  AOI22_X1 U514 ( .A1(data_in[5]), .A2(n827), .B1(n965), .B2(\mem[26][5] ), 
        .ZN(n960) );
  INV_X1 U515 ( .A(n959), .ZN(n671) );
  AOI22_X1 U516 ( .A1(data_in[6]), .A2(n827), .B1(n965), .B2(\mem[26][6] ), 
        .ZN(n959) );
  INV_X1 U517 ( .A(n958), .ZN(n670) );
  AOI22_X1 U518 ( .A1(data_in[7]), .A2(n827), .B1(n965), .B2(\mem[26][7] ), 
        .ZN(n958) );
  INV_X1 U519 ( .A(n957), .ZN(n669) );
  AOI22_X1 U520 ( .A1(data_in[0]), .A2(n826), .B1(n956), .B2(\mem[27][0] ), 
        .ZN(n957) );
  INV_X1 U521 ( .A(n955), .ZN(n668) );
  AOI22_X1 U522 ( .A1(data_in[1]), .A2(n826), .B1(n956), .B2(\mem[27][1] ), 
        .ZN(n955) );
  INV_X1 U523 ( .A(n954), .ZN(n667) );
  AOI22_X1 U524 ( .A1(data_in[2]), .A2(n826), .B1(n956), .B2(\mem[27][2] ), 
        .ZN(n954) );
  INV_X1 U525 ( .A(n953), .ZN(n666) );
  AOI22_X1 U526 ( .A1(data_in[3]), .A2(n826), .B1(n956), .B2(\mem[27][3] ), 
        .ZN(n953) );
  INV_X1 U527 ( .A(n952), .ZN(n665) );
  AOI22_X1 U528 ( .A1(data_in[4]), .A2(n826), .B1(n956), .B2(\mem[27][4] ), 
        .ZN(n952) );
  INV_X1 U529 ( .A(n951), .ZN(n664) );
  AOI22_X1 U530 ( .A1(data_in[5]), .A2(n826), .B1(n956), .B2(\mem[27][5] ), 
        .ZN(n951) );
  INV_X1 U531 ( .A(n950), .ZN(n663) );
  AOI22_X1 U532 ( .A1(data_in[6]), .A2(n826), .B1(n956), .B2(\mem[27][6] ), 
        .ZN(n950) );
  INV_X1 U533 ( .A(n949), .ZN(n662) );
  AOI22_X1 U534 ( .A1(data_in[7]), .A2(n826), .B1(n956), .B2(\mem[27][7] ), 
        .ZN(n949) );
  INV_X1 U535 ( .A(n948), .ZN(n661) );
  AOI22_X1 U536 ( .A1(data_in[0]), .A2(n825), .B1(n947), .B2(\mem[28][0] ), 
        .ZN(n948) );
  INV_X1 U537 ( .A(n946), .ZN(n660) );
  AOI22_X1 U538 ( .A1(data_in[1]), .A2(n825), .B1(n947), .B2(\mem[28][1] ), 
        .ZN(n946) );
  INV_X1 U539 ( .A(n945), .ZN(n659) );
  AOI22_X1 U540 ( .A1(data_in[2]), .A2(n825), .B1(n947), .B2(\mem[28][2] ), 
        .ZN(n945) );
  INV_X1 U541 ( .A(n944), .ZN(n658) );
  AOI22_X1 U542 ( .A1(data_in[3]), .A2(n825), .B1(n947), .B2(\mem[28][3] ), 
        .ZN(n944) );
  INV_X1 U543 ( .A(n943), .ZN(n657) );
  AOI22_X1 U544 ( .A1(data_in[4]), .A2(n825), .B1(n947), .B2(\mem[28][4] ), 
        .ZN(n943) );
  INV_X1 U545 ( .A(n942), .ZN(n656) );
  AOI22_X1 U546 ( .A1(data_in[5]), .A2(n825), .B1(n947), .B2(\mem[28][5] ), 
        .ZN(n942) );
  INV_X1 U547 ( .A(n941), .ZN(n655) );
  AOI22_X1 U548 ( .A1(data_in[6]), .A2(n825), .B1(n947), .B2(\mem[28][6] ), 
        .ZN(n941) );
  INV_X1 U549 ( .A(n940), .ZN(n654) );
  AOI22_X1 U550 ( .A1(data_in[7]), .A2(n825), .B1(n947), .B2(\mem[28][7] ), 
        .ZN(n940) );
  INV_X1 U551 ( .A(n939), .ZN(n653) );
  AOI22_X1 U552 ( .A1(data_in[0]), .A2(n824), .B1(n938), .B2(\mem[29][0] ), 
        .ZN(n939) );
  INV_X1 U553 ( .A(n937), .ZN(n652) );
  AOI22_X1 U554 ( .A1(data_in[1]), .A2(n824), .B1(n938), .B2(\mem[29][1] ), 
        .ZN(n937) );
  INV_X1 U555 ( .A(n936), .ZN(n651) );
  AOI22_X1 U556 ( .A1(data_in[2]), .A2(n824), .B1(n938), .B2(\mem[29][2] ), 
        .ZN(n936) );
  INV_X1 U557 ( .A(n935), .ZN(n650) );
  AOI22_X1 U558 ( .A1(data_in[3]), .A2(n824), .B1(n938), .B2(\mem[29][3] ), 
        .ZN(n935) );
  INV_X1 U559 ( .A(n934), .ZN(n649) );
  AOI22_X1 U560 ( .A1(data_in[4]), .A2(n824), .B1(n938), .B2(\mem[29][4] ), 
        .ZN(n934) );
  INV_X1 U561 ( .A(n933), .ZN(n648) );
  AOI22_X1 U562 ( .A1(data_in[5]), .A2(n824), .B1(n938), .B2(\mem[29][5] ), 
        .ZN(n933) );
  INV_X1 U563 ( .A(n932), .ZN(n647) );
  AOI22_X1 U564 ( .A1(data_in[6]), .A2(n824), .B1(n938), .B2(\mem[29][6] ), 
        .ZN(n932) );
  INV_X1 U565 ( .A(n931), .ZN(n646) );
  AOI22_X1 U566 ( .A1(data_in[7]), .A2(n824), .B1(n938), .B2(\mem[29][7] ), 
        .ZN(n931) );
  INV_X1 U567 ( .A(n930), .ZN(n645) );
  AOI22_X1 U568 ( .A1(data_in[0]), .A2(n823), .B1(n929), .B2(\mem[30][0] ), 
        .ZN(n930) );
  INV_X1 U569 ( .A(n928), .ZN(n644) );
  AOI22_X1 U570 ( .A1(data_in[1]), .A2(n823), .B1(n929), .B2(\mem[30][1] ), 
        .ZN(n928) );
  INV_X1 U571 ( .A(n927), .ZN(n643) );
  AOI22_X1 U572 ( .A1(data_in[2]), .A2(n823), .B1(n929), .B2(\mem[30][2] ), 
        .ZN(n927) );
  INV_X1 U573 ( .A(n926), .ZN(n642) );
  AOI22_X1 U574 ( .A1(data_in[3]), .A2(n823), .B1(n929), .B2(\mem[30][3] ), 
        .ZN(n926) );
  INV_X1 U575 ( .A(n925), .ZN(n641) );
  AOI22_X1 U576 ( .A1(data_in[4]), .A2(n823), .B1(n929), .B2(\mem[30][4] ), 
        .ZN(n925) );
  INV_X1 U577 ( .A(n924), .ZN(n640) );
  AOI22_X1 U578 ( .A1(data_in[5]), .A2(n823), .B1(n929), .B2(\mem[30][5] ), 
        .ZN(n924) );
  INV_X1 U579 ( .A(n923), .ZN(n639) );
  AOI22_X1 U580 ( .A1(data_in[6]), .A2(n823), .B1(n929), .B2(\mem[30][6] ), 
        .ZN(n923) );
  INV_X1 U581 ( .A(n922), .ZN(n638) );
  AOI22_X1 U582 ( .A1(data_in[7]), .A2(n823), .B1(n929), .B2(\mem[30][7] ), 
        .ZN(n922) );
  INV_X1 U583 ( .A(n921), .ZN(n637) );
  AOI22_X1 U584 ( .A1(data_in[0]), .A2(n822), .B1(n920), .B2(\mem[31][0] ), 
        .ZN(n921) );
  INV_X1 U585 ( .A(n919), .ZN(n636) );
  AOI22_X1 U586 ( .A1(data_in[1]), .A2(n822), .B1(n920), .B2(\mem[31][1] ), 
        .ZN(n919) );
  INV_X1 U587 ( .A(n918), .ZN(n635) );
  AOI22_X1 U588 ( .A1(data_in[2]), .A2(n822), .B1(n920), .B2(\mem[31][2] ), 
        .ZN(n918) );
  INV_X1 U589 ( .A(n917), .ZN(n634) );
  AOI22_X1 U590 ( .A1(data_in[3]), .A2(n822), .B1(n920), .B2(\mem[31][3] ), 
        .ZN(n917) );
  INV_X1 U591 ( .A(n916), .ZN(n633) );
  AOI22_X1 U592 ( .A1(data_in[4]), .A2(n822), .B1(n920), .B2(\mem[31][4] ), 
        .ZN(n916) );
  INV_X1 U593 ( .A(n915), .ZN(n632) );
  AOI22_X1 U594 ( .A1(data_in[5]), .A2(n822), .B1(n920), .B2(\mem[31][5] ), 
        .ZN(n915) );
  INV_X1 U595 ( .A(n914), .ZN(n631) );
  AOI22_X1 U596 ( .A1(data_in[6]), .A2(n822), .B1(n920), .B2(\mem[31][6] ), 
        .ZN(n914) );
  INV_X1 U597 ( .A(n913), .ZN(n630) );
  AOI22_X1 U598 ( .A1(data_in[7]), .A2(n822), .B1(n920), .B2(\mem[31][7] ), 
        .ZN(n913) );
  MUX2_X1 U599 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n613), .Z(n3) );
  MUX2_X1 U600 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n613), .Z(n4) );
  MUX2_X1 U601 ( .A(n4), .B(n3), .S(n610), .Z(n5) );
  MUX2_X1 U602 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n613), .Z(n6) );
  MUX2_X1 U603 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n613), .Z(n7) );
  MUX2_X1 U604 ( .A(n7), .B(n6), .S(n610), .Z(n8) );
  MUX2_X1 U605 ( .A(n8), .B(n5), .S(N12), .Z(n9) );
  MUX2_X1 U606 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n613), .Z(n10) );
  MUX2_X1 U607 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n613), .Z(n11) );
  MUX2_X1 U608 ( .A(n11), .B(n10), .S(n610), .Z(n12) );
  MUX2_X1 U609 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n613), .Z(n13) );
  MUX2_X1 U610 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n613), .Z(n14) );
  MUX2_X1 U611 ( .A(n14), .B(n13), .S(n610), .Z(n15) );
  MUX2_X1 U612 ( .A(n15), .B(n12), .S(n608), .Z(n16) );
  MUX2_X1 U613 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U614 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n614), .Z(n18) );
  MUX2_X1 U615 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n614), .Z(n19) );
  MUX2_X1 U616 ( .A(n19), .B(n18), .S(n610), .Z(n20) );
  MUX2_X1 U617 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n614), .Z(n21) );
  MUX2_X1 U618 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n614), .Z(n22) );
  MUX2_X1 U619 ( .A(n22), .B(n21), .S(N11), .Z(n23) );
  MUX2_X1 U620 ( .A(n23), .B(n20), .S(n609), .Z(n24) );
  MUX2_X1 U621 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n614), .Z(n25) );
  MUX2_X1 U622 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n614), .Z(n26) );
  MUX2_X1 U623 ( .A(n26), .B(n25), .S(N11), .Z(n27) );
  MUX2_X1 U624 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n614), .Z(n28) );
  MUX2_X1 U625 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n614), .Z(n29) );
  MUX2_X1 U626 ( .A(n29), .B(n28), .S(n612), .Z(n30) );
  MUX2_X1 U627 ( .A(n30), .B(n27), .S(n609), .Z(n31) );
  MUX2_X1 U628 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U629 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U630 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n614), .Z(n33) );
  MUX2_X1 U631 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n614), .Z(n34) );
  MUX2_X1 U632 ( .A(n34), .B(n33), .S(n611), .Z(n35) );
  MUX2_X1 U633 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n614), .Z(n36) );
  MUX2_X1 U634 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n614), .Z(n37) );
  MUX2_X1 U635 ( .A(n37), .B(n36), .S(N11), .Z(n38) );
  MUX2_X1 U636 ( .A(n38), .B(n35), .S(N12), .Z(n39) );
  MUX2_X1 U637 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n615), .Z(n40) );
  MUX2_X1 U638 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n615), .Z(n41) );
  MUX2_X1 U639 ( .A(n41), .B(n40), .S(n611), .Z(n42) );
  MUX2_X1 U640 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n615), .Z(n43) );
  MUX2_X1 U641 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n615), .Z(n44) );
  MUX2_X1 U642 ( .A(n44), .B(n43), .S(n612), .Z(n45) );
  MUX2_X1 U643 ( .A(n45), .B(n42), .S(n609), .Z(n46) );
  MUX2_X1 U644 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U645 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n615), .Z(n48) );
  MUX2_X1 U646 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n615), .Z(n49) );
  MUX2_X1 U647 ( .A(n49), .B(n48), .S(n612), .Z(n50) );
  MUX2_X1 U648 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n615), .Z(n51) );
  MUX2_X1 U649 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n615), .Z(n52) );
  MUX2_X1 U650 ( .A(n52), .B(n51), .S(n610), .Z(n53) );
  MUX2_X1 U651 ( .A(n53), .B(n50), .S(n608), .Z(n54) );
  MUX2_X1 U652 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n615), .Z(n55) );
  MUX2_X1 U653 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n615), .Z(n56) );
  MUX2_X1 U654 ( .A(n56), .B(n55), .S(N11), .Z(n57) );
  MUX2_X1 U655 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n615), .Z(n58) );
  MUX2_X1 U656 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n615), .Z(n59) );
  MUX2_X1 U657 ( .A(n59), .B(n58), .S(n611), .Z(n60) );
  MUX2_X1 U658 ( .A(n60), .B(n57), .S(N12), .Z(n61) );
  MUX2_X1 U659 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U660 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U661 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n616), .Z(n63) );
  MUX2_X1 U662 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n616), .Z(n64) );
  MUX2_X1 U663 ( .A(n64), .B(n63), .S(n610), .Z(n65) );
  MUX2_X1 U664 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n616), .Z(n66) );
  MUX2_X1 U665 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n616), .Z(n67) );
  MUX2_X1 U666 ( .A(n67), .B(n66), .S(n610), .Z(n68) );
  MUX2_X1 U667 ( .A(n68), .B(n65), .S(n608), .Z(n69) );
  MUX2_X1 U668 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n616), .Z(n70) );
  MUX2_X1 U669 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n616), .Z(n71) );
  MUX2_X1 U670 ( .A(n71), .B(n70), .S(n610), .Z(n72) );
  MUX2_X1 U671 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n616), .Z(n73) );
  MUX2_X1 U672 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n616), .Z(n74) );
  MUX2_X1 U673 ( .A(n74), .B(n73), .S(n610), .Z(n75) );
  MUX2_X1 U674 ( .A(n75), .B(n72), .S(n608), .Z(n76) );
  MUX2_X1 U675 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U676 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n616), .Z(n78) );
  MUX2_X1 U677 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n616), .Z(n79) );
  MUX2_X1 U678 ( .A(n79), .B(n78), .S(n610), .Z(n80) );
  MUX2_X1 U679 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n616), .Z(n81) );
  MUX2_X1 U680 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n616), .Z(n82) );
  MUX2_X1 U681 ( .A(n82), .B(n81), .S(n612), .Z(n83) );
  MUX2_X1 U682 ( .A(n83), .B(n80), .S(n608), .Z(n84) );
  MUX2_X1 U683 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n619), .Z(n85) );
  MUX2_X1 U684 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n613), .Z(n86) );
  MUX2_X1 U685 ( .A(n86), .B(n85), .S(n611), .Z(n87) );
  MUX2_X1 U686 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n618), .Z(n88) );
  MUX2_X1 U687 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n617), .Z(n89) );
  MUX2_X1 U688 ( .A(n89), .B(n88), .S(n610), .Z(n90) );
  MUX2_X1 U689 ( .A(n90), .B(n87), .S(n608), .Z(n91) );
  MUX2_X1 U690 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U691 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U692 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n618), .Z(n93) );
  MUX2_X1 U693 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n618), .Z(n94) );
  MUX2_X1 U694 ( .A(n94), .B(n93), .S(n610), .Z(n95) );
  MUX2_X1 U695 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n617), .Z(n96) );
  MUX2_X1 U696 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n617), .Z(n97) );
  MUX2_X1 U697 ( .A(n97), .B(n96), .S(n610), .Z(n98) );
  MUX2_X1 U698 ( .A(n98), .B(n95), .S(n608), .Z(n99) );
  MUX2_X1 U699 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n617), .Z(n100) );
  MUX2_X1 U700 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n617), .Z(n101) );
  MUX2_X1 U701 ( .A(n101), .B(n100), .S(n610), .Z(n102) );
  MUX2_X1 U702 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n616), .Z(n103) );
  MUX2_X1 U703 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n615), .Z(n104) );
  MUX2_X1 U704 ( .A(n104), .B(n103), .S(n612), .Z(n105) );
  MUX2_X1 U705 ( .A(n105), .B(n102), .S(n608), .Z(n106) );
  MUX2_X1 U706 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U707 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n613), .Z(n108) );
  MUX2_X1 U708 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n615), .Z(n109) );
  MUX2_X1 U709 ( .A(n109), .B(n108), .S(n611), .Z(n110) );
  MUX2_X1 U710 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n614), .Z(n111) );
  MUX2_X1 U711 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n112) );
  MUX2_X1 U712 ( .A(n112), .B(n111), .S(n611), .Z(n113) );
  MUX2_X1 U713 ( .A(n113), .B(n110), .S(n608), .Z(n114) );
  MUX2_X1 U714 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n619), .Z(n115) );
  MUX2_X1 U715 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n116) );
  MUX2_X1 U716 ( .A(n116), .B(n115), .S(n611), .Z(n117) );
  MUX2_X1 U717 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n118) );
  MUX2_X1 U718 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n119) );
  MUX2_X1 U719 ( .A(n119), .B(n118), .S(n611), .Z(n120) );
  MUX2_X1 U720 ( .A(n120), .B(n117), .S(n608), .Z(n121) );
  MUX2_X1 U721 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U722 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U723 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n613), .Z(n123) );
  MUX2_X1 U724 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n613), .Z(n124) );
  MUX2_X1 U725 ( .A(n124), .B(n123), .S(n611), .Z(n125) );
  MUX2_X1 U726 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n613), .Z(n126) );
  MUX2_X1 U727 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n619), .Z(n127) );
  MUX2_X1 U728 ( .A(n127), .B(n126), .S(n611), .Z(n128) );
  MUX2_X1 U729 ( .A(n128), .B(n125), .S(n608), .Z(n129) );
  MUX2_X1 U730 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n617), .Z(n130) );
  MUX2_X1 U731 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n617), .Z(n131) );
  MUX2_X1 U732 ( .A(n131), .B(n130), .S(n611), .Z(n132) );
  MUX2_X1 U733 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n617), .Z(n133) );
  MUX2_X1 U734 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n617), .Z(n134) );
  MUX2_X1 U735 ( .A(n134), .B(n133), .S(n611), .Z(n135) );
  MUX2_X1 U736 ( .A(n135), .B(n132), .S(n608), .Z(n136) );
  MUX2_X1 U737 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U738 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n617), .Z(n138) );
  MUX2_X1 U739 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n617), .Z(n139) );
  MUX2_X1 U740 ( .A(n139), .B(n138), .S(n611), .Z(n140) );
  MUX2_X1 U741 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n617), .Z(n141) );
  MUX2_X1 U742 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n617), .Z(n142) );
  MUX2_X1 U743 ( .A(n142), .B(n141), .S(n611), .Z(n143) );
  MUX2_X1 U744 ( .A(n143), .B(n140), .S(n608), .Z(n144) );
  MUX2_X1 U745 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n617), .Z(n145) );
  MUX2_X1 U746 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n617), .Z(n146) );
  MUX2_X1 U747 ( .A(n146), .B(n145), .S(n611), .Z(n147) );
  MUX2_X1 U748 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n617), .Z(n148) );
  MUX2_X1 U749 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n617), .Z(n149) );
  MUX2_X1 U750 ( .A(n149), .B(n148), .S(n611), .Z(n150) );
  MUX2_X1 U751 ( .A(n150), .B(n147), .S(n608), .Z(n151) );
  MUX2_X1 U752 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U753 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U754 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n618), .Z(n153) );
  MUX2_X1 U755 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n618), .Z(n154) );
  MUX2_X1 U756 ( .A(n154), .B(n153), .S(n612), .Z(n155) );
  MUX2_X1 U757 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n618), .Z(n156) );
  MUX2_X1 U758 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n618), .Z(n157) );
  MUX2_X1 U759 ( .A(n157), .B(n156), .S(n612), .Z(n158) );
  MUX2_X1 U760 ( .A(n158), .B(n155), .S(n609), .Z(n159) );
  MUX2_X1 U761 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n618), .Z(n160) );
  MUX2_X1 U762 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n618), .Z(n161) );
  MUX2_X1 U763 ( .A(n161), .B(n160), .S(n612), .Z(n162) );
  MUX2_X1 U764 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n618), .Z(n163) );
  MUX2_X1 U765 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n618), .Z(n164) );
  MUX2_X1 U766 ( .A(n164), .B(n163), .S(n612), .Z(n165) );
  MUX2_X1 U767 ( .A(n165), .B(n162), .S(n609), .Z(n166) );
  MUX2_X1 U768 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U769 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n618), .Z(n168) );
  MUX2_X1 U770 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n618), .Z(n169) );
  MUX2_X1 U771 ( .A(n169), .B(n168), .S(n612), .Z(n170) );
  MUX2_X1 U772 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n618), .Z(n171) );
  MUX2_X1 U773 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n618), .Z(n172) );
  MUX2_X1 U774 ( .A(n172), .B(n171), .S(n612), .Z(n173) );
  MUX2_X1 U775 ( .A(n173), .B(n170), .S(n609), .Z(n174) );
  MUX2_X1 U776 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n613), .Z(n175) );
  MUX2_X1 U777 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n619), .Z(n176) );
  MUX2_X1 U778 ( .A(n176), .B(n175), .S(n612), .Z(n177) );
  MUX2_X1 U779 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n619), .Z(n178) );
  MUX2_X1 U780 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n615), .Z(n179) );
  MUX2_X1 U781 ( .A(n179), .B(n178), .S(n612), .Z(n180) );
  MUX2_X1 U782 ( .A(n180), .B(n177), .S(n609), .Z(n181) );
  MUX2_X1 U783 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U784 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U785 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n619), .Z(n183) );
  MUX2_X1 U786 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n614), .Z(n184) );
  MUX2_X1 U787 ( .A(n184), .B(n183), .S(n612), .Z(n185) );
  MUX2_X1 U788 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n619), .Z(n186) );
  MUX2_X1 U789 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n619), .Z(n187) );
  MUX2_X1 U790 ( .A(n187), .B(n186), .S(n612), .Z(n188) );
  MUX2_X1 U791 ( .A(n188), .B(n185), .S(n609), .Z(n189) );
  MUX2_X1 U792 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n619), .Z(n190) );
  MUX2_X1 U793 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n616), .Z(n191) );
  MUX2_X1 U794 ( .A(n191), .B(n190), .S(n612), .Z(n192) );
  MUX2_X1 U795 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n615), .Z(n193) );
  MUX2_X1 U796 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n613), .Z(n194) );
  MUX2_X1 U797 ( .A(n194), .B(n193), .S(n612), .Z(n195) );
  MUX2_X1 U798 ( .A(n195), .B(n192), .S(n609), .Z(n196) );
  MUX2_X1 U799 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U800 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n619), .Z(n198) );
  MUX2_X1 U801 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n619), .Z(n199) );
  MUX2_X1 U802 ( .A(n199), .B(n198), .S(n611), .Z(n200) );
  MUX2_X1 U803 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n619), .Z(n201) );
  MUX2_X1 U804 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n616), .Z(n202) );
  MUX2_X1 U805 ( .A(n202), .B(n201), .S(n612), .Z(n203) );
  MUX2_X1 U806 ( .A(n203), .B(n200), .S(n609), .Z(n204) );
  MUX2_X1 U807 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n619), .Z(n205) );
  MUX2_X1 U808 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n619), .Z(n206) );
  MUX2_X1 U809 ( .A(n206), .B(n205), .S(n611), .Z(n207) );
  MUX2_X1 U810 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n619), .Z(n208) );
  MUX2_X1 U811 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n613), .Z(n209) );
  MUX2_X1 U812 ( .A(n209), .B(n208), .S(n610), .Z(n210) );
  MUX2_X1 U813 ( .A(n210), .B(n207), .S(n609), .Z(n211) );
  MUX2_X1 U814 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U815 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U816 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n619), .Z(n213) );
  MUX2_X1 U817 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n619), .Z(n214) );
  MUX2_X1 U818 ( .A(n214), .B(n213), .S(n612), .Z(n215) );
  MUX2_X1 U819 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n616), .Z(n216) );
  MUX2_X1 U820 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n618), .Z(n217) );
  MUX2_X1 U821 ( .A(n217), .B(n216), .S(n612), .Z(n218) );
  MUX2_X1 U822 ( .A(n218), .B(n215), .S(n609), .Z(n219) );
  MUX2_X1 U823 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n614), .Z(n220) );
  MUX2_X1 U824 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n615), .Z(n221) );
  MUX2_X1 U825 ( .A(n221), .B(n220), .S(N11), .Z(n222) );
  MUX2_X1 U826 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n619), .Z(n223) );
  MUX2_X1 U827 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n614), .Z(n224) );
  MUX2_X1 U828 ( .A(n224), .B(n223), .S(n611), .Z(n225) );
  MUX2_X1 U829 ( .A(n225), .B(n222), .S(n609), .Z(n226) );
  MUX2_X1 U830 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U831 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n613), .Z(n228) );
  MUX2_X1 U832 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n618), .Z(n229) );
  MUX2_X1 U833 ( .A(n229), .B(n228), .S(n610), .Z(n595) );
  MUX2_X1 U834 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n613), .Z(n596) );
  MUX2_X1 U835 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n619), .Z(n597) );
  MUX2_X1 U836 ( .A(n597), .B(n596), .S(n611), .Z(n598) );
  MUX2_X1 U837 ( .A(n598), .B(n595), .S(n609), .Z(n599) );
  MUX2_X1 U838 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n616), .Z(n600) );
  MUX2_X1 U839 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n601) );
  MUX2_X1 U840 ( .A(n601), .B(n600), .S(n610), .Z(n602) );
  MUX2_X1 U841 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n614), .Z(n603) );
  MUX2_X1 U842 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n604) );
  MUX2_X1 U843 ( .A(n604), .B(n603), .S(n612), .Z(n605) );
  MUX2_X1 U844 ( .A(n605), .B(n602), .S(n609), .Z(n606) );
  MUX2_X1 U845 ( .A(n606), .B(n599), .S(N13), .Z(n607) );
  MUX2_X1 U846 ( .A(n607), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U847 ( .A(N11), .Z(n610) );
  INV_X1 U848 ( .A(N10), .ZN(n620) );
  INV_X1 U849 ( .A(N11), .ZN(n621) );
  INV_X1 U850 ( .A(data_in[0]), .ZN(n622) );
  INV_X1 U851 ( .A(data_in[1]), .ZN(n623) );
  INV_X1 U852 ( .A(data_in[2]), .ZN(n624) );
  INV_X1 U853 ( .A(data_in[3]), .ZN(n625) );
  INV_X1 U854 ( .A(data_in[4]), .ZN(n626) );
  INV_X1 U855 ( .A(data_in[5]), .ZN(n627) );
  INV_X1 U856 ( .A(data_in[6]), .ZN(n628) );
  INV_X1 U857 ( .A(data_in[7]), .ZN(n629) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_18 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n627), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n628), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n629), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n630), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n631), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n632), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n633), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n634), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n635), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n636), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n637), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n638), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n639), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n640), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n641), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n642), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n643), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n644), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n645), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n646), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n647), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n648), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n649), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n650), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n651), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n652), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n653), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n654), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n655), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n656), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n657), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n658), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n659), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n660), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n661), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n662), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n663), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n664), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n665), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n666), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n667), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n668), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n669), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n670), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n671), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n672), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n673), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n674), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n675), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n676), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n677), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n678), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n679), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n680), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n681), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n682), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n683), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n684), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n685), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n686), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n687), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n688), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n689), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n690), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n691), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n692), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n693), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n694), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n695), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n696), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n697), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n698), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n699), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n700), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n701), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n702), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n703), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n704), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n705), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n706), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n707), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n708), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n709), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n710), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n711), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n712), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n713), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n714), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n715), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n716), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n717), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n718), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n719), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n720), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n721), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n722), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n723), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n724), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n725), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n726), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n727), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n728), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n729), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n730), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n731), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n732), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n733), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n734), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n735), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n736), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n737), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n738), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n739), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n740), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n741), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n742), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n743), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n744), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n745), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n746), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n747), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n748), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n749), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n750), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n751), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n752), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n753), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n754), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n755), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n756), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n757), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n758), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n759), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n760), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n761), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n762), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n763), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n764), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n765), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n766), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n767), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n768), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n769), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n770), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n771), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n772), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n773), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n774), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n775), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n776), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n777), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n778), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n779), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n780), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n781), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n782), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n783), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n784), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n785), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n786), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n787), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n788), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n789), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n790), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n791), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n792), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n793), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n794), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n795), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n796), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n797), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n798), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n799), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n800), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n801), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n802), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n803), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n804), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n805), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n806), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n807), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n808), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n809), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n810), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n811), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n812), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n813), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n814), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n815), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n816), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n817), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n818), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n846), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n847), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n848), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n849), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n850), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n851), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n852), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n853), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n854), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n855), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n856), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n857), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n858), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n859), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n860), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n861), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n862), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n863), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n864), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n865), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n866), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n867), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n868), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n869), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n870), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n871), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n872), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n873), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n874), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n875), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n876), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n877), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n878), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n879), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n880), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n881), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n882), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n883), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n884), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n885), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n886), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n887), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n888), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n889), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n890), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n891), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n892), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n893), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n894), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n895), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n896), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n897), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n898), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n899), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n900), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n901), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n902), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n903), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n904), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n905), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n906), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n907), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n908), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n909), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  BUF_X1 U3 ( .A(n616), .Z(n611) );
  BUF_X1 U4 ( .A(n616), .Z(n614) );
  BUF_X1 U5 ( .A(n616), .Z(n615) );
  BUF_X1 U6 ( .A(n616), .Z(n612) );
  BUF_X1 U7 ( .A(N10), .Z(n613) );
  BUF_X1 U8 ( .A(N11), .Z(n609) );
  BUF_X1 U9 ( .A(N11), .Z(n610) );
  BUF_X1 U10 ( .A(N10), .Z(n616) );
  NOR3_X1 U11 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1201) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(n617), .ZN(n1190) );
  NOR3_X1 U13 ( .A1(N10), .A2(N12), .A3(n618), .ZN(n1180) );
  NOR3_X1 U14 ( .A1(n617), .A2(N12), .A3(n618), .ZN(n1170) );
  INV_X1 U15 ( .A(n1127), .ZN(n842) );
  INV_X1 U16 ( .A(n1117), .ZN(n841) );
  INV_X1 U17 ( .A(n1108), .ZN(n840) );
  INV_X1 U18 ( .A(n1099), .ZN(n839) );
  INV_X1 U19 ( .A(n1054), .ZN(n834) );
  INV_X1 U20 ( .A(n1044), .ZN(n833) );
  INV_X1 U21 ( .A(n1035), .ZN(n832) );
  INV_X1 U22 ( .A(n1026), .ZN(n831) );
  INV_X1 U23 ( .A(n981), .ZN(n826) );
  INV_X1 U24 ( .A(n971), .ZN(n825) );
  INV_X1 U25 ( .A(n962), .ZN(n824) );
  INV_X1 U26 ( .A(n953), .ZN(n823) );
  INV_X1 U27 ( .A(n1090), .ZN(n838) );
  INV_X1 U28 ( .A(n1081), .ZN(n837) );
  INV_X1 U29 ( .A(n1072), .ZN(n836) );
  INV_X1 U30 ( .A(n1063), .ZN(n835) );
  INV_X1 U31 ( .A(n944), .ZN(n822) );
  INV_X1 U32 ( .A(n935), .ZN(n821) );
  INV_X1 U33 ( .A(n926), .ZN(n820) );
  INV_X1 U34 ( .A(n917), .ZN(n819) );
  INV_X1 U35 ( .A(n1017), .ZN(n830) );
  INV_X1 U36 ( .A(n1008), .ZN(n829) );
  INV_X1 U37 ( .A(n999), .ZN(n828) );
  INV_X1 U38 ( .A(n990), .ZN(n827) );
  BUF_X1 U39 ( .A(N12), .Z(n606) );
  BUF_X1 U40 ( .A(N12), .Z(n607) );
  INV_X1 U41 ( .A(N13), .ZN(n844) );
  AND3_X1 U42 ( .A1(n617), .A2(n618), .A3(N12), .ZN(n1160) );
  AND3_X1 U43 ( .A1(N10), .A2(n618), .A3(N12), .ZN(n1150) );
  AND3_X1 U44 ( .A1(N11), .A2(n617), .A3(N12), .ZN(n1140) );
  AND3_X1 U45 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1130) );
  INV_X1 U46 ( .A(N14), .ZN(n845) );
  NAND2_X1 U47 ( .A1(n1190), .A2(n1200), .ZN(n1199) );
  NAND2_X1 U48 ( .A1(n1180), .A2(n1200), .ZN(n1189) );
  NAND2_X1 U49 ( .A1(n1170), .A2(n1200), .ZN(n1179) );
  NAND2_X1 U50 ( .A1(n1160), .A2(n1200), .ZN(n1169) );
  NAND2_X1 U51 ( .A1(n1150), .A2(n1200), .ZN(n1159) );
  NAND2_X1 U52 ( .A1(n1140), .A2(n1200), .ZN(n1149) );
  NAND2_X1 U53 ( .A1(n1130), .A2(n1200), .ZN(n1139) );
  NAND2_X1 U54 ( .A1(n1201), .A2(n1200), .ZN(n1210) );
  NAND2_X1 U55 ( .A1(n1119), .A2(n1201), .ZN(n1127) );
  NAND2_X1 U56 ( .A1(n1119), .A2(n1190), .ZN(n1117) );
  NAND2_X1 U57 ( .A1(n1119), .A2(n1180), .ZN(n1108) );
  NAND2_X1 U58 ( .A1(n1119), .A2(n1170), .ZN(n1099) );
  NAND2_X1 U59 ( .A1(n1046), .A2(n1201), .ZN(n1054) );
  NAND2_X1 U60 ( .A1(n1046), .A2(n1190), .ZN(n1044) );
  NAND2_X1 U61 ( .A1(n1046), .A2(n1180), .ZN(n1035) );
  NAND2_X1 U62 ( .A1(n1046), .A2(n1170), .ZN(n1026) );
  NAND2_X1 U63 ( .A1(n973), .A2(n1201), .ZN(n981) );
  NAND2_X1 U64 ( .A1(n973), .A2(n1190), .ZN(n971) );
  NAND2_X1 U65 ( .A1(n973), .A2(n1180), .ZN(n962) );
  NAND2_X1 U66 ( .A1(n973), .A2(n1170), .ZN(n953) );
  NAND2_X1 U67 ( .A1(n1119), .A2(n1160), .ZN(n1090) );
  NAND2_X1 U68 ( .A1(n1119), .A2(n1150), .ZN(n1081) );
  NAND2_X1 U69 ( .A1(n1119), .A2(n1140), .ZN(n1072) );
  NAND2_X1 U70 ( .A1(n1119), .A2(n1130), .ZN(n1063) );
  NAND2_X1 U71 ( .A1(n1046), .A2(n1160), .ZN(n1017) );
  NAND2_X1 U72 ( .A1(n1046), .A2(n1150), .ZN(n1008) );
  NAND2_X1 U73 ( .A1(n1046), .A2(n1140), .ZN(n999) );
  NAND2_X1 U74 ( .A1(n1046), .A2(n1130), .ZN(n990) );
  NAND2_X1 U75 ( .A1(n973), .A2(n1160), .ZN(n944) );
  NAND2_X1 U76 ( .A1(n973), .A2(n1150), .ZN(n935) );
  NAND2_X1 U77 ( .A1(n973), .A2(n1140), .ZN(n926) );
  NAND2_X1 U78 ( .A1(n973), .A2(n1130), .ZN(n917) );
  AND3_X1 U79 ( .A1(n844), .A2(n845), .A3(n1129), .ZN(n1200) );
  AND3_X1 U80 ( .A1(N13), .A2(n1129), .A3(N14), .ZN(n973) );
  AND3_X1 U81 ( .A1(n1129), .A2(n845), .A3(N13), .ZN(n1119) );
  AND3_X1 U82 ( .A1(n1129), .A2(n844), .A3(N14), .ZN(n1046) );
  NOR2_X1 U83 ( .A1(n843), .A2(addr[5]), .ZN(n1129) );
  INV_X1 U84 ( .A(wr_en), .ZN(n843) );
  OAI21_X1 U85 ( .B1(n619), .B2(n1169), .A(n1168), .ZN(n877) );
  NAND2_X1 U86 ( .A1(\mem[4][0] ), .A2(n1169), .ZN(n1168) );
  OAI21_X1 U87 ( .B1(n620), .B2(n1169), .A(n1167), .ZN(n876) );
  NAND2_X1 U88 ( .A1(\mem[4][1] ), .A2(n1169), .ZN(n1167) );
  OAI21_X1 U89 ( .B1(n621), .B2(n1169), .A(n1166), .ZN(n875) );
  NAND2_X1 U90 ( .A1(\mem[4][2] ), .A2(n1169), .ZN(n1166) );
  OAI21_X1 U91 ( .B1(n622), .B2(n1169), .A(n1165), .ZN(n874) );
  NAND2_X1 U92 ( .A1(\mem[4][3] ), .A2(n1169), .ZN(n1165) );
  OAI21_X1 U93 ( .B1(n623), .B2(n1169), .A(n1164), .ZN(n873) );
  NAND2_X1 U94 ( .A1(\mem[4][4] ), .A2(n1169), .ZN(n1164) );
  OAI21_X1 U95 ( .B1(n624), .B2(n1169), .A(n1163), .ZN(n872) );
  NAND2_X1 U96 ( .A1(\mem[4][5] ), .A2(n1169), .ZN(n1163) );
  OAI21_X1 U97 ( .B1(n625), .B2(n1169), .A(n1162), .ZN(n871) );
  NAND2_X1 U98 ( .A1(\mem[4][6] ), .A2(n1169), .ZN(n1162) );
  OAI21_X1 U99 ( .B1(n626), .B2(n1169), .A(n1161), .ZN(n870) );
  NAND2_X1 U100 ( .A1(\mem[4][7] ), .A2(n1169), .ZN(n1161) );
  OAI21_X1 U101 ( .B1(n619), .B2(n1149), .A(n1148), .ZN(n861) );
  NAND2_X1 U102 ( .A1(\mem[6][0] ), .A2(n1149), .ZN(n1148) );
  OAI21_X1 U103 ( .B1(n620), .B2(n1149), .A(n1147), .ZN(n860) );
  NAND2_X1 U104 ( .A1(\mem[6][1] ), .A2(n1149), .ZN(n1147) );
  OAI21_X1 U105 ( .B1(n621), .B2(n1149), .A(n1146), .ZN(n859) );
  NAND2_X1 U106 ( .A1(\mem[6][2] ), .A2(n1149), .ZN(n1146) );
  OAI21_X1 U107 ( .B1(n622), .B2(n1149), .A(n1145), .ZN(n858) );
  NAND2_X1 U108 ( .A1(\mem[6][3] ), .A2(n1149), .ZN(n1145) );
  OAI21_X1 U109 ( .B1(n623), .B2(n1149), .A(n1144), .ZN(n857) );
  NAND2_X1 U110 ( .A1(\mem[6][4] ), .A2(n1149), .ZN(n1144) );
  OAI21_X1 U111 ( .B1(n624), .B2(n1149), .A(n1143), .ZN(n856) );
  NAND2_X1 U112 ( .A1(\mem[6][5] ), .A2(n1149), .ZN(n1143) );
  OAI21_X1 U113 ( .B1(n625), .B2(n1149), .A(n1142), .ZN(n855) );
  NAND2_X1 U114 ( .A1(\mem[6][6] ), .A2(n1149), .ZN(n1142) );
  OAI21_X1 U115 ( .B1(n626), .B2(n1149), .A(n1141), .ZN(n854) );
  NAND2_X1 U116 ( .A1(\mem[6][7] ), .A2(n1149), .ZN(n1141) );
  OAI21_X1 U117 ( .B1(n619), .B2(n1139), .A(n1138), .ZN(n853) );
  NAND2_X1 U118 ( .A1(\mem[7][0] ), .A2(n1139), .ZN(n1138) );
  OAI21_X1 U119 ( .B1(n620), .B2(n1139), .A(n1137), .ZN(n852) );
  NAND2_X1 U120 ( .A1(\mem[7][1] ), .A2(n1139), .ZN(n1137) );
  OAI21_X1 U121 ( .B1(n621), .B2(n1139), .A(n1136), .ZN(n851) );
  NAND2_X1 U122 ( .A1(\mem[7][2] ), .A2(n1139), .ZN(n1136) );
  OAI21_X1 U123 ( .B1(n622), .B2(n1139), .A(n1135), .ZN(n850) );
  NAND2_X1 U124 ( .A1(\mem[7][3] ), .A2(n1139), .ZN(n1135) );
  OAI21_X1 U125 ( .B1(n623), .B2(n1139), .A(n1134), .ZN(n849) );
  NAND2_X1 U126 ( .A1(\mem[7][4] ), .A2(n1139), .ZN(n1134) );
  OAI21_X1 U127 ( .B1(n624), .B2(n1139), .A(n1133), .ZN(n848) );
  NAND2_X1 U128 ( .A1(\mem[7][5] ), .A2(n1139), .ZN(n1133) );
  OAI21_X1 U129 ( .B1(n625), .B2(n1139), .A(n1132), .ZN(n847) );
  NAND2_X1 U130 ( .A1(\mem[7][6] ), .A2(n1139), .ZN(n1132) );
  OAI21_X1 U131 ( .B1(n626), .B2(n1139), .A(n1131), .ZN(n846) );
  NAND2_X1 U132 ( .A1(\mem[7][7] ), .A2(n1139), .ZN(n1131) );
  OAI21_X1 U133 ( .B1(n619), .B2(n1199), .A(n1198), .ZN(n901) );
  NAND2_X1 U134 ( .A1(\mem[1][0] ), .A2(n1199), .ZN(n1198) );
  OAI21_X1 U135 ( .B1(n620), .B2(n1199), .A(n1197), .ZN(n900) );
  NAND2_X1 U136 ( .A1(\mem[1][1] ), .A2(n1199), .ZN(n1197) );
  OAI21_X1 U137 ( .B1(n621), .B2(n1199), .A(n1196), .ZN(n899) );
  NAND2_X1 U138 ( .A1(\mem[1][2] ), .A2(n1199), .ZN(n1196) );
  OAI21_X1 U139 ( .B1(n622), .B2(n1199), .A(n1195), .ZN(n898) );
  NAND2_X1 U140 ( .A1(\mem[1][3] ), .A2(n1199), .ZN(n1195) );
  OAI21_X1 U141 ( .B1(n623), .B2(n1199), .A(n1194), .ZN(n897) );
  NAND2_X1 U142 ( .A1(\mem[1][4] ), .A2(n1199), .ZN(n1194) );
  OAI21_X1 U143 ( .B1(n624), .B2(n1199), .A(n1193), .ZN(n896) );
  NAND2_X1 U144 ( .A1(\mem[1][5] ), .A2(n1199), .ZN(n1193) );
  OAI21_X1 U145 ( .B1(n625), .B2(n1199), .A(n1192), .ZN(n895) );
  NAND2_X1 U146 ( .A1(\mem[1][6] ), .A2(n1199), .ZN(n1192) );
  OAI21_X1 U147 ( .B1(n626), .B2(n1199), .A(n1191), .ZN(n894) );
  NAND2_X1 U148 ( .A1(\mem[1][7] ), .A2(n1199), .ZN(n1191) );
  OAI21_X1 U149 ( .B1(n619), .B2(n1189), .A(n1188), .ZN(n893) );
  NAND2_X1 U150 ( .A1(\mem[2][0] ), .A2(n1189), .ZN(n1188) );
  OAI21_X1 U151 ( .B1(n620), .B2(n1189), .A(n1187), .ZN(n892) );
  NAND2_X1 U152 ( .A1(\mem[2][1] ), .A2(n1189), .ZN(n1187) );
  OAI21_X1 U153 ( .B1(n621), .B2(n1189), .A(n1186), .ZN(n891) );
  NAND2_X1 U154 ( .A1(\mem[2][2] ), .A2(n1189), .ZN(n1186) );
  OAI21_X1 U155 ( .B1(n622), .B2(n1189), .A(n1185), .ZN(n890) );
  NAND2_X1 U156 ( .A1(\mem[2][3] ), .A2(n1189), .ZN(n1185) );
  OAI21_X1 U157 ( .B1(n623), .B2(n1189), .A(n1184), .ZN(n889) );
  NAND2_X1 U158 ( .A1(\mem[2][4] ), .A2(n1189), .ZN(n1184) );
  OAI21_X1 U159 ( .B1(n624), .B2(n1189), .A(n1183), .ZN(n888) );
  NAND2_X1 U160 ( .A1(\mem[2][5] ), .A2(n1189), .ZN(n1183) );
  OAI21_X1 U161 ( .B1(n625), .B2(n1189), .A(n1182), .ZN(n887) );
  NAND2_X1 U162 ( .A1(\mem[2][6] ), .A2(n1189), .ZN(n1182) );
  OAI21_X1 U163 ( .B1(n626), .B2(n1189), .A(n1181), .ZN(n886) );
  NAND2_X1 U164 ( .A1(\mem[2][7] ), .A2(n1189), .ZN(n1181) );
  OAI21_X1 U165 ( .B1(n619), .B2(n1179), .A(n1178), .ZN(n885) );
  NAND2_X1 U166 ( .A1(\mem[3][0] ), .A2(n1179), .ZN(n1178) );
  OAI21_X1 U167 ( .B1(n620), .B2(n1179), .A(n1177), .ZN(n884) );
  NAND2_X1 U168 ( .A1(\mem[3][1] ), .A2(n1179), .ZN(n1177) );
  OAI21_X1 U169 ( .B1(n621), .B2(n1179), .A(n1176), .ZN(n883) );
  NAND2_X1 U170 ( .A1(\mem[3][2] ), .A2(n1179), .ZN(n1176) );
  OAI21_X1 U171 ( .B1(n622), .B2(n1179), .A(n1175), .ZN(n882) );
  NAND2_X1 U172 ( .A1(\mem[3][3] ), .A2(n1179), .ZN(n1175) );
  OAI21_X1 U173 ( .B1(n623), .B2(n1179), .A(n1174), .ZN(n881) );
  NAND2_X1 U174 ( .A1(\mem[3][4] ), .A2(n1179), .ZN(n1174) );
  OAI21_X1 U175 ( .B1(n624), .B2(n1179), .A(n1173), .ZN(n880) );
  NAND2_X1 U176 ( .A1(\mem[3][5] ), .A2(n1179), .ZN(n1173) );
  OAI21_X1 U177 ( .B1(n625), .B2(n1179), .A(n1172), .ZN(n879) );
  NAND2_X1 U178 ( .A1(\mem[3][6] ), .A2(n1179), .ZN(n1172) );
  OAI21_X1 U179 ( .B1(n626), .B2(n1179), .A(n1171), .ZN(n878) );
  NAND2_X1 U180 ( .A1(\mem[3][7] ), .A2(n1179), .ZN(n1171) );
  OAI21_X1 U181 ( .B1(n619), .B2(n1159), .A(n1158), .ZN(n869) );
  NAND2_X1 U182 ( .A1(\mem[5][0] ), .A2(n1159), .ZN(n1158) );
  OAI21_X1 U183 ( .B1(n620), .B2(n1159), .A(n1157), .ZN(n868) );
  NAND2_X1 U184 ( .A1(\mem[5][1] ), .A2(n1159), .ZN(n1157) );
  OAI21_X1 U185 ( .B1(n621), .B2(n1159), .A(n1156), .ZN(n867) );
  NAND2_X1 U186 ( .A1(\mem[5][2] ), .A2(n1159), .ZN(n1156) );
  OAI21_X1 U187 ( .B1(n622), .B2(n1159), .A(n1155), .ZN(n866) );
  NAND2_X1 U188 ( .A1(\mem[5][3] ), .A2(n1159), .ZN(n1155) );
  OAI21_X1 U189 ( .B1(n623), .B2(n1159), .A(n1154), .ZN(n865) );
  NAND2_X1 U190 ( .A1(\mem[5][4] ), .A2(n1159), .ZN(n1154) );
  OAI21_X1 U191 ( .B1(n624), .B2(n1159), .A(n1153), .ZN(n864) );
  NAND2_X1 U192 ( .A1(\mem[5][5] ), .A2(n1159), .ZN(n1153) );
  OAI21_X1 U193 ( .B1(n625), .B2(n1159), .A(n1152), .ZN(n863) );
  NAND2_X1 U194 ( .A1(\mem[5][6] ), .A2(n1159), .ZN(n1152) );
  OAI21_X1 U195 ( .B1(n626), .B2(n1159), .A(n1151), .ZN(n862) );
  NAND2_X1 U196 ( .A1(\mem[5][7] ), .A2(n1159), .ZN(n1151) );
  OAI21_X1 U197 ( .B1(n1210), .B2(n619), .A(n1209), .ZN(n909) );
  NAND2_X1 U198 ( .A1(\mem[0][0] ), .A2(n1210), .ZN(n1209) );
  OAI21_X1 U199 ( .B1(n1210), .B2(n620), .A(n1208), .ZN(n908) );
  NAND2_X1 U200 ( .A1(\mem[0][1] ), .A2(n1210), .ZN(n1208) );
  OAI21_X1 U201 ( .B1(n1210), .B2(n621), .A(n1207), .ZN(n907) );
  NAND2_X1 U202 ( .A1(\mem[0][2] ), .A2(n1210), .ZN(n1207) );
  OAI21_X1 U203 ( .B1(n1210), .B2(n622), .A(n1206), .ZN(n906) );
  NAND2_X1 U204 ( .A1(\mem[0][3] ), .A2(n1210), .ZN(n1206) );
  OAI21_X1 U205 ( .B1(n1210), .B2(n623), .A(n1205), .ZN(n905) );
  NAND2_X1 U206 ( .A1(\mem[0][4] ), .A2(n1210), .ZN(n1205) );
  OAI21_X1 U207 ( .B1(n1210), .B2(n624), .A(n1204), .ZN(n904) );
  NAND2_X1 U208 ( .A1(\mem[0][5] ), .A2(n1210), .ZN(n1204) );
  OAI21_X1 U209 ( .B1(n1210), .B2(n625), .A(n1203), .ZN(n903) );
  NAND2_X1 U210 ( .A1(\mem[0][6] ), .A2(n1210), .ZN(n1203) );
  OAI21_X1 U211 ( .B1(n1210), .B2(n626), .A(n1202), .ZN(n902) );
  NAND2_X1 U212 ( .A1(\mem[0][7] ), .A2(n1210), .ZN(n1202) );
  INV_X1 U213 ( .A(n1128), .ZN(n818) );
  AOI22_X1 U214 ( .A1(data_in[0]), .A2(n842), .B1(n1127), .B2(\mem[8][0] ), 
        .ZN(n1128) );
  INV_X1 U215 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U216 ( .A1(data_in[1]), .A2(n842), .B1(n1127), .B2(\mem[8][1] ), 
        .ZN(n1126) );
  INV_X1 U217 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U218 ( .A1(data_in[2]), .A2(n842), .B1(n1127), .B2(\mem[8][2] ), 
        .ZN(n1125) );
  INV_X1 U219 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U220 ( .A1(data_in[3]), .A2(n842), .B1(n1127), .B2(\mem[8][3] ), 
        .ZN(n1124) );
  INV_X1 U221 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U222 ( .A1(data_in[4]), .A2(n842), .B1(n1127), .B2(\mem[8][4] ), 
        .ZN(n1123) );
  INV_X1 U223 ( .A(n1122), .ZN(n813) );
  AOI22_X1 U224 ( .A1(data_in[5]), .A2(n842), .B1(n1127), .B2(\mem[8][5] ), 
        .ZN(n1122) );
  INV_X1 U225 ( .A(n1121), .ZN(n812) );
  AOI22_X1 U226 ( .A1(data_in[6]), .A2(n842), .B1(n1127), .B2(\mem[8][6] ), 
        .ZN(n1121) );
  INV_X1 U227 ( .A(n1120), .ZN(n811) );
  AOI22_X1 U228 ( .A1(data_in[7]), .A2(n842), .B1(n1127), .B2(\mem[8][7] ), 
        .ZN(n1120) );
  INV_X1 U229 ( .A(n1118), .ZN(n810) );
  AOI22_X1 U230 ( .A1(data_in[0]), .A2(n841), .B1(n1117), .B2(\mem[9][0] ), 
        .ZN(n1118) );
  INV_X1 U231 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U232 ( .A1(data_in[1]), .A2(n841), .B1(n1117), .B2(\mem[9][1] ), 
        .ZN(n1116) );
  INV_X1 U233 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U234 ( .A1(data_in[2]), .A2(n841), .B1(n1117), .B2(\mem[9][2] ), 
        .ZN(n1115) );
  INV_X1 U235 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U236 ( .A1(data_in[3]), .A2(n841), .B1(n1117), .B2(\mem[9][3] ), 
        .ZN(n1114) );
  INV_X1 U237 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U238 ( .A1(data_in[4]), .A2(n841), .B1(n1117), .B2(\mem[9][4] ), 
        .ZN(n1113) );
  INV_X1 U239 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U240 ( .A1(data_in[5]), .A2(n841), .B1(n1117), .B2(\mem[9][5] ), 
        .ZN(n1112) );
  INV_X1 U241 ( .A(n1111), .ZN(n804) );
  AOI22_X1 U242 ( .A1(data_in[6]), .A2(n841), .B1(n1117), .B2(\mem[9][6] ), 
        .ZN(n1111) );
  INV_X1 U243 ( .A(n1110), .ZN(n803) );
  AOI22_X1 U244 ( .A1(data_in[7]), .A2(n841), .B1(n1117), .B2(\mem[9][7] ), 
        .ZN(n1110) );
  INV_X1 U245 ( .A(n1109), .ZN(n802) );
  AOI22_X1 U246 ( .A1(data_in[0]), .A2(n840), .B1(n1108), .B2(\mem[10][0] ), 
        .ZN(n1109) );
  INV_X1 U247 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U248 ( .A1(data_in[1]), .A2(n840), .B1(n1108), .B2(\mem[10][1] ), 
        .ZN(n1107) );
  INV_X1 U249 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U250 ( .A1(data_in[2]), .A2(n840), .B1(n1108), .B2(\mem[10][2] ), 
        .ZN(n1106) );
  INV_X1 U251 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U252 ( .A1(data_in[3]), .A2(n840), .B1(n1108), .B2(\mem[10][3] ), 
        .ZN(n1105) );
  INV_X1 U253 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U254 ( .A1(data_in[4]), .A2(n840), .B1(n1108), .B2(\mem[10][4] ), 
        .ZN(n1104) );
  INV_X1 U255 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U256 ( .A1(data_in[5]), .A2(n840), .B1(n1108), .B2(\mem[10][5] ), 
        .ZN(n1103) );
  INV_X1 U257 ( .A(n1102), .ZN(n796) );
  AOI22_X1 U258 ( .A1(data_in[6]), .A2(n840), .B1(n1108), .B2(\mem[10][6] ), 
        .ZN(n1102) );
  INV_X1 U259 ( .A(n1101), .ZN(n795) );
  AOI22_X1 U260 ( .A1(data_in[7]), .A2(n840), .B1(n1108), .B2(\mem[10][7] ), 
        .ZN(n1101) );
  INV_X1 U261 ( .A(n1100), .ZN(n794) );
  AOI22_X1 U262 ( .A1(data_in[0]), .A2(n839), .B1(n1099), .B2(\mem[11][0] ), 
        .ZN(n1100) );
  INV_X1 U263 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U264 ( .A1(data_in[1]), .A2(n839), .B1(n1099), .B2(\mem[11][1] ), 
        .ZN(n1098) );
  INV_X1 U265 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U266 ( .A1(data_in[2]), .A2(n839), .B1(n1099), .B2(\mem[11][2] ), 
        .ZN(n1097) );
  INV_X1 U267 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U268 ( .A1(data_in[3]), .A2(n839), .B1(n1099), .B2(\mem[11][3] ), 
        .ZN(n1096) );
  INV_X1 U269 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U270 ( .A1(data_in[4]), .A2(n839), .B1(n1099), .B2(\mem[11][4] ), 
        .ZN(n1095) );
  INV_X1 U271 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U272 ( .A1(data_in[5]), .A2(n839), .B1(n1099), .B2(\mem[11][5] ), 
        .ZN(n1094) );
  INV_X1 U273 ( .A(n1093), .ZN(n788) );
  AOI22_X1 U274 ( .A1(data_in[6]), .A2(n839), .B1(n1099), .B2(\mem[11][6] ), 
        .ZN(n1093) );
  INV_X1 U275 ( .A(n1092), .ZN(n787) );
  AOI22_X1 U276 ( .A1(data_in[7]), .A2(n839), .B1(n1099), .B2(\mem[11][7] ), 
        .ZN(n1092) );
  INV_X1 U277 ( .A(n1091), .ZN(n786) );
  AOI22_X1 U278 ( .A1(data_in[0]), .A2(n838), .B1(n1090), .B2(\mem[12][0] ), 
        .ZN(n1091) );
  INV_X1 U279 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U280 ( .A1(data_in[1]), .A2(n838), .B1(n1090), .B2(\mem[12][1] ), 
        .ZN(n1089) );
  INV_X1 U281 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U282 ( .A1(data_in[2]), .A2(n838), .B1(n1090), .B2(\mem[12][2] ), 
        .ZN(n1088) );
  INV_X1 U283 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U284 ( .A1(data_in[3]), .A2(n838), .B1(n1090), .B2(\mem[12][3] ), 
        .ZN(n1087) );
  INV_X1 U285 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U286 ( .A1(data_in[4]), .A2(n838), .B1(n1090), .B2(\mem[12][4] ), 
        .ZN(n1086) );
  INV_X1 U287 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U288 ( .A1(data_in[5]), .A2(n838), .B1(n1090), .B2(\mem[12][5] ), 
        .ZN(n1085) );
  INV_X1 U289 ( .A(n1084), .ZN(n780) );
  AOI22_X1 U290 ( .A1(data_in[6]), .A2(n838), .B1(n1090), .B2(\mem[12][6] ), 
        .ZN(n1084) );
  INV_X1 U291 ( .A(n1083), .ZN(n779) );
  AOI22_X1 U292 ( .A1(data_in[7]), .A2(n838), .B1(n1090), .B2(\mem[12][7] ), 
        .ZN(n1083) );
  INV_X1 U293 ( .A(n1082), .ZN(n778) );
  AOI22_X1 U294 ( .A1(data_in[0]), .A2(n837), .B1(n1081), .B2(\mem[13][0] ), 
        .ZN(n1082) );
  INV_X1 U295 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U296 ( .A1(data_in[1]), .A2(n837), .B1(n1081), .B2(\mem[13][1] ), 
        .ZN(n1080) );
  INV_X1 U297 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U298 ( .A1(data_in[2]), .A2(n837), .B1(n1081), .B2(\mem[13][2] ), 
        .ZN(n1079) );
  INV_X1 U299 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U300 ( .A1(data_in[3]), .A2(n837), .B1(n1081), .B2(\mem[13][3] ), 
        .ZN(n1078) );
  INV_X1 U301 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U302 ( .A1(data_in[4]), .A2(n837), .B1(n1081), .B2(\mem[13][4] ), 
        .ZN(n1077) );
  INV_X1 U303 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U304 ( .A1(data_in[5]), .A2(n837), .B1(n1081), .B2(\mem[13][5] ), 
        .ZN(n1076) );
  INV_X1 U305 ( .A(n1075), .ZN(n772) );
  AOI22_X1 U306 ( .A1(data_in[6]), .A2(n837), .B1(n1081), .B2(\mem[13][6] ), 
        .ZN(n1075) );
  INV_X1 U307 ( .A(n1074), .ZN(n771) );
  AOI22_X1 U308 ( .A1(data_in[7]), .A2(n837), .B1(n1081), .B2(\mem[13][7] ), 
        .ZN(n1074) );
  INV_X1 U309 ( .A(n1073), .ZN(n770) );
  AOI22_X1 U310 ( .A1(data_in[0]), .A2(n836), .B1(n1072), .B2(\mem[14][0] ), 
        .ZN(n1073) );
  INV_X1 U311 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U312 ( .A1(data_in[1]), .A2(n836), .B1(n1072), .B2(\mem[14][1] ), 
        .ZN(n1071) );
  INV_X1 U313 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U314 ( .A1(data_in[2]), .A2(n836), .B1(n1072), .B2(\mem[14][2] ), 
        .ZN(n1070) );
  INV_X1 U315 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U316 ( .A1(data_in[3]), .A2(n836), .B1(n1072), .B2(\mem[14][3] ), 
        .ZN(n1069) );
  INV_X1 U317 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U318 ( .A1(data_in[4]), .A2(n836), .B1(n1072), .B2(\mem[14][4] ), 
        .ZN(n1068) );
  INV_X1 U319 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U320 ( .A1(data_in[5]), .A2(n836), .B1(n1072), .B2(\mem[14][5] ), 
        .ZN(n1067) );
  INV_X1 U321 ( .A(n1066), .ZN(n764) );
  AOI22_X1 U322 ( .A1(data_in[6]), .A2(n836), .B1(n1072), .B2(\mem[14][6] ), 
        .ZN(n1066) );
  INV_X1 U323 ( .A(n1065), .ZN(n763) );
  AOI22_X1 U324 ( .A1(data_in[7]), .A2(n836), .B1(n1072), .B2(\mem[14][7] ), 
        .ZN(n1065) );
  INV_X1 U325 ( .A(n1064), .ZN(n762) );
  AOI22_X1 U326 ( .A1(data_in[0]), .A2(n835), .B1(n1063), .B2(\mem[15][0] ), 
        .ZN(n1064) );
  INV_X1 U327 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U328 ( .A1(data_in[1]), .A2(n835), .B1(n1063), .B2(\mem[15][1] ), 
        .ZN(n1062) );
  INV_X1 U329 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U330 ( .A1(data_in[2]), .A2(n835), .B1(n1063), .B2(\mem[15][2] ), 
        .ZN(n1061) );
  INV_X1 U331 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U332 ( .A1(data_in[3]), .A2(n835), .B1(n1063), .B2(\mem[15][3] ), 
        .ZN(n1060) );
  INV_X1 U333 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U334 ( .A1(data_in[4]), .A2(n835), .B1(n1063), .B2(\mem[15][4] ), 
        .ZN(n1059) );
  INV_X1 U335 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U336 ( .A1(data_in[5]), .A2(n835), .B1(n1063), .B2(\mem[15][5] ), 
        .ZN(n1058) );
  INV_X1 U337 ( .A(n1057), .ZN(n756) );
  AOI22_X1 U338 ( .A1(data_in[6]), .A2(n835), .B1(n1063), .B2(\mem[15][6] ), 
        .ZN(n1057) );
  INV_X1 U339 ( .A(n1056), .ZN(n755) );
  AOI22_X1 U340 ( .A1(data_in[7]), .A2(n835), .B1(n1063), .B2(\mem[15][7] ), 
        .ZN(n1056) );
  INV_X1 U341 ( .A(n1055), .ZN(n754) );
  AOI22_X1 U342 ( .A1(data_in[0]), .A2(n834), .B1(n1054), .B2(\mem[16][0] ), 
        .ZN(n1055) );
  INV_X1 U343 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U344 ( .A1(data_in[1]), .A2(n834), .B1(n1054), .B2(\mem[16][1] ), 
        .ZN(n1053) );
  INV_X1 U345 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U346 ( .A1(data_in[2]), .A2(n834), .B1(n1054), .B2(\mem[16][2] ), 
        .ZN(n1052) );
  INV_X1 U347 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U348 ( .A1(data_in[3]), .A2(n834), .B1(n1054), .B2(\mem[16][3] ), 
        .ZN(n1051) );
  INV_X1 U349 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U350 ( .A1(data_in[4]), .A2(n834), .B1(n1054), .B2(\mem[16][4] ), 
        .ZN(n1050) );
  INV_X1 U351 ( .A(n1049), .ZN(n749) );
  AOI22_X1 U352 ( .A1(data_in[5]), .A2(n834), .B1(n1054), .B2(\mem[16][5] ), 
        .ZN(n1049) );
  INV_X1 U353 ( .A(n1048), .ZN(n748) );
  AOI22_X1 U354 ( .A1(data_in[6]), .A2(n834), .B1(n1054), .B2(\mem[16][6] ), 
        .ZN(n1048) );
  INV_X1 U355 ( .A(n1047), .ZN(n747) );
  AOI22_X1 U356 ( .A1(data_in[7]), .A2(n834), .B1(n1054), .B2(\mem[16][7] ), 
        .ZN(n1047) );
  INV_X1 U357 ( .A(n1045), .ZN(n746) );
  AOI22_X1 U358 ( .A1(data_in[0]), .A2(n833), .B1(n1044), .B2(\mem[17][0] ), 
        .ZN(n1045) );
  INV_X1 U359 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U360 ( .A1(data_in[1]), .A2(n833), .B1(n1044), .B2(\mem[17][1] ), 
        .ZN(n1043) );
  INV_X1 U361 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U362 ( .A1(data_in[2]), .A2(n833), .B1(n1044), .B2(\mem[17][2] ), 
        .ZN(n1042) );
  INV_X1 U363 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U364 ( .A1(data_in[3]), .A2(n833), .B1(n1044), .B2(\mem[17][3] ), 
        .ZN(n1041) );
  INV_X1 U365 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U366 ( .A1(data_in[4]), .A2(n833), .B1(n1044), .B2(\mem[17][4] ), 
        .ZN(n1040) );
  INV_X1 U367 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U368 ( .A1(data_in[5]), .A2(n833), .B1(n1044), .B2(\mem[17][5] ), 
        .ZN(n1039) );
  INV_X1 U369 ( .A(n1038), .ZN(n740) );
  AOI22_X1 U370 ( .A1(data_in[6]), .A2(n833), .B1(n1044), .B2(\mem[17][6] ), 
        .ZN(n1038) );
  INV_X1 U371 ( .A(n1037), .ZN(n739) );
  AOI22_X1 U372 ( .A1(data_in[7]), .A2(n833), .B1(n1044), .B2(\mem[17][7] ), 
        .ZN(n1037) );
  INV_X1 U373 ( .A(n1036), .ZN(n738) );
  AOI22_X1 U374 ( .A1(data_in[0]), .A2(n832), .B1(n1035), .B2(\mem[18][0] ), 
        .ZN(n1036) );
  INV_X1 U375 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U376 ( .A1(data_in[1]), .A2(n832), .B1(n1035), .B2(\mem[18][1] ), 
        .ZN(n1034) );
  INV_X1 U377 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U378 ( .A1(data_in[2]), .A2(n832), .B1(n1035), .B2(\mem[18][2] ), 
        .ZN(n1033) );
  INV_X1 U379 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U380 ( .A1(data_in[3]), .A2(n832), .B1(n1035), .B2(\mem[18][3] ), 
        .ZN(n1032) );
  INV_X1 U381 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U382 ( .A1(data_in[4]), .A2(n832), .B1(n1035), .B2(\mem[18][4] ), 
        .ZN(n1031) );
  INV_X1 U383 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U384 ( .A1(data_in[5]), .A2(n832), .B1(n1035), .B2(\mem[18][5] ), 
        .ZN(n1030) );
  INV_X1 U385 ( .A(n1029), .ZN(n732) );
  AOI22_X1 U386 ( .A1(data_in[6]), .A2(n832), .B1(n1035), .B2(\mem[18][6] ), 
        .ZN(n1029) );
  INV_X1 U387 ( .A(n1028), .ZN(n731) );
  AOI22_X1 U388 ( .A1(data_in[7]), .A2(n832), .B1(n1035), .B2(\mem[18][7] ), 
        .ZN(n1028) );
  INV_X1 U389 ( .A(n1027), .ZN(n730) );
  AOI22_X1 U390 ( .A1(data_in[0]), .A2(n831), .B1(n1026), .B2(\mem[19][0] ), 
        .ZN(n1027) );
  INV_X1 U391 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U392 ( .A1(data_in[1]), .A2(n831), .B1(n1026), .B2(\mem[19][1] ), 
        .ZN(n1025) );
  INV_X1 U393 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U394 ( .A1(data_in[2]), .A2(n831), .B1(n1026), .B2(\mem[19][2] ), 
        .ZN(n1024) );
  INV_X1 U395 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U396 ( .A1(data_in[3]), .A2(n831), .B1(n1026), .B2(\mem[19][3] ), 
        .ZN(n1023) );
  INV_X1 U397 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U398 ( .A1(data_in[4]), .A2(n831), .B1(n1026), .B2(\mem[19][4] ), 
        .ZN(n1022) );
  INV_X1 U399 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U400 ( .A1(data_in[5]), .A2(n831), .B1(n1026), .B2(\mem[19][5] ), 
        .ZN(n1021) );
  INV_X1 U401 ( .A(n1020), .ZN(n724) );
  AOI22_X1 U402 ( .A1(data_in[6]), .A2(n831), .B1(n1026), .B2(\mem[19][6] ), 
        .ZN(n1020) );
  INV_X1 U403 ( .A(n1019), .ZN(n723) );
  AOI22_X1 U404 ( .A1(data_in[7]), .A2(n831), .B1(n1026), .B2(\mem[19][7] ), 
        .ZN(n1019) );
  INV_X1 U405 ( .A(n1018), .ZN(n722) );
  AOI22_X1 U406 ( .A1(data_in[0]), .A2(n830), .B1(n1017), .B2(\mem[20][0] ), 
        .ZN(n1018) );
  INV_X1 U407 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U408 ( .A1(data_in[1]), .A2(n830), .B1(n1017), .B2(\mem[20][1] ), 
        .ZN(n1016) );
  INV_X1 U409 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U410 ( .A1(data_in[2]), .A2(n830), .B1(n1017), .B2(\mem[20][2] ), 
        .ZN(n1015) );
  INV_X1 U411 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U412 ( .A1(data_in[3]), .A2(n830), .B1(n1017), .B2(\mem[20][3] ), 
        .ZN(n1014) );
  INV_X1 U413 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U414 ( .A1(data_in[4]), .A2(n830), .B1(n1017), .B2(\mem[20][4] ), 
        .ZN(n1013) );
  INV_X1 U415 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U416 ( .A1(data_in[5]), .A2(n830), .B1(n1017), .B2(\mem[20][5] ), 
        .ZN(n1012) );
  INV_X1 U417 ( .A(n1011), .ZN(n716) );
  AOI22_X1 U418 ( .A1(data_in[6]), .A2(n830), .B1(n1017), .B2(\mem[20][6] ), 
        .ZN(n1011) );
  INV_X1 U419 ( .A(n1010), .ZN(n715) );
  AOI22_X1 U420 ( .A1(data_in[7]), .A2(n830), .B1(n1017), .B2(\mem[20][7] ), 
        .ZN(n1010) );
  INV_X1 U421 ( .A(n1009), .ZN(n714) );
  AOI22_X1 U422 ( .A1(data_in[0]), .A2(n829), .B1(n1008), .B2(\mem[21][0] ), 
        .ZN(n1009) );
  INV_X1 U423 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U424 ( .A1(data_in[1]), .A2(n829), .B1(n1008), .B2(\mem[21][1] ), 
        .ZN(n1007) );
  INV_X1 U425 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U426 ( .A1(data_in[2]), .A2(n829), .B1(n1008), .B2(\mem[21][2] ), 
        .ZN(n1006) );
  INV_X1 U427 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U428 ( .A1(data_in[3]), .A2(n829), .B1(n1008), .B2(\mem[21][3] ), 
        .ZN(n1005) );
  INV_X1 U429 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U430 ( .A1(data_in[4]), .A2(n829), .B1(n1008), .B2(\mem[21][4] ), 
        .ZN(n1004) );
  INV_X1 U431 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U432 ( .A1(data_in[5]), .A2(n829), .B1(n1008), .B2(\mem[21][5] ), 
        .ZN(n1003) );
  INV_X1 U433 ( .A(n1002), .ZN(n708) );
  AOI22_X1 U434 ( .A1(data_in[6]), .A2(n829), .B1(n1008), .B2(\mem[21][6] ), 
        .ZN(n1002) );
  INV_X1 U435 ( .A(n1001), .ZN(n707) );
  AOI22_X1 U436 ( .A1(data_in[7]), .A2(n829), .B1(n1008), .B2(\mem[21][7] ), 
        .ZN(n1001) );
  INV_X1 U437 ( .A(n1000), .ZN(n706) );
  AOI22_X1 U438 ( .A1(data_in[0]), .A2(n828), .B1(n999), .B2(\mem[22][0] ), 
        .ZN(n1000) );
  INV_X1 U439 ( .A(n998), .ZN(n705) );
  AOI22_X1 U440 ( .A1(data_in[1]), .A2(n828), .B1(n999), .B2(\mem[22][1] ), 
        .ZN(n998) );
  INV_X1 U441 ( .A(n997), .ZN(n704) );
  AOI22_X1 U442 ( .A1(data_in[2]), .A2(n828), .B1(n999), .B2(\mem[22][2] ), 
        .ZN(n997) );
  INV_X1 U443 ( .A(n996), .ZN(n703) );
  AOI22_X1 U444 ( .A1(data_in[3]), .A2(n828), .B1(n999), .B2(\mem[22][3] ), 
        .ZN(n996) );
  INV_X1 U445 ( .A(n995), .ZN(n702) );
  AOI22_X1 U446 ( .A1(data_in[4]), .A2(n828), .B1(n999), .B2(\mem[22][4] ), 
        .ZN(n995) );
  INV_X1 U447 ( .A(n994), .ZN(n701) );
  AOI22_X1 U448 ( .A1(data_in[5]), .A2(n828), .B1(n999), .B2(\mem[22][5] ), 
        .ZN(n994) );
  INV_X1 U449 ( .A(n993), .ZN(n700) );
  AOI22_X1 U450 ( .A1(data_in[6]), .A2(n828), .B1(n999), .B2(\mem[22][6] ), 
        .ZN(n993) );
  INV_X1 U451 ( .A(n992), .ZN(n699) );
  AOI22_X1 U452 ( .A1(data_in[7]), .A2(n828), .B1(n999), .B2(\mem[22][7] ), 
        .ZN(n992) );
  INV_X1 U453 ( .A(n991), .ZN(n698) );
  AOI22_X1 U454 ( .A1(data_in[0]), .A2(n827), .B1(n990), .B2(\mem[23][0] ), 
        .ZN(n991) );
  INV_X1 U455 ( .A(n989), .ZN(n697) );
  AOI22_X1 U456 ( .A1(data_in[1]), .A2(n827), .B1(n990), .B2(\mem[23][1] ), 
        .ZN(n989) );
  INV_X1 U457 ( .A(n988), .ZN(n696) );
  AOI22_X1 U458 ( .A1(data_in[2]), .A2(n827), .B1(n990), .B2(\mem[23][2] ), 
        .ZN(n988) );
  INV_X1 U459 ( .A(n987), .ZN(n695) );
  AOI22_X1 U460 ( .A1(data_in[3]), .A2(n827), .B1(n990), .B2(\mem[23][3] ), 
        .ZN(n987) );
  INV_X1 U461 ( .A(n986), .ZN(n694) );
  AOI22_X1 U462 ( .A1(data_in[4]), .A2(n827), .B1(n990), .B2(\mem[23][4] ), 
        .ZN(n986) );
  INV_X1 U463 ( .A(n985), .ZN(n693) );
  AOI22_X1 U464 ( .A1(data_in[5]), .A2(n827), .B1(n990), .B2(\mem[23][5] ), 
        .ZN(n985) );
  INV_X1 U465 ( .A(n984), .ZN(n692) );
  AOI22_X1 U466 ( .A1(data_in[6]), .A2(n827), .B1(n990), .B2(\mem[23][6] ), 
        .ZN(n984) );
  INV_X1 U467 ( .A(n983), .ZN(n691) );
  AOI22_X1 U468 ( .A1(data_in[7]), .A2(n827), .B1(n990), .B2(\mem[23][7] ), 
        .ZN(n983) );
  INV_X1 U469 ( .A(n982), .ZN(n690) );
  AOI22_X1 U470 ( .A1(data_in[0]), .A2(n826), .B1(n981), .B2(\mem[24][0] ), 
        .ZN(n982) );
  INV_X1 U471 ( .A(n980), .ZN(n689) );
  AOI22_X1 U472 ( .A1(data_in[1]), .A2(n826), .B1(n981), .B2(\mem[24][1] ), 
        .ZN(n980) );
  INV_X1 U473 ( .A(n979), .ZN(n688) );
  AOI22_X1 U474 ( .A1(data_in[2]), .A2(n826), .B1(n981), .B2(\mem[24][2] ), 
        .ZN(n979) );
  INV_X1 U475 ( .A(n978), .ZN(n687) );
  AOI22_X1 U476 ( .A1(data_in[3]), .A2(n826), .B1(n981), .B2(\mem[24][3] ), 
        .ZN(n978) );
  INV_X1 U477 ( .A(n977), .ZN(n686) );
  AOI22_X1 U478 ( .A1(data_in[4]), .A2(n826), .B1(n981), .B2(\mem[24][4] ), 
        .ZN(n977) );
  INV_X1 U479 ( .A(n976), .ZN(n685) );
  AOI22_X1 U480 ( .A1(data_in[5]), .A2(n826), .B1(n981), .B2(\mem[24][5] ), 
        .ZN(n976) );
  INV_X1 U481 ( .A(n975), .ZN(n684) );
  AOI22_X1 U482 ( .A1(data_in[6]), .A2(n826), .B1(n981), .B2(\mem[24][6] ), 
        .ZN(n975) );
  INV_X1 U483 ( .A(n974), .ZN(n683) );
  AOI22_X1 U484 ( .A1(data_in[7]), .A2(n826), .B1(n981), .B2(\mem[24][7] ), 
        .ZN(n974) );
  INV_X1 U485 ( .A(n972), .ZN(n682) );
  AOI22_X1 U486 ( .A1(data_in[0]), .A2(n825), .B1(n971), .B2(\mem[25][0] ), 
        .ZN(n972) );
  INV_X1 U487 ( .A(n970), .ZN(n681) );
  AOI22_X1 U488 ( .A1(data_in[1]), .A2(n825), .B1(n971), .B2(\mem[25][1] ), 
        .ZN(n970) );
  INV_X1 U489 ( .A(n969), .ZN(n680) );
  AOI22_X1 U490 ( .A1(data_in[2]), .A2(n825), .B1(n971), .B2(\mem[25][2] ), 
        .ZN(n969) );
  INV_X1 U491 ( .A(n968), .ZN(n679) );
  AOI22_X1 U492 ( .A1(data_in[3]), .A2(n825), .B1(n971), .B2(\mem[25][3] ), 
        .ZN(n968) );
  INV_X1 U493 ( .A(n967), .ZN(n678) );
  AOI22_X1 U494 ( .A1(data_in[4]), .A2(n825), .B1(n971), .B2(\mem[25][4] ), 
        .ZN(n967) );
  INV_X1 U495 ( .A(n966), .ZN(n677) );
  AOI22_X1 U496 ( .A1(data_in[5]), .A2(n825), .B1(n971), .B2(\mem[25][5] ), 
        .ZN(n966) );
  INV_X1 U497 ( .A(n965), .ZN(n676) );
  AOI22_X1 U498 ( .A1(data_in[6]), .A2(n825), .B1(n971), .B2(\mem[25][6] ), 
        .ZN(n965) );
  INV_X1 U499 ( .A(n964), .ZN(n675) );
  AOI22_X1 U500 ( .A1(data_in[7]), .A2(n825), .B1(n971), .B2(\mem[25][7] ), 
        .ZN(n964) );
  INV_X1 U501 ( .A(n963), .ZN(n674) );
  AOI22_X1 U502 ( .A1(data_in[0]), .A2(n824), .B1(n962), .B2(\mem[26][0] ), 
        .ZN(n963) );
  INV_X1 U503 ( .A(n961), .ZN(n673) );
  AOI22_X1 U504 ( .A1(data_in[1]), .A2(n824), .B1(n962), .B2(\mem[26][1] ), 
        .ZN(n961) );
  INV_X1 U505 ( .A(n960), .ZN(n672) );
  AOI22_X1 U506 ( .A1(data_in[2]), .A2(n824), .B1(n962), .B2(\mem[26][2] ), 
        .ZN(n960) );
  INV_X1 U507 ( .A(n959), .ZN(n671) );
  AOI22_X1 U508 ( .A1(data_in[3]), .A2(n824), .B1(n962), .B2(\mem[26][3] ), 
        .ZN(n959) );
  INV_X1 U509 ( .A(n958), .ZN(n670) );
  AOI22_X1 U510 ( .A1(data_in[4]), .A2(n824), .B1(n962), .B2(\mem[26][4] ), 
        .ZN(n958) );
  INV_X1 U511 ( .A(n957), .ZN(n669) );
  AOI22_X1 U512 ( .A1(data_in[5]), .A2(n824), .B1(n962), .B2(\mem[26][5] ), 
        .ZN(n957) );
  INV_X1 U513 ( .A(n956), .ZN(n668) );
  AOI22_X1 U514 ( .A1(data_in[6]), .A2(n824), .B1(n962), .B2(\mem[26][6] ), 
        .ZN(n956) );
  INV_X1 U515 ( .A(n955), .ZN(n667) );
  AOI22_X1 U516 ( .A1(data_in[7]), .A2(n824), .B1(n962), .B2(\mem[26][7] ), 
        .ZN(n955) );
  INV_X1 U517 ( .A(n954), .ZN(n666) );
  AOI22_X1 U518 ( .A1(data_in[0]), .A2(n823), .B1(n953), .B2(\mem[27][0] ), 
        .ZN(n954) );
  INV_X1 U519 ( .A(n952), .ZN(n665) );
  AOI22_X1 U520 ( .A1(data_in[1]), .A2(n823), .B1(n953), .B2(\mem[27][1] ), 
        .ZN(n952) );
  INV_X1 U521 ( .A(n951), .ZN(n664) );
  AOI22_X1 U522 ( .A1(data_in[2]), .A2(n823), .B1(n953), .B2(\mem[27][2] ), 
        .ZN(n951) );
  INV_X1 U523 ( .A(n950), .ZN(n663) );
  AOI22_X1 U524 ( .A1(data_in[3]), .A2(n823), .B1(n953), .B2(\mem[27][3] ), 
        .ZN(n950) );
  INV_X1 U525 ( .A(n949), .ZN(n662) );
  AOI22_X1 U526 ( .A1(data_in[4]), .A2(n823), .B1(n953), .B2(\mem[27][4] ), 
        .ZN(n949) );
  INV_X1 U527 ( .A(n948), .ZN(n661) );
  AOI22_X1 U528 ( .A1(data_in[5]), .A2(n823), .B1(n953), .B2(\mem[27][5] ), 
        .ZN(n948) );
  INV_X1 U529 ( .A(n947), .ZN(n660) );
  AOI22_X1 U530 ( .A1(data_in[6]), .A2(n823), .B1(n953), .B2(\mem[27][6] ), 
        .ZN(n947) );
  INV_X1 U531 ( .A(n946), .ZN(n659) );
  AOI22_X1 U532 ( .A1(data_in[7]), .A2(n823), .B1(n953), .B2(\mem[27][7] ), 
        .ZN(n946) );
  INV_X1 U533 ( .A(n945), .ZN(n658) );
  AOI22_X1 U534 ( .A1(data_in[0]), .A2(n822), .B1(n944), .B2(\mem[28][0] ), 
        .ZN(n945) );
  INV_X1 U535 ( .A(n943), .ZN(n657) );
  AOI22_X1 U536 ( .A1(data_in[1]), .A2(n822), .B1(n944), .B2(\mem[28][1] ), 
        .ZN(n943) );
  INV_X1 U537 ( .A(n942), .ZN(n656) );
  AOI22_X1 U538 ( .A1(data_in[2]), .A2(n822), .B1(n944), .B2(\mem[28][2] ), 
        .ZN(n942) );
  INV_X1 U539 ( .A(n941), .ZN(n655) );
  AOI22_X1 U540 ( .A1(data_in[3]), .A2(n822), .B1(n944), .B2(\mem[28][3] ), 
        .ZN(n941) );
  INV_X1 U541 ( .A(n940), .ZN(n654) );
  AOI22_X1 U542 ( .A1(data_in[4]), .A2(n822), .B1(n944), .B2(\mem[28][4] ), 
        .ZN(n940) );
  INV_X1 U543 ( .A(n939), .ZN(n653) );
  AOI22_X1 U544 ( .A1(data_in[5]), .A2(n822), .B1(n944), .B2(\mem[28][5] ), 
        .ZN(n939) );
  INV_X1 U545 ( .A(n938), .ZN(n652) );
  AOI22_X1 U546 ( .A1(data_in[6]), .A2(n822), .B1(n944), .B2(\mem[28][6] ), 
        .ZN(n938) );
  INV_X1 U547 ( .A(n937), .ZN(n651) );
  AOI22_X1 U548 ( .A1(data_in[7]), .A2(n822), .B1(n944), .B2(\mem[28][7] ), 
        .ZN(n937) );
  INV_X1 U549 ( .A(n936), .ZN(n650) );
  AOI22_X1 U550 ( .A1(data_in[0]), .A2(n821), .B1(n935), .B2(\mem[29][0] ), 
        .ZN(n936) );
  INV_X1 U551 ( .A(n934), .ZN(n649) );
  AOI22_X1 U552 ( .A1(data_in[1]), .A2(n821), .B1(n935), .B2(\mem[29][1] ), 
        .ZN(n934) );
  INV_X1 U553 ( .A(n933), .ZN(n648) );
  AOI22_X1 U554 ( .A1(data_in[2]), .A2(n821), .B1(n935), .B2(\mem[29][2] ), 
        .ZN(n933) );
  INV_X1 U555 ( .A(n932), .ZN(n647) );
  AOI22_X1 U556 ( .A1(data_in[3]), .A2(n821), .B1(n935), .B2(\mem[29][3] ), 
        .ZN(n932) );
  INV_X1 U557 ( .A(n931), .ZN(n646) );
  AOI22_X1 U558 ( .A1(data_in[4]), .A2(n821), .B1(n935), .B2(\mem[29][4] ), 
        .ZN(n931) );
  INV_X1 U559 ( .A(n930), .ZN(n645) );
  AOI22_X1 U560 ( .A1(data_in[5]), .A2(n821), .B1(n935), .B2(\mem[29][5] ), 
        .ZN(n930) );
  INV_X1 U561 ( .A(n929), .ZN(n644) );
  AOI22_X1 U562 ( .A1(data_in[6]), .A2(n821), .B1(n935), .B2(\mem[29][6] ), 
        .ZN(n929) );
  INV_X1 U563 ( .A(n928), .ZN(n643) );
  AOI22_X1 U564 ( .A1(data_in[7]), .A2(n821), .B1(n935), .B2(\mem[29][7] ), 
        .ZN(n928) );
  INV_X1 U565 ( .A(n927), .ZN(n642) );
  AOI22_X1 U566 ( .A1(data_in[0]), .A2(n820), .B1(n926), .B2(\mem[30][0] ), 
        .ZN(n927) );
  INV_X1 U567 ( .A(n925), .ZN(n641) );
  AOI22_X1 U568 ( .A1(data_in[1]), .A2(n820), .B1(n926), .B2(\mem[30][1] ), 
        .ZN(n925) );
  INV_X1 U569 ( .A(n924), .ZN(n640) );
  AOI22_X1 U570 ( .A1(data_in[2]), .A2(n820), .B1(n926), .B2(\mem[30][2] ), 
        .ZN(n924) );
  INV_X1 U571 ( .A(n923), .ZN(n639) );
  AOI22_X1 U572 ( .A1(data_in[3]), .A2(n820), .B1(n926), .B2(\mem[30][3] ), 
        .ZN(n923) );
  INV_X1 U573 ( .A(n922), .ZN(n638) );
  AOI22_X1 U574 ( .A1(data_in[4]), .A2(n820), .B1(n926), .B2(\mem[30][4] ), 
        .ZN(n922) );
  INV_X1 U575 ( .A(n921), .ZN(n637) );
  AOI22_X1 U576 ( .A1(data_in[5]), .A2(n820), .B1(n926), .B2(\mem[30][5] ), 
        .ZN(n921) );
  INV_X1 U577 ( .A(n920), .ZN(n636) );
  AOI22_X1 U578 ( .A1(data_in[6]), .A2(n820), .B1(n926), .B2(\mem[30][6] ), 
        .ZN(n920) );
  INV_X1 U579 ( .A(n919), .ZN(n635) );
  AOI22_X1 U580 ( .A1(data_in[7]), .A2(n820), .B1(n926), .B2(\mem[30][7] ), 
        .ZN(n919) );
  INV_X1 U581 ( .A(n918), .ZN(n634) );
  AOI22_X1 U582 ( .A1(data_in[0]), .A2(n819), .B1(n917), .B2(\mem[31][0] ), 
        .ZN(n918) );
  INV_X1 U583 ( .A(n916), .ZN(n633) );
  AOI22_X1 U584 ( .A1(data_in[1]), .A2(n819), .B1(n917), .B2(\mem[31][1] ), 
        .ZN(n916) );
  INV_X1 U585 ( .A(n915), .ZN(n632) );
  AOI22_X1 U586 ( .A1(data_in[2]), .A2(n819), .B1(n917), .B2(\mem[31][2] ), 
        .ZN(n915) );
  INV_X1 U587 ( .A(n914), .ZN(n631) );
  AOI22_X1 U588 ( .A1(data_in[3]), .A2(n819), .B1(n917), .B2(\mem[31][3] ), 
        .ZN(n914) );
  INV_X1 U589 ( .A(n913), .ZN(n630) );
  AOI22_X1 U590 ( .A1(data_in[4]), .A2(n819), .B1(n917), .B2(\mem[31][4] ), 
        .ZN(n913) );
  INV_X1 U591 ( .A(n912), .ZN(n629) );
  AOI22_X1 U592 ( .A1(data_in[5]), .A2(n819), .B1(n917), .B2(\mem[31][5] ), 
        .ZN(n912) );
  INV_X1 U593 ( .A(n911), .ZN(n628) );
  AOI22_X1 U594 ( .A1(data_in[6]), .A2(n819), .B1(n917), .B2(\mem[31][6] ), 
        .ZN(n911) );
  INV_X1 U595 ( .A(n910), .ZN(n627) );
  AOI22_X1 U596 ( .A1(data_in[7]), .A2(n819), .B1(n917), .B2(\mem[31][7] ), 
        .ZN(n910) );
  MUX2_X1 U597 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n611), .Z(n1) );
  MUX2_X1 U598 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n611), .Z(n2) );
  MUX2_X1 U599 ( .A(n2), .B(n1), .S(n608), .Z(n3) );
  MUX2_X1 U600 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n611), .Z(n4) );
  MUX2_X1 U601 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n611), .Z(n5) );
  MUX2_X1 U602 ( .A(n5), .B(n4), .S(n608), .Z(n6) );
  MUX2_X1 U603 ( .A(n6), .B(n3), .S(n606), .Z(n7) );
  MUX2_X1 U604 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n611), .Z(n8) );
  MUX2_X1 U605 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n611), .Z(n9) );
  MUX2_X1 U606 ( .A(n9), .B(n8), .S(n608), .Z(n10) );
  MUX2_X1 U607 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n611), .Z(n11) );
  MUX2_X1 U608 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n611), .Z(n12) );
  MUX2_X1 U609 ( .A(n12), .B(n11), .S(n608), .Z(n13) );
  MUX2_X1 U610 ( .A(n13), .B(n10), .S(N12), .Z(n14) );
  MUX2_X1 U611 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U612 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n614), .Z(n16) );
  MUX2_X1 U613 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n615), .Z(n17) );
  MUX2_X1 U614 ( .A(n17), .B(n16), .S(n608), .Z(n18) );
  MUX2_X1 U615 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(N10), .Z(n19) );
  MUX2_X1 U616 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n20) );
  MUX2_X1 U617 ( .A(n20), .B(n19), .S(n609), .Z(n21) );
  MUX2_X1 U618 ( .A(n21), .B(n18), .S(N12), .Z(n22) );
  MUX2_X1 U619 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n611), .Z(n23) );
  MUX2_X1 U620 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n616), .Z(n24) );
  MUX2_X1 U621 ( .A(n24), .B(n23), .S(n608), .Z(n25) );
  MUX2_X1 U622 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n26) );
  MUX2_X1 U623 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n27) );
  MUX2_X1 U624 ( .A(n27), .B(n26), .S(n610), .Z(n28) );
  MUX2_X1 U625 ( .A(n28), .B(n25), .S(n607), .Z(n29) );
  MUX2_X1 U626 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U627 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U628 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n612), .Z(n31) );
  MUX2_X1 U629 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n616), .Z(n32) );
  MUX2_X1 U630 ( .A(n32), .B(n31), .S(n608), .Z(n33) );
  MUX2_X1 U631 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n613), .Z(n34) );
  MUX2_X1 U632 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n616), .Z(n35) );
  MUX2_X1 U633 ( .A(n35), .B(n34), .S(n608), .Z(n36) );
  MUX2_X1 U634 ( .A(n36), .B(n33), .S(n607), .Z(n37) );
  MUX2_X1 U635 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n611), .Z(n38) );
  MUX2_X1 U636 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n614), .Z(n39) );
  MUX2_X1 U637 ( .A(n39), .B(n38), .S(n608), .Z(n40) );
  MUX2_X1 U638 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n615), .Z(n41) );
  MUX2_X1 U639 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n616), .Z(n42) );
  MUX2_X1 U640 ( .A(n42), .B(n41), .S(N11), .Z(n43) );
  MUX2_X1 U641 ( .A(n43), .B(n40), .S(N12), .Z(n44) );
  MUX2_X1 U642 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U643 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n611), .Z(n46) );
  MUX2_X1 U644 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n611), .Z(n47) );
  MUX2_X1 U645 ( .A(n47), .B(n46), .S(n608), .Z(n48) );
  MUX2_X1 U646 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n612), .Z(n49) );
  MUX2_X1 U647 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n614), .Z(n50) );
  MUX2_X1 U648 ( .A(n50), .B(n49), .S(n610), .Z(n51) );
  MUX2_X1 U649 ( .A(n51), .B(n48), .S(n606), .Z(n52) );
  MUX2_X1 U650 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n611), .Z(n53) );
  MUX2_X1 U651 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n615), .Z(n54) );
  MUX2_X1 U652 ( .A(n54), .B(n53), .S(n608), .Z(n55) );
  MUX2_X1 U653 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n612), .Z(n56) );
  MUX2_X1 U654 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n616), .Z(n57) );
  MUX2_X1 U655 ( .A(n57), .B(n56), .S(n608), .Z(n58) );
  MUX2_X1 U656 ( .A(n58), .B(n55), .S(n606), .Z(n59) );
  MUX2_X1 U657 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U658 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U659 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n612), .Z(n61) );
  MUX2_X1 U660 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n612), .Z(n62) );
  MUX2_X1 U661 ( .A(n62), .B(n61), .S(n609), .Z(n63) );
  MUX2_X1 U662 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n612), .Z(n64) );
  MUX2_X1 U663 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n612), .Z(n65) );
  MUX2_X1 U664 ( .A(n65), .B(n64), .S(n609), .Z(n66) );
  MUX2_X1 U665 ( .A(n66), .B(n63), .S(n606), .Z(n67) );
  MUX2_X1 U666 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n612), .Z(n68) );
  MUX2_X1 U667 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n612), .Z(n69) );
  MUX2_X1 U668 ( .A(n69), .B(n68), .S(n609), .Z(n70) );
  MUX2_X1 U669 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n612), .Z(n71) );
  MUX2_X1 U670 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n612), .Z(n72) );
  MUX2_X1 U671 ( .A(n72), .B(n71), .S(n609), .Z(n73) );
  MUX2_X1 U672 ( .A(n73), .B(n70), .S(n606), .Z(n74) );
  MUX2_X1 U673 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U674 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n612), .Z(n76) );
  MUX2_X1 U675 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n612), .Z(n77) );
  MUX2_X1 U676 ( .A(n77), .B(n76), .S(n609), .Z(n78) );
  MUX2_X1 U677 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n612), .Z(n79) );
  MUX2_X1 U678 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n612), .Z(n80) );
  MUX2_X1 U679 ( .A(n80), .B(n79), .S(n609), .Z(n81) );
  MUX2_X1 U680 ( .A(n81), .B(n78), .S(n606), .Z(n82) );
  MUX2_X1 U681 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n613), .Z(n83) );
  MUX2_X1 U682 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n613), .Z(n84) );
  MUX2_X1 U683 ( .A(n84), .B(n83), .S(n609), .Z(n85) );
  MUX2_X1 U684 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n613), .Z(n86) );
  MUX2_X1 U685 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n613), .Z(n87) );
  MUX2_X1 U686 ( .A(n87), .B(n86), .S(n609), .Z(n88) );
  MUX2_X1 U687 ( .A(n88), .B(n85), .S(n606), .Z(n89) );
  MUX2_X1 U688 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U689 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U690 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n613), .Z(n91) );
  MUX2_X1 U691 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n613), .Z(n92) );
  MUX2_X1 U692 ( .A(n92), .B(n91), .S(n609), .Z(n93) );
  MUX2_X1 U693 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n613), .Z(n94) );
  MUX2_X1 U694 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n613), .Z(n95) );
  MUX2_X1 U695 ( .A(n95), .B(n94), .S(n609), .Z(n96) );
  MUX2_X1 U696 ( .A(n96), .B(n93), .S(n606), .Z(n97) );
  MUX2_X1 U697 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n613), .Z(n98) );
  MUX2_X1 U698 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n613), .Z(n99) );
  MUX2_X1 U699 ( .A(n99), .B(n98), .S(n609), .Z(n100) );
  MUX2_X1 U700 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n613), .Z(n101) );
  MUX2_X1 U701 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n613), .Z(n102) );
  MUX2_X1 U702 ( .A(n102), .B(n101), .S(n609), .Z(n103) );
  MUX2_X1 U703 ( .A(n103), .B(n100), .S(n606), .Z(n104) );
  MUX2_X1 U704 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U705 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n616), .Z(n106) );
  MUX2_X1 U706 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n616), .Z(n107) );
  MUX2_X1 U707 ( .A(n107), .B(n106), .S(n610), .Z(n108) );
  MUX2_X1 U708 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n616), .Z(n109) );
  MUX2_X1 U709 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n611), .Z(n110) );
  MUX2_X1 U710 ( .A(n110), .B(n109), .S(n610), .Z(n111) );
  MUX2_X1 U711 ( .A(n111), .B(n108), .S(n606), .Z(n112) );
  MUX2_X1 U712 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n616), .Z(n113) );
  MUX2_X1 U713 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n612), .Z(n114) );
  MUX2_X1 U714 ( .A(n114), .B(n113), .S(n610), .Z(n115) );
  MUX2_X1 U715 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n615), .Z(n116) );
  MUX2_X1 U716 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n614), .Z(n117) );
  MUX2_X1 U717 ( .A(n117), .B(n116), .S(n610), .Z(n118) );
  MUX2_X1 U718 ( .A(n118), .B(n115), .S(n606), .Z(n119) );
  MUX2_X1 U719 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U720 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U721 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n616), .Z(n121) );
  MUX2_X1 U722 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n616), .Z(n122) );
  MUX2_X1 U723 ( .A(n122), .B(n121), .S(n610), .Z(n123) );
  MUX2_X1 U724 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n616), .Z(n124) );
  MUX2_X1 U725 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n616), .Z(n125) );
  MUX2_X1 U726 ( .A(n125), .B(n124), .S(n610), .Z(n126) );
  MUX2_X1 U727 ( .A(n126), .B(n123), .S(n606), .Z(n127) );
  MUX2_X1 U728 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n615), .Z(n128) );
  MUX2_X1 U729 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(N10), .Z(n129) );
  MUX2_X1 U730 ( .A(n129), .B(n128), .S(n610), .Z(n130) );
  MUX2_X1 U731 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n612), .Z(n131) );
  MUX2_X1 U732 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n616), .Z(n132) );
  MUX2_X1 U733 ( .A(n132), .B(n131), .S(n610), .Z(n133) );
  MUX2_X1 U734 ( .A(n133), .B(n130), .S(n606), .Z(n134) );
  MUX2_X1 U735 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U736 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n616), .Z(n136) );
  MUX2_X1 U737 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n616), .Z(n137) );
  MUX2_X1 U738 ( .A(n137), .B(n136), .S(n610), .Z(n138) );
  MUX2_X1 U739 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n611), .Z(n139) );
  MUX2_X1 U740 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n616), .Z(n140) );
  MUX2_X1 U741 ( .A(n140), .B(n139), .S(n610), .Z(n141) );
  MUX2_X1 U742 ( .A(n141), .B(n138), .S(n606), .Z(n142) );
  MUX2_X1 U743 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n611), .Z(n143) );
  MUX2_X1 U744 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n616), .Z(n144) );
  MUX2_X1 U745 ( .A(n144), .B(n143), .S(n610), .Z(n145) );
  MUX2_X1 U746 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n616), .Z(n146) );
  MUX2_X1 U747 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n616), .Z(n147) );
  MUX2_X1 U748 ( .A(n147), .B(n146), .S(n610), .Z(n148) );
  MUX2_X1 U749 ( .A(n148), .B(n145), .S(n606), .Z(n149) );
  MUX2_X1 U750 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U751 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U752 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n613), .Z(n151) );
  MUX2_X1 U753 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n613), .Z(n152) );
  MUX2_X1 U754 ( .A(n152), .B(n151), .S(n608), .Z(n153) );
  MUX2_X1 U755 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n613), .Z(n154) );
  MUX2_X1 U756 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n613), .Z(n155) );
  MUX2_X1 U757 ( .A(n155), .B(n154), .S(n608), .Z(n156) );
  MUX2_X1 U758 ( .A(n156), .B(n153), .S(n607), .Z(n157) );
  MUX2_X1 U759 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n613), .Z(n158) );
  MUX2_X1 U760 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n613), .Z(n159) );
  MUX2_X1 U761 ( .A(n159), .B(n158), .S(n610), .Z(n160) );
  MUX2_X1 U762 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n613), .Z(n161) );
  MUX2_X1 U763 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n611), .Z(n162) );
  MUX2_X1 U764 ( .A(n162), .B(n161), .S(n609), .Z(n163) );
  MUX2_X1 U765 ( .A(n163), .B(n160), .S(n607), .Z(n164) );
  MUX2_X1 U766 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U767 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n613), .Z(n166) );
  MUX2_X1 U768 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n613), .Z(n167) );
  MUX2_X1 U769 ( .A(n167), .B(n166), .S(n609), .Z(n168) );
  MUX2_X1 U770 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n613), .Z(n169) );
  MUX2_X1 U771 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n612), .Z(n170) );
  MUX2_X1 U772 ( .A(n170), .B(n169), .S(n610), .Z(n171) );
  MUX2_X1 U773 ( .A(n171), .B(n168), .S(n607), .Z(n172) );
  MUX2_X1 U774 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n614), .Z(n173) );
  MUX2_X1 U775 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n614), .Z(n174) );
  MUX2_X1 U776 ( .A(n174), .B(n173), .S(N11), .Z(n175) );
  MUX2_X1 U777 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n614), .Z(n176) );
  MUX2_X1 U778 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n614), .Z(n177) );
  MUX2_X1 U779 ( .A(n177), .B(n176), .S(n608), .Z(n178) );
  MUX2_X1 U780 ( .A(n178), .B(n175), .S(n607), .Z(n179) );
  MUX2_X1 U781 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U782 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U783 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n614), .Z(n181) );
  MUX2_X1 U784 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n614), .Z(n182) );
  MUX2_X1 U785 ( .A(n182), .B(n181), .S(n610), .Z(n183) );
  MUX2_X1 U786 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n614), .Z(n184) );
  MUX2_X1 U787 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n614), .Z(n185) );
  MUX2_X1 U788 ( .A(n185), .B(n184), .S(n610), .Z(n186) );
  MUX2_X1 U789 ( .A(n186), .B(n183), .S(n607), .Z(n187) );
  MUX2_X1 U790 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n614), .Z(n188) );
  MUX2_X1 U791 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n614), .Z(n189) );
  MUX2_X1 U792 ( .A(n189), .B(n188), .S(n608), .Z(n190) );
  MUX2_X1 U793 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n614), .Z(n191) );
  MUX2_X1 U794 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n614), .Z(n192) );
  MUX2_X1 U795 ( .A(n192), .B(n191), .S(n608), .Z(n193) );
  MUX2_X1 U796 ( .A(n193), .B(n190), .S(n607), .Z(n194) );
  MUX2_X1 U797 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U798 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n615), .Z(n196) );
  MUX2_X1 U799 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n615), .Z(n197) );
  MUX2_X1 U800 ( .A(n197), .B(n196), .S(n610), .Z(n198) );
  MUX2_X1 U801 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n615), .Z(n199) );
  MUX2_X1 U802 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n615), .Z(n200) );
  MUX2_X1 U803 ( .A(n200), .B(n199), .S(n610), .Z(n201) );
  MUX2_X1 U804 ( .A(n201), .B(n198), .S(n607), .Z(n202) );
  MUX2_X1 U805 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n615), .Z(n203) );
  MUX2_X1 U806 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n615), .Z(n204) );
  MUX2_X1 U807 ( .A(n204), .B(n203), .S(N11), .Z(n205) );
  MUX2_X1 U808 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n615), .Z(n206) );
  MUX2_X1 U809 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n615), .Z(n207) );
  MUX2_X1 U810 ( .A(n207), .B(n206), .S(n609), .Z(n208) );
  MUX2_X1 U811 ( .A(n208), .B(n205), .S(n607), .Z(n209) );
  MUX2_X1 U812 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U813 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U814 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n615), .Z(n211) );
  MUX2_X1 U815 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n615), .Z(n212) );
  MUX2_X1 U816 ( .A(n212), .B(n211), .S(n609), .Z(n213) );
  MUX2_X1 U817 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n615), .Z(n214) );
  MUX2_X1 U818 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n615), .Z(n215) );
  MUX2_X1 U819 ( .A(n215), .B(n214), .S(N11), .Z(n216) );
  MUX2_X1 U820 ( .A(n216), .B(n213), .S(n607), .Z(n217) );
  MUX2_X1 U821 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n615), .Z(n218) );
  MUX2_X1 U822 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n611), .Z(n219) );
  MUX2_X1 U823 ( .A(n219), .B(n218), .S(n608), .Z(n220) );
  MUX2_X1 U824 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n615), .Z(n221) );
  MUX2_X1 U825 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n612), .Z(n222) );
  MUX2_X1 U826 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U827 ( .A(n223), .B(n220), .S(n607), .Z(n224) );
  MUX2_X1 U828 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U829 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n614), .Z(n226) );
  MUX2_X1 U830 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n611), .Z(n227) );
  MUX2_X1 U831 ( .A(n227), .B(n226), .S(n609), .Z(n228) );
  MUX2_X1 U832 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n614), .Z(n229) );
  MUX2_X1 U833 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n611), .Z(n595) );
  MUX2_X1 U834 ( .A(n595), .B(n229), .S(n609), .Z(n596) );
  MUX2_X1 U835 ( .A(n596), .B(n228), .S(n607), .Z(n597) );
  MUX2_X1 U836 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n615), .Z(n598) );
  MUX2_X1 U837 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n612), .Z(n599) );
  MUX2_X1 U838 ( .A(n599), .B(n598), .S(n609), .Z(n600) );
  MUX2_X1 U839 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n614), .Z(n601) );
  MUX2_X1 U840 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n614), .Z(n602) );
  MUX2_X1 U841 ( .A(n602), .B(n601), .S(n610), .Z(n603) );
  MUX2_X1 U842 ( .A(n603), .B(n600), .S(n607), .Z(n604) );
  MUX2_X1 U843 ( .A(n604), .B(n597), .S(N13), .Z(n605) );
  MUX2_X1 U844 ( .A(n605), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U845 ( .A(N11), .Z(n608) );
  INV_X1 U846 ( .A(N10), .ZN(n617) );
  INV_X1 U847 ( .A(N11), .ZN(n618) );
  INV_X1 U848 ( .A(data_in[0]), .ZN(n619) );
  INV_X1 U849 ( .A(data_in[1]), .ZN(n620) );
  INV_X1 U850 ( .A(data_in[2]), .ZN(n621) );
  INV_X1 U851 ( .A(data_in[3]), .ZN(n622) );
  INV_X1 U852 ( .A(data_in[4]), .ZN(n623) );
  INV_X1 U853 ( .A(data_in[5]), .ZN(n624) );
  INV_X1 U854 ( .A(data_in[6]), .ZN(n625) );
  INV_X1 U855 ( .A(data_in[7]), .ZN(n626) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_17 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n628), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n629), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n630), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n631), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n632), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n633), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n634), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n635), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n636), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n637), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n638), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n639), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n640), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n641), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n642), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n643), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n644), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n645), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n646), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n647), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n648), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n649), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n650), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n651), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n652), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n653), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n654), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n655), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n656), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n657), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n658), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n659), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n660), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n661), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n662), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n663), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n664), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n665), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n666), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n667), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n668), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n669), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n670), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n671), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n672), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n673), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n674), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n675), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n676), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n677), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n678), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n679), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n680), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n681), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n682), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n683), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n684), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n685), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n686), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n687), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n688), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n689), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n690), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n691), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n692), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n693), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n694), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n695), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n696), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n697), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n698), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n699), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n700), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n701), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n702), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n703), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n704), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n705), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n706), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n707), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n708), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n709), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n710), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n711), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n712), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n713), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n714), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n715), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n716), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n717), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n718), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n719), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n720), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n721), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n722), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n723), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n724), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n725), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n726), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n727), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n728), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n729), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n730), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n731), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n732), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n733), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n734), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n735), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n736), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n737), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n738), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n739), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n740), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n741), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n742), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n743), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n744), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n745), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n746), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n747), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n748), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n749), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n750), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n751), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n752), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n753), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n754), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n755), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n756), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n757), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n758), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n759), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n760), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n761), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n762), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n763), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n764), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n765), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n766), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n767), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n768), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n769), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n770), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n771), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n772), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n773), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n774), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n775), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n776), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n777), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n778), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n779), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n780), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n781), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n782), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n783), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n784), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n785), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n786), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n787), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n788), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n789), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n790), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n791), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n792), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n793), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n794), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n795), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n796), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n797), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n798), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n799), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n800), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n801), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n802), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n803), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n804), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n805), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n806), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n807), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n808), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n809), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n810), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n811), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n812), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n813), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n814), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n815), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n816), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n817), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n818), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n819), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n847), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n848), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n849), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n850), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n851), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n852), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n853), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n854), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n855), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n856), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n857), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n858), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n859), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n860), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n861), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n862), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n863), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n864), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n865), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n866), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n867), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n868), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n869), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n870), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n871), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n872), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n873), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n874), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n875), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n876), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n877), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n878), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n879), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n880), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n881), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n882), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n883), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n884), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n885), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n886), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n887), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n888), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n889), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n890), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n891), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n892), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n893), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n894), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n895), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n896), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n897), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n898), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n899), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n900), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n901), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n902), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n903), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n904), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n905), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n906), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n907), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n908), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n909), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n910), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  BUF_X1 U3 ( .A(n617), .Z(n614) );
  BUF_X1 U4 ( .A(n617), .Z(n615) );
  BUF_X1 U5 ( .A(n617), .Z(n616) );
  BUF_X1 U6 ( .A(n617), .Z(n612) );
  BUF_X1 U7 ( .A(n617), .Z(n613) );
  BUF_X1 U8 ( .A(N11), .Z(n609) );
  BUF_X1 U9 ( .A(N11), .Z(n610) );
  BUF_X1 U10 ( .A(N10), .Z(n617) );
  NOR3_X1 U11 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1202) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(n618), .ZN(n1191) );
  NOR3_X1 U13 ( .A1(N10), .A2(N12), .A3(n619), .ZN(n1181) );
  NOR3_X1 U14 ( .A1(n618), .A2(N12), .A3(n619), .ZN(n1171) );
  INV_X1 U15 ( .A(n1128), .ZN(n843) );
  INV_X1 U16 ( .A(n1118), .ZN(n842) );
  INV_X1 U17 ( .A(n1109), .ZN(n841) );
  INV_X1 U18 ( .A(n1100), .ZN(n840) );
  INV_X1 U19 ( .A(n1055), .ZN(n835) );
  INV_X1 U20 ( .A(n1045), .ZN(n834) );
  INV_X1 U21 ( .A(n1036), .ZN(n833) );
  INV_X1 U22 ( .A(n1027), .ZN(n832) );
  INV_X1 U23 ( .A(n982), .ZN(n827) );
  INV_X1 U24 ( .A(n972), .ZN(n826) );
  INV_X1 U25 ( .A(n963), .ZN(n825) );
  INV_X1 U26 ( .A(n954), .ZN(n824) );
  INV_X1 U27 ( .A(n945), .ZN(n823) );
  INV_X1 U28 ( .A(n936), .ZN(n822) );
  INV_X1 U29 ( .A(n927), .ZN(n821) );
  INV_X1 U30 ( .A(n918), .ZN(n820) );
  INV_X1 U31 ( .A(n1091), .ZN(n839) );
  INV_X1 U32 ( .A(n1082), .ZN(n838) );
  INV_X1 U33 ( .A(n1073), .ZN(n837) );
  INV_X1 U34 ( .A(n1064), .ZN(n836) );
  INV_X1 U35 ( .A(n1018), .ZN(n831) );
  INV_X1 U36 ( .A(n1009), .ZN(n830) );
  INV_X1 U37 ( .A(n1000), .ZN(n829) );
  INV_X1 U38 ( .A(n991), .ZN(n828) );
  BUF_X1 U39 ( .A(N12), .Z(n606) );
  BUF_X1 U40 ( .A(N12), .Z(n607) );
  INV_X1 U41 ( .A(N13), .ZN(n845) );
  AND3_X1 U42 ( .A1(n618), .A2(n619), .A3(N12), .ZN(n1161) );
  AND3_X1 U43 ( .A1(N10), .A2(n619), .A3(N12), .ZN(n1151) );
  AND3_X1 U44 ( .A1(N11), .A2(n618), .A3(N12), .ZN(n1141) );
  AND3_X1 U45 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1131) );
  INV_X1 U46 ( .A(N14), .ZN(n846) );
  NAND2_X1 U47 ( .A1(n1191), .A2(n1201), .ZN(n1200) );
  NAND2_X1 U48 ( .A1(n1181), .A2(n1201), .ZN(n1190) );
  NAND2_X1 U49 ( .A1(n1171), .A2(n1201), .ZN(n1180) );
  NAND2_X1 U50 ( .A1(n1161), .A2(n1201), .ZN(n1170) );
  NAND2_X1 U51 ( .A1(n1151), .A2(n1201), .ZN(n1160) );
  NAND2_X1 U52 ( .A1(n1141), .A2(n1201), .ZN(n1150) );
  NAND2_X1 U53 ( .A1(n1131), .A2(n1201), .ZN(n1140) );
  NAND2_X1 U54 ( .A1(n1202), .A2(n1201), .ZN(n1211) );
  NAND2_X1 U55 ( .A1(n1120), .A2(n1202), .ZN(n1128) );
  NAND2_X1 U56 ( .A1(n1120), .A2(n1191), .ZN(n1118) );
  NAND2_X1 U57 ( .A1(n1120), .A2(n1181), .ZN(n1109) );
  NAND2_X1 U58 ( .A1(n1120), .A2(n1171), .ZN(n1100) );
  NAND2_X1 U59 ( .A1(n1047), .A2(n1202), .ZN(n1055) );
  NAND2_X1 U60 ( .A1(n1047), .A2(n1191), .ZN(n1045) );
  NAND2_X1 U61 ( .A1(n1047), .A2(n1181), .ZN(n1036) );
  NAND2_X1 U62 ( .A1(n1047), .A2(n1171), .ZN(n1027) );
  NAND2_X1 U63 ( .A1(n974), .A2(n1202), .ZN(n982) );
  NAND2_X1 U64 ( .A1(n974), .A2(n1191), .ZN(n972) );
  NAND2_X1 U65 ( .A1(n974), .A2(n1181), .ZN(n963) );
  NAND2_X1 U66 ( .A1(n974), .A2(n1171), .ZN(n954) );
  NAND2_X1 U67 ( .A1(n1120), .A2(n1161), .ZN(n1091) );
  NAND2_X1 U68 ( .A1(n1120), .A2(n1151), .ZN(n1082) );
  NAND2_X1 U69 ( .A1(n1120), .A2(n1141), .ZN(n1073) );
  NAND2_X1 U70 ( .A1(n1120), .A2(n1131), .ZN(n1064) );
  NAND2_X1 U71 ( .A1(n1047), .A2(n1161), .ZN(n1018) );
  NAND2_X1 U72 ( .A1(n1047), .A2(n1151), .ZN(n1009) );
  NAND2_X1 U73 ( .A1(n1047), .A2(n1141), .ZN(n1000) );
  NAND2_X1 U74 ( .A1(n1047), .A2(n1131), .ZN(n991) );
  NAND2_X1 U75 ( .A1(n974), .A2(n1161), .ZN(n945) );
  NAND2_X1 U76 ( .A1(n974), .A2(n1151), .ZN(n936) );
  NAND2_X1 U77 ( .A1(n974), .A2(n1141), .ZN(n927) );
  NAND2_X1 U78 ( .A1(n974), .A2(n1131), .ZN(n918) );
  AND3_X1 U79 ( .A1(n845), .A2(n846), .A3(n1130), .ZN(n1201) );
  AND3_X1 U80 ( .A1(N13), .A2(n1130), .A3(N14), .ZN(n974) );
  AND3_X1 U81 ( .A1(n1130), .A2(n846), .A3(N13), .ZN(n1120) );
  AND3_X1 U82 ( .A1(n1130), .A2(n845), .A3(N14), .ZN(n1047) );
  NOR2_X1 U83 ( .A1(n844), .A2(addr[5]), .ZN(n1130) );
  INV_X1 U84 ( .A(wr_en), .ZN(n844) );
  OAI21_X1 U85 ( .B1(n620), .B2(n1170), .A(n1169), .ZN(n878) );
  NAND2_X1 U86 ( .A1(\mem[4][0] ), .A2(n1170), .ZN(n1169) );
  OAI21_X1 U87 ( .B1(n621), .B2(n1170), .A(n1168), .ZN(n877) );
  NAND2_X1 U88 ( .A1(\mem[4][1] ), .A2(n1170), .ZN(n1168) );
  OAI21_X1 U89 ( .B1(n622), .B2(n1170), .A(n1167), .ZN(n876) );
  NAND2_X1 U90 ( .A1(\mem[4][2] ), .A2(n1170), .ZN(n1167) );
  OAI21_X1 U91 ( .B1(n623), .B2(n1170), .A(n1166), .ZN(n875) );
  NAND2_X1 U92 ( .A1(\mem[4][3] ), .A2(n1170), .ZN(n1166) );
  OAI21_X1 U93 ( .B1(n624), .B2(n1170), .A(n1165), .ZN(n874) );
  NAND2_X1 U94 ( .A1(\mem[4][4] ), .A2(n1170), .ZN(n1165) );
  OAI21_X1 U95 ( .B1(n625), .B2(n1170), .A(n1164), .ZN(n873) );
  NAND2_X1 U96 ( .A1(\mem[4][5] ), .A2(n1170), .ZN(n1164) );
  OAI21_X1 U97 ( .B1(n626), .B2(n1170), .A(n1163), .ZN(n872) );
  NAND2_X1 U98 ( .A1(\mem[4][6] ), .A2(n1170), .ZN(n1163) );
  OAI21_X1 U99 ( .B1(n627), .B2(n1170), .A(n1162), .ZN(n871) );
  NAND2_X1 U100 ( .A1(\mem[4][7] ), .A2(n1170), .ZN(n1162) );
  OAI21_X1 U101 ( .B1(n620), .B2(n1150), .A(n1149), .ZN(n862) );
  NAND2_X1 U102 ( .A1(\mem[6][0] ), .A2(n1150), .ZN(n1149) );
  OAI21_X1 U103 ( .B1(n621), .B2(n1150), .A(n1148), .ZN(n861) );
  NAND2_X1 U104 ( .A1(\mem[6][1] ), .A2(n1150), .ZN(n1148) );
  OAI21_X1 U105 ( .B1(n622), .B2(n1150), .A(n1147), .ZN(n860) );
  NAND2_X1 U106 ( .A1(\mem[6][2] ), .A2(n1150), .ZN(n1147) );
  OAI21_X1 U107 ( .B1(n623), .B2(n1150), .A(n1146), .ZN(n859) );
  NAND2_X1 U108 ( .A1(\mem[6][3] ), .A2(n1150), .ZN(n1146) );
  OAI21_X1 U109 ( .B1(n624), .B2(n1150), .A(n1145), .ZN(n858) );
  NAND2_X1 U110 ( .A1(\mem[6][4] ), .A2(n1150), .ZN(n1145) );
  OAI21_X1 U111 ( .B1(n625), .B2(n1150), .A(n1144), .ZN(n857) );
  NAND2_X1 U112 ( .A1(\mem[6][5] ), .A2(n1150), .ZN(n1144) );
  OAI21_X1 U113 ( .B1(n626), .B2(n1150), .A(n1143), .ZN(n856) );
  NAND2_X1 U114 ( .A1(\mem[6][6] ), .A2(n1150), .ZN(n1143) );
  OAI21_X1 U115 ( .B1(n627), .B2(n1150), .A(n1142), .ZN(n855) );
  NAND2_X1 U116 ( .A1(\mem[6][7] ), .A2(n1150), .ZN(n1142) );
  OAI21_X1 U117 ( .B1(n620), .B2(n1140), .A(n1139), .ZN(n854) );
  NAND2_X1 U118 ( .A1(\mem[7][0] ), .A2(n1140), .ZN(n1139) );
  OAI21_X1 U119 ( .B1(n621), .B2(n1140), .A(n1138), .ZN(n853) );
  NAND2_X1 U120 ( .A1(\mem[7][1] ), .A2(n1140), .ZN(n1138) );
  OAI21_X1 U121 ( .B1(n622), .B2(n1140), .A(n1137), .ZN(n852) );
  NAND2_X1 U122 ( .A1(\mem[7][2] ), .A2(n1140), .ZN(n1137) );
  OAI21_X1 U123 ( .B1(n623), .B2(n1140), .A(n1136), .ZN(n851) );
  NAND2_X1 U124 ( .A1(\mem[7][3] ), .A2(n1140), .ZN(n1136) );
  OAI21_X1 U125 ( .B1(n624), .B2(n1140), .A(n1135), .ZN(n850) );
  NAND2_X1 U126 ( .A1(\mem[7][4] ), .A2(n1140), .ZN(n1135) );
  OAI21_X1 U127 ( .B1(n625), .B2(n1140), .A(n1134), .ZN(n849) );
  NAND2_X1 U128 ( .A1(\mem[7][5] ), .A2(n1140), .ZN(n1134) );
  OAI21_X1 U129 ( .B1(n626), .B2(n1140), .A(n1133), .ZN(n848) );
  NAND2_X1 U130 ( .A1(\mem[7][6] ), .A2(n1140), .ZN(n1133) );
  OAI21_X1 U131 ( .B1(n627), .B2(n1140), .A(n1132), .ZN(n847) );
  NAND2_X1 U132 ( .A1(\mem[7][7] ), .A2(n1140), .ZN(n1132) );
  OAI21_X1 U133 ( .B1(n620), .B2(n1200), .A(n1199), .ZN(n902) );
  NAND2_X1 U134 ( .A1(\mem[1][0] ), .A2(n1200), .ZN(n1199) );
  OAI21_X1 U135 ( .B1(n621), .B2(n1200), .A(n1198), .ZN(n901) );
  NAND2_X1 U136 ( .A1(\mem[1][1] ), .A2(n1200), .ZN(n1198) );
  OAI21_X1 U137 ( .B1(n622), .B2(n1200), .A(n1197), .ZN(n900) );
  NAND2_X1 U138 ( .A1(\mem[1][2] ), .A2(n1200), .ZN(n1197) );
  OAI21_X1 U139 ( .B1(n623), .B2(n1200), .A(n1196), .ZN(n899) );
  NAND2_X1 U140 ( .A1(\mem[1][3] ), .A2(n1200), .ZN(n1196) );
  OAI21_X1 U141 ( .B1(n624), .B2(n1200), .A(n1195), .ZN(n898) );
  NAND2_X1 U142 ( .A1(\mem[1][4] ), .A2(n1200), .ZN(n1195) );
  OAI21_X1 U143 ( .B1(n625), .B2(n1200), .A(n1194), .ZN(n897) );
  NAND2_X1 U144 ( .A1(\mem[1][5] ), .A2(n1200), .ZN(n1194) );
  OAI21_X1 U145 ( .B1(n626), .B2(n1200), .A(n1193), .ZN(n896) );
  NAND2_X1 U146 ( .A1(\mem[1][6] ), .A2(n1200), .ZN(n1193) );
  OAI21_X1 U147 ( .B1(n627), .B2(n1200), .A(n1192), .ZN(n895) );
  NAND2_X1 U148 ( .A1(\mem[1][7] ), .A2(n1200), .ZN(n1192) );
  OAI21_X1 U149 ( .B1(n620), .B2(n1190), .A(n1189), .ZN(n894) );
  NAND2_X1 U150 ( .A1(\mem[2][0] ), .A2(n1190), .ZN(n1189) );
  OAI21_X1 U151 ( .B1(n621), .B2(n1190), .A(n1188), .ZN(n893) );
  NAND2_X1 U152 ( .A1(\mem[2][1] ), .A2(n1190), .ZN(n1188) );
  OAI21_X1 U153 ( .B1(n622), .B2(n1190), .A(n1187), .ZN(n892) );
  NAND2_X1 U154 ( .A1(\mem[2][2] ), .A2(n1190), .ZN(n1187) );
  OAI21_X1 U155 ( .B1(n623), .B2(n1190), .A(n1186), .ZN(n891) );
  NAND2_X1 U156 ( .A1(\mem[2][3] ), .A2(n1190), .ZN(n1186) );
  OAI21_X1 U157 ( .B1(n624), .B2(n1190), .A(n1185), .ZN(n890) );
  NAND2_X1 U158 ( .A1(\mem[2][4] ), .A2(n1190), .ZN(n1185) );
  OAI21_X1 U159 ( .B1(n625), .B2(n1190), .A(n1184), .ZN(n889) );
  NAND2_X1 U160 ( .A1(\mem[2][5] ), .A2(n1190), .ZN(n1184) );
  OAI21_X1 U161 ( .B1(n626), .B2(n1190), .A(n1183), .ZN(n888) );
  NAND2_X1 U162 ( .A1(\mem[2][6] ), .A2(n1190), .ZN(n1183) );
  OAI21_X1 U163 ( .B1(n627), .B2(n1190), .A(n1182), .ZN(n887) );
  NAND2_X1 U164 ( .A1(\mem[2][7] ), .A2(n1190), .ZN(n1182) );
  OAI21_X1 U165 ( .B1(n620), .B2(n1180), .A(n1179), .ZN(n886) );
  NAND2_X1 U166 ( .A1(\mem[3][0] ), .A2(n1180), .ZN(n1179) );
  OAI21_X1 U167 ( .B1(n621), .B2(n1180), .A(n1178), .ZN(n885) );
  NAND2_X1 U168 ( .A1(\mem[3][1] ), .A2(n1180), .ZN(n1178) );
  OAI21_X1 U169 ( .B1(n622), .B2(n1180), .A(n1177), .ZN(n884) );
  NAND2_X1 U170 ( .A1(\mem[3][2] ), .A2(n1180), .ZN(n1177) );
  OAI21_X1 U171 ( .B1(n623), .B2(n1180), .A(n1176), .ZN(n883) );
  NAND2_X1 U172 ( .A1(\mem[3][3] ), .A2(n1180), .ZN(n1176) );
  OAI21_X1 U173 ( .B1(n624), .B2(n1180), .A(n1175), .ZN(n882) );
  NAND2_X1 U174 ( .A1(\mem[3][4] ), .A2(n1180), .ZN(n1175) );
  OAI21_X1 U175 ( .B1(n625), .B2(n1180), .A(n1174), .ZN(n881) );
  NAND2_X1 U176 ( .A1(\mem[3][5] ), .A2(n1180), .ZN(n1174) );
  OAI21_X1 U177 ( .B1(n626), .B2(n1180), .A(n1173), .ZN(n880) );
  NAND2_X1 U178 ( .A1(\mem[3][6] ), .A2(n1180), .ZN(n1173) );
  OAI21_X1 U179 ( .B1(n627), .B2(n1180), .A(n1172), .ZN(n879) );
  NAND2_X1 U180 ( .A1(\mem[3][7] ), .A2(n1180), .ZN(n1172) );
  OAI21_X1 U181 ( .B1(n620), .B2(n1160), .A(n1159), .ZN(n870) );
  NAND2_X1 U182 ( .A1(\mem[5][0] ), .A2(n1160), .ZN(n1159) );
  OAI21_X1 U183 ( .B1(n621), .B2(n1160), .A(n1158), .ZN(n869) );
  NAND2_X1 U184 ( .A1(\mem[5][1] ), .A2(n1160), .ZN(n1158) );
  OAI21_X1 U185 ( .B1(n622), .B2(n1160), .A(n1157), .ZN(n868) );
  NAND2_X1 U186 ( .A1(\mem[5][2] ), .A2(n1160), .ZN(n1157) );
  OAI21_X1 U187 ( .B1(n623), .B2(n1160), .A(n1156), .ZN(n867) );
  NAND2_X1 U188 ( .A1(\mem[5][3] ), .A2(n1160), .ZN(n1156) );
  OAI21_X1 U189 ( .B1(n624), .B2(n1160), .A(n1155), .ZN(n866) );
  NAND2_X1 U190 ( .A1(\mem[5][4] ), .A2(n1160), .ZN(n1155) );
  OAI21_X1 U191 ( .B1(n625), .B2(n1160), .A(n1154), .ZN(n865) );
  NAND2_X1 U192 ( .A1(\mem[5][5] ), .A2(n1160), .ZN(n1154) );
  OAI21_X1 U193 ( .B1(n626), .B2(n1160), .A(n1153), .ZN(n864) );
  NAND2_X1 U194 ( .A1(\mem[5][6] ), .A2(n1160), .ZN(n1153) );
  OAI21_X1 U195 ( .B1(n627), .B2(n1160), .A(n1152), .ZN(n863) );
  NAND2_X1 U196 ( .A1(\mem[5][7] ), .A2(n1160), .ZN(n1152) );
  OAI21_X1 U197 ( .B1(n1211), .B2(n620), .A(n1210), .ZN(n910) );
  NAND2_X1 U198 ( .A1(\mem[0][0] ), .A2(n1211), .ZN(n1210) );
  OAI21_X1 U199 ( .B1(n1211), .B2(n621), .A(n1209), .ZN(n909) );
  NAND2_X1 U200 ( .A1(\mem[0][1] ), .A2(n1211), .ZN(n1209) );
  OAI21_X1 U201 ( .B1(n1211), .B2(n622), .A(n1208), .ZN(n908) );
  NAND2_X1 U202 ( .A1(\mem[0][2] ), .A2(n1211), .ZN(n1208) );
  OAI21_X1 U203 ( .B1(n1211), .B2(n623), .A(n1207), .ZN(n907) );
  NAND2_X1 U204 ( .A1(\mem[0][3] ), .A2(n1211), .ZN(n1207) );
  OAI21_X1 U205 ( .B1(n1211), .B2(n624), .A(n1206), .ZN(n906) );
  NAND2_X1 U206 ( .A1(\mem[0][4] ), .A2(n1211), .ZN(n1206) );
  OAI21_X1 U207 ( .B1(n1211), .B2(n625), .A(n1205), .ZN(n905) );
  NAND2_X1 U208 ( .A1(\mem[0][5] ), .A2(n1211), .ZN(n1205) );
  OAI21_X1 U209 ( .B1(n1211), .B2(n626), .A(n1204), .ZN(n904) );
  NAND2_X1 U210 ( .A1(\mem[0][6] ), .A2(n1211), .ZN(n1204) );
  OAI21_X1 U211 ( .B1(n1211), .B2(n627), .A(n1203), .ZN(n903) );
  NAND2_X1 U212 ( .A1(\mem[0][7] ), .A2(n1211), .ZN(n1203) );
  INV_X1 U213 ( .A(n1129), .ZN(n819) );
  AOI22_X1 U214 ( .A1(data_in[0]), .A2(n843), .B1(n1128), .B2(\mem[8][0] ), 
        .ZN(n1129) );
  INV_X1 U215 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U216 ( .A1(data_in[1]), .A2(n843), .B1(n1128), .B2(\mem[8][1] ), 
        .ZN(n1127) );
  INV_X1 U217 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U218 ( .A1(data_in[2]), .A2(n843), .B1(n1128), .B2(\mem[8][2] ), 
        .ZN(n1126) );
  INV_X1 U219 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U220 ( .A1(data_in[3]), .A2(n843), .B1(n1128), .B2(\mem[8][3] ), 
        .ZN(n1125) );
  INV_X1 U221 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U222 ( .A1(data_in[4]), .A2(n843), .B1(n1128), .B2(\mem[8][4] ), 
        .ZN(n1124) );
  INV_X1 U223 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U224 ( .A1(data_in[5]), .A2(n843), .B1(n1128), .B2(\mem[8][5] ), 
        .ZN(n1123) );
  INV_X1 U225 ( .A(n1122), .ZN(n813) );
  AOI22_X1 U226 ( .A1(data_in[6]), .A2(n843), .B1(n1128), .B2(\mem[8][6] ), 
        .ZN(n1122) );
  INV_X1 U227 ( .A(n1121), .ZN(n812) );
  AOI22_X1 U228 ( .A1(data_in[7]), .A2(n843), .B1(n1128), .B2(\mem[8][7] ), 
        .ZN(n1121) );
  INV_X1 U229 ( .A(n1119), .ZN(n811) );
  AOI22_X1 U230 ( .A1(data_in[0]), .A2(n842), .B1(n1118), .B2(\mem[9][0] ), 
        .ZN(n1119) );
  INV_X1 U231 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U232 ( .A1(data_in[1]), .A2(n842), .B1(n1118), .B2(\mem[9][1] ), 
        .ZN(n1117) );
  INV_X1 U233 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U234 ( .A1(data_in[2]), .A2(n842), .B1(n1118), .B2(\mem[9][2] ), 
        .ZN(n1116) );
  INV_X1 U235 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U236 ( .A1(data_in[3]), .A2(n842), .B1(n1118), .B2(\mem[9][3] ), 
        .ZN(n1115) );
  INV_X1 U237 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U238 ( .A1(data_in[4]), .A2(n842), .B1(n1118), .B2(\mem[9][4] ), 
        .ZN(n1114) );
  INV_X1 U239 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U240 ( .A1(data_in[5]), .A2(n842), .B1(n1118), .B2(\mem[9][5] ), 
        .ZN(n1113) );
  INV_X1 U241 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U242 ( .A1(data_in[6]), .A2(n842), .B1(n1118), .B2(\mem[9][6] ), 
        .ZN(n1112) );
  INV_X1 U243 ( .A(n1111), .ZN(n804) );
  AOI22_X1 U244 ( .A1(data_in[7]), .A2(n842), .B1(n1118), .B2(\mem[9][7] ), 
        .ZN(n1111) );
  INV_X1 U245 ( .A(n1110), .ZN(n803) );
  AOI22_X1 U246 ( .A1(data_in[0]), .A2(n841), .B1(n1109), .B2(\mem[10][0] ), 
        .ZN(n1110) );
  INV_X1 U247 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U248 ( .A1(data_in[1]), .A2(n841), .B1(n1109), .B2(\mem[10][1] ), 
        .ZN(n1108) );
  INV_X1 U249 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U250 ( .A1(data_in[2]), .A2(n841), .B1(n1109), .B2(\mem[10][2] ), 
        .ZN(n1107) );
  INV_X1 U251 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U252 ( .A1(data_in[3]), .A2(n841), .B1(n1109), .B2(\mem[10][3] ), 
        .ZN(n1106) );
  INV_X1 U253 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U254 ( .A1(data_in[4]), .A2(n841), .B1(n1109), .B2(\mem[10][4] ), 
        .ZN(n1105) );
  INV_X1 U255 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U256 ( .A1(data_in[5]), .A2(n841), .B1(n1109), .B2(\mem[10][5] ), 
        .ZN(n1104) );
  INV_X1 U257 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U258 ( .A1(data_in[6]), .A2(n841), .B1(n1109), .B2(\mem[10][6] ), 
        .ZN(n1103) );
  INV_X1 U259 ( .A(n1102), .ZN(n796) );
  AOI22_X1 U260 ( .A1(data_in[7]), .A2(n841), .B1(n1109), .B2(\mem[10][7] ), 
        .ZN(n1102) );
  INV_X1 U261 ( .A(n1101), .ZN(n795) );
  AOI22_X1 U262 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[11][0] ), 
        .ZN(n1101) );
  INV_X1 U263 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U264 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[11][1] ), 
        .ZN(n1099) );
  INV_X1 U265 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U266 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[11][2] ), 
        .ZN(n1098) );
  INV_X1 U267 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U268 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[11][3] ), 
        .ZN(n1097) );
  INV_X1 U269 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U270 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[11][4] ), 
        .ZN(n1096) );
  INV_X1 U271 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U272 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[11][5] ), 
        .ZN(n1095) );
  INV_X1 U273 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U274 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[11][6] ), 
        .ZN(n1094) );
  INV_X1 U275 ( .A(n1093), .ZN(n788) );
  AOI22_X1 U276 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[11][7] ), 
        .ZN(n1093) );
  INV_X1 U277 ( .A(n1092), .ZN(n787) );
  AOI22_X1 U278 ( .A1(data_in[0]), .A2(n839), .B1(n1091), .B2(\mem[12][0] ), 
        .ZN(n1092) );
  INV_X1 U279 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U280 ( .A1(data_in[1]), .A2(n839), .B1(n1091), .B2(\mem[12][1] ), 
        .ZN(n1090) );
  INV_X1 U281 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U282 ( .A1(data_in[2]), .A2(n839), .B1(n1091), .B2(\mem[12][2] ), 
        .ZN(n1089) );
  INV_X1 U283 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U284 ( .A1(data_in[3]), .A2(n839), .B1(n1091), .B2(\mem[12][3] ), 
        .ZN(n1088) );
  INV_X1 U285 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U286 ( .A1(data_in[4]), .A2(n839), .B1(n1091), .B2(\mem[12][4] ), 
        .ZN(n1087) );
  INV_X1 U287 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U288 ( .A1(data_in[5]), .A2(n839), .B1(n1091), .B2(\mem[12][5] ), 
        .ZN(n1086) );
  INV_X1 U289 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U290 ( .A1(data_in[6]), .A2(n839), .B1(n1091), .B2(\mem[12][6] ), 
        .ZN(n1085) );
  INV_X1 U291 ( .A(n1084), .ZN(n780) );
  AOI22_X1 U292 ( .A1(data_in[7]), .A2(n839), .B1(n1091), .B2(\mem[12][7] ), 
        .ZN(n1084) );
  INV_X1 U293 ( .A(n1083), .ZN(n779) );
  AOI22_X1 U294 ( .A1(data_in[0]), .A2(n838), .B1(n1082), .B2(\mem[13][0] ), 
        .ZN(n1083) );
  INV_X1 U295 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U296 ( .A1(data_in[1]), .A2(n838), .B1(n1082), .B2(\mem[13][1] ), 
        .ZN(n1081) );
  INV_X1 U297 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U298 ( .A1(data_in[2]), .A2(n838), .B1(n1082), .B2(\mem[13][2] ), 
        .ZN(n1080) );
  INV_X1 U299 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U300 ( .A1(data_in[3]), .A2(n838), .B1(n1082), .B2(\mem[13][3] ), 
        .ZN(n1079) );
  INV_X1 U301 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U302 ( .A1(data_in[4]), .A2(n838), .B1(n1082), .B2(\mem[13][4] ), 
        .ZN(n1078) );
  INV_X1 U303 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U304 ( .A1(data_in[5]), .A2(n838), .B1(n1082), .B2(\mem[13][5] ), 
        .ZN(n1077) );
  INV_X1 U305 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U306 ( .A1(data_in[6]), .A2(n838), .B1(n1082), .B2(\mem[13][6] ), 
        .ZN(n1076) );
  INV_X1 U307 ( .A(n1075), .ZN(n772) );
  AOI22_X1 U308 ( .A1(data_in[7]), .A2(n838), .B1(n1082), .B2(\mem[13][7] ), 
        .ZN(n1075) );
  INV_X1 U309 ( .A(n1074), .ZN(n771) );
  AOI22_X1 U310 ( .A1(data_in[0]), .A2(n837), .B1(n1073), .B2(\mem[14][0] ), 
        .ZN(n1074) );
  INV_X1 U311 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U312 ( .A1(data_in[1]), .A2(n837), .B1(n1073), .B2(\mem[14][1] ), 
        .ZN(n1072) );
  INV_X1 U313 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U314 ( .A1(data_in[2]), .A2(n837), .B1(n1073), .B2(\mem[14][2] ), 
        .ZN(n1071) );
  INV_X1 U315 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U316 ( .A1(data_in[3]), .A2(n837), .B1(n1073), .B2(\mem[14][3] ), 
        .ZN(n1070) );
  INV_X1 U317 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U318 ( .A1(data_in[4]), .A2(n837), .B1(n1073), .B2(\mem[14][4] ), 
        .ZN(n1069) );
  INV_X1 U319 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U320 ( .A1(data_in[5]), .A2(n837), .B1(n1073), .B2(\mem[14][5] ), 
        .ZN(n1068) );
  INV_X1 U321 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U322 ( .A1(data_in[6]), .A2(n837), .B1(n1073), .B2(\mem[14][6] ), 
        .ZN(n1067) );
  INV_X1 U323 ( .A(n1066), .ZN(n764) );
  AOI22_X1 U324 ( .A1(data_in[7]), .A2(n837), .B1(n1073), .B2(\mem[14][7] ), 
        .ZN(n1066) );
  INV_X1 U325 ( .A(n1065), .ZN(n763) );
  AOI22_X1 U326 ( .A1(data_in[0]), .A2(n836), .B1(n1064), .B2(\mem[15][0] ), 
        .ZN(n1065) );
  INV_X1 U327 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U328 ( .A1(data_in[1]), .A2(n836), .B1(n1064), .B2(\mem[15][1] ), 
        .ZN(n1063) );
  INV_X1 U329 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U330 ( .A1(data_in[2]), .A2(n836), .B1(n1064), .B2(\mem[15][2] ), 
        .ZN(n1062) );
  INV_X1 U331 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U332 ( .A1(data_in[3]), .A2(n836), .B1(n1064), .B2(\mem[15][3] ), 
        .ZN(n1061) );
  INV_X1 U333 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U334 ( .A1(data_in[4]), .A2(n836), .B1(n1064), .B2(\mem[15][4] ), 
        .ZN(n1060) );
  INV_X1 U335 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U336 ( .A1(data_in[5]), .A2(n836), .B1(n1064), .B2(\mem[15][5] ), 
        .ZN(n1059) );
  INV_X1 U337 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U338 ( .A1(data_in[6]), .A2(n836), .B1(n1064), .B2(\mem[15][6] ), 
        .ZN(n1058) );
  INV_X1 U339 ( .A(n1057), .ZN(n756) );
  AOI22_X1 U340 ( .A1(data_in[7]), .A2(n836), .B1(n1064), .B2(\mem[15][7] ), 
        .ZN(n1057) );
  INV_X1 U341 ( .A(n1056), .ZN(n755) );
  AOI22_X1 U342 ( .A1(data_in[0]), .A2(n835), .B1(n1055), .B2(\mem[16][0] ), 
        .ZN(n1056) );
  INV_X1 U343 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U344 ( .A1(data_in[1]), .A2(n835), .B1(n1055), .B2(\mem[16][1] ), 
        .ZN(n1054) );
  INV_X1 U345 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U346 ( .A1(data_in[2]), .A2(n835), .B1(n1055), .B2(\mem[16][2] ), 
        .ZN(n1053) );
  INV_X1 U347 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U348 ( .A1(data_in[3]), .A2(n835), .B1(n1055), .B2(\mem[16][3] ), 
        .ZN(n1052) );
  INV_X1 U349 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U350 ( .A1(data_in[4]), .A2(n835), .B1(n1055), .B2(\mem[16][4] ), 
        .ZN(n1051) );
  INV_X1 U351 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U352 ( .A1(data_in[5]), .A2(n835), .B1(n1055), .B2(\mem[16][5] ), 
        .ZN(n1050) );
  INV_X1 U353 ( .A(n1049), .ZN(n749) );
  AOI22_X1 U354 ( .A1(data_in[6]), .A2(n835), .B1(n1055), .B2(\mem[16][6] ), 
        .ZN(n1049) );
  INV_X1 U355 ( .A(n1048), .ZN(n748) );
  AOI22_X1 U356 ( .A1(data_in[7]), .A2(n835), .B1(n1055), .B2(\mem[16][7] ), 
        .ZN(n1048) );
  INV_X1 U357 ( .A(n1046), .ZN(n747) );
  AOI22_X1 U358 ( .A1(data_in[0]), .A2(n834), .B1(n1045), .B2(\mem[17][0] ), 
        .ZN(n1046) );
  INV_X1 U359 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U360 ( .A1(data_in[1]), .A2(n834), .B1(n1045), .B2(\mem[17][1] ), 
        .ZN(n1044) );
  INV_X1 U361 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U362 ( .A1(data_in[2]), .A2(n834), .B1(n1045), .B2(\mem[17][2] ), 
        .ZN(n1043) );
  INV_X1 U363 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U364 ( .A1(data_in[3]), .A2(n834), .B1(n1045), .B2(\mem[17][3] ), 
        .ZN(n1042) );
  INV_X1 U365 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U366 ( .A1(data_in[4]), .A2(n834), .B1(n1045), .B2(\mem[17][4] ), 
        .ZN(n1041) );
  INV_X1 U367 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U368 ( .A1(data_in[5]), .A2(n834), .B1(n1045), .B2(\mem[17][5] ), 
        .ZN(n1040) );
  INV_X1 U369 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U370 ( .A1(data_in[6]), .A2(n834), .B1(n1045), .B2(\mem[17][6] ), 
        .ZN(n1039) );
  INV_X1 U371 ( .A(n1038), .ZN(n740) );
  AOI22_X1 U372 ( .A1(data_in[7]), .A2(n834), .B1(n1045), .B2(\mem[17][7] ), 
        .ZN(n1038) );
  INV_X1 U373 ( .A(n1037), .ZN(n739) );
  AOI22_X1 U374 ( .A1(data_in[0]), .A2(n833), .B1(n1036), .B2(\mem[18][0] ), 
        .ZN(n1037) );
  INV_X1 U375 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U376 ( .A1(data_in[1]), .A2(n833), .B1(n1036), .B2(\mem[18][1] ), 
        .ZN(n1035) );
  INV_X1 U377 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U378 ( .A1(data_in[2]), .A2(n833), .B1(n1036), .B2(\mem[18][2] ), 
        .ZN(n1034) );
  INV_X1 U379 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U380 ( .A1(data_in[3]), .A2(n833), .B1(n1036), .B2(\mem[18][3] ), 
        .ZN(n1033) );
  INV_X1 U381 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U382 ( .A1(data_in[4]), .A2(n833), .B1(n1036), .B2(\mem[18][4] ), 
        .ZN(n1032) );
  INV_X1 U383 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U384 ( .A1(data_in[5]), .A2(n833), .B1(n1036), .B2(\mem[18][5] ), 
        .ZN(n1031) );
  INV_X1 U385 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U386 ( .A1(data_in[6]), .A2(n833), .B1(n1036), .B2(\mem[18][6] ), 
        .ZN(n1030) );
  INV_X1 U387 ( .A(n1029), .ZN(n732) );
  AOI22_X1 U388 ( .A1(data_in[7]), .A2(n833), .B1(n1036), .B2(\mem[18][7] ), 
        .ZN(n1029) );
  INV_X1 U389 ( .A(n1028), .ZN(n731) );
  AOI22_X1 U390 ( .A1(data_in[0]), .A2(n832), .B1(n1027), .B2(\mem[19][0] ), 
        .ZN(n1028) );
  INV_X1 U391 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U392 ( .A1(data_in[1]), .A2(n832), .B1(n1027), .B2(\mem[19][1] ), 
        .ZN(n1026) );
  INV_X1 U393 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U394 ( .A1(data_in[2]), .A2(n832), .B1(n1027), .B2(\mem[19][2] ), 
        .ZN(n1025) );
  INV_X1 U395 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U396 ( .A1(data_in[3]), .A2(n832), .B1(n1027), .B2(\mem[19][3] ), 
        .ZN(n1024) );
  INV_X1 U397 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U398 ( .A1(data_in[4]), .A2(n832), .B1(n1027), .B2(\mem[19][4] ), 
        .ZN(n1023) );
  INV_X1 U399 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U400 ( .A1(data_in[5]), .A2(n832), .B1(n1027), .B2(\mem[19][5] ), 
        .ZN(n1022) );
  INV_X1 U401 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U402 ( .A1(data_in[6]), .A2(n832), .B1(n1027), .B2(\mem[19][6] ), 
        .ZN(n1021) );
  INV_X1 U403 ( .A(n1020), .ZN(n724) );
  AOI22_X1 U404 ( .A1(data_in[7]), .A2(n832), .B1(n1027), .B2(\mem[19][7] ), 
        .ZN(n1020) );
  INV_X1 U405 ( .A(n1019), .ZN(n723) );
  AOI22_X1 U406 ( .A1(data_in[0]), .A2(n831), .B1(n1018), .B2(\mem[20][0] ), 
        .ZN(n1019) );
  INV_X1 U407 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U408 ( .A1(data_in[1]), .A2(n831), .B1(n1018), .B2(\mem[20][1] ), 
        .ZN(n1017) );
  INV_X1 U409 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U410 ( .A1(data_in[2]), .A2(n831), .B1(n1018), .B2(\mem[20][2] ), 
        .ZN(n1016) );
  INV_X1 U411 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U412 ( .A1(data_in[3]), .A2(n831), .B1(n1018), .B2(\mem[20][3] ), 
        .ZN(n1015) );
  INV_X1 U413 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U414 ( .A1(data_in[4]), .A2(n831), .B1(n1018), .B2(\mem[20][4] ), 
        .ZN(n1014) );
  INV_X1 U415 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U416 ( .A1(data_in[5]), .A2(n831), .B1(n1018), .B2(\mem[20][5] ), 
        .ZN(n1013) );
  INV_X1 U417 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U418 ( .A1(data_in[6]), .A2(n831), .B1(n1018), .B2(\mem[20][6] ), 
        .ZN(n1012) );
  INV_X1 U419 ( .A(n1011), .ZN(n716) );
  AOI22_X1 U420 ( .A1(data_in[7]), .A2(n831), .B1(n1018), .B2(\mem[20][7] ), 
        .ZN(n1011) );
  INV_X1 U421 ( .A(n1010), .ZN(n715) );
  AOI22_X1 U422 ( .A1(data_in[0]), .A2(n830), .B1(n1009), .B2(\mem[21][0] ), 
        .ZN(n1010) );
  INV_X1 U423 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U424 ( .A1(data_in[1]), .A2(n830), .B1(n1009), .B2(\mem[21][1] ), 
        .ZN(n1008) );
  INV_X1 U425 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U426 ( .A1(data_in[2]), .A2(n830), .B1(n1009), .B2(\mem[21][2] ), 
        .ZN(n1007) );
  INV_X1 U427 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U428 ( .A1(data_in[3]), .A2(n830), .B1(n1009), .B2(\mem[21][3] ), 
        .ZN(n1006) );
  INV_X1 U429 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U430 ( .A1(data_in[4]), .A2(n830), .B1(n1009), .B2(\mem[21][4] ), 
        .ZN(n1005) );
  INV_X1 U431 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U432 ( .A1(data_in[5]), .A2(n830), .B1(n1009), .B2(\mem[21][5] ), 
        .ZN(n1004) );
  INV_X1 U433 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U434 ( .A1(data_in[6]), .A2(n830), .B1(n1009), .B2(\mem[21][6] ), 
        .ZN(n1003) );
  INV_X1 U435 ( .A(n1002), .ZN(n708) );
  AOI22_X1 U436 ( .A1(data_in[7]), .A2(n830), .B1(n1009), .B2(\mem[21][7] ), 
        .ZN(n1002) );
  INV_X1 U437 ( .A(n1001), .ZN(n707) );
  AOI22_X1 U438 ( .A1(data_in[0]), .A2(n829), .B1(n1000), .B2(\mem[22][0] ), 
        .ZN(n1001) );
  INV_X1 U439 ( .A(n999), .ZN(n706) );
  AOI22_X1 U440 ( .A1(data_in[1]), .A2(n829), .B1(n1000), .B2(\mem[22][1] ), 
        .ZN(n999) );
  INV_X1 U441 ( .A(n998), .ZN(n705) );
  AOI22_X1 U442 ( .A1(data_in[2]), .A2(n829), .B1(n1000), .B2(\mem[22][2] ), 
        .ZN(n998) );
  INV_X1 U443 ( .A(n997), .ZN(n704) );
  AOI22_X1 U444 ( .A1(data_in[3]), .A2(n829), .B1(n1000), .B2(\mem[22][3] ), 
        .ZN(n997) );
  INV_X1 U445 ( .A(n996), .ZN(n703) );
  AOI22_X1 U446 ( .A1(data_in[4]), .A2(n829), .B1(n1000), .B2(\mem[22][4] ), 
        .ZN(n996) );
  INV_X1 U447 ( .A(n995), .ZN(n702) );
  AOI22_X1 U448 ( .A1(data_in[5]), .A2(n829), .B1(n1000), .B2(\mem[22][5] ), 
        .ZN(n995) );
  INV_X1 U449 ( .A(n994), .ZN(n701) );
  AOI22_X1 U450 ( .A1(data_in[6]), .A2(n829), .B1(n1000), .B2(\mem[22][6] ), 
        .ZN(n994) );
  INV_X1 U451 ( .A(n993), .ZN(n700) );
  AOI22_X1 U452 ( .A1(data_in[7]), .A2(n829), .B1(n1000), .B2(\mem[22][7] ), 
        .ZN(n993) );
  INV_X1 U453 ( .A(n992), .ZN(n699) );
  AOI22_X1 U454 ( .A1(data_in[0]), .A2(n828), .B1(n991), .B2(\mem[23][0] ), 
        .ZN(n992) );
  INV_X1 U455 ( .A(n990), .ZN(n698) );
  AOI22_X1 U456 ( .A1(data_in[1]), .A2(n828), .B1(n991), .B2(\mem[23][1] ), 
        .ZN(n990) );
  INV_X1 U457 ( .A(n989), .ZN(n697) );
  AOI22_X1 U458 ( .A1(data_in[2]), .A2(n828), .B1(n991), .B2(\mem[23][2] ), 
        .ZN(n989) );
  INV_X1 U459 ( .A(n988), .ZN(n696) );
  AOI22_X1 U460 ( .A1(data_in[3]), .A2(n828), .B1(n991), .B2(\mem[23][3] ), 
        .ZN(n988) );
  INV_X1 U461 ( .A(n987), .ZN(n695) );
  AOI22_X1 U462 ( .A1(data_in[4]), .A2(n828), .B1(n991), .B2(\mem[23][4] ), 
        .ZN(n987) );
  INV_X1 U463 ( .A(n986), .ZN(n694) );
  AOI22_X1 U464 ( .A1(data_in[5]), .A2(n828), .B1(n991), .B2(\mem[23][5] ), 
        .ZN(n986) );
  INV_X1 U465 ( .A(n985), .ZN(n693) );
  AOI22_X1 U466 ( .A1(data_in[6]), .A2(n828), .B1(n991), .B2(\mem[23][6] ), 
        .ZN(n985) );
  INV_X1 U467 ( .A(n984), .ZN(n692) );
  AOI22_X1 U468 ( .A1(data_in[7]), .A2(n828), .B1(n991), .B2(\mem[23][7] ), 
        .ZN(n984) );
  INV_X1 U469 ( .A(n983), .ZN(n691) );
  AOI22_X1 U470 ( .A1(data_in[0]), .A2(n827), .B1(n982), .B2(\mem[24][0] ), 
        .ZN(n983) );
  INV_X1 U471 ( .A(n981), .ZN(n690) );
  AOI22_X1 U472 ( .A1(data_in[1]), .A2(n827), .B1(n982), .B2(\mem[24][1] ), 
        .ZN(n981) );
  INV_X1 U473 ( .A(n980), .ZN(n689) );
  AOI22_X1 U474 ( .A1(data_in[2]), .A2(n827), .B1(n982), .B2(\mem[24][2] ), 
        .ZN(n980) );
  INV_X1 U475 ( .A(n979), .ZN(n688) );
  AOI22_X1 U476 ( .A1(data_in[3]), .A2(n827), .B1(n982), .B2(\mem[24][3] ), 
        .ZN(n979) );
  INV_X1 U477 ( .A(n978), .ZN(n687) );
  AOI22_X1 U478 ( .A1(data_in[4]), .A2(n827), .B1(n982), .B2(\mem[24][4] ), 
        .ZN(n978) );
  INV_X1 U479 ( .A(n977), .ZN(n686) );
  AOI22_X1 U480 ( .A1(data_in[5]), .A2(n827), .B1(n982), .B2(\mem[24][5] ), 
        .ZN(n977) );
  INV_X1 U481 ( .A(n976), .ZN(n685) );
  AOI22_X1 U482 ( .A1(data_in[6]), .A2(n827), .B1(n982), .B2(\mem[24][6] ), 
        .ZN(n976) );
  INV_X1 U483 ( .A(n975), .ZN(n684) );
  AOI22_X1 U484 ( .A1(data_in[7]), .A2(n827), .B1(n982), .B2(\mem[24][7] ), 
        .ZN(n975) );
  INV_X1 U485 ( .A(n973), .ZN(n683) );
  AOI22_X1 U486 ( .A1(data_in[0]), .A2(n826), .B1(n972), .B2(\mem[25][0] ), 
        .ZN(n973) );
  INV_X1 U487 ( .A(n971), .ZN(n682) );
  AOI22_X1 U488 ( .A1(data_in[1]), .A2(n826), .B1(n972), .B2(\mem[25][1] ), 
        .ZN(n971) );
  INV_X1 U489 ( .A(n970), .ZN(n681) );
  AOI22_X1 U490 ( .A1(data_in[2]), .A2(n826), .B1(n972), .B2(\mem[25][2] ), 
        .ZN(n970) );
  INV_X1 U491 ( .A(n969), .ZN(n680) );
  AOI22_X1 U492 ( .A1(data_in[3]), .A2(n826), .B1(n972), .B2(\mem[25][3] ), 
        .ZN(n969) );
  INV_X1 U493 ( .A(n968), .ZN(n679) );
  AOI22_X1 U494 ( .A1(data_in[4]), .A2(n826), .B1(n972), .B2(\mem[25][4] ), 
        .ZN(n968) );
  INV_X1 U495 ( .A(n967), .ZN(n678) );
  AOI22_X1 U496 ( .A1(data_in[5]), .A2(n826), .B1(n972), .B2(\mem[25][5] ), 
        .ZN(n967) );
  INV_X1 U497 ( .A(n966), .ZN(n677) );
  AOI22_X1 U498 ( .A1(data_in[6]), .A2(n826), .B1(n972), .B2(\mem[25][6] ), 
        .ZN(n966) );
  INV_X1 U499 ( .A(n965), .ZN(n676) );
  AOI22_X1 U500 ( .A1(data_in[7]), .A2(n826), .B1(n972), .B2(\mem[25][7] ), 
        .ZN(n965) );
  INV_X1 U501 ( .A(n964), .ZN(n675) );
  AOI22_X1 U502 ( .A1(data_in[0]), .A2(n825), .B1(n963), .B2(\mem[26][0] ), 
        .ZN(n964) );
  INV_X1 U503 ( .A(n962), .ZN(n674) );
  AOI22_X1 U504 ( .A1(data_in[1]), .A2(n825), .B1(n963), .B2(\mem[26][1] ), 
        .ZN(n962) );
  INV_X1 U505 ( .A(n961), .ZN(n673) );
  AOI22_X1 U506 ( .A1(data_in[2]), .A2(n825), .B1(n963), .B2(\mem[26][2] ), 
        .ZN(n961) );
  INV_X1 U507 ( .A(n960), .ZN(n672) );
  AOI22_X1 U508 ( .A1(data_in[3]), .A2(n825), .B1(n963), .B2(\mem[26][3] ), 
        .ZN(n960) );
  INV_X1 U509 ( .A(n959), .ZN(n671) );
  AOI22_X1 U510 ( .A1(data_in[4]), .A2(n825), .B1(n963), .B2(\mem[26][4] ), 
        .ZN(n959) );
  INV_X1 U511 ( .A(n958), .ZN(n670) );
  AOI22_X1 U512 ( .A1(data_in[5]), .A2(n825), .B1(n963), .B2(\mem[26][5] ), 
        .ZN(n958) );
  INV_X1 U513 ( .A(n957), .ZN(n669) );
  AOI22_X1 U514 ( .A1(data_in[6]), .A2(n825), .B1(n963), .B2(\mem[26][6] ), 
        .ZN(n957) );
  INV_X1 U515 ( .A(n956), .ZN(n668) );
  AOI22_X1 U516 ( .A1(data_in[7]), .A2(n825), .B1(n963), .B2(\mem[26][7] ), 
        .ZN(n956) );
  INV_X1 U517 ( .A(n955), .ZN(n667) );
  AOI22_X1 U518 ( .A1(data_in[0]), .A2(n824), .B1(n954), .B2(\mem[27][0] ), 
        .ZN(n955) );
  INV_X1 U519 ( .A(n953), .ZN(n666) );
  AOI22_X1 U520 ( .A1(data_in[1]), .A2(n824), .B1(n954), .B2(\mem[27][1] ), 
        .ZN(n953) );
  INV_X1 U521 ( .A(n952), .ZN(n665) );
  AOI22_X1 U522 ( .A1(data_in[2]), .A2(n824), .B1(n954), .B2(\mem[27][2] ), 
        .ZN(n952) );
  INV_X1 U523 ( .A(n951), .ZN(n664) );
  AOI22_X1 U524 ( .A1(data_in[3]), .A2(n824), .B1(n954), .B2(\mem[27][3] ), 
        .ZN(n951) );
  INV_X1 U525 ( .A(n950), .ZN(n663) );
  AOI22_X1 U526 ( .A1(data_in[4]), .A2(n824), .B1(n954), .B2(\mem[27][4] ), 
        .ZN(n950) );
  INV_X1 U527 ( .A(n949), .ZN(n662) );
  AOI22_X1 U528 ( .A1(data_in[5]), .A2(n824), .B1(n954), .B2(\mem[27][5] ), 
        .ZN(n949) );
  INV_X1 U529 ( .A(n948), .ZN(n661) );
  AOI22_X1 U530 ( .A1(data_in[6]), .A2(n824), .B1(n954), .B2(\mem[27][6] ), 
        .ZN(n948) );
  INV_X1 U531 ( .A(n947), .ZN(n660) );
  AOI22_X1 U532 ( .A1(data_in[7]), .A2(n824), .B1(n954), .B2(\mem[27][7] ), 
        .ZN(n947) );
  INV_X1 U533 ( .A(n946), .ZN(n659) );
  AOI22_X1 U534 ( .A1(data_in[0]), .A2(n823), .B1(n945), .B2(\mem[28][0] ), 
        .ZN(n946) );
  INV_X1 U535 ( .A(n944), .ZN(n658) );
  AOI22_X1 U536 ( .A1(data_in[1]), .A2(n823), .B1(n945), .B2(\mem[28][1] ), 
        .ZN(n944) );
  INV_X1 U537 ( .A(n943), .ZN(n657) );
  AOI22_X1 U538 ( .A1(data_in[2]), .A2(n823), .B1(n945), .B2(\mem[28][2] ), 
        .ZN(n943) );
  INV_X1 U539 ( .A(n942), .ZN(n656) );
  AOI22_X1 U540 ( .A1(data_in[3]), .A2(n823), .B1(n945), .B2(\mem[28][3] ), 
        .ZN(n942) );
  INV_X1 U541 ( .A(n941), .ZN(n655) );
  AOI22_X1 U542 ( .A1(data_in[4]), .A2(n823), .B1(n945), .B2(\mem[28][4] ), 
        .ZN(n941) );
  INV_X1 U543 ( .A(n940), .ZN(n654) );
  AOI22_X1 U544 ( .A1(data_in[5]), .A2(n823), .B1(n945), .B2(\mem[28][5] ), 
        .ZN(n940) );
  INV_X1 U545 ( .A(n939), .ZN(n653) );
  AOI22_X1 U546 ( .A1(data_in[6]), .A2(n823), .B1(n945), .B2(\mem[28][6] ), 
        .ZN(n939) );
  INV_X1 U547 ( .A(n938), .ZN(n652) );
  AOI22_X1 U548 ( .A1(data_in[7]), .A2(n823), .B1(n945), .B2(\mem[28][7] ), 
        .ZN(n938) );
  INV_X1 U549 ( .A(n937), .ZN(n651) );
  AOI22_X1 U550 ( .A1(data_in[0]), .A2(n822), .B1(n936), .B2(\mem[29][0] ), 
        .ZN(n937) );
  INV_X1 U551 ( .A(n935), .ZN(n650) );
  AOI22_X1 U552 ( .A1(data_in[1]), .A2(n822), .B1(n936), .B2(\mem[29][1] ), 
        .ZN(n935) );
  INV_X1 U553 ( .A(n934), .ZN(n649) );
  AOI22_X1 U554 ( .A1(data_in[2]), .A2(n822), .B1(n936), .B2(\mem[29][2] ), 
        .ZN(n934) );
  INV_X1 U555 ( .A(n933), .ZN(n648) );
  AOI22_X1 U556 ( .A1(data_in[3]), .A2(n822), .B1(n936), .B2(\mem[29][3] ), 
        .ZN(n933) );
  INV_X1 U557 ( .A(n932), .ZN(n647) );
  AOI22_X1 U558 ( .A1(data_in[4]), .A2(n822), .B1(n936), .B2(\mem[29][4] ), 
        .ZN(n932) );
  INV_X1 U559 ( .A(n931), .ZN(n646) );
  AOI22_X1 U560 ( .A1(data_in[5]), .A2(n822), .B1(n936), .B2(\mem[29][5] ), 
        .ZN(n931) );
  INV_X1 U561 ( .A(n930), .ZN(n645) );
  AOI22_X1 U562 ( .A1(data_in[6]), .A2(n822), .B1(n936), .B2(\mem[29][6] ), 
        .ZN(n930) );
  INV_X1 U563 ( .A(n929), .ZN(n644) );
  AOI22_X1 U564 ( .A1(data_in[7]), .A2(n822), .B1(n936), .B2(\mem[29][7] ), 
        .ZN(n929) );
  INV_X1 U565 ( .A(n928), .ZN(n643) );
  AOI22_X1 U566 ( .A1(data_in[0]), .A2(n821), .B1(n927), .B2(\mem[30][0] ), 
        .ZN(n928) );
  INV_X1 U567 ( .A(n926), .ZN(n642) );
  AOI22_X1 U568 ( .A1(data_in[1]), .A2(n821), .B1(n927), .B2(\mem[30][1] ), 
        .ZN(n926) );
  INV_X1 U569 ( .A(n925), .ZN(n641) );
  AOI22_X1 U570 ( .A1(data_in[2]), .A2(n821), .B1(n927), .B2(\mem[30][2] ), 
        .ZN(n925) );
  INV_X1 U571 ( .A(n924), .ZN(n640) );
  AOI22_X1 U572 ( .A1(data_in[3]), .A2(n821), .B1(n927), .B2(\mem[30][3] ), 
        .ZN(n924) );
  INV_X1 U573 ( .A(n923), .ZN(n639) );
  AOI22_X1 U574 ( .A1(data_in[4]), .A2(n821), .B1(n927), .B2(\mem[30][4] ), 
        .ZN(n923) );
  INV_X1 U575 ( .A(n922), .ZN(n638) );
  AOI22_X1 U576 ( .A1(data_in[5]), .A2(n821), .B1(n927), .B2(\mem[30][5] ), 
        .ZN(n922) );
  INV_X1 U577 ( .A(n921), .ZN(n637) );
  AOI22_X1 U578 ( .A1(data_in[6]), .A2(n821), .B1(n927), .B2(\mem[30][6] ), 
        .ZN(n921) );
  INV_X1 U579 ( .A(n920), .ZN(n636) );
  AOI22_X1 U580 ( .A1(data_in[7]), .A2(n821), .B1(n927), .B2(\mem[30][7] ), 
        .ZN(n920) );
  INV_X1 U581 ( .A(n919), .ZN(n635) );
  AOI22_X1 U582 ( .A1(data_in[0]), .A2(n820), .B1(n918), .B2(\mem[31][0] ), 
        .ZN(n919) );
  INV_X1 U583 ( .A(n917), .ZN(n634) );
  AOI22_X1 U584 ( .A1(data_in[1]), .A2(n820), .B1(n918), .B2(\mem[31][1] ), 
        .ZN(n917) );
  INV_X1 U585 ( .A(n916), .ZN(n633) );
  AOI22_X1 U586 ( .A1(data_in[2]), .A2(n820), .B1(n918), .B2(\mem[31][2] ), 
        .ZN(n916) );
  INV_X1 U587 ( .A(n915), .ZN(n632) );
  AOI22_X1 U588 ( .A1(data_in[3]), .A2(n820), .B1(n918), .B2(\mem[31][3] ), 
        .ZN(n915) );
  INV_X1 U589 ( .A(n914), .ZN(n631) );
  AOI22_X1 U590 ( .A1(data_in[4]), .A2(n820), .B1(n918), .B2(\mem[31][4] ), 
        .ZN(n914) );
  INV_X1 U591 ( .A(n913), .ZN(n630) );
  AOI22_X1 U592 ( .A1(data_in[5]), .A2(n820), .B1(n918), .B2(\mem[31][5] ), 
        .ZN(n913) );
  INV_X1 U593 ( .A(n912), .ZN(n629) );
  AOI22_X1 U594 ( .A1(data_in[6]), .A2(n820), .B1(n918), .B2(\mem[31][6] ), 
        .ZN(n912) );
  INV_X1 U595 ( .A(n911), .ZN(n628) );
  AOI22_X1 U596 ( .A1(data_in[7]), .A2(n820), .B1(n918), .B2(\mem[31][7] ), 
        .ZN(n911) );
  MUX2_X1 U597 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n611), .Z(n1) );
  MUX2_X1 U598 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n611), .Z(n2) );
  MUX2_X1 U599 ( .A(n2), .B(n1), .S(n608), .Z(n3) );
  MUX2_X1 U600 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n611), .Z(n4) );
  MUX2_X1 U601 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n611), .Z(n5) );
  MUX2_X1 U602 ( .A(n5), .B(n4), .S(n608), .Z(n6) );
  MUX2_X1 U603 ( .A(n6), .B(n3), .S(N12), .Z(n7) );
  MUX2_X1 U604 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n611), .Z(n8) );
  MUX2_X1 U605 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n611), .Z(n9) );
  MUX2_X1 U606 ( .A(n9), .B(n8), .S(n608), .Z(n10) );
  MUX2_X1 U607 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n611), .Z(n11) );
  MUX2_X1 U608 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n611), .Z(n12) );
  MUX2_X1 U609 ( .A(n12), .B(n11), .S(n608), .Z(n13) );
  MUX2_X1 U610 ( .A(n13), .B(n10), .S(n606), .Z(n14) );
  MUX2_X1 U611 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U612 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n615), .Z(n16) );
  MUX2_X1 U613 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n617), .Z(n17) );
  MUX2_X1 U614 ( .A(n17), .B(n16), .S(n609), .Z(n18) );
  MUX2_X1 U615 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n614), .Z(n19) );
  MUX2_X1 U616 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n615), .Z(n20) );
  MUX2_X1 U617 ( .A(n20), .B(n19), .S(n609), .Z(n21) );
  MUX2_X1 U618 ( .A(n21), .B(n18), .S(n607), .Z(n22) );
  MUX2_X1 U619 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n617), .Z(n23) );
  MUX2_X1 U620 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n617), .Z(n24) );
  MUX2_X1 U621 ( .A(n24), .B(n23), .S(n609), .Z(n25) );
  MUX2_X1 U622 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n616), .Z(n26) );
  MUX2_X1 U623 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n617), .Z(n27) );
  MUX2_X1 U624 ( .A(n27), .B(n26), .S(n609), .Z(n28) );
  MUX2_X1 U625 ( .A(n28), .B(n25), .S(n607), .Z(n29) );
  MUX2_X1 U626 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U627 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U628 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n611), .Z(n31) );
  MUX2_X1 U629 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n611), .Z(n32) );
  MUX2_X1 U630 ( .A(n32), .B(n31), .S(n609), .Z(n33) );
  MUX2_X1 U631 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n611), .Z(n34) );
  MUX2_X1 U632 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n613), .Z(n35) );
  MUX2_X1 U633 ( .A(n35), .B(n34), .S(n609), .Z(n36) );
  MUX2_X1 U634 ( .A(n36), .B(n33), .S(n607), .Z(n37) );
  MUX2_X1 U635 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n613), .Z(n38) );
  MUX2_X1 U636 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(N10), .Z(n39) );
  MUX2_X1 U637 ( .A(n39), .B(n38), .S(n609), .Z(n40) );
  MUX2_X1 U638 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n613), .Z(n41) );
  MUX2_X1 U639 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(N10), .Z(n42) );
  MUX2_X1 U640 ( .A(n42), .B(n41), .S(n609), .Z(n43) );
  MUX2_X1 U641 ( .A(n43), .B(n40), .S(N12), .Z(n44) );
  MUX2_X1 U642 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U643 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(N10), .Z(n46) );
  MUX2_X1 U644 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n617), .Z(n47) );
  MUX2_X1 U645 ( .A(n47), .B(n46), .S(n609), .Z(n48) );
  MUX2_X1 U646 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n614), .Z(n49) );
  MUX2_X1 U647 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(N10), .Z(n50) );
  MUX2_X1 U648 ( .A(n50), .B(n49), .S(n609), .Z(n51) );
  MUX2_X1 U649 ( .A(n51), .B(n48), .S(n606), .Z(n52) );
  MUX2_X1 U650 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n617), .Z(n53) );
  MUX2_X1 U651 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n54) );
  MUX2_X1 U652 ( .A(n54), .B(n53), .S(n609), .Z(n55) );
  MUX2_X1 U653 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(N10), .Z(n56) );
  MUX2_X1 U654 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n616), .Z(n57) );
  MUX2_X1 U655 ( .A(n57), .B(n56), .S(n609), .Z(n58) );
  MUX2_X1 U656 ( .A(n58), .B(n55), .S(N12), .Z(n59) );
  MUX2_X1 U657 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U658 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U659 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n612), .Z(n61) );
  MUX2_X1 U660 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n612), .Z(n62) );
  MUX2_X1 U661 ( .A(n62), .B(n61), .S(n610), .Z(n63) );
  MUX2_X1 U662 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n612), .Z(n64) );
  MUX2_X1 U663 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n612), .Z(n65) );
  MUX2_X1 U664 ( .A(n65), .B(n64), .S(n610), .Z(n66) );
  MUX2_X1 U665 ( .A(n66), .B(n63), .S(n606), .Z(n67) );
  MUX2_X1 U666 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n612), .Z(n68) );
  MUX2_X1 U667 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n612), .Z(n69) );
  MUX2_X1 U668 ( .A(n69), .B(n68), .S(n610), .Z(n70) );
  MUX2_X1 U669 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n612), .Z(n71) );
  MUX2_X1 U670 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n612), .Z(n72) );
  MUX2_X1 U671 ( .A(n72), .B(n71), .S(n610), .Z(n73) );
  MUX2_X1 U672 ( .A(n73), .B(n70), .S(n606), .Z(n74) );
  MUX2_X1 U673 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U674 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n612), .Z(n76) );
  MUX2_X1 U675 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n612), .Z(n77) );
  MUX2_X1 U676 ( .A(n77), .B(n76), .S(n610), .Z(n78) );
  MUX2_X1 U677 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n612), .Z(n79) );
  MUX2_X1 U678 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n612), .Z(n80) );
  MUX2_X1 U679 ( .A(n80), .B(n79), .S(n610), .Z(n81) );
  MUX2_X1 U680 ( .A(n81), .B(n78), .S(n606), .Z(n82) );
  MUX2_X1 U681 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n613), .Z(n83) );
  MUX2_X1 U682 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n613), .Z(n84) );
  MUX2_X1 U683 ( .A(n84), .B(n83), .S(n610), .Z(n85) );
  MUX2_X1 U684 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n613), .Z(n86) );
  MUX2_X1 U685 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n613), .Z(n87) );
  MUX2_X1 U686 ( .A(n87), .B(n86), .S(n610), .Z(n88) );
  MUX2_X1 U687 ( .A(n88), .B(n85), .S(n606), .Z(n89) );
  MUX2_X1 U688 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U689 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U690 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n613), .Z(n91) );
  MUX2_X1 U691 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n613), .Z(n92) );
  MUX2_X1 U692 ( .A(n92), .B(n91), .S(n610), .Z(n93) );
  MUX2_X1 U693 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n613), .Z(n94) );
  MUX2_X1 U694 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n613), .Z(n95) );
  MUX2_X1 U695 ( .A(n95), .B(n94), .S(n610), .Z(n96) );
  MUX2_X1 U696 ( .A(n96), .B(n93), .S(n606), .Z(n97) );
  MUX2_X1 U697 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n613), .Z(n98) );
  MUX2_X1 U698 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n613), .Z(n99) );
  MUX2_X1 U699 ( .A(n99), .B(n98), .S(n610), .Z(n100) );
  MUX2_X1 U700 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n613), .Z(n101) );
  MUX2_X1 U701 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n613), .Z(n102) );
  MUX2_X1 U702 ( .A(n102), .B(n101), .S(n610), .Z(n103) );
  MUX2_X1 U703 ( .A(n103), .B(n100), .S(n606), .Z(n104) );
  MUX2_X1 U704 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U705 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n616), .Z(n106) );
  MUX2_X1 U706 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n612), .Z(n107) );
  MUX2_X1 U707 ( .A(n107), .B(n106), .S(n610), .Z(n108) );
  MUX2_X1 U708 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n612), .Z(n109) );
  MUX2_X1 U709 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n613), .Z(n110) );
  MUX2_X1 U710 ( .A(n110), .B(n109), .S(n610), .Z(n111) );
  MUX2_X1 U711 ( .A(n111), .B(n108), .S(n606), .Z(n112) );
  MUX2_X1 U712 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n614), .Z(n113) );
  MUX2_X1 U713 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n615), .Z(n114) );
  MUX2_X1 U714 ( .A(n114), .B(n113), .S(n608), .Z(n115) );
  MUX2_X1 U715 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n616), .Z(n116) );
  MUX2_X1 U716 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n614), .Z(n117) );
  MUX2_X1 U717 ( .A(n117), .B(n116), .S(n609), .Z(n118) );
  MUX2_X1 U718 ( .A(n118), .B(n115), .S(n606), .Z(n119) );
  MUX2_X1 U719 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U720 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U721 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n615), .Z(n121) );
  MUX2_X1 U722 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n611), .Z(n122) );
  MUX2_X1 U723 ( .A(n122), .B(n121), .S(n608), .Z(n123) );
  MUX2_X1 U724 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n617), .Z(n124) );
  MUX2_X1 U725 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n612), .Z(n125) );
  MUX2_X1 U726 ( .A(n125), .B(n124), .S(n608), .Z(n126) );
  MUX2_X1 U727 ( .A(n126), .B(n123), .S(n606), .Z(n127) );
  MUX2_X1 U728 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n617), .Z(n128) );
  MUX2_X1 U729 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n617), .Z(n129) );
  MUX2_X1 U730 ( .A(n129), .B(n128), .S(n609), .Z(n130) );
  MUX2_X1 U731 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n617), .Z(n131) );
  MUX2_X1 U732 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n617), .Z(n132) );
  MUX2_X1 U733 ( .A(n132), .B(n131), .S(n609), .Z(n133) );
  MUX2_X1 U734 ( .A(n133), .B(n130), .S(n606), .Z(n134) );
  MUX2_X1 U735 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U736 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n611), .Z(n136) );
  MUX2_X1 U737 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n617), .Z(n137) );
  MUX2_X1 U738 ( .A(n137), .B(n136), .S(n610), .Z(n138) );
  MUX2_X1 U739 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n614), .Z(n139) );
  MUX2_X1 U740 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n613), .Z(n140) );
  MUX2_X1 U741 ( .A(n140), .B(n139), .S(n608), .Z(n141) );
  MUX2_X1 U742 ( .A(n141), .B(n138), .S(n606), .Z(n142) );
  MUX2_X1 U743 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n617), .Z(n143) );
  MUX2_X1 U744 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n617), .Z(n144) );
  MUX2_X1 U745 ( .A(n144), .B(n143), .S(n609), .Z(n145) );
  MUX2_X1 U746 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n617), .Z(n146) );
  MUX2_X1 U747 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n617), .Z(n147) );
  MUX2_X1 U748 ( .A(n147), .B(n146), .S(n610), .Z(n148) );
  MUX2_X1 U749 ( .A(n148), .B(n145), .S(n606), .Z(n149) );
  MUX2_X1 U750 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U751 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U752 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n612), .Z(n151) );
  MUX2_X1 U753 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n616), .Z(n152) );
  MUX2_X1 U754 ( .A(n152), .B(n151), .S(N11), .Z(n153) );
  MUX2_X1 U755 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n613), .Z(n154) );
  MUX2_X1 U756 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n616), .Z(n155) );
  MUX2_X1 U757 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U758 ( .A(n156), .B(n153), .S(n607), .Z(n157) );
  MUX2_X1 U759 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n612), .Z(n158) );
  MUX2_X1 U760 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n611), .Z(n159) );
  MUX2_X1 U761 ( .A(n159), .B(n158), .S(n608), .Z(n160) );
  MUX2_X1 U762 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n612), .Z(n161) );
  MUX2_X1 U763 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n617), .Z(n162) );
  MUX2_X1 U764 ( .A(n162), .B(n161), .S(N11), .Z(n163) );
  MUX2_X1 U765 ( .A(n163), .B(n160), .S(n607), .Z(n164) );
  MUX2_X1 U766 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U767 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n611), .Z(n166) );
  MUX2_X1 U768 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n617), .Z(n167) );
  MUX2_X1 U769 ( .A(n167), .B(n166), .S(n610), .Z(n168) );
  MUX2_X1 U770 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n615), .Z(n169) );
  MUX2_X1 U771 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n617), .Z(n170) );
  MUX2_X1 U772 ( .A(n170), .B(n169), .S(n610), .Z(n171) );
  MUX2_X1 U773 ( .A(n171), .B(n168), .S(n607), .Z(n172) );
  MUX2_X1 U774 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n614), .Z(n173) );
  MUX2_X1 U775 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n614), .Z(n174) );
  MUX2_X1 U776 ( .A(n174), .B(n173), .S(n609), .Z(n175) );
  MUX2_X1 U777 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n614), .Z(n176) );
  MUX2_X1 U778 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n614), .Z(n177) );
  MUX2_X1 U779 ( .A(n177), .B(n176), .S(n609), .Z(n178) );
  MUX2_X1 U780 ( .A(n178), .B(n175), .S(n607), .Z(n179) );
  MUX2_X1 U781 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U782 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U783 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n614), .Z(n181) );
  MUX2_X1 U784 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n614), .Z(n182) );
  MUX2_X1 U785 ( .A(n182), .B(n181), .S(n609), .Z(n183) );
  MUX2_X1 U786 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n614), .Z(n184) );
  MUX2_X1 U787 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n614), .Z(n185) );
  MUX2_X1 U788 ( .A(n185), .B(n184), .S(n610), .Z(n186) );
  MUX2_X1 U789 ( .A(n186), .B(n183), .S(n607), .Z(n187) );
  MUX2_X1 U790 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n614), .Z(n188) );
  MUX2_X1 U791 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n614), .Z(n189) );
  MUX2_X1 U792 ( .A(n189), .B(n188), .S(N11), .Z(n190) );
  MUX2_X1 U793 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n614), .Z(n191) );
  MUX2_X1 U794 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n614), .Z(n192) );
  MUX2_X1 U795 ( .A(n192), .B(n191), .S(n608), .Z(n193) );
  MUX2_X1 U796 ( .A(n193), .B(n190), .S(n607), .Z(n194) );
  MUX2_X1 U797 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U798 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n615), .Z(n196) );
  MUX2_X1 U799 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n615), .Z(n197) );
  MUX2_X1 U800 ( .A(n197), .B(n196), .S(n608), .Z(n198) );
  MUX2_X1 U801 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n615), .Z(n199) );
  MUX2_X1 U802 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n615), .Z(n200) );
  MUX2_X1 U803 ( .A(n200), .B(n199), .S(N11), .Z(n201) );
  MUX2_X1 U804 ( .A(n201), .B(n198), .S(n607), .Z(n202) );
  MUX2_X1 U805 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n615), .Z(n203) );
  MUX2_X1 U806 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n615), .Z(n204) );
  MUX2_X1 U807 ( .A(n204), .B(n203), .S(n608), .Z(n205) );
  MUX2_X1 U808 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n615), .Z(n206) );
  MUX2_X1 U809 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n615), .Z(n207) );
  MUX2_X1 U810 ( .A(n207), .B(n206), .S(n610), .Z(n208) );
  MUX2_X1 U811 ( .A(n208), .B(n205), .S(n607), .Z(n209) );
  MUX2_X1 U812 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U813 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U814 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n615), .Z(n211) );
  MUX2_X1 U815 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n615), .Z(n212) );
  MUX2_X1 U816 ( .A(n212), .B(n211), .S(n608), .Z(n213) );
  MUX2_X1 U817 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n615), .Z(n214) );
  MUX2_X1 U818 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n615), .Z(n215) );
  MUX2_X1 U819 ( .A(n215), .B(n214), .S(n608), .Z(n216) );
  MUX2_X1 U820 ( .A(n216), .B(n213), .S(n607), .Z(n217) );
  MUX2_X1 U821 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n616), .Z(n218) );
  MUX2_X1 U822 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n616), .Z(n219) );
  MUX2_X1 U823 ( .A(n219), .B(n218), .S(n608), .Z(n220) );
  MUX2_X1 U824 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n616), .Z(n221) );
  MUX2_X1 U825 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n616), .Z(n222) );
  MUX2_X1 U826 ( .A(n222), .B(n221), .S(n609), .Z(n223) );
  MUX2_X1 U827 ( .A(n223), .B(n220), .S(n607), .Z(n224) );
  MUX2_X1 U828 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U829 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n616), .Z(n226) );
  MUX2_X1 U830 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n616), .Z(n227) );
  MUX2_X1 U831 ( .A(n227), .B(n226), .S(n608), .Z(n228) );
  MUX2_X1 U832 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n616), .Z(n229) );
  MUX2_X1 U833 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n616), .Z(n595) );
  MUX2_X1 U834 ( .A(n595), .B(n229), .S(n610), .Z(n596) );
  MUX2_X1 U835 ( .A(n596), .B(n228), .S(n607), .Z(n597) );
  MUX2_X1 U836 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n616), .Z(n598) );
  MUX2_X1 U837 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n616), .Z(n599) );
  MUX2_X1 U838 ( .A(n599), .B(n598), .S(n608), .Z(n600) );
  MUX2_X1 U839 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n616), .Z(n601) );
  MUX2_X1 U840 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n616), .Z(n602) );
  MUX2_X1 U841 ( .A(n602), .B(n601), .S(n608), .Z(n603) );
  MUX2_X1 U842 ( .A(n603), .B(n600), .S(n607), .Z(n604) );
  MUX2_X1 U843 ( .A(n604), .B(n597), .S(N13), .Z(n605) );
  MUX2_X1 U844 ( .A(n605), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U845 ( .A(N11), .Z(n608) );
  CLKBUF_X1 U846 ( .A(n617), .Z(n611) );
  INV_X1 U847 ( .A(N10), .ZN(n618) );
  INV_X1 U848 ( .A(N11), .ZN(n619) );
  INV_X1 U849 ( .A(data_in[0]), .ZN(n620) );
  INV_X1 U850 ( .A(data_in[1]), .ZN(n621) );
  INV_X1 U851 ( .A(data_in[2]), .ZN(n622) );
  INV_X1 U852 ( .A(data_in[3]), .ZN(n623) );
  INV_X1 U853 ( .A(data_in[4]), .ZN(n624) );
  INV_X1 U854 ( .A(data_in[5]), .ZN(n625) );
  INV_X1 U855 ( .A(data_in[6]), .ZN(n626) );
  INV_X1 U856 ( .A(data_in[7]), .ZN(n627) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_16 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n629), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n630), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n631), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n632), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n633), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n634), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n635), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n636), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n637), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n638), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n639), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n640), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n641), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n642), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n643), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n644), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n645), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n646), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n647), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n648), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n649), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n650), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n651), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n652), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n653), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n654), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n655), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n656), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n657), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n658), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n659), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n660), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n661), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n662), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n663), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n664), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n665), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n666), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n667), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n668), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n669), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n670), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n671), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n672), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n673), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n674), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n675), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n676), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n677), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n678), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n679), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n680), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n681), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n682), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n683), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n684), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n685), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n686), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n687), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n688), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n689), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n690), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n691), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n692), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n693), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n694), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n695), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n696), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n697), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n698), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n699), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n700), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n701), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n702), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n703), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n704), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n705), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n706), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n707), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n708), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n709), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n710), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n711), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n712), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n713), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n714), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n715), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n716), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n717), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n718), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n719), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n720), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n721), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n722), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n723), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n724), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n725), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n726), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n727), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n728), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n729), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n730), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n731), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n732), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n733), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n734), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n735), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n736), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n737), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n738), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n739), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n740), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n741), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n742), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n743), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n744), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n745), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n746), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n747), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n748), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n749), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n750), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n751), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n752), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n753), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n754), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n755), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n756), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n757), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n758), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n759), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n760), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n761), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n762), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n763), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n764), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n765), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n766), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n767), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n768), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n769), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n770), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n771), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n772), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n773), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n774), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n775), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n776), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n777), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n778), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n779), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n780), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n781), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n782), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n783), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n784), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n785), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n786), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n787), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n788), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n789), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n790), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n791), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n792), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n793), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n794), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n795), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n796), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n797), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n798), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n799), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n800), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n801), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n802), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n803), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n804), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n805), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n806), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n807), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n808), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n809), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n810), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n811), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n812), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n813), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n814), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n815), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n816), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n817), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n818), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n819), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n820), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n848), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n849), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n850), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n851), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n852), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n853), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n854), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n855), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n856), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n857), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n858), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n859), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n860), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n861), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n862), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n863), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n864), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n865), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n866), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n867), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n868), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n869), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n870), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n871), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n872), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n873), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n874), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n875), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n876), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n877), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n878), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n879), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n880), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n881), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n882), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n883), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n884), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n885), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n886), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n887), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n888), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n889), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n890), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n891), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n892), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n893), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n894), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n895), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n896), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n897), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n898), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n899), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n900), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n901), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n902), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n903), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n904), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n905), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n906), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n907), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n908), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n909), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n910), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n911), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(n618), .Z(n617) );
  BUF_X1 U5 ( .A(n618), .Z(n614) );
  BUF_X1 U6 ( .A(N10), .Z(n615) );
  BUF_X1 U7 ( .A(n618), .Z(n616) );
  BUF_X1 U8 ( .A(n618), .Z(n613) );
  BUF_X1 U9 ( .A(N11), .Z(n611) );
  BUF_X1 U10 ( .A(N11), .Z(n612) );
  BUF_X1 U11 ( .A(N10), .Z(n618) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1203) );
  NOR3_X1 U13 ( .A1(N11), .A2(N12), .A3(n619), .ZN(n1192) );
  NOR3_X1 U14 ( .A1(N10), .A2(N12), .A3(n620), .ZN(n1182) );
  NOR3_X1 U15 ( .A1(n619), .A2(N12), .A3(n620), .ZN(n1172) );
  INV_X1 U16 ( .A(n1129), .ZN(n844) );
  INV_X1 U17 ( .A(n1119), .ZN(n843) );
  INV_X1 U18 ( .A(n1110), .ZN(n842) );
  INV_X1 U19 ( .A(n1101), .ZN(n841) );
  INV_X1 U20 ( .A(n1056), .ZN(n836) );
  INV_X1 U21 ( .A(n1046), .ZN(n835) );
  INV_X1 U22 ( .A(n1037), .ZN(n834) );
  INV_X1 U23 ( .A(n1028), .ZN(n833) );
  INV_X1 U24 ( .A(n983), .ZN(n828) );
  INV_X1 U25 ( .A(n973), .ZN(n827) );
  INV_X1 U26 ( .A(n964), .ZN(n826) );
  INV_X1 U27 ( .A(n955), .ZN(n825) );
  INV_X1 U28 ( .A(n946), .ZN(n824) );
  INV_X1 U29 ( .A(n937), .ZN(n823) );
  INV_X1 U30 ( .A(n928), .ZN(n822) );
  INV_X1 U31 ( .A(n919), .ZN(n821) );
  INV_X1 U32 ( .A(n1092), .ZN(n840) );
  INV_X1 U33 ( .A(n1083), .ZN(n839) );
  INV_X1 U34 ( .A(n1074), .ZN(n838) );
  INV_X1 U35 ( .A(n1065), .ZN(n837) );
  INV_X1 U36 ( .A(n1019), .ZN(n832) );
  INV_X1 U37 ( .A(n1010), .ZN(n831) );
  INV_X1 U38 ( .A(n1001), .ZN(n830) );
  INV_X1 U39 ( .A(n992), .ZN(n829) );
  BUF_X1 U40 ( .A(N12), .Z(n608) );
  BUF_X1 U41 ( .A(N12), .Z(n609) );
  INV_X1 U42 ( .A(N13), .ZN(n846) );
  AND3_X1 U43 ( .A1(n619), .A2(n620), .A3(N12), .ZN(n1162) );
  AND3_X1 U44 ( .A1(N10), .A2(n620), .A3(N12), .ZN(n1152) );
  AND3_X1 U45 ( .A1(N11), .A2(n619), .A3(N12), .ZN(n1142) );
  AND3_X1 U46 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1132) );
  INV_X1 U47 ( .A(N14), .ZN(n847) );
  NAND2_X1 U48 ( .A1(n1192), .A2(n1202), .ZN(n1201) );
  NAND2_X1 U49 ( .A1(n1182), .A2(n1202), .ZN(n1191) );
  NAND2_X1 U50 ( .A1(n1172), .A2(n1202), .ZN(n1181) );
  NAND2_X1 U51 ( .A1(n1162), .A2(n1202), .ZN(n1171) );
  NAND2_X1 U52 ( .A1(n1152), .A2(n1202), .ZN(n1161) );
  NAND2_X1 U53 ( .A1(n1142), .A2(n1202), .ZN(n1151) );
  NAND2_X1 U54 ( .A1(n1132), .A2(n1202), .ZN(n1141) );
  NAND2_X1 U55 ( .A1(n1203), .A2(n1202), .ZN(n1212) );
  NAND2_X1 U56 ( .A1(n1121), .A2(n1203), .ZN(n1129) );
  NAND2_X1 U57 ( .A1(n1121), .A2(n1192), .ZN(n1119) );
  NAND2_X1 U58 ( .A1(n1121), .A2(n1182), .ZN(n1110) );
  NAND2_X1 U59 ( .A1(n1121), .A2(n1172), .ZN(n1101) );
  NAND2_X1 U60 ( .A1(n1048), .A2(n1203), .ZN(n1056) );
  NAND2_X1 U61 ( .A1(n1048), .A2(n1192), .ZN(n1046) );
  NAND2_X1 U62 ( .A1(n1048), .A2(n1182), .ZN(n1037) );
  NAND2_X1 U63 ( .A1(n1048), .A2(n1172), .ZN(n1028) );
  NAND2_X1 U64 ( .A1(n975), .A2(n1203), .ZN(n983) );
  NAND2_X1 U65 ( .A1(n975), .A2(n1192), .ZN(n973) );
  NAND2_X1 U66 ( .A1(n975), .A2(n1182), .ZN(n964) );
  NAND2_X1 U67 ( .A1(n975), .A2(n1172), .ZN(n955) );
  NAND2_X1 U68 ( .A1(n1121), .A2(n1162), .ZN(n1092) );
  NAND2_X1 U69 ( .A1(n1121), .A2(n1152), .ZN(n1083) );
  NAND2_X1 U70 ( .A1(n1121), .A2(n1142), .ZN(n1074) );
  NAND2_X1 U71 ( .A1(n1121), .A2(n1132), .ZN(n1065) );
  NAND2_X1 U72 ( .A1(n1048), .A2(n1162), .ZN(n1019) );
  NAND2_X1 U73 ( .A1(n1048), .A2(n1152), .ZN(n1010) );
  NAND2_X1 U74 ( .A1(n1048), .A2(n1142), .ZN(n1001) );
  NAND2_X1 U75 ( .A1(n1048), .A2(n1132), .ZN(n992) );
  NAND2_X1 U76 ( .A1(n975), .A2(n1162), .ZN(n946) );
  NAND2_X1 U77 ( .A1(n975), .A2(n1152), .ZN(n937) );
  NAND2_X1 U78 ( .A1(n975), .A2(n1142), .ZN(n928) );
  NAND2_X1 U79 ( .A1(n975), .A2(n1132), .ZN(n919) );
  AND3_X1 U80 ( .A1(n846), .A2(n847), .A3(n1131), .ZN(n1202) );
  AND3_X1 U81 ( .A1(N13), .A2(n1131), .A3(N14), .ZN(n975) );
  AND3_X1 U82 ( .A1(n1131), .A2(n847), .A3(N13), .ZN(n1121) );
  AND3_X1 U83 ( .A1(n1131), .A2(n846), .A3(N14), .ZN(n1048) );
  NOR2_X1 U84 ( .A1(n845), .A2(addr[5]), .ZN(n1131) );
  INV_X1 U85 ( .A(wr_en), .ZN(n845) );
  OAI21_X1 U86 ( .B1(n621), .B2(n1171), .A(n1170), .ZN(n879) );
  NAND2_X1 U87 ( .A1(\mem[4][0] ), .A2(n1171), .ZN(n1170) );
  OAI21_X1 U88 ( .B1(n622), .B2(n1171), .A(n1169), .ZN(n878) );
  NAND2_X1 U89 ( .A1(\mem[4][1] ), .A2(n1171), .ZN(n1169) );
  OAI21_X1 U90 ( .B1(n623), .B2(n1171), .A(n1168), .ZN(n877) );
  NAND2_X1 U91 ( .A1(\mem[4][2] ), .A2(n1171), .ZN(n1168) );
  OAI21_X1 U92 ( .B1(n624), .B2(n1171), .A(n1167), .ZN(n876) );
  NAND2_X1 U93 ( .A1(\mem[4][3] ), .A2(n1171), .ZN(n1167) );
  OAI21_X1 U94 ( .B1(n625), .B2(n1171), .A(n1166), .ZN(n875) );
  NAND2_X1 U95 ( .A1(\mem[4][4] ), .A2(n1171), .ZN(n1166) );
  OAI21_X1 U96 ( .B1(n626), .B2(n1171), .A(n1165), .ZN(n874) );
  NAND2_X1 U97 ( .A1(\mem[4][5] ), .A2(n1171), .ZN(n1165) );
  OAI21_X1 U98 ( .B1(n627), .B2(n1171), .A(n1164), .ZN(n873) );
  NAND2_X1 U99 ( .A1(\mem[4][6] ), .A2(n1171), .ZN(n1164) );
  OAI21_X1 U100 ( .B1(n628), .B2(n1171), .A(n1163), .ZN(n872) );
  NAND2_X1 U101 ( .A1(\mem[4][7] ), .A2(n1171), .ZN(n1163) );
  OAI21_X1 U102 ( .B1(n621), .B2(n1151), .A(n1150), .ZN(n863) );
  NAND2_X1 U103 ( .A1(\mem[6][0] ), .A2(n1151), .ZN(n1150) );
  OAI21_X1 U104 ( .B1(n622), .B2(n1151), .A(n1149), .ZN(n862) );
  NAND2_X1 U105 ( .A1(\mem[6][1] ), .A2(n1151), .ZN(n1149) );
  OAI21_X1 U106 ( .B1(n623), .B2(n1151), .A(n1148), .ZN(n861) );
  NAND2_X1 U107 ( .A1(\mem[6][2] ), .A2(n1151), .ZN(n1148) );
  OAI21_X1 U108 ( .B1(n624), .B2(n1151), .A(n1147), .ZN(n860) );
  NAND2_X1 U109 ( .A1(\mem[6][3] ), .A2(n1151), .ZN(n1147) );
  OAI21_X1 U110 ( .B1(n625), .B2(n1151), .A(n1146), .ZN(n859) );
  NAND2_X1 U111 ( .A1(\mem[6][4] ), .A2(n1151), .ZN(n1146) );
  OAI21_X1 U112 ( .B1(n626), .B2(n1151), .A(n1145), .ZN(n858) );
  NAND2_X1 U113 ( .A1(\mem[6][5] ), .A2(n1151), .ZN(n1145) );
  OAI21_X1 U114 ( .B1(n627), .B2(n1151), .A(n1144), .ZN(n857) );
  NAND2_X1 U115 ( .A1(\mem[6][6] ), .A2(n1151), .ZN(n1144) );
  OAI21_X1 U116 ( .B1(n628), .B2(n1151), .A(n1143), .ZN(n856) );
  NAND2_X1 U117 ( .A1(\mem[6][7] ), .A2(n1151), .ZN(n1143) );
  OAI21_X1 U118 ( .B1(n621), .B2(n1141), .A(n1140), .ZN(n855) );
  NAND2_X1 U119 ( .A1(\mem[7][0] ), .A2(n1141), .ZN(n1140) );
  OAI21_X1 U120 ( .B1(n622), .B2(n1141), .A(n1139), .ZN(n854) );
  NAND2_X1 U121 ( .A1(\mem[7][1] ), .A2(n1141), .ZN(n1139) );
  OAI21_X1 U122 ( .B1(n623), .B2(n1141), .A(n1138), .ZN(n853) );
  NAND2_X1 U123 ( .A1(\mem[7][2] ), .A2(n1141), .ZN(n1138) );
  OAI21_X1 U124 ( .B1(n624), .B2(n1141), .A(n1137), .ZN(n852) );
  NAND2_X1 U125 ( .A1(\mem[7][3] ), .A2(n1141), .ZN(n1137) );
  OAI21_X1 U126 ( .B1(n625), .B2(n1141), .A(n1136), .ZN(n851) );
  NAND2_X1 U127 ( .A1(\mem[7][4] ), .A2(n1141), .ZN(n1136) );
  OAI21_X1 U128 ( .B1(n626), .B2(n1141), .A(n1135), .ZN(n850) );
  NAND2_X1 U129 ( .A1(\mem[7][5] ), .A2(n1141), .ZN(n1135) );
  OAI21_X1 U130 ( .B1(n627), .B2(n1141), .A(n1134), .ZN(n849) );
  NAND2_X1 U131 ( .A1(\mem[7][6] ), .A2(n1141), .ZN(n1134) );
  OAI21_X1 U132 ( .B1(n628), .B2(n1141), .A(n1133), .ZN(n848) );
  NAND2_X1 U133 ( .A1(\mem[7][7] ), .A2(n1141), .ZN(n1133) );
  OAI21_X1 U134 ( .B1(n621), .B2(n1201), .A(n1200), .ZN(n903) );
  NAND2_X1 U135 ( .A1(\mem[1][0] ), .A2(n1201), .ZN(n1200) );
  OAI21_X1 U136 ( .B1(n622), .B2(n1201), .A(n1199), .ZN(n902) );
  NAND2_X1 U137 ( .A1(\mem[1][1] ), .A2(n1201), .ZN(n1199) );
  OAI21_X1 U138 ( .B1(n623), .B2(n1201), .A(n1198), .ZN(n901) );
  NAND2_X1 U139 ( .A1(\mem[1][2] ), .A2(n1201), .ZN(n1198) );
  OAI21_X1 U140 ( .B1(n624), .B2(n1201), .A(n1197), .ZN(n900) );
  NAND2_X1 U141 ( .A1(\mem[1][3] ), .A2(n1201), .ZN(n1197) );
  OAI21_X1 U142 ( .B1(n625), .B2(n1201), .A(n1196), .ZN(n899) );
  NAND2_X1 U143 ( .A1(\mem[1][4] ), .A2(n1201), .ZN(n1196) );
  OAI21_X1 U144 ( .B1(n626), .B2(n1201), .A(n1195), .ZN(n898) );
  NAND2_X1 U145 ( .A1(\mem[1][5] ), .A2(n1201), .ZN(n1195) );
  OAI21_X1 U146 ( .B1(n627), .B2(n1201), .A(n1194), .ZN(n897) );
  NAND2_X1 U147 ( .A1(\mem[1][6] ), .A2(n1201), .ZN(n1194) );
  OAI21_X1 U148 ( .B1(n628), .B2(n1201), .A(n1193), .ZN(n896) );
  NAND2_X1 U149 ( .A1(\mem[1][7] ), .A2(n1201), .ZN(n1193) );
  OAI21_X1 U150 ( .B1(n621), .B2(n1191), .A(n1190), .ZN(n895) );
  NAND2_X1 U151 ( .A1(\mem[2][0] ), .A2(n1191), .ZN(n1190) );
  OAI21_X1 U152 ( .B1(n622), .B2(n1191), .A(n1189), .ZN(n894) );
  NAND2_X1 U153 ( .A1(\mem[2][1] ), .A2(n1191), .ZN(n1189) );
  OAI21_X1 U154 ( .B1(n623), .B2(n1191), .A(n1188), .ZN(n893) );
  NAND2_X1 U155 ( .A1(\mem[2][2] ), .A2(n1191), .ZN(n1188) );
  OAI21_X1 U156 ( .B1(n624), .B2(n1191), .A(n1187), .ZN(n892) );
  NAND2_X1 U157 ( .A1(\mem[2][3] ), .A2(n1191), .ZN(n1187) );
  OAI21_X1 U158 ( .B1(n625), .B2(n1191), .A(n1186), .ZN(n891) );
  NAND2_X1 U159 ( .A1(\mem[2][4] ), .A2(n1191), .ZN(n1186) );
  OAI21_X1 U160 ( .B1(n626), .B2(n1191), .A(n1185), .ZN(n890) );
  NAND2_X1 U161 ( .A1(\mem[2][5] ), .A2(n1191), .ZN(n1185) );
  OAI21_X1 U162 ( .B1(n627), .B2(n1191), .A(n1184), .ZN(n889) );
  NAND2_X1 U163 ( .A1(\mem[2][6] ), .A2(n1191), .ZN(n1184) );
  OAI21_X1 U164 ( .B1(n628), .B2(n1191), .A(n1183), .ZN(n888) );
  NAND2_X1 U165 ( .A1(\mem[2][7] ), .A2(n1191), .ZN(n1183) );
  OAI21_X1 U166 ( .B1(n621), .B2(n1181), .A(n1180), .ZN(n887) );
  NAND2_X1 U167 ( .A1(\mem[3][0] ), .A2(n1181), .ZN(n1180) );
  OAI21_X1 U168 ( .B1(n622), .B2(n1181), .A(n1179), .ZN(n886) );
  NAND2_X1 U169 ( .A1(\mem[3][1] ), .A2(n1181), .ZN(n1179) );
  OAI21_X1 U170 ( .B1(n623), .B2(n1181), .A(n1178), .ZN(n885) );
  NAND2_X1 U171 ( .A1(\mem[3][2] ), .A2(n1181), .ZN(n1178) );
  OAI21_X1 U172 ( .B1(n624), .B2(n1181), .A(n1177), .ZN(n884) );
  NAND2_X1 U173 ( .A1(\mem[3][3] ), .A2(n1181), .ZN(n1177) );
  OAI21_X1 U174 ( .B1(n625), .B2(n1181), .A(n1176), .ZN(n883) );
  NAND2_X1 U175 ( .A1(\mem[3][4] ), .A2(n1181), .ZN(n1176) );
  OAI21_X1 U176 ( .B1(n626), .B2(n1181), .A(n1175), .ZN(n882) );
  NAND2_X1 U177 ( .A1(\mem[3][5] ), .A2(n1181), .ZN(n1175) );
  OAI21_X1 U178 ( .B1(n627), .B2(n1181), .A(n1174), .ZN(n881) );
  NAND2_X1 U179 ( .A1(\mem[3][6] ), .A2(n1181), .ZN(n1174) );
  OAI21_X1 U180 ( .B1(n628), .B2(n1181), .A(n1173), .ZN(n880) );
  NAND2_X1 U181 ( .A1(\mem[3][7] ), .A2(n1181), .ZN(n1173) );
  OAI21_X1 U182 ( .B1(n621), .B2(n1161), .A(n1160), .ZN(n871) );
  NAND2_X1 U183 ( .A1(\mem[5][0] ), .A2(n1161), .ZN(n1160) );
  OAI21_X1 U184 ( .B1(n622), .B2(n1161), .A(n1159), .ZN(n870) );
  NAND2_X1 U185 ( .A1(\mem[5][1] ), .A2(n1161), .ZN(n1159) );
  OAI21_X1 U186 ( .B1(n623), .B2(n1161), .A(n1158), .ZN(n869) );
  NAND2_X1 U187 ( .A1(\mem[5][2] ), .A2(n1161), .ZN(n1158) );
  OAI21_X1 U188 ( .B1(n624), .B2(n1161), .A(n1157), .ZN(n868) );
  NAND2_X1 U189 ( .A1(\mem[5][3] ), .A2(n1161), .ZN(n1157) );
  OAI21_X1 U190 ( .B1(n625), .B2(n1161), .A(n1156), .ZN(n867) );
  NAND2_X1 U191 ( .A1(\mem[5][4] ), .A2(n1161), .ZN(n1156) );
  OAI21_X1 U192 ( .B1(n626), .B2(n1161), .A(n1155), .ZN(n866) );
  NAND2_X1 U193 ( .A1(\mem[5][5] ), .A2(n1161), .ZN(n1155) );
  OAI21_X1 U194 ( .B1(n627), .B2(n1161), .A(n1154), .ZN(n865) );
  NAND2_X1 U195 ( .A1(\mem[5][6] ), .A2(n1161), .ZN(n1154) );
  OAI21_X1 U196 ( .B1(n628), .B2(n1161), .A(n1153), .ZN(n864) );
  NAND2_X1 U197 ( .A1(\mem[5][7] ), .A2(n1161), .ZN(n1153) );
  OAI21_X1 U198 ( .B1(n1212), .B2(n621), .A(n1211), .ZN(n911) );
  NAND2_X1 U199 ( .A1(\mem[0][0] ), .A2(n1212), .ZN(n1211) );
  OAI21_X1 U200 ( .B1(n1212), .B2(n622), .A(n1210), .ZN(n910) );
  NAND2_X1 U201 ( .A1(\mem[0][1] ), .A2(n1212), .ZN(n1210) );
  OAI21_X1 U202 ( .B1(n1212), .B2(n623), .A(n1209), .ZN(n909) );
  NAND2_X1 U203 ( .A1(\mem[0][2] ), .A2(n1212), .ZN(n1209) );
  OAI21_X1 U204 ( .B1(n1212), .B2(n624), .A(n1208), .ZN(n908) );
  NAND2_X1 U205 ( .A1(\mem[0][3] ), .A2(n1212), .ZN(n1208) );
  OAI21_X1 U206 ( .B1(n1212), .B2(n625), .A(n1207), .ZN(n907) );
  NAND2_X1 U207 ( .A1(\mem[0][4] ), .A2(n1212), .ZN(n1207) );
  OAI21_X1 U208 ( .B1(n1212), .B2(n626), .A(n1206), .ZN(n906) );
  NAND2_X1 U209 ( .A1(\mem[0][5] ), .A2(n1212), .ZN(n1206) );
  OAI21_X1 U210 ( .B1(n1212), .B2(n627), .A(n1205), .ZN(n905) );
  NAND2_X1 U211 ( .A1(\mem[0][6] ), .A2(n1212), .ZN(n1205) );
  OAI21_X1 U212 ( .B1(n1212), .B2(n628), .A(n1204), .ZN(n904) );
  NAND2_X1 U213 ( .A1(\mem[0][7] ), .A2(n1212), .ZN(n1204) );
  INV_X1 U214 ( .A(n1130), .ZN(n820) );
  AOI22_X1 U215 ( .A1(data_in[0]), .A2(n844), .B1(n1129), .B2(\mem[8][0] ), 
        .ZN(n1130) );
  INV_X1 U216 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U217 ( .A1(data_in[1]), .A2(n844), .B1(n1129), .B2(\mem[8][1] ), 
        .ZN(n1128) );
  INV_X1 U218 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U219 ( .A1(data_in[2]), .A2(n844), .B1(n1129), .B2(\mem[8][2] ), 
        .ZN(n1127) );
  INV_X1 U220 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U221 ( .A1(data_in[3]), .A2(n844), .B1(n1129), .B2(\mem[8][3] ), 
        .ZN(n1126) );
  INV_X1 U222 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U223 ( .A1(data_in[4]), .A2(n844), .B1(n1129), .B2(\mem[8][4] ), 
        .ZN(n1125) );
  INV_X1 U224 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U225 ( .A1(data_in[5]), .A2(n844), .B1(n1129), .B2(\mem[8][5] ), 
        .ZN(n1124) );
  INV_X1 U226 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U227 ( .A1(data_in[6]), .A2(n844), .B1(n1129), .B2(\mem[8][6] ), 
        .ZN(n1123) );
  INV_X1 U228 ( .A(n1122), .ZN(n813) );
  AOI22_X1 U229 ( .A1(data_in[7]), .A2(n844), .B1(n1129), .B2(\mem[8][7] ), 
        .ZN(n1122) );
  INV_X1 U230 ( .A(n1120), .ZN(n812) );
  AOI22_X1 U231 ( .A1(data_in[0]), .A2(n843), .B1(n1119), .B2(\mem[9][0] ), 
        .ZN(n1120) );
  INV_X1 U232 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U233 ( .A1(data_in[1]), .A2(n843), .B1(n1119), .B2(\mem[9][1] ), 
        .ZN(n1118) );
  INV_X1 U234 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U235 ( .A1(data_in[2]), .A2(n843), .B1(n1119), .B2(\mem[9][2] ), 
        .ZN(n1117) );
  INV_X1 U236 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U237 ( .A1(data_in[3]), .A2(n843), .B1(n1119), .B2(\mem[9][3] ), 
        .ZN(n1116) );
  INV_X1 U238 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U239 ( .A1(data_in[4]), .A2(n843), .B1(n1119), .B2(\mem[9][4] ), 
        .ZN(n1115) );
  INV_X1 U240 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U241 ( .A1(data_in[5]), .A2(n843), .B1(n1119), .B2(\mem[9][5] ), 
        .ZN(n1114) );
  INV_X1 U242 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U243 ( .A1(data_in[6]), .A2(n843), .B1(n1119), .B2(\mem[9][6] ), 
        .ZN(n1113) );
  INV_X1 U244 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U245 ( .A1(data_in[7]), .A2(n843), .B1(n1119), .B2(\mem[9][7] ), 
        .ZN(n1112) );
  INV_X1 U246 ( .A(n1111), .ZN(n804) );
  AOI22_X1 U247 ( .A1(data_in[0]), .A2(n842), .B1(n1110), .B2(\mem[10][0] ), 
        .ZN(n1111) );
  INV_X1 U248 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U249 ( .A1(data_in[1]), .A2(n842), .B1(n1110), .B2(\mem[10][1] ), 
        .ZN(n1109) );
  INV_X1 U250 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U251 ( .A1(data_in[2]), .A2(n842), .B1(n1110), .B2(\mem[10][2] ), 
        .ZN(n1108) );
  INV_X1 U252 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U253 ( .A1(data_in[3]), .A2(n842), .B1(n1110), .B2(\mem[10][3] ), 
        .ZN(n1107) );
  INV_X1 U254 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U255 ( .A1(data_in[4]), .A2(n842), .B1(n1110), .B2(\mem[10][4] ), 
        .ZN(n1106) );
  INV_X1 U256 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U257 ( .A1(data_in[5]), .A2(n842), .B1(n1110), .B2(\mem[10][5] ), 
        .ZN(n1105) );
  INV_X1 U258 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U259 ( .A1(data_in[6]), .A2(n842), .B1(n1110), .B2(\mem[10][6] ), 
        .ZN(n1104) );
  INV_X1 U260 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U261 ( .A1(data_in[7]), .A2(n842), .B1(n1110), .B2(\mem[10][7] ), 
        .ZN(n1103) );
  INV_X1 U262 ( .A(n1102), .ZN(n796) );
  AOI22_X1 U263 ( .A1(data_in[0]), .A2(n841), .B1(n1101), .B2(\mem[11][0] ), 
        .ZN(n1102) );
  INV_X1 U264 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U265 ( .A1(data_in[1]), .A2(n841), .B1(n1101), .B2(\mem[11][1] ), 
        .ZN(n1100) );
  INV_X1 U266 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U267 ( .A1(data_in[2]), .A2(n841), .B1(n1101), .B2(\mem[11][2] ), 
        .ZN(n1099) );
  INV_X1 U268 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U269 ( .A1(data_in[3]), .A2(n841), .B1(n1101), .B2(\mem[11][3] ), 
        .ZN(n1098) );
  INV_X1 U270 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U271 ( .A1(data_in[4]), .A2(n841), .B1(n1101), .B2(\mem[11][4] ), 
        .ZN(n1097) );
  INV_X1 U272 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U273 ( .A1(data_in[5]), .A2(n841), .B1(n1101), .B2(\mem[11][5] ), 
        .ZN(n1096) );
  INV_X1 U274 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U275 ( .A1(data_in[6]), .A2(n841), .B1(n1101), .B2(\mem[11][6] ), 
        .ZN(n1095) );
  INV_X1 U276 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U277 ( .A1(data_in[7]), .A2(n841), .B1(n1101), .B2(\mem[11][7] ), 
        .ZN(n1094) );
  INV_X1 U278 ( .A(n1093), .ZN(n788) );
  AOI22_X1 U279 ( .A1(data_in[0]), .A2(n840), .B1(n1092), .B2(\mem[12][0] ), 
        .ZN(n1093) );
  INV_X1 U280 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U281 ( .A1(data_in[1]), .A2(n840), .B1(n1092), .B2(\mem[12][1] ), 
        .ZN(n1091) );
  INV_X1 U282 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U283 ( .A1(data_in[2]), .A2(n840), .B1(n1092), .B2(\mem[12][2] ), 
        .ZN(n1090) );
  INV_X1 U284 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U285 ( .A1(data_in[3]), .A2(n840), .B1(n1092), .B2(\mem[12][3] ), 
        .ZN(n1089) );
  INV_X1 U286 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U287 ( .A1(data_in[4]), .A2(n840), .B1(n1092), .B2(\mem[12][4] ), 
        .ZN(n1088) );
  INV_X1 U288 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U289 ( .A1(data_in[5]), .A2(n840), .B1(n1092), .B2(\mem[12][5] ), 
        .ZN(n1087) );
  INV_X1 U290 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U291 ( .A1(data_in[6]), .A2(n840), .B1(n1092), .B2(\mem[12][6] ), 
        .ZN(n1086) );
  INV_X1 U292 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U293 ( .A1(data_in[7]), .A2(n840), .B1(n1092), .B2(\mem[12][7] ), 
        .ZN(n1085) );
  INV_X1 U294 ( .A(n1084), .ZN(n780) );
  AOI22_X1 U295 ( .A1(data_in[0]), .A2(n839), .B1(n1083), .B2(\mem[13][0] ), 
        .ZN(n1084) );
  INV_X1 U296 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U297 ( .A1(data_in[1]), .A2(n839), .B1(n1083), .B2(\mem[13][1] ), 
        .ZN(n1082) );
  INV_X1 U298 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U299 ( .A1(data_in[2]), .A2(n839), .B1(n1083), .B2(\mem[13][2] ), 
        .ZN(n1081) );
  INV_X1 U300 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U301 ( .A1(data_in[3]), .A2(n839), .B1(n1083), .B2(\mem[13][3] ), 
        .ZN(n1080) );
  INV_X1 U302 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U303 ( .A1(data_in[4]), .A2(n839), .B1(n1083), .B2(\mem[13][4] ), 
        .ZN(n1079) );
  INV_X1 U304 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U305 ( .A1(data_in[5]), .A2(n839), .B1(n1083), .B2(\mem[13][5] ), 
        .ZN(n1078) );
  INV_X1 U306 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U307 ( .A1(data_in[6]), .A2(n839), .B1(n1083), .B2(\mem[13][6] ), 
        .ZN(n1077) );
  INV_X1 U308 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U309 ( .A1(data_in[7]), .A2(n839), .B1(n1083), .B2(\mem[13][7] ), 
        .ZN(n1076) );
  INV_X1 U310 ( .A(n1075), .ZN(n772) );
  AOI22_X1 U311 ( .A1(data_in[0]), .A2(n838), .B1(n1074), .B2(\mem[14][0] ), 
        .ZN(n1075) );
  INV_X1 U312 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U313 ( .A1(data_in[1]), .A2(n838), .B1(n1074), .B2(\mem[14][1] ), 
        .ZN(n1073) );
  INV_X1 U314 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U315 ( .A1(data_in[2]), .A2(n838), .B1(n1074), .B2(\mem[14][2] ), 
        .ZN(n1072) );
  INV_X1 U316 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U317 ( .A1(data_in[3]), .A2(n838), .B1(n1074), .B2(\mem[14][3] ), 
        .ZN(n1071) );
  INV_X1 U318 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U319 ( .A1(data_in[4]), .A2(n838), .B1(n1074), .B2(\mem[14][4] ), 
        .ZN(n1070) );
  INV_X1 U320 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U321 ( .A1(data_in[5]), .A2(n838), .B1(n1074), .B2(\mem[14][5] ), 
        .ZN(n1069) );
  INV_X1 U322 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U323 ( .A1(data_in[6]), .A2(n838), .B1(n1074), .B2(\mem[14][6] ), 
        .ZN(n1068) );
  INV_X1 U324 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U325 ( .A1(data_in[7]), .A2(n838), .B1(n1074), .B2(\mem[14][7] ), 
        .ZN(n1067) );
  INV_X1 U326 ( .A(n1066), .ZN(n764) );
  AOI22_X1 U327 ( .A1(data_in[0]), .A2(n837), .B1(n1065), .B2(\mem[15][0] ), 
        .ZN(n1066) );
  INV_X1 U328 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U329 ( .A1(data_in[1]), .A2(n837), .B1(n1065), .B2(\mem[15][1] ), 
        .ZN(n1064) );
  INV_X1 U330 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U331 ( .A1(data_in[2]), .A2(n837), .B1(n1065), .B2(\mem[15][2] ), 
        .ZN(n1063) );
  INV_X1 U332 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U333 ( .A1(data_in[3]), .A2(n837), .B1(n1065), .B2(\mem[15][3] ), 
        .ZN(n1062) );
  INV_X1 U334 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U335 ( .A1(data_in[4]), .A2(n837), .B1(n1065), .B2(\mem[15][4] ), 
        .ZN(n1061) );
  INV_X1 U336 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U337 ( .A1(data_in[5]), .A2(n837), .B1(n1065), .B2(\mem[15][5] ), 
        .ZN(n1060) );
  INV_X1 U338 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U339 ( .A1(data_in[6]), .A2(n837), .B1(n1065), .B2(\mem[15][6] ), 
        .ZN(n1059) );
  INV_X1 U340 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U341 ( .A1(data_in[7]), .A2(n837), .B1(n1065), .B2(\mem[15][7] ), 
        .ZN(n1058) );
  INV_X1 U342 ( .A(n1057), .ZN(n756) );
  AOI22_X1 U343 ( .A1(data_in[0]), .A2(n836), .B1(n1056), .B2(\mem[16][0] ), 
        .ZN(n1057) );
  INV_X1 U344 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U345 ( .A1(data_in[1]), .A2(n836), .B1(n1056), .B2(\mem[16][1] ), 
        .ZN(n1055) );
  INV_X1 U346 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U347 ( .A1(data_in[2]), .A2(n836), .B1(n1056), .B2(\mem[16][2] ), 
        .ZN(n1054) );
  INV_X1 U348 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U349 ( .A1(data_in[3]), .A2(n836), .B1(n1056), .B2(\mem[16][3] ), 
        .ZN(n1053) );
  INV_X1 U350 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U351 ( .A1(data_in[4]), .A2(n836), .B1(n1056), .B2(\mem[16][4] ), 
        .ZN(n1052) );
  INV_X1 U352 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U353 ( .A1(data_in[5]), .A2(n836), .B1(n1056), .B2(\mem[16][5] ), 
        .ZN(n1051) );
  INV_X1 U354 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U355 ( .A1(data_in[6]), .A2(n836), .B1(n1056), .B2(\mem[16][6] ), 
        .ZN(n1050) );
  INV_X1 U356 ( .A(n1049), .ZN(n749) );
  AOI22_X1 U357 ( .A1(data_in[7]), .A2(n836), .B1(n1056), .B2(\mem[16][7] ), 
        .ZN(n1049) );
  INV_X1 U358 ( .A(n1047), .ZN(n748) );
  AOI22_X1 U359 ( .A1(data_in[0]), .A2(n835), .B1(n1046), .B2(\mem[17][0] ), 
        .ZN(n1047) );
  INV_X1 U360 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U361 ( .A1(data_in[1]), .A2(n835), .B1(n1046), .B2(\mem[17][1] ), 
        .ZN(n1045) );
  INV_X1 U362 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U363 ( .A1(data_in[2]), .A2(n835), .B1(n1046), .B2(\mem[17][2] ), 
        .ZN(n1044) );
  INV_X1 U364 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[3]), .A2(n835), .B1(n1046), .B2(\mem[17][3] ), 
        .ZN(n1043) );
  INV_X1 U366 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[4]), .A2(n835), .B1(n1046), .B2(\mem[17][4] ), 
        .ZN(n1042) );
  INV_X1 U368 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[5]), .A2(n835), .B1(n1046), .B2(\mem[17][5] ), 
        .ZN(n1041) );
  INV_X1 U370 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[6]), .A2(n835), .B1(n1046), .B2(\mem[17][6] ), 
        .ZN(n1040) );
  INV_X1 U372 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[7]), .A2(n835), .B1(n1046), .B2(\mem[17][7] ), 
        .ZN(n1039) );
  INV_X1 U374 ( .A(n1038), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[0]), .A2(n834), .B1(n1037), .B2(\mem[18][0] ), 
        .ZN(n1038) );
  INV_X1 U376 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[1]), .A2(n834), .B1(n1037), .B2(\mem[18][1] ), 
        .ZN(n1036) );
  INV_X1 U378 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[2]), .A2(n834), .B1(n1037), .B2(\mem[18][2] ), 
        .ZN(n1035) );
  INV_X1 U380 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U381 ( .A1(data_in[3]), .A2(n834), .B1(n1037), .B2(\mem[18][3] ), 
        .ZN(n1034) );
  INV_X1 U382 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U383 ( .A1(data_in[4]), .A2(n834), .B1(n1037), .B2(\mem[18][4] ), 
        .ZN(n1033) );
  INV_X1 U384 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U385 ( .A1(data_in[5]), .A2(n834), .B1(n1037), .B2(\mem[18][5] ), 
        .ZN(n1032) );
  INV_X1 U386 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U387 ( .A1(data_in[6]), .A2(n834), .B1(n1037), .B2(\mem[18][6] ), 
        .ZN(n1031) );
  INV_X1 U388 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U389 ( .A1(data_in[7]), .A2(n834), .B1(n1037), .B2(\mem[18][7] ), 
        .ZN(n1030) );
  INV_X1 U390 ( .A(n1029), .ZN(n732) );
  AOI22_X1 U391 ( .A1(data_in[0]), .A2(n833), .B1(n1028), .B2(\mem[19][0] ), 
        .ZN(n1029) );
  INV_X1 U392 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U393 ( .A1(data_in[1]), .A2(n833), .B1(n1028), .B2(\mem[19][1] ), 
        .ZN(n1027) );
  INV_X1 U394 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U395 ( .A1(data_in[2]), .A2(n833), .B1(n1028), .B2(\mem[19][2] ), 
        .ZN(n1026) );
  INV_X1 U396 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U397 ( .A1(data_in[3]), .A2(n833), .B1(n1028), .B2(\mem[19][3] ), 
        .ZN(n1025) );
  INV_X1 U398 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U399 ( .A1(data_in[4]), .A2(n833), .B1(n1028), .B2(\mem[19][4] ), 
        .ZN(n1024) );
  INV_X1 U400 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U401 ( .A1(data_in[5]), .A2(n833), .B1(n1028), .B2(\mem[19][5] ), 
        .ZN(n1023) );
  INV_X1 U402 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U403 ( .A1(data_in[6]), .A2(n833), .B1(n1028), .B2(\mem[19][6] ), 
        .ZN(n1022) );
  INV_X1 U404 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U405 ( .A1(data_in[7]), .A2(n833), .B1(n1028), .B2(\mem[19][7] ), 
        .ZN(n1021) );
  INV_X1 U406 ( .A(n1020), .ZN(n724) );
  AOI22_X1 U407 ( .A1(data_in[0]), .A2(n832), .B1(n1019), .B2(\mem[20][0] ), 
        .ZN(n1020) );
  INV_X1 U408 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U409 ( .A1(data_in[1]), .A2(n832), .B1(n1019), .B2(\mem[20][1] ), 
        .ZN(n1018) );
  INV_X1 U410 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U411 ( .A1(data_in[2]), .A2(n832), .B1(n1019), .B2(\mem[20][2] ), 
        .ZN(n1017) );
  INV_X1 U412 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U413 ( .A1(data_in[3]), .A2(n832), .B1(n1019), .B2(\mem[20][3] ), 
        .ZN(n1016) );
  INV_X1 U414 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U415 ( .A1(data_in[4]), .A2(n832), .B1(n1019), .B2(\mem[20][4] ), 
        .ZN(n1015) );
  INV_X1 U416 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U417 ( .A1(data_in[5]), .A2(n832), .B1(n1019), .B2(\mem[20][5] ), 
        .ZN(n1014) );
  INV_X1 U418 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U419 ( .A1(data_in[6]), .A2(n832), .B1(n1019), .B2(\mem[20][6] ), 
        .ZN(n1013) );
  INV_X1 U420 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U421 ( .A1(data_in[7]), .A2(n832), .B1(n1019), .B2(\mem[20][7] ), 
        .ZN(n1012) );
  INV_X1 U422 ( .A(n1011), .ZN(n716) );
  AOI22_X1 U423 ( .A1(data_in[0]), .A2(n831), .B1(n1010), .B2(\mem[21][0] ), 
        .ZN(n1011) );
  INV_X1 U424 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U425 ( .A1(data_in[1]), .A2(n831), .B1(n1010), .B2(\mem[21][1] ), 
        .ZN(n1009) );
  INV_X1 U426 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U427 ( .A1(data_in[2]), .A2(n831), .B1(n1010), .B2(\mem[21][2] ), 
        .ZN(n1008) );
  INV_X1 U428 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U429 ( .A1(data_in[3]), .A2(n831), .B1(n1010), .B2(\mem[21][3] ), 
        .ZN(n1007) );
  INV_X1 U430 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U431 ( .A1(data_in[4]), .A2(n831), .B1(n1010), .B2(\mem[21][4] ), 
        .ZN(n1006) );
  INV_X1 U432 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U433 ( .A1(data_in[5]), .A2(n831), .B1(n1010), .B2(\mem[21][5] ), 
        .ZN(n1005) );
  INV_X1 U434 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U435 ( .A1(data_in[6]), .A2(n831), .B1(n1010), .B2(\mem[21][6] ), 
        .ZN(n1004) );
  INV_X1 U436 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U437 ( .A1(data_in[7]), .A2(n831), .B1(n1010), .B2(\mem[21][7] ), 
        .ZN(n1003) );
  INV_X1 U438 ( .A(n1002), .ZN(n708) );
  AOI22_X1 U439 ( .A1(data_in[0]), .A2(n830), .B1(n1001), .B2(\mem[22][0] ), 
        .ZN(n1002) );
  INV_X1 U440 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U441 ( .A1(data_in[1]), .A2(n830), .B1(n1001), .B2(\mem[22][1] ), 
        .ZN(n1000) );
  INV_X1 U442 ( .A(n999), .ZN(n706) );
  AOI22_X1 U443 ( .A1(data_in[2]), .A2(n830), .B1(n1001), .B2(\mem[22][2] ), 
        .ZN(n999) );
  INV_X1 U444 ( .A(n998), .ZN(n705) );
  AOI22_X1 U445 ( .A1(data_in[3]), .A2(n830), .B1(n1001), .B2(\mem[22][3] ), 
        .ZN(n998) );
  INV_X1 U446 ( .A(n997), .ZN(n704) );
  AOI22_X1 U447 ( .A1(data_in[4]), .A2(n830), .B1(n1001), .B2(\mem[22][4] ), 
        .ZN(n997) );
  INV_X1 U448 ( .A(n996), .ZN(n703) );
  AOI22_X1 U449 ( .A1(data_in[5]), .A2(n830), .B1(n1001), .B2(\mem[22][5] ), 
        .ZN(n996) );
  INV_X1 U450 ( .A(n995), .ZN(n702) );
  AOI22_X1 U451 ( .A1(data_in[6]), .A2(n830), .B1(n1001), .B2(\mem[22][6] ), 
        .ZN(n995) );
  INV_X1 U452 ( .A(n994), .ZN(n701) );
  AOI22_X1 U453 ( .A1(data_in[7]), .A2(n830), .B1(n1001), .B2(\mem[22][7] ), 
        .ZN(n994) );
  INV_X1 U454 ( .A(n993), .ZN(n700) );
  AOI22_X1 U455 ( .A1(data_in[0]), .A2(n829), .B1(n992), .B2(\mem[23][0] ), 
        .ZN(n993) );
  INV_X1 U456 ( .A(n991), .ZN(n699) );
  AOI22_X1 U457 ( .A1(data_in[1]), .A2(n829), .B1(n992), .B2(\mem[23][1] ), 
        .ZN(n991) );
  INV_X1 U458 ( .A(n990), .ZN(n698) );
  AOI22_X1 U459 ( .A1(data_in[2]), .A2(n829), .B1(n992), .B2(\mem[23][2] ), 
        .ZN(n990) );
  INV_X1 U460 ( .A(n989), .ZN(n697) );
  AOI22_X1 U461 ( .A1(data_in[3]), .A2(n829), .B1(n992), .B2(\mem[23][3] ), 
        .ZN(n989) );
  INV_X1 U462 ( .A(n988), .ZN(n696) );
  AOI22_X1 U463 ( .A1(data_in[4]), .A2(n829), .B1(n992), .B2(\mem[23][4] ), 
        .ZN(n988) );
  INV_X1 U464 ( .A(n987), .ZN(n695) );
  AOI22_X1 U465 ( .A1(data_in[5]), .A2(n829), .B1(n992), .B2(\mem[23][5] ), 
        .ZN(n987) );
  INV_X1 U466 ( .A(n986), .ZN(n694) );
  AOI22_X1 U467 ( .A1(data_in[6]), .A2(n829), .B1(n992), .B2(\mem[23][6] ), 
        .ZN(n986) );
  INV_X1 U468 ( .A(n985), .ZN(n693) );
  AOI22_X1 U469 ( .A1(data_in[7]), .A2(n829), .B1(n992), .B2(\mem[23][7] ), 
        .ZN(n985) );
  INV_X1 U470 ( .A(n984), .ZN(n692) );
  AOI22_X1 U471 ( .A1(data_in[0]), .A2(n828), .B1(n983), .B2(\mem[24][0] ), 
        .ZN(n984) );
  INV_X1 U472 ( .A(n982), .ZN(n691) );
  AOI22_X1 U473 ( .A1(data_in[1]), .A2(n828), .B1(n983), .B2(\mem[24][1] ), 
        .ZN(n982) );
  INV_X1 U474 ( .A(n981), .ZN(n690) );
  AOI22_X1 U475 ( .A1(data_in[2]), .A2(n828), .B1(n983), .B2(\mem[24][2] ), 
        .ZN(n981) );
  INV_X1 U476 ( .A(n980), .ZN(n689) );
  AOI22_X1 U477 ( .A1(data_in[3]), .A2(n828), .B1(n983), .B2(\mem[24][3] ), 
        .ZN(n980) );
  INV_X1 U478 ( .A(n979), .ZN(n688) );
  AOI22_X1 U479 ( .A1(data_in[4]), .A2(n828), .B1(n983), .B2(\mem[24][4] ), 
        .ZN(n979) );
  INV_X1 U480 ( .A(n978), .ZN(n687) );
  AOI22_X1 U481 ( .A1(data_in[5]), .A2(n828), .B1(n983), .B2(\mem[24][5] ), 
        .ZN(n978) );
  INV_X1 U482 ( .A(n977), .ZN(n686) );
  AOI22_X1 U483 ( .A1(data_in[6]), .A2(n828), .B1(n983), .B2(\mem[24][6] ), 
        .ZN(n977) );
  INV_X1 U484 ( .A(n976), .ZN(n685) );
  AOI22_X1 U485 ( .A1(data_in[7]), .A2(n828), .B1(n983), .B2(\mem[24][7] ), 
        .ZN(n976) );
  INV_X1 U486 ( .A(n974), .ZN(n684) );
  AOI22_X1 U487 ( .A1(data_in[0]), .A2(n827), .B1(n973), .B2(\mem[25][0] ), 
        .ZN(n974) );
  INV_X1 U488 ( .A(n972), .ZN(n683) );
  AOI22_X1 U489 ( .A1(data_in[1]), .A2(n827), .B1(n973), .B2(\mem[25][1] ), 
        .ZN(n972) );
  INV_X1 U490 ( .A(n971), .ZN(n682) );
  AOI22_X1 U491 ( .A1(data_in[2]), .A2(n827), .B1(n973), .B2(\mem[25][2] ), 
        .ZN(n971) );
  INV_X1 U492 ( .A(n970), .ZN(n681) );
  AOI22_X1 U493 ( .A1(data_in[3]), .A2(n827), .B1(n973), .B2(\mem[25][3] ), 
        .ZN(n970) );
  INV_X1 U494 ( .A(n969), .ZN(n680) );
  AOI22_X1 U495 ( .A1(data_in[4]), .A2(n827), .B1(n973), .B2(\mem[25][4] ), 
        .ZN(n969) );
  INV_X1 U496 ( .A(n968), .ZN(n679) );
  AOI22_X1 U497 ( .A1(data_in[5]), .A2(n827), .B1(n973), .B2(\mem[25][5] ), 
        .ZN(n968) );
  INV_X1 U498 ( .A(n967), .ZN(n678) );
  AOI22_X1 U499 ( .A1(data_in[6]), .A2(n827), .B1(n973), .B2(\mem[25][6] ), 
        .ZN(n967) );
  INV_X1 U500 ( .A(n966), .ZN(n677) );
  AOI22_X1 U501 ( .A1(data_in[7]), .A2(n827), .B1(n973), .B2(\mem[25][7] ), 
        .ZN(n966) );
  INV_X1 U502 ( .A(n965), .ZN(n676) );
  AOI22_X1 U503 ( .A1(data_in[0]), .A2(n826), .B1(n964), .B2(\mem[26][0] ), 
        .ZN(n965) );
  INV_X1 U504 ( .A(n963), .ZN(n675) );
  AOI22_X1 U505 ( .A1(data_in[1]), .A2(n826), .B1(n964), .B2(\mem[26][1] ), 
        .ZN(n963) );
  INV_X1 U506 ( .A(n962), .ZN(n674) );
  AOI22_X1 U507 ( .A1(data_in[2]), .A2(n826), .B1(n964), .B2(\mem[26][2] ), 
        .ZN(n962) );
  INV_X1 U508 ( .A(n961), .ZN(n673) );
  AOI22_X1 U509 ( .A1(data_in[3]), .A2(n826), .B1(n964), .B2(\mem[26][3] ), 
        .ZN(n961) );
  INV_X1 U510 ( .A(n960), .ZN(n672) );
  AOI22_X1 U511 ( .A1(data_in[4]), .A2(n826), .B1(n964), .B2(\mem[26][4] ), 
        .ZN(n960) );
  INV_X1 U512 ( .A(n959), .ZN(n671) );
  AOI22_X1 U513 ( .A1(data_in[5]), .A2(n826), .B1(n964), .B2(\mem[26][5] ), 
        .ZN(n959) );
  INV_X1 U514 ( .A(n958), .ZN(n670) );
  AOI22_X1 U515 ( .A1(data_in[6]), .A2(n826), .B1(n964), .B2(\mem[26][6] ), 
        .ZN(n958) );
  INV_X1 U516 ( .A(n957), .ZN(n669) );
  AOI22_X1 U517 ( .A1(data_in[7]), .A2(n826), .B1(n964), .B2(\mem[26][7] ), 
        .ZN(n957) );
  INV_X1 U518 ( .A(n956), .ZN(n668) );
  AOI22_X1 U519 ( .A1(data_in[0]), .A2(n825), .B1(n955), .B2(\mem[27][0] ), 
        .ZN(n956) );
  INV_X1 U520 ( .A(n954), .ZN(n667) );
  AOI22_X1 U521 ( .A1(data_in[1]), .A2(n825), .B1(n955), .B2(\mem[27][1] ), 
        .ZN(n954) );
  INV_X1 U522 ( .A(n953), .ZN(n666) );
  AOI22_X1 U523 ( .A1(data_in[2]), .A2(n825), .B1(n955), .B2(\mem[27][2] ), 
        .ZN(n953) );
  INV_X1 U524 ( .A(n952), .ZN(n665) );
  AOI22_X1 U525 ( .A1(data_in[3]), .A2(n825), .B1(n955), .B2(\mem[27][3] ), 
        .ZN(n952) );
  INV_X1 U526 ( .A(n951), .ZN(n664) );
  AOI22_X1 U527 ( .A1(data_in[4]), .A2(n825), .B1(n955), .B2(\mem[27][4] ), 
        .ZN(n951) );
  INV_X1 U528 ( .A(n950), .ZN(n663) );
  AOI22_X1 U529 ( .A1(data_in[5]), .A2(n825), .B1(n955), .B2(\mem[27][5] ), 
        .ZN(n950) );
  INV_X1 U530 ( .A(n949), .ZN(n662) );
  AOI22_X1 U531 ( .A1(data_in[6]), .A2(n825), .B1(n955), .B2(\mem[27][6] ), 
        .ZN(n949) );
  INV_X1 U532 ( .A(n948), .ZN(n661) );
  AOI22_X1 U533 ( .A1(data_in[7]), .A2(n825), .B1(n955), .B2(\mem[27][7] ), 
        .ZN(n948) );
  INV_X1 U534 ( .A(n947), .ZN(n660) );
  AOI22_X1 U535 ( .A1(data_in[0]), .A2(n824), .B1(n946), .B2(\mem[28][0] ), 
        .ZN(n947) );
  INV_X1 U536 ( .A(n945), .ZN(n659) );
  AOI22_X1 U537 ( .A1(data_in[1]), .A2(n824), .B1(n946), .B2(\mem[28][1] ), 
        .ZN(n945) );
  INV_X1 U538 ( .A(n944), .ZN(n658) );
  AOI22_X1 U539 ( .A1(data_in[2]), .A2(n824), .B1(n946), .B2(\mem[28][2] ), 
        .ZN(n944) );
  INV_X1 U540 ( .A(n943), .ZN(n657) );
  AOI22_X1 U541 ( .A1(data_in[3]), .A2(n824), .B1(n946), .B2(\mem[28][3] ), 
        .ZN(n943) );
  INV_X1 U542 ( .A(n942), .ZN(n656) );
  AOI22_X1 U543 ( .A1(data_in[4]), .A2(n824), .B1(n946), .B2(\mem[28][4] ), 
        .ZN(n942) );
  INV_X1 U544 ( .A(n941), .ZN(n655) );
  AOI22_X1 U545 ( .A1(data_in[5]), .A2(n824), .B1(n946), .B2(\mem[28][5] ), 
        .ZN(n941) );
  INV_X1 U546 ( .A(n940), .ZN(n654) );
  AOI22_X1 U547 ( .A1(data_in[6]), .A2(n824), .B1(n946), .B2(\mem[28][6] ), 
        .ZN(n940) );
  INV_X1 U548 ( .A(n939), .ZN(n653) );
  AOI22_X1 U549 ( .A1(data_in[7]), .A2(n824), .B1(n946), .B2(\mem[28][7] ), 
        .ZN(n939) );
  INV_X1 U550 ( .A(n938), .ZN(n652) );
  AOI22_X1 U551 ( .A1(data_in[0]), .A2(n823), .B1(n937), .B2(\mem[29][0] ), 
        .ZN(n938) );
  INV_X1 U552 ( .A(n936), .ZN(n651) );
  AOI22_X1 U553 ( .A1(data_in[1]), .A2(n823), .B1(n937), .B2(\mem[29][1] ), 
        .ZN(n936) );
  INV_X1 U554 ( .A(n935), .ZN(n650) );
  AOI22_X1 U555 ( .A1(data_in[2]), .A2(n823), .B1(n937), .B2(\mem[29][2] ), 
        .ZN(n935) );
  INV_X1 U556 ( .A(n934), .ZN(n649) );
  AOI22_X1 U557 ( .A1(data_in[3]), .A2(n823), .B1(n937), .B2(\mem[29][3] ), 
        .ZN(n934) );
  INV_X1 U558 ( .A(n933), .ZN(n648) );
  AOI22_X1 U559 ( .A1(data_in[4]), .A2(n823), .B1(n937), .B2(\mem[29][4] ), 
        .ZN(n933) );
  INV_X1 U560 ( .A(n932), .ZN(n647) );
  AOI22_X1 U561 ( .A1(data_in[5]), .A2(n823), .B1(n937), .B2(\mem[29][5] ), 
        .ZN(n932) );
  INV_X1 U562 ( .A(n931), .ZN(n646) );
  AOI22_X1 U563 ( .A1(data_in[6]), .A2(n823), .B1(n937), .B2(\mem[29][6] ), 
        .ZN(n931) );
  INV_X1 U564 ( .A(n930), .ZN(n645) );
  AOI22_X1 U565 ( .A1(data_in[7]), .A2(n823), .B1(n937), .B2(\mem[29][7] ), 
        .ZN(n930) );
  INV_X1 U566 ( .A(n929), .ZN(n644) );
  AOI22_X1 U567 ( .A1(data_in[0]), .A2(n822), .B1(n928), .B2(\mem[30][0] ), 
        .ZN(n929) );
  INV_X1 U568 ( .A(n927), .ZN(n643) );
  AOI22_X1 U569 ( .A1(data_in[1]), .A2(n822), .B1(n928), .B2(\mem[30][1] ), 
        .ZN(n927) );
  INV_X1 U570 ( .A(n926), .ZN(n642) );
  AOI22_X1 U571 ( .A1(data_in[2]), .A2(n822), .B1(n928), .B2(\mem[30][2] ), 
        .ZN(n926) );
  INV_X1 U572 ( .A(n925), .ZN(n641) );
  AOI22_X1 U573 ( .A1(data_in[3]), .A2(n822), .B1(n928), .B2(\mem[30][3] ), 
        .ZN(n925) );
  INV_X1 U574 ( .A(n924), .ZN(n640) );
  AOI22_X1 U575 ( .A1(data_in[4]), .A2(n822), .B1(n928), .B2(\mem[30][4] ), 
        .ZN(n924) );
  INV_X1 U576 ( .A(n923), .ZN(n639) );
  AOI22_X1 U577 ( .A1(data_in[5]), .A2(n822), .B1(n928), .B2(\mem[30][5] ), 
        .ZN(n923) );
  INV_X1 U578 ( .A(n922), .ZN(n638) );
  AOI22_X1 U579 ( .A1(data_in[6]), .A2(n822), .B1(n928), .B2(\mem[30][6] ), 
        .ZN(n922) );
  INV_X1 U580 ( .A(n921), .ZN(n637) );
  AOI22_X1 U581 ( .A1(data_in[7]), .A2(n822), .B1(n928), .B2(\mem[30][7] ), 
        .ZN(n921) );
  INV_X1 U582 ( .A(n920), .ZN(n636) );
  AOI22_X1 U583 ( .A1(data_in[0]), .A2(n821), .B1(n919), .B2(\mem[31][0] ), 
        .ZN(n920) );
  INV_X1 U584 ( .A(n918), .ZN(n635) );
  AOI22_X1 U585 ( .A1(data_in[1]), .A2(n821), .B1(n919), .B2(\mem[31][1] ), 
        .ZN(n918) );
  INV_X1 U586 ( .A(n917), .ZN(n634) );
  AOI22_X1 U587 ( .A1(data_in[2]), .A2(n821), .B1(n919), .B2(\mem[31][2] ), 
        .ZN(n917) );
  INV_X1 U588 ( .A(n916), .ZN(n633) );
  AOI22_X1 U589 ( .A1(data_in[3]), .A2(n821), .B1(n919), .B2(\mem[31][3] ), 
        .ZN(n916) );
  INV_X1 U590 ( .A(n915), .ZN(n632) );
  AOI22_X1 U591 ( .A1(data_in[4]), .A2(n821), .B1(n919), .B2(\mem[31][4] ), 
        .ZN(n915) );
  INV_X1 U592 ( .A(n914), .ZN(n631) );
  AOI22_X1 U593 ( .A1(data_in[5]), .A2(n821), .B1(n919), .B2(\mem[31][5] ), 
        .ZN(n914) );
  INV_X1 U594 ( .A(n913), .ZN(n630) );
  AOI22_X1 U595 ( .A1(data_in[6]), .A2(n821), .B1(n919), .B2(\mem[31][6] ), 
        .ZN(n913) );
  INV_X1 U596 ( .A(n912), .ZN(n629) );
  AOI22_X1 U597 ( .A1(data_in[7]), .A2(n821), .B1(n919), .B2(\mem[31][7] ), 
        .ZN(n912) );
  MUX2_X1 U598 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n615), .Z(n3) );
  MUX2_X1 U599 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n615), .Z(n4) );
  MUX2_X1 U600 ( .A(n4), .B(n3), .S(n610), .Z(n5) );
  MUX2_X1 U601 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n615), .Z(n6) );
  MUX2_X1 U602 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n615), .Z(n7) );
  MUX2_X1 U603 ( .A(n7), .B(n6), .S(n610), .Z(n8) );
  MUX2_X1 U604 ( .A(n8), .B(n5), .S(n608), .Z(n9) );
  MUX2_X1 U605 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n615), .Z(n10) );
  MUX2_X1 U606 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n615), .Z(n11) );
  MUX2_X1 U607 ( .A(n11), .B(n10), .S(n610), .Z(n12) );
  MUX2_X1 U608 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n615), .Z(n13) );
  MUX2_X1 U609 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n615), .Z(n14) );
  MUX2_X1 U610 ( .A(n14), .B(n13), .S(n610), .Z(n15) );
  MUX2_X1 U611 ( .A(n15), .B(n12), .S(N12), .Z(n16) );
  MUX2_X1 U612 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U613 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n613), .Z(n18) );
  MUX2_X1 U614 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n613), .Z(n19) );
  MUX2_X1 U615 ( .A(n19), .B(n18), .S(n610), .Z(n20) );
  MUX2_X1 U616 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n613), .Z(n21) );
  MUX2_X1 U617 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n613), .Z(n22) );
  MUX2_X1 U618 ( .A(n22), .B(n21), .S(n611), .Z(n23) );
  MUX2_X1 U619 ( .A(n23), .B(n20), .S(N12), .Z(n24) );
  MUX2_X1 U620 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n613), .Z(n25) );
  MUX2_X1 U621 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n613), .Z(n26) );
  MUX2_X1 U622 ( .A(n26), .B(n25), .S(n610), .Z(n27) );
  MUX2_X1 U623 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n613), .Z(n28) );
  MUX2_X1 U624 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n613), .Z(n29) );
  MUX2_X1 U625 ( .A(n29), .B(n28), .S(N11), .Z(n30) );
  MUX2_X1 U626 ( .A(n30), .B(n27), .S(n609), .Z(n31) );
  MUX2_X1 U627 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U628 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U629 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n613), .Z(n33) );
  MUX2_X1 U630 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n613), .Z(n34) );
  MUX2_X1 U631 ( .A(n34), .B(n33), .S(n610), .Z(n35) );
  MUX2_X1 U632 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n613), .Z(n36) );
  MUX2_X1 U633 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n613), .Z(n37) );
  MUX2_X1 U634 ( .A(n37), .B(n36), .S(n610), .Z(n38) );
  MUX2_X1 U635 ( .A(n38), .B(n35), .S(n609), .Z(n39) );
  MUX2_X1 U636 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n614), .Z(n40) );
  MUX2_X1 U637 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n616), .Z(n41) );
  MUX2_X1 U638 ( .A(n41), .B(n40), .S(n610), .Z(n42) );
  MUX2_X1 U639 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n613), .Z(n43) );
  MUX2_X1 U640 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n616), .Z(n44) );
  MUX2_X1 U641 ( .A(n44), .B(n43), .S(n611), .Z(n45) );
  MUX2_X1 U642 ( .A(n45), .B(n42), .S(n608), .Z(n46) );
  MUX2_X1 U643 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U644 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n617), .Z(n48) );
  MUX2_X1 U645 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n617), .Z(n49) );
  MUX2_X1 U646 ( .A(n49), .B(n48), .S(n610), .Z(n50) );
  MUX2_X1 U647 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n617), .Z(n51) );
  MUX2_X1 U648 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n613), .Z(n52) );
  MUX2_X1 U649 ( .A(n52), .B(n51), .S(n612), .Z(n53) );
  MUX2_X1 U650 ( .A(n53), .B(n50), .S(N12), .Z(n54) );
  MUX2_X1 U651 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n613), .Z(n55) );
  MUX2_X1 U652 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n614), .Z(n56) );
  MUX2_X1 U653 ( .A(n56), .B(n55), .S(n610), .Z(n57) );
  MUX2_X1 U654 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n613), .Z(n58) );
  MUX2_X1 U655 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n617), .Z(n59) );
  MUX2_X1 U656 ( .A(n59), .B(n58), .S(n610), .Z(n60) );
  MUX2_X1 U657 ( .A(n60), .B(n57), .S(n608), .Z(n61) );
  MUX2_X1 U658 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U659 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U660 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n616), .Z(n63) );
  MUX2_X1 U661 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n616), .Z(n64) );
  MUX2_X1 U662 ( .A(n64), .B(n63), .S(n611), .Z(n65) );
  MUX2_X1 U663 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n618), .Z(n66) );
  MUX2_X1 U664 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n614), .Z(n67) );
  MUX2_X1 U665 ( .A(n67), .B(n66), .S(n611), .Z(n68) );
  MUX2_X1 U666 ( .A(n68), .B(n65), .S(n608), .Z(n69) );
  MUX2_X1 U667 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n614), .Z(n70) );
  MUX2_X1 U668 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n614), .Z(n71) );
  MUX2_X1 U669 ( .A(n71), .B(n70), .S(n611), .Z(n72) );
  MUX2_X1 U670 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n616), .Z(n73) );
  MUX2_X1 U671 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n616), .Z(n74) );
  MUX2_X1 U672 ( .A(n74), .B(n73), .S(n611), .Z(n75) );
  MUX2_X1 U673 ( .A(n75), .B(n72), .S(n608), .Z(n76) );
  MUX2_X1 U674 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U675 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n613), .Z(n78) );
  MUX2_X1 U676 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n613), .Z(n79) );
  MUX2_X1 U677 ( .A(n79), .B(n78), .S(n611), .Z(n80) );
  MUX2_X1 U678 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n617), .Z(n81) );
  MUX2_X1 U679 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n617), .Z(n82) );
  MUX2_X1 U680 ( .A(n82), .B(n81), .S(n611), .Z(n83) );
  MUX2_X1 U681 ( .A(n83), .B(n80), .S(n608), .Z(n84) );
  MUX2_X1 U682 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n618), .Z(n85) );
  MUX2_X1 U683 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n614), .Z(n86) );
  MUX2_X1 U684 ( .A(n86), .B(n85), .S(n611), .Z(n87) );
  MUX2_X1 U685 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n618), .Z(n88) );
  MUX2_X1 U686 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n617), .Z(n89) );
  MUX2_X1 U687 ( .A(n89), .B(n88), .S(n611), .Z(n90) );
  MUX2_X1 U688 ( .A(n90), .B(n87), .S(n608), .Z(n91) );
  MUX2_X1 U689 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U690 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U691 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n616), .Z(n93) );
  MUX2_X1 U692 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n618), .Z(n94) );
  MUX2_X1 U693 ( .A(n94), .B(n93), .S(n611), .Z(n95) );
  MUX2_X1 U694 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n618), .Z(n96) );
  MUX2_X1 U695 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n618), .Z(n97) );
  MUX2_X1 U696 ( .A(n97), .B(n96), .S(n611), .Z(n98) );
  MUX2_X1 U697 ( .A(n98), .B(n95), .S(n608), .Z(n99) );
  MUX2_X1 U698 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n618), .Z(n100) );
  MUX2_X1 U699 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n618), .Z(n101) );
  MUX2_X1 U700 ( .A(n101), .B(n100), .S(n611), .Z(n102) );
  MUX2_X1 U701 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n618), .Z(n103) );
  MUX2_X1 U702 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n613), .Z(n104) );
  MUX2_X1 U703 ( .A(n104), .B(n103), .S(n611), .Z(n105) );
  MUX2_X1 U704 ( .A(n105), .B(n102), .S(n608), .Z(n106) );
  MUX2_X1 U705 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U706 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n614), .Z(n108) );
  MUX2_X1 U707 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n614), .Z(n109) );
  MUX2_X1 U708 ( .A(n109), .B(n108), .S(n612), .Z(n110) );
  MUX2_X1 U709 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n614), .Z(n111) );
  MUX2_X1 U710 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n614), .Z(n112) );
  MUX2_X1 U711 ( .A(n112), .B(n111), .S(n612), .Z(n113) );
  MUX2_X1 U712 ( .A(n113), .B(n110), .S(n608), .Z(n114) );
  MUX2_X1 U713 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n614), .Z(n115) );
  MUX2_X1 U714 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n614), .Z(n116) );
  MUX2_X1 U715 ( .A(n116), .B(n115), .S(n612), .Z(n117) );
  MUX2_X1 U716 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n614), .Z(n118) );
  MUX2_X1 U717 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n614), .Z(n119) );
  MUX2_X1 U718 ( .A(n119), .B(n118), .S(n612), .Z(n120) );
  MUX2_X1 U719 ( .A(n120), .B(n117), .S(n608), .Z(n121) );
  MUX2_X1 U720 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U721 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U722 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n614), .Z(n123) );
  MUX2_X1 U723 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n614), .Z(n124) );
  MUX2_X1 U724 ( .A(n124), .B(n123), .S(n612), .Z(n125) );
  MUX2_X1 U725 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n614), .Z(n126) );
  MUX2_X1 U726 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n614), .Z(n127) );
  MUX2_X1 U727 ( .A(n127), .B(n126), .S(n612), .Z(n128) );
  MUX2_X1 U728 ( .A(n128), .B(n125), .S(n608), .Z(n129) );
  MUX2_X1 U729 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n615), .Z(n130) );
  MUX2_X1 U730 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n615), .Z(n131) );
  MUX2_X1 U731 ( .A(n131), .B(n130), .S(n612), .Z(n132) );
  MUX2_X1 U732 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n615), .Z(n133) );
  MUX2_X1 U733 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n615), .Z(n134) );
  MUX2_X1 U734 ( .A(n134), .B(n133), .S(n612), .Z(n135) );
  MUX2_X1 U735 ( .A(n135), .B(n132), .S(n608), .Z(n136) );
  MUX2_X1 U736 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U737 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n615), .Z(n138) );
  MUX2_X1 U738 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n615), .Z(n139) );
  MUX2_X1 U739 ( .A(n139), .B(n138), .S(n612), .Z(n140) );
  MUX2_X1 U740 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n615), .Z(n141) );
  MUX2_X1 U741 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n615), .Z(n142) );
  MUX2_X1 U742 ( .A(n142), .B(n141), .S(n612), .Z(n143) );
  MUX2_X1 U743 ( .A(n143), .B(n140), .S(n608), .Z(n144) );
  MUX2_X1 U744 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n615), .Z(n145) );
  MUX2_X1 U745 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n615), .Z(n146) );
  MUX2_X1 U746 ( .A(n146), .B(n145), .S(n612), .Z(n147) );
  MUX2_X1 U747 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n615), .Z(n148) );
  MUX2_X1 U748 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n615), .Z(n149) );
  MUX2_X1 U749 ( .A(n149), .B(n148), .S(n612), .Z(n150) );
  MUX2_X1 U750 ( .A(n150), .B(n147), .S(n608), .Z(n151) );
  MUX2_X1 U751 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U752 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U753 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n616), .Z(n153) );
  MUX2_X1 U754 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n616), .Z(n154) );
  MUX2_X1 U755 ( .A(n154), .B(n153), .S(n610), .Z(n155) );
  MUX2_X1 U756 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n616), .Z(n156) );
  MUX2_X1 U757 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n616), .Z(n157) );
  MUX2_X1 U758 ( .A(n157), .B(n156), .S(n612), .Z(n158) );
  MUX2_X1 U759 ( .A(n158), .B(n155), .S(n609), .Z(n159) );
  MUX2_X1 U760 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n616), .Z(n160) );
  MUX2_X1 U761 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n616), .Z(n161) );
  MUX2_X1 U762 ( .A(n161), .B(n160), .S(N11), .Z(n162) );
  MUX2_X1 U763 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n616), .Z(n163) );
  MUX2_X1 U764 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n616), .Z(n164) );
  MUX2_X1 U765 ( .A(n164), .B(n163), .S(n612), .Z(n165) );
  MUX2_X1 U766 ( .A(n165), .B(n162), .S(n609), .Z(n166) );
  MUX2_X1 U767 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U768 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n616), .Z(n168) );
  MUX2_X1 U769 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n616), .Z(n169) );
  MUX2_X1 U770 ( .A(n169), .B(n168), .S(n612), .Z(n170) );
  MUX2_X1 U771 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n616), .Z(n171) );
  MUX2_X1 U772 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n616), .Z(n172) );
  MUX2_X1 U773 ( .A(n172), .B(n171), .S(n612), .Z(n173) );
  MUX2_X1 U774 ( .A(n173), .B(n170), .S(n609), .Z(n174) );
  MUX2_X1 U775 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n618), .Z(n175) );
  MUX2_X1 U776 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n618), .Z(n176) );
  MUX2_X1 U777 ( .A(n176), .B(n175), .S(n611), .Z(n177) );
  MUX2_X1 U778 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n618), .Z(n178) );
  MUX2_X1 U779 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n179) );
  MUX2_X1 U780 ( .A(n179), .B(n178), .S(n611), .Z(n180) );
  MUX2_X1 U781 ( .A(n180), .B(n177), .S(n609), .Z(n181) );
  MUX2_X1 U782 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U783 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U784 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n613), .Z(n183) );
  MUX2_X1 U785 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n618), .Z(n184) );
  MUX2_X1 U786 ( .A(n184), .B(n183), .S(n611), .Z(n185) );
  MUX2_X1 U787 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n618), .Z(n186) );
  MUX2_X1 U788 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n614), .Z(n187) );
  MUX2_X1 U789 ( .A(n187), .B(n186), .S(n610), .Z(n188) );
  MUX2_X1 U790 ( .A(n188), .B(n185), .S(n609), .Z(n189) );
  MUX2_X1 U791 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n618), .Z(n190) );
  MUX2_X1 U792 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n618), .Z(n191) );
  MUX2_X1 U793 ( .A(n191), .B(n190), .S(n611), .Z(n192) );
  MUX2_X1 U794 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n616), .Z(n193) );
  MUX2_X1 U795 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n617), .Z(n194) );
  MUX2_X1 U796 ( .A(n194), .B(n193), .S(n610), .Z(n195) );
  MUX2_X1 U797 ( .A(n195), .B(n192), .S(n609), .Z(n196) );
  MUX2_X1 U798 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U799 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n614), .Z(n198) );
  MUX2_X1 U800 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n618), .Z(n199) );
  MUX2_X1 U801 ( .A(n199), .B(n198), .S(n612), .Z(n200) );
  MUX2_X1 U802 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n618), .Z(n201) );
  MUX2_X1 U803 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n202) );
  MUX2_X1 U804 ( .A(n202), .B(n201), .S(n612), .Z(n203) );
  MUX2_X1 U805 ( .A(n203), .B(n200), .S(n609), .Z(n204) );
  MUX2_X1 U806 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n618), .Z(n205) );
  MUX2_X1 U807 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n206) );
  MUX2_X1 U808 ( .A(n206), .B(n205), .S(N11), .Z(n207) );
  MUX2_X1 U809 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n208) );
  MUX2_X1 U810 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n209) );
  MUX2_X1 U811 ( .A(n209), .B(n208), .S(n611), .Z(n210) );
  MUX2_X1 U812 ( .A(n210), .B(n207), .S(n609), .Z(n211) );
  MUX2_X1 U813 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U814 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U815 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n615), .Z(n213) );
  MUX2_X1 U816 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n615), .Z(n214) );
  MUX2_X1 U817 ( .A(n214), .B(n213), .S(n611), .Z(n215) );
  MUX2_X1 U818 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n615), .Z(n216) );
  MUX2_X1 U819 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n618), .Z(n217) );
  MUX2_X1 U820 ( .A(n217), .B(n216), .S(N11), .Z(n218) );
  MUX2_X1 U821 ( .A(n218), .B(n215), .S(n609), .Z(n219) );
  MUX2_X1 U822 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n617), .Z(n220) );
  MUX2_X1 U823 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n617), .Z(n221) );
  MUX2_X1 U824 ( .A(n221), .B(n220), .S(n610), .Z(n222) );
  MUX2_X1 U825 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n617), .Z(n223) );
  MUX2_X1 U826 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n617), .Z(n224) );
  MUX2_X1 U827 ( .A(n224), .B(n223), .S(N11), .Z(n225) );
  MUX2_X1 U828 ( .A(n225), .B(n222), .S(n609), .Z(n226) );
  MUX2_X1 U829 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U830 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n617), .Z(n228) );
  MUX2_X1 U831 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n617), .Z(n229) );
  MUX2_X1 U832 ( .A(n229), .B(n228), .S(n610), .Z(n595) );
  MUX2_X1 U833 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n617), .Z(n596) );
  MUX2_X1 U834 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n617), .Z(n597) );
  MUX2_X1 U835 ( .A(n597), .B(n596), .S(n610), .Z(n598) );
  MUX2_X1 U836 ( .A(n598), .B(n595), .S(n609), .Z(n599) );
  MUX2_X1 U837 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n617), .Z(n600) );
  MUX2_X1 U838 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n617), .Z(n601) );
  MUX2_X1 U839 ( .A(n601), .B(n600), .S(n611), .Z(n602) );
  MUX2_X1 U840 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n617), .Z(n603) );
  MUX2_X1 U841 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n617), .Z(n604) );
  MUX2_X1 U842 ( .A(n604), .B(n603), .S(n612), .Z(n605) );
  MUX2_X1 U843 ( .A(n605), .B(n602), .S(n609), .Z(n606) );
  MUX2_X1 U844 ( .A(n606), .B(n599), .S(N13), .Z(n607) );
  MUX2_X1 U845 ( .A(n607), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U846 ( .A(N11), .Z(n610) );
  INV_X1 U847 ( .A(N10), .ZN(n619) );
  INV_X1 U848 ( .A(N11), .ZN(n620) );
  INV_X1 U849 ( .A(data_in[0]), .ZN(n621) );
  INV_X1 U850 ( .A(data_in[1]), .ZN(n622) );
  INV_X1 U851 ( .A(data_in[2]), .ZN(n623) );
  INV_X1 U852 ( .A(data_in[3]), .ZN(n624) );
  INV_X1 U853 ( .A(data_in[4]), .ZN(n625) );
  INV_X1 U854 ( .A(data_in[5]), .ZN(n626) );
  INV_X1 U855 ( .A(data_in[6]), .ZN(n627) );
  INV_X1 U856 ( .A(data_in[7]), .ZN(n628) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_15 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n633), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n634), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n635), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n636), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n637), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n638), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n639), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n640), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n641), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n642), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n643), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n644), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n645), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n646), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n647), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n648), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n649), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n650), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n651), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n652), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n653), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n654), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n655), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n656), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n657), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n658), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n659), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n660), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n661), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n662), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n663), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n664), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n665), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n666), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n667), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n668), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n669), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n670), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n671), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n672), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n673), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n674), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n675), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n676), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n677), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n678), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n679), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n680), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n681), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n682), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n683), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n684), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n685), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n686), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n687), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n688), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n689), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n690), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n691), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n692), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n693), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n694), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n695), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n696), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n697), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n698), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n699), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n700), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n701), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n702), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n703), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n704), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n705), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n706), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n707), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n708), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n709), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n710), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n711), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n712), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n713), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n714), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n715), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n716), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n717), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n718), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n719), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n720), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n721), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n722), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n723), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n724), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n725), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n726), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n727), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n728), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n729), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n730), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n731), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n732), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n733), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n734), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n735), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n736), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n737), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n738), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n739), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n740), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n741), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n742), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n743), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n744), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n745), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n746), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n747), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n748), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n749), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n750), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n751), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n752), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n753), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n754), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n755), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n756), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n757), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n758), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n759), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n760), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n761), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n762), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n763), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n764), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n765), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n766), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n767), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n768), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n769), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n770), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n771), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n772), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n773), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n774), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n775), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n776), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n777), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n778), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n779), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n780), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n781), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n782), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n783), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n784), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n785), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n786), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n787), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n788), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n789), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n790), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n791), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n792), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n793), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n794), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n795), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n796), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n797), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n798), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n799), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n800), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n801), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n802), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n803), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n804), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n805), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n806), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n807), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n808), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n809), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n810), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n811), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n812), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n813), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n814), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n815), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n816), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n817), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n818), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n819), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n820), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n821), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n822), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n823), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n824), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n852), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n853), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n854), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n855), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n856), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n857), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n858), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n859), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n860), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n861), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n862), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n863), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n864), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n865), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n866), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n867), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n868), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n869), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n870), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n871), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n872), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n873), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n874), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n875), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n876), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n877), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n878), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n879), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n880), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n881), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n882), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n883), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n884), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n885), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n886), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n887), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n888), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n889), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n890), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n891), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n892), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n893), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n894), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n895), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n896), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n897), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n898), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n899), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n900), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n901), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n902), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n903), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n904), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n905), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n906), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n907), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n908), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n909), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n910), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n911), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n912), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n913), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n914), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n915), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  BUF_X1 U3 ( .A(n621), .Z(n613) );
  CLKBUF_X1 U4 ( .A(N10), .Z(n621) );
  INV_X2 U5 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U6 ( .A(n622), .Z(n618) );
  BUF_X1 U7 ( .A(n622), .Z(n619) );
  BUF_X1 U8 ( .A(n622), .Z(n620) );
  BUF_X1 U9 ( .A(n621), .Z(n615) );
  BUF_X1 U10 ( .A(n621), .Z(n614) );
  BUF_X1 U11 ( .A(n621), .Z(n616) );
  BUF_X1 U12 ( .A(n621), .Z(n617) );
  BUF_X1 U13 ( .A(N11), .Z(n611) );
  BUF_X1 U14 ( .A(N11), .Z(n612) );
  BUF_X1 U15 ( .A(N10), .Z(n622) );
  NOR3_X1 U16 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1207) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(n623), .ZN(n1196) );
  NOR3_X1 U18 ( .A1(N10), .A2(N12), .A3(n624), .ZN(n1186) );
  NOR3_X1 U19 ( .A1(n623), .A2(N12), .A3(n624), .ZN(n1176) );
  INV_X1 U20 ( .A(n1133), .ZN(n848) );
  INV_X1 U21 ( .A(n1123), .ZN(n847) );
  INV_X1 U22 ( .A(n1114), .ZN(n846) );
  INV_X1 U23 ( .A(n1105), .ZN(n845) );
  INV_X1 U24 ( .A(n1060), .ZN(n840) );
  INV_X1 U25 ( .A(n1050), .ZN(n839) );
  INV_X1 U26 ( .A(n1041), .ZN(n838) );
  INV_X1 U27 ( .A(n1032), .ZN(n837) );
  INV_X1 U28 ( .A(n987), .ZN(n832) );
  INV_X1 U29 ( .A(n977), .ZN(n831) );
  INV_X1 U30 ( .A(n968), .ZN(n830) );
  INV_X1 U31 ( .A(n959), .ZN(n829) );
  INV_X1 U32 ( .A(n950), .ZN(n828) );
  INV_X1 U33 ( .A(n941), .ZN(n827) );
  INV_X1 U34 ( .A(n932), .ZN(n826) );
  INV_X1 U35 ( .A(n923), .ZN(n825) );
  INV_X1 U36 ( .A(n1096), .ZN(n844) );
  INV_X1 U37 ( .A(n1087), .ZN(n843) );
  INV_X1 U38 ( .A(n1078), .ZN(n842) );
  INV_X1 U39 ( .A(n1069), .ZN(n841) );
  INV_X1 U40 ( .A(n1023), .ZN(n836) );
  INV_X1 U41 ( .A(n1014), .ZN(n835) );
  INV_X1 U42 ( .A(n1005), .ZN(n834) );
  INV_X1 U43 ( .A(n996), .ZN(n833) );
  BUF_X1 U44 ( .A(N12), .Z(n608) );
  BUF_X1 U45 ( .A(N12), .Z(n609) );
  INV_X1 U46 ( .A(N13), .ZN(n850) );
  AND3_X1 U47 ( .A1(n623), .A2(n624), .A3(N12), .ZN(n1166) );
  AND3_X1 U48 ( .A1(N10), .A2(n624), .A3(N12), .ZN(n1156) );
  AND3_X1 U49 ( .A1(N11), .A2(n623), .A3(N12), .ZN(n1146) );
  AND3_X1 U50 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1136) );
  INV_X1 U51 ( .A(N14), .ZN(n851) );
  NAND2_X1 U52 ( .A1(n1196), .A2(n1206), .ZN(n1205) );
  NAND2_X1 U53 ( .A1(n1186), .A2(n1206), .ZN(n1195) );
  NAND2_X1 U54 ( .A1(n1176), .A2(n1206), .ZN(n1185) );
  NAND2_X1 U55 ( .A1(n1166), .A2(n1206), .ZN(n1175) );
  NAND2_X1 U56 ( .A1(n1156), .A2(n1206), .ZN(n1165) );
  NAND2_X1 U57 ( .A1(n1146), .A2(n1206), .ZN(n1155) );
  NAND2_X1 U58 ( .A1(n1136), .A2(n1206), .ZN(n1145) );
  NAND2_X1 U59 ( .A1(n1207), .A2(n1206), .ZN(n1216) );
  NAND2_X1 U60 ( .A1(n1125), .A2(n1207), .ZN(n1133) );
  NAND2_X1 U61 ( .A1(n1125), .A2(n1196), .ZN(n1123) );
  NAND2_X1 U62 ( .A1(n1125), .A2(n1186), .ZN(n1114) );
  NAND2_X1 U63 ( .A1(n1125), .A2(n1176), .ZN(n1105) );
  NAND2_X1 U64 ( .A1(n1052), .A2(n1207), .ZN(n1060) );
  NAND2_X1 U65 ( .A1(n1052), .A2(n1196), .ZN(n1050) );
  NAND2_X1 U66 ( .A1(n1052), .A2(n1186), .ZN(n1041) );
  NAND2_X1 U67 ( .A1(n1052), .A2(n1176), .ZN(n1032) );
  NAND2_X1 U68 ( .A1(n979), .A2(n1207), .ZN(n987) );
  NAND2_X1 U69 ( .A1(n979), .A2(n1196), .ZN(n977) );
  NAND2_X1 U70 ( .A1(n979), .A2(n1186), .ZN(n968) );
  NAND2_X1 U71 ( .A1(n979), .A2(n1176), .ZN(n959) );
  NAND2_X1 U72 ( .A1(n1125), .A2(n1166), .ZN(n1096) );
  NAND2_X1 U73 ( .A1(n1125), .A2(n1156), .ZN(n1087) );
  NAND2_X1 U74 ( .A1(n1125), .A2(n1146), .ZN(n1078) );
  NAND2_X1 U75 ( .A1(n1125), .A2(n1136), .ZN(n1069) );
  NAND2_X1 U76 ( .A1(n1052), .A2(n1166), .ZN(n1023) );
  NAND2_X1 U77 ( .A1(n1052), .A2(n1156), .ZN(n1014) );
  NAND2_X1 U78 ( .A1(n1052), .A2(n1146), .ZN(n1005) );
  NAND2_X1 U79 ( .A1(n1052), .A2(n1136), .ZN(n996) );
  NAND2_X1 U80 ( .A1(n979), .A2(n1166), .ZN(n950) );
  NAND2_X1 U81 ( .A1(n979), .A2(n1156), .ZN(n941) );
  NAND2_X1 U82 ( .A1(n979), .A2(n1146), .ZN(n932) );
  NAND2_X1 U83 ( .A1(n979), .A2(n1136), .ZN(n923) );
  AND3_X1 U84 ( .A1(n850), .A2(n851), .A3(n1135), .ZN(n1206) );
  AND3_X1 U85 ( .A1(N13), .A2(n1135), .A3(N14), .ZN(n979) );
  AND3_X1 U86 ( .A1(n1135), .A2(n851), .A3(N13), .ZN(n1125) );
  AND3_X1 U87 ( .A1(n1135), .A2(n850), .A3(N14), .ZN(n1052) );
  NOR2_X1 U88 ( .A1(n849), .A2(addr[5]), .ZN(n1135) );
  INV_X1 U89 ( .A(wr_en), .ZN(n849) );
  OAI21_X1 U90 ( .B1(n625), .B2(n1175), .A(n1174), .ZN(n883) );
  NAND2_X1 U91 ( .A1(\mem[4][0] ), .A2(n1175), .ZN(n1174) );
  OAI21_X1 U92 ( .B1(n626), .B2(n1175), .A(n1173), .ZN(n882) );
  NAND2_X1 U93 ( .A1(\mem[4][1] ), .A2(n1175), .ZN(n1173) );
  OAI21_X1 U94 ( .B1(n627), .B2(n1175), .A(n1172), .ZN(n881) );
  NAND2_X1 U95 ( .A1(\mem[4][2] ), .A2(n1175), .ZN(n1172) );
  OAI21_X1 U96 ( .B1(n628), .B2(n1175), .A(n1171), .ZN(n880) );
  NAND2_X1 U97 ( .A1(\mem[4][3] ), .A2(n1175), .ZN(n1171) );
  OAI21_X1 U98 ( .B1(n629), .B2(n1175), .A(n1170), .ZN(n879) );
  NAND2_X1 U99 ( .A1(\mem[4][4] ), .A2(n1175), .ZN(n1170) );
  OAI21_X1 U100 ( .B1(n630), .B2(n1175), .A(n1169), .ZN(n878) );
  NAND2_X1 U101 ( .A1(\mem[4][5] ), .A2(n1175), .ZN(n1169) );
  OAI21_X1 U102 ( .B1(n631), .B2(n1175), .A(n1168), .ZN(n877) );
  NAND2_X1 U103 ( .A1(\mem[4][6] ), .A2(n1175), .ZN(n1168) );
  OAI21_X1 U104 ( .B1(n632), .B2(n1175), .A(n1167), .ZN(n876) );
  NAND2_X1 U105 ( .A1(\mem[4][7] ), .A2(n1175), .ZN(n1167) );
  OAI21_X1 U106 ( .B1(n625), .B2(n1155), .A(n1154), .ZN(n867) );
  NAND2_X1 U107 ( .A1(\mem[6][0] ), .A2(n1155), .ZN(n1154) );
  OAI21_X1 U108 ( .B1(n626), .B2(n1155), .A(n1153), .ZN(n866) );
  NAND2_X1 U109 ( .A1(\mem[6][1] ), .A2(n1155), .ZN(n1153) );
  OAI21_X1 U110 ( .B1(n627), .B2(n1155), .A(n1152), .ZN(n865) );
  NAND2_X1 U111 ( .A1(\mem[6][2] ), .A2(n1155), .ZN(n1152) );
  OAI21_X1 U112 ( .B1(n628), .B2(n1155), .A(n1151), .ZN(n864) );
  NAND2_X1 U113 ( .A1(\mem[6][3] ), .A2(n1155), .ZN(n1151) );
  OAI21_X1 U114 ( .B1(n629), .B2(n1155), .A(n1150), .ZN(n863) );
  NAND2_X1 U115 ( .A1(\mem[6][4] ), .A2(n1155), .ZN(n1150) );
  OAI21_X1 U116 ( .B1(n630), .B2(n1155), .A(n1149), .ZN(n862) );
  NAND2_X1 U117 ( .A1(\mem[6][5] ), .A2(n1155), .ZN(n1149) );
  OAI21_X1 U118 ( .B1(n631), .B2(n1155), .A(n1148), .ZN(n861) );
  NAND2_X1 U119 ( .A1(\mem[6][6] ), .A2(n1155), .ZN(n1148) );
  OAI21_X1 U120 ( .B1(n632), .B2(n1155), .A(n1147), .ZN(n860) );
  NAND2_X1 U121 ( .A1(\mem[6][7] ), .A2(n1155), .ZN(n1147) );
  OAI21_X1 U122 ( .B1(n625), .B2(n1145), .A(n1144), .ZN(n859) );
  NAND2_X1 U123 ( .A1(\mem[7][0] ), .A2(n1145), .ZN(n1144) );
  OAI21_X1 U124 ( .B1(n626), .B2(n1145), .A(n1143), .ZN(n858) );
  NAND2_X1 U125 ( .A1(\mem[7][1] ), .A2(n1145), .ZN(n1143) );
  OAI21_X1 U126 ( .B1(n627), .B2(n1145), .A(n1142), .ZN(n857) );
  NAND2_X1 U127 ( .A1(\mem[7][2] ), .A2(n1145), .ZN(n1142) );
  OAI21_X1 U128 ( .B1(n628), .B2(n1145), .A(n1141), .ZN(n856) );
  NAND2_X1 U129 ( .A1(\mem[7][3] ), .A2(n1145), .ZN(n1141) );
  OAI21_X1 U130 ( .B1(n629), .B2(n1145), .A(n1140), .ZN(n855) );
  NAND2_X1 U131 ( .A1(\mem[7][4] ), .A2(n1145), .ZN(n1140) );
  OAI21_X1 U132 ( .B1(n630), .B2(n1145), .A(n1139), .ZN(n854) );
  NAND2_X1 U133 ( .A1(\mem[7][5] ), .A2(n1145), .ZN(n1139) );
  OAI21_X1 U134 ( .B1(n631), .B2(n1145), .A(n1138), .ZN(n853) );
  NAND2_X1 U135 ( .A1(\mem[7][6] ), .A2(n1145), .ZN(n1138) );
  OAI21_X1 U136 ( .B1(n632), .B2(n1145), .A(n1137), .ZN(n852) );
  NAND2_X1 U137 ( .A1(\mem[7][7] ), .A2(n1145), .ZN(n1137) );
  OAI21_X1 U138 ( .B1(n625), .B2(n1205), .A(n1204), .ZN(n907) );
  NAND2_X1 U139 ( .A1(\mem[1][0] ), .A2(n1205), .ZN(n1204) );
  OAI21_X1 U140 ( .B1(n626), .B2(n1205), .A(n1203), .ZN(n906) );
  NAND2_X1 U141 ( .A1(\mem[1][1] ), .A2(n1205), .ZN(n1203) );
  OAI21_X1 U142 ( .B1(n627), .B2(n1205), .A(n1202), .ZN(n905) );
  NAND2_X1 U143 ( .A1(\mem[1][2] ), .A2(n1205), .ZN(n1202) );
  OAI21_X1 U144 ( .B1(n628), .B2(n1205), .A(n1201), .ZN(n904) );
  NAND2_X1 U145 ( .A1(\mem[1][3] ), .A2(n1205), .ZN(n1201) );
  OAI21_X1 U146 ( .B1(n629), .B2(n1205), .A(n1200), .ZN(n903) );
  NAND2_X1 U147 ( .A1(\mem[1][4] ), .A2(n1205), .ZN(n1200) );
  OAI21_X1 U148 ( .B1(n630), .B2(n1205), .A(n1199), .ZN(n902) );
  NAND2_X1 U149 ( .A1(\mem[1][5] ), .A2(n1205), .ZN(n1199) );
  OAI21_X1 U150 ( .B1(n631), .B2(n1205), .A(n1198), .ZN(n901) );
  NAND2_X1 U151 ( .A1(\mem[1][6] ), .A2(n1205), .ZN(n1198) );
  OAI21_X1 U152 ( .B1(n632), .B2(n1205), .A(n1197), .ZN(n900) );
  NAND2_X1 U153 ( .A1(\mem[1][7] ), .A2(n1205), .ZN(n1197) );
  OAI21_X1 U154 ( .B1(n625), .B2(n1195), .A(n1194), .ZN(n899) );
  NAND2_X1 U155 ( .A1(\mem[2][0] ), .A2(n1195), .ZN(n1194) );
  OAI21_X1 U156 ( .B1(n626), .B2(n1195), .A(n1193), .ZN(n898) );
  NAND2_X1 U157 ( .A1(\mem[2][1] ), .A2(n1195), .ZN(n1193) );
  OAI21_X1 U158 ( .B1(n627), .B2(n1195), .A(n1192), .ZN(n897) );
  NAND2_X1 U159 ( .A1(\mem[2][2] ), .A2(n1195), .ZN(n1192) );
  OAI21_X1 U160 ( .B1(n628), .B2(n1195), .A(n1191), .ZN(n896) );
  NAND2_X1 U161 ( .A1(\mem[2][3] ), .A2(n1195), .ZN(n1191) );
  OAI21_X1 U162 ( .B1(n629), .B2(n1195), .A(n1190), .ZN(n895) );
  NAND2_X1 U163 ( .A1(\mem[2][4] ), .A2(n1195), .ZN(n1190) );
  OAI21_X1 U164 ( .B1(n630), .B2(n1195), .A(n1189), .ZN(n894) );
  NAND2_X1 U165 ( .A1(\mem[2][5] ), .A2(n1195), .ZN(n1189) );
  OAI21_X1 U166 ( .B1(n631), .B2(n1195), .A(n1188), .ZN(n893) );
  NAND2_X1 U167 ( .A1(\mem[2][6] ), .A2(n1195), .ZN(n1188) );
  OAI21_X1 U168 ( .B1(n632), .B2(n1195), .A(n1187), .ZN(n892) );
  NAND2_X1 U169 ( .A1(\mem[2][7] ), .A2(n1195), .ZN(n1187) );
  OAI21_X1 U170 ( .B1(n625), .B2(n1185), .A(n1184), .ZN(n891) );
  NAND2_X1 U171 ( .A1(\mem[3][0] ), .A2(n1185), .ZN(n1184) );
  OAI21_X1 U172 ( .B1(n626), .B2(n1185), .A(n1183), .ZN(n890) );
  NAND2_X1 U173 ( .A1(\mem[3][1] ), .A2(n1185), .ZN(n1183) );
  OAI21_X1 U174 ( .B1(n627), .B2(n1185), .A(n1182), .ZN(n889) );
  NAND2_X1 U175 ( .A1(\mem[3][2] ), .A2(n1185), .ZN(n1182) );
  OAI21_X1 U176 ( .B1(n628), .B2(n1185), .A(n1181), .ZN(n888) );
  NAND2_X1 U177 ( .A1(\mem[3][3] ), .A2(n1185), .ZN(n1181) );
  OAI21_X1 U178 ( .B1(n629), .B2(n1185), .A(n1180), .ZN(n887) );
  NAND2_X1 U179 ( .A1(\mem[3][4] ), .A2(n1185), .ZN(n1180) );
  OAI21_X1 U180 ( .B1(n630), .B2(n1185), .A(n1179), .ZN(n886) );
  NAND2_X1 U181 ( .A1(\mem[3][5] ), .A2(n1185), .ZN(n1179) );
  OAI21_X1 U182 ( .B1(n631), .B2(n1185), .A(n1178), .ZN(n885) );
  NAND2_X1 U183 ( .A1(\mem[3][6] ), .A2(n1185), .ZN(n1178) );
  OAI21_X1 U184 ( .B1(n632), .B2(n1185), .A(n1177), .ZN(n884) );
  NAND2_X1 U185 ( .A1(\mem[3][7] ), .A2(n1185), .ZN(n1177) );
  OAI21_X1 U186 ( .B1(n625), .B2(n1165), .A(n1164), .ZN(n875) );
  NAND2_X1 U187 ( .A1(\mem[5][0] ), .A2(n1165), .ZN(n1164) );
  OAI21_X1 U188 ( .B1(n626), .B2(n1165), .A(n1163), .ZN(n874) );
  NAND2_X1 U189 ( .A1(\mem[5][1] ), .A2(n1165), .ZN(n1163) );
  OAI21_X1 U190 ( .B1(n627), .B2(n1165), .A(n1162), .ZN(n873) );
  NAND2_X1 U191 ( .A1(\mem[5][2] ), .A2(n1165), .ZN(n1162) );
  OAI21_X1 U192 ( .B1(n628), .B2(n1165), .A(n1161), .ZN(n872) );
  NAND2_X1 U193 ( .A1(\mem[5][3] ), .A2(n1165), .ZN(n1161) );
  OAI21_X1 U194 ( .B1(n629), .B2(n1165), .A(n1160), .ZN(n871) );
  NAND2_X1 U195 ( .A1(\mem[5][4] ), .A2(n1165), .ZN(n1160) );
  OAI21_X1 U196 ( .B1(n630), .B2(n1165), .A(n1159), .ZN(n870) );
  NAND2_X1 U197 ( .A1(\mem[5][5] ), .A2(n1165), .ZN(n1159) );
  OAI21_X1 U198 ( .B1(n631), .B2(n1165), .A(n1158), .ZN(n869) );
  NAND2_X1 U199 ( .A1(\mem[5][6] ), .A2(n1165), .ZN(n1158) );
  OAI21_X1 U200 ( .B1(n632), .B2(n1165), .A(n1157), .ZN(n868) );
  NAND2_X1 U201 ( .A1(\mem[5][7] ), .A2(n1165), .ZN(n1157) );
  OAI21_X1 U202 ( .B1(n1216), .B2(n625), .A(n1215), .ZN(n915) );
  NAND2_X1 U203 ( .A1(\mem[0][0] ), .A2(n1216), .ZN(n1215) );
  OAI21_X1 U204 ( .B1(n1216), .B2(n626), .A(n1214), .ZN(n914) );
  NAND2_X1 U205 ( .A1(\mem[0][1] ), .A2(n1216), .ZN(n1214) );
  OAI21_X1 U206 ( .B1(n1216), .B2(n627), .A(n1213), .ZN(n913) );
  NAND2_X1 U207 ( .A1(\mem[0][2] ), .A2(n1216), .ZN(n1213) );
  OAI21_X1 U208 ( .B1(n1216), .B2(n628), .A(n1212), .ZN(n912) );
  NAND2_X1 U209 ( .A1(\mem[0][3] ), .A2(n1216), .ZN(n1212) );
  OAI21_X1 U210 ( .B1(n1216), .B2(n629), .A(n1211), .ZN(n911) );
  NAND2_X1 U211 ( .A1(\mem[0][4] ), .A2(n1216), .ZN(n1211) );
  OAI21_X1 U212 ( .B1(n1216), .B2(n630), .A(n1210), .ZN(n910) );
  NAND2_X1 U213 ( .A1(\mem[0][5] ), .A2(n1216), .ZN(n1210) );
  OAI21_X1 U214 ( .B1(n1216), .B2(n631), .A(n1209), .ZN(n909) );
  NAND2_X1 U215 ( .A1(\mem[0][6] ), .A2(n1216), .ZN(n1209) );
  OAI21_X1 U216 ( .B1(n1216), .B2(n632), .A(n1208), .ZN(n908) );
  NAND2_X1 U217 ( .A1(\mem[0][7] ), .A2(n1216), .ZN(n1208) );
  INV_X1 U218 ( .A(n1134), .ZN(n824) );
  AOI22_X1 U219 ( .A1(data_in[0]), .A2(n848), .B1(n1133), .B2(\mem[8][0] ), 
        .ZN(n1134) );
  INV_X1 U220 ( .A(n1132), .ZN(n823) );
  AOI22_X1 U221 ( .A1(data_in[1]), .A2(n848), .B1(n1133), .B2(\mem[8][1] ), 
        .ZN(n1132) );
  INV_X1 U222 ( .A(n1131), .ZN(n822) );
  AOI22_X1 U223 ( .A1(data_in[2]), .A2(n848), .B1(n1133), .B2(\mem[8][2] ), 
        .ZN(n1131) );
  INV_X1 U224 ( .A(n1130), .ZN(n821) );
  AOI22_X1 U225 ( .A1(data_in[3]), .A2(n848), .B1(n1133), .B2(\mem[8][3] ), 
        .ZN(n1130) );
  INV_X1 U226 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U227 ( .A1(data_in[4]), .A2(n848), .B1(n1133), .B2(\mem[8][4] ), 
        .ZN(n1129) );
  INV_X1 U228 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U229 ( .A1(data_in[5]), .A2(n848), .B1(n1133), .B2(\mem[8][5] ), 
        .ZN(n1128) );
  INV_X1 U230 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U231 ( .A1(data_in[6]), .A2(n848), .B1(n1133), .B2(\mem[8][6] ), 
        .ZN(n1127) );
  INV_X1 U232 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n848), .B1(n1133), .B2(\mem[8][7] ), 
        .ZN(n1126) );
  INV_X1 U234 ( .A(n1124), .ZN(n816) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n847), .B1(n1123), .B2(\mem[9][0] ), 
        .ZN(n1124) );
  INV_X1 U236 ( .A(n1122), .ZN(n815) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n847), .B1(n1123), .B2(\mem[9][1] ), 
        .ZN(n1122) );
  INV_X1 U238 ( .A(n1121), .ZN(n814) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n847), .B1(n1123), .B2(\mem[9][2] ), 
        .ZN(n1121) );
  INV_X1 U240 ( .A(n1120), .ZN(n813) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n847), .B1(n1123), .B2(\mem[9][3] ), 
        .ZN(n1120) );
  INV_X1 U242 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n847), .B1(n1123), .B2(\mem[9][4] ), 
        .ZN(n1119) );
  INV_X1 U244 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n847), .B1(n1123), .B2(\mem[9][5] ), 
        .ZN(n1118) );
  INV_X1 U246 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n847), .B1(n1123), .B2(\mem[9][6] ), 
        .ZN(n1117) );
  INV_X1 U248 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n847), .B1(n1123), .B2(\mem[9][7] ), 
        .ZN(n1116) );
  INV_X1 U250 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n846), .B1(n1114), .B2(\mem[10][0] ), 
        .ZN(n1115) );
  INV_X1 U252 ( .A(n1113), .ZN(n807) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n846), .B1(n1114), .B2(\mem[10][1] ), 
        .ZN(n1113) );
  INV_X1 U254 ( .A(n1112), .ZN(n806) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n846), .B1(n1114), .B2(\mem[10][2] ), 
        .ZN(n1112) );
  INV_X1 U256 ( .A(n1111), .ZN(n805) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n846), .B1(n1114), .B2(\mem[10][3] ), 
        .ZN(n1111) );
  INV_X1 U258 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n846), .B1(n1114), .B2(\mem[10][4] ), 
        .ZN(n1110) );
  INV_X1 U260 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n846), .B1(n1114), .B2(\mem[10][5] ), 
        .ZN(n1109) );
  INV_X1 U262 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n846), .B1(n1114), .B2(\mem[10][6] ), 
        .ZN(n1108) );
  INV_X1 U264 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n846), .B1(n1114), .B2(\mem[10][7] ), 
        .ZN(n1107) );
  INV_X1 U266 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n845), .B1(n1105), .B2(\mem[11][0] ), 
        .ZN(n1106) );
  INV_X1 U268 ( .A(n1104), .ZN(n799) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n845), .B1(n1105), .B2(\mem[11][1] ), 
        .ZN(n1104) );
  INV_X1 U270 ( .A(n1103), .ZN(n798) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n845), .B1(n1105), .B2(\mem[11][2] ), 
        .ZN(n1103) );
  INV_X1 U272 ( .A(n1102), .ZN(n797) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n845), .B1(n1105), .B2(\mem[11][3] ), 
        .ZN(n1102) );
  INV_X1 U274 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n845), .B1(n1105), .B2(\mem[11][4] ), 
        .ZN(n1101) );
  INV_X1 U276 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n845), .B1(n1105), .B2(\mem[11][5] ), 
        .ZN(n1100) );
  INV_X1 U278 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n845), .B1(n1105), .B2(\mem[11][6] ), 
        .ZN(n1099) );
  INV_X1 U280 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n845), .B1(n1105), .B2(\mem[11][7] ), 
        .ZN(n1098) );
  INV_X1 U282 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n844), .B1(n1096), .B2(\mem[12][0] ), 
        .ZN(n1097) );
  INV_X1 U284 ( .A(n1095), .ZN(n791) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n844), .B1(n1096), .B2(\mem[12][1] ), 
        .ZN(n1095) );
  INV_X1 U286 ( .A(n1094), .ZN(n790) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n844), .B1(n1096), .B2(\mem[12][2] ), 
        .ZN(n1094) );
  INV_X1 U288 ( .A(n1093), .ZN(n789) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n844), .B1(n1096), .B2(\mem[12][3] ), 
        .ZN(n1093) );
  INV_X1 U290 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n844), .B1(n1096), .B2(\mem[12][4] ), 
        .ZN(n1092) );
  INV_X1 U292 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n844), .B1(n1096), .B2(\mem[12][5] ), 
        .ZN(n1091) );
  INV_X1 U294 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n844), .B1(n1096), .B2(\mem[12][6] ), 
        .ZN(n1090) );
  INV_X1 U296 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n844), .B1(n1096), .B2(\mem[12][7] ), 
        .ZN(n1089) );
  INV_X1 U298 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n843), .B1(n1087), .B2(\mem[13][0] ), 
        .ZN(n1088) );
  INV_X1 U300 ( .A(n1086), .ZN(n783) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n843), .B1(n1087), .B2(\mem[13][1] ), 
        .ZN(n1086) );
  INV_X1 U302 ( .A(n1085), .ZN(n782) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n843), .B1(n1087), .B2(\mem[13][2] ), 
        .ZN(n1085) );
  INV_X1 U304 ( .A(n1084), .ZN(n781) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n843), .B1(n1087), .B2(\mem[13][3] ), 
        .ZN(n1084) );
  INV_X1 U306 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n843), .B1(n1087), .B2(\mem[13][4] ), 
        .ZN(n1083) );
  INV_X1 U308 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n843), .B1(n1087), .B2(\mem[13][5] ), 
        .ZN(n1082) );
  INV_X1 U310 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n843), .B1(n1087), .B2(\mem[13][6] ), 
        .ZN(n1081) );
  INV_X1 U312 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n843), .B1(n1087), .B2(\mem[13][7] ), 
        .ZN(n1080) );
  INV_X1 U314 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n842), .B1(n1078), .B2(\mem[14][0] ), 
        .ZN(n1079) );
  INV_X1 U316 ( .A(n1077), .ZN(n775) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n842), .B1(n1078), .B2(\mem[14][1] ), 
        .ZN(n1077) );
  INV_X1 U318 ( .A(n1076), .ZN(n774) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n842), .B1(n1078), .B2(\mem[14][2] ), 
        .ZN(n1076) );
  INV_X1 U320 ( .A(n1075), .ZN(n773) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n842), .B1(n1078), .B2(\mem[14][3] ), 
        .ZN(n1075) );
  INV_X1 U322 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n842), .B1(n1078), .B2(\mem[14][4] ), 
        .ZN(n1074) );
  INV_X1 U324 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n842), .B1(n1078), .B2(\mem[14][5] ), 
        .ZN(n1073) );
  INV_X1 U326 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n842), .B1(n1078), .B2(\mem[14][6] ), 
        .ZN(n1072) );
  INV_X1 U328 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n842), .B1(n1078), .B2(\mem[14][7] ), 
        .ZN(n1071) );
  INV_X1 U330 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U331 ( .A1(data_in[0]), .A2(n841), .B1(n1069), .B2(\mem[15][0] ), 
        .ZN(n1070) );
  INV_X1 U332 ( .A(n1068), .ZN(n767) );
  AOI22_X1 U333 ( .A1(data_in[1]), .A2(n841), .B1(n1069), .B2(\mem[15][1] ), 
        .ZN(n1068) );
  INV_X1 U334 ( .A(n1067), .ZN(n766) );
  AOI22_X1 U335 ( .A1(data_in[2]), .A2(n841), .B1(n1069), .B2(\mem[15][2] ), 
        .ZN(n1067) );
  INV_X1 U336 ( .A(n1066), .ZN(n765) );
  AOI22_X1 U337 ( .A1(data_in[3]), .A2(n841), .B1(n1069), .B2(\mem[15][3] ), 
        .ZN(n1066) );
  INV_X1 U338 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U339 ( .A1(data_in[4]), .A2(n841), .B1(n1069), .B2(\mem[15][4] ), 
        .ZN(n1065) );
  INV_X1 U340 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U341 ( .A1(data_in[5]), .A2(n841), .B1(n1069), .B2(\mem[15][5] ), 
        .ZN(n1064) );
  INV_X1 U342 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U343 ( .A1(data_in[6]), .A2(n841), .B1(n1069), .B2(\mem[15][6] ), 
        .ZN(n1063) );
  INV_X1 U344 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U345 ( .A1(data_in[7]), .A2(n841), .B1(n1069), .B2(\mem[15][7] ), 
        .ZN(n1062) );
  INV_X1 U346 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U347 ( .A1(data_in[0]), .A2(n840), .B1(n1060), .B2(\mem[16][0] ), 
        .ZN(n1061) );
  INV_X1 U348 ( .A(n1059), .ZN(n759) );
  AOI22_X1 U349 ( .A1(data_in[1]), .A2(n840), .B1(n1060), .B2(\mem[16][1] ), 
        .ZN(n1059) );
  INV_X1 U350 ( .A(n1058), .ZN(n758) );
  AOI22_X1 U351 ( .A1(data_in[2]), .A2(n840), .B1(n1060), .B2(\mem[16][2] ), 
        .ZN(n1058) );
  INV_X1 U352 ( .A(n1057), .ZN(n757) );
  AOI22_X1 U353 ( .A1(data_in[3]), .A2(n840), .B1(n1060), .B2(\mem[16][3] ), 
        .ZN(n1057) );
  INV_X1 U354 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U355 ( .A1(data_in[4]), .A2(n840), .B1(n1060), .B2(\mem[16][4] ), 
        .ZN(n1056) );
  INV_X1 U356 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U357 ( .A1(data_in[5]), .A2(n840), .B1(n1060), .B2(\mem[16][5] ), 
        .ZN(n1055) );
  INV_X1 U358 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U359 ( .A1(data_in[6]), .A2(n840), .B1(n1060), .B2(\mem[16][6] ), 
        .ZN(n1054) );
  INV_X1 U360 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U361 ( .A1(data_in[7]), .A2(n840), .B1(n1060), .B2(\mem[16][7] ), 
        .ZN(n1053) );
  INV_X1 U362 ( .A(n1051), .ZN(n752) );
  AOI22_X1 U363 ( .A1(data_in[0]), .A2(n839), .B1(n1050), .B2(\mem[17][0] ), 
        .ZN(n1051) );
  INV_X1 U364 ( .A(n1049), .ZN(n751) );
  AOI22_X1 U365 ( .A1(data_in[1]), .A2(n839), .B1(n1050), .B2(\mem[17][1] ), 
        .ZN(n1049) );
  INV_X1 U366 ( .A(n1048), .ZN(n750) );
  AOI22_X1 U367 ( .A1(data_in[2]), .A2(n839), .B1(n1050), .B2(\mem[17][2] ), 
        .ZN(n1048) );
  INV_X1 U368 ( .A(n1047), .ZN(n749) );
  AOI22_X1 U369 ( .A1(data_in[3]), .A2(n839), .B1(n1050), .B2(\mem[17][3] ), 
        .ZN(n1047) );
  INV_X1 U370 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U371 ( .A1(data_in[4]), .A2(n839), .B1(n1050), .B2(\mem[17][4] ), 
        .ZN(n1046) );
  INV_X1 U372 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U373 ( .A1(data_in[5]), .A2(n839), .B1(n1050), .B2(\mem[17][5] ), 
        .ZN(n1045) );
  INV_X1 U374 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U375 ( .A1(data_in[6]), .A2(n839), .B1(n1050), .B2(\mem[17][6] ), 
        .ZN(n1044) );
  INV_X1 U376 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U377 ( .A1(data_in[7]), .A2(n839), .B1(n1050), .B2(\mem[17][7] ), 
        .ZN(n1043) );
  INV_X1 U378 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U379 ( .A1(data_in[0]), .A2(n838), .B1(n1041), .B2(\mem[18][0] ), 
        .ZN(n1042) );
  INV_X1 U380 ( .A(n1040), .ZN(n743) );
  AOI22_X1 U381 ( .A1(data_in[1]), .A2(n838), .B1(n1041), .B2(\mem[18][1] ), 
        .ZN(n1040) );
  INV_X1 U382 ( .A(n1039), .ZN(n742) );
  AOI22_X1 U383 ( .A1(data_in[2]), .A2(n838), .B1(n1041), .B2(\mem[18][2] ), 
        .ZN(n1039) );
  INV_X1 U384 ( .A(n1038), .ZN(n741) );
  AOI22_X1 U385 ( .A1(data_in[3]), .A2(n838), .B1(n1041), .B2(\mem[18][3] ), 
        .ZN(n1038) );
  INV_X1 U386 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U387 ( .A1(data_in[4]), .A2(n838), .B1(n1041), .B2(\mem[18][4] ), 
        .ZN(n1037) );
  INV_X1 U388 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U389 ( .A1(data_in[5]), .A2(n838), .B1(n1041), .B2(\mem[18][5] ), 
        .ZN(n1036) );
  INV_X1 U390 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U391 ( .A1(data_in[6]), .A2(n838), .B1(n1041), .B2(\mem[18][6] ), 
        .ZN(n1035) );
  INV_X1 U392 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U393 ( .A1(data_in[7]), .A2(n838), .B1(n1041), .B2(\mem[18][7] ), 
        .ZN(n1034) );
  INV_X1 U394 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U395 ( .A1(data_in[0]), .A2(n837), .B1(n1032), .B2(\mem[19][0] ), 
        .ZN(n1033) );
  INV_X1 U396 ( .A(n1031), .ZN(n735) );
  AOI22_X1 U397 ( .A1(data_in[1]), .A2(n837), .B1(n1032), .B2(\mem[19][1] ), 
        .ZN(n1031) );
  INV_X1 U398 ( .A(n1030), .ZN(n734) );
  AOI22_X1 U399 ( .A1(data_in[2]), .A2(n837), .B1(n1032), .B2(\mem[19][2] ), 
        .ZN(n1030) );
  INV_X1 U400 ( .A(n1029), .ZN(n733) );
  AOI22_X1 U401 ( .A1(data_in[3]), .A2(n837), .B1(n1032), .B2(\mem[19][3] ), 
        .ZN(n1029) );
  INV_X1 U402 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U403 ( .A1(data_in[4]), .A2(n837), .B1(n1032), .B2(\mem[19][4] ), 
        .ZN(n1028) );
  INV_X1 U404 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U405 ( .A1(data_in[5]), .A2(n837), .B1(n1032), .B2(\mem[19][5] ), 
        .ZN(n1027) );
  INV_X1 U406 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U407 ( .A1(data_in[6]), .A2(n837), .B1(n1032), .B2(\mem[19][6] ), 
        .ZN(n1026) );
  INV_X1 U408 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U409 ( .A1(data_in[7]), .A2(n837), .B1(n1032), .B2(\mem[19][7] ), 
        .ZN(n1025) );
  INV_X1 U410 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U411 ( .A1(data_in[0]), .A2(n836), .B1(n1023), .B2(\mem[20][0] ), 
        .ZN(n1024) );
  INV_X1 U412 ( .A(n1022), .ZN(n727) );
  AOI22_X1 U413 ( .A1(data_in[1]), .A2(n836), .B1(n1023), .B2(\mem[20][1] ), 
        .ZN(n1022) );
  INV_X1 U414 ( .A(n1021), .ZN(n726) );
  AOI22_X1 U415 ( .A1(data_in[2]), .A2(n836), .B1(n1023), .B2(\mem[20][2] ), 
        .ZN(n1021) );
  INV_X1 U416 ( .A(n1020), .ZN(n725) );
  AOI22_X1 U417 ( .A1(data_in[3]), .A2(n836), .B1(n1023), .B2(\mem[20][3] ), 
        .ZN(n1020) );
  INV_X1 U418 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U419 ( .A1(data_in[4]), .A2(n836), .B1(n1023), .B2(\mem[20][4] ), 
        .ZN(n1019) );
  INV_X1 U420 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U421 ( .A1(data_in[5]), .A2(n836), .B1(n1023), .B2(\mem[20][5] ), 
        .ZN(n1018) );
  INV_X1 U422 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U423 ( .A1(data_in[6]), .A2(n836), .B1(n1023), .B2(\mem[20][6] ), 
        .ZN(n1017) );
  INV_X1 U424 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U425 ( .A1(data_in[7]), .A2(n836), .B1(n1023), .B2(\mem[20][7] ), 
        .ZN(n1016) );
  INV_X1 U426 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U427 ( .A1(data_in[0]), .A2(n835), .B1(n1014), .B2(\mem[21][0] ), 
        .ZN(n1015) );
  INV_X1 U428 ( .A(n1013), .ZN(n719) );
  AOI22_X1 U429 ( .A1(data_in[1]), .A2(n835), .B1(n1014), .B2(\mem[21][1] ), 
        .ZN(n1013) );
  INV_X1 U430 ( .A(n1012), .ZN(n718) );
  AOI22_X1 U431 ( .A1(data_in[2]), .A2(n835), .B1(n1014), .B2(\mem[21][2] ), 
        .ZN(n1012) );
  INV_X1 U432 ( .A(n1011), .ZN(n717) );
  AOI22_X1 U433 ( .A1(data_in[3]), .A2(n835), .B1(n1014), .B2(\mem[21][3] ), 
        .ZN(n1011) );
  INV_X1 U434 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U435 ( .A1(data_in[4]), .A2(n835), .B1(n1014), .B2(\mem[21][4] ), 
        .ZN(n1010) );
  INV_X1 U436 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U437 ( .A1(data_in[5]), .A2(n835), .B1(n1014), .B2(\mem[21][5] ), 
        .ZN(n1009) );
  INV_X1 U438 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U439 ( .A1(data_in[6]), .A2(n835), .B1(n1014), .B2(\mem[21][6] ), 
        .ZN(n1008) );
  INV_X1 U440 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U441 ( .A1(data_in[7]), .A2(n835), .B1(n1014), .B2(\mem[21][7] ), 
        .ZN(n1007) );
  INV_X1 U442 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U443 ( .A1(data_in[0]), .A2(n834), .B1(n1005), .B2(\mem[22][0] ), 
        .ZN(n1006) );
  INV_X1 U444 ( .A(n1004), .ZN(n711) );
  AOI22_X1 U445 ( .A1(data_in[1]), .A2(n834), .B1(n1005), .B2(\mem[22][1] ), 
        .ZN(n1004) );
  INV_X1 U446 ( .A(n1003), .ZN(n710) );
  AOI22_X1 U447 ( .A1(data_in[2]), .A2(n834), .B1(n1005), .B2(\mem[22][2] ), 
        .ZN(n1003) );
  INV_X1 U448 ( .A(n1002), .ZN(n709) );
  AOI22_X1 U449 ( .A1(data_in[3]), .A2(n834), .B1(n1005), .B2(\mem[22][3] ), 
        .ZN(n1002) );
  INV_X1 U450 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U451 ( .A1(data_in[4]), .A2(n834), .B1(n1005), .B2(\mem[22][4] ), 
        .ZN(n1001) );
  INV_X1 U452 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U453 ( .A1(data_in[5]), .A2(n834), .B1(n1005), .B2(\mem[22][5] ), 
        .ZN(n1000) );
  INV_X1 U454 ( .A(n999), .ZN(n706) );
  AOI22_X1 U455 ( .A1(data_in[6]), .A2(n834), .B1(n1005), .B2(\mem[22][6] ), 
        .ZN(n999) );
  INV_X1 U456 ( .A(n998), .ZN(n705) );
  AOI22_X1 U457 ( .A1(data_in[7]), .A2(n834), .B1(n1005), .B2(\mem[22][7] ), 
        .ZN(n998) );
  INV_X1 U458 ( .A(n997), .ZN(n704) );
  AOI22_X1 U459 ( .A1(data_in[0]), .A2(n833), .B1(n996), .B2(\mem[23][0] ), 
        .ZN(n997) );
  INV_X1 U460 ( .A(n995), .ZN(n703) );
  AOI22_X1 U461 ( .A1(data_in[1]), .A2(n833), .B1(n996), .B2(\mem[23][1] ), 
        .ZN(n995) );
  INV_X1 U462 ( .A(n994), .ZN(n702) );
  AOI22_X1 U463 ( .A1(data_in[2]), .A2(n833), .B1(n996), .B2(\mem[23][2] ), 
        .ZN(n994) );
  INV_X1 U464 ( .A(n993), .ZN(n701) );
  AOI22_X1 U465 ( .A1(data_in[3]), .A2(n833), .B1(n996), .B2(\mem[23][3] ), 
        .ZN(n993) );
  INV_X1 U466 ( .A(n992), .ZN(n700) );
  AOI22_X1 U467 ( .A1(data_in[4]), .A2(n833), .B1(n996), .B2(\mem[23][4] ), 
        .ZN(n992) );
  INV_X1 U468 ( .A(n991), .ZN(n699) );
  AOI22_X1 U469 ( .A1(data_in[5]), .A2(n833), .B1(n996), .B2(\mem[23][5] ), 
        .ZN(n991) );
  INV_X1 U470 ( .A(n990), .ZN(n698) );
  AOI22_X1 U471 ( .A1(data_in[6]), .A2(n833), .B1(n996), .B2(\mem[23][6] ), 
        .ZN(n990) );
  INV_X1 U472 ( .A(n989), .ZN(n697) );
  AOI22_X1 U473 ( .A1(data_in[7]), .A2(n833), .B1(n996), .B2(\mem[23][7] ), 
        .ZN(n989) );
  INV_X1 U474 ( .A(n988), .ZN(n696) );
  AOI22_X1 U475 ( .A1(data_in[0]), .A2(n832), .B1(n987), .B2(\mem[24][0] ), 
        .ZN(n988) );
  INV_X1 U476 ( .A(n986), .ZN(n695) );
  AOI22_X1 U477 ( .A1(data_in[1]), .A2(n832), .B1(n987), .B2(\mem[24][1] ), 
        .ZN(n986) );
  INV_X1 U478 ( .A(n985), .ZN(n694) );
  AOI22_X1 U479 ( .A1(data_in[2]), .A2(n832), .B1(n987), .B2(\mem[24][2] ), 
        .ZN(n985) );
  INV_X1 U480 ( .A(n984), .ZN(n693) );
  AOI22_X1 U481 ( .A1(data_in[3]), .A2(n832), .B1(n987), .B2(\mem[24][3] ), 
        .ZN(n984) );
  INV_X1 U482 ( .A(n983), .ZN(n692) );
  AOI22_X1 U483 ( .A1(data_in[4]), .A2(n832), .B1(n987), .B2(\mem[24][4] ), 
        .ZN(n983) );
  INV_X1 U484 ( .A(n982), .ZN(n691) );
  AOI22_X1 U485 ( .A1(data_in[5]), .A2(n832), .B1(n987), .B2(\mem[24][5] ), 
        .ZN(n982) );
  INV_X1 U486 ( .A(n981), .ZN(n690) );
  AOI22_X1 U487 ( .A1(data_in[6]), .A2(n832), .B1(n987), .B2(\mem[24][6] ), 
        .ZN(n981) );
  INV_X1 U488 ( .A(n980), .ZN(n689) );
  AOI22_X1 U489 ( .A1(data_in[7]), .A2(n832), .B1(n987), .B2(\mem[24][7] ), 
        .ZN(n980) );
  INV_X1 U490 ( .A(n978), .ZN(n688) );
  AOI22_X1 U491 ( .A1(data_in[0]), .A2(n831), .B1(n977), .B2(\mem[25][0] ), 
        .ZN(n978) );
  INV_X1 U492 ( .A(n976), .ZN(n687) );
  AOI22_X1 U493 ( .A1(data_in[1]), .A2(n831), .B1(n977), .B2(\mem[25][1] ), 
        .ZN(n976) );
  INV_X1 U494 ( .A(n975), .ZN(n686) );
  AOI22_X1 U495 ( .A1(data_in[2]), .A2(n831), .B1(n977), .B2(\mem[25][2] ), 
        .ZN(n975) );
  INV_X1 U496 ( .A(n974), .ZN(n685) );
  AOI22_X1 U497 ( .A1(data_in[3]), .A2(n831), .B1(n977), .B2(\mem[25][3] ), 
        .ZN(n974) );
  INV_X1 U498 ( .A(n973), .ZN(n684) );
  AOI22_X1 U499 ( .A1(data_in[4]), .A2(n831), .B1(n977), .B2(\mem[25][4] ), 
        .ZN(n973) );
  INV_X1 U500 ( .A(n972), .ZN(n683) );
  AOI22_X1 U501 ( .A1(data_in[5]), .A2(n831), .B1(n977), .B2(\mem[25][5] ), 
        .ZN(n972) );
  INV_X1 U502 ( .A(n971), .ZN(n682) );
  AOI22_X1 U503 ( .A1(data_in[6]), .A2(n831), .B1(n977), .B2(\mem[25][6] ), 
        .ZN(n971) );
  INV_X1 U504 ( .A(n970), .ZN(n681) );
  AOI22_X1 U505 ( .A1(data_in[7]), .A2(n831), .B1(n977), .B2(\mem[25][7] ), 
        .ZN(n970) );
  INV_X1 U506 ( .A(n969), .ZN(n680) );
  AOI22_X1 U507 ( .A1(data_in[0]), .A2(n830), .B1(n968), .B2(\mem[26][0] ), 
        .ZN(n969) );
  INV_X1 U508 ( .A(n967), .ZN(n679) );
  AOI22_X1 U509 ( .A1(data_in[1]), .A2(n830), .B1(n968), .B2(\mem[26][1] ), 
        .ZN(n967) );
  INV_X1 U510 ( .A(n966), .ZN(n678) );
  AOI22_X1 U511 ( .A1(data_in[2]), .A2(n830), .B1(n968), .B2(\mem[26][2] ), 
        .ZN(n966) );
  INV_X1 U512 ( .A(n965), .ZN(n677) );
  AOI22_X1 U513 ( .A1(data_in[3]), .A2(n830), .B1(n968), .B2(\mem[26][3] ), 
        .ZN(n965) );
  INV_X1 U514 ( .A(n964), .ZN(n676) );
  AOI22_X1 U515 ( .A1(data_in[4]), .A2(n830), .B1(n968), .B2(\mem[26][4] ), 
        .ZN(n964) );
  INV_X1 U516 ( .A(n963), .ZN(n675) );
  AOI22_X1 U517 ( .A1(data_in[5]), .A2(n830), .B1(n968), .B2(\mem[26][5] ), 
        .ZN(n963) );
  INV_X1 U518 ( .A(n962), .ZN(n674) );
  AOI22_X1 U519 ( .A1(data_in[6]), .A2(n830), .B1(n968), .B2(\mem[26][6] ), 
        .ZN(n962) );
  INV_X1 U520 ( .A(n961), .ZN(n673) );
  AOI22_X1 U521 ( .A1(data_in[7]), .A2(n830), .B1(n968), .B2(\mem[26][7] ), 
        .ZN(n961) );
  INV_X1 U522 ( .A(n960), .ZN(n672) );
  AOI22_X1 U523 ( .A1(data_in[0]), .A2(n829), .B1(n959), .B2(\mem[27][0] ), 
        .ZN(n960) );
  INV_X1 U524 ( .A(n958), .ZN(n671) );
  AOI22_X1 U525 ( .A1(data_in[1]), .A2(n829), .B1(n959), .B2(\mem[27][1] ), 
        .ZN(n958) );
  INV_X1 U526 ( .A(n957), .ZN(n670) );
  AOI22_X1 U527 ( .A1(data_in[2]), .A2(n829), .B1(n959), .B2(\mem[27][2] ), 
        .ZN(n957) );
  INV_X1 U528 ( .A(n956), .ZN(n669) );
  AOI22_X1 U529 ( .A1(data_in[3]), .A2(n829), .B1(n959), .B2(\mem[27][3] ), 
        .ZN(n956) );
  INV_X1 U530 ( .A(n955), .ZN(n668) );
  AOI22_X1 U531 ( .A1(data_in[4]), .A2(n829), .B1(n959), .B2(\mem[27][4] ), 
        .ZN(n955) );
  INV_X1 U532 ( .A(n954), .ZN(n667) );
  AOI22_X1 U533 ( .A1(data_in[5]), .A2(n829), .B1(n959), .B2(\mem[27][5] ), 
        .ZN(n954) );
  INV_X1 U534 ( .A(n953), .ZN(n666) );
  AOI22_X1 U535 ( .A1(data_in[6]), .A2(n829), .B1(n959), .B2(\mem[27][6] ), 
        .ZN(n953) );
  INV_X1 U536 ( .A(n952), .ZN(n665) );
  AOI22_X1 U537 ( .A1(data_in[7]), .A2(n829), .B1(n959), .B2(\mem[27][7] ), 
        .ZN(n952) );
  INV_X1 U538 ( .A(n951), .ZN(n664) );
  AOI22_X1 U539 ( .A1(data_in[0]), .A2(n828), .B1(n950), .B2(\mem[28][0] ), 
        .ZN(n951) );
  INV_X1 U540 ( .A(n949), .ZN(n663) );
  AOI22_X1 U541 ( .A1(data_in[1]), .A2(n828), .B1(n950), .B2(\mem[28][1] ), 
        .ZN(n949) );
  INV_X1 U542 ( .A(n948), .ZN(n662) );
  AOI22_X1 U543 ( .A1(data_in[2]), .A2(n828), .B1(n950), .B2(\mem[28][2] ), 
        .ZN(n948) );
  INV_X1 U544 ( .A(n947), .ZN(n661) );
  AOI22_X1 U545 ( .A1(data_in[3]), .A2(n828), .B1(n950), .B2(\mem[28][3] ), 
        .ZN(n947) );
  INV_X1 U546 ( .A(n946), .ZN(n660) );
  AOI22_X1 U547 ( .A1(data_in[4]), .A2(n828), .B1(n950), .B2(\mem[28][4] ), 
        .ZN(n946) );
  INV_X1 U548 ( .A(n945), .ZN(n659) );
  AOI22_X1 U549 ( .A1(data_in[5]), .A2(n828), .B1(n950), .B2(\mem[28][5] ), 
        .ZN(n945) );
  INV_X1 U550 ( .A(n944), .ZN(n658) );
  AOI22_X1 U551 ( .A1(data_in[6]), .A2(n828), .B1(n950), .B2(\mem[28][6] ), 
        .ZN(n944) );
  INV_X1 U552 ( .A(n943), .ZN(n657) );
  AOI22_X1 U553 ( .A1(data_in[7]), .A2(n828), .B1(n950), .B2(\mem[28][7] ), 
        .ZN(n943) );
  INV_X1 U554 ( .A(n942), .ZN(n656) );
  AOI22_X1 U555 ( .A1(data_in[0]), .A2(n827), .B1(n941), .B2(\mem[29][0] ), 
        .ZN(n942) );
  INV_X1 U556 ( .A(n940), .ZN(n655) );
  AOI22_X1 U557 ( .A1(data_in[1]), .A2(n827), .B1(n941), .B2(\mem[29][1] ), 
        .ZN(n940) );
  INV_X1 U558 ( .A(n939), .ZN(n654) );
  AOI22_X1 U559 ( .A1(data_in[2]), .A2(n827), .B1(n941), .B2(\mem[29][2] ), 
        .ZN(n939) );
  INV_X1 U560 ( .A(n938), .ZN(n653) );
  AOI22_X1 U561 ( .A1(data_in[3]), .A2(n827), .B1(n941), .B2(\mem[29][3] ), 
        .ZN(n938) );
  INV_X1 U562 ( .A(n937), .ZN(n652) );
  AOI22_X1 U563 ( .A1(data_in[4]), .A2(n827), .B1(n941), .B2(\mem[29][4] ), 
        .ZN(n937) );
  INV_X1 U564 ( .A(n936), .ZN(n651) );
  AOI22_X1 U565 ( .A1(data_in[5]), .A2(n827), .B1(n941), .B2(\mem[29][5] ), 
        .ZN(n936) );
  INV_X1 U566 ( .A(n935), .ZN(n650) );
  AOI22_X1 U567 ( .A1(data_in[6]), .A2(n827), .B1(n941), .B2(\mem[29][6] ), 
        .ZN(n935) );
  INV_X1 U568 ( .A(n934), .ZN(n649) );
  AOI22_X1 U569 ( .A1(data_in[7]), .A2(n827), .B1(n941), .B2(\mem[29][7] ), 
        .ZN(n934) );
  INV_X1 U570 ( .A(n933), .ZN(n648) );
  AOI22_X1 U571 ( .A1(data_in[0]), .A2(n826), .B1(n932), .B2(\mem[30][0] ), 
        .ZN(n933) );
  INV_X1 U572 ( .A(n931), .ZN(n647) );
  AOI22_X1 U573 ( .A1(data_in[1]), .A2(n826), .B1(n932), .B2(\mem[30][1] ), 
        .ZN(n931) );
  INV_X1 U574 ( .A(n930), .ZN(n646) );
  AOI22_X1 U575 ( .A1(data_in[2]), .A2(n826), .B1(n932), .B2(\mem[30][2] ), 
        .ZN(n930) );
  INV_X1 U576 ( .A(n929), .ZN(n645) );
  AOI22_X1 U577 ( .A1(data_in[3]), .A2(n826), .B1(n932), .B2(\mem[30][3] ), 
        .ZN(n929) );
  INV_X1 U578 ( .A(n928), .ZN(n644) );
  AOI22_X1 U579 ( .A1(data_in[4]), .A2(n826), .B1(n932), .B2(\mem[30][4] ), 
        .ZN(n928) );
  INV_X1 U580 ( .A(n927), .ZN(n643) );
  AOI22_X1 U581 ( .A1(data_in[5]), .A2(n826), .B1(n932), .B2(\mem[30][5] ), 
        .ZN(n927) );
  INV_X1 U582 ( .A(n926), .ZN(n642) );
  AOI22_X1 U583 ( .A1(data_in[6]), .A2(n826), .B1(n932), .B2(\mem[30][6] ), 
        .ZN(n926) );
  INV_X1 U584 ( .A(n925), .ZN(n641) );
  AOI22_X1 U585 ( .A1(data_in[7]), .A2(n826), .B1(n932), .B2(\mem[30][7] ), 
        .ZN(n925) );
  INV_X1 U586 ( .A(n924), .ZN(n640) );
  AOI22_X1 U587 ( .A1(data_in[0]), .A2(n825), .B1(n923), .B2(\mem[31][0] ), 
        .ZN(n924) );
  INV_X1 U588 ( .A(n922), .ZN(n639) );
  AOI22_X1 U589 ( .A1(data_in[1]), .A2(n825), .B1(n923), .B2(\mem[31][1] ), 
        .ZN(n922) );
  INV_X1 U590 ( .A(n921), .ZN(n638) );
  AOI22_X1 U591 ( .A1(data_in[2]), .A2(n825), .B1(n923), .B2(\mem[31][2] ), 
        .ZN(n921) );
  INV_X1 U592 ( .A(n920), .ZN(n637) );
  AOI22_X1 U593 ( .A1(data_in[3]), .A2(n825), .B1(n923), .B2(\mem[31][3] ), 
        .ZN(n920) );
  INV_X1 U594 ( .A(n919), .ZN(n636) );
  AOI22_X1 U595 ( .A1(data_in[4]), .A2(n825), .B1(n923), .B2(\mem[31][4] ), 
        .ZN(n919) );
  INV_X1 U596 ( .A(n918), .ZN(n635) );
  AOI22_X1 U597 ( .A1(data_in[5]), .A2(n825), .B1(n923), .B2(\mem[31][5] ), 
        .ZN(n918) );
  INV_X1 U598 ( .A(n917), .ZN(n634) );
  AOI22_X1 U599 ( .A1(data_in[6]), .A2(n825), .B1(n923), .B2(\mem[31][6] ), 
        .ZN(n917) );
  INV_X1 U600 ( .A(n916), .ZN(n633) );
  AOI22_X1 U601 ( .A1(data_in[7]), .A2(n825), .B1(n923), .B2(\mem[31][7] ), 
        .ZN(n916) );
  MUX2_X1 U602 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n613), .Z(n3) );
  MUX2_X1 U603 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n613), .Z(n4) );
  MUX2_X1 U604 ( .A(n4), .B(n3), .S(n610), .Z(n5) );
  MUX2_X1 U605 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n613), .Z(n6) );
  MUX2_X1 U606 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n613), .Z(n7) );
  MUX2_X1 U607 ( .A(n7), .B(n6), .S(n610), .Z(n8) );
  MUX2_X1 U608 ( .A(n8), .B(n5), .S(n608), .Z(n9) );
  MUX2_X1 U609 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n613), .Z(n10) );
  MUX2_X1 U610 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n613), .Z(n11) );
  MUX2_X1 U611 ( .A(n11), .B(n10), .S(n610), .Z(n12) );
  MUX2_X1 U612 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n613), .Z(n13) );
  MUX2_X1 U613 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n613), .Z(n14) );
  MUX2_X1 U614 ( .A(n14), .B(n13), .S(n610), .Z(n15) );
  MUX2_X1 U615 ( .A(n15), .B(n12), .S(N12), .Z(n16) );
  MUX2_X1 U616 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U617 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n614), .Z(n18) );
  MUX2_X1 U618 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n614), .Z(n19) );
  MUX2_X1 U619 ( .A(n19), .B(n18), .S(n611), .Z(n20) );
  MUX2_X1 U620 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n614), .Z(n21) );
  MUX2_X1 U621 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n614), .Z(n22) );
  MUX2_X1 U622 ( .A(n22), .B(n21), .S(n611), .Z(n23) );
  MUX2_X1 U623 ( .A(n23), .B(n20), .S(N12), .Z(n24) );
  MUX2_X1 U624 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n614), .Z(n25) );
  MUX2_X1 U625 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n614), .Z(n26) );
  MUX2_X1 U626 ( .A(n26), .B(n25), .S(n611), .Z(n27) );
  MUX2_X1 U627 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n614), .Z(n28) );
  MUX2_X1 U628 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n614), .Z(n29) );
  MUX2_X1 U629 ( .A(n29), .B(n28), .S(n611), .Z(n30) );
  MUX2_X1 U630 ( .A(n30), .B(n27), .S(n609), .Z(n31) );
  MUX2_X1 U631 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U632 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U633 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n614), .Z(n33) );
  MUX2_X1 U634 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n614), .Z(n34) );
  MUX2_X1 U635 ( .A(n34), .B(n33), .S(n611), .Z(n35) );
  MUX2_X1 U636 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n614), .Z(n36) );
  MUX2_X1 U637 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n614), .Z(n37) );
  MUX2_X1 U638 ( .A(n37), .B(n36), .S(n611), .Z(n38) );
  MUX2_X1 U639 ( .A(n38), .B(n35), .S(n609), .Z(n39) );
  MUX2_X1 U640 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n615), .Z(n40) );
  MUX2_X1 U641 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n615), .Z(n41) );
  MUX2_X1 U642 ( .A(n41), .B(n40), .S(n611), .Z(n42) );
  MUX2_X1 U643 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n615), .Z(n43) );
  MUX2_X1 U644 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n615), .Z(n44) );
  MUX2_X1 U645 ( .A(n44), .B(n43), .S(n611), .Z(n45) );
  MUX2_X1 U646 ( .A(n45), .B(n42), .S(N12), .Z(n46) );
  MUX2_X1 U647 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U648 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n615), .Z(n48) );
  MUX2_X1 U649 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n615), .Z(n49) );
  MUX2_X1 U650 ( .A(n49), .B(n48), .S(n611), .Z(n50) );
  MUX2_X1 U651 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n615), .Z(n51) );
  MUX2_X1 U652 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n615), .Z(n52) );
  MUX2_X1 U653 ( .A(n52), .B(n51), .S(n611), .Z(n53) );
  MUX2_X1 U654 ( .A(n53), .B(n50), .S(n608), .Z(n54) );
  MUX2_X1 U655 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n615), .Z(n55) );
  MUX2_X1 U656 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n615), .Z(n56) );
  MUX2_X1 U657 ( .A(n56), .B(n55), .S(n611), .Z(n57) );
  MUX2_X1 U658 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n615), .Z(n58) );
  MUX2_X1 U659 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n615), .Z(n59) );
  MUX2_X1 U660 ( .A(n59), .B(n58), .S(n611), .Z(n60) );
  MUX2_X1 U661 ( .A(n60), .B(n57), .S(n608), .Z(n61) );
  MUX2_X1 U662 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U663 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U664 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n616), .Z(n63) );
  MUX2_X1 U665 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n616), .Z(n64) );
  MUX2_X1 U666 ( .A(n64), .B(n63), .S(n612), .Z(n65) );
  MUX2_X1 U667 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n616), .Z(n66) );
  MUX2_X1 U668 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n616), .Z(n67) );
  MUX2_X1 U669 ( .A(n67), .B(n66), .S(n612), .Z(n68) );
  MUX2_X1 U670 ( .A(n68), .B(n65), .S(n608), .Z(n69) );
  MUX2_X1 U671 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n616), .Z(n70) );
  MUX2_X1 U672 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n616), .Z(n71) );
  MUX2_X1 U673 ( .A(n71), .B(n70), .S(n612), .Z(n72) );
  MUX2_X1 U674 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n616), .Z(n73) );
  MUX2_X1 U675 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n616), .Z(n74) );
  MUX2_X1 U676 ( .A(n74), .B(n73), .S(n612), .Z(n75) );
  MUX2_X1 U677 ( .A(n75), .B(n72), .S(n608), .Z(n76) );
  MUX2_X1 U678 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U679 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n616), .Z(n78) );
  MUX2_X1 U680 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n616), .Z(n79) );
  MUX2_X1 U681 ( .A(n79), .B(n78), .S(n612), .Z(n80) );
  MUX2_X1 U682 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n616), .Z(n81) );
  MUX2_X1 U683 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n616), .Z(n82) );
  MUX2_X1 U684 ( .A(n82), .B(n81), .S(n612), .Z(n83) );
  MUX2_X1 U685 ( .A(n83), .B(n80), .S(n608), .Z(n84) );
  MUX2_X1 U686 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n617), .Z(n85) );
  MUX2_X1 U687 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n617), .Z(n86) );
  MUX2_X1 U688 ( .A(n86), .B(n85), .S(n612), .Z(n87) );
  MUX2_X1 U689 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n617), .Z(n88) );
  MUX2_X1 U690 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n617), .Z(n89) );
  MUX2_X1 U691 ( .A(n89), .B(n88), .S(n612), .Z(n90) );
  MUX2_X1 U692 ( .A(n90), .B(n87), .S(n608), .Z(n91) );
  MUX2_X1 U693 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U694 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U695 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n617), .Z(n93) );
  MUX2_X1 U696 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n617), .Z(n94) );
  MUX2_X1 U697 ( .A(n94), .B(n93), .S(n612), .Z(n95) );
  MUX2_X1 U698 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n617), .Z(n96) );
  MUX2_X1 U699 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n617), .Z(n97) );
  MUX2_X1 U700 ( .A(n97), .B(n96), .S(n612), .Z(n98) );
  MUX2_X1 U701 ( .A(n98), .B(n95), .S(n608), .Z(n99) );
  MUX2_X1 U702 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n617), .Z(n100) );
  MUX2_X1 U703 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n617), .Z(n101) );
  MUX2_X1 U704 ( .A(n101), .B(n100), .S(n612), .Z(n102) );
  MUX2_X1 U705 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n617), .Z(n103) );
  MUX2_X1 U706 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n617), .Z(n104) );
  MUX2_X1 U707 ( .A(n104), .B(n103), .S(n612), .Z(n105) );
  MUX2_X1 U708 ( .A(n105), .B(n102), .S(n608), .Z(n106) );
  MUX2_X1 U709 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U710 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n618), .Z(n108) );
  MUX2_X1 U711 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n618), .Z(n109) );
  MUX2_X1 U712 ( .A(n109), .B(n108), .S(n611), .Z(n110) );
  MUX2_X1 U713 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n618), .Z(n111) );
  MUX2_X1 U714 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n618), .Z(n112) );
  MUX2_X1 U715 ( .A(n112), .B(n111), .S(n612), .Z(n113) );
  MUX2_X1 U716 ( .A(n113), .B(n110), .S(n608), .Z(n114) );
  MUX2_X1 U717 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n618), .Z(n115) );
  MUX2_X1 U718 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n618), .Z(n116) );
  MUX2_X1 U719 ( .A(n116), .B(n115), .S(n611), .Z(n117) );
  MUX2_X1 U720 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n618), .Z(n118) );
  MUX2_X1 U721 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n618), .Z(n119) );
  MUX2_X1 U722 ( .A(n119), .B(n118), .S(n610), .Z(n120) );
  MUX2_X1 U723 ( .A(n120), .B(n117), .S(n608), .Z(n121) );
  MUX2_X1 U724 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U725 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U726 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n618), .Z(n123) );
  MUX2_X1 U727 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n618), .Z(n124) );
  MUX2_X1 U728 ( .A(n124), .B(n123), .S(n612), .Z(n125) );
  MUX2_X1 U729 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n618), .Z(n126) );
  MUX2_X1 U730 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n618), .Z(n127) );
  MUX2_X1 U731 ( .A(n127), .B(n126), .S(n612), .Z(n128) );
  MUX2_X1 U732 ( .A(n128), .B(n125), .S(n608), .Z(n129) );
  MUX2_X1 U733 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n619), .Z(n130) );
  MUX2_X1 U734 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n619), .Z(n131) );
  MUX2_X1 U735 ( .A(n131), .B(n130), .S(N11), .Z(n132) );
  MUX2_X1 U736 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n619), .Z(n133) );
  MUX2_X1 U737 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n619), .Z(n134) );
  MUX2_X1 U738 ( .A(n134), .B(n133), .S(n610), .Z(n135) );
  MUX2_X1 U739 ( .A(n135), .B(n132), .S(n608), .Z(n136) );
  MUX2_X1 U740 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U741 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n619), .Z(n138) );
  MUX2_X1 U742 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n619), .Z(n139) );
  MUX2_X1 U743 ( .A(n139), .B(n138), .S(n610), .Z(n140) );
  MUX2_X1 U744 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n619), .Z(n141) );
  MUX2_X1 U745 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n619), .Z(n142) );
  MUX2_X1 U746 ( .A(n142), .B(n141), .S(n611), .Z(n143) );
  MUX2_X1 U747 ( .A(n143), .B(n140), .S(n608), .Z(n144) );
  MUX2_X1 U748 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n619), .Z(n145) );
  MUX2_X1 U749 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n619), .Z(n146) );
  MUX2_X1 U750 ( .A(n146), .B(n145), .S(n610), .Z(n147) );
  MUX2_X1 U751 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n619), .Z(n148) );
  MUX2_X1 U752 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n619), .Z(n149) );
  MUX2_X1 U753 ( .A(n149), .B(n148), .S(n612), .Z(n150) );
  MUX2_X1 U754 ( .A(n150), .B(n147), .S(n608), .Z(n151) );
  MUX2_X1 U755 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U756 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U757 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n620), .Z(n153) );
  MUX2_X1 U758 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n620), .Z(n154) );
  MUX2_X1 U759 ( .A(n154), .B(n153), .S(n611), .Z(n155) );
  MUX2_X1 U760 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n620), .Z(n156) );
  MUX2_X1 U761 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n620), .Z(n157) );
  MUX2_X1 U762 ( .A(n157), .B(n156), .S(n610), .Z(n158) );
  MUX2_X1 U763 ( .A(n158), .B(n155), .S(n609), .Z(n159) );
  MUX2_X1 U764 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n620), .Z(n160) );
  MUX2_X1 U765 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n620), .Z(n161) );
  MUX2_X1 U766 ( .A(n161), .B(n160), .S(n611), .Z(n162) );
  MUX2_X1 U767 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n620), .Z(n163) );
  MUX2_X1 U768 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n620), .Z(n164) );
  MUX2_X1 U769 ( .A(n164), .B(n163), .S(n610), .Z(n165) );
  MUX2_X1 U770 ( .A(n165), .B(n162), .S(n609), .Z(n166) );
  MUX2_X1 U771 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U772 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n620), .Z(n168) );
  MUX2_X1 U773 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n620), .Z(n169) );
  MUX2_X1 U774 ( .A(n169), .B(n168), .S(n612), .Z(n170) );
  MUX2_X1 U775 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n620), .Z(n171) );
  MUX2_X1 U776 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n620), .Z(n172) );
  MUX2_X1 U777 ( .A(n172), .B(n171), .S(N11), .Z(n173) );
  MUX2_X1 U778 ( .A(n173), .B(n170), .S(n609), .Z(n174) );
  MUX2_X1 U779 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n620), .Z(n175) );
  MUX2_X1 U780 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n622), .Z(n176) );
  MUX2_X1 U781 ( .A(n176), .B(n175), .S(N11), .Z(n177) );
  MUX2_X1 U782 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n622), .Z(n178) );
  MUX2_X1 U783 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n622), .Z(n179) );
  MUX2_X1 U784 ( .A(n179), .B(n178), .S(n612), .Z(n180) );
  MUX2_X1 U785 ( .A(n180), .B(n177), .S(n609), .Z(n181) );
  MUX2_X1 U786 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U787 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U788 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n622), .Z(n183) );
  MUX2_X1 U789 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n622), .Z(n184) );
  MUX2_X1 U790 ( .A(n184), .B(n183), .S(n611), .Z(n185) );
  MUX2_X1 U791 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n622), .Z(n186) );
  MUX2_X1 U792 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n615), .Z(n187) );
  MUX2_X1 U793 ( .A(n187), .B(n186), .S(N11), .Z(n188) );
  MUX2_X1 U794 ( .A(n188), .B(n185), .S(n609), .Z(n189) );
  MUX2_X1 U795 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n622), .Z(n190) );
  MUX2_X1 U796 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n614), .Z(n191) );
  MUX2_X1 U797 ( .A(n191), .B(n190), .S(N11), .Z(n192) );
  MUX2_X1 U798 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n616), .Z(n193) );
  MUX2_X1 U799 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n617), .Z(n194) );
  MUX2_X1 U800 ( .A(n194), .B(n193), .S(n612), .Z(n195) );
  MUX2_X1 U801 ( .A(n195), .B(n192), .S(n609), .Z(n196) );
  MUX2_X1 U802 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U803 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n621), .Z(n198) );
  MUX2_X1 U804 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n618), .Z(n199) );
  MUX2_X1 U805 ( .A(n199), .B(n198), .S(n610), .Z(n200) );
  MUX2_X1 U806 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n621), .Z(n201) );
  MUX2_X1 U807 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n621), .Z(n202) );
  MUX2_X1 U808 ( .A(n202), .B(n201), .S(n611), .Z(n203) );
  MUX2_X1 U809 ( .A(n203), .B(n200), .S(n609), .Z(n204) );
  MUX2_X1 U810 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n621), .Z(n205) );
  MUX2_X1 U811 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n622), .Z(n206) );
  MUX2_X1 U812 ( .A(n206), .B(n205), .S(n610), .Z(n207) );
  MUX2_X1 U813 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n622), .Z(n208) );
  MUX2_X1 U814 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n622), .Z(n209) );
  MUX2_X1 U815 ( .A(n209), .B(n208), .S(n612), .Z(n210) );
  MUX2_X1 U816 ( .A(n210), .B(n207), .S(n609), .Z(n211) );
  MUX2_X1 U817 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U818 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U819 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n613), .Z(n213) );
  MUX2_X1 U820 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n621), .Z(n214) );
  MUX2_X1 U821 ( .A(n214), .B(n213), .S(n610), .Z(n215) );
  MUX2_X1 U822 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n621), .Z(n216) );
  MUX2_X1 U823 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n619), .Z(n217) );
  MUX2_X1 U824 ( .A(n217), .B(n216), .S(n610), .Z(n218) );
  MUX2_X1 U825 ( .A(n218), .B(n215), .S(n609), .Z(n219) );
  MUX2_X1 U826 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n613), .Z(n220) );
  MUX2_X1 U827 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n622), .Z(n221) );
  MUX2_X1 U828 ( .A(n221), .B(n220), .S(n610), .Z(n222) );
  MUX2_X1 U829 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(N10), .Z(n223) );
  MUX2_X1 U830 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n224) );
  MUX2_X1 U831 ( .A(n224), .B(n223), .S(n611), .Z(n225) );
  MUX2_X1 U832 ( .A(n225), .B(n222), .S(n609), .Z(n226) );
  MUX2_X1 U833 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U834 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n613), .Z(n228) );
  MUX2_X1 U835 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n621), .Z(n229) );
  MUX2_X1 U836 ( .A(n229), .B(n228), .S(n610), .Z(n595) );
  MUX2_X1 U837 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(N10), .Z(n596) );
  MUX2_X1 U838 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n597) );
  MUX2_X1 U839 ( .A(n597), .B(n596), .S(n612), .Z(n598) );
  MUX2_X1 U840 ( .A(n598), .B(n595), .S(n609), .Z(n599) );
  MUX2_X1 U841 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n613), .Z(n600) );
  MUX2_X1 U842 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n622), .Z(n601) );
  MUX2_X1 U843 ( .A(n601), .B(n600), .S(n610), .Z(n602) );
  MUX2_X1 U844 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n621), .Z(n603) );
  MUX2_X1 U845 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n604) );
  MUX2_X1 U846 ( .A(n604), .B(n603), .S(n610), .Z(n605) );
  MUX2_X1 U847 ( .A(n605), .B(n602), .S(n609), .Z(n606) );
  MUX2_X1 U848 ( .A(n606), .B(n599), .S(N13), .Z(n607) );
  MUX2_X1 U849 ( .A(n607), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U850 ( .A(N11), .Z(n610) );
  INV_X1 U851 ( .A(N10), .ZN(n623) );
  INV_X1 U852 ( .A(N11), .ZN(n624) );
  INV_X1 U853 ( .A(data_in[0]), .ZN(n625) );
  INV_X1 U854 ( .A(data_in[1]), .ZN(n626) );
  INV_X1 U855 ( .A(data_in[2]), .ZN(n627) );
  INV_X1 U856 ( .A(data_in[3]), .ZN(n628) );
  INV_X1 U857 ( .A(data_in[4]), .ZN(n629) );
  INV_X1 U858 ( .A(data_in[5]), .ZN(n630) );
  INV_X1 U859 ( .A(data_in[6]), .ZN(n631) );
  INV_X1 U860 ( .A(data_in[7]), .ZN(n632) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_14 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n627), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n628), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n629), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n630), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n631), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n632), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n633), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n634), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n635), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n636), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n637), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n638), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n639), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n640), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n641), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n642), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n643), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n644), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n645), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n646), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n647), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n648), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n649), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n650), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n651), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n652), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n653), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n654), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n655), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n656), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n657), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n658), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n659), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n660), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n661), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n662), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n663), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n664), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n665), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n666), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n667), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n668), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n669), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n670), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n671), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n672), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n673), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n674), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n675), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n676), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n677), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n678), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n679), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n680), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n681), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n682), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n683), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n684), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n685), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n686), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n687), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n688), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n689), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n690), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n691), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n692), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n693), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n694), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n695), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n696), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n697), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n698), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n699), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n700), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n701), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n702), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n703), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n704), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n705), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n706), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n707), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n708), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n709), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n710), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n711), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n712), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n713), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n714), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n715), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n716), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n717), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n718), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n719), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n720), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n721), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n722), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n723), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n724), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n725), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n726), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n727), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n728), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n729), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n730), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n731), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n732), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n733), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n734), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n735), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n736), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n737), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n738), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n739), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n740), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n741), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n742), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n743), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n744), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n745), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n746), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n747), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n748), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n749), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n750), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n751), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n752), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n753), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n754), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n755), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n756), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n757), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n758), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n759), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n760), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n761), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n762), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n763), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n764), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n765), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n766), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n767), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n768), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n769), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n770), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n771), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n772), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n773), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n774), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n775), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n776), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n777), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n778), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n779), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n780), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n781), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n782), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n783), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n784), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n785), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n786), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n787), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n788), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n789), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n790), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n791), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n792), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n793), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n794), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n795), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n796), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n797), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n798), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n799), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n800), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n801), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n802), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n803), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n804), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n805), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n806), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n807), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n808), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n809), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n810), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n811), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n812), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n813), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n814), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n815), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n816), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n817), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n818), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n846), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n847), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n848), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n849), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n850), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n851), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n852), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n853), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n854), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n855), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n856), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n857), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n858), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n859), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n860), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n861), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n862), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n863), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n864), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n865), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n866), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n867), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n868), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n869), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n870), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n871), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n872), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n873), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n874), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n875), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n876), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n877), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n878), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n879), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n880), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n881), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n882), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n883), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n884), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n885), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n886), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n887), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n888), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n889), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n890), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n891), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n892), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n893), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n894), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n895), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n896), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n897), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n898), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n899), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n900), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n901), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n902), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n903), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n904), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n905), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n906), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n907), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n908), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n909), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X2 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n616), .Z(n613) );
  BUF_X1 U4 ( .A(n616), .Z(n614) );
  BUF_X1 U5 ( .A(n616), .Z(n615) );
  BUF_X1 U6 ( .A(N10), .Z(n611) );
  BUF_X1 U7 ( .A(n616), .Z(n612) );
  BUF_X1 U8 ( .A(N11), .Z(n609) );
  BUF_X1 U9 ( .A(N11), .Z(n610) );
  BUF_X1 U10 ( .A(N10), .Z(n616) );
  NOR3_X1 U11 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1201) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(n617), .ZN(n1190) );
  NOR3_X1 U13 ( .A1(N10), .A2(N12), .A3(n618), .ZN(n1180) );
  NOR3_X1 U14 ( .A1(n617), .A2(N12), .A3(n618), .ZN(n1170) );
  INV_X1 U15 ( .A(n1127), .ZN(n842) );
  INV_X1 U16 ( .A(n1117), .ZN(n841) );
  INV_X1 U17 ( .A(n1108), .ZN(n840) );
  INV_X1 U18 ( .A(n1099), .ZN(n839) );
  INV_X1 U19 ( .A(n1054), .ZN(n834) );
  INV_X1 U20 ( .A(n1044), .ZN(n833) );
  INV_X1 U21 ( .A(n1035), .ZN(n832) );
  INV_X1 U22 ( .A(n1026), .ZN(n831) );
  INV_X1 U23 ( .A(n981), .ZN(n826) );
  INV_X1 U24 ( .A(n971), .ZN(n825) );
  INV_X1 U25 ( .A(n962), .ZN(n824) );
  INV_X1 U26 ( .A(n953), .ZN(n823) );
  INV_X1 U27 ( .A(n944), .ZN(n822) );
  INV_X1 U28 ( .A(n935), .ZN(n821) );
  INV_X1 U29 ( .A(n926), .ZN(n820) );
  INV_X1 U30 ( .A(n917), .ZN(n819) );
  INV_X1 U31 ( .A(n1090), .ZN(n838) );
  INV_X1 U32 ( .A(n1081), .ZN(n837) );
  INV_X1 U33 ( .A(n1072), .ZN(n836) );
  INV_X1 U34 ( .A(n1063), .ZN(n835) );
  INV_X1 U35 ( .A(n1017), .ZN(n830) );
  INV_X1 U36 ( .A(n1008), .ZN(n829) );
  INV_X1 U37 ( .A(n999), .ZN(n828) );
  INV_X1 U38 ( .A(n990), .ZN(n827) );
  BUF_X1 U39 ( .A(N12), .Z(n606) );
  BUF_X1 U40 ( .A(N12), .Z(n607) );
  INV_X1 U41 ( .A(N13), .ZN(n844) );
  AND3_X1 U42 ( .A1(n617), .A2(n618), .A3(N12), .ZN(n1160) );
  AND3_X1 U43 ( .A1(N10), .A2(n618), .A3(N12), .ZN(n1150) );
  AND3_X1 U44 ( .A1(N11), .A2(n617), .A3(N12), .ZN(n1140) );
  AND3_X1 U45 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1130) );
  INV_X1 U46 ( .A(N14), .ZN(n845) );
  NAND2_X1 U47 ( .A1(n1190), .A2(n1200), .ZN(n1199) );
  NAND2_X1 U48 ( .A1(n1180), .A2(n1200), .ZN(n1189) );
  NAND2_X1 U49 ( .A1(n1170), .A2(n1200), .ZN(n1179) );
  NAND2_X1 U50 ( .A1(n1160), .A2(n1200), .ZN(n1169) );
  NAND2_X1 U51 ( .A1(n1150), .A2(n1200), .ZN(n1159) );
  NAND2_X1 U52 ( .A1(n1140), .A2(n1200), .ZN(n1149) );
  NAND2_X1 U53 ( .A1(n1130), .A2(n1200), .ZN(n1139) );
  NAND2_X1 U54 ( .A1(n1201), .A2(n1200), .ZN(n1210) );
  NAND2_X1 U55 ( .A1(n1119), .A2(n1201), .ZN(n1127) );
  NAND2_X1 U56 ( .A1(n1119), .A2(n1190), .ZN(n1117) );
  NAND2_X1 U57 ( .A1(n1119), .A2(n1180), .ZN(n1108) );
  NAND2_X1 U58 ( .A1(n1119), .A2(n1170), .ZN(n1099) );
  NAND2_X1 U59 ( .A1(n1046), .A2(n1201), .ZN(n1054) );
  NAND2_X1 U60 ( .A1(n1046), .A2(n1190), .ZN(n1044) );
  NAND2_X1 U61 ( .A1(n1046), .A2(n1180), .ZN(n1035) );
  NAND2_X1 U62 ( .A1(n1046), .A2(n1170), .ZN(n1026) );
  NAND2_X1 U63 ( .A1(n973), .A2(n1201), .ZN(n981) );
  NAND2_X1 U64 ( .A1(n973), .A2(n1190), .ZN(n971) );
  NAND2_X1 U65 ( .A1(n973), .A2(n1180), .ZN(n962) );
  NAND2_X1 U66 ( .A1(n973), .A2(n1170), .ZN(n953) );
  NAND2_X1 U67 ( .A1(n1119), .A2(n1160), .ZN(n1090) );
  NAND2_X1 U68 ( .A1(n1119), .A2(n1150), .ZN(n1081) );
  NAND2_X1 U69 ( .A1(n1119), .A2(n1140), .ZN(n1072) );
  NAND2_X1 U70 ( .A1(n1119), .A2(n1130), .ZN(n1063) );
  NAND2_X1 U71 ( .A1(n1046), .A2(n1160), .ZN(n1017) );
  NAND2_X1 U72 ( .A1(n1046), .A2(n1150), .ZN(n1008) );
  NAND2_X1 U73 ( .A1(n1046), .A2(n1140), .ZN(n999) );
  NAND2_X1 U74 ( .A1(n1046), .A2(n1130), .ZN(n990) );
  NAND2_X1 U75 ( .A1(n973), .A2(n1160), .ZN(n944) );
  NAND2_X1 U76 ( .A1(n973), .A2(n1150), .ZN(n935) );
  NAND2_X1 U77 ( .A1(n973), .A2(n1140), .ZN(n926) );
  NAND2_X1 U78 ( .A1(n973), .A2(n1130), .ZN(n917) );
  AND3_X1 U79 ( .A1(n844), .A2(n845), .A3(n1129), .ZN(n1200) );
  AND3_X1 U80 ( .A1(N13), .A2(n1129), .A3(N14), .ZN(n973) );
  AND3_X1 U81 ( .A1(n1129), .A2(n845), .A3(N13), .ZN(n1119) );
  AND3_X1 U82 ( .A1(n1129), .A2(n844), .A3(N14), .ZN(n1046) );
  NOR2_X1 U83 ( .A1(n843), .A2(addr[5]), .ZN(n1129) );
  INV_X1 U84 ( .A(wr_en), .ZN(n843) );
  OAI21_X1 U85 ( .B1(n619), .B2(n1169), .A(n1168), .ZN(n877) );
  NAND2_X1 U86 ( .A1(\mem[4][0] ), .A2(n1169), .ZN(n1168) );
  OAI21_X1 U87 ( .B1(n620), .B2(n1169), .A(n1167), .ZN(n876) );
  NAND2_X1 U88 ( .A1(\mem[4][1] ), .A2(n1169), .ZN(n1167) );
  OAI21_X1 U89 ( .B1(n621), .B2(n1169), .A(n1166), .ZN(n875) );
  NAND2_X1 U90 ( .A1(\mem[4][2] ), .A2(n1169), .ZN(n1166) );
  OAI21_X1 U91 ( .B1(n622), .B2(n1169), .A(n1165), .ZN(n874) );
  NAND2_X1 U92 ( .A1(\mem[4][3] ), .A2(n1169), .ZN(n1165) );
  OAI21_X1 U93 ( .B1(n623), .B2(n1169), .A(n1164), .ZN(n873) );
  NAND2_X1 U94 ( .A1(\mem[4][4] ), .A2(n1169), .ZN(n1164) );
  OAI21_X1 U95 ( .B1(n624), .B2(n1169), .A(n1163), .ZN(n872) );
  NAND2_X1 U96 ( .A1(\mem[4][5] ), .A2(n1169), .ZN(n1163) );
  OAI21_X1 U97 ( .B1(n625), .B2(n1169), .A(n1162), .ZN(n871) );
  NAND2_X1 U98 ( .A1(\mem[4][6] ), .A2(n1169), .ZN(n1162) );
  OAI21_X1 U99 ( .B1(n626), .B2(n1169), .A(n1161), .ZN(n870) );
  NAND2_X1 U100 ( .A1(\mem[4][7] ), .A2(n1169), .ZN(n1161) );
  OAI21_X1 U101 ( .B1(n619), .B2(n1149), .A(n1148), .ZN(n861) );
  NAND2_X1 U102 ( .A1(\mem[6][0] ), .A2(n1149), .ZN(n1148) );
  OAI21_X1 U103 ( .B1(n620), .B2(n1149), .A(n1147), .ZN(n860) );
  NAND2_X1 U104 ( .A1(\mem[6][1] ), .A2(n1149), .ZN(n1147) );
  OAI21_X1 U105 ( .B1(n621), .B2(n1149), .A(n1146), .ZN(n859) );
  NAND2_X1 U106 ( .A1(\mem[6][2] ), .A2(n1149), .ZN(n1146) );
  OAI21_X1 U107 ( .B1(n622), .B2(n1149), .A(n1145), .ZN(n858) );
  NAND2_X1 U108 ( .A1(\mem[6][3] ), .A2(n1149), .ZN(n1145) );
  OAI21_X1 U109 ( .B1(n623), .B2(n1149), .A(n1144), .ZN(n857) );
  NAND2_X1 U110 ( .A1(\mem[6][4] ), .A2(n1149), .ZN(n1144) );
  OAI21_X1 U111 ( .B1(n624), .B2(n1149), .A(n1143), .ZN(n856) );
  NAND2_X1 U112 ( .A1(\mem[6][5] ), .A2(n1149), .ZN(n1143) );
  OAI21_X1 U113 ( .B1(n625), .B2(n1149), .A(n1142), .ZN(n855) );
  NAND2_X1 U114 ( .A1(\mem[6][6] ), .A2(n1149), .ZN(n1142) );
  OAI21_X1 U115 ( .B1(n626), .B2(n1149), .A(n1141), .ZN(n854) );
  NAND2_X1 U116 ( .A1(\mem[6][7] ), .A2(n1149), .ZN(n1141) );
  OAI21_X1 U117 ( .B1(n619), .B2(n1139), .A(n1138), .ZN(n853) );
  NAND2_X1 U118 ( .A1(\mem[7][0] ), .A2(n1139), .ZN(n1138) );
  OAI21_X1 U119 ( .B1(n620), .B2(n1139), .A(n1137), .ZN(n852) );
  NAND2_X1 U120 ( .A1(\mem[7][1] ), .A2(n1139), .ZN(n1137) );
  OAI21_X1 U121 ( .B1(n621), .B2(n1139), .A(n1136), .ZN(n851) );
  NAND2_X1 U122 ( .A1(\mem[7][2] ), .A2(n1139), .ZN(n1136) );
  OAI21_X1 U123 ( .B1(n622), .B2(n1139), .A(n1135), .ZN(n850) );
  NAND2_X1 U124 ( .A1(\mem[7][3] ), .A2(n1139), .ZN(n1135) );
  OAI21_X1 U125 ( .B1(n623), .B2(n1139), .A(n1134), .ZN(n849) );
  NAND2_X1 U126 ( .A1(\mem[7][4] ), .A2(n1139), .ZN(n1134) );
  OAI21_X1 U127 ( .B1(n624), .B2(n1139), .A(n1133), .ZN(n848) );
  NAND2_X1 U128 ( .A1(\mem[7][5] ), .A2(n1139), .ZN(n1133) );
  OAI21_X1 U129 ( .B1(n625), .B2(n1139), .A(n1132), .ZN(n847) );
  NAND2_X1 U130 ( .A1(\mem[7][6] ), .A2(n1139), .ZN(n1132) );
  OAI21_X1 U131 ( .B1(n626), .B2(n1139), .A(n1131), .ZN(n846) );
  NAND2_X1 U132 ( .A1(\mem[7][7] ), .A2(n1139), .ZN(n1131) );
  OAI21_X1 U133 ( .B1(n619), .B2(n1199), .A(n1198), .ZN(n901) );
  NAND2_X1 U134 ( .A1(\mem[1][0] ), .A2(n1199), .ZN(n1198) );
  OAI21_X1 U135 ( .B1(n620), .B2(n1199), .A(n1197), .ZN(n900) );
  NAND2_X1 U136 ( .A1(\mem[1][1] ), .A2(n1199), .ZN(n1197) );
  OAI21_X1 U137 ( .B1(n621), .B2(n1199), .A(n1196), .ZN(n899) );
  NAND2_X1 U138 ( .A1(\mem[1][2] ), .A2(n1199), .ZN(n1196) );
  OAI21_X1 U139 ( .B1(n622), .B2(n1199), .A(n1195), .ZN(n898) );
  NAND2_X1 U140 ( .A1(\mem[1][3] ), .A2(n1199), .ZN(n1195) );
  OAI21_X1 U141 ( .B1(n623), .B2(n1199), .A(n1194), .ZN(n897) );
  NAND2_X1 U142 ( .A1(\mem[1][4] ), .A2(n1199), .ZN(n1194) );
  OAI21_X1 U143 ( .B1(n624), .B2(n1199), .A(n1193), .ZN(n896) );
  NAND2_X1 U144 ( .A1(\mem[1][5] ), .A2(n1199), .ZN(n1193) );
  OAI21_X1 U145 ( .B1(n625), .B2(n1199), .A(n1192), .ZN(n895) );
  NAND2_X1 U146 ( .A1(\mem[1][6] ), .A2(n1199), .ZN(n1192) );
  OAI21_X1 U147 ( .B1(n626), .B2(n1199), .A(n1191), .ZN(n894) );
  NAND2_X1 U148 ( .A1(\mem[1][7] ), .A2(n1199), .ZN(n1191) );
  OAI21_X1 U149 ( .B1(n619), .B2(n1189), .A(n1188), .ZN(n893) );
  NAND2_X1 U150 ( .A1(\mem[2][0] ), .A2(n1189), .ZN(n1188) );
  OAI21_X1 U151 ( .B1(n620), .B2(n1189), .A(n1187), .ZN(n892) );
  NAND2_X1 U152 ( .A1(\mem[2][1] ), .A2(n1189), .ZN(n1187) );
  OAI21_X1 U153 ( .B1(n621), .B2(n1189), .A(n1186), .ZN(n891) );
  NAND2_X1 U154 ( .A1(\mem[2][2] ), .A2(n1189), .ZN(n1186) );
  OAI21_X1 U155 ( .B1(n622), .B2(n1189), .A(n1185), .ZN(n890) );
  NAND2_X1 U156 ( .A1(\mem[2][3] ), .A2(n1189), .ZN(n1185) );
  OAI21_X1 U157 ( .B1(n623), .B2(n1189), .A(n1184), .ZN(n889) );
  NAND2_X1 U158 ( .A1(\mem[2][4] ), .A2(n1189), .ZN(n1184) );
  OAI21_X1 U159 ( .B1(n624), .B2(n1189), .A(n1183), .ZN(n888) );
  NAND2_X1 U160 ( .A1(\mem[2][5] ), .A2(n1189), .ZN(n1183) );
  OAI21_X1 U161 ( .B1(n625), .B2(n1189), .A(n1182), .ZN(n887) );
  NAND2_X1 U162 ( .A1(\mem[2][6] ), .A2(n1189), .ZN(n1182) );
  OAI21_X1 U163 ( .B1(n626), .B2(n1189), .A(n1181), .ZN(n886) );
  NAND2_X1 U164 ( .A1(\mem[2][7] ), .A2(n1189), .ZN(n1181) );
  OAI21_X1 U165 ( .B1(n619), .B2(n1179), .A(n1178), .ZN(n885) );
  NAND2_X1 U166 ( .A1(\mem[3][0] ), .A2(n1179), .ZN(n1178) );
  OAI21_X1 U167 ( .B1(n620), .B2(n1179), .A(n1177), .ZN(n884) );
  NAND2_X1 U168 ( .A1(\mem[3][1] ), .A2(n1179), .ZN(n1177) );
  OAI21_X1 U169 ( .B1(n621), .B2(n1179), .A(n1176), .ZN(n883) );
  NAND2_X1 U170 ( .A1(\mem[3][2] ), .A2(n1179), .ZN(n1176) );
  OAI21_X1 U171 ( .B1(n622), .B2(n1179), .A(n1175), .ZN(n882) );
  NAND2_X1 U172 ( .A1(\mem[3][3] ), .A2(n1179), .ZN(n1175) );
  OAI21_X1 U173 ( .B1(n623), .B2(n1179), .A(n1174), .ZN(n881) );
  NAND2_X1 U174 ( .A1(\mem[3][4] ), .A2(n1179), .ZN(n1174) );
  OAI21_X1 U175 ( .B1(n624), .B2(n1179), .A(n1173), .ZN(n880) );
  NAND2_X1 U176 ( .A1(\mem[3][5] ), .A2(n1179), .ZN(n1173) );
  OAI21_X1 U177 ( .B1(n625), .B2(n1179), .A(n1172), .ZN(n879) );
  NAND2_X1 U178 ( .A1(\mem[3][6] ), .A2(n1179), .ZN(n1172) );
  OAI21_X1 U179 ( .B1(n626), .B2(n1179), .A(n1171), .ZN(n878) );
  NAND2_X1 U180 ( .A1(\mem[3][7] ), .A2(n1179), .ZN(n1171) );
  OAI21_X1 U181 ( .B1(n619), .B2(n1159), .A(n1158), .ZN(n869) );
  NAND2_X1 U182 ( .A1(\mem[5][0] ), .A2(n1159), .ZN(n1158) );
  OAI21_X1 U183 ( .B1(n620), .B2(n1159), .A(n1157), .ZN(n868) );
  NAND2_X1 U184 ( .A1(\mem[5][1] ), .A2(n1159), .ZN(n1157) );
  OAI21_X1 U185 ( .B1(n621), .B2(n1159), .A(n1156), .ZN(n867) );
  NAND2_X1 U186 ( .A1(\mem[5][2] ), .A2(n1159), .ZN(n1156) );
  OAI21_X1 U187 ( .B1(n622), .B2(n1159), .A(n1155), .ZN(n866) );
  NAND2_X1 U188 ( .A1(\mem[5][3] ), .A2(n1159), .ZN(n1155) );
  OAI21_X1 U189 ( .B1(n623), .B2(n1159), .A(n1154), .ZN(n865) );
  NAND2_X1 U190 ( .A1(\mem[5][4] ), .A2(n1159), .ZN(n1154) );
  OAI21_X1 U191 ( .B1(n624), .B2(n1159), .A(n1153), .ZN(n864) );
  NAND2_X1 U192 ( .A1(\mem[5][5] ), .A2(n1159), .ZN(n1153) );
  OAI21_X1 U193 ( .B1(n625), .B2(n1159), .A(n1152), .ZN(n863) );
  NAND2_X1 U194 ( .A1(\mem[5][6] ), .A2(n1159), .ZN(n1152) );
  OAI21_X1 U195 ( .B1(n626), .B2(n1159), .A(n1151), .ZN(n862) );
  NAND2_X1 U196 ( .A1(\mem[5][7] ), .A2(n1159), .ZN(n1151) );
  OAI21_X1 U197 ( .B1(n1210), .B2(n619), .A(n1209), .ZN(n909) );
  NAND2_X1 U198 ( .A1(\mem[0][0] ), .A2(n1210), .ZN(n1209) );
  OAI21_X1 U199 ( .B1(n1210), .B2(n620), .A(n1208), .ZN(n908) );
  NAND2_X1 U200 ( .A1(\mem[0][1] ), .A2(n1210), .ZN(n1208) );
  OAI21_X1 U201 ( .B1(n1210), .B2(n621), .A(n1207), .ZN(n907) );
  NAND2_X1 U202 ( .A1(\mem[0][2] ), .A2(n1210), .ZN(n1207) );
  OAI21_X1 U203 ( .B1(n1210), .B2(n622), .A(n1206), .ZN(n906) );
  NAND2_X1 U204 ( .A1(\mem[0][3] ), .A2(n1210), .ZN(n1206) );
  OAI21_X1 U205 ( .B1(n1210), .B2(n623), .A(n1205), .ZN(n905) );
  NAND2_X1 U206 ( .A1(\mem[0][4] ), .A2(n1210), .ZN(n1205) );
  OAI21_X1 U207 ( .B1(n1210), .B2(n624), .A(n1204), .ZN(n904) );
  NAND2_X1 U208 ( .A1(\mem[0][5] ), .A2(n1210), .ZN(n1204) );
  OAI21_X1 U209 ( .B1(n1210), .B2(n625), .A(n1203), .ZN(n903) );
  NAND2_X1 U210 ( .A1(\mem[0][6] ), .A2(n1210), .ZN(n1203) );
  OAI21_X1 U211 ( .B1(n1210), .B2(n626), .A(n1202), .ZN(n902) );
  NAND2_X1 U212 ( .A1(\mem[0][7] ), .A2(n1210), .ZN(n1202) );
  INV_X1 U213 ( .A(n1128), .ZN(n818) );
  AOI22_X1 U214 ( .A1(data_in[0]), .A2(n842), .B1(n1127), .B2(\mem[8][0] ), 
        .ZN(n1128) );
  INV_X1 U215 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U216 ( .A1(data_in[1]), .A2(n842), .B1(n1127), .B2(\mem[8][1] ), 
        .ZN(n1126) );
  INV_X1 U217 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U218 ( .A1(data_in[2]), .A2(n842), .B1(n1127), .B2(\mem[8][2] ), 
        .ZN(n1125) );
  INV_X1 U219 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U220 ( .A1(data_in[3]), .A2(n842), .B1(n1127), .B2(\mem[8][3] ), 
        .ZN(n1124) );
  INV_X1 U221 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U222 ( .A1(data_in[4]), .A2(n842), .B1(n1127), .B2(\mem[8][4] ), 
        .ZN(n1123) );
  INV_X1 U223 ( .A(n1122), .ZN(n813) );
  AOI22_X1 U224 ( .A1(data_in[5]), .A2(n842), .B1(n1127), .B2(\mem[8][5] ), 
        .ZN(n1122) );
  INV_X1 U225 ( .A(n1121), .ZN(n812) );
  AOI22_X1 U226 ( .A1(data_in[6]), .A2(n842), .B1(n1127), .B2(\mem[8][6] ), 
        .ZN(n1121) );
  INV_X1 U227 ( .A(n1120), .ZN(n811) );
  AOI22_X1 U228 ( .A1(data_in[7]), .A2(n842), .B1(n1127), .B2(\mem[8][7] ), 
        .ZN(n1120) );
  INV_X1 U229 ( .A(n1118), .ZN(n810) );
  AOI22_X1 U230 ( .A1(data_in[0]), .A2(n841), .B1(n1117), .B2(\mem[9][0] ), 
        .ZN(n1118) );
  INV_X1 U231 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U232 ( .A1(data_in[1]), .A2(n841), .B1(n1117), .B2(\mem[9][1] ), 
        .ZN(n1116) );
  INV_X1 U233 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U234 ( .A1(data_in[2]), .A2(n841), .B1(n1117), .B2(\mem[9][2] ), 
        .ZN(n1115) );
  INV_X1 U235 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U236 ( .A1(data_in[3]), .A2(n841), .B1(n1117), .B2(\mem[9][3] ), 
        .ZN(n1114) );
  INV_X1 U237 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U238 ( .A1(data_in[4]), .A2(n841), .B1(n1117), .B2(\mem[9][4] ), 
        .ZN(n1113) );
  INV_X1 U239 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U240 ( .A1(data_in[5]), .A2(n841), .B1(n1117), .B2(\mem[9][5] ), 
        .ZN(n1112) );
  INV_X1 U241 ( .A(n1111), .ZN(n804) );
  AOI22_X1 U242 ( .A1(data_in[6]), .A2(n841), .B1(n1117), .B2(\mem[9][6] ), 
        .ZN(n1111) );
  INV_X1 U243 ( .A(n1110), .ZN(n803) );
  AOI22_X1 U244 ( .A1(data_in[7]), .A2(n841), .B1(n1117), .B2(\mem[9][7] ), 
        .ZN(n1110) );
  INV_X1 U245 ( .A(n1109), .ZN(n802) );
  AOI22_X1 U246 ( .A1(data_in[0]), .A2(n840), .B1(n1108), .B2(\mem[10][0] ), 
        .ZN(n1109) );
  INV_X1 U247 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U248 ( .A1(data_in[1]), .A2(n840), .B1(n1108), .B2(\mem[10][1] ), 
        .ZN(n1107) );
  INV_X1 U249 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U250 ( .A1(data_in[2]), .A2(n840), .B1(n1108), .B2(\mem[10][2] ), 
        .ZN(n1106) );
  INV_X1 U251 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U252 ( .A1(data_in[3]), .A2(n840), .B1(n1108), .B2(\mem[10][3] ), 
        .ZN(n1105) );
  INV_X1 U253 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U254 ( .A1(data_in[4]), .A2(n840), .B1(n1108), .B2(\mem[10][4] ), 
        .ZN(n1104) );
  INV_X1 U255 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U256 ( .A1(data_in[5]), .A2(n840), .B1(n1108), .B2(\mem[10][5] ), 
        .ZN(n1103) );
  INV_X1 U257 ( .A(n1102), .ZN(n796) );
  AOI22_X1 U258 ( .A1(data_in[6]), .A2(n840), .B1(n1108), .B2(\mem[10][6] ), 
        .ZN(n1102) );
  INV_X1 U259 ( .A(n1101), .ZN(n795) );
  AOI22_X1 U260 ( .A1(data_in[7]), .A2(n840), .B1(n1108), .B2(\mem[10][7] ), 
        .ZN(n1101) );
  INV_X1 U261 ( .A(n1100), .ZN(n794) );
  AOI22_X1 U262 ( .A1(data_in[0]), .A2(n839), .B1(n1099), .B2(\mem[11][0] ), 
        .ZN(n1100) );
  INV_X1 U263 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U264 ( .A1(data_in[1]), .A2(n839), .B1(n1099), .B2(\mem[11][1] ), 
        .ZN(n1098) );
  INV_X1 U265 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U266 ( .A1(data_in[2]), .A2(n839), .B1(n1099), .B2(\mem[11][2] ), 
        .ZN(n1097) );
  INV_X1 U267 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U268 ( .A1(data_in[3]), .A2(n839), .B1(n1099), .B2(\mem[11][3] ), 
        .ZN(n1096) );
  INV_X1 U269 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U270 ( .A1(data_in[4]), .A2(n839), .B1(n1099), .B2(\mem[11][4] ), 
        .ZN(n1095) );
  INV_X1 U271 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U272 ( .A1(data_in[5]), .A2(n839), .B1(n1099), .B2(\mem[11][5] ), 
        .ZN(n1094) );
  INV_X1 U273 ( .A(n1093), .ZN(n788) );
  AOI22_X1 U274 ( .A1(data_in[6]), .A2(n839), .B1(n1099), .B2(\mem[11][6] ), 
        .ZN(n1093) );
  INV_X1 U275 ( .A(n1092), .ZN(n787) );
  AOI22_X1 U276 ( .A1(data_in[7]), .A2(n839), .B1(n1099), .B2(\mem[11][7] ), 
        .ZN(n1092) );
  INV_X1 U277 ( .A(n1091), .ZN(n786) );
  AOI22_X1 U278 ( .A1(data_in[0]), .A2(n838), .B1(n1090), .B2(\mem[12][0] ), 
        .ZN(n1091) );
  INV_X1 U279 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U280 ( .A1(data_in[1]), .A2(n838), .B1(n1090), .B2(\mem[12][1] ), 
        .ZN(n1089) );
  INV_X1 U281 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U282 ( .A1(data_in[2]), .A2(n838), .B1(n1090), .B2(\mem[12][2] ), 
        .ZN(n1088) );
  INV_X1 U283 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U284 ( .A1(data_in[3]), .A2(n838), .B1(n1090), .B2(\mem[12][3] ), 
        .ZN(n1087) );
  INV_X1 U285 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U286 ( .A1(data_in[4]), .A2(n838), .B1(n1090), .B2(\mem[12][4] ), 
        .ZN(n1086) );
  INV_X1 U287 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U288 ( .A1(data_in[5]), .A2(n838), .B1(n1090), .B2(\mem[12][5] ), 
        .ZN(n1085) );
  INV_X1 U289 ( .A(n1084), .ZN(n780) );
  AOI22_X1 U290 ( .A1(data_in[6]), .A2(n838), .B1(n1090), .B2(\mem[12][6] ), 
        .ZN(n1084) );
  INV_X1 U291 ( .A(n1083), .ZN(n779) );
  AOI22_X1 U292 ( .A1(data_in[7]), .A2(n838), .B1(n1090), .B2(\mem[12][7] ), 
        .ZN(n1083) );
  INV_X1 U293 ( .A(n1082), .ZN(n778) );
  AOI22_X1 U294 ( .A1(data_in[0]), .A2(n837), .B1(n1081), .B2(\mem[13][0] ), 
        .ZN(n1082) );
  INV_X1 U295 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U296 ( .A1(data_in[1]), .A2(n837), .B1(n1081), .B2(\mem[13][1] ), 
        .ZN(n1080) );
  INV_X1 U297 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U298 ( .A1(data_in[2]), .A2(n837), .B1(n1081), .B2(\mem[13][2] ), 
        .ZN(n1079) );
  INV_X1 U299 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U300 ( .A1(data_in[3]), .A2(n837), .B1(n1081), .B2(\mem[13][3] ), 
        .ZN(n1078) );
  INV_X1 U301 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U302 ( .A1(data_in[4]), .A2(n837), .B1(n1081), .B2(\mem[13][4] ), 
        .ZN(n1077) );
  INV_X1 U303 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U304 ( .A1(data_in[5]), .A2(n837), .B1(n1081), .B2(\mem[13][5] ), 
        .ZN(n1076) );
  INV_X1 U305 ( .A(n1075), .ZN(n772) );
  AOI22_X1 U306 ( .A1(data_in[6]), .A2(n837), .B1(n1081), .B2(\mem[13][6] ), 
        .ZN(n1075) );
  INV_X1 U307 ( .A(n1074), .ZN(n771) );
  AOI22_X1 U308 ( .A1(data_in[7]), .A2(n837), .B1(n1081), .B2(\mem[13][7] ), 
        .ZN(n1074) );
  INV_X1 U309 ( .A(n1073), .ZN(n770) );
  AOI22_X1 U310 ( .A1(data_in[0]), .A2(n836), .B1(n1072), .B2(\mem[14][0] ), 
        .ZN(n1073) );
  INV_X1 U311 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U312 ( .A1(data_in[1]), .A2(n836), .B1(n1072), .B2(\mem[14][1] ), 
        .ZN(n1071) );
  INV_X1 U313 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U314 ( .A1(data_in[2]), .A2(n836), .B1(n1072), .B2(\mem[14][2] ), 
        .ZN(n1070) );
  INV_X1 U315 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U316 ( .A1(data_in[3]), .A2(n836), .B1(n1072), .B2(\mem[14][3] ), 
        .ZN(n1069) );
  INV_X1 U317 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U318 ( .A1(data_in[4]), .A2(n836), .B1(n1072), .B2(\mem[14][4] ), 
        .ZN(n1068) );
  INV_X1 U319 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U320 ( .A1(data_in[5]), .A2(n836), .B1(n1072), .B2(\mem[14][5] ), 
        .ZN(n1067) );
  INV_X1 U321 ( .A(n1066), .ZN(n764) );
  AOI22_X1 U322 ( .A1(data_in[6]), .A2(n836), .B1(n1072), .B2(\mem[14][6] ), 
        .ZN(n1066) );
  INV_X1 U323 ( .A(n1065), .ZN(n763) );
  AOI22_X1 U324 ( .A1(data_in[7]), .A2(n836), .B1(n1072), .B2(\mem[14][7] ), 
        .ZN(n1065) );
  INV_X1 U325 ( .A(n1064), .ZN(n762) );
  AOI22_X1 U326 ( .A1(data_in[0]), .A2(n835), .B1(n1063), .B2(\mem[15][0] ), 
        .ZN(n1064) );
  INV_X1 U327 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U328 ( .A1(data_in[1]), .A2(n835), .B1(n1063), .B2(\mem[15][1] ), 
        .ZN(n1062) );
  INV_X1 U329 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U330 ( .A1(data_in[2]), .A2(n835), .B1(n1063), .B2(\mem[15][2] ), 
        .ZN(n1061) );
  INV_X1 U331 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U332 ( .A1(data_in[3]), .A2(n835), .B1(n1063), .B2(\mem[15][3] ), 
        .ZN(n1060) );
  INV_X1 U333 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U334 ( .A1(data_in[4]), .A2(n835), .B1(n1063), .B2(\mem[15][4] ), 
        .ZN(n1059) );
  INV_X1 U335 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U336 ( .A1(data_in[5]), .A2(n835), .B1(n1063), .B2(\mem[15][5] ), 
        .ZN(n1058) );
  INV_X1 U337 ( .A(n1057), .ZN(n756) );
  AOI22_X1 U338 ( .A1(data_in[6]), .A2(n835), .B1(n1063), .B2(\mem[15][6] ), 
        .ZN(n1057) );
  INV_X1 U339 ( .A(n1056), .ZN(n755) );
  AOI22_X1 U340 ( .A1(data_in[7]), .A2(n835), .B1(n1063), .B2(\mem[15][7] ), 
        .ZN(n1056) );
  INV_X1 U341 ( .A(n1055), .ZN(n754) );
  AOI22_X1 U342 ( .A1(data_in[0]), .A2(n834), .B1(n1054), .B2(\mem[16][0] ), 
        .ZN(n1055) );
  INV_X1 U343 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U344 ( .A1(data_in[1]), .A2(n834), .B1(n1054), .B2(\mem[16][1] ), 
        .ZN(n1053) );
  INV_X1 U345 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U346 ( .A1(data_in[2]), .A2(n834), .B1(n1054), .B2(\mem[16][2] ), 
        .ZN(n1052) );
  INV_X1 U347 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U348 ( .A1(data_in[3]), .A2(n834), .B1(n1054), .B2(\mem[16][3] ), 
        .ZN(n1051) );
  INV_X1 U349 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U350 ( .A1(data_in[4]), .A2(n834), .B1(n1054), .B2(\mem[16][4] ), 
        .ZN(n1050) );
  INV_X1 U351 ( .A(n1049), .ZN(n749) );
  AOI22_X1 U352 ( .A1(data_in[5]), .A2(n834), .B1(n1054), .B2(\mem[16][5] ), 
        .ZN(n1049) );
  INV_X1 U353 ( .A(n1048), .ZN(n748) );
  AOI22_X1 U354 ( .A1(data_in[6]), .A2(n834), .B1(n1054), .B2(\mem[16][6] ), 
        .ZN(n1048) );
  INV_X1 U355 ( .A(n1047), .ZN(n747) );
  AOI22_X1 U356 ( .A1(data_in[7]), .A2(n834), .B1(n1054), .B2(\mem[16][7] ), 
        .ZN(n1047) );
  INV_X1 U357 ( .A(n1045), .ZN(n746) );
  AOI22_X1 U358 ( .A1(data_in[0]), .A2(n833), .B1(n1044), .B2(\mem[17][0] ), 
        .ZN(n1045) );
  INV_X1 U359 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U360 ( .A1(data_in[1]), .A2(n833), .B1(n1044), .B2(\mem[17][1] ), 
        .ZN(n1043) );
  INV_X1 U361 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U362 ( .A1(data_in[2]), .A2(n833), .B1(n1044), .B2(\mem[17][2] ), 
        .ZN(n1042) );
  INV_X1 U363 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U364 ( .A1(data_in[3]), .A2(n833), .B1(n1044), .B2(\mem[17][3] ), 
        .ZN(n1041) );
  INV_X1 U365 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U366 ( .A1(data_in[4]), .A2(n833), .B1(n1044), .B2(\mem[17][4] ), 
        .ZN(n1040) );
  INV_X1 U367 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U368 ( .A1(data_in[5]), .A2(n833), .B1(n1044), .B2(\mem[17][5] ), 
        .ZN(n1039) );
  INV_X1 U369 ( .A(n1038), .ZN(n740) );
  AOI22_X1 U370 ( .A1(data_in[6]), .A2(n833), .B1(n1044), .B2(\mem[17][6] ), 
        .ZN(n1038) );
  INV_X1 U371 ( .A(n1037), .ZN(n739) );
  AOI22_X1 U372 ( .A1(data_in[7]), .A2(n833), .B1(n1044), .B2(\mem[17][7] ), 
        .ZN(n1037) );
  INV_X1 U373 ( .A(n1036), .ZN(n738) );
  AOI22_X1 U374 ( .A1(data_in[0]), .A2(n832), .B1(n1035), .B2(\mem[18][0] ), 
        .ZN(n1036) );
  INV_X1 U375 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U376 ( .A1(data_in[1]), .A2(n832), .B1(n1035), .B2(\mem[18][1] ), 
        .ZN(n1034) );
  INV_X1 U377 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U378 ( .A1(data_in[2]), .A2(n832), .B1(n1035), .B2(\mem[18][2] ), 
        .ZN(n1033) );
  INV_X1 U379 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U380 ( .A1(data_in[3]), .A2(n832), .B1(n1035), .B2(\mem[18][3] ), 
        .ZN(n1032) );
  INV_X1 U381 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U382 ( .A1(data_in[4]), .A2(n832), .B1(n1035), .B2(\mem[18][4] ), 
        .ZN(n1031) );
  INV_X1 U383 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U384 ( .A1(data_in[5]), .A2(n832), .B1(n1035), .B2(\mem[18][5] ), 
        .ZN(n1030) );
  INV_X1 U385 ( .A(n1029), .ZN(n732) );
  AOI22_X1 U386 ( .A1(data_in[6]), .A2(n832), .B1(n1035), .B2(\mem[18][6] ), 
        .ZN(n1029) );
  INV_X1 U387 ( .A(n1028), .ZN(n731) );
  AOI22_X1 U388 ( .A1(data_in[7]), .A2(n832), .B1(n1035), .B2(\mem[18][7] ), 
        .ZN(n1028) );
  INV_X1 U389 ( .A(n1027), .ZN(n730) );
  AOI22_X1 U390 ( .A1(data_in[0]), .A2(n831), .B1(n1026), .B2(\mem[19][0] ), 
        .ZN(n1027) );
  INV_X1 U391 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U392 ( .A1(data_in[1]), .A2(n831), .B1(n1026), .B2(\mem[19][1] ), 
        .ZN(n1025) );
  INV_X1 U393 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U394 ( .A1(data_in[2]), .A2(n831), .B1(n1026), .B2(\mem[19][2] ), 
        .ZN(n1024) );
  INV_X1 U395 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U396 ( .A1(data_in[3]), .A2(n831), .B1(n1026), .B2(\mem[19][3] ), 
        .ZN(n1023) );
  INV_X1 U397 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U398 ( .A1(data_in[4]), .A2(n831), .B1(n1026), .B2(\mem[19][4] ), 
        .ZN(n1022) );
  INV_X1 U399 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U400 ( .A1(data_in[5]), .A2(n831), .B1(n1026), .B2(\mem[19][5] ), 
        .ZN(n1021) );
  INV_X1 U401 ( .A(n1020), .ZN(n724) );
  AOI22_X1 U402 ( .A1(data_in[6]), .A2(n831), .B1(n1026), .B2(\mem[19][6] ), 
        .ZN(n1020) );
  INV_X1 U403 ( .A(n1019), .ZN(n723) );
  AOI22_X1 U404 ( .A1(data_in[7]), .A2(n831), .B1(n1026), .B2(\mem[19][7] ), 
        .ZN(n1019) );
  INV_X1 U405 ( .A(n1018), .ZN(n722) );
  AOI22_X1 U406 ( .A1(data_in[0]), .A2(n830), .B1(n1017), .B2(\mem[20][0] ), 
        .ZN(n1018) );
  INV_X1 U407 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U408 ( .A1(data_in[1]), .A2(n830), .B1(n1017), .B2(\mem[20][1] ), 
        .ZN(n1016) );
  INV_X1 U409 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U410 ( .A1(data_in[2]), .A2(n830), .B1(n1017), .B2(\mem[20][2] ), 
        .ZN(n1015) );
  INV_X1 U411 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U412 ( .A1(data_in[3]), .A2(n830), .B1(n1017), .B2(\mem[20][3] ), 
        .ZN(n1014) );
  INV_X1 U413 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U414 ( .A1(data_in[4]), .A2(n830), .B1(n1017), .B2(\mem[20][4] ), 
        .ZN(n1013) );
  INV_X1 U415 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U416 ( .A1(data_in[5]), .A2(n830), .B1(n1017), .B2(\mem[20][5] ), 
        .ZN(n1012) );
  INV_X1 U417 ( .A(n1011), .ZN(n716) );
  AOI22_X1 U418 ( .A1(data_in[6]), .A2(n830), .B1(n1017), .B2(\mem[20][6] ), 
        .ZN(n1011) );
  INV_X1 U419 ( .A(n1010), .ZN(n715) );
  AOI22_X1 U420 ( .A1(data_in[7]), .A2(n830), .B1(n1017), .B2(\mem[20][7] ), 
        .ZN(n1010) );
  INV_X1 U421 ( .A(n1009), .ZN(n714) );
  AOI22_X1 U422 ( .A1(data_in[0]), .A2(n829), .B1(n1008), .B2(\mem[21][0] ), 
        .ZN(n1009) );
  INV_X1 U423 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U424 ( .A1(data_in[1]), .A2(n829), .B1(n1008), .B2(\mem[21][1] ), 
        .ZN(n1007) );
  INV_X1 U425 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U426 ( .A1(data_in[2]), .A2(n829), .B1(n1008), .B2(\mem[21][2] ), 
        .ZN(n1006) );
  INV_X1 U427 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U428 ( .A1(data_in[3]), .A2(n829), .B1(n1008), .B2(\mem[21][3] ), 
        .ZN(n1005) );
  INV_X1 U429 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U430 ( .A1(data_in[4]), .A2(n829), .B1(n1008), .B2(\mem[21][4] ), 
        .ZN(n1004) );
  INV_X1 U431 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U432 ( .A1(data_in[5]), .A2(n829), .B1(n1008), .B2(\mem[21][5] ), 
        .ZN(n1003) );
  INV_X1 U433 ( .A(n1002), .ZN(n708) );
  AOI22_X1 U434 ( .A1(data_in[6]), .A2(n829), .B1(n1008), .B2(\mem[21][6] ), 
        .ZN(n1002) );
  INV_X1 U435 ( .A(n1001), .ZN(n707) );
  AOI22_X1 U436 ( .A1(data_in[7]), .A2(n829), .B1(n1008), .B2(\mem[21][7] ), 
        .ZN(n1001) );
  INV_X1 U437 ( .A(n1000), .ZN(n706) );
  AOI22_X1 U438 ( .A1(data_in[0]), .A2(n828), .B1(n999), .B2(\mem[22][0] ), 
        .ZN(n1000) );
  INV_X1 U439 ( .A(n998), .ZN(n705) );
  AOI22_X1 U440 ( .A1(data_in[1]), .A2(n828), .B1(n999), .B2(\mem[22][1] ), 
        .ZN(n998) );
  INV_X1 U441 ( .A(n997), .ZN(n704) );
  AOI22_X1 U442 ( .A1(data_in[2]), .A2(n828), .B1(n999), .B2(\mem[22][2] ), 
        .ZN(n997) );
  INV_X1 U443 ( .A(n996), .ZN(n703) );
  AOI22_X1 U444 ( .A1(data_in[3]), .A2(n828), .B1(n999), .B2(\mem[22][3] ), 
        .ZN(n996) );
  INV_X1 U445 ( .A(n995), .ZN(n702) );
  AOI22_X1 U446 ( .A1(data_in[4]), .A2(n828), .B1(n999), .B2(\mem[22][4] ), 
        .ZN(n995) );
  INV_X1 U447 ( .A(n994), .ZN(n701) );
  AOI22_X1 U448 ( .A1(data_in[5]), .A2(n828), .B1(n999), .B2(\mem[22][5] ), 
        .ZN(n994) );
  INV_X1 U449 ( .A(n993), .ZN(n700) );
  AOI22_X1 U450 ( .A1(data_in[6]), .A2(n828), .B1(n999), .B2(\mem[22][6] ), 
        .ZN(n993) );
  INV_X1 U451 ( .A(n992), .ZN(n699) );
  AOI22_X1 U452 ( .A1(data_in[7]), .A2(n828), .B1(n999), .B2(\mem[22][7] ), 
        .ZN(n992) );
  INV_X1 U453 ( .A(n991), .ZN(n698) );
  AOI22_X1 U454 ( .A1(data_in[0]), .A2(n827), .B1(n990), .B2(\mem[23][0] ), 
        .ZN(n991) );
  INV_X1 U455 ( .A(n989), .ZN(n697) );
  AOI22_X1 U456 ( .A1(data_in[1]), .A2(n827), .B1(n990), .B2(\mem[23][1] ), 
        .ZN(n989) );
  INV_X1 U457 ( .A(n988), .ZN(n696) );
  AOI22_X1 U458 ( .A1(data_in[2]), .A2(n827), .B1(n990), .B2(\mem[23][2] ), 
        .ZN(n988) );
  INV_X1 U459 ( .A(n987), .ZN(n695) );
  AOI22_X1 U460 ( .A1(data_in[3]), .A2(n827), .B1(n990), .B2(\mem[23][3] ), 
        .ZN(n987) );
  INV_X1 U461 ( .A(n986), .ZN(n694) );
  AOI22_X1 U462 ( .A1(data_in[4]), .A2(n827), .B1(n990), .B2(\mem[23][4] ), 
        .ZN(n986) );
  INV_X1 U463 ( .A(n985), .ZN(n693) );
  AOI22_X1 U464 ( .A1(data_in[5]), .A2(n827), .B1(n990), .B2(\mem[23][5] ), 
        .ZN(n985) );
  INV_X1 U465 ( .A(n984), .ZN(n692) );
  AOI22_X1 U466 ( .A1(data_in[6]), .A2(n827), .B1(n990), .B2(\mem[23][6] ), 
        .ZN(n984) );
  INV_X1 U467 ( .A(n983), .ZN(n691) );
  AOI22_X1 U468 ( .A1(data_in[7]), .A2(n827), .B1(n990), .B2(\mem[23][7] ), 
        .ZN(n983) );
  INV_X1 U469 ( .A(n982), .ZN(n690) );
  AOI22_X1 U470 ( .A1(data_in[0]), .A2(n826), .B1(n981), .B2(\mem[24][0] ), 
        .ZN(n982) );
  INV_X1 U471 ( .A(n980), .ZN(n689) );
  AOI22_X1 U472 ( .A1(data_in[1]), .A2(n826), .B1(n981), .B2(\mem[24][1] ), 
        .ZN(n980) );
  INV_X1 U473 ( .A(n979), .ZN(n688) );
  AOI22_X1 U474 ( .A1(data_in[2]), .A2(n826), .B1(n981), .B2(\mem[24][2] ), 
        .ZN(n979) );
  INV_X1 U475 ( .A(n978), .ZN(n687) );
  AOI22_X1 U476 ( .A1(data_in[3]), .A2(n826), .B1(n981), .B2(\mem[24][3] ), 
        .ZN(n978) );
  INV_X1 U477 ( .A(n977), .ZN(n686) );
  AOI22_X1 U478 ( .A1(data_in[4]), .A2(n826), .B1(n981), .B2(\mem[24][4] ), 
        .ZN(n977) );
  INV_X1 U479 ( .A(n976), .ZN(n685) );
  AOI22_X1 U480 ( .A1(data_in[5]), .A2(n826), .B1(n981), .B2(\mem[24][5] ), 
        .ZN(n976) );
  INV_X1 U481 ( .A(n975), .ZN(n684) );
  AOI22_X1 U482 ( .A1(data_in[6]), .A2(n826), .B1(n981), .B2(\mem[24][6] ), 
        .ZN(n975) );
  INV_X1 U483 ( .A(n974), .ZN(n683) );
  AOI22_X1 U484 ( .A1(data_in[7]), .A2(n826), .B1(n981), .B2(\mem[24][7] ), 
        .ZN(n974) );
  INV_X1 U485 ( .A(n972), .ZN(n682) );
  AOI22_X1 U486 ( .A1(data_in[0]), .A2(n825), .B1(n971), .B2(\mem[25][0] ), 
        .ZN(n972) );
  INV_X1 U487 ( .A(n970), .ZN(n681) );
  AOI22_X1 U488 ( .A1(data_in[1]), .A2(n825), .B1(n971), .B2(\mem[25][1] ), 
        .ZN(n970) );
  INV_X1 U489 ( .A(n969), .ZN(n680) );
  AOI22_X1 U490 ( .A1(data_in[2]), .A2(n825), .B1(n971), .B2(\mem[25][2] ), 
        .ZN(n969) );
  INV_X1 U491 ( .A(n968), .ZN(n679) );
  AOI22_X1 U492 ( .A1(data_in[3]), .A2(n825), .B1(n971), .B2(\mem[25][3] ), 
        .ZN(n968) );
  INV_X1 U493 ( .A(n967), .ZN(n678) );
  AOI22_X1 U494 ( .A1(data_in[4]), .A2(n825), .B1(n971), .B2(\mem[25][4] ), 
        .ZN(n967) );
  INV_X1 U495 ( .A(n966), .ZN(n677) );
  AOI22_X1 U496 ( .A1(data_in[5]), .A2(n825), .B1(n971), .B2(\mem[25][5] ), 
        .ZN(n966) );
  INV_X1 U497 ( .A(n965), .ZN(n676) );
  AOI22_X1 U498 ( .A1(data_in[6]), .A2(n825), .B1(n971), .B2(\mem[25][6] ), 
        .ZN(n965) );
  INV_X1 U499 ( .A(n964), .ZN(n675) );
  AOI22_X1 U500 ( .A1(data_in[7]), .A2(n825), .B1(n971), .B2(\mem[25][7] ), 
        .ZN(n964) );
  INV_X1 U501 ( .A(n963), .ZN(n674) );
  AOI22_X1 U502 ( .A1(data_in[0]), .A2(n824), .B1(n962), .B2(\mem[26][0] ), 
        .ZN(n963) );
  INV_X1 U503 ( .A(n961), .ZN(n673) );
  AOI22_X1 U504 ( .A1(data_in[1]), .A2(n824), .B1(n962), .B2(\mem[26][1] ), 
        .ZN(n961) );
  INV_X1 U505 ( .A(n960), .ZN(n672) );
  AOI22_X1 U506 ( .A1(data_in[2]), .A2(n824), .B1(n962), .B2(\mem[26][2] ), 
        .ZN(n960) );
  INV_X1 U507 ( .A(n959), .ZN(n671) );
  AOI22_X1 U508 ( .A1(data_in[3]), .A2(n824), .B1(n962), .B2(\mem[26][3] ), 
        .ZN(n959) );
  INV_X1 U509 ( .A(n958), .ZN(n670) );
  AOI22_X1 U510 ( .A1(data_in[4]), .A2(n824), .B1(n962), .B2(\mem[26][4] ), 
        .ZN(n958) );
  INV_X1 U511 ( .A(n957), .ZN(n669) );
  AOI22_X1 U512 ( .A1(data_in[5]), .A2(n824), .B1(n962), .B2(\mem[26][5] ), 
        .ZN(n957) );
  INV_X1 U513 ( .A(n956), .ZN(n668) );
  AOI22_X1 U514 ( .A1(data_in[6]), .A2(n824), .B1(n962), .B2(\mem[26][6] ), 
        .ZN(n956) );
  INV_X1 U515 ( .A(n955), .ZN(n667) );
  AOI22_X1 U516 ( .A1(data_in[7]), .A2(n824), .B1(n962), .B2(\mem[26][7] ), 
        .ZN(n955) );
  INV_X1 U517 ( .A(n954), .ZN(n666) );
  AOI22_X1 U518 ( .A1(data_in[0]), .A2(n823), .B1(n953), .B2(\mem[27][0] ), 
        .ZN(n954) );
  INV_X1 U519 ( .A(n952), .ZN(n665) );
  AOI22_X1 U520 ( .A1(data_in[1]), .A2(n823), .B1(n953), .B2(\mem[27][1] ), 
        .ZN(n952) );
  INV_X1 U521 ( .A(n951), .ZN(n664) );
  AOI22_X1 U522 ( .A1(data_in[2]), .A2(n823), .B1(n953), .B2(\mem[27][2] ), 
        .ZN(n951) );
  INV_X1 U523 ( .A(n950), .ZN(n663) );
  AOI22_X1 U524 ( .A1(data_in[3]), .A2(n823), .B1(n953), .B2(\mem[27][3] ), 
        .ZN(n950) );
  INV_X1 U525 ( .A(n949), .ZN(n662) );
  AOI22_X1 U526 ( .A1(data_in[4]), .A2(n823), .B1(n953), .B2(\mem[27][4] ), 
        .ZN(n949) );
  INV_X1 U527 ( .A(n948), .ZN(n661) );
  AOI22_X1 U528 ( .A1(data_in[5]), .A2(n823), .B1(n953), .B2(\mem[27][5] ), 
        .ZN(n948) );
  INV_X1 U529 ( .A(n947), .ZN(n660) );
  AOI22_X1 U530 ( .A1(data_in[6]), .A2(n823), .B1(n953), .B2(\mem[27][6] ), 
        .ZN(n947) );
  INV_X1 U531 ( .A(n946), .ZN(n659) );
  AOI22_X1 U532 ( .A1(data_in[7]), .A2(n823), .B1(n953), .B2(\mem[27][7] ), 
        .ZN(n946) );
  INV_X1 U533 ( .A(n945), .ZN(n658) );
  AOI22_X1 U534 ( .A1(data_in[0]), .A2(n822), .B1(n944), .B2(\mem[28][0] ), 
        .ZN(n945) );
  INV_X1 U535 ( .A(n943), .ZN(n657) );
  AOI22_X1 U536 ( .A1(data_in[1]), .A2(n822), .B1(n944), .B2(\mem[28][1] ), 
        .ZN(n943) );
  INV_X1 U537 ( .A(n942), .ZN(n656) );
  AOI22_X1 U538 ( .A1(data_in[2]), .A2(n822), .B1(n944), .B2(\mem[28][2] ), 
        .ZN(n942) );
  INV_X1 U539 ( .A(n941), .ZN(n655) );
  AOI22_X1 U540 ( .A1(data_in[3]), .A2(n822), .B1(n944), .B2(\mem[28][3] ), 
        .ZN(n941) );
  INV_X1 U541 ( .A(n940), .ZN(n654) );
  AOI22_X1 U542 ( .A1(data_in[4]), .A2(n822), .B1(n944), .B2(\mem[28][4] ), 
        .ZN(n940) );
  INV_X1 U543 ( .A(n939), .ZN(n653) );
  AOI22_X1 U544 ( .A1(data_in[5]), .A2(n822), .B1(n944), .B2(\mem[28][5] ), 
        .ZN(n939) );
  INV_X1 U545 ( .A(n938), .ZN(n652) );
  AOI22_X1 U546 ( .A1(data_in[6]), .A2(n822), .B1(n944), .B2(\mem[28][6] ), 
        .ZN(n938) );
  INV_X1 U547 ( .A(n937), .ZN(n651) );
  AOI22_X1 U548 ( .A1(data_in[7]), .A2(n822), .B1(n944), .B2(\mem[28][7] ), 
        .ZN(n937) );
  INV_X1 U549 ( .A(n936), .ZN(n650) );
  AOI22_X1 U550 ( .A1(data_in[0]), .A2(n821), .B1(n935), .B2(\mem[29][0] ), 
        .ZN(n936) );
  INV_X1 U551 ( .A(n934), .ZN(n649) );
  AOI22_X1 U552 ( .A1(data_in[1]), .A2(n821), .B1(n935), .B2(\mem[29][1] ), 
        .ZN(n934) );
  INV_X1 U553 ( .A(n933), .ZN(n648) );
  AOI22_X1 U554 ( .A1(data_in[2]), .A2(n821), .B1(n935), .B2(\mem[29][2] ), 
        .ZN(n933) );
  INV_X1 U555 ( .A(n932), .ZN(n647) );
  AOI22_X1 U556 ( .A1(data_in[3]), .A2(n821), .B1(n935), .B2(\mem[29][3] ), 
        .ZN(n932) );
  INV_X1 U557 ( .A(n931), .ZN(n646) );
  AOI22_X1 U558 ( .A1(data_in[4]), .A2(n821), .B1(n935), .B2(\mem[29][4] ), 
        .ZN(n931) );
  INV_X1 U559 ( .A(n930), .ZN(n645) );
  AOI22_X1 U560 ( .A1(data_in[5]), .A2(n821), .B1(n935), .B2(\mem[29][5] ), 
        .ZN(n930) );
  INV_X1 U561 ( .A(n929), .ZN(n644) );
  AOI22_X1 U562 ( .A1(data_in[6]), .A2(n821), .B1(n935), .B2(\mem[29][6] ), 
        .ZN(n929) );
  INV_X1 U563 ( .A(n928), .ZN(n643) );
  AOI22_X1 U564 ( .A1(data_in[7]), .A2(n821), .B1(n935), .B2(\mem[29][7] ), 
        .ZN(n928) );
  INV_X1 U565 ( .A(n927), .ZN(n642) );
  AOI22_X1 U566 ( .A1(data_in[0]), .A2(n820), .B1(n926), .B2(\mem[30][0] ), 
        .ZN(n927) );
  INV_X1 U567 ( .A(n925), .ZN(n641) );
  AOI22_X1 U568 ( .A1(data_in[1]), .A2(n820), .B1(n926), .B2(\mem[30][1] ), 
        .ZN(n925) );
  INV_X1 U569 ( .A(n924), .ZN(n640) );
  AOI22_X1 U570 ( .A1(data_in[2]), .A2(n820), .B1(n926), .B2(\mem[30][2] ), 
        .ZN(n924) );
  INV_X1 U571 ( .A(n923), .ZN(n639) );
  AOI22_X1 U572 ( .A1(data_in[3]), .A2(n820), .B1(n926), .B2(\mem[30][3] ), 
        .ZN(n923) );
  INV_X1 U573 ( .A(n922), .ZN(n638) );
  AOI22_X1 U574 ( .A1(data_in[4]), .A2(n820), .B1(n926), .B2(\mem[30][4] ), 
        .ZN(n922) );
  INV_X1 U575 ( .A(n921), .ZN(n637) );
  AOI22_X1 U576 ( .A1(data_in[5]), .A2(n820), .B1(n926), .B2(\mem[30][5] ), 
        .ZN(n921) );
  INV_X1 U577 ( .A(n920), .ZN(n636) );
  AOI22_X1 U578 ( .A1(data_in[6]), .A2(n820), .B1(n926), .B2(\mem[30][6] ), 
        .ZN(n920) );
  INV_X1 U579 ( .A(n919), .ZN(n635) );
  AOI22_X1 U580 ( .A1(data_in[7]), .A2(n820), .B1(n926), .B2(\mem[30][7] ), 
        .ZN(n919) );
  INV_X1 U581 ( .A(n918), .ZN(n634) );
  AOI22_X1 U582 ( .A1(data_in[0]), .A2(n819), .B1(n917), .B2(\mem[31][0] ), 
        .ZN(n918) );
  INV_X1 U583 ( .A(n916), .ZN(n633) );
  AOI22_X1 U584 ( .A1(data_in[1]), .A2(n819), .B1(n917), .B2(\mem[31][1] ), 
        .ZN(n916) );
  INV_X1 U585 ( .A(n915), .ZN(n632) );
  AOI22_X1 U586 ( .A1(data_in[2]), .A2(n819), .B1(n917), .B2(\mem[31][2] ), 
        .ZN(n915) );
  INV_X1 U587 ( .A(n914), .ZN(n631) );
  AOI22_X1 U588 ( .A1(data_in[3]), .A2(n819), .B1(n917), .B2(\mem[31][3] ), 
        .ZN(n914) );
  INV_X1 U589 ( .A(n913), .ZN(n630) );
  AOI22_X1 U590 ( .A1(data_in[4]), .A2(n819), .B1(n917), .B2(\mem[31][4] ), 
        .ZN(n913) );
  INV_X1 U591 ( .A(n912), .ZN(n629) );
  AOI22_X1 U592 ( .A1(data_in[5]), .A2(n819), .B1(n917), .B2(\mem[31][5] ), 
        .ZN(n912) );
  INV_X1 U593 ( .A(n911), .ZN(n628) );
  AOI22_X1 U594 ( .A1(data_in[6]), .A2(n819), .B1(n917), .B2(\mem[31][6] ), 
        .ZN(n911) );
  INV_X1 U595 ( .A(n910), .ZN(n627) );
  AOI22_X1 U596 ( .A1(data_in[7]), .A2(n819), .B1(n917), .B2(\mem[31][7] ), 
        .ZN(n910) );
  MUX2_X1 U597 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n612), .Z(n1) );
  MUX2_X1 U598 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n613), .Z(n2) );
  MUX2_X1 U599 ( .A(n2), .B(n1), .S(n608), .Z(n3) );
  MUX2_X1 U600 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n613), .Z(n4) );
  MUX2_X1 U601 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n613), .Z(n5) );
  MUX2_X1 U602 ( .A(n5), .B(n4), .S(n608), .Z(n6) );
  MUX2_X1 U603 ( .A(n6), .B(n3), .S(n607), .Z(n7) );
  MUX2_X1 U604 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n612), .Z(n8) );
  MUX2_X1 U605 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n615), .Z(n9) );
  MUX2_X1 U606 ( .A(n9), .B(n8), .S(n608), .Z(n10) );
  MUX2_X1 U607 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n614), .Z(n11) );
  MUX2_X1 U608 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n612), .Z(n12) );
  MUX2_X1 U609 ( .A(n12), .B(n11), .S(n608), .Z(n13) );
  MUX2_X1 U610 ( .A(n13), .B(n10), .S(N12), .Z(n14) );
  MUX2_X1 U611 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U612 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n615), .Z(n16) );
  MUX2_X1 U613 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n616), .Z(n17) );
  MUX2_X1 U614 ( .A(n17), .B(n16), .S(n608), .Z(n18) );
  MUX2_X1 U615 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(N10), .Z(n19) );
  MUX2_X1 U616 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n20) );
  MUX2_X1 U617 ( .A(n20), .B(n19), .S(n610), .Z(n21) );
  MUX2_X1 U618 ( .A(n21), .B(n18), .S(N12), .Z(n22) );
  MUX2_X1 U619 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n615), .Z(n23) );
  MUX2_X1 U620 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n24) );
  MUX2_X1 U621 ( .A(n24), .B(n23), .S(n608), .Z(n25) );
  MUX2_X1 U622 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n616), .Z(n26) );
  MUX2_X1 U623 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n616), .Z(n27) );
  MUX2_X1 U624 ( .A(n27), .B(n26), .S(n609), .Z(n28) );
  MUX2_X1 U625 ( .A(n28), .B(n25), .S(n606), .Z(n29) );
  MUX2_X1 U626 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U627 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U628 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n611), .Z(n31) );
  MUX2_X1 U629 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n613), .Z(n32) );
  MUX2_X1 U630 ( .A(n32), .B(n31), .S(n608), .Z(n33) );
  MUX2_X1 U631 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n612), .Z(n34) );
  MUX2_X1 U632 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n616), .Z(n35) );
  MUX2_X1 U633 ( .A(n35), .B(n34), .S(n608), .Z(n36) );
  MUX2_X1 U634 ( .A(n36), .B(n33), .S(n606), .Z(n37) );
  MUX2_X1 U635 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n614), .Z(n38) );
  MUX2_X1 U636 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n614), .Z(n39) );
  MUX2_X1 U637 ( .A(n39), .B(n38), .S(n608), .Z(n40) );
  MUX2_X1 U638 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n616), .Z(n41) );
  MUX2_X1 U639 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(N10), .Z(n42) );
  MUX2_X1 U640 ( .A(n42), .B(n41), .S(n609), .Z(n43) );
  MUX2_X1 U641 ( .A(n43), .B(n40), .S(n607), .Z(n44) );
  MUX2_X1 U642 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U643 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n615), .Z(n46) );
  MUX2_X1 U644 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n614), .Z(n47) );
  MUX2_X1 U645 ( .A(n47), .B(n46), .S(n608), .Z(n48) );
  MUX2_X1 U646 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n615), .Z(n49) );
  MUX2_X1 U647 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n615), .Z(n50) );
  MUX2_X1 U648 ( .A(n50), .B(n49), .S(n610), .Z(n51) );
  MUX2_X1 U649 ( .A(n51), .B(n48), .S(N12), .Z(n52) );
  MUX2_X1 U650 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n612), .Z(n53) );
  MUX2_X1 U651 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n614), .Z(n54) );
  MUX2_X1 U652 ( .A(n54), .B(n53), .S(n608), .Z(n55) );
  MUX2_X1 U653 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n615), .Z(n56) );
  MUX2_X1 U654 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n614), .Z(n57) );
  MUX2_X1 U655 ( .A(n57), .B(n56), .S(n608), .Z(n58) );
  MUX2_X1 U656 ( .A(n58), .B(n55), .S(n607), .Z(n59) );
  MUX2_X1 U657 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U658 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U659 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n611), .Z(n61) );
  MUX2_X1 U660 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n611), .Z(n62) );
  MUX2_X1 U661 ( .A(n62), .B(n61), .S(n609), .Z(n63) );
  MUX2_X1 U662 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n611), .Z(n64) );
  MUX2_X1 U663 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n611), .Z(n65) );
  MUX2_X1 U664 ( .A(n65), .B(n64), .S(n609), .Z(n66) );
  MUX2_X1 U665 ( .A(n66), .B(n63), .S(n606), .Z(n67) );
  MUX2_X1 U666 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n611), .Z(n68) );
  MUX2_X1 U667 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n611), .Z(n69) );
  MUX2_X1 U668 ( .A(n69), .B(n68), .S(n609), .Z(n70) );
  MUX2_X1 U669 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n611), .Z(n71) );
  MUX2_X1 U670 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n611), .Z(n72) );
  MUX2_X1 U671 ( .A(n72), .B(n71), .S(n609), .Z(n73) );
  MUX2_X1 U672 ( .A(n73), .B(n70), .S(n606), .Z(n74) );
  MUX2_X1 U673 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U674 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n611), .Z(n76) );
  MUX2_X1 U675 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n611), .Z(n77) );
  MUX2_X1 U676 ( .A(n77), .B(n76), .S(n609), .Z(n78) );
  MUX2_X1 U677 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n611), .Z(n79) );
  MUX2_X1 U678 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n611), .Z(n80) );
  MUX2_X1 U679 ( .A(n80), .B(n79), .S(n609), .Z(n81) );
  MUX2_X1 U680 ( .A(n81), .B(n78), .S(n606), .Z(n82) );
  MUX2_X1 U681 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n612), .Z(n83) );
  MUX2_X1 U682 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n612), .Z(n84) );
  MUX2_X1 U683 ( .A(n84), .B(n83), .S(n609), .Z(n85) );
  MUX2_X1 U684 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n612), .Z(n86) );
  MUX2_X1 U685 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n612), .Z(n87) );
  MUX2_X1 U686 ( .A(n87), .B(n86), .S(n609), .Z(n88) );
  MUX2_X1 U687 ( .A(n88), .B(n85), .S(n606), .Z(n89) );
  MUX2_X1 U688 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U689 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U690 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n612), .Z(n91) );
  MUX2_X1 U691 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n612), .Z(n92) );
  MUX2_X1 U692 ( .A(n92), .B(n91), .S(n609), .Z(n93) );
  MUX2_X1 U693 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n612), .Z(n94) );
  MUX2_X1 U694 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n612), .Z(n95) );
  MUX2_X1 U695 ( .A(n95), .B(n94), .S(n609), .Z(n96) );
  MUX2_X1 U696 ( .A(n96), .B(n93), .S(n606), .Z(n97) );
  MUX2_X1 U697 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n612), .Z(n98) );
  MUX2_X1 U698 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n612), .Z(n99) );
  MUX2_X1 U699 ( .A(n99), .B(n98), .S(n609), .Z(n100) );
  MUX2_X1 U700 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n612), .Z(n101) );
  MUX2_X1 U701 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n612), .Z(n102) );
  MUX2_X1 U702 ( .A(n102), .B(n101), .S(n609), .Z(n103) );
  MUX2_X1 U703 ( .A(n103), .B(n100), .S(n606), .Z(n104) );
  MUX2_X1 U704 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U705 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n613), .Z(n106) );
  MUX2_X1 U706 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n616), .Z(n107) );
  MUX2_X1 U707 ( .A(n107), .B(n106), .S(n610), .Z(n108) );
  MUX2_X1 U708 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n616), .Z(n109) );
  MUX2_X1 U709 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n616), .Z(n110) );
  MUX2_X1 U710 ( .A(n110), .B(n109), .S(n610), .Z(n111) );
  MUX2_X1 U711 ( .A(n111), .B(n108), .S(n606), .Z(n112) );
  MUX2_X1 U712 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n616), .Z(n113) );
  MUX2_X1 U713 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n616), .Z(n114) );
  MUX2_X1 U714 ( .A(n114), .B(n113), .S(n610), .Z(n115) );
  MUX2_X1 U715 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n616), .Z(n116) );
  MUX2_X1 U716 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n616), .Z(n117) );
  MUX2_X1 U717 ( .A(n117), .B(n116), .S(n610), .Z(n118) );
  MUX2_X1 U718 ( .A(n118), .B(n115), .S(n606), .Z(n119) );
  MUX2_X1 U719 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U720 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U721 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n614), .Z(n121) );
  MUX2_X1 U722 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n613), .Z(n122) );
  MUX2_X1 U723 ( .A(n122), .B(n121), .S(n610), .Z(n123) );
  MUX2_X1 U724 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n612), .Z(n124) );
  MUX2_X1 U725 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n614), .Z(n125) );
  MUX2_X1 U726 ( .A(n125), .B(n124), .S(n610), .Z(n126) );
  MUX2_X1 U727 ( .A(n126), .B(n123), .S(n606), .Z(n127) );
  MUX2_X1 U728 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n612), .Z(n128) );
  MUX2_X1 U729 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n616), .Z(n129) );
  MUX2_X1 U730 ( .A(n129), .B(n128), .S(n610), .Z(n130) );
  MUX2_X1 U731 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(N10), .Z(n131) );
  MUX2_X1 U732 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n616), .Z(n132) );
  MUX2_X1 U733 ( .A(n132), .B(n131), .S(n610), .Z(n133) );
  MUX2_X1 U734 ( .A(n133), .B(n130), .S(n606), .Z(n134) );
  MUX2_X1 U735 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U736 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n615), .Z(n136) );
  MUX2_X1 U737 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n616), .Z(n137) );
  MUX2_X1 U738 ( .A(n137), .B(n136), .S(n610), .Z(n138) );
  MUX2_X1 U739 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n613), .Z(n139) );
  MUX2_X1 U740 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n616), .Z(n140) );
  MUX2_X1 U741 ( .A(n140), .B(n139), .S(n610), .Z(n141) );
  MUX2_X1 U742 ( .A(n141), .B(n138), .S(n606), .Z(n142) );
  MUX2_X1 U743 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n616), .Z(n143) );
  MUX2_X1 U744 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n616), .Z(n144) );
  MUX2_X1 U745 ( .A(n144), .B(n143), .S(n610), .Z(n145) );
  MUX2_X1 U746 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n616), .Z(n146) );
  MUX2_X1 U747 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n616), .Z(n147) );
  MUX2_X1 U748 ( .A(n147), .B(n146), .S(n610), .Z(n148) );
  MUX2_X1 U749 ( .A(n148), .B(n145), .S(n606), .Z(n149) );
  MUX2_X1 U750 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U751 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U752 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n611), .Z(n151) );
  MUX2_X1 U753 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n611), .Z(n152) );
  MUX2_X1 U754 ( .A(n152), .B(n151), .S(n609), .Z(n153) );
  MUX2_X1 U755 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n611), .Z(n154) );
  MUX2_X1 U756 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n611), .Z(n155) );
  MUX2_X1 U757 ( .A(n155), .B(n154), .S(n609), .Z(n156) );
  MUX2_X1 U758 ( .A(n156), .B(n153), .S(n607), .Z(n157) );
  MUX2_X1 U759 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n611), .Z(n158) );
  MUX2_X1 U760 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n611), .Z(n159) );
  MUX2_X1 U761 ( .A(n159), .B(n158), .S(n610), .Z(n160) );
  MUX2_X1 U762 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n611), .Z(n161) );
  MUX2_X1 U763 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n613), .Z(n162) );
  MUX2_X1 U764 ( .A(n162), .B(n161), .S(n610), .Z(n163) );
  MUX2_X1 U765 ( .A(n163), .B(n160), .S(n607), .Z(n164) );
  MUX2_X1 U766 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U767 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n611), .Z(n166) );
  MUX2_X1 U768 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n611), .Z(n167) );
  MUX2_X1 U769 ( .A(n167), .B(n166), .S(n608), .Z(n168) );
  MUX2_X1 U770 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n611), .Z(n169) );
  MUX2_X1 U771 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n612), .Z(n170) );
  MUX2_X1 U772 ( .A(n170), .B(n169), .S(N11), .Z(n171) );
  MUX2_X1 U773 ( .A(n171), .B(n168), .S(n607), .Z(n172) );
  MUX2_X1 U774 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n613), .Z(n173) );
  MUX2_X1 U775 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n613), .Z(n174) );
  MUX2_X1 U776 ( .A(n174), .B(n173), .S(n608), .Z(n175) );
  MUX2_X1 U777 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n613), .Z(n176) );
  MUX2_X1 U778 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n613), .Z(n177) );
  MUX2_X1 U779 ( .A(n177), .B(n176), .S(n609), .Z(n178) );
  MUX2_X1 U780 ( .A(n178), .B(n175), .S(n607), .Z(n179) );
  MUX2_X1 U781 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U782 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U783 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n613), .Z(n181) );
  MUX2_X1 U784 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n613), .Z(n182) );
  MUX2_X1 U785 ( .A(n182), .B(n181), .S(n608), .Z(n183) );
  MUX2_X1 U786 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n613), .Z(n184) );
  MUX2_X1 U787 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n613), .Z(n185) );
  MUX2_X1 U788 ( .A(n185), .B(n184), .S(n608), .Z(n186) );
  MUX2_X1 U789 ( .A(n186), .B(n183), .S(n607), .Z(n187) );
  MUX2_X1 U790 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n613), .Z(n188) );
  MUX2_X1 U791 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n613), .Z(n189) );
  MUX2_X1 U792 ( .A(n189), .B(n188), .S(n609), .Z(n190) );
  MUX2_X1 U793 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n613), .Z(n191) );
  MUX2_X1 U794 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n613), .Z(n192) );
  MUX2_X1 U795 ( .A(n192), .B(n191), .S(n608), .Z(n193) );
  MUX2_X1 U796 ( .A(n193), .B(n190), .S(n607), .Z(n194) );
  MUX2_X1 U797 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U798 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n614), .Z(n196) );
  MUX2_X1 U799 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n614), .Z(n197) );
  MUX2_X1 U800 ( .A(n197), .B(n196), .S(n610), .Z(n198) );
  MUX2_X1 U801 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n614), .Z(n199) );
  MUX2_X1 U802 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n614), .Z(n200) );
  MUX2_X1 U803 ( .A(n200), .B(n199), .S(n609), .Z(n201) );
  MUX2_X1 U804 ( .A(n201), .B(n198), .S(n607), .Z(n202) );
  MUX2_X1 U805 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n614), .Z(n203) );
  MUX2_X1 U806 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n614), .Z(n204) );
  MUX2_X1 U807 ( .A(n204), .B(n203), .S(N11), .Z(n205) );
  MUX2_X1 U808 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n614), .Z(n206) );
  MUX2_X1 U809 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n614), .Z(n207) );
  MUX2_X1 U810 ( .A(n207), .B(n206), .S(n610), .Z(n208) );
  MUX2_X1 U811 ( .A(n208), .B(n205), .S(n607), .Z(n209) );
  MUX2_X1 U812 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U813 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U814 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n614), .Z(n211) );
  MUX2_X1 U815 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n614), .Z(n212) );
  MUX2_X1 U816 ( .A(n212), .B(n211), .S(n610), .Z(n213) );
  MUX2_X1 U817 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n614), .Z(n214) );
  MUX2_X1 U818 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n614), .Z(n215) );
  MUX2_X1 U819 ( .A(n215), .B(n214), .S(N11), .Z(n216) );
  MUX2_X1 U820 ( .A(n216), .B(n213), .S(n607), .Z(n217) );
  MUX2_X1 U821 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n615), .Z(n218) );
  MUX2_X1 U822 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n615), .Z(n219) );
  MUX2_X1 U823 ( .A(n219), .B(n218), .S(n608), .Z(n220) );
  MUX2_X1 U824 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n615), .Z(n221) );
  MUX2_X1 U825 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n615), .Z(n222) );
  MUX2_X1 U826 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U827 ( .A(n223), .B(n220), .S(n607), .Z(n224) );
  MUX2_X1 U828 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U829 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n615), .Z(n226) );
  MUX2_X1 U830 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n615), .Z(n227) );
  MUX2_X1 U831 ( .A(n227), .B(n226), .S(n609), .Z(n228) );
  MUX2_X1 U832 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n615), .Z(n229) );
  MUX2_X1 U833 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n615), .Z(n595) );
  MUX2_X1 U834 ( .A(n595), .B(n229), .S(N11), .Z(n596) );
  MUX2_X1 U835 ( .A(n596), .B(n228), .S(n607), .Z(n597) );
  MUX2_X1 U836 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n615), .Z(n598) );
  MUX2_X1 U837 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n615), .Z(n599) );
  MUX2_X1 U838 ( .A(n599), .B(n598), .S(n610), .Z(n600) );
  MUX2_X1 U839 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n615), .Z(n601) );
  MUX2_X1 U840 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n615), .Z(n602) );
  MUX2_X1 U841 ( .A(n602), .B(n601), .S(n610), .Z(n603) );
  MUX2_X1 U842 ( .A(n603), .B(n600), .S(n607), .Z(n604) );
  MUX2_X1 U843 ( .A(n604), .B(n597), .S(N13), .Z(n605) );
  MUX2_X1 U844 ( .A(n605), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U845 ( .A(N11), .Z(n608) );
  INV_X1 U846 ( .A(N10), .ZN(n617) );
  INV_X1 U847 ( .A(N11), .ZN(n618) );
  INV_X1 U848 ( .A(data_in[0]), .ZN(n619) );
  INV_X1 U849 ( .A(data_in[1]), .ZN(n620) );
  INV_X1 U850 ( .A(data_in[2]), .ZN(n621) );
  INV_X1 U851 ( .A(data_in[3]), .ZN(n622) );
  INV_X1 U852 ( .A(data_in[4]), .ZN(n623) );
  INV_X1 U853 ( .A(data_in[5]), .ZN(n624) );
  INV_X1 U854 ( .A(data_in[6]), .ZN(n625) );
  INV_X1 U855 ( .A(data_in[7]), .ZN(n626) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_13 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .QN(n2) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n630), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n631), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n632), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n633), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n634), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n635), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n636), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n637), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n638), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n639), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n640), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n641), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n642), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n643), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n644), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n645), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n646), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n647), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n648), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n649), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n650), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n651), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n652), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n653), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n654), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n655), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n656), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n657), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n658), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n659), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n660), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n661), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n662), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n663), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n664), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n665), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n666), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n667), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n668), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n669), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n670), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n671), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n672), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n673), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n674), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n675), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n676), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n677), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n678), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n679), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n680), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n681), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n682), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n683), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n684), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n685), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n686), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n687), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n688), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n689), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n690), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n691), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n692), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n693), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n694), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n695), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n696), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n697), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n698), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n699), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n700), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n701), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n702), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n703), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n704), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n705), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n706), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n707), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n708), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n709), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n710), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n711), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n712), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n713), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n714), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n715), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n716), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n717), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n718), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n719), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n720), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n721), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n722), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n723), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n724), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n725), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n726), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n727), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n728), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n729), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n730), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n731), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n732), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n733), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n734), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n735), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n736), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n737), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n738), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n739), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n740), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n741), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n742), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n743), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n744), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n745), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n746), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n747), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n748), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n749), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n750), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n751), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n752), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n753), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n754), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n755), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n756), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n757), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n758), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n759), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n760), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n761), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n762), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n763), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n764), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n765), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n766), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n767), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n768), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n769), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n770), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n771), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n772), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n773), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n774), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n775), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n776), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n777), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n778), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n779), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n780), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n781), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n782), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n783), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n784), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n785), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n786), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n787), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n788), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n789), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n790), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n791), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n792), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n793), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n794), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n795), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n796), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n797), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n798), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n799), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n800), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n801), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n802), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n803), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n804), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n805), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n806), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n807), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n808), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n809), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n810), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n811), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n812), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n813), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n814), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n815), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n816), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n817), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n818), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n819), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n820), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n821), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n849), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n850), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n851), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n852), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n853), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n854), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n855), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n856), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n857), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n858), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n859), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n860), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n861), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n862), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n863), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n864), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n865), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n866), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n867), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n868), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n869), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n870), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n871), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n872), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n873), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n874), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n875), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n876), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n877), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n878), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n879), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n880), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n881), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n882), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n883), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n884), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n885), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n886), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n887), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n888), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n889), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n890), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n891), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n892), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n893), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n894), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n895), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n896), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n897), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n898), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n899), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n900), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n901), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n902), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n903), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n904), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n905), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n906), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n907), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n908), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n909), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n910), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n911), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n912), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  INV_X2 U3 ( .A(n2), .ZN(data_out[5]) );
  BUF_X1 U4 ( .A(n619), .Z(n617) );
  BUF_X1 U5 ( .A(n619), .Z(n618) );
  BUF_X1 U6 ( .A(N10), .Z(n614) );
  BUF_X1 U7 ( .A(n619), .Z(n615) );
  BUF_X1 U8 ( .A(n619), .Z(n616) );
  BUF_X1 U9 ( .A(N11), .Z(n612) );
  BUF_X1 U10 ( .A(N11), .Z(n613) );
  BUF_X1 U11 ( .A(N10), .Z(n619) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1204) );
  NOR3_X1 U13 ( .A1(N11), .A2(N12), .A3(n620), .ZN(n1193) );
  NOR3_X1 U14 ( .A1(N10), .A2(N12), .A3(n621), .ZN(n1183) );
  NOR3_X1 U15 ( .A1(n620), .A2(N12), .A3(n621), .ZN(n1173) );
  INV_X1 U16 ( .A(n1130), .ZN(n845) );
  INV_X1 U17 ( .A(n1120), .ZN(n844) );
  INV_X1 U18 ( .A(n1111), .ZN(n843) );
  INV_X1 U19 ( .A(n1102), .ZN(n842) );
  INV_X1 U20 ( .A(n1057), .ZN(n837) );
  INV_X1 U21 ( .A(n1047), .ZN(n836) );
  INV_X1 U22 ( .A(n1038), .ZN(n835) );
  INV_X1 U23 ( .A(n1029), .ZN(n834) );
  INV_X1 U24 ( .A(n984), .ZN(n829) );
  INV_X1 U25 ( .A(n974), .ZN(n828) );
  INV_X1 U26 ( .A(n965), .ZN(n827) );
  INV_X1 U27 ( .A(n956), .ZN(n826) );
  INV_X1 U28 ( .A(n947), .ZN(n825) );
  INV_X1 U29 ( .A(n938), .ZN(n824) );
  INV_X1 U30 ( .A(n929), .ZN(n823) );
  INV_X1 U31 ( .A(n920), .ZN(n822) );
  INV_X1 U32 ( .A(n1093), .ZN(n841) );
  INV_X1 U33 ( .A(n1084), .ZN(n840) );
  INV_X1 U34 ( .A(n1075), .ZN(n839) );
  INV_X1 U35 ( .A(n1066), .ZN(n838) );
  INV_X1 U36 ( .A(n1020), .ZN(n833) );
  INV_X1 U37 ( .A(n1011), .ZN(n832) );
  INV_X1 U38 ( .A(n1002), .ZN(n831) );
  INV_X1 U39 ( .A(n993), .ZN(n830) );
  BUF_X1 U40 ( .A(N12), .Z(n609) );
  BUF_X1 U41 ( .A(N12), .Z(n610) );
  INV_X1 U42 ( .A(N13), .ZN(n847) );
  AND3_X1 U43 ( .A1(n620), .A2(n621), .A3(N12), .ZN(n1163) );
  AND3_X1 U44 ( .A1(N10), .A2(n621), .A3(N12), .ZN(n1153) );
  AND3_X1 U45 ( .A1(N11), .A2(n620), .A3(N12), .ZN(n1143) );
  AND3_X1 U46 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1133) );
  INV_X1 U47 ( .A(N14), .ZN(n848) );
  NAND2_X1 U48 ( .A1(n1193), .A2(n1203), .ZN(n1202) );
  NAND2_X1 U49 ( .A1(n1183), .A2(n1203), .ZN(n1192) );
  NAND2_X1 U50 ( .A1(n1173), .A2(n1203), .ZN(n1182) );
  NAND2_X1 U51 ( .A1(n1163), .A2(n1203), .ZN(n1172) );
  NAND2_X1 U52 ( .A1(n1153), .A2(n1203), .ZN(n1162) );
  NAND2_X1 U53 ( .A1(n1143), .A2(n1203), .ZN(n1152) );
  NAND2_X1 U54 ( .A1(n1133), .A2(n1203), .ZN(n1142) );
  NAND2_X1 U55 ( .A1(n1204), .A2(n1203), .ZN(n1213) );
  NAND2_X1 U56 ( .A1(n1122), .A2(n1204), .ZN(n1130) );
  NAND2_X1 U57 ( .A1(n1122), .A2(n1193), .ZN(n1120) );
  NAND2_X1 U58 ( .A1(n1122), .A2(n1183), .ZN(n1111) );
  NAND2_X1 U59 ( .A1(n1122), .A2(n1173), .ZN(n1102) );
  NAND2_X1 U60 ( .A1(n1049), .A2(n1204), .ZN(n1057) );
  NAND2_X1 U61 ( .A1(n1049), .A2(n1193), .ZN(n1047) );
  NAND2_X1 U62 ( .A1(n1049), .A2(n1183), .ZN(n1038) );
  NAND2_X1 U63 ( .A1(n1049), .A2(n1173), .ZN(n1029) );
  NAND2_X1 U64 ( .A1(n976), .A2(n1204), .ZN(n984) );
  NAND2_X1 U65 ( .A1(n976), .A2(n1193), .ZN(n974) );
  NAND2_X1 U66 ( .A1(n976), .A2(n1183), .ZN(n965) );
  NAND2_X1 U67 ( .A1(n976), .A2(n1173), .ZN(n956) );
  NAND2_X1 U68 ( .A1(n1122), .A2(n1163), .ZN(n1093) );
  NAND2_X1 U69 ( .A1(n1122), .A2(n1153), .ZN(n1084) );
  NAND2_X1 U70 ( .A1(n1122), .A2(n1143), .ZN(n1075) );
  NAND2_X1 U71 ( .A1(n1122), .A2(n1133), .ZN(n1066) );
  NAND2_X1 U72 ( .A1(n1049), .A2(n1163), .ZN(n1020) );
  NAND2_X1 U73 ( .A1(n1049), .A2(n1153), .ZN(n1011) );
  NAND2_X1 U74 ( .A1(n1049), .A2(n1143), .ZN(n1002) );
  NAND2_X1 U75 ( .A1(n1049), .A2(n1133), .ZN(n993) );
  NAND2_X1 U76 ( .A1(n976), .A2(n1163), .ZN(n947) );
  NAND2_X1 U77 ( .A1(n976), .A2(n1153), .ZN(n938) );
  NAND2_X1 U78 ( .A1(n976), .A2(n1143), .ZN(n929) );
  NAND2_X1 U79 ( .A1(n976), .A2(n1133), .ZN(n920) );
  AND3_X1 U80 ( .A1(n847), .A2(n848), .A3(n1132), .ZN(n1203) );
  AND3_X1 U81 ( .A1(N13), .A2(n1132), .A3(N14), .ZN(n976) );
  AND3_X1 U82 ( .A1(n1132), .A2(n848), .A3(N13), .ZN(n1122) );
  AND3_X1 U83 ( .A1(n1132), .A2(n847), .A3(N14), .ZN(n1049) );
  NOR2_X1 U84 ( .A1(n846), .A2(addr[5]), .ZN(n1132) );
  INV_X1 U85 ( .A(wr_en), .ZN(n846) );
  OAI21_X1 U86 ( .B1(n622), .B2(n1172), .A(n1171), .ZN(n880) );
  NAND2_X1 U87 ( .A1(\mem[4][0] ), .A2(n1172), .ZN(n1171) );
  OAI21_X1 U88 ( .B1(n623), .B2(n1172), .A(n1170), .ZN(n879) );
  NAND2_X1 U89 ( .A1(\mem[4][1] ), .A2(n1172), .ZN(n1170) );
  OAI21_X1 U90 ( .B1(n624), .B2(n1172), .A(n1169), .ZN(n878) );
  NAND2_X1 U91 ( .A1(\mem[4][2] ), .A2(n1172), .ZN(n1169) );
  OAI21_X1 U92 ( .B1(n625), .B2(n1172), .A(n1168), .ZN(n877) );
  NAND2_X1 U93 ( .A1(\mem[4][3] ), .A2(n1172), .ZN(n1168) );
  OAI21_X1 U94 ( .B1(n626), .B2(n1172), .A(n1167), .ZN(n876) );
  NAND2_X1 U95 ( .A1(\mem[4][4] ), .A2(n1172), .ZN(n1167) );
  OAI21_X1 U96 ( .B1(n627), .B2(n1172), .A(n1166), .ZN(n875) );
  NAND2_X1 U97 ( .A1(\mem[4][5] ), .A2(n1172), .ZN(n1166) );
  OAI21_X1 U98 ( .B1(n628), .B2(n1172), .A(n1165), .ZN(n874) );
  NAND2_X1 U99 ( .A1(\mem[4][6] ), .A2(n1172), .ZN(n1165) );
  OAI21_X1 U100 ( .B1(n629), .B2(n1172), .A(n1164), .ZN(n873) );
  NAND2_X1 U101 ( .A1(\mem[4][7] ), .A2(n1172), .ZN(n1164) );
  OAI21_X1 U102 ( .B1(n622), .B2(n1152), .A(n1151), .ZN(n864) );
  NAND2_X1 U103 ( .A1(\mem[6][0] ), .A2(n1152), .ZN(n1151) );
  OAI21_X1 U104 ( .B1(n623), .B2(n1152), .A(n1150), .ZN(n863) );
  NAND2_X1 U105 ( .A1(\mem[6][1] ), .A2(n1152), .ZN(n1150) );
  OAI21_X1 U106 ( .B1(n624), .B2(n1152), .A(n1149), .ZN(n862) );
  NAND2_X1 U107 ( .A1(\mem[6][2] ), .A2(n1152), .ZN(n1149) );
  OAI21_X1 U108 ( .B1(n625), .B2(n1152), .A(n1148), .ZN(n861) );
  NAND2_X1 U109 ( .A1(\mem[6][3] ), .A2(n1152), .ZN(n1148) );
  OAI21_X1 U110 ( .B1(n626), .B2(n1152), .A(n1147), .ZN(n860) );
  NAND2_X1 U111 ( .A1(\mem[6][4] ), .A2(n1152), .ZN(n1147) );
  OAI21_X1 U112 ( .B1(n627), .B2(n1152), .A(n1146), .ZN(n859) );
  NAND2_X1 U113 ( .A1(\mem[6][5] ), .A2(n1152), .ZN(n1146) );
  OAI21_X1 U114 ( .B1(n628), .B2(n1152), .A(n1145), .ZN(n858) );
  NAND2_X1 U115 ( .A1(\mem[6][6] ), .A2(n1152), .ZN(n1145) );
  OAI21_X1 U116 ( .B1(n629), .B2(n1152), .A(n1144), .ZN(n857) );
  NAND2_X1 U117 ( .A1(\mem[6][7] ), .A2(n1152), .ZN(n1144) );
  OAI21_X1 U118 ( .B1(n622), .B2(n1142), .A(n1141), .ZN(n856) );
  NAND2_X1 U119 ( .A1(\mem[7][0] ), .A2(n1142), .ZN(n1141) );
  OAI21_X1 U120 ( .B1(n623), .B2(n1142), .A(n1140), .ZN(n855) );
  NAND2_X1 U121 ( .A1(\mem[7][1] ), .A2(n1142), .ZN(n1140) );
  OAI21_X1 U122 ( .B1(n624), .B2(n1142), .A(n1139), .ZN(n854) );
  NAND2_X1 U123 ( .A1(\mem[7][2] ), .A2(n1142), .ZN(n1139) );
  OAI21_X1 U124 ( .B1(n625), .B2(n1142), .A(n1138), .ZN(n853) );
  NAND2_X1 U125 ( .A1(\mem[7][3] ), .A2(n1142), .ZN(n1138) );
  OAI21_X1 U126 ( .B1(n626), .B2(n1142), .A(n1137), .ZN(n852) );
  NAND2_X1 U127 ( .A1(\mem[7][4] ), .A2(n1142), .ZN(n1137) );
  OAI21_X1 U128 ( .B1(n627), .B2(n1142), .A(n1136), .ZN(n851) );
  NAND2_X1 U129 ( .A1(\mem[7][5] ), .A2(n1142), .ZN(n1136) );
  OAI21_X1 U130 ( .B1(n628), .B2(n1142), .A(n1135), .ZN(n850) );
  NAND2_X1 U131 ( .A1(\mem[7][6] ), .A2(n1142), .ZN(n1135) );
  OAI21_X1 U132 ( .B1(n629), .B2(n1142), .A(n1134), .ZN(n849) );
  NAND2_X1 U133 ( .A1(\mem[7][7] ), .A2(n1142), .ZN(n1134) );
  OAI21_X1 U134 ( .B1(n622), .B2(n1202), .A(n1201), .ZN(n904) );
  NAND2_X1 U135 ( .A1(\mem[1][0] ), .A2(n1202), .ZN(n1201) );
  OAI21_X1 U136 ( .B1(n623), .B2(n1202), .A(n1200), .ZN(n903) );
  NAND2_X1 U137 ( .A1(\mem[1][1] ), .A2(n1202), .ZN(n1200) );
  OAI21_X1 U138 ( .B1(n624), .B2(n1202), .A(n1199), .ZN(n902) );
  NAND2_X1 U139 ( .A1(\mem[1][2] ), .A2(n1202), .ZN(n1199) );
  OAI21_X1 U140 ( .B1(n625), .B2(n1202), .A(n1198), .ZN(n901) );
  NAND2_X1 U141 ( .A1(\mem[1][3] ), .A2(n1202), .ZN(n1198) );
  OAI21_X1 U142 ( .B1(n626), .B2(n1202), .A(n1197), .ZN(n900) );
  NAND2_X1 U143 ( .A1(\mem[1][4] ), .A2(n1202), .ZN(n1197) );
  OAI21_X1 U144 ( .B1(n627), .B2(n1202), .A(n1196), .ZN(n899) );
  NAND2_X1 U145 ( .A1(\mem[1][5] ), .A2(n1202), .ZN(n1196) );
  OAI21_X1 U146 ( .B1(n628), .B2(n1202), .A(n1195), .ZN(n898) );
  NAND2_X1 U147 ( .A1(\mem[1][6] ), .A2(n1202), .ZN(n1195) );
  OAI21_X1 U148 ( .B1(n629), .B2(n1202), .A(n1194), .ZN(n897) );
  NAND2_X1 U149 ( .A1(\mem[1][7] ), .A2(n1202), .ZN(n1194) );
  OAI21_X1 U150 ( .B1(n622), .B2(n1192), .A(n1191), .ZN(n896) );
  NAND2_X1 U151 ( .A1(\mem[2][0] ), .A2(n1192), .ZN(n1191) );
  OAI21_X1 U152 ( .B1(n623), .B2(n1192), .A(n1190), .ZN(n895) );
  NAND2_X1 U153 ( .A1(\mem[2][1] ), .A2(n1192), .ZN(n1190) );
  OAI21_X1 U154 ( .B1(n624), .B2(n1192), .A(n1189), .ZN(n894) );
  NAND2_X1 U155 ( .A1(\mem[2][2] ), .A2(n1192), .ZN(n1189) );
  OAI21_X1 U156 ( .B1(n625), .B2(n1192), .A(n1188), .ZN(n893) );
  NAND2_X1 U157 ( .A1(\mem[2][3] ), .A2(n1192), .ZN(n1188) );
  OAI21_X1 U158 ( .B1(n626), .B2(n1192), .A(n1187), .ZN(n892) );
  NAND2_X1 U159 ( .A1(\mem[2][4] ), .A2(n1192), .ZN(n1187) );
  OAI21_X1 U160 ( .B1(n627), .B2(n1192), .A(n1186), .ZN(n891) );
  NAND2_X1 U161 ( .A1(\mem[2][5] ), .A2(n1192), .ZN(n1186) );
  OAI21_X1 U162 ( .B1(n628), .B2(n1192), .A(n1185), .ZN(n890) );
  NAND2_X1 U163 ( .A1(\mem[2][6] ), .A2(n1192), .ZN(n1185) );
  OAI21_X1 U164 ( .B1(n629), .B2(n1192), .A(n1184), .ZN(n889) );
  NAND2_X1 U165 ( .A1(\mem[2][7] ), .A2(n1192), .ZN(n1184) );
  OAI21_X1 U166 ( .B1(n622), .B2(n1182), .A(n1181), .ZN(n888) );
  NAND2_X1 U167 ( .A1(\mem[3][0] ), .A2(n1182), .ZN(n1181) );
  OAI21_X1 U168 ( .B1(n623), .B2(n1182), .A(n1180), .ZN(n887) );
  NAND2_X1 U169 ( .A1(\mem[3][1] ), .A2(n1182), .ZN(n1180) );
  OAI21_X1 U170 ( .B1(n624), .B2(n1182), .A(n1179), .ZN(n886) );
  NAND2_X1 U171 ( .A1(\mem[3][2] ), .A2(n1182), .ZN(n1179) );
  OAI21_X1 U172 ( .B1(n625), .B2(n1182), .A(n1178), .ZN(n885) );
  NAND2_X1 U173 ( .A1(\mem[3][3] ), .A2(n1182), .ZN(n1178) );
  OAI21_X1 U174 ( .B1(n626), .B2(n1182), .A(n1177), .ZN(n884) );
  NAND2_X1 U175 ( .A1(\mem[3][4] ), .A2(n1182), .ZN(n1177) );
  OAI21_X1 U176 ( .B1(n627), .B2(n1182), .A(n1176), .ZN(n883) );
  NAND2_X1 U177 ( .A1(\mem[3][5] ), .A2(n1182), .ZN(n1176) );
  OAI21_X1 U178 ( .B1(n628), .B2(n1182), .A(n1175), .ZN(n882) );
  NAND2_X1 U179 ( .A1(\mem[3][6] ), .A2(n1182), .ZN(n1175) );
  OAI21_X1 U180 ( .B1(n629), .B2(n1182), .A(n1174), .ZN(n881) );
  NAND2_X1 U181 ( .A1(\mem[3][7] ), .A2(n1182), .ZN(n1174) );
  OAI21_X1 U182 ( .B1(n622), .B2(n1162), .A(n1161), .ZN(n872) );
  NAND2_X1 U183 ( .A1(\mem[5][0] ), .A2(n1162), .ZN(n1161) );
  OAI21_X1 U184 ( .B1(n623), .B2(n1162), .A(n1160), .ZN(n871) );
  NAND2_X1 U185 ( .A1(\mem[5][1] ), .A2(n1162), .ZN(n1160) );
  OAI21_X1 U186 ( .B1(n624), .B2(n1162), .A(n1159), .ZN(n870) );
  NAND2_X1 U187 ( .A1(\mem[5][2] ), .A2(n1162), .ZN(n1159) );
  OAI21_X1 U188 ( .B1(n625), .B2(n1162), .A(n1158), .ZN(n869) );
  NAND2_X1 U189 ( .A1(\mem[5][3] ), .A2(n1162), .ZN(n1158) );
  OAI21_X1 U190 ( .B1(n626), .B2(n1162), .A(n1157), .ZN(n868) );
  NAND2_X1 U191 ( .A1(\mem[5][4] ), .A2(n1162), .ZN(n1157) );
  OAI21_X1 U192 ( .B1(n627), .B2(n1162), .A(n1156), .ZN(n867) );
  NAND2_X1 U193 ( .A1(\mem[5][5] ), .A2(n1162), .ZN(n1156) );
  OAI21_X1 U194 ( .B1(n628), .B2(n1162), .A(n1155), .ZN(n866) );
  NAND2_X1 U195 ( .A1(\mem[5][6] ), .A2(n1162), .ZN(n1155) );
  OAI21_X1 U196 ( .B1(n629), .B2(n1162), .A(n1154), .ZN(n865) );
  NAND2_X1 U197 ( .A1(\mem[5][7] ), .A2(n1162), .ZN(n1154) );
  OAI21_X1 U198 ( .B1(n1213), .B2(n622), .A(n1212), .ZN(n912) );
  NAND2_X1 U199 ( .A1(\mem[0][0] ), .A2(n1213), .ZN(n1212) );
  OAI21_X1 U200 ( .B1(n1213), .B2(n623), .A(n1211), .ZN(n911) );
  NAND2_X1 U201 ( .A1(\mem[0][1] ), .A2(n1213), .ZN(n1211) );
  OAI21_X1 U202 ( .B1(n1213), .B2(n624), .A(n1210), .ZN(n910) );
  NAND2_X1 U203 ( .A1(\mem[0][2] ), .A2(n1213), .ZN(n1210) );
  OAI21_X1 U204 ( .B1(n1213), .B2(n625), .A(n1209), .ZN(n909) );
  NAND2_X1 U205 ( .A1(\mem[0][3] ), .A2(n1213), .ZN(n1209) );
  OAI21_X1 U206 ( .B1(n1213), .B2(n626), .A(n1208), .ZN(n908) );
  NAND2_X1 U207 ( .A1(\mem[0][4] ), .A2(n1213), .ZN(n1208) );
  OAI21_X1 U208 ( .B1(n1213), .B2(n627), .A(n1207), .ZN(n907) );
  NAND2_X1 U209 ( .A1(\mem[0][5] ), .A2(n1213), .ZN(n1207) );
  OAI21_X1 U210 ( .B1(n1213), .B2(n628), .A(n1206), .ZN(n906) );
  NAND2_X1 U211 ( .A1(\mem[0][6] ), .A2(n1213), .ZN(n1206) );
  OAI21_X1 U212 ( .B1(n1213), .B2(n629), .A(n1205), .ZN(n905) );
  NAND2_X1 U213 ( .A1(\mem[0][7] ), .A2(n1213), .ZN(n1205) );
  INV_X1 U214 ( .A(n1131), .ZN(n821) );
  AOI22_X1 U215 ( .A1(data_in[0]), .A2(n845), .B1(n1130), .B2(\mem[8][0] ), 
        .ZN(n1131) );
  INV_X1 U216 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U217 ( .A1(data_in[1]), .A2(n845), .B1(n1130), .B2(\mem[8][1] ), 
        .ZN(n1129) );
  INV_X1 U218 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U219 ( .A1(data_in[2]), .A2(n845), .B1(n1130), .B2(\mem[8][2] ), 
        .ZN(n1128) );
  INV_X1 U220 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U221 ( .A1(data_in[3]), .A2(n845), .B1(n1130), .B2(\mem[8][3] ), 
        .ZN(n1127) );
  INV_X1 U222 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U223 ( .A1(data_in[4]), .A2(n845), .B1(n1130), .B2(\mem[8][4] ), 
        .ZN(n1126) );
  INV_X1 U224 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U225 ( .A1(data_in[5]), .A2(n845), .B1(n1130), .B2(\mem[8][5] ), 
        .ZN(n1125) );
  INV_X1 U226 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U227 ( .A1(data_in[6]), .A2(n845), .B1(n1130), .B2(\mem[8][6] ), 
        .ZN(n1124) );
  INV_X1 U228 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U229 ( .A1(data_in[7]), .A2(n845), .B1(n1130), .B2(\mem[8][7] ), 
        .ZN(n1123) );
  INV_X1 U230 ( .A(n1121), .ZN(n813) );
  AOI22_X1 U231 ( .A1(data_in[0]), .A2(n844), .B1(n1120), .B2(\mem[9][0] ), 
        .ZN(n1121) );
  INV_X1 U232 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U233 ( .A1(data_in[1]), .A2(n844), .B1(n1120), .B2(\mem[9][1] ), 
        .ZN(n1119) );
  INV_X1 U234 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U235 ( .A1(data_in[2]), .A2(n844), .B1(n1120), .B2(\mem[9][2] ), 
        .ZN(n1118) );
  INV_X1 U236 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U237 ( .A1(data_in[3]), .A2(n844), .B1(n1120), .B2(\mem[9][3] ), 
        .ZN(n1117) );
  INV_X1 U238 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U239 ( .A1(data_in[4]), .A2(n844), .B1(n1120), .B2(\mem[9][4] ), 
        .ZN(n1116) );
  INV_X1 U240 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U241 ( .A1(data_in[5]), .A2(n844), .B1(n1120), .B2(\mem[9][5] ), 
        .ZN(n1115) );
  INV_X1 U242 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U243 ( .A1(data_in[6]), .A2(n844), .B1(n1120), .B2(\mem[9][6] ), 
        .ZN(n1114) );
  INV_X1 U244 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U245 ( .A1(data_in[7]), .A2(n844), .B1(n1120), .B2(\mem[9][7] ), 
        .ZN(n1113) );
  INV_X1 U246 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U247 ( .A1(data_in[0]), .A2(n843), .B1(n1111), .B2(\mem[10][0] ), 
        .ZN(n1112) );
  INV_X1 U248 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U249 ( .A1(data_in[1]), .A2(n843), .B1(n1111), .B2(\mem[10][1] ), 
        .ZN(n1110) );
  INV_X1 U250 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U251 ( .A1(data_in[2]), .A2(n843), .B1(n1111), .B2(\mem[10][2] ), 
        .ZN(n1109) );
  INV_X1 U252 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U253 ( .A1(data_in[3]), .A2(n843), .B1(n1111), .B2(\mem[10][3] ), 
        .ZN(n1108) );
  INV_X1 U254 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U255 ( .A1(data_in[4]), .A2(n843), .B1(n1111), .B2(\mem[10][4] ), 
        .ZN(n1107) );
  INV_X1 U256 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U257 ( .A1(data_in[5]), .A2(n843), .B1(n1111), .B2(\mem[10][5] ), 
        .ZN(n1106) );
  INV_X1 U258 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U259 ( .A1(data_in[6]), .A2(n843), .B1(n1111), .B2(\mem[10][6] ), 
        .ZN(n1105) );
  INV_X1 U260 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U261 ( .A1(data_in[7]), .A2(n843), .B1(n1111), .B2(\mem[10][7] ), 
        .ZN(n1104) );
  INV_X1 U262 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U263 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[11][0] ), 
        .ZN(n1103) );
  INV_X1 U264 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U265 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[11][1] ), 
        .ZN(n1101) );
  INV_X1 U266 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U267 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[11][2] ), 
        .ZN(n1100) );
  INV_X1 U268 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U269 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[11][3] ), 
        .ZN(n1099) );
  INV_X1 U270 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U271 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[11][4] ), 
        .ZN(n1098) );
  INV_X1 U272 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U273 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[11][5] ), 
        .ZN(n1097) );
  INV_X1 U274 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U275 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[11][6] ), 
        .ZN(n1096) );
  INV_X1 U276 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U277 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[11][7] ), 
        .ZN(n1095) );
  INV_X1 U278 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U279 ( .A1(data_in[0]), .A2(n841), .B1(n1093), .B2(\mem[12][0] ), 
        .ZN(n1094) );
  INV_X1 U280 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U281 ( .A1(data_in[1]), .A2(n841), .B1(n1093), .B2(\mem[12][1] ), 
        .ZN(n1092) );
  INV_X1 U282 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U283 ( .A1(data_in[2]), .A2(n841), .B1(n1093), .B2(\mem[12][2] ), 
        .ZN(n1091) );
  INV_X1 U284 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U285 ( .A1(data_in[3]), .A2(n841), .B1(n1093), .B2(\mem[12][3] ), 
        .ZN(n1090) );
  INV_X1 U286 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U287 ( .A1(data_in[4]), .A2(n841), .B1(n1093), .B2(\mem[12][4] ), 
        .ZN(n1089) );
  INV_X1 U288 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U289 ( .A1(data_in[5]), .A2(n841), .B1(n1093), .B2(\mem[12][5] ), 
        .ZN(n1088) );
  INV_X1 U290 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U291 ( .A1(data_in[6]), .A2(n841), .B1(n1093), .B2(\mem[12][6] ), 
        .ZN(n1087) );
  INV_X1 U292 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U293 ( .A1(data_in[7]), .A2(n841), .B1(n1093), .B2(\mem[12][7] ), 
        .ZN(n1086) );
  INV_X1 U294 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U295 ( .A1(data_in[0]), .A2(n840), .B1(n1084), .B2(\mem[13][0] ), 
        .ZN(n1085) );
  INV_X1 U296 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U297 ( .A1(data_in[1]), .A2(n840), .B1(n1084), .B2(\mem[13][1] ), 
        .ZN(n1083) );
  INV_X1 U298 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U299 ( .A1(data_in[2]), .A2(n840), .B1(n1084), .B2(\mem[13][2] ), 
        .ZN(n1082) );
  INV_X1 U300 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U301 ( .A1(data_in[3]), .A2(n840), .B1(n1084), .B2(\mem[13][3] ), 
        .ZN(n1081) );
  INV_X1 U302 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U303 ( .A1(data_in[4]), .A2(n840), .B1(n1084), .B2(\mem[13][4] ), 
        .ZN(n1080) );
  INV_X1 U304 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U305 ( .A1(data_in[5]), .A2(n840), .B1(n1084), .B2(\mem[13][5] ), 
        .ZN(n1079) );
  INV_X1 U306 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U307 ( .A1(data_in[6]), .A2(n840), .B1(n1084), .B2(\mem[13][6] ), 
        .ZN(n1078) );
  INV_X1 U308 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U309 ( .A1(data_in[7]), .A2(n840), .B1(n1084), .B2(\mem[13][7] ), 
        .ZN(n1077) );
  INV_X1 U310 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U311 ( .A1(data_in[0]), .A2(n839), .B1(n1075), .B2(\mem[14][0] ), 
        .ZN(n1076) );
  INV_X1 U312 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U313 ( .A1(data_in[1]), .A2(n839), .B1(n1075), .B2(\mem[14][1] ), 
        .ZN(n1074) );
  INV_X1 U314 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U315 ( .A1(data_in[2]), .A2(n839), .B1(n1075), .B2(\mem[14][2] ), 
        .ZN(n1073) );
  INV_X1 U316 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U317 ( .A1(data_in[3]), .A2(n839), .B1(n1075), .B2(\mem[14][3] ), 
        .ZN(n1072) );
  INV_X1 U318 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U319 ( .A1(data_in[4]), .A2(n839), .B1(n1075), .B2(\mem[14][4] ), 
        .ZN(n1071) );
  INV_X1 U320 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U321 ( .A1(data_in[5]), .A2(n839), .B1(n1075), .B2(\mem[14][5] ), 
        .ZN(n1070) );
  INV_X1 U322 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U323 ( .A1(data_in[6]), .A2(n839), .B1(n1075), .B2(\mem[14][6] ), 
        .ZN(n1069) );
  INV_X1 U324 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U325 ( .A1(data_in[7]), .A2(n839), .B1(n1075), .B2(\mem[14][7] ), 
        .ZN(n1068) );
  INV_X1 U326 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U327 ( .A1(data_in[0]), .A2(n838), .B1(n1066), .B2(\mem[15][0] ), 
        .ZN(n1067) );
  INV_X1 U328 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U329 ( .A1(data_in[1]), .A2(n838), .B1(n1066), .B2(\mem[15][1] ), 
        .ZN(n1065) );
  INV_X1 U330 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U331 ( .A1(data_in[2]), .A2(n838), .B1(n1066), .B2(\mem[15][2] ), 
        .ZN(n1064) );
  INV_X1 U332 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U333 ( .A1(data_in[3]), .A2(n838), .B1(n1066), .B2(\mem[15][3] ), 
        .ZN(n1063) );
  INV_X1 U334 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U335 ( .A1(data_in[4]), .A2(n838), .B1(n1066), .B2(\mem[15][4] ), 
        .ZN(n1062) );
  INV_X1 U336 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U337 ( .A1(data_in[5]), .A2(n838), .B1(n1066), .B2(\mem[15][5] ), 
        .ZN(n1061) );
  INV_X1 U338 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U339 ( .A1(data_in[6]), .A2(n838), .B1(n1066), .B2(\mem[15][6] ), 
        .ZN(n1060) );
  INV_X1 U340 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U341 ( .A1(data_in[7]), .A2(n838), .B1(n1066), .B2(\mem[15][7] ), 
        .ZN(n1059) );
  INV_X1 U342 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U343 ( .A1(data_in[0]), .A2(n837), .B1(n1057), .B2(\mem[16][0] ), 
        .ZN(n1058) );
  INV_X1 U344 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U345 ( .A1(data_in[1]), .A2(n837), .B1(n1057), .B2(\mem[16][1] ), 
        .ZN(n1056) );
  INV_X1 U346 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U347 ( .A1(data_in[2]), .A2(n837), .B1(n1057), .B2(\mem[16][2] ), 
        .ZN(n1055) );
  INV_X1 U348 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U349 ( .A1(data_in[3]), .A2(n837), .B1(n1057), .B2(\mem[16][3] ), 
        .ZN(n1054) );
  INV_X1 U350 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U351 ( .A1(data_in[4]), .A2(n837), .B1(n1057), .B2(\mem[16][4] ), 
        .ZN(n1053) );
  INV_X1 U352 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U353 ( .A1(data_in[5]), .A2(n837), .B1(n1057), .B2(\mem[16][5] ), 
        .ZN(n1052) );
  INV_X1 U354 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U355 ( .A1(data_in[6]), .A2(n837), .B1(n1057), .B2(\mem[16][6] ), 
        .ZN(n1051) );
  INV_X1 U356 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U357 ( .A1(data_in[7]), .A2(n837), .B1(n1057), .B2(\mem[16][7] ), 
        .ZN(n1050) );
  INV_X1 U358 ( .A(n1048), .ZN(n749) );
  AOI22_X1 U359 ( .A1(data_in[0]), .A2(n836), .B1(n1047), .B2(\mem[17][0] ), 
        .ZN(n1048) );
  INV_X1 U360 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U361 ( .A1(data_in[1]), .A2(n836), .B1(n1047), .B2(\mem[17][1] ), 
        .ZN(n1046) );
  INV_X1 U362 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U363 ( .A1(data_in[2]), .A2(n836), .B1(n1047), .B2(\mem[17][2] ), 
        .ZN(n1045) );
  INV_X1 U364 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U365 ( .A1(data_in[3]), .A2(n836), .B1(n1047), .B2(\mem[17][3] ), 
        .ZN(n1044) );
  INV_X1 U366 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U367 ( .A1(data_in[4]), .A2(n836), .B1(n1047), .B2(\mem[17][4] ), 
        .ZN(n1043) );
  INV_X1 U368 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U369 ( .A1(data_in[5]), .A2(n836), .B1(n1047), .B2(\mem[17][5] ), 
        .ZN(n1042) );
  INV_X1 U370 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U371 ( .A1(data_in[6]), .A2(n836), .B1(n1047), .B2(\mem[17][6] ), 
        .ZN(n1041) );
  INV_X1 U372 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U373 ( .A1(data_in[7]), .A2(n836), .B1(n1047), .B2(\mem[17][7] ), 
        .ZN(n1040) );
  INV_X1 U374 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U375 ( .A1(data_in[0]), .A2(n835), .B1(n1038), .B2(\mem[18][0] ), 
        .ZN(n1039) );
  INV_X1 U376 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U377 ( .A1(data_in[1]), .A2(n835), .B1(n1038), .B2(\mem[18][1] ), 
        .ZN(n1037) );
  INV_X1 U378 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U379 ( .A1(data_in[2]), .A2(n835), .B1(n1038), .B2(\mem[18][2] ), 
        .ZN(n1036) );
  INV_X1 U380 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U381 ( .A1(data_in[3]), .A2(n835), .B1(n1038), .B2(\mem[18][3] ), 
        .ZN(n1035) );
  INV_X1 U382 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U383 ( .A1(data_in[4]), .A2(n835), .B1(n1038), .B2(\mem[18][4] ), 
        .ZN(n1034) );
  INV_X1 U384 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U385 ( .A1(data_in[5]), .A2(n835), .B1(n1038), .B2(\mem[18][5] ), 
        .ZN(n1033) );
  INV_X1 U386 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U387 ( .A1(data_in[6]), .A2(n835), .B1(n1038), .B2(\mem[18][6] ), 
        .ZN(n1032) );
  INV_X1 U388 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U389 ( .A1(data_in[7]), .A2(n835), .B1(n1038), .B2(\mem[18][7] ), 
        .ZN(n1031) );
  INV_X1 U390 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U391 ( .A1(data_in[0]), .A2(n834), .B1(n1029), .B2(\mem[19][0] ), 
        .ZN(n1030) );
  INV_X1 U392 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U393 ( .A1(data_in[1]), .A2(n834), .B1(n1029), .B2(\mem[19][1] ), 
        .ZN(n1028) );
  INV_X1 U394 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U395 ( .A1(data_in[2]), .A2(n834), .B1(n1029), .B2(\mem[19][2] ), 
        .ZN(n1027) );
  INV_X1 U396 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U397 ( .A1(data_in[3]), .A2(n834), .B1(n1029), .B2(\mem[19][3] ), 
        .ZN(n1026) );
  INV_X1 U398 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U399 ( .A1(data_in[4]), .A2(n834), .B1(n1029), .B2(\mem[19][4] ), 
        .ZN(n1025) );
  INV_X1 U400 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U401 ( .A1(data_in[5]), .A2(n834), .B1(n1029), .B2(\mem[19][5] ), 
        .ZN(n1024) );
  INV_X1 U402 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U403 ( .A1(data_in[6]), .A2(n834), .B1(n1029), .B2(\mem[19][6] ), 
        .ZN(n1023) );
  INV_X1 U404 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U405 ( .A1(data_in[7]), .A2(n834), .B1(n1029), .B2(\mem[19][7] ), 
        .ZN(n1022) );
  INV_X1 U406 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U407 ( .A1(data_in[0]), .A2(n833), .B1(n1020), .B2(\mem[20][0] ), 
        .ZN(n1021) );
  INV_X1 U408 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U409 ( .A1(data_in[1]), .A2(n833), .B1(n1020), .B2(\mem[20][1] ), 
        .ZN(n1019) );
  INV_X1 U410 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U411 ( .A1(data_in[2]), .A2(n833), .B1(n1020), .B2(\mem[20][2] ), 
        .ZN(n1018) );
  INV_X1 U412 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U413 ( .A1(data_in[3]), .A2(n833), .B1(n1020), .B2(\mem[20][3] ), 
        .ZN(n1017) );
  INV_X1 U414 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U415 ( .A1(data_in[4]), .A2(n833), .B1(n1020), .B2(\mem[20][4] ), 
        .ZN(n1016) );
  INV_X1 U416 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U417 ( .A1(data_in[5]), .A2(n833), .B1(n1020), .B2(\mem[20][5] ), 
        .ZN(n1015) );
  INV_X1 U418 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U419 ( .A1(data_in[6]), .A2(n833), .B1(n1020), .B2(\mem[20][6] ), 
        .ZN(n1014) );
  INV_X1 U420 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U421 ( .A1(data_in[7]), .A2(n833), .B1(n1020), .B2(\mem[20][7] ), 
        .ZN(n1013) );
  INV_X1 U422 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U423 ( .A1(data_in[0]), .A2(n832), .B1(n1011), .B2(\mem[21][0] ), 
        .ZN(n1012) );
  INV_X1 U424 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U425 ( .A1(data_in[1]), .A2(n832), .B1(n1011), .B2(\mem[21][1] ), 
        .ZN(n1010) );
  INV_X1 U426 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U427 ( .A1(data_in[2]), .A2(n832), .B1(n1011), .B2(\mem[21][2] ), 
        .ZN(n1009) );
  INV_X1 U428 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U429 ( .A1(data_in[3]), .A2(n832), .B1(n1011), .B2(\mem[21][3] ), 
        .ZN(n1008) );
  INV_X1 U430 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U431 ( .A1(data_in[4]), .A2(n832), .B1(n1011), .B2(\mem[21][4] ), 
        .ZN(n1007) );
  INV_X1 U432 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U433 ( .A1(data_in[5]), .A2(n832), .B1(n1011), .B2(\mem[21][5] ), 
        .ZN(n1006) );
  INV_X1 U434 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U435 ( .A1(data_in[6]), .A2(n832), .B1(n1011), .B2(\mem[21][6] ), 
        .ZN(n1005) );
  INV_X1 U436 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U437 ( .A1(data_in[7]), .A2(n832), .B1(n1011), .B2(\mem[21][7] ), 
        .ZN(n1004) );
  INV_X1 U438 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U439 ( .A1(data_in[0]), .A2(n831), .B1(n1002), .B2(\mem[22][0] ), 
        .ZN(n1003) );
  INV_X1 U440 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U441 ( .A1(data_in[1]), .A2(n831), .B1(n1002), .B2(\mem[22][1] ), 
        .ZN(n1001) );
  INV_X1 U442 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U443 ( .A1(data_in[2]), .A2(n831), .B1(n1002), .B2(\mem[22][2] ), 
        .ZN(n1000) );
  INV_X1 U444 ( .A(n999), .ZN(n706) );
  AOI22_X1 U445 ( .A1(data_in[3]), .A2(n831), .B1(n1002), .B2(\mem[22][3] ), 
        .ZN(n999) );
  INV_X1 U446 ( .A(n998), .ZN(n705) );
  AOI22_X1 U447 ( .A1(data_in[4]), .A2(n831), .B1(n1002), .B2(\mem[22][4] ), 
        .ZN(n998) );
  INV_X1 U448 ( .A(n997), .ZN(n704) );
  AOI22_X1 U449 ( .A1(data_in[5]), .A2(n831), .B1(n1002), .B2(\mem[22][5] ), 
        .ZN(n997) );
  INV_X1 U450 ( .A(n996), .ZN(n703) );
  AOI22_X1 U451 ( .A1(data_in[6]), .A2(n831), .B1(n1002), .B2(\mem[22][6] ), 
        .ZN(n996) );
  INV_X1 U452 ( .A(n995), .ZN(n702) );
  AOI22_X1 U453 ( .A1(data_in[7]), .A2(n831), .B1(n1002), .B2(\mem[22][7] ), 
        .ZN(n995) );
  INV_X1 U454 ( .A(n994), .ZN(n701) );
  AOI22_X1 U455 ( .A1(data_in[0]), .A2(n830), .B1(n993), .B2(\mem[23][0] ), 
        .ZN(n994) );
  INV_X1 U456 ( .A(n992), .ZN(n700) );
  AOI22_X1 U457 ( .A1(data_in[1]), .A2(n830), .B1(n993), .B2(\mem[23][1] ), 
        .ZN(n992) );
  INV_X1 U458 ( .A(n991), .ZN(n699) );
  AOI22_X1 U459 ( .A1(data_in[2]), .A2(n830), .B1(n993), .B2(\mem[23][2] ), 
        .ZN(n991) );
  INV_X1 U460 ( .A(n990), .ZN(n698) );
  AOI22_X1 U461 ( .A1(data_in[3]), .A2(n830), .B1(n993), .B2(\mem[23][3] ), 
        .ZN(n990) );
  INV_X1 U462 ( .A(n989), .ZN(n697) );
  AOI22_X1 U463 ( .A1(data_in[4]), .A2(n830), .B1(n993), .B2(\mem[23][4] ), 
        .ZN(n989) );
  INV_X1 U464 ( .A(n988), .ZN(n696) );
  AOI22_X1 U465 ( .A1(data_in[5]), .A2(n830), .B1(n993), .B2(\mem[23][5] ), 
        .ZN(n988) );
  INV_X1 U466 ( .A(n987), .ZN(n695) );
  AOI22_X1 U467 ( .A1(data_in[6]), .A2(n830), .B1(n993), .B2(\mem[23][6] ), 
        .ZN(n987) );
  INV_X1 U468 ( .A(n986), .ZN(n694) );
  AOI22_X1 U469 ( .A1(data_in[7]), .A2(n830), .B1(n993), .B2(\mem[23][7] ), 
        .ZN(n986) );
  INV_X1 U470 ( .A(n985), .ZN(n693) );
  AOI22_X1 U471 ( .A1(data_in[0]), .A2(n829), .B1(n984), .B2(\mem[24][0] ), 
        .ZN(n985) );
  INV_X1 U472 ( .A(n983), .ZN(n692) );
  AOI22_X1 U473 ( .A1(data_in[1]), .A2(n829), .B1(n984), .B2(\mem[24][1] ), 
        .ZN(n983) );
  INV_X1 U474 ( .A(n982), .ZN(n691) );
  AOI22_X1 U475 ( .A1(data_in[2]), .A2(n829), .B1(n984), .B2(\mem[24][2] ), 
        .ZN(n982) );
  INV_X1 U476 ( .A(n981), .ZN(n690) );
  AOI22_X1 U477 ( .A1(data_in[3]), .A2(n829), .B1(n984), .B2(\mem[24][3] ), 
        .ZN(n981) );
  INV_X1 U478 ( .A(n980), .ZN(n689) );
  AOI22_X1 U479 ( .A1(data_in[4]), .A2(n829), .B1(n984), .B2(\mem[24][4] ), 
        .ZN(n980) );
  INV_X1 U480 ( .A(n979), .ZN(n688) );
  AOI22_X1 U481 ( .A1(data_in[5]), .A2(n829), .B1(n984), .B2(\mem[24][5] ), 
        .ZN(n979) );
  INV_X1 U482 ( .A(n978), .ZN(n687) );
  AOI22_X1 U483 ( .A1(data_in[6]), .A2(n829), .B1(n984), .B2(\mem[24][6] ), 
        .ZN(n978) );
  INV_X1 U484 ( .A(n977), .ZN(n686) );
  AOI22_X1 U485 ( .A1(data_in[7]), .A2(n829), .B1(n984), .B2(\mem[24][7] ), 
        .ZN(n977) );
  INV_X1 U486 ( .A(n975), .ZN(n685) );
  AOI22_X1 U487 ( .A1(data_in[0]), .A2(n828), .B1(n974), .B2(\mem[25][0] ), 
        .ZN(n975) );
  INV_X1 U488 ( .A(n973), .ZN(n684) );
  AOI22_X1 U489 ( .A1(data_in[1]), .A2(n828), .B1(n974), .B2(\mem[25][1] ), 
        .ZN(n973) );
  INV_X1 U490 ( .A(n972), .ZN(n683) );
  AOI22_X1 U491 ( .A1(data_in[2]), .A2(n828), .B1(n974), .B2(\mem[25][2] ), 
        .ZN(n972) );
  INV_X1 U492 ( .A(n971), .ZN(n682) );
  AOI22_X1 U493 ( .A1(data_in[3]), .A2(n828), .B1(n974), .B2(\mem[25][3] ), 
        .ZN(n971) );
  INV_X1 U494 ( .A(n970), .ZN(n681) );
  AOI22_X1 U495 ( .A1(data_in[4]), .A2(n828), .B1(n974), .B2(\mem[25][4] ), 
        .ZN(n970) );
  INV_X1 U496 ( .A(n969), .ZN(n680) );
  AOI22_X1 U497 ( .A1(data_in[5]), .A2(n828), .B1(n974), .B2(\mem[25][5] ), 
        .ZN(n969) );
  INV_X1 U498 ( .A(n968), .ZN(n679) );
  AOI22_X1 U499 ( .A1(data_in[6]), .A2(n828), .B1(n974), .B2(\mem[25][6] ), 
        .ZN(n968) );
  INV_X1 U500 ( .A(n967), .ZN(n678) );
  AOI22_X1 U501 ( .A1(data_in[7]), .A2(n828), .B1(n974), .B2(\mem[25][7] ), 
        .ZN(n967) );
  INV_X1 U502 ( .A(n966), .ZN(n677) );
  AOI22_X1 U503 ( .A1(data_in[0]), .A2(n827), .B1(n965), .B2(\mem[26][0] ), 
        .ZN(n966) );
  INV_X1 U504 ( .A(n964), .ZN(n676) );
  AOI22_X1 U505 ( .A1(data_in[1]), .A2(n827), .B1(n965), .B2(\mem[26][1] ), 
        .ZN(n964) );
  INV_X1 U506 ( .A(n963), .ZN(n675) );
  AOI22_X1 U507 ( .A1(data_in[2]), .A2(n827), .B1(n965), .B2(\mem[26][2] ), 
        .ZN(n963) );
  INV_X1 U508 ( .A(n962), .ZN(n674) );
  AOI22_X1 U509 ( .A1(data_in[3]), .A2(n827), .B1(n965), .B2(\mem[26][3] ), 
        .ZN(n962) );
  INV_X1 U510 ( .A(n961), .ZN(n673) );
  AOI22_X1 U511 ( .A1(data_in[4]), .A2(n827), .B1(n965), .B2(\mem[26][4] ), 
        .ZN(n961) );
  INV_X1 U512 ( .A(n960), .ZN(n672) );
  AOI22_X1 U513 ( .A1(data_in[5]), .A2(n827), .B1(n965), .B2(\mem[26][5] ), 
        .ZN(n960) );
  INV_X1 U514 ( .A(n959), .ZN(n671) );
  AOI22_X1 U515 ( .A1(data_in[6]), .A2(n827), .B1(n965), .B2(\mem[26][6] ), 
        .ZN(n959) );
  INV_X1 U516 ( .A(n958), .ZN(n670) );
  AOI22_X1 U517 ( .A1(data_in[7]), .A2(n827), .B1(n965), .B2(\mem[26][7] ), 
        .ZN(n958) );
  INV_X1 U518 ( .A(n957), .ZN(n669) );
  AOI22_X1 U519 ( .A1(data_in[0]), .A2(n826), .B1(n956), .B2(\mem[27][0] ), 
        .ZN(n957) );
  INV_X1 U520 ( .A(n955), .ZN(n668) );
  AOI22_X1 U521 ( .A1(data_in[1]), .A2(n826), .B1(n956), .B2(\mem[27][1] ), 
        .ZN(n955) );
  INV_X1 U522 ( .A(n954), .ZN(n667) );
  AOI22_X1 U523 ( .A1(data_in[2]), .A2(n826), .B1(n956), .B2(\mem[27][2] ), 
        .ZN(n954) );
  INV_X1 U524 ( .A(n953), .ZN(n666) );
  AOI22_X1 U525 ( .A1(data_in[3]), .A2(n826), .B1(n956), .B2(\mem[27][3] ), 
        .ZN(n953) );
  INV_X1 U526 ( .A(n952), .ZN(n665) );
  AOI22_X1 U527 ( .A1(data_in[4]), .A2(n826), .B1(n956), .B2(\mem[27][4] ), 
        .ZN(n952) );
  INV_X1 U528 ( .A(n951), .ZN(n664) );
  AOI22_X1 U529 ( .A1(data_in[5]), .A2(n826), .B1(n956), .B2(\mem[27][5] ), 
        .ZN(n951) );
  INV_X1 U530 ( .A(n950), .ZN(n663) );
  AOI22_X1 U531 ( .A1(data_in[6]), .A2(n826), .B1(n956), .B2(\mem[27][6] ), 
        .ZN(n950) );
  INV_X1 U532 ( .A(n949), .ZN(n662) );
  AOI22_X1 U533 ( .A1(data_in[7]), .A2(n826), .B1(n956), .B2(\mem[27][7] ), 
        .ZN(n949) );
  INV_X1 U534 ( .A(n948), .ZN(n661) );
  AOI22_X1 U535 ( .A1(data_in[0]), .A2(n825), .B1(n947), .B2(\mem[28][0] ), 
        .ZN(n948) );
  INV_X1 U536 ( .A(n946), .ZN(n660) );
  AOI22_X1 U537 ( .A1(data_in[1]), .A2(n825), .B1(n947), .B2(\mem[28][1] ), 
        .ZN(n946) );
  INV_X1 U538 ( .A(n945), .ZN(n659) );
  AOI22_X1 U539 ( .A1(data_in[2]), .A2(n825), .B1(n947), .B2(\mem[28][2] ), 
        .ZN(n945) );
  INV_X1 U540 ( .A(n944), .ZN(n658) );
  AOI22_X1 U541 ( .A1(data_in[3]), .A2(n825), .B1(n947), .B2(\mem[28][3] ), 
        .ZN(n944) );
  INV_X1 U542 ( .A(n943), .ZN(n657) );
  AOI22_X1 U543 ( .A1(data_in[4]), .A2(n825), .B1(n947), .B2(\mem[28][4] ), 
        .ZN(n943) );
  INV_X1 U544 ( .A(n942), .ZN(n656) );
  AOI22_X1 U545 ( .A1(data_in[5]), .A2(n825), .B1(n947), .B2(\mem[28][5] ), 
        .ZN(n942) );
  INV_X1 U546 ( .A(n941), .ZN(n655) );
  AOI22_X1 U547 ( .A1(data_in[6]), .A2(n825), .B1(n947), .B2(\mem[28][6] ), 
        .ZN(n941) );
  INV_X1 U548 ( .A(n940), .ZN(n654) );
  AOI22_X1 U549 ( .A1(data_in[7]), .A2(n825), .B1(n947), .B2(\mem[28][7] ), 
        .ZN(n940) );
  INV_X1 U550 ( .A(n939), .ZN(n653) );
  AOI22_X1 U551 ( .A1(data_in[0]), .A2(n824), .B1(n938), .B2(\mem[29][0] ), 
        .ZN(n939) );
  INV_X1 U552 ( .A(n937), .ZN(n652) );
  AOI22_X1 U553 ( .A1(data_in[1]), .A2(n824), .B1(n938), .B2(\mem[29][1] ), 
        .ZN(n937) );
  INV_X1 U554 ( .A(n936), .ZN(n651) );
  AOI22_X1 U555 ( .A1(data_in[2]), .A2(n824), .B1(n938), .B2(\mem[29][2] ), 
        .ZN(n936) );
  INV_X1 U556 ( .A(n935), .ZN(n650) );
  AOI22_X1 U557 ( .A1(data_in[3]), .A2(n824), .B1(n938), .B2(\mem[29][3] ), 
        .ZN(n935) );
  INV_X1 U558 ( .A(n934), .ZN(n649) );
  AOI22_X1 U559 ( .A1(data_in[4]), .A2(n824), .B1(n938), .B2(\mem[29][4] ), 
        .ZN(n934) );
  INV_X1 U560 ( .A(n933), .ZN(n648) );
  AOI22_X1 U561 ( .A1(data_in[5]), .A2(n824), .B1(n938), .B2(\mem[29][5] ), 
        .ZN(n933) );
  INV_X1 U562 ( .A(n932), .ZN(n647) );
  AOI22_X1 U563 ( .A1(data_in[6]), .A2(n824), .B1(n938), .B2(\mem[29][6] ), 
        .ZN(n932) );
  INV_X1 U564 ( .A(n931), .ZN(n646) );
  AOI22_X1 U565 ( .A1(data_in[7]), .A2(n824), .B1(n938), .B2(\mem[29][7] ), 
        .ZN(n931) );
  INV_X1 U566 ( .A(n930), .ZN(n645) );
  AOI22_X1 U567 ( .A1(data_in[0]), .A2(n823), .B1(n929), .B2(\mem[30][0] ), 
        .ZN(n930) );
  INV_X1 U568 ( .A(n928), .ZN(n644) );
  AOI22_X1 U569 ( .A1(data_in[1]), .A2(n823), .B1(n929), .B2(\mem[30][1] ), 
        .ZN(n928) );
  INV_X1 U570 ( .A(n927), .ZN(n643) );
  AOI22_X1 U571 ( .A1(data_in[2]), .A2(n823), .B1(n929), .B2(\mem[30][2] ), 
        .ZN(n927) );
  INV_X1 U572 ( .A(n926), .ZN(n642) );
  AOI22_X1 U573 ( .A1(data_in[3]), .A2(n823), .B1(n929), .B2(\mem[30][3] ), 
        .ZN(n926) );
  INV_X1 U574 ( .A(n925), .ZN(n641) );
  AOI22_X1 U575 ( .A1(data_in[4]), .A2(n823), .B1(n929), .B2(\mem[30][4] ), 
        .ZN(n925) );
  INV_X1 U576 ( .A(n924), .ZN(n640) );
  AOI22_X1 U577 ( .A1(data_in[5]), .A2(n823), .B1(n929), .B2(\mem[30][5] ), 
        .ZN(n924) );
  INV_X1 U578 ( .A(n923), .ZN(n639) );
  AOI22_X1 U579 ( .A1(data_in[6]), .A2(n823), .B1(n929), .B2(\mem[30][6] ), 
        .ZN(n923) );
  INV_X1 U580 ( .A(n922), .ZN(n638) );
  AOI22_X1 U581 ( .A1(data_in[7]), .A2(n823), .B1(n929), .B2(\mem[30][7] ), 
        .ZN(n922) );
  INV_X1 U582 ( .A(n921), .ZN(n637) );
  AOI22_X1 U583 ( .A1(data_in[0]), .A2(n822), .B1(n920), .B2(\mem[31][0] ), 
        .ZN(n921) );
  INV_X1 U584 ( .A(n919), .ZN(n636) );
  AOI22_X1 U585 ( .A1(data_in[1]), .A2(n822), .B1(n920), .B2(\mem[31][1] ), 
        .ZN(n919) );
  INV_X1 U586 ( .A(n918), .ZN(n635) );
  AOI22_X1 U587 ( .A1(data_in[2]), .A2(n822), .B1(n920), .B2(\mem[31][2] ), 
        .ZN(n918) );
  INV_X1 U588 ( .A(n917), .ZN(n634) );
  AOI22_X1 U589 ( .A1(data_in[3]), .A2(n822), .B1(n920), .B2(\mem[31][3] ), 
        .ZN(n917) );
  INV_X1 U590 ( .A(n916), .ZN(n633) );
  AOI22_X1 U591 ( .A1(data_in[4]), .A2(n822), .B1(n920), .B2(\mem[31][4] ), 
        .ZN(n916) );
  INV_X1 U592 ( .A(n915), .ZN(n632) );
  AOI22_X1 U593 ( .A1(data_in[5]), .A2(n822), .B1(n920), .B2(\mem[31][5] ), 
        .ZN(n915) );
  INV_X1 U594 ( .A(n914), .ZN(n631) );
  AOI22_X1 U595 ( .A1(data_in[6]), .A2(n822), .B1(n920), .B2(\mem[31][6] ), 
        .ZN(n914) );
  INV_X1 U596 ( .A(n913), .ZN(n630) );
  AOI22_X1 U597 ( .A1(data_in[7]), .A2(n822), .B1(n920), .B2(\mem[31][7] ), 
        .ZN(n913) );
  MUX2_X1 U598 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n618), .Z(n4) );
  MUX2_X1 U599 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n618), .Z(n5) );
  MUX2_X1 U600 ( .A(n5), .B(n4), .S(n611), .Z(n6) );
  MUX2_X1 U601 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n617), .Z(n7) );
  MUX2_X1 U602 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n616), .Z(n8) );
  MUX2_X1 U603 ( .A(n8), .B(n7), .S(n611), .Z(n9) );
  MUX2_X1 U604 ( .A(n9), .B(n6), .S(n609), .Z(n10) );
  MUX2_X1 U605 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n617), .Z(n11) );
  MUX2_X1 U606 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n618), .Z(n12) );
  MUX2_X1 U607 ( .A(n12), .B(n11), .S(n611), .Z(n13) );
  MUX2_X1 U608 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n615), .Z(n14) );
  MUX2_X1 U609 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n615), .Z(n15) );
  MUX2_X1 U610 ( .A(n15), .B(n14), .S(n611), .Z(n16) );
  MUX2_X1 U611 ( .A(n16), .B(n13), .S(N12), .Z(n17) );
  MUX2_X1 U612 ( .A(n17), .B(n10), .S(N13), .Z(n18) );
  MUX2_X1 U613 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n614), .Z(n19) );
  MUX2_X1 U614 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n614), .Z(n20) );
  MUX2_X1 U615 ( .A(n20), .B(n19), .S(n613), .Z(n21) );
  MUX2_X1 U616 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n614), .Z(n22) );
  MUX2_X1 U617 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n614), .Z(n23) );
  MUX2_X1 U618 ( .A(n23), .B(n22), .S(N11), .Z(n24) );
  MUX2_X1 U619 ( .A(n24), .B(n21), .S(N12), .Z(n25) );
  MUX2_X1 U620 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n614), .Z(n26) );
  MUX2_X1 U621 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n614), .Z(n27) );
  MUX2_X1 U622 ( .A(n27), .B(n26), .S(n613), .Z(n28) );
  MUX2_X1 U623 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n614), .Z(n29) );
  MUX2_X1 U624 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n614), .Z(n30) );
  MUX2_X1 U625 ( .A(n30), .B(n29), .S(n613), .Z(n31) );
  MUX2_X1 U626 ( .A(n31), .B(n28), .S(n610), .Z(n32) );
  MUX2_X1 U627 ( .A(n32), .B(n25), .S(N13), .Z(n33) );
  MUX2_X1 U628 ( .A(n33), .B(n18), .S(N14), .Z(N22) );
  MUX2_X1 U629 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n614), .Z(n34) );
  MUX2_X1 U630 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n614), .Z(n35) );
  MUX2_X1 U631 ( .A(n35), .B(n34), .S(n612), .Z(n36) );
  MUX2_X1 U632 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n614), .Z(n37) );
  MUX2_X1 U633 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n614), .Z(n38) );
  MUX2_X1 U634 ( .A(n38), .B(n37), .S(n613), .Z(n39) );
  MUX2_X1 U635 ( .A(n39), .B(n36), .S(n610), .Z(n40) );
  MUX2_X1 U636 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n615), .Z(n41) );
  MUX2_X1 U637 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n619), .Z(n42) );
  MUX2_X1 U638 ( .A(n42), .B(n41), .S(n611), .Z(n43) );
  MUX2_X1 U639 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n619), .Z(n44) );
  MUX2_X1 U640 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(N10), .Z(n45) );
  MUX2_X1 U641 ( .A(n45), .B(n44), .S(N11), .Z(n46) );
  MUX2_X1 U642 ( .A(n46), .B(n43), .S(n609), .Z(n47) );
  MUX2_X1 U643 ( .A(n47), .B(n40), .S(N13), .Z(n48) );
  MUX2_X1 U644 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n616), .Z(n49) );
  MUX2_X1 U645 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n617), .Z(n50) );
  MUX2_X1 U646 ( .A(n50), .B(n49), .S(n611), .Z(n51) );
  MUX2_X1 U647 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n619), .Z(n52) );
  MUX2_X1 U648 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(N10), .Z(n53) );
  MUX2_X1 U649 ( .A(n53), .B(n52), .S(N11), .Z(n54) );
  MUX2_X1 U650 ( .A(n54), .B(n51), .S(N12), .Z(n55) );
  MUX2_X1 U651 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n619), .Z(n56) );
  MUX2_X1 U652 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n57) );
  MUX2_X1 U653 ( .A(n57), .B(n56), .S(n612), .Z(n58) );
  MUX2_X1 U654 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(N10), .Z(n59) );
  MUX2_X1 U655 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(N10), .Z(n60) );
  MUX2_X1 U656 ( .A(n60), .B(n59), .S(n612), .Z(n61) );
  MUX2_X1 U657 ( .A(n61), .B(n58), .S(n609), .Z(n62) );
  MUX2_X1 U658 ( .A(n62), .B(n55), .S(N13), .Z(n63) );
  MUX2_X1 U659 ( .A(n63), .B(n48), .S(N14), .Z(N21) );
  MUX2_X1 U660 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n615), .Z(n64) );
  MUX2_X1 U661 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n615), .Z(n65) );
  MUX2_X1 U662 ( .A(n65), .B(n64), .S(n611), .Z(n66) );
  MUX2_X1 U663 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n615), .Z(n67) );
  MUX2_X1 U664 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n615), .Z(n68) );
  MUX2_X1 U665 ( .A(n68), .B(n67), .S(n611), .Z(n69) );
  MUX2_X1 U666 ( .A(n69), .B(n66), .S(n609), .Z(n70) );
  MUX2_X1 U667 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n615), .Z(n71) );
  MUX2_X1 U668 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n615), .Z(n72) );
  MUX2_X1 U669 ( .A(n72), .B(n71), .S(n611), .Z(n73) );
  MUX2_X1 U670 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n615), .Z(n74) );
  MUX2_X1 U671 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n615), .Z(n75) );
  MUX2_X1 U672 ( .A(n75), .B(n74), .S(n611), .Z(n76) );
  MUX2_X1 U673 ( .A(n76), .B(n73), .S(n609), .Z(n77) );
  MUX2_X1 U674 ( .A(n77), .B(n70), .S(N13), .Z(n78) );
  MUX2_X1 U675 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n615), .Z(n79) );
  MUX2_X1 U676 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n615), .Z(n80) );
  MUX2_X1 U677 ( .A(n80), .B(n79), .S(n611), .Z(n81) );
  MUX2_X1 U678 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n615), .Z(n82) );
  MUX2_X1 U679 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n615), .Z(n83) );
  MUX2_X1 U680 ( .A(n83), .B(n82), .S(n613), .Z(n84) );
  MUX2_X1 U681 ( .A(n84), .B(n81), .S(n609), .Z(n85) );
  MUX2_X1 U682 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n616), .Z(n86) );
  MUX2_X1 U683 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n616), .Z(n87) );
  MUX2_X1 U684 ( .A(n87), .B(n86), .S(n612), .Z(n88) );
  MUX2_X1 U685 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n616), .Z(n89) );
  MUX2_X1 U686 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n616), .Z(n90) );
  MUX2_X1 U687 ( .A(n90), .B(n89), .S(n611), .Z(n91) );
  MUX2_X1 U688 ( .A(n91), .B(n88), .S(n609), .Z(n92) );
  MUX2_X1 U689 ( .A(n92), .B(n85), .S(N13), .Z(n93) );
  MUX2_X1 U690 ( .A(n93), .B(n78), .S(N14), .Z(N20) );
  MUX2_X1 U691 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n616), .Z(n94) );
  MUX2_X1 U692 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n616), .Z(n95) );
  MUX2_X1 U693 ( .A(n95), .B(n94), .S(n611), .Z(n96) );
  MUX2_X1 U694 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n616), .Z(n97) );
  MUX2_X1 U695 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n616), .Z(n98) );
  MUX2_X1 U696 ( .A(n98), .B(n97), .S(n611), .Z(n99) );
  MUX2_X1 U697 ( .A(n99), .B(n96), .S(n609), .Z(n100) );
  MUX2_X1 U698 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n616), .Z(n101) );
  MUX2_X1 U699 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n616), .Z(n102) );
  MUX2_X1 U700 ( .A(n102), .B(n101), .S(n611), .Z(n103) );
  MUX2_X1 U701 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n616), .Z(n104) );
  MUX2_X1 U702 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n616), .Z(n105) );
  MUX2_X1 U703 ( .A(n105), .B(n104), .S(N11), .Z(n106) );
  MUX2_X1 U704 ( .A(n106), .B(n103), .S(n609), .Z(n107) );
  MUX2_X1 U705 ( .A(n107), .B(n100), .S(N13), .Z(n108) );
  MUX2_X1 U706 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n619), .Z(n109) );
  MUX2_X1 U707 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n619), .Z(n110) );
  MUX2_X1 U708 ( .A(n110), .B(n109), .S(n612), .Z(n111) );
  MUX2_X1 U709 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n619), .Z(n112) );
  MUX2_X1 U710 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n618), .Z(n113) );
  MUX2_X1 U711 ( .A(n113), .B(n112), .S(n612), .Z(n114) );
  MUX2_X1 U712 ( .A(n114), .B(n111), .S(n609), .Z(n115) );
  MUX2_X1 U713 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n619), .Z(n116) );
  MUX2_X1 U714 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n615), .Z(n117) );
  MUX2_X1 U715 ( .A(n117), .B(n116), .S(n612), .Z(n118) );
  MUX2_X1 U716 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n617), .Z(n119) );
  MUX2_X1 U717 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n616), .Z(n120) );
  MUX2_X1 U718 ( .A(n120), .B(n119), .S(n612), .Z(n121) );
  MUX2_X1 U719 ( .A(n121), .B(n118), .S(n609), .Z(n122) );
  MUX2_X1 U720 ( .A(n122), .B(n115), .S(N13), .Z(n123) );
  MUX2_X1 U721 ( .A(n123), .B(n108), .S(N14), .Z(N19) );
  MUX2_X1 U722 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n616), .Z(n124) );
  MUX2_X1 U723 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n619), .Z(n125) );
  MUX2_X1 U724 ( .A(n125), .B(n124), .S(n612), .Z(n126) );
  MUX2_X1 U725 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n619), .Z(n127) );
  MUX2_X1 U726 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n619), .Z(n128) );
  MUX2_X1 U727 ( .A(n128), .B(n127), .S(n612), .Z(n129) );
  MUX2_X1 U728 ( .A(n129), .B(n126), .S(n609), .Z(n130) );
  MUX2_X1 U729 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n617), .Z(n131) );
  MUX2_X1 U730 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n619), .Z(n132) );
  MUX2_X1 U731 ( .A(n132), .B(n131), .S(n612), .Z(n133) );
  MUX2_X1 U732 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n616), .Z(n134) );
  MUX2_X1 U733 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n619), .Z(n135) );
  MUX2_X1 U734 ( .A(n135), .B(n134), .S(n612), .Z(n136) );
  MUX2_X1 U735 ( .A(n136), .B(n133), .S(n609), .Z(n137) );
  MUX2_X1 U736 ( .A(n137), .B(n130), .S(N13), .Z(n138) );
  MUX2_X1 U737 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n619), .Z(n139) );
  MUX2_X1 U738 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n617), .Z(n140) );
  MUX2_X1 U739 ( .A(n140), .B(n139), .S(n612), .Z(n141) );
  MUX2_X1 U740 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n618), .Z(n142) );
  MUX2_X1 U741 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n619), .Z(n143) );
  MUX2_X1 U742 ( .A(n143), .B(n142), .S(n612), .Z(n144) );
  MUX2_X1 U743 ( .A(n144), .B(n141), .S(n609), .Z(n145) );
  MUX2_X1 U744 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n615), .Z(n146) );
  MUX2_X1 U745 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n619), .Z(n147) );
  MUX2_X1 U746 ( .A(n147), .B(n146), .S(n612), .Z(n148) );
  MUX2_X1 U747 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n619), .Z(n149) );
  MUX2_X1 U748 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n619), .Z(n150) );
  MUX2_X1 U749 ( .A(n150), .B(n149), .S(n612), .Z(n151) );
  MUX2_X1 U750 ( .A(n151), .B(n148), .S(n609), .Z(n152) );
  MUX2_X1 U751 ( .A(n152), .B(n145), .S(N13), .Z(n153) );
  MUX2_X1 U752 ( .A(n153), .B(n138), .S(N14), .Z(N18) );
  MUX2_X1 U753 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n614), .Z(n154) );
  MUX2_X1 U754 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n614), .Z(n155) );
  MUX2_X1 U755 ( .A(n155), .B(n154), .S(n613), .Z(n156) );
  MUX2_X1 U756 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n614), .Z(n157) );
  MUX2_X1 U757 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n614), .Z(n158) );
  MUX2_X1 U758 ( .A(n158), .B(n157), .S(n613), .Z(n159) );
  MUX2_X1 U759 ( .A(n159), .B(n156), .S(n610), .Z(n160) );
  MUX2_X1 U760 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n614), .Z(n161) );
  MUX2_X1 U761 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n614), .Z(n162) );
  MUX2_X1 U762 ( .A(n162), .B(n161), .S(n613), .Z(n163) );
  MUX2_X1 U763 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n614), .Z(n164) );
  MUX2_X1 U764 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n619), .Z(n165) );
  MUX2_X1 U765 ( .A(n165), .B(n164), .S(n613), .Z(n166) );
  MUX2_X1 U766 ( .A(n166), .B(n163), .S(n610), .Z(n167) );
  MUX2_X1 U767 ( .A(n167), .B(n160), .S(N13), .Z(n168) );
  MUX2_X1 U768 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n614), .Z(n169) );
  MUX2_X1 U769 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n614), .Z(n170) );
  MUX2_X1 U770 ( .A(n170), .B(n169), .S(n613), .Z(n171) );
  MUX2_X1 U771 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n614), .Z(n172) );
  MUX2_X1 U772 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n614), .Z(n173) );
  MUX2_X1 U773 ( .A(n173), .B(n172), .S(n613), .Z(n174) );
  MUX2_X1 U774 ( .A(n174), .B(n171), .S(n610), .Z(n175) );
  MUX2_X1 U775 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n617), .Z(n176) );
  MUX2_X1 U776 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n617), .Z(n177) );
  MUX2_X1 U777 ( .A(n177), .B(n176), .S(n613), .Z(n178) );
  MUX2_X1 U778 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n617), .Z(n179) );
  MUX2_X1 U779 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n617), .Z(n180) );
  MUX2_X1 U780 ( .A(n180), .B(n179), .S(n613), .Z(n181) );
  MUX2_X1 U781 ( .A(n181), .B(n178), .S(n610), .Z(n182) );
  MUX2_X1 U782 ( .A(n182), .B(n175), .S(N13), .Z(n183) );
  MUX2_X1 U783 ( .A(n183), .B(n168), .S(N14), .Z(N17) );
  MUX2_X1 U784 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n617), .Z(n184) );
  MUX2_X1 U785 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n617), .Z(n185) );
  MUX2_X1 U786 ( .A(n185), .B(n184), .S(n613), .Z(n186) );
  MUX2_X1 U787 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n617), .Z(n187) );
  MUX2_X1 U788 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n617), .Z(n188) );
  MUX2_X1 U789 ( .A(n188), .B(n187), .S(n613), .Z(n189) );
  MUX2_X1 U790 ( .A(n189), .B(n186), .S(n610), .Z(n190) );
  MUX2_X1 U791 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n617), .Z(n191) );
  MUX2_X1 U792 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n617), .Z(n192) );
  MUX2_X1 U793 ( .A(n192), .B(n191), .S(n613), .Z(n193) );
  MUX2_X1 U794 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n617), .Z(n194) );
  MUX2_X1 U795 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n617), .Z(n195) );
  MUX2_X1 U796 ( .A(n195), .B(n194), .S(n613), .Z(n196) );
  MUX2_X1 U797 ( .A(n196), .B(n193), .S(n610), .Z(n197) );
  MUX2_X1 U798 ( .A(n197), .B(n190), .S(N13), .Z(n198) );
  MUX2_X1 U799 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n618), .Z(n199) );
  MUX2_X1 U800 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n618), .Z(n200) );
  MUX2_X1 U801 ( .A(n200), .B(n199), .S(n613), .Z(n201) );
  MUX2_X1 U802 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n618), .Z(n202) );
  MUX2_X1 U803 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n618), .Z(n203) );
  MUX2_X1 U804 ( .A(n203), .B(n202), .S(n613), .Z(n204) );
  MUX2_X1 U805 ( .A(n204), .B(n201), .S(n610), .Z(n205) );
  MUX2_X1 U806 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n618), .Z(n206) );
  MUX2_X1 U807 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n618), .Z(n207) );
  MUX2_X1 U808 ( .A(n207), .B(n206), .S(n612), .Z(n208) );
  MUX2_X1 U809 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n618), .Z(n209) );
  MUX2_X1 U810 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n618), .Z(n210) );
  MUX2_X1 U811 ( .A(n210), .B(n209), .S(n611), .Z(n211) );
  MUX2_X1 U812 ( .A(n211), .B(n208), .S(n610), .Z(n212) );
  MUX2_X1 U813 ( .A(n212), .B(n205), .S(N13), .Z(n213) );
  MUX2_X1 U814 ( .A(n213), .B(n198), .S(N14), .Z(N16) );
  MUX2_X1 U815 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n618), .Z(n214) );
  MUX2_X1 U816 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n618), .Z(n215) );
  MUX2_X1 U817 ( .A(n215), .B(n214), .S(n612), .Z(n216) );
  MUX2_X1 U818 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n618), .Z(n217) );
  MUX2_X1 U819 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n618), .Z(n218) );
  MUX2_X1 U820 ( .A(n218), .B(n217), .S(N11), .Z(n219) );
  MUX2_X1 U821 ( .A(n219), .B(n216), .S(n610), .Z(n220) );
  MUX2_X1 U822 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n618), .Z(n221) );
  MUX2_X1 U823 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n615), .Z(n222) );
  MUX2_X1 U824 ( .A(n222), .B(n221), .S(n611), .Z(n223) );
  MUX2_X1 U825 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n617), .Z(n224) );
  MUX2_X1 U826 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n618), .Z(n225) );
  MUX2_X1 U827 ( .A(n225), .B(n224), .S(n613), .Z(n226) );
  MUX2_X1 U828 ( .A(n226), .B(n223), .S(n610), .Z(n227) );
  MUX2_X1 U829 ( .A(n227), .B(n220), .S(N13), .Z(n228) );
  MUX2_X1 U830 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n619), .Z(n229) );
  MUX2_X1 U831 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n615), .Z(n595) );
  MUX2_X1 U832 ( .A(n595), .B(n229), .S(n612), .Z(n596) );
  MUX2_X1 U833 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n616), .Z(n597) );
  MUX2_X1 U834 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n616), .Z(n598) );
  MUX2_X1 U835 ( .A(n598), .B(n597), .S(n612), .Z(n599) );
  MUX2_X1 U836 ( .A(n599), .B(n596), .S(n610), .Z(n600) );
  MUX2_X1 U837 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n617), .Z(n601) );
  MUX2_X1 U838 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n616), .Z(n602) );
  MUX2_X1 U839 ( .A(n602), .B(n601), .S(n611), .Z(n603) );
  MUX2_X1 U840 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n618), .Z(n604) );
  MUX2_X1 U841 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n615), .Z(n605) );
  MUX2_X1 U842 ( .A(n605), .B(n604), .S(n613), .Z(n606) );
  MUX2_X1 U843 ( .A(n606), .B(n603), .S(n610), .Z(n607) );
  MUX2_X1 U844 ( .A(n607), .B(n600), .S(N13), .Z(n608) );
  MUX2_X1 U845 ( .A(n608), .B(n228), .S(N14), .Z(N15) );
  CLKBUF_X1 U846 ( .A(N11), .Z(n611) );
  INV_X1 U847 ( .A(N10), .ZN(n620) );
  INV_X1 U848 ( .A(N11), .ZN(n621) );
  INV_X1 U849 ( .A(data_in[0]), .ZN(n622) );
  INV_X1 U850 ( .A(data_in[1]), .ZN(n623) );
  INV_X1 U851 ( .A(data_in[2]), .ZN(n624) );
  INV_X1 U852 ( .A(data_in[3]), .ZN(n625) );
  INV_X1 U853 ( .A(data_in[4]), .ZN(n626) );
  INV_X1 U854 ( .A(data_in[5]), .ZN(n627) );
  INV_X1 U855 ( .A(data_in[6]), .ZN(n628) );
  INV_X1 U856 ( .A(data_in[7]), .ZN(n629) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_12 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n632), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n633), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n634), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n635), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n636), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n637), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n638), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n639), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n640), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n641), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n642), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n643), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n644), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n645), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n646), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n647), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n648), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n649), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n650), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n651), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n652), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n653), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n654), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n655), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n656), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n657), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n658), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n659), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n660), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n661), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n662), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n663), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n664), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n665), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n666), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n667), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n668), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n669), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n670), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n671), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n672), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n673), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n674), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n675), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n676), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n677), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n678), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n679), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n680), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n681), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n682), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n683), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n684), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n685), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n686), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n687), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n688), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n689), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n690), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n691), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n692), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n693), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n694), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n695), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n696), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n697), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n698), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n699), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n700), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n701), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n702), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n703), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n704), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n705), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n706), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n707), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n708), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n709), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n710), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n711), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n712), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n713), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n714), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n715), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n716), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n717), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n718), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n719), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n720), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n721), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n722), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n723), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n724), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n725), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n726), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n727), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n728), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n729), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n730), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n731), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n732), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n733), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n734), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n735), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n736), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n737), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n738), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n739), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n740), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n741), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n742), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n743), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n744), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n745), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n746), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n747), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n748), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n749), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n750), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n751), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n752), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n753), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n754), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n755), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n756), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n757), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n758), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n759), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n760), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n761), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n762), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n763), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n764), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n765), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n766), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n767), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n768), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n769), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n770), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n771), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n772), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n773), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n774), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n775), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n776), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n777), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n778), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n779), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n780), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n781), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n782), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n783), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n784), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n785), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n786), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n787), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n788), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n789), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n790), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n791), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n792), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n793), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n794), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n795), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n796), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n797), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n798), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n799), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n800), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n801), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n802), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n803), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n804), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n805), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n806), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n807), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n808), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n809), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n810), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n811), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n812), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n813), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n814), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n815), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n816), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n817), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n818), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n819), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n820), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n821), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n822), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n823), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n851), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n852), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n853), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n854), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n855), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n856), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n857), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n858), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n859), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n860), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n861), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n862), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n863), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n864), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n865), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n866), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n867), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n868), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n869), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n870), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n871), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n872), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n873), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n874), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n875), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n876), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n877), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n878), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n879), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n880), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n881), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n882), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n883), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n884), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n885), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n886), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n887), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n888), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n889), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n890), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n891), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n892), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n893), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n894), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n895), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n896), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n897), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n898), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n899), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n900), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n901), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n902), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n903), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n904), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n905), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n906), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n907), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n908), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n909), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n910), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n911), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n912), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n913), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n914), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  CLKBUF_X1 U3 ( .A(N10), .Z(n621) );
  BUF_X1 U4 ( .A(n620), .Z(n612) );
  BUF_X1 U5 ( .A(n621), .Z(n618) );
  BUF_X1 U6 ( .A(n621), .Z(n619) );
  BUF_X1 U7 ( .A(n621), .Z(n617) );
  BUF_X1 U8 ( .A(n620), .Z(n614) );
  BUF_X1 U9 ( .A(n620), .Z(n613) );
  BUF_X1 U10 ( .A(n620), .Z(n615) );
  BUF_X1 U11 ( .A(n620), .Z(n616) );
  BUF_X1 U12 ( .A(N11), .Z(n610) );
  BUF_X1 U13 ( .A(N11), .Z(n611) );
  BUF_X1 U14 ( .A(N10), .Z(n620) );
  NOR3_X1 U15 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1206) );
  NOR3_X1 U16 ( .A1(N11), .A2(N12), .A3(n622), .ZN(n1195) );
  NOR3_X1 U17 ( .A1(N10), .A2(N12), .A3(n623), .ZN(n1185) );
  NOR3_X1 U18 ( .A1(n622), .A2(N12), .A3(n623), .ZN(n1175) );
  INV_X1 U19 ( .A(n1132), .ZN(n847) );
  INV_X1 U20 ( .A(n1122), .ZN(n846) );
  INV_X1 U21 ( .A(n1113), .ZN(n845) );
  INV_X1 U22 ( .A(n1104), .ZN(n844) );
  INV_X1 U23 ( .A(n1059), .ZN(n839) );
  INV_X1 U24 ( .A(n1049), .ZN(n838) );
  INV_X1 U25 ( .A(n1040), .ZN(n837) );
  INV_X1 U26 ( .A(n1031), .ZN(n836) );
  INV_X1 U27 ( .A(n986), .ZN(n831) );
  INV_X1 U28 ( .A(n976), .ZN(n830) );
  INV_X1 U29 ( .A(n967), .ZN(n829) );
  INV_X1 U30 ( .A(n958), .ZN(n828) );
  INV_X1 U31 ( .A(n949), .ZN(n827) );
  INV_X1 U32 ( .A(n940), .ZN(n826) );
  INV_X1 U33 ( .A(n931), .ZN(n825) );
  INV_X1 U34 ( .A(n922), .ZN(n824) );
  INV_X1 U35 ( .A(n1095), .ZN(n843) );
  INV_X1 U36 ( .A(n1086), .ZN(n842) );
  INV_X1 U37 ( .A(n1077), .ZN(n841) );
  INV_X1 U38 ( .A(n1068), .ZN(n840) );
  INV_X1 U39 ( .A(n1022), .ZN(n835) );
  INV_X1 U40 ( .A(n1013), .ZN(n834) );
  INV_X1 U41 ( .A(n1004), .ZN(n833) );
  INV_X1 U42 ( .A(n995), .ZN(n832) );
  BUF_X1 U43 ( .A(N12), .Z(n607) );
  BUF_X1 U44 ( .A(N12), .Z(n608) );
  INV_X1 U45 ( .A(N13), .ZN(n849) );
  AND3_X1 U46 ( .A1(n622), .A2(n623), .A3(N12), .ZN(n1165) );
  AND3_X1 U47 ( .A1(N10), .A2(n623), .A3(N12), .ZN(n1155) );
  AND3_X1 U48 ( .A1(N11), .A2(n622), .A3(N12), .ZN(n1145) );
  AND3_X1 U49 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1135) );
  INV_X1 U50 ( .A(N14), .ZN(n850) );
  NAND2_X1 U51 ( .A1(n1195), .A2(n1205), .ZN(n1204) );
  NAND2_X1 U52 ( .A1(n1185), .A2(n1205), .ZN(n1194) );
  NAND2_X1 U53 ( .A1(n1175), .A2(n1205), .ZN(n1184) );
  NAND2_X1 U54 ( .A1(n1165), .A2(n1205), .ZN(n1174) );
  NAND2_X1 U55 ( .A1(n1155), .A2(n1205), .ZN(n1164) );
  NAND2_X1 U56 ( .A1(n1145), .A2(n1205), .ZN(n1154) );
  NAND2_X1 U57 ( .A1(n1135), .A2(n1205), .ZN(n1144) );
  NAND2_X1 U58 ( .A1(n1206), .A2(n1205), .ZN(n1215) );
  NAND2_X1 U59 ( .A1(n1124), .A2(n1206), .ZN(n1132) );
  NAND2_X1 U60 ( .A1(n1124), .A2(n1195), .ZN(n1122) );
  NAND2_X1 U61 ( .A1(n1124), .A2(n1185), .ZN(n1113) );
  NAND2_X1 U62 ( .A1(n1124), .A2(n1175), .ZN(n1104) );
  NAND2_X1 U63 ( .A1(n1051), .A2(n1206), .ZN(n1059) );
  NAND2_X1 U64 ( .A1(n1051), .A2(n1195), .ZN(n1049) );
  NAND2_X1 U65 ( .A1(n1051), .A2(n1185), .ZN(n1040) );
  NAND2_X1 U66 ( .A1(n1051), .A2(n1175), .ZN(n1031) );
  NAND2_X1 U67 ( .A1(n978), .A2(n1206), .ZN(n986) );
  NAND2_X1 U68 ( .A1(n978), .A2(n1195), .ZN(n976) );
  NAND2_X1 U69 ( .A1(n978), .A2(n1185), .ZN(n967) );
  NAND2_X1 U70 ( .A1(n978), .A2(n1175), .ZN(n958) );
  NAND2_X1 U71 ( .A1(n1124), .A2(n1165), .ZN(n1095) );
  NAND2_X1 U72 ( .A1(n1124), .A2(n1155), .ZN(n1086) );
  NAND2_X1 U73 ( .A1(n1124), .A2(n1145), .ZN(n1077) );
  NAND2_X1 U74 ( .A1(n1124), .A2(n1135), .ZN(n1068) );
  NAND2_X1 U75 ( .A1(n1051), .A2(n1165), .ZN(n1022) );
  NAND2_X1 U76 ( .A1(n1051), .A2(n1155), .ZN(n1013) );
  NAND2_X1 U77 ( .A1(n1051), .A2(n1145), .ZN(n1004) );
  NAND2_X1 U78 ( .A1(n1051), .A2(n1135), .ZN(n995) );
  NAND2_X1 U79 ( .A1(n978), .A2(n1165), .ZN(n949) );
  NAND2_X1 U80 ( .A1(n978), .A2(n1155), .ZN(n940) );
  NAND2_X1 U81 ( .A1(n978), .A2(n1145), .ZN(n931) );
  NAND2_X1 U82 ( .A1(n978), .A2(n1135), .ZN(n922) );
  AND3_X1 U83 ( .A1(n849), .A2(n850), .A3(n1134), .ZN(n1205) );
  AND3_X1 U84 ( .A1(N13), .A2(n1134), .A3(N14), .ZN(n978) );
  AND3_X1 U85 ( .A1(n1134), .A2(n850), .A3(N13), .ZN(n1124) );
  AND3_X1 U86 ( .A1(n1134), .A2(n849), .A3(N14), .ZN(n1051) );
  NOR2_X1 U87 ( .A1(n848), .A2(addr[5]), .ZN(n1134) );
  INV_X1 U88 ( .A(wr_en), .ZN(n848) );
  OAI21_X1 U89 ( .B1(n624), .B2(n1174), .A(n1173), .ZN(n882) );
  NAND2_X1 U90 ( .A1(\mem[4][0] ), .A2(n1174), .ZN(n1173) );
  OAI21_X1 U91 ( .B1(n625), .B2(n1174), .A(n1172), .ZN(n881) );
  NAND2_X1 U92 ( .A1(\mem[4][1] ), .A2(n1174), .ZN(n1172) );
  OAI21_X1 U93 ( .B1(n626), .B2(n1174), .A(n1171), .ZN(n880) );
  NAND2_X1 U94 ( .A1(\mem[4][2] ), .A2(n1174), .ZN(n1171) );
  OAI21_X1 U95 ( .B1(n627), .B2(n1174), .A(n1170), .ZN(n879) );
  NAND2_X1 U96 ( .A1(\mem[4][3] ), .A2(n1174), .ZN(n1170) );
  OAI21_X1 U97 ( .B1(n628), .B2(n1174), .A(n1169), .ZN(n878) );
  NAND2_X1 U98 ( .A1(\mem[4][4] ), .A2(n1174), .ZN(n1169) );
  OAI21_X1 U99 ( .B1(n629), .B2(n1174), .A(n1168), .ZN(n877) );
  NAND2_X1 U100 ( .A1(\mem[4][5] ), .A2(n1174), .ZN(n1168) );
  OAI21_X1 U101 ( .B1(n630), .B2(n1174), .A(n1167), .ZN(n876) );
  NAND2_X1 U102 ( .A1(\mem[4][6] ), .A2(n1174), .ZN(n1167) );
  OAI21_X1 U103 ( .B1(n631), .B2(n1174), .A(n1166), .ZN(n875) );
  NAND2_X1 U104 ( .A1(\mem[4][7] ), .A2(n1174), .ZN(n1166) );
  OAI21_X1 U105 ( .B1(n624), .B2(n1154), .A(n1153), .ZN(n866) );
  NAND2_X1 U106 ( .A1(\mem[6][0] ), .A2(n1154), .ZN(n1153) );
  OAI21_X1 U107 ( .B1(n625), .B2(n1154), .A(n1152), .ZN(n865) );
  NAND2_X1 U108 ( .A1(\mem[6][1] ), .A2(n1154), .ZN(n1152) );
  OAI21_X1 U109 ( .B1(n626), .B2(n1154), .A(n1151), .ZN(n864) );
  NAND2_X1 U110 ( .A1(\mem[6][2] ), .A2(n1154), .ZN(n1151) );
  OAI21_X1 U111 ( .B1(n627), .B2(n1154), .A(n1150), .ZN(n863) );
  NAND2_X1 U112 ( .A1(\mem[6][3] ), .A2(n1154), .ZN(n1150) );
  OAI21_X1 U113 ( .B1(n628), .B2(n1154), .A(n1149), .ZN(n862) );
  NAND2_X1 U114 ( .A1(\mem[6][4] ), .A2(n1154), .ZN(n1149) );
  OAI21_X1 U115 ( .B1(n629), .B2(n1154), .A(n1148), .ZN(n861) );
  NAND2_X1 U116 ( .A1(\mem[6][5] ), .A2(n1154), .ZN(n1148) );
  OAI21_X1 U117 ( .B1(n630), .B2(n1154), .A(n1147), .ZN(n860) );
  NAND2_X1 U118 ( .A1(\mem[6][6] ), .A2(n1154), .ZN(n1147) );
  OAI21_X1 U119 ( .B1(n631), .B2(n1154), .A(n1146), .ZN(n859) );
  NAND2_X1 U120 ( .A1(\mem[6][7] ), .A2(n1154), .ZN(n1146) );
  OAI21_X1 U121 ( .B1(n624), .B2(n1144), .A(n1143), .ZN(n858) );
  NAND2_X1 U122 ( .A1(\mem[7][0] ), .A2(n1144), .ZN(n1143) );
  OAI21_X1 U123 ( .B1(n625), .B2(n1144), .A(n1142), .ZN(n857) );
  NAND2_X1 U124 ( .A1(\mem[7][1] ), .A2(n1144), .ZN(n1142) );
  OAI21_X1 U125 ( .B1(n626), .B2(n1144), .A(n1141), .ZN(n856) );
  NAND2_X1 U126 ( .A1(\mem[7][2] ), .A2(n1144), .ZN(n1141) );
  OAI21_X1 U127 ( .B1(n627), .B2(n1144), .A(n1140), .ZN(n855) );
  NAND2_X1 U128 ( .A1(\mem[7][3] ), .A2(n1144), .ZN(n1140) );
  OAI21_X1 U129 ( .B1(n628), .B2(n1144), .A(n1139), .ZN(n854) );
  NAND2_X1 U130 ( .A1(\mem[7][4] ), .A2(n1144), .ZN(n1139) );
  OAI21_X1 U131 ( .B1(n629), .B2(n1144), .A(n1138), .ZN(n853) );
  NAND2_X1 U132 ( .A1(\mem[7][5] ), .A2(n1144), .ZN(n1138) );
  OAI21_X1 U133 ( .B1(n630), .B2(n1144), .A(n1137), .ZN(n852) );
  NAND2_X1 U134 ( .A1(\mem[7][6] ), .A2(n1144), .ZN(n1137) );
  OAI21_X1 U135 ( .B1(n631), .B2(n1144), .A(n1136), .ZN(n851) );
  NAND2_X1 U136 ( .A1(\mem[7][7] ), .A2(n1144), .ZN(n1136) );
  OAI21_X1 U137 ( .B1(n624), .B2(n1204), .A(n1203), .ZN(n906) );
  NAND2_X1 U138 ( .A1(\mem[1][0] ), .A2(n1204), .ZN(n1203) );
  OAI21_X1 U139 ( .B1(n625), .B2(n1204), .A(n1202), .ZN(n905) );
  NAND2_X1 U140 ( .A1(\mem[1][1] ), .A2(n1204), .ZN(n1202) );
  OAI21_X1 U141 ( .B1(n626), .B2(n1204), .A(n1201), .ZN(n904) );
  NAND2_X1 U142 ( .A1(\mem[1][2] ), .A2(n1204), .ZN(n1201) );
  OAI21_X1 U143 ( .B1(n627), .B2(n1204), .A(n1200), .ZN(n903) );
  NAND2_X1 U144 ( .A1(\mem[1][3] ), .A2(n1204), .ZN(n1200) );
  OAI21_X1 U145 ( .B1(n628), .B2(n1204), .A(n1199), .ZN(n902) );
  NAND2_X1 U146 ( .A1(\mem[1][4] ), .A2(n1204), .ZN(n1199) );
  OAI21_X1 U147 ( .B1(n629), .B2(n1204), .A(n1198), .ZN(n901) );
  NAND2_X1 U148 ( .A1(\mem[1][5] ), .A2(n1204), .ZN(n1198) );
  OAI21_X1 U149 ( .B1(n630), .B2(n1204), .A(n1197), .ZN(n900) );
  NAND2_X1 U150 ( .A1(\mem[1][6] ), .A2(n1204), .ZN(n1197) );
  OAI21_X1 U151 ( .B1(n631), .B2(n1204), .A(n1196), .ZN(n899) );
  NAND2_X1 U152 ( .A1(\mem[1][7] ), .A2(n1204), .ZN(n1196) );
  OAI21_X1 U153 ( .B1(n624), .B2(n1194), .A(n1193), .ZN(n898) );
  NAND2_X1 U154 ( .A1(\mem[2][0] ), .A2(n1194), .ZN(n1193) );
  OAI21_X1 U155 ( .B1(n625), .B2(n1194), .A(n1192), .ZN(n897) );
  NAND2_X1 U156 ( .A1(\mem[2][1] ), .A2(n1194), .ZN(n1192) );
  OAI21_X1 U157 ( .B1(n626), .B2(n1194), .A(n1191), .ZN(n896) );
  NAND2_X1 U158 ( .A1(\mem[2][2] ), .A2(n1194), .ZN(n1191) );
  OAI21_X1 U159 ( .B1(n627), .B2(n1194), .A(n1190), .ZN(n895) );
  NAND2_X1 U160 ( .A1(\mem[2][3] ), .A2(n1194), .ZN(n1190) );
  OAI21_X1 U161 ( .B1(n628), .B2(n1194), .A(n1189), .ZN(n894) );
  NAND2_X1 U162 ( .A1(\mem[2][4] ), .A2(n1194), .ZN(n1189) );
  OAI21_X1 U163 ( .B1(n629), .B2(n1194), .A(n1188), .ZN(n893) );
  NAND2_X1 U164 ( .A1(\mem[2][5] ), .A2(n1194), .ZN(n1188) );
  OAI21_X1 U165 ( .B1(n630), .B2(n1194), .A(n1187), .ZN(n892) );
  NAND2_X1 U166 ( .A1(\mem[2][6] ), .A2(n1194), .ZN(n1187) );
  OAI21_X1 U167 ( .B1(n631), .B2(n1194), .A(n1186), .ZN(n891) );
  NAND2_X1 U168 ( .A1(\mem[2][7] ), .A2(n1194), .ZN(n1186) );
  OAI21_X1 U169 ( .B1(n624), .B2(n1184), .A(n1183), .ZN(n890) );
  NAND2_X1 U170 ( .A1(\mem[3][0] ), .A2(n1184), .ZN(n1183) );
  OAI21_X1 U171 ( .B1(n625), .B2(n1184), .A(n1182), .ZN(n889) );
  NAND2_X1 U172 ( .A1(\mem[3][1] ), .A2(n1184), .ZN(n1182) );
  OAI21_X1 U173 ( .B1(n626), .B2(n1184), .A(n1181), .ZN(n888) );
  NAND2_X1 U174 ( .A1(\mem[3][2] ), .A2(n1184), .ZN(n1181) );
  OAI21_X1 U175 ( .B1(n627), .B2(n1184), .A(n1180), .ZN(n887) );
  NAND2_X1 U176 ( .A1(\mem[3][3] ), .A2(n1184), .ZN(n1180) );
  OAI21_X1 U177 ( .B1(n628), .B2(n1184), .A(n1179), .ZN(n886) );
  NAND2_X1 U178 ( .A1(\mem[3][4] ), .A2(n1184), .ZN(n1179) );
  OAI21_X1 U179 ( .B1(n629), .B2(n1184), .A(n1178), .ZN(n885) );
  NAND2_X1 U180 ( .A1(\mem[3][5] ), .A2(n1184), .ZN(n1178) );
  OAI21_X1 U181 ( .B1(n630), .B2(n1184), .A(n1177), .ZN(n884) );
  NAND2_X1 U182 ( .A1(\mem[3][6] ), .A2(n1184), .ZN(n1177) );
  OAI21_X1 U183 ( .B1(n631), .B2(n1184), .A(n1176), .ZN(n883) );
  NAND2_X1 U184 ( .A1(\mem[3][7] ), .A2(n1184), .ZN(n1176) );
  OAI21_X1 U185 ( .B1(n624), .B2(n1164), .A(n1163), .ZN(n874) );
  NAND2_X1 U186 ( .A1(\mem[5][0] ), .A2(n1164), .ZN(n1163) );
  OAI21_X1 U187 ( .B1(n625), .B2(n1164), .A(n1162), .ZN(n873) );
  NAND2_X1 U188 ( .A1(\mem[5][1] ), .A2(n1164), .ZN(n1162) );
  OAI21_X1 U189 ( .B1(n626), .B2(n1164), .A(n1161), .ZN(n872) );
  NAND2_X1 U190 ( .A1(\mem[5][2] ), .A2(n1164), .ZN(n1161) );
  OAI21_X1 U191 ( .B1(n627), .B2(n1164), .A(n1160), .ZN(n871) );
  NAND2_X1 U192 ( .A1(\mem[5][3] ), .A2(n1164), .ZN(n1160) );
  OAI21_X1 U193 ( .B1(n628), .B2(n1164), .A(n1159), .ZN(n870) );
  NAND2_X1 U194 ( .A1(\mem[5][4] ), .A2(n1164), .ZN(n1159) );
  OAI21_X1 U195 ( .B1(n629), .B2(n1164), .A(n1158), .ZN(n869) );
  NAND2_X1 U196 ( .A1(\mem[5][5] ), .A2(n1164), .ZN(n1158) );
  OAI21_X1 U197 ( .B1(n630), .B2(n1164), .A(n1157), .ZN(n868) );
  NAND2_X1 U198 ( .A1(\mem[5][6] ), .A2(n1164), .ZN(n1157) );
  OAI21_X1 U199 ( .B1(n631), .B2(n1164), .A(n1156), .ZN(n867) );
  NAND2_X1 U200 ( .A1(\mem[5][7] ), .A2(n1164), .ZN(n1156) );
  OAI21_X1 U201 ( .B1(n1215), .B2(n624), .A(n1214), .ZN(n914) );
  NAND2_X1 U202 ( .A1(\mem[0][0] ), .A2(n1215), .ZN(n1214) );
  OAI21_X1 U203 ( .B1(n1215), .B2(n625), .A(n1213), .ZN(n913) );
  NAND2_X1 U204 ( .A1(\mem[0][1] ), .A2(n1215), .ZN(n1213) );
  OAI21_X1 U205 ( .B1(n1215), .B2(n626), .A(n1212), .ZN(n912) );
  NAND2_X1 U206 ( .A1(\mem[0][2] ), .A2(n1215), .ZN(n1212) );
  OAI21_X1 U207 ( .B1(n1215), .B2(n627), .A(n1211), .ZN(n911) );
  NAND2_X1 U208 ( .A1(\mem[0][3] ), .A2(n1215), .ZN(n1211) );
  OAI21_X1 U209 ( .B1(n1215), .B2(n628), .A(n1210), .ZN(n910) );
  NAND2_X1 U210 ( .A1(\mem[0][4] ), .A2(n1215), .ZN(n1210) );
  OAI21_X1 U211 ( .B1(n1215), .B2(n629), .A(n1209), .ZN(n909) );
  NAND2_X1 U212 ( .A1(\mem[0][5] ), .A2(n1215), .ZN(n1209) );
  OAI21_X1 U213 ( .B1(n1215), .B2(n630), .A(n1208), .ZN(n908) );
  NAND2_X1 U214 ( .A1(\mem[0][6] ), .A2(n1215), .ZN(n1208) );
  OAI21_X1 U215 ( .B1(n1215), .B2(n631), .A(n1207), .ZN(n907) );
  NAND2_X1 U216 ( .A1(\mem[0][7] ), .A2(n1215), .ZN(n1207) );
  INV_X1 U217 ( .A(n1133), .ZN(n823) );
  AOI22_X1 U218 ( .A1(data_in[0]), .A2(n847), .B1(n1132), .B2(\mem[8][0] ), 
        .ZN(n1133) );
  INV_X1 U219 ( .A(n1131), .ZN(n822) );
  AOI22_X1 U220 ( .A1(data_in[1]), .A2(n847), .B1(n1132), .B2(\mem[8][1] ), 
        .ZN(n1131) );
  INV_X1 U221 ( .A(n1130), .ZN(n821) );
  AOI22_X1 U222 ( .A1(data_in[2]), .A2(n847), .B1(n1132), .B2(\mem[8][2] ), 
        .ZN(n1130) );
  INV_X1 U223 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U224 ( .A1(data_in[3]), .A2(n847), .B1(n1132), .B2(\mem[8][3] ), 
        .ZN(n1129) );
  INV_X1 U225 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U226 ( .A1(data_in[4]), .A2(n847), .B1(n1132), .B2(\mem[8][4] ), 
        .ZN(n1128) );
  INV_X1 U227 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U228 ( .A1(data_in[5]), .A2(n847), .B1(n1132), .B2(\mem[8][5] ), 
        .ZN(n1127) );
  INV_X1 U229 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U230 ( .A1(data_in[6]), .A2(n847), .B1(n1132), .B2(\mem[8][6] ), 
        .ZN(n1126) );
  INV_X1 U231 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U232 ( .A1(data_in[7]), .A2(n847), .B1(n1132), .B2(\mem[8][7] ), 
        .ZN(n1125) );
  INV_X1 U233 ( .A(n1123), .ZN(n815) );
  AOI22_X1 U234 ( .A1(data_in[0]), .A2(n846), .B1(n1122), .B2(\mem[9][0] ), 
        .ZN(n1123) );
  INV_X1 U235 ( .A(n1121), .ZN(n814) );
  AOI22_X1 U236 ( .A1(data_in[1]), .A2(n846), .B1(n1122), .B2(\mem[9][1] ), 
        .ZN(n1121) );
  INV_X1 U237 ( .A(n1120), .ZN(n813) );
  AOI22_X1 U238 ( .A1(data_in[2]), .A2(n846), .B1(n1122), .B2(\mem[9][2] ), 
        .ZN(n1120) );
  INV_X1 U239 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U240 ( .A1(data_in[3]), .A2(n846), .B1(n1122), .B2(\mem[9][3] ), 
        .ZN(n1119) );
  INV_X1 U241 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U242 ( .A1(data_in[4]), .A2(n846), .B1(n1122), .B2(\mem[9][4] ), 
        .ZN(n1118) );
  INV_X1 U243 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U244 ( .A1(data_in[5]), .A2(n846), .B1(n1122), .B2(\mem[9][5] ), 
        .ZN(n1117) );
  INV_X1 U245 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U246 ( .A1(data_in[6]), .A2(n846), .B1(n1122), .B2(\mem[9][6] ), 
        .ZN(n1116) );
  INV_X1 U247 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U248 ( .A1(data_in[7]), .A2(n846), .B1(n1122), .B2(\mem[9][7] ), 
        .ZN(n1115) );
  INV_X1 U249 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U250 ( .A1(data_in[0]), .A2(n845), .B1(n1113), .B2(\mem[10][0] ), 
        .ZN(n1114) );
  INV_X1 U251 ( .A(n1112), .ZN(n806) );
  AOI22_X1 U252 ( .A1(data_in[1]), .A2(n845), .B1(n1113), .B2(\mem[10][1] ), 
        .ZN(n1112) );
  INV_X1 U253 ( .A(n1111), .ZN(n805) );
  AOI22_X1 U254 ( .A1(data_in[2]), .A2(n845), .B1(n1113), .B2(\mem[10][2] ), 
        .ZN(n1111) );
  INV_X1 U255 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U256 ( .A1(data_in[3]), .A2(n845), .B1(n1113), .B2(\mem[10][3] ), 
        .ZN(n1110) );
  INV_X1 U257 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U258 ( .A1(data_in[4]), .A2(n845), .B1(n1113), .B2(\mem[10][4] ), 
        .ZN(n1109) );
  INV_X1 U259 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U260 ( .A1(data_in[5]), .A2(n845), .B1(n1113), .B2(\mem[10][5] ), 
        .ZN(n1108) );
  INV_X1 U261 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U262 ( .A1(data_in[6]), .A2(n845), .B1(n1113), .B2(\mem[10][6] ), 
        .ZN(n1107) );
  INV_X1 U263 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U264 ( .A1(data_in[7]), .A2(n845), .B1(n1113), .B2(\mem[10][7] ), 
        .ZN(n1106) );
  INV_X1 U265 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U266 ( .A1(data_in[0]), .A2(n844), .B1(n1104), .B2(\mem[11][0] ), 
        .ZN(n1105) );
  INV_X1 U267 ( .A(n1103), .ZN(n798) );
  AOI22_X1 U268 ( .A1(data_in[1]), .A2(n844), .B1(n1104), .B2(\mem[11][1] ), 
        .ZN(n1103) );
  INV_X1 U269 ( .A(n1102), .ZN(n797) );
  AOI22_X1 U270 ( .A1(data_in[2]), .A2(n844), .B1(n1104), .B2(\mem[11][2] ), 
        .ZN(n1102) );
  INV_X1 U271 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U272 ( .A1(data_in[3]), .A2(n844), .B1(n1104), .B2(\mem[11][3] ), 
        .ZN(n1101) );
  INV_X1 U273 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U274 ( .A1(data_in[4]), .A2(n844), .B1(n1104), .B2(\mem[11][4] ), 
        .ZN(n1100) );
  INV_X1 U275 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U276 ( .A1(data_in[5]), .A2(n844), .B1(n1104), .B2(\mem[11][5] ), 
        .ZN(n1099) );
  INV_X1 U277 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U278 ( .A1(data_in[6]), .A2(n844), .B1(n1104), .B2(\mem[11][6] ), 
        .ZN(n1098) );
  INV_X1 U279 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U280 ( .A1(data_in[7]), .A2(n844), .B1(n1104), .B2(\mem[11][7] ), 
        .ZN(n1097) );
  INV_X1 U281 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U282 ( .A1(data_in[0]), .A2(n843), .B1(n1095), .B2(\mem[12][0] ), 
        .ZN(n1096) );
  INV_X1 U283 ( .A(n1094), .ZN(n790) );
  AOI22_X1 U284 ( .A1(data_in[1]), .A2(n843), .B1(n1095), .B2(\mem[12][1] ), 
        .ZN(n1094) );
  INV_X1 U285 ( .A(n1093), .ZN(n789) );
  AOI22_X1 U286 ( .A1(data_in[2]), .A2(n843), .B1(n1095), .B2(\mem[12][2] ), 
        .ZN(n1093) );
  INV_X1 U287 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U288 ( .A1(data_in[3]), .A2(n843), .B1(n1095), .B2(\mem[12][3] ), 
        .ZN(n1092) );
  INV_X1 U289 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U290 ( .A1(data_in[4]), .A2(n843), .B1(n1095), .B2(\mem[12][4] ), 
        .ZN(n1091) );
  INV_X1 U291 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U292 ( .A1(data_in[5]), .A2(n843), .B1(n1095), .B2(\mem[12][5] ), 
        .ZN(n1090) );
  INV_X1 U293 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U294 ( .A1(data_in[6]), .A2(n843), .B1(n1095), .B2(\mem[12][6] ), 
        .ZN(n1089) );
  INV_X1 U295 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U296 ( .A1(data_in[7]), .A2(n843), .B1(n1095), .B2(\mem[12][7] ), 
        .ZN(n1088) );
  INV_X1 U297 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U298 ( .A1(data_in[0]), .A2(n842), .B1(n1086), .B2(\mem[13][0] ), 
        .ZN(n1087) );
  INV_X1 U299 ( .A(n1085), .ZN(n782) );
  AOI22_X1 U300 ( .A1(data_in[1]), .A2(n842), .B1(n1086), .B2(\mem[13][1] ), 
        .ZN(n1085) );
  INV_X1 U301 ( .A(n1084), .ZN(n781) );
  AOI22_X1 U302 ( .A1(data_in[2]), .A2(n842), .B1(n1086), .B2(\mem[13][2] ), 
        .ZN(n1084) );
  INV_X1 U303 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U304 ( .A1(data_in[3]), .A2(n842), .B1(n1086), .B2(\mem[13][3] ), 
        .ZN(n1083) );
  INV_X1 U305 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U306 ( .A1(data_in[4]), .A2(n842), .B1(n1086), .B2(\mem[13][4] ), 
        .ZN(n1082) );
  INV_X1 U307 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U308 ( .A1(data_in[5]), .A2(n842), .B1(n1086), .B2(\mem[13][5] ), 
        .ZN(n1081) );
  INV_X1 U309 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U310 ( .A1(data_in[6]), .A2(n842), .B1(n1086), .B2(\mem[13][6] ), 
        .ZN(n1080) );
  INV_X1 U311 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U312 ( .A1(data_in[7]), .A2(n842), .B1(n1086), .B2(\mem[13][7] ), 
        .ZN(n1079) );
  INV_X1 U313 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U314 ( .A1(data_in[0]), .A2(n841), .B1(n1077), .B2(\mem[14][0] ), 
        .ZN(n1078) );
  INV_X1 U315 ( .A(n1076), .ZN(n774) );
  AOI22_X1 U316 ( .A1(data_in[1]), .A2(n841), .B1(n1077), .B2(\mem[14][1] ), 
        .ZN(n1076) );
  INV_X1 U317 ( .A(n1075), .ZN(n773) );
  AOI22_X1 U318 ( .A1(data_in[2]), .A2(n841), .B1(n1077), .B2(\mem[14][2] ), 
        .ZN(n1075) );
  INV_X1 U319 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U320 ( .A1(data_in[3]), .A2(n841), .B1(n1077), .B2(\mem[14][3] ), 
        .ZN(n1074) );
  INV_X1 U321 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U322 ( .A1(data_in[4]), .A2(n841), .B1(n1077), .B2(\mem[14][4] ), 
        .ZN(n1073) );
  INV_X1 U323 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U324 ( .A1(data_in[5]), .A2(n841), .B1(n1077), .B2(\mem[14][5] ), 
        .ZN(n1072) );
  INV_X1 U325 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U326 ( .A1(data_in[6]), .A2(n841), .B1(n1077), .B2(\mem[14][6] ), 
        .ZN(n1071) );
  INV_X1 U327 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U328 ( .A1(data_in[7]), .A2(n841), .B1(n1077), .B2(\mem[14][7] ), 
        .ZN(n1070) );
  INV_X1 U329 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U330 ( .A1(data_in[0]), .A2(n840), .B1(n1068), .B2(\mem[15][0] ), 
        .ZN(n1069) );
  INV_X1 U331 ( .A(n1067), .ZN(n766) );
  AOI22_X1 U332 ( .A1(data_in[1]), .A2(n840), .B1(n1068), .B2(\mem[15][1] ), 
        .ZN(n1067) );
  INV_X1 U333 ( .A(n1066), .ZN(n765) );
  AOI22_X1 U334 ( .A1(data_in[2]), .A2(n840), .B1(n1068), .B2(\mem[15][2] ), 
        .ZN(n1066) );
  INV_X1 U335 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U336 ( .A1(data_in[3]), .A2(n840), .B1(n1068), .B2(\mem[15][3] ), 
        .ZN(n1065) );
  INV_X1 U337 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U338 ( .A1(data_in[4]), .A2(n840), .B1(n1068), .B2(\mem[15][4] ), 
        .ZN(n1064) );
  INV_X1 U339 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U340 ( .A1(data_in[5]), .A2(n840), .B1(n1068), .B2(\mem[15][5] ), 
        .ZN(n1063) );
  INV_X1 U341 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U342 ( .A1(data_in[6]), .A2(n840), .B1(n1068), .B2(\mem[15][6] ), 
        .ZN(n1062) );
  INV_X1 U343 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U344 ( .A1(data_in[7]), .A2(n840), .B1(n1068), .B2(\mem[15][7] ), 
        .ZN(n1061) );
  INV_X1 U345 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U346 ( .A1(data_in[0]), .A2(n839), .B1(n1059), .B2(\mem[16][0] ), 
        .ZN(n1060) );
  INV_X1 U347 ( .A(n1058), .ZN(n758) );
  AOI22_X1 U348 ( .A1(data_in[1]), .A2(n839), .B1(n1059), .B2(\mem[16][1] ), 
        .ZN(n1058) );
  INV_X1 U349 ( .A(n1057), .ZN(n757) );
  AOI22_X1 U350 ( .A1(data_in[2]), .A2(n839), .B1(n1059), .B2(\mem[16][2] ), 
        .ZN(n1057) );
  INV_X1 U351 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U352 ( .A1(data_in[3]), .A2(n839), .B1(n1059), .B2(\mem[16][3] ), 
        .ZN(n1056) );
  INV_X1 U353 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U354 ( .A1(data_in[4]), .A2(n839), .B1(n1059), .B2(\mem[16][4] ), 
        .ZN(n1055) );
  INV_X1 U355 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U356 ( .A1(data_in[5]), .A2(n839), .B1(n1059), .B2(\mem[16][5] ), 
        .ZN(n1054) );
  INV_X1 U357 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U358 ( .A1(data_in[6]), .A2(n839), .B1(n1059), .B2(\mem[16][6] ), 
        .ZN(n1053) );
  INV_X1 U359 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U360 ( .A1(data_in[7]), .A2(n839), .B1(n1059), .B2(\mem[16][7] ), 
        .ZN(n1052) );
  INV_X1 U361 ( .A(n1050), .ZN(n751) );
  AOI22_X1 U362 ( .A1(data_in[0]), .A2(n838), .B1(n1049), .B2(\mem[17][0] ), 
        .ZN(n1050) );
  INV_X1 U363 ( .A(n1048), .ZN(n750) );
  AOI22_X1 U364 ( .A1(data_in[1]), .A2(n838), .B1(n1049), .B2(\mem[17][1] ), 
        .ZN(n1048) );
  INV_X1 U365 ( .A(n1047), .ZN(n749) );
  AOI22_X1 U366 ( .A1(data_in[2]), .A2(n838), .B1(n1049), .B2(\mem[17][2] ), 
        .ZN(n1047) );
  INV_X1 U367 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U368 ( .A1(data_in[3]), .A2(n838), .B1(n1049), .B2(\mem[17][3] ), 
        .ZN(n1046) );
  INV_X1 U369 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U370 ( .A1(data_in[4]), .A2(n838), .B1(n1049), .B2(\mem[17][4] ), 
        .ZN(n1045) );
  INV_X1 U371 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U372 ( .A1(data_in[5]), .A2(n838), .B1(n1049), .B2(\mem[17][5] ), 
        .ZN(n1044) );
  INV_X1 U373 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U374 ( .A1(data_in[6]), .A2(n838), .B1(n1049), .B2(\mem[17][6] ), 
        .ZN(n1043) );
  INV_X1 U375 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U376 ( .A1(data_in[7]), .A2(n838), .B1(n1049), .B2(\mem[17][7] ), 
        .ZN(n1042) );
  INV_X1 U377 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U378 ( .A1(data_in[0]), .A2(n837), .B1(n1040), .B2(\mem[18][0] ), 
        .ZN(n1041) );
  INV_X1 U379 ( .A(n1039), .ZN(n742) );
  AOI22_X1 U380 ( .A1(data_in[1]), .A2(n837), .B1(n1040), .B2(\mem[18][1] ), 
        .ZN(n1039) );
  INV_X1 U381 ( .A(n1038), .ZN(n741) );
  AOI22_X1 U382 ( .A1(data_in[2]), .A2(n837), .B1(n1040), .B2(\mem[18][2] ), 
        .ZN(n1038) );
  INV_X1 U383 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U384 ( .A1(data_in[3]), .A2(n837), .B1(n1040), .B2(\mem[18][3] ), 
        .ZN(n1037) );
  INV_X1 U385 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U386 ( .A1(data_in[4]), .A2(n837), .B1(n1040), .B2(\mem[18][4] ), 
        .ZN(n1036) );
  INV_X1 U387 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U388 ( .A1(data_in[5]), .A2(n837), .B1(n1040), .B2(\mem[18][5] ), 
        .ZN(n1035) );
  INV_X1 U389 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U390 ( .A1(data_in[6]), .A2(n837), .B1(n1040), .B2(\mem[18][6] ), 
        .ZN(n1034) );
  INV_X1 U391 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U392 ( .A1(data_in[7]), .A2(n837), .B1(n1040), .B2(\mem[18][7] ), 
        .ZN(n1033) );
  INV_X1 U393 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U394 ( .A1(data_in[0]), .A2(n836), .B1(n1031), .B2(\mem[19][0] ), 
        .ZN(n1032) );
  INV_X1 U395 ( .A(n1030), .ZN(n734) );
  AOI22_X1 U396 ( .A1(data_in[1]), .A2(n836), .B1(n1031), .B2(\mem[19][1] ), 
        .ZN(n1030) );
  INV_X1 U397 ( .A(n1029), .ZN(n733) );
  AOI22_X1 U398 ( .A1(data_in[2]), .A2(n836), .B1(n1031), .B2(\mem[19][2] ), 
        .ZN(n1029) );
  INV_X1 U399 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U400 ( .A1(data_in[3]), .A2(n836), .B1(n1031), .B2(\mem[19][3] ), 
        .ZN(n1028) );
  INV_X1 U401 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U402 ( .A1(data_in[4]), .A2(n836), .B1(n1031), .B2(\mem[19][4] ), 
        .ZN(n1027) );
  INV_X1 U403 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U404 ( .A1(data_in[5]), .A2(n836), .B1(n1031), .B2(\mem[19][5] ), 
        .ZN(n1026) );
  INV_X1 U405 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U406 ( .A1(data_in[6]), .A2(n836), .B1(n1031), .B2(\mem[19][6] ), 
        .ZN(n1025) );
  INV_X1 U407 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U408 ( .A1(data_in[7]), .A2(n836), .B1(n1031), .B2(\mem[19][7] ), 
        .ZN(n1024) );
  INV_X1 U409 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U410 ( .A1(data_in[0]), .A2(n835), .B1(n1022), .B2(\mem[20][0] ), 
        .ZN(n1023) );
  INV_X1 U411 ( .A(n1021), .ZN(n726) );
  AOI22_X1 U412 ( .A1(data_in[1]), .A2(n835), .B1(n1022), .B2(\mem[20][1] ), 
        .ZN(n1021) );
  INV_X1 U413 ( .A(n1020), .ZN(n725) );
  AOI22_X1 U414 ( .A1(data_in[2]), .A2(n835), .B1(n1022), .B2(\mem[20][2] ), 
        .ZN(n1020) );
  INV_X1 U415 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U416 ( .A1(data_in[3]), .A2(n835), .B1(n1022), .B2(\mem[20][3] ), 
        .ZN(n1019) );
  INV_X1 U417 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U418 ( .A1(data_in[4]), .A2(n835), .B1(n1022), .B2(\mem[20][4] ), 
        .ZN(n1018) );
  INV_X1 U419 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U420 ( .A1(data_in[5]), .A2(n835), .B1(n1022), .B2(\mem[20][5] ), 
        .ZN(n1017) );
  INV_X1 U421 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U422 ( .A1(data_in[6]), .A2(n835), .B1(n1022), .B2(\mem[20][6] ), 
        .ZN(n1016) );
  INV_X1 U423 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U424 ( .A1(data_in[7]), .A2(n835), .B1(n1022), .B2(\mem[20][7] ), 
        .ZN(n1015) );
  INV_X1 U425 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U426 ( .A1(data_in[0]), .A2(n834), .B1(n1013), .B2(\mem[21][0] ), 
        .ZN(n1014) );
  INV_X1 U427 ( .A(n1012), .ZN(n718) );
  AOI22_X1 U428 ( .A1(data_in[1]), .A2(n834), .B1(n1013), .B2(\mem[21][1] ), 
        .ZN(n1012) );
  INV_X1 U429 ( .A(n1011), .ZN(n717) );
  AOI22_X1 U430 ( .A1(data_in[2]), .A2(n834), .B1(n1013), .B2(\mem[21][2] ), 
        .ZN(n1011) );
  INV_X1 U431 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U432 ( .A1(data_in[3]), .A2(n834), .B1(n1013), .B2(\mem[21][3] ), 
        .ZN(n1010) );
  INV_X1 U433 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U434 ( .A1(data_in[4]), .A2(n834), .B1(n1013), .B2(\mem[21][4] ), 
        .ZN(n1009) );
  INV_X1 U435 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U436 ( .A1(data_in[5]), .A2(n834), .B1(n1013), .B2(\mem[21][5] ), 
        .ZN(n1008) );
  INV_X1 U437 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U438 ( .A1(data_in[6]), .A2(n834), .B1(n1013), .B2(\mem[21][6] ), 
        .ZN(n1007) );
  INV_X1 U439 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U440 ( .A1(data_in[7]), .A2(n834), .B1(n1013), .B2(\mem[21][7] ), 
        .ZN(n1006) );
  INV_X1 U441 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U442 ( .A1(data_in[0]), .A2(n833), .B1(n1004), .B2(\mem[22][0] ), 
        .ZN(n1005) );
  INV_X1 U443 ( .A(n1003), .ZN(n710) );
  AOI22_X1 U444 ( .A1(data_in[1]), .A2(n833), .B1(n1004), .B2(\mem[22][1] ), 
        .ZN(n1003) );
  INV_X1 U445 ( .A(n1002), .ZN(n709) );
  AOI22_X1 U446 ( .A1(data_in[2]), .A2(n833), .B1(n1004), .B2(\mem[22][2] ), 
        .ZN(n1002) );
  INV_X1 U447 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U448 ( .A1(data_in[3]), .A2(n833), .B1(n1004), .B2(\mem[22][3] ), 
        .ZN(n1001) );
  INV_X1 U449 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U450 ( .A1(data_in[4]), .A2(n833), .B1(n1004), .B2(\mem[22][4] ), 
        .ZN(n1000) );
  INV_X1 U451 ( .A(n999), .ZN(n706) );
  AOI22_X1 U452 ( .A1(data_in[5]), .A2(n833), .B1(n1004), .B2(\mem[22][5] ), 
        .ZN(n999) );
  INV_X1 U453 ( .A(n998), .ZN(n705) );
  AOI22_X1 U454 ( .A1(data_in[6]), .A2(n833), .B1(n1004), .B2(\mem[22][6] ), 
        .ZN(n998) );
  INV_X1 U455 ( .A(n997), .ZN(n704) );
  AOI22_X1 U456 ( .A1(data_in[7]), .A2(n833), .B1(n1004), .B2(\mem[22][7] ), 
        .ZN(n997) );
  INV_X1 U457 ( .A(n996), .ZN(n703) );
  AOI22_X1 U458 ( .A1(data_in[0]), .A2(n832), .B1(n995), .B2(\mem[23][0] ), 
        .ZN(n996) );
  INV_X1 U459 ( .A(n994), .ZN(n702) );
  AOI22_X1 U460 ( .A1(data_in[1]), .A2(n832), .B1(n995), .B2(\mem[23][1] ), 
        .ZN(n994) );
  INV_X1 U461 ( .A(n993), .ZN(n701) );
  AOI22_X1 U462 ( .A1(data_in[2]), .A2(n832), .B1(n995), .B2(\mem[23][2] ), 
        .ZN(n993) );
  INV_X1 U463 ( .A(n992), .ZN(n700) );
  AOI22_X1 U464 ( .A1(data_in[3]), .A2(n832), .B1(n995), .B2(\mem[23][3] ), 
        .ZN(n992) );
  INV_X1 U465 ( .A(n991), .ZN(n699) );
  AOI22_X1 U466 ( .A1(data_in[4]), .A2(n832), .B1(n995), .B2(\mem[23][4] ), 
        .ZN(n991) );
  INV_X1 U467 ( .A(n990), .ZN(n698) );
  AOI22_X1 U468 ( .A1(data_in[5]), .A2(n832), .B1(n995), .B2(\mem[23][5] ), 
        .ZN(n990) );
  INV_X1 U469 ( .A(n989), .ZN(n697) );
  AOI22_X1 U470 ( .A1(data_in[6]), .A2(n832), .B1(n995), .B2(\mem[23][6] ), 
        .ZN(n989) );
  INV_X1 U471 ( .A(n988), .ZN(n696) );
  AOI22_X1 U472 ( .A1(data_in[7]), .A2(n832), .B1(n995), .B2(\mem[23][7] ), 
        .ZN(n988) );
  INV_X1 U473 ( .A(n987), .ZN(n695) );
  AOI22_X1 U474 ( .A1(data_in[0]), .A2(n831), .B1(n986), .B2(\mem[24][0] ), 
        .ZN(n987) );
  INV_X1 U475 ( .A(n985), .ZN(n694) );
  AOI22_X1 U476 ( .A1(data_in[1]), .A2(n831), .B1(n986), .B2(\mem[24][1] ), 
        .ZN(n985) );
  INV_X1 U477 ( .A(n984), .ZN(n693) );
  AOI22_X1 U478 ( .A1(data_in[2]), .A2(n831), .B1(n986), .B2(\mem[24][2] ), 
        .ZN(n984) );
  INV_X1 U479 ( .A(n983), .ZN(n692) );
  AOI22_X1 U480 ( .A1(data_in[3]), .A2(n831), .B1(n986), .B2(\mem[24][3] ), 
        .ZN(n983) );
  INV_X1 U481 ( .A(n982), .ZN(n691) );
  AOI22_X1 U482 ( .A1(data_in[4]), .A2(n831), .B1(n986), .B2(\mem[24][4] ), 
        .ZN(n982) );
  INV_X1 U483 ( .A(n981), .ZN(n690) );
  AOI22_X1 U484 ( .A1(data_in[5]), .A2(n831), .B1(n986), .B2(\mem[24][5] ), 
        .ZN(n981) );
  INV_X1 U485 ( .A(n980), .ZN(n689) );
  AOI22_X1 U486 ( .A1(data_in[6]), .A2(n831), .B1(n986), .B2(\mem[24][6] ), 
        .ZN(n980) );
  INV_X1 U487 ( .A(n979), .ZN(n688) );
  AOI22_X1 U488 ( .A1(data_in[7]), .A2(n831), .B1(n986), .B2(\mem[24][7] ), 
        .ZN(n979) );
  INV_X1 U489 ( .A(n977), .ZN(n687) );
  AOI22_X1 U490 ( .A1(data_in[0]), .A2(n830), .B1(n976), .B2(\mem[25][0] ), 
        .ZN(n977) );
  INV_X1 U491 ( .A(n975), .ZN(n686) );
  AOI22_X1 U492 ( .A1(data_in[1]), .A2(n830), .B1(n976), .B2(\mem[25][1] ), 
        .ZN(n975) );
  INV_X1 U493 ( .A(n974), .ZN(n685) );
  AOI22_X1 U494 ( .A1(data_in[2]), .A2(n830), .B1(n976), .B2(\mem[25][2] ), 
        .ZN(n974) );
  INV_X1 U495 ( .A(n973), .ZN(n684) );
  AOI22_X1 U496 ( .A1(data_in[3]), .A2(n830), .B1(n976), .B2(\mem[25][3] ), 
        .ZN(n973) );
  INV_X1 U497 ( .A(n972), .ZN(n683) );
  AOI22_X1 U498 ( .A1(data_in[4]), .A2(n830), .B1(n976), .B2(\mem[25][4] ), 
        .ZN(n972) );
  INV_X1 U499 ( .A(n971), .ZN(n682) );
  AOI22_X1 U500 ( .A1(data_in[5]), .A2(n830), .B1(n976), .B2(\mem[25][5] ), 
        .ZN(n971) );
  INV_X1 U501 ( .A(n970), .ZN(n681) );
  AOI22_X1 U502 ( .A1(data_in[6]), .A2(n830), .B1(n976), .B2(\mem[25][6] ), 
        .ZN(n970) );
  INV_X1 U503 ( .A(n969), .ZN(n680) );
  AOI22_X1 U504 ( .A1(data_in[7]), .A2(n830), .B1(n976), .B2(\mem[25][7] ), 
        .ZN(n969) );
  INV_X1 U505 ( .A(n968), .ZN(n679) );
  AOI22_X1 U506 ( .A1(data_in[0]), .A2(n829), .B1(n967), .B2(\mem[26][0] ), 
        .ZN(n968) );
  INV_X1 U507 ( .A(n966), .ZN(n678) );
  AOI22_X1 U508 ( .A1(data_in[1]), .A2(n829), .B1(n967), .B2(\mem[26][1] ), 
        .ZN(n966) );
  INV_X1 U509 ( .A(n965), .ZN(n677) );
  AOI22_X1 U510 ( .A1(data_in[2]), .A2(n829), .B1(n967), .B2(\mem[26][2] ), 
        .ZN(n965) );
  INV_X1 U511 ( .A(n964), .ZN(n676) );
  AOI22_X1 U512 ( .A1(data_in[3]), .A2(n829), .B1(n967), .B2(\mem[26][3] ), 
        .ZN(n964) );
  INV_X1 U513 ( .A(n963), .ZN(n675) );
  AOI22_X1 U514 ( .A1(data_in[4]), .A2(n829), .B1(n967), .B2(\mem[26][4] ), 
        .ZN(n963) );
  INV_X1 U515 ( .A(n962), .ZN(n674) );
  AOI22_X1 U516 ( .A1(data_in[5]), .A2(n829), .B1(n967), .B2(\mem[26][5] ), 
        .ZN(n962) );
  INV_X1 U517 ( .A(n961), .ZN(n673) );
  AOI22_X1 U518 ( .A1(data_in[6]), .A2(n829), .B1(n967), .B2(\mem[26][6] ), 
        .ZN(n961) );
  INV_X1 U519 ( .A(n960), .ZN(n672) );
  AOI22_X1 U520 ( .A1(data_in[7]), .A2(n829), .B1(n967), .B2(\mem[26][7] ), 
        .ZN(n960) );
  INV_X1 U521 ( .A(n959), .ZN(n671) );
  AOI22_X1 U522 ( .A1(data_in[0]), .A2(n828), .B1(n958), .B2(\mem[27][0] ), 
        .ZN(n959) );
  INV_X1 U523 ( .A(n957), .ZN(n670) );
  AOI22_X1 U524 ( .A1(data_in[1]), .A2(n828), .B1(n958), .B2(\mem[27][1] ), 
        .ZN(n957) );
  INV_X1 U525 ( .A(n956), .ZN(n669) );
  AOI22_X1 U526 ( .A1(data_in[2]), .A2(n828), .B1(n958), .B2(\mem[27][2] ), 
        .ZN(n956) );
  INV_X1 U527 ( .A(n955), .ZN(n668) );
  AOI22_X1 U528 ( .A1(data_in[3]), .A2(n828), .B1(n958), .B2(\mem[27][3] ), 
        .ZN(n955) );
  INV_X1 U529 ( .A(n954), .ZN(n667) );
  AOI22_X1 U530 ( .A1(data_in[4]), .A2(n828), .B1(n958), .B2(\mem[27][4] ), 
        .ZN(n954) );
  INV_X1 U531 ( .A(n953), .ZN(n666) );
  AOI22_X1 U532 ( .A1(data_in[5]), .A2(n828), .B1(n958), .B2(\mem[27][5] ), 
        .ZN(n953) );
  INV_X1 U533 ( .A(n952), .ZN(n665) );
  AOI22_X1 U534 ( .A1(data_in[6]), .A2(n828), .B1(n958), .B2(\mem[27][6] ), 
        .ZN(n952) );
  INV_X1 U535 ( .A(n951), .ZN(n664) );
  AOI22_X1 U536 ( .A1(data_in[7]), .A2(n828), .B1(n958), .B2(\mem[27][7] ), 
        .ZN(n951) );
  INV_X1 U537 ( .A(n950), .ZN(n663) );
  AOI22_X1 U538 ( .A1(data_in[0]), .A2(n827), .B1(n949), .B2(\mem[28][0] ), 
        .ZN(n950) );
  INV_X1 U539 ( .A(n948), .ZN(n662) );
  AOI22_X1 U540 ( .A1(data_in[1]), .A2(n827), .B1(n949), .B2(\mem[28][1] ), 
        .ZN(n948) );
  INV_X1 U541 ( .A(n947), .ZN(n661) );
  AOI22_X1 U542 ( .A1(data_in[2]), .A2(n827), .B1(n949), .B2(\mem[28][2] ), 
        .ZN(n947) );
  INV_X1 U543 ( .A(n946), .ZN(n660) );
  AOI22_X1 U544 ( .A1(data_in[3]), .A2(n827), .B1(n949), .B2(\mem[28][3] ), 
        .ZN(n946) );
  INV_X1 U545 ( .A(n945), .ZN(n659) );
  AOI22_X1 U546 ( .A1(data_in[4]), .A2(n827), .B1(n949), .B2(\mem[28][4] ), 
        .ZN(n945) );
  INV_X1 U547 ( .A(n944), .ZN(n658) );
  AOI22_X1 U548 ( .A1(data_in[5]), .A2(n827), .B1(n949), .B2(\mem[28][5] ), 
        .ZN(n944) );
  INV_X1 U549 ( .A(n943), .ZN(n657) );
  AOI22_X1 U550 ( .A1(data_in[6]), .A2(n827), .B1(n949), .B2(\mem[28][6] ), 
        .ZN(n943) );
  INV_X1 U551 ( .A(n942), .ZN(n656) );
  AOI22_X1 U552 ( .A1(data_in[7]), .A2(n827), .B1(n949), .B2(\mem[28][7] ), 
        .ZN(n942) );
  INV_X1 U553 ( .A(n941), .ZN(n655) );
  AOI22_X1 U554 ( .A1(data_in[0]), .A2(n826), .B1(n940), .B2(\mem[29][0] ), 
        .ZN(n941) );
  INV_X1 U555 ( .A(n939), .ZN(n654) );
  AOI22_X1 U556 ( .A1(data_in[1]), .A2(n826), .B1(n940), .B2(\mem[29][1] ), 
        .ZN(n939) );
  INV_X1 U557 ( .A(n938), .ZN(n653) );
  AOI22_X1 U558 ( .A1(data_in[2]), .A2(n826), .B1(n940), .B2(\mem[29][2] ), 
        .ZN(n938) );
  INV_X1 U559 ( .A(n937), .ZN(n652) );
  AOI22_X1 U560 ( .A1(data_in[3]), .A2(n826), .B1(n940), .B2(\mem[29][3] ), 
        .ZN(n937) );
  INV_X1 U561 ( .A(n936), .ZN(n651) );
  AOI22_X1 U562 ( .A1(data_in[4]), .A2(n826), .B1(n940), .B2(\mem[29][4] ), 
        .ZN(n936) );
  INV_X1 U563 ( .A(n935), .ZN(n650) );
  AOI22_X1 U564 ( .A1(data_in[5]), .A2(n826), .B1(n940), .B2(\mem[29][5] ), 
        .ZN(n935) );
  INV_X1 U565 ( .A(n934), .ZN(n649) );
  AOI22_X1 U566 ( .A1(data_in[6]), .A2(n826), .B1(n940), .B2(\mem[29][6] ), 
        .ZN(n934) );
  INV_X1 U567 ( .A(n933), .ZN(n648) );
  AOI22_X1 U568 ( .A1(data_in[7]), .A2(n826), .B1(n940), .B2(\mem[29][7] ), 
        .ZN(n933) );
  INV_X1 U569 ( .A(n932), .ZN(n647) );
  AOI22_X1 U570 ( .A1(data_in[0]), .A2(n825), .B1(n931), .B2(\mem[30][0] ), 
        .ZN(n932) );
  INV_X1 U571 ( .A(n930), .ZN(n646) );
  AOI22_X1 U572 ( .A1(data_in[1]), .A2(n825), .B1(n931), .B2(\mem[30][1] ), 
        .ZN(n930) );
  INV_X1 U573 ( .A(n929), .ZN(n645) );
  AOI22_X1 U574 ( .A1(data_in[2]), .A2(n825), .B1(n931), .B2(\mem[30][2] ), 
        .ZN(n929) );
  INV_X1 U575 ( .A(n928), .ZN(n644) );
  AOI22_X1 U576 ( .A1(data_in[3]), .A2(n825), .B1(n931), .B2(\mem[30][3] ), 
        .ZN(n928) );
  INV_X1 U577 ( .A(n927), .ZN(n643) );
  AOI22_X1 U578 ( .A1(data_in[4]), .A2(n825), .B1(n931), .B2(\mem[30][4] ), 
        .ZN(n927) );
  INV_X1 U579 ( .A(n926), .ZN(n642) );
  AOI22_X1 U580 ( .A1(data_in[5]), .A2(n825), .B1(n931), .B2(\mem[30][5] ), 
        .ZN(n926) );
  INV_X1 U581 ( .A(n925), .ZN(n641) );
  AOI22_X1 U582 ( .A1(data_in[6]), .A2(n825), .B1(n931), .B2(\mem[30][6] ), 
        .ZN(n925) );
  INV_X1 U583 ( .A(n924), .ZN(n640) );
  AOI22_X1 U584 ( .A1(data_in[7]), .A2(n825), .B1(n931), .B2(\mem[30][7] ), 
        .ZN(n924) );
  INV_X1 U585 ( .A(n923), .ZN(n639) );
  AOI22_X1 U586 ( .A1(data_in[0]), .A2(n824), .B1(n922), .B2(\mem[31][0] ), 
        .ZN(n923) );
  INV_X1 U587 ( .A(n921), .ZN(n638) );
  AOI22_X1 U588 ( .A1(data_in[1]), .A2(n824), .B1(n922), .B2(\mem[31][1] ), 
        .ZN(n921) );
  INV_X1 U589 ( .A(n920), .ZN(n637) );
  AOI22_X1 U590 ( .A1(data_in[2]), .A2(n824), .B1(n922), .B2(\mem[31][2] ), 
        .ZN(n920) );
  INV_X1 U591 ( .A(n919), .ZN(n636) );
  AOI22_X1 U592 ( .A1(data_in[3]), .A2(n824), .B1(n922), .B2(\mem[31][3] ), 
        .ZN(n919) );
  INV_X1 U593 ( .A(n918), .ZN(n635) );
  AOI22_X1 U594 ( .A1(data_in[4]), .A2(n824), .B1(n922), .B2(\mem[31][4] ), 
        .ZN(n918) );
  INV_X1 U595 ( .A(n917), .ZN(n634) );
  AOI22_X1 U596 ( .A1(data_in[5]), .A2(n824), .B1(n922), .B2(\mem[31][5] ), 
        .ZN(n917) );
  INV_X1 U597 ( .A(n916), .ZN(n633) );
  AOI22_X1 U598 ( .A1(data_in[6]), .A2(n824), .B1(n922), .B2(\mem[31][6] ), 
        .ZN(n916) );
  INV_X1 U599 ( .A(n915), .ZN(n632) );
  AOI22_X1 U600 ( .A1(data_in[7]), .A2(n824), .B1(n922), .B2(\mem[31][7] ), 
        .ZN(n915) );
  MUX2_X1 U601 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n612), .Z(n2) );
  MUX2_X1 U602 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n612), .Z(n3) );
  MUX2_X1 U603 ( .A(n3), .B(n2), .S(n609), .Z(n4) );
  MUX2_X1 U604 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n612), .Z(n5) );
  MUX2_X1 U605 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n612), .Z(n6) );
  MUX2_X1 U606 ( .A(n6), .B(n5), .S(n609), .Z(n7) );
  MUX2_X1 U607 ( .A(n7), .B(n4), .S(N12), .Z(n8) );
  MUX2_X1 U608 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n612), .Z(n9) );
  MUX2_X1 U609 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n612), .Z(n10) );
  MUX2_X1 U610 ( .A(n10), .B(n9), .S(n609), .Z(n11) );
  MUX2_X1 U611 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n612), .Z(n12) );
  MUX2_X1 U612 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n612), .Z(n13) );
  MUX2_X1 U613 ( .A(n13), .B(n12), .S(n609), .Z(n14) );
  MUX2_X1 U614 ( .A(n14), .B(n11), .S(n607), .Z(n15) );
  MUX2_X1 U615 ( .A(n15), .B(n8), .S(N13), .Z(n16) );
  MUX2_X1 U616 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n613), .Z(n17) );
  MUX2_X1 U617 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n613), .Z(n18) );
  MUX2_X1 U618 ( .A(n18), .B(n17), .S(n610), .Z(n19) );
  MUX2_X1 U619 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n613), .Z(n20) );
  MUX2_X1 U620 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n613), .Z(n21) );
  MUX2_X1 U621 ( .A(n21), .B(n20), .S(n610), .Z(n22) );
  MUX2_X1 U622 ( .A(n22), .B(n19), .S(n608), .Z(n23) );
  MUX2_X1 U623 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n613), .Z(n24) );
  MUX2_X1 U624 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n613), .Z(n25) );
  MUX2_X1 U625 ( .A(n25), .B(n24), .S(n610), .Z(n26) );
  MUX2_X1 U626 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n613), .Z(n27) );
  MUX2_X1 U627 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n613), .Z(n28) );
  MUX2_X1 U628 ( .A(n28), .B(n27), .S(n610), .Z(n29) );
  MUX2_X1 U629 ( .A(n29), .B(n26), .S(n608), .Z(n30) );
  MUX2_X1 U630 ( .A(n30), .B(n23), .S(N13), .Z(n31) );
  MUX2_X1 U631 ( .A(n31), .B(n16), .S(N14), .Z(N22) );
  MUX2_X1 U632 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n613), .Z(n32) );
  MUX2_X1 U633 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n613), .Z(n33) );
  MUX2_X1 U634 ( .A(n33), .B(n32), .S(n610), .Z(n34) );
  MUX2_X1 U635 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n613), .Z(n35) );
  MUX2_X1 U636 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n613), .Z(n36) );
  MUX2_X1 U637 ( .A(n36), .B(n35), .S(n610), .Z(n37) );
  MUX2_X1 U638 ( .A(n37), .B(n34), .S(N12), .Z(n38) );
  MUX2_X1 U639 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n614), .Z(n39) );
  MUX2_X1 U640 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n614), .Z(n40) );
  MUX2_X1 U641 ( .A(n40), .B(n39), .S(n610), .Z(n41) );
  MUX2_X1 U642 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n614), .Z(n42) );
  MUX2_X1 U643 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n614), .Z(n43) );
  MUX2_X1 U644 ( .A(n43), .B(n42), .S(n610), .Z(n44) );
  MUX2_X1 U645 ( .A(n44), .B(n41), .S(n608), .Z(n45) );
  MUX2_X1 U646 ( .A(n45), .B(n38), .S(N13), .Z(n46) );
  MUX2_X1 U647 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n614), .Z(n47) );
  MUX2_X1 U648 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n614), .Z(n48) );
  MUX2_X1 U649 ( .A(n48), .B(n47), .S(n610), .Z(n49) );
  MUX2_X1 U650 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n614), .Z(n50) );
  MUX2_X1 U651 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n614), .Z(n51) );
  MUX2_X1 U652 ( .A(n51), .B(n50), .S(n610), .Z(n52) );
  MUX2_X1 U653 ( .A(n52), .B(n49), .S(n607), .Z(n53) );
  MUX2_X1 U654 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n614), .Z(n54) );
  MUX2_X1 U655 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n614), .Z(n55) );
  MUX2_X1 U656 ( .A(n55), .B(n54), .S(n610), .Z(n56) );
  MUX2_X1 U657 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n614), .Z(n57) );
  MUX2_X1 U658 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n614), .Z(n58) );
  MUX2_X1 U659 ( .A(n58), .B(n57), .S(n610), .Z(n59) );
  MUX2_X1 U660 ( .A(n59), .B(n56), .S(N12), .Z(n60) );
  MUX2_X1 U661 ( .A(n60), .B(n53), .S(N13), .Z(n61) );
  MUX2_X1 U662 ( .A(n61), .B(n46), .S(N14), .Z(N21) );
  MUX2_X1 U663 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n615), .Z(n62) );
  MUX2_X1 U664 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n615), .Z(n63) );
  MUX2_X1 U665 ( .A(n63), .B(n62), .S(n611), .Z(n64) );
  MUX2_X1 U666 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n615), .Z(n65) );
  MUX2_X1 U667 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n615), .Z(n66) );
  MUX2_X1 U668 ( .A(n66), .B(n65), .S(n611), .Z(n67) );
  MUX2_X1 U669 ( .A(n67), .B(n64), .S(n607), .Z(n68) );
  MUX2_X1 U670 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n615), .Z(n69) );
  MUX2_X1 U671 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n615), .Z(n70) );
  MUX2_X1 U672 ( .A(n70), .B(n69), .S(n611), .Z(n71) );
  MUX2_X1 U673 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n615), .Z(n72) );
  MUX2_X1 U674 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n615), .Z(n73) );
  MUX2_X1 U675 ( .A(n73), .B(n72), .S(n611), .Z(n74) );
  MUX2_X1 U676 ( .A(n74), .B(n71), .S(n607), .Z(n75) );
  MUX2_X1 U677 ( .A(n75), .B(n68), .S(N13), .Z(n76) );
  MUX2_X1 U678 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n615), .Z(n77) );
  MUX2_X1 U679 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n615), .Z(n78) );
  MUX2_X1 U680 ( .A(n78), .B(n77), .S(n611), .Z(n79) );
  MUX2_X1 U681 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n615), .Z(n80) );
  MUX2_X1 U682 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n615), .Z(n81) );
  MUX2_X1 U683 ( .A(n81), .B(n80), .S(n611), .Z(n82) );
  MUX2_X1 U684 ( .A(n82), .B(n79), .S(n607), .Z(n83) );
  MUX2_X1 U685 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n616), .Z(n84) );
  MUX2_X1 U686 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n616), .Z(n85) );
  MUX2_X1 U687 ( .A(n85), .B(n84), .S(n611), .Z(n86) );
  MUX2_X1 U688 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n616), .Z(n87) );
  MUX2_X1 U689 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n616), .Z(n88) );
  MUX2_X1 U690 ( .A(n88), .B(n87), .S(n611), .Z(n89) );
  MUX2_X1 U691 ( .A(n89), .B(n86), .S(n607), .Z(n90) );
  MUX2_X1 U692 ( .A(n90), .B(n83), .S(N13), .Z(n91) );
  MUX2_X1 U693 ( .A(n91), .B(n76), .S(N14), .Z(N20) );
  MUX2_X1 U694 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n616), .Z(n92) );
  MUX2_X1 U695 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n616), .Z(n93) );
  MUX2_X1 U696 ( .A(n93), .B(n92), .S(n611), .Z(n94) );
  MUX2_X1 U697 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n616), .Z(n95) );
  MUX2_X1 U698 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n616), .Z(n96) );
  MUX2_X1 U699 ( .A(n96), .B(n95), .S(n611), .Z(n97) );
  MUX2_X1 U700 ( .A(n97), .B(n94), .S(n607), .Z(n98) );
  MUX2_X1 U701 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n616), .Z(n99) );
  MUX2_X1 U702 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n616), .Z(n100) );
  MUX2_X1 U703 ( .A(n100), .B(n99), .S(n611), .Z(n101) );
  MUX2_X1 U704 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n616), .Z(n102) );
  MUX2_X1 U705 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n616), .Z(n103) );
  MUX2_X1 U706 ( .A(n103), .B(n102), .S(n611), .Z(n104) );
  MUX2_X1 U707 ( .A(n104), .B(n101), .S(n607), .Z(n105) );
  MUX2_X1 U708 ( .A(n105), .B(n98), .S(N13), .Z(n106) );
  MUX2_X1 U709 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n615), .Z(n107) );
  MUX2_X1 U710 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n621), .Z(n108) );
  MUX2_X1 U711 ( .A(n108), .B(n107), .S(n611), .Z(n109) );
  MUX2_X1 U712 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n620), .Z(n110) );
  MUX2_X1 U713 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n111) );
  MUX2_X1 U714 ( .A(n111), .B(n110), .S(n611), .Z(n112) );
  MUX2_X1 U715 ( .A(n112), .B(n109), .S(n607), .Z(n113) );
  MUX2_X1 U716 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n620), .Z(n114) );
  MUX2_X1 U717 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n620), .Z(n115) );
  MUX2_X1 U718 ( .A(n115), .B(n114), .S(n610), .Z(n116) );
  MUX2_X1 U719 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n621), .Z(n117) );
  MUX2_X1 U720 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n621), .Z(n118) );
  MUX2_X1 U721 ( .A(n118), .B(n117), .S(n610), .Z(n119) );
  MUX2_X1 U722 ( .A(n119), .B(n116), .S(n607), .Z(n120) );
  MUX2_X1 U723 ( .A(n120), .B(n113), .S(N13), .Z(n121) );
  MUX2_X1 U724 ( .A(n121), .B(n106), .S(N14), .Z(N19) );
  MUX2_X1 U725 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n612), .Z(n122) );
  MUX2_X1 U726 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n620), .Z(n123) );
  MUX2_X1 U727 ( .A(n123), .B(n122), .S(n610), .Z(n124) );
  MUX2_X1 U728 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n616), .Z(n125) );
  MUX2_X1 U729 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n620), .Z(n126) );
  MUX2_X1 U730 ( .A(n126), .B(n125), .S(N11), .Z(n127) );
  MUX2_X1 U731 ( .A(n127), .B(n124), .S(n607), .Z(n128) );
  MUX2_X1 U732 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n612), .Z(n129) );
  MUX2_X1 U733 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n621), .Z(n130) );
  MUX2_X1 U734 ( .A(n130), .B(n129), .S(n609), .Z(n131) );
  MUX2_X1 U735 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n621), .Z(n132) );
  MUX2_X1 U736 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(N10), .Z(n133) );
  MUX2_X1 U737 ( .A(n133), .B(n132), .S(n611), .Z(n134) );
  MUX2_X1 U738 ( .A(n134), .B(n131), .S(n607), .Z(n135) );
  MUX2_X1 U739 ( .A(n135), .B(n128), .S(N13), .Z(n136) );
  MUX2_X1 U740 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n612), .Z(n137) );
  MUX2_X1 U741 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n620), .Z(n138) );
  MUX2_X1 U742 ( .A(n138), .B(n137), .S(n610), .Z(n139) );
  MUX2_X1 U743 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n612), .Z(n140) );
  MUX2_X1 U744 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n141) );
  MUX2_X1 U745 ( .A(n141), .B(n140), .S(n610), .Z(n142) );
  MUX2_X1 U746 ( .A(n142), .B(n139), .S(n607), .Z(n143) );
  MUX2_X1 U747 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n612), .Z(n144) );
  MUX2_X1 U748 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n145) );
  MUX2_X1 U749 ( .A(n145), .B(n144), .S(n609), .Z(n146) );
  MUX2_X1 U750 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n620), .Z(n147) );
  MUX2_X1 U751 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n148) );
  MUX2_X1 U752 ( .A(n148), .B(n147), .S(n609), .Z(n149) );
  MUX2_X1 U753 ( .A(n149), .B(n146), .S(n607), .Z(n150) );
  MUX2_X1 U754 ( .A(n150), .B(n143), .S(N13), .Z(n151) );
  MUX2_X1 U755 ( .A(n151), .B(n136), .S(N14), .Z(N18) );
  MUX2_X1 U756 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n617), .Z(n152) );
  MUX2_X1 U757 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n617), .Z(n153) );
  MUX2_X1 U758 ( .A(n153), .B(n152), .S(n611), .Z(n154) );
  MUX2_X1 U759 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n617), .Z(n155) );
  MUX2_X1 U760 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n617), .Z(n156) );
  MUX2_X1 U761 ( .A(n156), .B(n155), .S(n611), .Z(n157) );
  MUX2_X1 U762 ( .A(n157), .B(n154), .S(n608), .Z(n158) );
  MUX2_X1 U763 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n617), .Z(n159) );
  MUX2_X1 U764 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n617), .Z(n160) );
  MUX2_X1 U765 ( .A(n160), .B(n159), .S(n609), .Z(n161) );
  MUX2_X1 U766 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n617), .Z(n162) );
  MUX2_X1 U767 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n617), .Z(n163) );
  MUX2_X1 U768 ( .A(n163), .B(n162), .S(N11), .Z(n164) );
  MUX2_X1 U769 ( .A(n164), .B(n161), .S(n608), .Z(n165) );
  MUX2_X1 U770 ( .A(n165), .B(n158), .S(N13), .Z(n166) );
  MUX2_X1 U771 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n617), .Z(n167) );
  MUX2_X1 U772 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n617), .Z(n168) );
  MUX2_X1 U773 ( .A(n168), .B(n167), .S(n610), .Z(n169) );
  MUX2_X1 U774 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n617), .Z(n170) );
  MUX2_X1 U775 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n617), .Z(n171) );
  MUX2_X1 U776 ( .A(n171), .B(n170), .S(n610), .Z(n172) );
  MUX2_X1 U777 ( .A(n172), .B(n169), .S(n608), .Z(n173) );
  MUX2_X1 U778 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n618), .Z(n174) );
  MUX2_X1 U779 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n618), .Z(n175) );
  MUX2_X1 U780 ( .A(n175), .B(n174), .S(N11), .Z(n176) );
  MUX2_X1 U781 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n618), .Z(n177) );
  MUX2_X1 U782 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n618), .Z(n178) );
  MUX2_X1 U783 ( .A(n178), .B(n177), .S(n611), .Z(n179) );
  MUX2_X1 U784 ( .A(n179), .B(n176), .S(n608), .Z(n180) );
  MUX2_X1 U785 ( .A(n180), .B(n173), .S(N13), .Z(n181) );
  MUX2_X1 U786 ( .A(n181), .B(n166), .S(N14), .Z(N17) );
  MUX2_X1 U787 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n618), .Z(n182) );
  MUX2_X1 U788 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n618), .Z(n183) );
  MUX2_X1 U789 ( .A(n183), .B(n182), .S(n609), .Z(n184) );
  MUX2_X1 U790 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n618), .Z(n185) );
  MUX2_X1 U791 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n618), .Z(n186) );
  MUX2_X1 U792 ( .A(n186), .B(n185), .S(N11), .Z(n187) );
  MUX2_X1 U793 ( .A(n187), .B(n184), .S(n608), .Z(n188) );
  MUX2_X1 U794 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n618), .Z(n189) );
  MUX2_X1 U795 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n618), .Z(n190) );
  MUX2_X1 U796 ( .A(n190), .B(n189), .S(n611), .Z(n191) );
  MUX2_X1 U797 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n618), .Z(n192) );
  MUX2_X1 U798 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n618), .Z(n193) );
  MUX2_X1 U799 ( .A(n193), .B(n192), .S(N11), .Z(n194) );
  MUX2_X1 U800 ( .A(n194), .B(n191), .S(n608), .Z(n195) );
  MUX2_X1 U801 ( .A(n195), .B(n188), .S(N13), .Z(n196) );
  MUX2_X1 U802 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n619), .Z(n197) );
  MUX2_X1 U803 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n619), .Z(n198) );
  MUX2_X1 U804 ( .A(n198), .B(n197), .S(n609), .Z(n199) );
  MUX2_X1 U805 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n619), .Z(n200) );
  MUX2_X1 U806 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n619), .Z(n201) );
  MUX2_X1 U807 ( .A(n201), .B(n200), .S(n611), .Z(n202) );
  MUX2_X1 U808 ( .A(n202), .B(n199), .S(n608), .Z(n203) );
  MUX2_X1 U809 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n619), .Z(n204) );
  MUX2_X1 U810 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n619), .Z(n205) );
  MUX2_X1 U811 ( .A(n205), .B(n204), .S(n609), .Z(n206) );
  MUX2_X1 U812 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n619), .Z(n207) );
  MUX2_X1 U813 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n619), .Z(n208) );
  MUX2_X1 U814 ( .A(n208), .B(n207), .S(n610), .Z(n209) );
  MUX2_X1 U815 ( .A(n209), .B(n206), .S(n608), .Z(n210) );
  MUX2_X1 U816 ( .A(n210), .B(n203), .S(N13), .Z(n211) );
  MUX2_X1 U817 ( .A(n211), .B(n196), .S(N14), .Z(N16) );
  MUX2_X1 U818 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n619), .Z(n212) );
  MUX2_X1 U819 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n619), .Z(n213) );
  MUX2_X1 U820 ( .A(n213), .B(n212), .S(n609), .Z(n214) );
  MUX2_X1 U821 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n619), .Z(n215) );
  MUX2_X1 U822 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n619), .Z(n216) );
  MUX2_X1 U823 ( .A(n216), .B(n215), .S(n609), .Z(n217) );
  MUX2_X1 U824 ( .A(n217), .B(n214), .S(n608), .Z(n218) );
  MUX2_X1 U825 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n614), .Z(n219) );
  MUX2_X1 U826 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n621), .Z(n220) );
  MUX2_X1 U827 ( .A(n220), .B(n219), .S(n609), .Z(n221) );
  MUX2_X1 U828 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n621), .Z(n222) );
  MUX2_X1 U829 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n621), .Z(n223) );
  MUX2_X1 U830 ( .A(n223), .B(n222), .S(n611), .Z(n224) );
  MUX2_X1 U831 ( .A(n224), .B(n221), .S(n608), .Z(n225) );
  MUX2_X1 U832 ( .A(n225), .B(n218), .S(N13), .Z(n226) );
  MUX2_X1 U833 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n621), .Z(n227) );
  MUX2_X1 U834 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n620), .Z(n228) );
  MUX2_X1 U835 ( .A(n228), .B(n227), .S(n609), .Z(n229) );
  MUX2_X1 U836 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n613), .Z(n595) );
  MUX2_X1 U837 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n621), .Z(n596) );
  MUX2_X1 U838 ( .A(n596), .B(n595), .S(n609), .Z(n597) );
  MUX2_X1 U839 ( .A(n597), .B(n229), .S(n608), .Z(n598) );
  MUX2_X1 U840 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n621), .Z(n599) );
  MUX2_X1 U841 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n620), .Z(n600) );
  MUX2_X1 U842 ( .A(n600), .B(n599), .S(n609), .Z(n601) );
  MUX2_X1 U843 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n620), .Z(n602) );
  MUX2_X1 U844 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n620), .Z(n603) );
  MUX2_X1 U845 ( .A(n603), .B(n602), .S(n609), .Z(n604) );
  MUX2_X1 U846 ( .A(n604), .B(n601), .S(n608), .Z(n605) );
  MUX2_X1 U847 ( .A(n605), .B(n598), .S(N13), .Z(n606) );
  MUX2_X1 U848 ( .A(n606), .B(n226), .S(N14), .Z(N15) );
  CLKBUF_X1 U849 ( .A(N11), .Z(n609) );
  INV_X1 U850 ( .A(N10), .ZN(n622) );
  INV_X1 U851 ( .A(N11), .ZN(n623) );
  INV_X1 U852 ( .A(data_in[0]), .ZN(n624) );
  INV_X1 U853 ( .A(data_in[1]), .ZN(n625) );
  INV_X1 U854 ( .A(data_in[2]), .ZN(n626) );
  INV_X1 U855 ( .A(data_in[3]), .ZN(n627) );
  INV_X1 U856 ( .A(data_in[4]), .ZN(n628) );
  INV_X1 U857 ( .A(data_in[5]), .ZN(n629) );
  INV_X1 U858 ( .A(data_in[6]), .ZN(n630) );
  INV_X1 U859 ( .A(data_in[7]), .ZN(n631) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_11 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n628), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n629), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n630), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n631), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n632), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n633), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n634), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n635), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n636), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n637), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n638), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n639), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n640), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n641), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n642), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n643), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n644), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n645), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n646), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n647), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n648), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n649), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n650), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n651), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n652), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n653), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n654), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n655), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n656), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n657), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n658), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n659), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n660), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n661), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n662), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n663), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n664), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n665), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n666), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n667), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n668), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n669), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n670), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n671), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n672), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n673), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n674), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n675), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n676), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n677), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n678), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n679), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n680), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n681), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n682), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n683), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n684), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n685), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n686), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n687), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n688), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n689), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n690), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n691), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n692), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n693), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n694), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n695), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n696), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n697), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n698), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n699), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n700), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n701), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n702), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n703), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n704), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n705), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n706), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n707), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n708), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n709), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n710), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n711), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n712), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n713), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n714), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n715), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n716), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n717), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n718), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n719), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n720), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n721), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n722), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n723), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n724), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n725), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n726), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n727), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n728), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n729), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n730), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n731), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n732), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n733), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n734), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n735), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n736), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n737), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n738), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n739), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n740), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n741), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n742), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n743), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n744), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n745), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n746), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n747), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n748), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n749), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n750), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n751), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n752), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n753), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n754), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n755), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n756), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n757), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n758), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n759), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n760), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n761), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n762), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n763), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n764), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n765), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n766), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n767), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n768), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n769), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n770), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n771), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n772), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n773), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n774), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n775), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n776), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n777), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n778), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n779), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n780), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n781), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n782), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n783), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n784), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n785), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n786), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n787), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n788), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n789), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n790), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n791), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n792), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n793), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n794), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n795), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n796), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n797), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n798), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n799), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n800), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n801), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n802), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n803), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n804), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n805), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n806), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n807), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n808), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n809), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n810), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n811), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n812), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n813), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n814), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n815), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n816), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n817), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n818), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n819), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n847), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n848), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n849), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n850), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n851), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n852), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n853), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n854), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n855), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n856), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n857), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n858), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n859), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n860), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n861), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n862), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n863), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n864), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n865), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n866), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n867), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n868), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n869), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n870), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n871), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n872), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n873), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n874), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n875), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n876), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n877), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n878), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n879), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n880), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n881), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n882), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n883), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n884), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n885), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n886), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n887), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n888), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n889), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n890), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n891), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n892), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n893), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n894), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n895), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n896), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n897), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n898), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n899), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n900), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n901), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n902), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n903), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n904), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n905), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n906), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n907), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n908), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n909), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n910), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  CLKBUF_X1 U3 ( .A(N10), .Z(n617) );
  BUF_X1 U4 ( .A(N10), .Z(n611) );
  BUF_X1 U5 ( .A(n617), .Z(n616) );
  BUF_X1 U6 ( .A(N10), .Z(n613) );
  BUF_X1 U7 ( .A(N10), .Z(n612) );
  BUF_X1 U8 ( .A(N10), .Z(n614) );
  BUF_X1 U9 ( .A(n617), .Z(n615) );
  BUF_X1 U10 ( .A(N11), .Z(n609) );
  BUF_X1 U11 ( .A(N11), .Z(n610) );
  NOR3_X1 U12 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1202) );
  NOR3_X1 U13 ( .A1(N11), .A2(N12), .A3(n618), .ZN(n1191) );
  NOR3_X1 U14 ( .A1(N10), .A2(N12), .A3(n619), .ZN(n1181) );
  NOR3_X1 U15 ( .A1(n618), .A2(N12), .A3(n619), .ZN(n1171) );
  INV_X1 U16 ( .A(n1128), .ZN(n843) );
  INV_X1 U17 ( .A(n1118), .ZN(n842) );
  INV_X1 U18 ( .A(n1109), .ZN(n841) );
  INV_X1 U19 ( .A(n1100), .ZN(n840) );
  INV_X1 U20 ( .A(n1055), .ZN(n835) );
  INV_X1 U21 ( .A(n1045), .ZN(n834) );
  INV_X1 U22 ( .A(n1036), .ZN(n833) );
  INV_X1 U23 ( .A(n1027), .ZN(n832) );
  INV_X1 U24 ( .A(n982), .ZN(n827) );
  INV_X1 U25 ( .A(n972), .ZN(n826) );
  INV_X1 U26 ( .A(n963), .ZN(n825) );
  INV_X1 U27 ( .A(n954), .ZN(n824) );
  INV_X1 U28 ( .A(n945), .ZN(n823) );
  INV_X1 U29 ( .A(n936), .ZN(n822) );
  INV_X1 U30 ( .A(n927), .ZN(n821) );
  INV_X1 U31 ( .A(n918), .ZN(n820) );
  INV_X1 U32 ( .A(n1091), .ZN(n839) );
  INV_X1 U33 ( .A(n1082), .ZN(n838) );
  INV_X1 U34 ( .A(n1073), .ZN(n837) );
  INV_X1 U35 ( .A(n1064), .ZN(n836) );
  INV_X1 U36 ( .A(n1018), .ZN(n831) );
  INV_X1 U37 ( .A(n1009), .ZN(n830) );
  INV_X1 U38 ( .A(n1000), .ZN(n829) );
  INV_X1 U39 ( .A(n991), .ZN(n828) );
  BUF_X1 U40 ( .A(N12), .Z(n607) );
  INV_X1 U41 ( .A(N13), .ZN(n845) );
  AND3_X1 U42 ( .A1(n618), .A2(n619), .A3(N12), .ZN(n1161) );
  AND3_X1 U43 ( .A1(N10), .A2(n619), .A3(N12), .ZN(n1151) );
  AND3_X1 U44 ( .A1(N11), .A2(n618), .A3(N12), .ZN(n1141) );
  AND3_X1 U45 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1131) );
  BUF_X1 U46 ( .A(N12), .Z(n606) );
  INV_X1 U47 ( .A(N14), .ZN(n846) );
  NAND2_X1 U48 ( .A1(n1191), .A2(n1201), .ZN(n1200) );
  NAND2_X1 U49 ( .A1(n1181), .A2(n1201), .ZN(n1190) );
  NAND2_X1 U50 ( .A1(n1171), .A2(n1201), .ZN(n1180) );
  NAND2_X1 U51 ( .A1(n1161), .A2(n1201), .ZN(n1170) );
  NAND2_X1 U52 ( .A1(n1151), .A2(n1201), .ZN(n1160) );
  NAND2_X1 U53 ( .A1(n1141), .A2(n1201), .ZN(n1150) );
  NAND2_X1 U54 ( .A1(n1131), .A2(n1201), .ZN(n1140) );
  NAND2_X1 U55 ( .A1(n1202), .A2(n1201), .ZN(n1211) );
  NAND2_X1 U56 ( .A1(n1120), .A2(n1202), .ZN(n1128) );
  NAND2_X1 U57 ( .A1(n1120), .A2(n1191), .ZN(n1118) );
  NAND2_X1 U58 ( .A1(n1120), .A2(n1181), .ZN(n1109) );
  NAND2_X1 U59 ( .A1(n1120), .A2(n1171), .ZN(n1100) );
  NAND2_X1 U60 ( .A1(n1047), .A2(n1202), .ZN(n1055) );
  NAND2_X1 U61 ( .A1(n1047), .A2(n1191), .ZN(n1045) );
  NAND2_X1 U62 ( .A1(n1047), .A2(n1181), .ZN(n1036) );
  NAND2_X1 U63 ( .A1(n1047), .A2(n1171), .ZN(n1027) );
  NAND2_X1 U64 ( .A1(n974), .A2(n1202), .ZN(n982) );
  NAND2_X1 U65 ( .A1(n974), .A2(n1191), .ZN(n972) );
  NAND2_X1 U66 ( .A1(n974), .A2(n1181), .ZN(n963) );
  NAND2_X1 U67 ( .A1(n974), .A2(n1171), .ZN(n954) );
  NAND2_X1 U68 ( .A1(n1120), .A2(n1161), .ZN(n1091) );
  NAND2_X1 U69 ( .A1(n1120), .A2(n1151), .ZN(n1082) );
  NAND2_X1 U70 ( .A1(n1120), .A2(n1141), .ZN(n1073) );
  NAND2_X1 U71 ( .A1(n1120), .A2(n1131), .ZN(n1064) );
  NAND2_X1 U72 ( .A1(n1047), .A2(n1161), .ZN(n1018) );
  NAND2_X1 U73 ( .A1(n1047), .A2(n1151), .ZN(n1009) );
  NAND2_X1 U74 ( .A1(n1047), .A2(n1141), .ZN(n1000) );
  NAND2_X1 U75 ( .A1(n1047), .A2(n1131), .ZN(n991) );
  NAND2_X1 U76 ( .A1(n974), .A2(n1161), .ZN(n945) );
  NAND2_X1 U77 ( .A1(n974), .A2(n1151), .ZN(n936) );
  NAND2_X1 U78 ( .A1(n974), .A2(n1141), .ZN(n927) );
  NAND2_X1 U79 ( .A1(n974), .A2(n1131), .ZN(n918) );
  AND3_X1 U80 ( .A1(n845), .A2(n846), .A3(n1130), .ZN(n1201) );
  AND3_X1 U81 ( .A1(N13), .A2(n1130), .A3(N14), .ZN(n974) );
  AND3_X1 U82 ( .A1(n1130), .A2(n846), .A3(N13), .ZN(n1120) );
  AND3_X1 U83 ( .A1(n1130), .A2(n845), .A3(N14), .ZN(n1047) );
  NOR2_X1 U84 ( .A1(n844), .A2(addr[5]), .ZN(n1130) );
  INV_X1 U85 ( .A(wr_en), .ZN(n844) );
  OAI21_X1 U86 ( .B1(n620), .B2(n1170), .A(n1169), .ZN(n878) );
  NAND2_X1 U87 ( .A1(\mem[4][0] ), .A2(n1170), .ZN(n1169) );
  OAI21_X1 U88 ( .B1(n621), .B2(n1170), .A(n1168), .ZN(n877) );
  NAND2_X1 U89 ( .A1(\mem[4][1] ), .A2(n1170), .ZN(n1168) );
  OAI21_X1 U90 ( .B1(n622), .B2(n1170), .A(n1167), .ZN(n876) );
  NAND2_X1 U91 ( .A1(\mem[4][2] ), .A2(n1170), .ZN(n1167) );
  OAI21_X1 U92 ( .B1(n623), .B2(n1170), .A(n1166), .ZN(n875) );
  NAND2_X1 U93 ( .A1(\mem[4][3] ), .A2(n1170), .ZN(n1166) );
  OAI21_X1 U94 ( .B1(n624), .B2(n1170), .A(n1165), .ZN(n874) );
  NAND2_X1 U95 ( .A1(\mem[4][4] ), .A2(n1170), .ZN(n1165) );
  OAI21_X1 U96 ( .B1(n625), .B2(n1170), .A(n1164), .ZN(n873) );
  NAND2_X1 U97 ( .A1(\mem[4][5] ), .A2(n1170), .ZN(n1164) );
  OAI21_X1 U98 ( .B1(n626), .B2(n1170), .A(n1163), .ZN(n872) );
  NAND2_X1 U99 ( .A1(\mem[4][6] ), .A2(n1170), .ZN(n1163) );
  OAI21_X1 U100 ( .B1(n627), .B2(n1170), .A(n1162), .ZN(n871) );
  NAND2_X1 U101 ( .A1(\mem[4][7] ), .A2(n1170), .ZN(n1162) );
  OAI21_X1 U102 ( .B1(n620), .B2(n1150), .A(n1149), .ZN(n862) );
  NAND2_X1 U103 ( .A1(\mem[6][0] ), .A2(n1150), .ZN(n1149) );
  OAI21_X1 U104 ( .B1(n621), .B2(n1150), .A(n1148), .ZN(n861) );
  NAND2_X1 U105 ( .A1(\mem[6][1] ), .A2(n1150), .ZN(n1148) );
  OAI21_X1 U106 ( .B1(n622), .B2(n1150), .A(n1147), .ZN(n860) );
  NAND2_X1 U107 ( .A1(\mem[6][2] ), .A2(n1150), .ZN(n1147) );
  OAI21_X1 U108 ( .B1(n623), .B2(n1150), .A(n1146), .ZN(n859) );
  NAND2_X1 U109 ( .A1(\mem[6][3] ), .A2(n1150), .ZN(n1146) );
  OAI21_X1 U110 ( .B1(n624), .B2(n1150), .A(n1145), .ZN(n858) );
  NAND2_X1 U111 ( .A1(\mem[6][4] ), .A2(n1150), .ZN(n1145) );
  OAI21_X1 U112 ( .B1(n625), .B2(n1150), .A(n1144), .ZN(n857) );
  NAND2_X1 U113 ( .A1(\mem[6][5] ), .A2(n1150), .ZN(n1144) );
  OAI21_X1 U114 ( .B1(n626), .B2(n1150), .A(n1143), .ZN(n856) );
  NAND2_X1 U115 ( .A1(\mem[6][6] ), .A2(n1150), .ZN(n1143) );
  OAI21_X1 U116 ( .B1(n627), .B2(n1150), .A(n1142), .ZN(n855) );
  NAND2_X1 U117 ( .A1(\mem[6][7] ), .A2(n1150), .ZN(n1142) );
  OAI21_X1 U118 ( .B1(n620), .B2(n1140), .A(n1139), .ZN(n854) );
  NAND2_X1 U119 ( .A1(\mem[7][0] ), .A2(n1140), .ZN(n1139) );
  OAI21_X1 U120 ( .B1(n621), .B2(n1140), .A(n1138), .ZN(n853) );
  NAND2_X1 U121 ( .A1(\mem[7][1] ), .A2(n1140), .ZN(n1138) );
  OAI21_X1 U122 ( .B1(n622), .B2(n1140), .A(n1137), .ZN(n852) );
  NAND2_X1 U123 ( .A1(\mem[7][2] ), .A2(n1140), .ZN(n1137) );
  OAI21_X1 U124 ( .B1(n623), .B2(n1140), .A(n1136), .ZN(n851) );
  NAND2_X1 U125 ( .A1(\mem[7][3] ), .A2(n1140), .ZN(n1136) );
  OAI21_X1 U126 ( .B1(n624), .B2(n1140), .A(n1135), .ZN(n850) );
  NAND2_X1 U127 ( .A1(\mem[7][4] ), .A2(n1140), .ZN(n1135) );
  OAI21_X1 U128 ( .B1(n625), .B2(n1140), .A(n1134), .ZN(n849) );
  NAND2_X1 U129 ( .A1(\mem[7][5] ), .A2(n1140), .ZN(n1134) );
  OAI21_X1 U130 ( .B1(n626), .B2(n1140), .A(n1133), .ZN(n848) );
  NAND2_X1 U131 ( .A1(\mem[7][6] ), .A2(n1140), .ZN(n1133) );
  OAI21_X1 U132 ( .B1(n627), .B2(n1140), .A(n1132), .ZN(n847) );
  NAND2_X1 U133 ( .A1(\mem[7][7] ), .A2(n1140), .ZN(n1132) );
  OAI21_X1 U134 ( .B1(n620), .B2(n1200), .A(n1199), .ZN(n902) );
  NAND2_X1 U135 ( .A1(\mem[1][0] ), .A2(n1200), .ZN(n1199) );
  OAI21_X1 U136 ( .B1(n621), .B2(n1200), .A(n1198), .ZN(n901) );
  NAND2_X1 U137 ( .A1(\mem[1][1] ), .A2(n1200), .ZN(n1198) );
  OAI21_X1 U138 ( .B1(n622), .B2(n1200), .A(n1197), .ZN(n900) );
  NAND2_X1 U139 ( .A1(\mem[1][2] ), .A2(n1200), .ZN(n1197) );
  OAI21_X1 U140 ( .B1(n623), .B2(n1200), .A(n1196), .ZN(n899) );
  NAND2_X1 U141 ( .A1(\mem[1][3] ), .A2(n1200), .ZN(n1196) );
  OAI21_X1 U142 ( .B1(n624), .B2(n1200), .A(n1195), .ZN(n898) );
  NAND2_X1 U143 ( .A1(\mem[1][4] ), .A2(n1200), .ZN(n1195) );
  OAI21_X1 U144 ( .B1(n625), .B2(n1200), .A(n1194), .ZN(n897) );
  NAND2_X1 U145 ( .A1(\mem[1][5] ), .A2(n1200), .ZN(n1194) );
  OAI21_X1 U146 ( .B1(n626), .B2(n1200), .A(n1193), .ZN(n896) );
  NAND2_X1 U147 ( .A1(\mem[1][6] ), .A2(n1200), .ZN(n1193) );
  OAI21_X1 U148 ( .B1(n627), .B2(n1200), .A(n1192), .ZN(n895) );
  NAND2_X1 U149 ( .A1(\mem[1][7] ), .A2(n1200), .ZN(n1192) );
  OAI21_X1 U150 ( .B1(n620), .B2(n1190), .A(n1189), .ZN(n894) );
  NAND2_X1 U151 ( .A1(\mem[2][0] ), .A2(n1190), .ZN(n1189) );
  OAI21_X1 U152 ( .B1(n621), .B2(n1190), .A(n1188), .ZN(n893) );
  NAND2_X1 U153 ( .A1(\mem[2][1] ), .A2(n1190), .ZN(n1188) );
  OAI21_X1 U154 ( .B1(n622), .B2(n1190), .A(n1187), .ZN(n892) );
  NAND2_X1 U155 ( .A1(\mem[2][2] ), .A2(n1190), .ZN(n1187) );
  OAI21_X1 U156 ( .B1(n623), .B2(n1190), .A(n1186), .ZN(n891) );
  NAND2_X1 U157 ( .A1(\mem[2][3] ), .A2(n1190), .ZN(n1186) );
  OAI21_X1 U158 ( .B1(n624), .B2(n1190), .A(n1185), .ZN(n890) );
  NAND2_X1 U159 ( .A1(\mem[2][4] ), .A2(n1190), .ZN(n1185) );
  OAI21_X1 U160 ( .B1(n625), .B2(n1190), .A(n1184), .ZN(n889) );
  NAND2_X1 U161 ( .A1(\mem[2][5] ), .A2(n1190), .ZN(n1184) );
  OAI21_X1 U162 ( .B1(n626), .B2(n1190), .A(n1183), .ZN(n888) );
  NAND2_X1 U163 ( .A1(\mem[2][6] ), .A2(n1190), .ZN(n1183) );
  OAI21_X1 U164 ( .B1(n627), .B2(n1190), .A(n1182), .ZN(n887) );
  NAND2_X1 U165 ( .A1(\mem[2][7] ), .A2(n1190), .ZN(n1182) );
  OAI21_X1 U166 ( .B1(n620), .B2(n1180), .A(n1179), .ZN(n886) );
  NAND2_X1 U167 ( .A1(\mem[3][0] ), .A2(n1180), .ZN(n1179) );
  OAI21_X1 U168 ( .B1(n621), .B2(n1180), .A(n1178), .ZN(n885) );
  NAND2_X1 U169 ( .A1(\mem[3][1] ), .A2(n1180), .ZN(n1178) );
  OAI21_X1 U170 ( .B1(n622), .B2(n1180), .A(n1177), .ZN(n884) );
  NAND2_X1 U171 ( .A1(\mem[3][2] ), .A2(n1180), .ZN(n1177) );
  OAI21_X1 U172 ( .B1(n623), .B2(n1180), .A(n1176), .ZN(n883) );
  NAND2_X1 U173 ( .A1(\mem[3][3] ), .A2(n1180), .ZN(n1176) );
  OAI21_X1 U174 ( .B1(n624), .B2(n1180), .A(n1175), .ZN(n882) );
  NAND2_X1 U175 ( .A1(\mem[3][4] ), .A2(n1180), .ZN(n1175) );
  OAI21_X1 U176 ( .B1(n625), .B2(n1180), .A(n1174), .ZN(n881) );
  NAND2_X1 U177 ( .A1(\mem[3][5] ), .A2(n1180), .ZN(n1174) );
  OAI21_X1 U178 ( .B1(n626), .B2(n1180), .A(n1173), .ZN(n880) );
  NAND2_X1 U179 ( .A1(\mem[3][6] ), .A2(n1180), .ZN(n1173) );
  OAI21_X1 U180 ( .B1(n627), .B2(n1180), .A(n1172), .ZN(n879) );
  NAND2_X1 U181 ( .A1(\mem[3][7] ), .A2(n1180), .ZN(n1172) );
  OAI21_X1 U182 ( .B1(n620), .B2(n1160), .A(n1159), .ZN(n870) );
  NAND2_X1 U183 ( .A1(\mem[5][0] ), .A2(n1160), .ZN(n1159) );
  OAI21_X1 U184 ( .B1(n621), .B2(n1160), .A(n1158), .ZN(n869) );
  NAND2_X1 U185 ( .A1(\mem[5][1] ), .A2(n1160), .ZN(n1158) );
  OAI21_X1 U186 ( .B1(n622), .B2(n1160), .A(n1157), .ZN(n868) );
  NAND2_X1 U187 ( .A1(\mem[5][2] ), .A2(n1160), .ZN(n1157) );
  OAI21_X1 U188 ( .B1(n623), .B2(n1160), .A(n1156), .ZN(n867) );
  NAND2_X1 U189 ( .A1(\mem[5][3] ), .A2(n1160), .ZN(n1156) );
  OAI21_X1 U190 ( .B1(n624), .B2(n1160), .A(n1155), .ZN(n866) );
  NAND2_X1 U191 ( .A1(\mem[5][4] ), .A2(n1160), .ZN(n1155) );
  OAI21_X1 U192 ( .B1(n625), .B2(n1160), .A(n1154), .ZN(n865) );
  NAND2_X1 U193 ( .A1(\mem[5][5] ), .A2(n1160), .ZN(n1154) );
  OAI21_X1 U194 ( .B1(n626), .B2(n1160), .A(n1153), .ZN(n864) );
  NAND2_X1 U195 ( .A1(\mem[5][6] ), .A2(n1160), .ZN(n1153) );
  OAI21_X1 U196 ( .B1(n627), .B2(n1160), .A(n1152), .ZN(n863) );
  NAND2_X1 U197 ( .A1(\mem[5][7] ), .A2(n1160), .ZN(n1152) );
  OAI21_X1 U198 ( .B1(n1211), .B2(n620), .A(n1210), .ZN(n910) );
  NAND2_X1 U199 ( .A1(\mem[0][0] ), .A2(n1211), .ZN(n1210) );
  OAI21_X1 U200 ( .B1(n1211), .B2(n621), .A(n1209), .ZN(n909) );
  NAND2_X1 U201 ( .A1(\mem[0][1] ), .A2(n1211), .ZN(n1209) );
  OAI21_X1 U202 ( .B1(n1211), .B2(n622), .A(n1208), .ZN(n908) );
  NAND2_X1 U203 ( .A1(\mem[0][2] ), .A2(n1211), .ZN(n1208) );
  OAI21_X1 U204 ( .B1(n1211), .B2(n623), .A(n1207), .ZN(n907) );
  NAND2_X1 U205 ( .A1(\mem[0][3] ), .A2(n1211), .ZN(n1207) );
  OAI21_X1 U206 ( .B1(n1211), .B2(n624), .A(n1206), .ZN(n906) );
  NAND2_X1 U207 ( .A1(\mem[0][4] ), .A2(n1211), .ZN(n1206) );
  OAI21_X1 U208 ( .B1(n1211), .B2(n625), .A(n1205), .ZN(n905) );
  NAND2_X1 U209 ( .A1(\mem[0][5] ), .A2(n1211), .ZN(n1205) );
  OAI21_X1 U210 ( .B1(n1211), .B2(n626), .A(n1204), .ZN(n904) );
  NAND2_X1 U211 ( .A1(\mem[0][6] ), .A2(n1211), .ZN(n1204) );
  OAI21_X1 U212 ( .B1(n1211), .B2(n627), .A(n1203), .ZN(n903) );
  NAND2_X1 U213 ( .A1(\mem[0][7] ), .A2(n1211), .ZN(n1203) );
  INV_X1 U214 ( .A(n1129), .ZN(n819) );
  AOI22_X1 U215 ( .A1(data_in[0]), .A2(n843), .B1(n1128), .B2(\mem[8][0] ), 
        .ZN(n1129) );
  INV_X1 U216 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U217 ( .A1(data_in[1]), .A2(n843), .B1(n1128), .B2(\mem[8][1] ), 
        .ZN(n1127) );
  INV_X1 U218 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U219 ( .A1(data_in[2]), .A2(n843), .B1(n1128), .B2(\mem[8][2] ), 
        .ZN(n1126) );
  INV_X1 U220 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U221 ( .A1(data_in[3]), .A2(n843), .B1(n1128), .B2(\mem[8][3] ), 
        .ZN(n1125) );
  INV_X1 U222 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U223 ( .A1(data_in[4]), .A2(n843), .B1(n1128), .B2(\mem[8][4] ), 
        .ZN(n1124) );
  INV_X1 U224 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U225 ( .A1(data_in[5]), .A2(n843), .B1(n1128), .B2(\mem[8][5] ), 
        .ZN(n1123) );
  INV_X1 U226 ( .A(n1122), .ZN(n813) );
  AOI22_X1 U227 ( .A1(data_in[6]), .A2(n843), .B1(n1128), .B2(\mem[8][6] ), 
        .ZN(n1122) );
  INV_X1 U228 ( .A(n1121), .ZN(n812) );
  AOI22_X1 U229 ( .A1(data_in[7]), .A2(n843), .B1(n1128), .B2(\mem[8][7] ), 
        .ZN(n1121) );
  INV_X1 U230 ( .A(n1119), .ZN(n811) );
  AOI22_X1 U231 ( .A1(data_in[0]), .A2(n842), .B1(n1118), .B2(\mem[9][0] ), 
        .ZN(n1119) );
  INV_X1 U232 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U233 ( .A1(data_in[1]), .A2(n842), .B1(n1118), .B2(\mem[9][1] ), 
        .ZN(n1117) );
  INV_X1 U234 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U235 ( .A1(data_in[2]), .A2(n842), .B1(n1118), .B2(\mem[9][2] ), 
        .ZN(n1116) );
  INV_X1 U236 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U237 ( .A1(data_in[3]), .A2(n842), .B1(n1118), .B2(\mem[9][3] ), 
        .ZN(n1115) );
  INV_X1 U238 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U239 ( .A1(data_in[4]), .A2(n842), .B1(n1118), .B2(\mem[9][4] ), 
        .ZN(n1114) );
  INV_X1 U240 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U241 ( .A1(data_in[5]), .A2(n842), .B1(n1118), .B2(\mem[9][5] ), 
        .ZN(n1113) );
  INV_X1 U242 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U243 ( .A1(data_in[6]), .A2(n842), .B1(n1118), .B2(\mem[9][6] ), 
        .ZN(n1112) );
  INV_X1 U244 ( .A(n1111), .ZN(n804) );
  AOI22_X1 U245 ( .A1(data_in[7]), .A2(n842), .B1(n1118), .B2(\mem[9][7] ), 
        .ZN(n1111) );
  INV_X1 U246 ( .A(n1110), .ZN(n803) );
  AOI22_X1 U247 ( .A1(data_in[0]), .A2(n841), .B1(n1109), .B2(\mem[10][0] ), 
        .ZN(n1110) );
  INV_X1 U248 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U249 ( .A1(data_in[1]), .A2(n841), .B1(n1109), .B2(\mem[10][1] ), 
        .ZN(n1108) );
  INV_X1 U250 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U251 ( .A1(data_in[2]), .A2(n841), .B1(n1109), .B2(\mem[10][2] ), 
        .ZN(n1107) );
  INV_X1 U252 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U253 ( .A1(data_in[3]), .A2(n841), .B1(n1109), .B2(\mem[10][3] ), 
        .ZN(n1106) );
  INV_X1 U254 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U255 ( .A1(data_in[4]), .A2(n841), .B1(n1109), .B2(\mem[10][4] ), 
        .ZN(n1105) );
  INV_X1 U256 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U257 ( .A1(data_in[5]), .A2(n841), .B1(n1109), .B2(\mem[10][5] ), 
        .ZN(n1104) );
  INV_X1 U258 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U259 ( .A1(data_in[6]), .A2(n841), .B1(n1109), .B2(\mem[10][6] ), 
        .ZN(n1103) );
  INV_X1 U260 ( .A(n1102), .ZN(n796) );
  AOI22_X1 U261 ( .A1(data_in[7]), .A2(n841), .B1(n1109), .B2(\mem[10][7] ), 
        .ZN(n1102) );
  INV_X1 U262 ( .A(n1101), .ZN(n795) );
  AOI22_X1 U263 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[11][0] ), 
        .ZN(n1101) );
  INV_X1 U264 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U265 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[11][1] ), 
        .ZN(n1099) );
  INV_X1 U266 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U267 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[11][2] ), 
        .ZN(n1098) );
  INV_X1 U268 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U269 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[11][3] ), 
        .ZN(n1097) );
  INV_X1 U270 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U271 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[11][4] ), 
        .ZN(n1096) );
  INV_X1 U272 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U273 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[11][5] ), 
        .ZN(n1095) );
  INV_X1 U274 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U275 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[11][6] ), 
        .ZN(n1094) );
  INV_X1 U276 ( .A(n1093), .ZN(n788) );
  AOI22_X1 U277 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[11][7] ), 
        .ZN(n1093) );
  INV_X1 U278 ( .A(n1092), .ZN(n787) );
  AOI22_X1 U279 ( .A1(data_in[0]), .A2(n839), .B1(n1091), .B2(\mem[12][0] ), 
        .ZN(n1092) );
  INV_X1 U280 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U281 ( .A1(data_in[1]), .A2(n839), .B1(n1091), .B2(\mem[12][1] ), 
        .ZN(n1090) );
  INV_X1 U282 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U283 ( .A1(data_in[2]), .A2(n839), .B1(n1091), .B2(\mem[12][2] ), 
        .ZN(n1089) );
  INV_X1 U284 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U285 ( .A1(data_in[3]), .A2(n839), .B1(n1091), .B2(\mem[12][3] ), 
        .ZN(n1088) );
  INV_X1 U286 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U287 ( .A1(data_in[4]), .A2(n839), .B1(n1091), .B2(\mem[12][4] ), 
        .ZN(n1087) );
  INV_X1 U288 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U289 ( .A1(data_in[5]), .A2(n839), .B1(n1091), .B2(\mem[12][5] ), 
        .ZN(n1086) );
  INV_X1 U290 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U291 ( .A1(data_in[6]), .A2(n839), .B1(n1091), .B2(\mem[12][6] ), 
        .ZN(n1085) );
  INV_X1 U292 ( .A(n1084), .ZN(n780) );
  AOI22_X1 U293 ( .A1(data_in[7]), .A2(n839), .B1(n1091), .B2(\mem[12][7] ), 
        .ZN(n1084) );
  INV_X1 U294 ( .A(n1083), .ZN(n779) );
  AOI22_X1 U295 ( .A1(data_in[0]), .A2(n838), .B1(n1082), .B2(\mem[13][0] ), 
        .ZN(n1083) );
  INV_X1 U296 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U297 ( .A1(data_in[1]), .A2(n838), .B1(n1082), .B2(\mem[13][1] ), 
        .ZN(n1081) );
  INV_X1 U298 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U299 ( .A1(data_in[2]), .A2(n838), .B1(n1082), .B2(\mem[13][2] ), 
        .ZN(n1080) );
  INV_X1 U300 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U301 ( .A1(data_in[3]), .A2(n838), .B1(n1082), .B2(\mem[13][3] ), 
        .ZN(n1079) );
  INV_X1 U302 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U303 ( .A1(data_in[4]), .A2(n838), .B1(n1082), .B2(\mem[13][4] ), 
        .ZN(n1078) );
  INV_X1 U304 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U305 ( .A1(data_in[5]), .A2(n838), .B1(n1082), .B2(\mem[13][5] ), 
        .ZN(n1077) );
  INV_X1 U306 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U307 ( .A1(data_in[6]), .A2(n838), .B1(n1082), .B2(\mem[13][6] ), 
        .ZN(n1076) );
  INV_X1 U308 ( .A(n1075), .ZN(n772) );
  AOI22_X1 U309 ( .A1(data_in[7]), .A2(n838), .B1(n1082), .B2(\mem[13][7] ), 
        .ZN(n1075) );
  INV_X1 U310 ( .A(n1074), .ZN(n771) );
  AOI22_X1 U311 ( .A1(data_in[0]), .A2(n837), .B1(n1073), .B2(\mem[14][0] ), 
        .ZN(n1074) );
  INV_X1 U312 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U313 ( .A1(data_in[1]), .A2(n837), .B1(n1073), .B2(\mem[14][1] ), 
        .ZN(n1072) );
  INV_X1 U314 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U315 ( .A1(data_in[2]), .A2(n837), .B1(n1073), .B2(\mem[14][2] ), 
        .ZN(n1071) );
  INV_X1 U316 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U317 ( .A1(data_in[3]), .A2(n837), .B1(n1073), .B2(\mem[14][3] ), 
        .ZN(n1070) );
  INV_X1 U318 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U319 ( .A1(data_in[4]), .A2(n837), .B1(n1073), .B2(\mem[14][4] ), 
        .ZN(n1069) );
  INV_X1 U320 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U321 ( .A1(data_in[5]), .A2(n837), .B1(n1073), .B2(\mem[14][5] ), 
        .ZN(n1068) );
  INV_X1 U322 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U323 ( .A1(data_in[6]), .A2(n837), .B1(n1073), .B2(\mem[14][6] ), 
        .ZN(n1067) );
  INV_X1 U324 ( .A(n1066), .ZN(n764) );
  AOI22_X1 U325 ( .A1(data_in[7]), .A2(n837), .B1(n1073), .B2(\mem[14][7] ), 
        .ZN(n1066) );
  INV_X1 U326 ( .A(n1065), .ZN(n763) );
  AOI22_X1 U327 ( .A1(data_in[0]), .A2(n836), .B1(n1064), .B2(\mem[15][0] ), 
        .ZN(n1065) );
  INV_X1 U328 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U329 ( .A1(data_in[1]), .A2(n836), .B1(n1064), .B2(\mem[15][1] ), 
        .ZN(n1063) );
  INV_X1 U330 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U331 ( .A1(data_in[2]), .A2(n836), .B1(n1064), .B2(\mem[15][2] ), 
        .ZN(n1062) );
  INV_X1 U332 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U333 ( .A1(data_in[3]), .A2(n836), .B1(n1064), .B2(\mem[15][3] ), 
        .ZN(n1061) );
  INV_X1 U334 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U335 ( .A1(data_in[4]), .A2(n836), .B1(n1064), .B2(\mem[15][4] ), 
        .ZN(n1060) );
  INV_X1 U336 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U337 ( .A1(data_in[5]), .A2(n836), .B1(n1064), .B2(\mem[15][5] ), 
        .ZN(n1059) );
  INV_X1 U338 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U339 ( .A1(data_in[6]), .A2(n836), .B1(n1064), .B2(\mem[15][6] ), 
        .ZN(n1058) );
  INV_X1 U340 ( .A(n1057), .ZN(n756) );
  AOI22_X1 U341 ( .A1(data_in[7]), .A2(n836), .B1(n1064), .B2(\mem[15][7] ), 
        .ZN(n1057) );
  INV_X1 U342 ( .A(n1056), .ZN(n755) );
  AOI22_X1 U343 ( .A1(data_in[0]), .A2(n835), .B1(n1055), .B2(\mem[16][0] ), 
        .ZN(n1056) );
  INV_X1 U344 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U345 ( .A1(data_in[1]), .A2(n835), .B1(n1055), .B2(\mem[16][1] ), 
        .ZN(n1054) );
  INV_X1 U346 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U347 ( .A1(data_in[2]), .A2(n835), .B1(n1055), .B2(\mem[16][2] ), 
        .ZN(n1053) );
  INV_X1 U348 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U349 ( .A1(data_in[3]), .A2(n835), .B1(n1055), .B2(\mem[16][3] ), 
        .ZN(n1052) );
  INV_X1 U350 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U351 ( .A1(data_in[4]), .A2(n835), .B1(n1055), .B2(\mem[16][4] ), 
        .ZN(n1051) );
  INV_X1 U352 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U353 ( .A1(data_in[5]), .A2(n835), .B1(n1055), .B2(\mem[16][5] ), 
        .ZN(n1050) );
  INV_X1 U354 ( .A(n1049), .ZN(n749) );
  AOI22_X1 U355 ( .A1(data_in[6]), .A2(n835), .B1(n1055), .B2(\mem[16][6] ), 
        .ZN(n1049) );
  INV_X1 U356 ( .A(n1048), .ZN(n748) );
  AOI22_X1 U357 ( .A1(data_in[7]), .A2(n835), .B1(n1055), .B2(\mem[16][7] ), 
        .ZN(n1048) );
  INV_X1 U358 ( .A(n1046), .ZN(n747) );
  AOI22_X1 U359 ( .A1(data_in[0]), .A2(n834), .B1(n1045), .B2(\mem[17][0] ), 
        .ZN(n1046) );
  INV_X1 U360 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U361 ( .A1(data_in[1]), .A2(n834), .B1(n1045), .B2(\mem[17][1] ), 
        .ZN(n1044) );
  INV_X1 U362 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U363 ( .A1(data_in[2]), .A2(n834), .B1(n1045), .B2(\mem[17][2] ), 
        .ZN(n1043) );
  INV_X1 U364 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U365 ( .A1(data_in[3]), .A2(n834), .B1(n1045), .B2(\mem[17][3] ), 
        .ZN(n1042) );
  INV_X1 U366 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U367 ( .A1(data_in[4]), .A2(n834), .B1(n1045), .B2(\mem[17][4] ), 
        .ZN(n1041) );
  INV_X1 U368 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U369 ( .A1(data_in[5]), .A2(n834), .B1(n1045), .B2(\mem[17][5] ), 
        .ZN(n1040) );
  INV_X1 U370 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U371 ( .A1(data_in[6]), .A2(n834), .B1(n1045), .B2(\mem[17][6] ), 
        .ZN(n1039) );
  INV_X1 U372 ( .A(n1038), .ZN(n740) );
  AOI22_X1 U373 ( .A1(data_in[7]), .A2(n834), .B1(n1045), .B2(\mem[17][7] ), 
        .ZN(n1038) );
  INV_X1 U374 ( .A(n1037), .ZN(n739) );
  AOI22_X1 U375 ( .A1(data_in[0]), .A2(n833), .B1(n1036), .B2(\mem[18][0] ), 
        .ZN(n1037) );
  INV_X1 U376 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U377 ( .A1(data_in[1]), .A2(n833), .B1(n1036), .B2(\mem[18][1] ), 
        .ZN(n1035) );
  INV_X1 U378 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U379 ( .A1(data_in[2]), .A2(n833), .B1(n1036), .B2(\mem[18][2] ), 
        .ZN(n1034) );
  INV_X1 U380 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U381 ( .A1(data_in[3]), .A2(n833), .B1(n1036), .B2(\mem[18][3] ), 
        .ZN(n1033) );
  INV_X1 U382 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U383 ( .A1(data_in[4]), .A2(n833), .B1(n1036), .B2(\mem[18][4] ), 
        .ZN(n1032) );
  INV_X1 U384 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U385 ( .A1(data_in[5]), .A2(n833), .B1(n1036), .B2(\mem[18][5] ), 
        .ZN(n1031) );
  INV_X1 U386 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U387 ( .A1(data_in[6]), .A2(n833), .B1(n1036), .B2(\mem[18][6] ), 
        .ZN(n1030) );
  INV_X1 U388 ( .A(n1029), .ZN(n732) );
  AOI22_X1 U389 ( .A1(data_in[7]), .A2(n833), .B1(n1036), .B2(\mem[18][7] ), 
        .ZN(n1029) );
  INV_X1 U390 ( .A(n1028), .ZN(n731) );
  AOI22_X1 U391 ( .A1(data_in[0]), .A2(n832), .B1(n1027), .B2(\mem[19][0] ), 
        .ZN(n1028) );
  INV_X1 U392 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U393 ( .A1(data_in[1]), .A2(n832), .B1(n1027), .B2(\mem[19][1] ), 
        .ZN(n1026) );
  INV_X1 U394 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U395 ( .A1(data_in[2]), .A2(n832), .B1(n1027), .B2(\mem[19][2] ), 
        .ZN(n1025) );
  INV_X1 U396 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U397 ( .A1(data_in[3]), .A2(n832), .B1(n1027), .B2(\mem[19][3] ), 
        .ZN(n1024) );
  INV_X1 U398 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U399 ( .A1(data_in[4]), .A2(n832), .B1(n1027), .B2(\mem[19][4] ), 
        .ZN(n1023) );
  INV_X1 U400 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U401 ( .A1(data_in[5]), .A2(n832), .B1(n1027), .B2(\mem[19][5] ), 
        .ZN(n1022) );
  INV_X1 U402 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U403 ( .A1(data_in[6]), .A2(n832), .B1(n1027), .B2(\mem[19][6] ), 
        .ZN(n1021) );
  INV_X1 U404 ( .A(n1020), .ZN(n724) );
  AOI22_X1 U405 ( .A1(data_in[7]), .A2(n832), .B1(n1027), .B2(\mem[19][7] ), 
        .ZN(n1020) );
  INV_X1 U406 ( .A(n1019), .ZN(n723) );
  AOI22_X1 U407 ( .A1(data_in[0]), .A2(n831), .B1(n1018), .B2(\mem[20][0] ), 
        .ZN(n1019) );
  INV_X1 U408 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U409 ( .A1(data_in[1]), .A2(n831), .B1(n1018), .B2(\mem[20][1] ), 
        .ZN(n1017) );
  INV_X1 U410 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U411 ( .A1(data_in[2]), .A2(n831), .B1(n1018), .B2(\mem[20][2] ), 
        .ZN(n1016) );
  INV_X1 U412 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U413 ( .A1(data_in[3]), .A2(n831), .B1(n1018), .B2(\mem[20][3] ), 
        .ZN(n1015) );
  INV_X1 U414 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U415 ( .A1(data_in[4]), .A2(n831), .B1(n1018), .B2(\mem[20][4] ), 
        .ZN(n1014) );
  INV_X1 U416 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U417 ( .A1(data_in[5]), .A2(n831), .B1(n1018), .B2(\mem[20][5] ), 
        .ZN(n1013) );
  INV_X1 U418 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U419 ( .A1(data_in[6]), .A2(n831), .B1(n1018), .B2(\mem[20][6] ), 
        .ZN(n1012) );
  INV_X1 U420 ( .A(n1011), .ZN(n716) );
  AOI22_X1 U421 ( .A1(data_in[7]), .A2(n831), .B1(n1018), .B2(\mem[20][7] ), 
        .ZN(n1011) );
  INV_X1 U422 ( .A(n1010), .ZN(n715) );
  AOI22_X1 U423 ( .A1(data_in[0]), .A2(n830), .B1(n1009), .B2(\mem[21][0] ), 
        .ZN(n1010) );
  INV_X1 U424 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U425 ( .A1(data_in[1]), .A2(n830), .B1(n1009), .B2(\mem[21][1] ), 
        .ZN(n1008) );
  INV_X1 U426 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U427 ( .A1(data_in[2]), .A2(n830), .B1(n1009), .B2(\mem[21][2] ), 
        .ZN(n1007) );
  INV_X1 U428 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U429 ( .A1(data_in[3]), .A2(n830), .B1(n1009), .B2(\mem[21][3] ), 
        .ZN(n1006) );
  INV_X1 U430 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U431 ( .A1(data_in[4]), .A2(n830), .B1(n1009), .B2(\mem[21][4] ), 
        .ZN(n1005) );
  INV_X1 U432 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U433 ( .A1(data_in[5]), .A2(n830), .B1(n1009), .B2(\mem[21][5] ), 
        .ZN(n1004) );
  INV_X1 U434 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U435 ( .A1(data_in[6]), .A2(n830), .B1(n1009), .B2(\mem[21][6] ), 
        .ZN(n1003) );
  INV_X1 U436 ( .A(n1002), .ZN(n708) );
  AOI22_X1 U437 ( .A1(data_in[7]), .A2(n830), .B1(n1009), .B2(\mem[21][7] ), 
        .ZN(n1002) );
  INV_X1 U438 ( .A(n1001), .ZN(n707) );
  AOI22_X1 U439 ( .A1(data_in[0]), .A2(n829), .B1(n1000), .B2(\mem[22][0] ), 
        .ZN(n1001) );
  INV_X1 U440 ( .A(n999), .ZN(n706) );
  AOI22_X1 U441 ( .A1(data_in[1]), .A2(n829), .B1(n1000), .B2(\mem[22][1] ), 
        .ZN(n999) );
  INV_X1 U442 ( .A(n998), .ZN(n705) );
  AOI22_X1 U443 ( .A1(data_in[2]), .A2(n829), .B1(n1000), .B2(\mem[22][2] ), 
        .ZN(n998) );
  INV_X1 U444 ( .A(n997), .ZN(n704) );
  AOI22_X1 U445 ( .A1(data_in[3]), .A2(n829), .B1(n1000), .B2(\mem[22][3] ), 
        .ZN(n997) );
  INV_X1 U446 ( .A(n996), .ZN(n703) );
  AOI22_X1 U447 ( .A1(data_in[4]), .A2(n829), .B1(n1000), .B2(\mem[22][4] ), 
        .ZN(n996) );
  INV_X1 U448 ( .A(n995), .ZN(n702) );
  AOI22_X1 U449 ( .A1(data_in[5]), .A2(n829), .B1(n1000), .B2(\mem[22][5] ), 
        .ZN(n995) );
  INV_X1 U450 ( .A(n994), .ZN(n701) );
  AOI22_X1 U451 ( .A1(data_in[6]), .A2(n829), .B1(n1000), .B2(\mem[22][6] ), 
        .ZN(n994) );
  INV_X1 U452 ( .A(n993), .ZN(n700) );
  AOI22_X1 U453 ( .A1(data_in[7]), .A2(n829), .B1(n1000), .B2(\mem[22][7] ), 
        .ZN(n993) );
  INV_X1 U454 ( .A(n992), .ZN(n699) );
  AOI22_X1 U455 ( .A1(data_in[0]), .A2(n828), .B1(n991), .B2(\mem[23][0] ), 
        .ZN(n992) );
  INV_X1 U456 ( .A(n990), .ZN(n698) );
  AOI22_X1 U457 ( .A1(data_in[1]), .A2(n828), .B1(n991), .B2(\mem[23][1] ), 
        .ZN(n990) );
  INV_X1 U458 ( .A(n989), .ZN(n697) );
  AOI22_X1 U459 ( .A1(data_in[2]), .A2(n828), .B1(n991), .B2(\mem[23][2] ), 
        .ZN(n989) );
  INV_X1 U460 ( .A(n988), .ZN(n696) );
  AOI22_X1 U461 ( .A1(data_in[3]), .A2(n828), .B1(n991), .B2(\mem[23][3] ), 
        .ZN(n988) );
  INV_X1 U462 ( .A(n987), .ZN(n695) );
  AOI22_X1 U463 ( .A1(data_in[4]), .A2(n828), .B1(n991), .B2(\mem[23][4] ), 
        .ZN(n987) );
  INV_X1 U464 ( .A(n986), .ZN(n694) );
  AOI22_X1 U465 ( .A1(data_in[5]), .A2(n828), .B1(n991), .B2(\mem[23][5] ), 
        .ZN(n986) );
  INV_X1 U466 ( .A(n985), .ZN(n693) );
  AOI22_X1 U467 ( .A1(data_in[6]), .A2(n828), .B1(n991), .B2(\mem[23][6] ), 
        .ZN(n985) );
  INV_X1 U468 ( .A(n984), .ZN(n692) );
  AOI22_X1 U469 ( .A1(data_in[7]), .A2(n828), .B1(n991), .B2(\mem[23][7] ), 
        .ZN(n984) );
  INV_X1 U470 ( .A(n983), .ZN(n691) );
  AOI22_X1 U471 ( .A1(data_in[0]), .A2(n827), .B1(n982), .B2(\mem[24][0] ), 
        .ZN(n983) );
  INV_X1 U472 ( .A(n981), .ZN(n690) );
  AOI22_X1 U473 ( .A1(data_in[1]), .A2(n827), .B1(n982), .B2(\mem[24][1] ), 
        .ZN(n981) );
  INV_X1 U474 ( .A(n980), .ZN(n689) );
  AOI22_X1 U475 ( .A1(data_in[2]), .A2(n827), .B1(n982), .B2(\mem[24][2] ), 
        .ZN(n980) );
  INV_X1 U476 ( .A(n979), .ZN(n688) );
  AOI22_X1 U477 ( .A1(data_in[3]), .A2(n827), .B1(n982), .B2(\mem[24][3] ), 
        .ZN(n979) );
  INV_X1 U478 ( .A(n978), .ZN(n687) );
  AOI22_X1 U479 ( .A1(data_in[4]), .A2(n827), .B1(n982), .B2(\mem[24][4] ), 
        .ZN(n978) );
  INV_X1 U480 ( .A(n977), .ZN(n686) );
  AOI22_X1 U481 ( .A1(data_in[5]), .A2(n827), .B1(n982), .B2(\mem[24][5] ), 
        .ZN(n977) );
  INV_X1 U482 ( .A(n976), .ZN(n685) );
  AOI22_X1 U483 ( .A1(data_in[6]), .A2(n827), .B1(n982), .B2(\mem[24][6] ), 
        .ZN(n976) );
  INV_X1 U484 ( .A(n975), .ZN(n684) );
  AOI22_X1 U485 ( .A1(data_in[7]), .A2(n827), .B1(n982), .B2(\mem[24][7] ), 
        .ZN(n975) );
  INV_X1 U486 ( .A(n973), .ZN(n683) );
  AOI22_X1 U487 ( .A1(data_in[0]), .A2(n826), .B1(n972), .B2(\mem[25][0] ), 
        .ZN(n973) );
  INV_X1 U488 ( .A(n971), .ZN(n682) );
  AOI22_X1 U489 ( .A1(data_in[1]), .A2(n826), .B1(n972), .B2(\mem[25][1] ), 
        .ZN(n971) );
  INV_X1 U490 ( .A(n970), .ZN(n681) );
  AOI22_X1 U491 ( .A1(data_in[2]), .A2(n826), .B1(n972), .B2(\mem[25][2] ), 
        .ZN(n970) );
  INV_X1 U492 ( .A(n969), .ZN(n680) );
  AOI22_X1 U493 ( .A1(data_in[3]), .A2(n826), .B1(n972), .B2(\mem[25][3] ), 
        .ZN(n969) );
  INV_X1 U494 ( .A(n968), .ZN(n679) );
  AOI22_X1 U495 ( .A1(data_in[4]), .A2(n826), .B1(n972), .B2(\mem[25][4] ), 
        .ZN(n968) );
  INV_X1 U496 ( .A(n967), .ZN(n678) );
  AOI22_X1 U497 ( .A1(data_in[5]), .A2(n826), .B1(n972), .B2(\mem[25][5] ), 
        .ZN(n967) );
  INV_X1 U498 ( .A(n966), .ZN(n677) );
  AOI22_X1 U499 ( .A1(data_in[6]), .A2(n826), .B1(n972), .B2(\mem[25][6] ), 
        .ZN(n966) );
  INV_X1 U500 ( .A(n965), .ZN(n676) );
  AOI22_X1 U501 ( .A1(data_in[7]), .A2(n826), .B1(n972), .B2(\mem[25][7] ), 
        .ZN(n965) );
  INV_X1 U502 ( .A(n964), .ZN(n675) );
  AOI22_X1 U503 ( .A1(data_in[0]), .A2(n825), .B1(n963), .B2(\mem[26][0] ), 
        .ZN(n964) );
  INV_X1 U504 ( .A(n962), .ZN(n674) );
  AOI22_X1 U505 ( .A1(data_in[1]), .A2(n825), .B1(n963), .B2(\mem[26][1] ), 
        .ZN(n962) );
  INV_X1 U506 ( .A(n961), .ZN(n673) );
  AOI22_X1 U507 ( .A1(data_in[2]), .A2(n825), .B1(n963), .B2(\mem[26][2] ), 
        .ZN(n961) );
  INV_X1 U508 ( .A(n960), .ZN(n672) );
  AOI22_X1 U509 ( .A1(data_in[3]), .A2(n825), .B1(n963), .B2(\mem[26][3] ), 
        .ZN(n960) );
  INV_X1 U510 ( .A(n959), .ZN(n671) );
  AOI22_X1 U511 ( .A1(data_in[4]), .A2(n825), .B1(n963), .B2(\mem[26][4] ), 
        .ZN(n959) );
  INV_X1 U512 ( .A(n958), .ZN(n670) );
  AOI22_X1 U513 ( .A1(data_in[5]), .A2(n825), .B1(n963), .B2(\mem[26][5] ), 
        .ZN(n958) );
  INV_X1 U514 ( .A(n957), .ZN(n669) );
  AOI22_X1 U515 ( .A1(data_in[6]), .A2(n825), .B1(n963), .B2(\mem[26][6] ), 
        .ZN(n957) );
  INV_X1 U516 ( .A(n956), .ZN(n668) );
  AOI22_X1 U517 ( .A1(data_in[7]), .A2(n825), .B1(n963), .B2(\mem[26][7] ), 
        .ZN(n956) );
  INV_X1 U518 ( .A(n955), .ZN(n667) );
  AOI22_X1 U519 ( .A1(data_in[0]), .A2(n824), .B1(n954), .B2(\mem[27][0] ), 
        .ZN(n955) );
  INV_X1 U520 ( .A(n953), .ZN(n666) );
  AOI22_X1 U521 ( .A1(data_in[1]), .A2(n824), .B1(n954), .B2(\mem[27][1] ), 
        .ZN(n953) );
  INV_X1 U522 ( .A(n952), .ZN(n665) );
  AOI22_X1 U523 ( .A1(data_in[2]), .A2(n824), .B1(n954), .B2(\mem[27][2] ), 
        .ZN(n952) );
  INV_X1 U524 ( .A(n951), .ZN(n664) );
  AOI22_X1 U525 ( .A1(data_in[3]), .A2(n824), .B1(n954), .B2(\mem[27][3] ), 
        .ZN(n951) );
  INV_X1 U526 ( .A(n950), .ZN(n663) );
  AOI22_X1 U527 ( .A1(data_in[4]), .A2(n824), .B1(n954), .B2(\mem[27][4] ), 
        .ZN(n950) );
  INV_X1 U528 ( .A(n949), .ZN(n662) );
  AOI22_X1 U529 ( .A1(data_in[5]), .A2(n824), .B1(n954), .B2(\mem[27][5] ), 
        .ZN(n949) );
  INV_X1 U530 ( .A(n948), .ZN(n661) );
  AOI22_X1 U531 ( .A1(data_in[6]), .A2(n824), .B1(n954), .B2(\mem[27][6] ), 
        .ZN(n948) );
  INV_X1 U532 ( .A(n947), .ZN(n660) );
  AOI22_X1 U533 ( .A1(data_in[7]), .A2(n824), .B1(n954), .B2(\mem[27][7] ), 
        .ZN(n947) );
  INV_X1 U534 ( .A(n946), .ZN(n659) );
  AOI22_X1 U535 ( .A1(data_in[0]), .A2(n823), .B1(n945), .B2(\mem[28][0] ), 
        .ZN(n946) );
  INV_X1 U536 ( .A(n944), .ZN(n658) );
  AOI22_X1 U537 ( .A1(data_in[1]), .A2(n823), .B1(n945), .B2(\mem[28][1] ), 
        .ZN(n944) );
  INV_X1 U538 ( .A(n943), .ZN(n657) );
  AOI22_X1 U539 ( .A1(data_in[2]), .A2(n823), .B1(n945), .B2(\mem[28][2] ), 
        .ZN(n943) );
  INV_X1 U540 ( .A(n942), .ZN(n656) );
  AOI22_X1 U541 ( .A1(data_in[3]), .A2(n823), .B1(n945), .B2(\mem[28][3] ), 
        .ZN(n942) );
  INV_X1 U542 ( .A(n941), .ZN(n655) );
  AOI22_X1 U543 ( .A1(data_in[4]), .A2(n823), .B1(n945), .B2(\mem[28][4] ), 
        .ZN(n941) );
  INV_X1 U544 ( .A(n940), .ZN(n654) );
  AOI22_X1 U545 ( .A1(data_in[5]), .A2(n823), .B1(n945), .B2(\mem[28][5] ), 
        .ZN(n940) );
  INV_X1 U546 ( .A(n939), .ZN(n653) );
  AOI22_X1 U547 ( .A1(data_in[6]), .A2(n823), .B1(n945), .B2(\mem[28][6] ), 
        .ZN(n939) );
  INV_X1 U548 ( .A(n938), .ZN(n652) );
  AOI22_X1 U549 ( .A1(data_in[7]), .A2(n823), .B1(n945), .B2(\mem[28][7] ), 
        .ZN(n938) );
  INV_X1 U550 ( .A(n937), .ZN(n651) );
  AOI22_X1 U551 ( .A1(data_in[0]), .A2(n822), .B1(n936), .B2(\mem[29][0] ), 
        .ZN(n937) );
  INV_X1 U552 ( .A(n935), .ZN(n650) );
  AOI22_X1 U553 ( .A1(data_in[1]), .A2(n822), .B1(n936), .B2(\mem[29][1] ), 
        .ZN(n935) );
  INV_X1 U554 ( .A(n934), .ZN(n649) );
  AOI22_X1 U555 ( .A1(data_in[2]), .A2(n822), .B1(n936), .B2(\mem[29][2] ), 
        .ZN(n934) );
  INV_X1 U556 ( .A(n933), .ZN(n648) );
  AOI22_X1 U557 ( .A1(data_in[3]), .A2(n822), .B1(n936), .B2(\mem[29][3] ), 
        .ZN(n933) );
  INV_X1 U558 ( .A(n932), .ZN(n647) );
  AOI22_X1 U559 ( .A1(data_in[4]), .A2(n822), .B1(n936), .B2(\mem[29][4] ), 
        .ZN(n932) );
  INV_X1 U560 ( .A(n931), .ZN(n646) );
  AOI22_X1 U561 ( .A1(data_in[5]), .A2(n822), .B1(n936), .B2(\mem[29][5] ), 
        .ZN(n931) );
  INV_X1 U562 ( .A(n930), .ZN(n645) );
  AOI22_X1 U563 ( .A1(data_in[6]), .A2(n822), .B1(n936), .B2(\mem[29][6] ), 
        .ZN(n930) );
  INV_X1 U564 ( .A(n929), .ZN(n644) );
  AOI22_X1 U565 ( .A1(data_in[7]), .A2(n822), .B1(n936), .B2(\mem[29][7] ), 
        .ZN(n929) );
  INV_X1 U566 ( .A(n928), .ZN(n643) );
  AOI22_X1 U567 ( .A1(data_in[0]), .A2(n821), .B1(n927), .B2(\mem[30][0] ), 
        .ZN(n928) );
  INV_X1 U568 ( .A(n926), .ZN(n642) );
  AOI22_X1 U569 ( .A1(data_in[1]), .A2(n821), .B1(n927), .B2(\mem[30][1] ), 
        .ZN(n926) );
  INV_X1 U570 ( .A(n925), .ZN(n641) );
  AOI22_X1 U571 ( .A1(data_in[2]), .A2(n821), .B1(n927), .B2(\mem[30][2] ), 
        .ZN(n925) );
  INV_X1 U572 ( .A(n924), .ZN(n640) );
  AOI22_X1 U573 ( .A1(data_in[3]), .A2(n821), .B1(n927), .B2(\mem[30][3] ), 
        .ZN(n924) );
  INV_X1 U574 ( .A(n923), .ZN(n639) );
  AOI22_X1 U575 ( .A1(data_in[4]), .A2(n821), .B1(n927), .B2(\mem[30][4] ), 
        .ZN(n923) );
  INV_X1 U576 ( .A(n922), .ZN(n638) );
  AOI22_X1 U577 ( .A1(data_in[5]), .A2(n821), .B1(n927), .B2(\mem[30][5] ), 
        .ZN(n922) );
  INV_X1 U578 ( .A(n921), .ZN(n637) );
  AOI22_X1 U579 ( .A1(data_in[6]), .A2(n821), .B1(n927), .B2(\mem[30][6] ), 
        .ZN(n921) );
  INV_X1 U580 ( .A(n920), .ZN(n636) );
  AOI22_X1 U581 ( .A1(data_in[7]), .A2(n821), .B1(n927), .B2(\mem[30][7] ), 
        .ZN(n920) );
  INV_X1 U582 ( .A(n919), .ZN(n635) );
  AOI22_X1 U583 ( .A1(data_in[0]), .A2(n820), .B1(n918), .B2(\mem[31][0] ), 
        .ZN(n919) );
  INV_X1 U584 ( .A(n917), .ZN(n634) );
  AOI22_X1 U585 ( .A1(data_in[1]), .A2(n820), .B1(n918), .B2(\mem[31][1] ), 
        .ZN(n917) );
  INV_X1 U586 ( .A(n916), .ZN(n633) );
  AOI22_X1 U587 ( .A1(data_in[2]), .A2(n820), .B1(n918), .B2(\mem[31][2] ), 
        .ZN(n916) );
  INV_X1 U588 ( .A(n915), .ZN(n632) );
  AOI22_X1 U589 ( .A1(data_in[3]), .A2(n820), .B1(n918), .B2(\mem[31][3] ), 
        .ZN(n915) );
  INV_X1 U590 ( .A(n914), .ZN(n631) );
  AOI22_X1 U591 ( .A1(data_in[4]), .A2(n820), .B1(n918), .B2(\mem[31][4] ), 
        .ZN(n914) );
  INV_X1 U592 ( .A(n913), .ZN(n630) );
  AOI22_X1 U593 ( .A1(data_in[5]), .A2(n820), .B1(n918), .B2(\mem[31][5] ), 
        .ZN(n913) );
  INV_X1 U594 ( .A(n912), .ZN(n629) );
  AOI22_X1 U595 ( .A1(data_in[6]), .A2(n820), .B1(n918), .B2(\mem[31][6] ), 
        .ZN(n912) );
  INV_X1 U596 ( .A(n911), .ZN(n628) );
  AOI22_X1 U597 ( .A1(data_in[7]), .A2(n820), .B1(n918), .B2(\mem[31][7] ), 
        .ZN(n911) );
  MUX2_X1 U598 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n611), .Z(n1) );
  MUX2_X1 U599 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n611), .Z(n2) );
  MUX2_X1 U600 ( .A(n2), .B(n1), .S(n608), .Z(n3) );
  MUX2_X1 U601 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n611), .Z(n4) );
  MUX2_X1 U602 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n611), .Z(n5) );
  MUX2_X1 U603 ( .A(n5), .B(n4), .S(n608), .Z(n6) );
  MUX2_X1 U604 ( .A(n6), .B(n3), .S(n606), .Z(n7) );
  MUX2_X1 U605 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n611), .Z(n8) );
  MUX2_X1 U606 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n611), .Z(n9) );
  MUX2_X1 U607 ( .A(n9), .B(n8), .S(n608), .Z(n10) );
  MUX2_X1 U608 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n611), .Z(n11) );
  MUX2_X1 U609 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n611), .Z(n12) );
  MUX2_X1 U610 ( .A(n12), .B(n11), .S(n608), .Z(n13) );
  MUX2_X1 U611 ( .A(n13), .B(n10), .S(n606), .Z(n14) );
  MUX2_X1 U612 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U613 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n612), .Z(n16) );
  MUX2_X1 U614 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n612), .Z(n17) );
  MUX2_X1 U615 ( .A(n17), .B(n16), .S(n609), .Z(n18) );
  MUX2_X1 U616 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n612), .Z(n19) );
  MUX2_X1 U617 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n612), .Z(n20) );
  MUX2_X1 U618 ( .A(n20), .B(n19), .S(n609), .Z(n21) );
  MUX2_X1 U619 ( .A(n21), .B(n18), .S(n606), .Z(n22) );
  MUX2_X1 U620 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n612), .Z(n23) );
  MUX2_X1 U621 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n612), .Z(n24) );
  MUX2_X1 U622 ( .A(n24), .B(n23), .S(n609), .Z(n25) );
  MUX2_X1 U623 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n612), .Z(n26) );
  MUX2_X1 U624 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n612), .Z(n27) );
  MUX2_X1 U625 ( .A(n27), .B(n26), .S(n609), .Z(n28) );
  MUX2_X1 U626 ( .A(n28), .B(n25), .S(n606), .Z(n29) );
  MUX2_X1 U627 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U628 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U629 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n612), .Z(n31) );
  MUX2_X1 U630 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n612), .Z(n32) );
  MUX2_X1 U631 ( .A(n32), .B(n31), .S(n609), .Z(n33) );
  MUX2_X1 U632 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n612), .Z(n34) );
  MUX2_X1 U633 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n612), .Z(n35) );
  MUX2_X1 U634 ( .A(n35), .B(n34), .S(n609), .Z(n36) );
  MUX2_X1 U635 ( .A(n36), .B(n33), .S(n606), .Z(n37) );
  MUX2_X1 U636 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n613), .Z(n38) );
  MUX2_X1 U637 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n613), .Z(n39) );
  MUX2_X1 U638 ( .A(n39), .B(n38), .S(n609), .Z(n40) );
  MUX2_X1 U639 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n613), .Z(n41) );
  MUX2_X1 U640 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n613), .Z(n42) );
  MUX2_X1 U641 ( .A(n42), .B(n41), .S(n609), .Z(n43) );
  MUX2_X1 U642 ( .A(n43), .B(n40), .S(n606), .Z(n44) );
  MUX2_X1 U643 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U644 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n613), .Z(n46) );
  MUX2_X1 U645 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n613), .Z(n47) );
  MUX2_X1 U646 ( .A(n47), .B(n46), .S(n609), .Z(n48) );
  MUX2_X1 U647 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n613), .Z(n49) );
  MUX2_X1 U648 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n613), .Z(n50) );
  MUX2_X1 U649 ( .A(n50), .B(n49), .S(n609), .Z(n51) );
  MUX2_X1 U650 ( .A(n51), .B(n48), .S(n606), .Z(n52) );
  MUX2_X1 U651 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n613), .Z(n53) );
  MUX2_X1 U652 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n613), .Z(n54) );
  MUX2_X1 U653 ( .A(n54), .B(n53), .S(n609), .Z(n55) );
  MUX2_X1 U654 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n613), .Z(n56) );
  MUX2_X1 U655 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n613), .Z(n57) );
  MUX2_X1 U656 ( .A(n57), .B(n56), .S(n609), .Z(n58) );
  MUX2_X1 U657 ( .A(n58), .B(n55), .S(n606), .Z(n59) );
  MUX2_X1 U658 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U659 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U660 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n614), .Z(n61) );
  MUX2_X1 U661 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n614), .Z(n62) );
  MUX2_X1 U662 ( .A(n62), .B(n61), .S(n610), .Z(n63) );
  MUX2_X1 U663 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n614), .Z(n64) );
  MUX2_X1 U664 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n614), .Z(n65) );
  MUX2_X1 U665 ( .A(n65), .B(n64), .S(n610), .Z(n66) );
  MUX2_X1 U666 ( .A(n66), .B(n63), .S(n607), .Z(n67) );
  MUX2_X1 U667 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n614), .Z(n68) );
  MUX2_X1 U668 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n614), .Z(n69) );
  MUX2_X1 U669 ( .A(n69), .B(n68), .S(n610), .Z(n70) );
  MUX2_X1 U670 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n614), .Z(n71) );
  MUX2_X1 U671 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n614), .Z(n72) );
  MUX2_X1 U672 ( .A(n72), .B(n71), .S(n610), .Z(n73) );
  MUX2_X1 U673 ( .A(n73), .B(n70), .S(n607), .Z(n74) );
  MUX2_X1 U674 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U675 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n614), .Z(n76) );
  MUX2_X1 U676 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n614), .Z(n77) );
  MUX2_X1 U677 ( .A(n77), .B(n76), .S(n610), .Z(n78) );
  MUX2_X1 U678 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n614), .Z(n79) );
  MUX2_X1 U679 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n614), .Z(n80) );
  MUX2_X1 U680 ( .A(n80), .B(n79), .S(n610), .Z(n81) );
  MUX2_X1 U681 ( .A(n81), .B(n78), .S(n607), .Z(n82) );
  MUX2_X1 U682 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n615), .Z(n83) );
  MUX2_X1 U683 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n615), .Z(n84) );
  MUX2_X1 U684 ( .A(n84), .B(n83), .S(n610), .Z(n85) );
  MUX2_X1 U685 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n615), .Z(n86) );
  MUX2_X1 U686 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n615), .Z(n87) );
  MUX2_X1 U687 ( .A(n87), .B(n86), .S(n610), .Z(n88) );
  MUX2_X1 U688 ( .A(n88), .B(n85), .S(n607), .Z(n89) );
  MUX2_X1 U689 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U690 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U691 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n615), .Z(n91) );
  MUX2_X1 U692 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n615), .Z(n92) );
  MUX2_X1 U693 ( .A(n92), .B(n91), .S(n610), .Z(n93) );
  MUX2_X1 U694 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n615), .Z(n94) );
  MUX2_X1 U695 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n615), .Z(n95) );
  MUX2_X1 U696 ( .A(n95), .B(n94), .S(n610), .Z(n96) );
  MUX2_X1 U697 ( .A(n96), .B(n93), .S(n607), .Z(n97) );
  MUX2_X1 U698 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n615), .Z(n98) );
  MUX2_X1 U699 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n615), .Z(n99) );
  MUX2_X1 U700 ( .A(n99), .B(n98), .S(n610), .Z(n100) );
  MUX2_X1 U701 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n615), .Z(n101) );
  MUX2_X1 U702 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n615), .Z(n102) );
  MUX2_X1 U703 ( .A(n102), .B(n101), .S(n610), .Z(n103) );
  MUX2_X1 U704 ( .A(n103), .B(n100), .S(n607), .Z(n104) );
  MUX2_X1 U705 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U706 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n613), .Z(n106) );
  MUX2_X1 U707 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n612), .Z(n107) );
  MUX2_X1 U708 ( .A(n107), .B(n106), .S(n610), .Z(n108) );
  MUX2_X1 U709 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n614), .Z(n109) );
  MUX2_X1 U710 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n611), .Z(n110) );
  MUX2_X1 U711 ( .A(n110), .B(n109), .S(n609), .Z(n111) );
  MUX2_X1 U712 ( .A(n111), .B(n108), .S(n607), .Z(n112) );
  MUX2_X1 U713 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n612), .Z(n113) );
  MUX2_X1 U714 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n611), .Z(n114) );
  MUX2_X1 U715 ( .A(n114), .B(n113), .S(n608), .Z(n115) );
  MUX2_X1 U716 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n614), .Z(n116) );
  MUX2_X1 U717 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n612), .Z(n117) );
  MUX2_X1 U718 ( .A(n117), .B(n116), .S(n610), .Z(n118) );
  MUX2_X1 U719 ( .A(n118), .B(n115), .S(n607), .Z(n119) );
  MUX2_X1 U720 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U721 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U722 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n613), .Z(n121) );
  MUX2_X1 U723 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n617), .Z(n122) );
  MUX2_X1 U724 ( .A(n122), .B(n121), .S(n608), .Z(n123) );
  MUX2_X1 U725 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n611), .Z(n124) );
  MUX2_X1 U726 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n125) );
  MUX2_X1 U727 ( .A(n125), .B(n124), .S(n608), .Z(n126) );
  MUX2_X1 U728 ( .A(n126), .B(n123), .S(n607), .Z(n127) );
  MUX2_X1 U729 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n611), .Z(n128) );
  MUX2_X1 U730 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n611), .Z(n129) );
  MUX2_X1 U731 ( .A(n129), .B(n128), .S(n610), .Z(n130) );
  MUX2_X1 U732 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n614), .Z(n131) );
  MUX2_X1 U733 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n614), .Z(n132) );
  MUX2_X1 U734 ( .A(n132), .B(n131), .S(n609), .Z(n133) );
  MUX2_X1 U735 ( .A(n133), .B(n130), .S(n607), .Z(n134) );
  MUX2_X1 U736 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U737 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n612), .Z(n136) );
  MUX2_X1 U738 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n612), .Z(n137) );
  MUX2_X1 U739 ( .A(n137), .B(n136), .S(n609), .Z(n138) );
  MUX2_X1 U740 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n611), .Z(n139) );
  MUX2_X1 U741 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n613), .Z(n140) );
  MUX2_X1 U742 ( .A(n140), .B(n139), .S(n608), .Z(n141) );
  MUX2_X1 U743 ( .A(n141), .B(n138), .S(n607), .Z(n142) );
  MUX2_X1 U744 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n613), .Z(n143) );
  MUX2_X1 U745 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n613), .Z(n144) );
  MUX2_X1 U746 ( .A(n144), .B(n143), .S(n609), .Z(n145) );
  MUX2_X1 U747 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n612), .Z(n146) );
  MUX2_X1 U748 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n614), .Z(n147) );
  MUX2_X1 U749 ( .A(n147), .B(n146), .S(n608), .Z(n148) );
  MUX2_X1 U750 ( .A(n148), .B(n145), .S(n607), .Z(n149) );
  MUX2_X1 U751 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U752 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U753 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n611), .Z(n151) );
  MUX2_X1 U754 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n612), .Z(n152) );
  MUX2_X1 U755 ( .A(n152), .B(n151), .S(n609), .Z(n153) );
  MUX2_X1 U756 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n613), .Z(n154) );
  MUX2_X1 U757 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n611), .Z(n155) );
  MUX2_X1 U758 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U759 ( .A(n156), .B(n153), .S(n606), .Z(n157) );
  MUX2_X1 U760 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n611), .Z(n158) );
  MUX2_X1 U761 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n611), .Z(n159) );
  MUX2_X1 U762 ( .A(n159), .B(n158), .S(n608), .Z(n160) );
  MUX2_X1 U763 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n614), .Z(n161) );
  MUX2_X1 U764 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n614), .Z(n162) );
  MUX2_X1 U765 ( .A(n162), .B(n161), .S(N11), .Z(n163) );
  MUX2_X1 U766 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U767 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U768 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n614), .Z(n166) );
  MUX2_X1 U769 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n612), .Z(n167) );
  MUX2_X1 U770 ( .A(n167), .B(n166), .S(n610), .Z(n168) );
  MUX2_X1 U771 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n613), .Z(n169) );
  MUX2_X1 U772 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n613), .Z(n170) );
  MUX2_X1 U773 ( .A(n170), .B(n169), .S(n610), .Z(n171) );
  MUX2_X1 U774 ( .A(n171), .B(n168), .S(n606), .Z(n172) );
  MUX2_X1 U775 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n616), .Z(n173) );
  MUX2_X1 U776 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n616), .Z(n174) );
  MUX2_X1 U777 ( .A(n174), .B(n173), .S(n610), .Z(n175) );
  MUX2_X1 U778 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n616), .Z(n176) );
  MUX2_X1 U779 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n616), .Z(n177) );
  MUX2_X1 U780 ( .A(n177), .B(n176), .S(n609), .Z(n178) );
  MUX2_X1 U781 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U782 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U783 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U784 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n616), .Z(n181) );
  MUX2_X1 U785 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n616), .Z(n182) );
  MUX2_X1 U786 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U787 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n616), .Z(n184) );
  MUX2_X1 U788 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n616), .Z(n185) );
  MUX2_X1 U789 ( .A(n185), .B(n184), .S(N11), .Z(n186) );
  MUX2_X1 U790 ( .A(n186), .B(n183), .S(n606), .Z(n187) );
  MUX2_X1 U791 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n616), .Z(n188) );
  MUX2_X1 U792 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n616), .Z(n189) );
  MUX2_X1 U793 ( .A(n189), .B(n188), .S(n609), .Z(n190) );
  MUX2_X1 U794 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n616), .Z(n191) );
  MUX2_X1 U795 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n616), .Z(n192) );
  MUX2_X1 U796 ( .A(n192), .B(n191), .S(n609), .Z(n193) );
  MUX2_X1 U797 ( .A(n193), .B(n190), .S(n606), .Z(n194) );
  MUX2_X1 U798 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U799 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n613), .Z(n196) );
  MUX2_X1 U800 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n611), .Z(n197) );
  MUX2_X1 U801 ( .A(n197), .B(n196), .S(n608), .Z(n198) );
  MUX2_X1 U802 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n617), .Z(n199) );
  MUX2_X1 U803 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n611), .Z(n200) );
  MUX2_X1 U804 ( .A(n200), .B(n199), .S(n609), .Z(n201) );
  MUX2_X1 U805 ( .A(n201), .B(n198), .S(n606), .Z(n202) );
  MUX2_X1 U806 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n611), .Z(n203) );
  MUX2_X1 U807 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n617), .Z(n204) );
  MUX2_X1 U808 ( .A(n204), .B(n203), .S(n608), .Z(n205) );
  MUX2_X1 U809 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n617), .Z(n206) );
  MUX2_X1 U810 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n617), .Z(n207) );
  MUX2_X1 U811 ( .A(n207), .B(n206), .S(n610), .Z(n208) );
  MUX2_X1 U812 ( .A(n208), .B(n205), .S(n607), .Z(n209) );
  MUX2_X1 U813 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U814 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U815 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n617), .Z(n211) );
  MUX2_X1 U816 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n612), .Z(n212) );
  MUX2_X1 U817 ( .A(n212), .B(n211), .S(n608), .Z(n213) );
  MUX2_X1 U818 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n614), .Z(n214) );
  MUX2_X1 U819 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n617), .Z(n215) );
  MUX2_X1 U820 ( .A(n215), .B(n214), .S(n608), .Z(n216) );
  MUX2_X1 U821 ( .A(n216), .B(n213), .S(n606), .Z(n217) );
  MUX2_X1 U822 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n613), .Z(n218) );
  MUX2_X1 U823 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n611), .Z(n219) );
  MUX2_X1 U824 ( .A(n219), .B(n218), .S(n608), .Z(n220) );
  MUX2_X1 U825 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n612), .Z(n221) );
  MUX2_X1 U826 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n222) );
  MUX2_X1 U827 ( .A(n222), .B(n221), .S(n610), .Z(n223) );
  MUX2_X1 U828 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U829 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U830 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n614), .Z(n226) );
  MUX2_X1 U831 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n612), .Z(n227) );
  MUX2_X1 U832 ( .A(n227), .B(n226), .S(n608), .Z(n228) );
  MUX2_X1 U833 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n611), .Z(n229) );
  MUX2_X1 U834 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n595) );
  MUX2_X1 U835 ( .A(n595), .B(n229), .S(N11), .Z(n596) );
  MUX2_X1 U836 ( .A(n596), .B(n228), .S(n607), .Z(n597) );
  MUX2_X1 U837 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n617), .Z(n598) );
  MUX2_X1 U838 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n614), .Z(n599) );
  MUX2_X1 U839 ( .A(n599), .B(n598), .S(n608), .Z(n600) );
  MUX2_X1 U840 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n617), .Z(n601) );
  MUX2_X1 U841 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n613), .Z(n602) );
  MUX2_X1 U842 ( .A(n602), .B(n601), .S(n608), .Z(n603) );
  MUX2_X1 U843 ( .A(n603), .B(n600), .S(n606), .Z(n604) );
  MUX2_X1 U844 ( .A(n604), .B(n597), .S(N13), .Z(n605) );
  MUX2_X1 U845 ( .A(n605), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U846 ( .A(N11), .Z(n608) );
  INV_X1 U847 ( .A(N10), .ZN(n618) );
  INV_X1 U848 ( .A(N11), .ZN(n619) );
  INV_X1 U849 ( .A(data_in[0]), .ZN(n620) );
  INV_X1 U850 ( .A(data_in[1]), .ZN(n621) );
  INV_X1 U851 ( .A(data_in[2]), .ZN(n622) );
  INV_X1 U852 ( .A(data_in[3]), .ZN(n623) );
  INV_X1 U853 ( .A(data_in[4]), .ZN(n624) );
  INV_X1 U854 ( .A(data_in[5]), .ZN(n625) );
  INV_X1 U855 ( .A(data_in[6]), .ZN(n626) );
  INV_X1 U856 ( .A(data_in[7]), .ZN(n627) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_10 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n633), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n634), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n635), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n636), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n637), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n638), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n639), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n640), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n641), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n642), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n643), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n644), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n645), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n646), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n647), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n648), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n649), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n650), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n651), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n652), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n653), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n654), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n655), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n656), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n657), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n658), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n659), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n660), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n661), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n662), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n663), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n664), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n665), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n666), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n667), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n668), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n669), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n670), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n671), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n672), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n673), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n674), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n675), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n676), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n677), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n678), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n679), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n680), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n681), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n682), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n683), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n684), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n685), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n686), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n687), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n688), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n689), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n690), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n691), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n692), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n693), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n694), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n695), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n696), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n697), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n698), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n699), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n700), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n701), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n702), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n703), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n704), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n705), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n706), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n707), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n708), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n709), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n710), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n711), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n712), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n713), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n714), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n715), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n716), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n717), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n718), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n719), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n720), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n721), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n722), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n723), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n724), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n725), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n726), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n727), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n728), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n729), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n730), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n731), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n732), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n733), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n734), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n735), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n736), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n737), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n738), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n739), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n740), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n741), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n742), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n743), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n744), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n745), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n746), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n747), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n748), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n749), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n750), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n751), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n752), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n753), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n754), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n755), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n756), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n757), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n758), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n759), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n760), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n761), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n762), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n763), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n764), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n765), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n766), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n767), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n768), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n769), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n770), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n771), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n772), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n773), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n774), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n775), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n776), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n777), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n778), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n779), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n780), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n781), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n782), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n783), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n784), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n785), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n786), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n787), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n788), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n789), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n790), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n791), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n792), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n793), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n794), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n795), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n796), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n797), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n798), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n799), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n800), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n801), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n802), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n803), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n804), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n805), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n806), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n807), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n808), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n809), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n810), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n811), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n812), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n813), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n814), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n815), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n816), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n817), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n818), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n819), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n820), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n821), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n822), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n823), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n824), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n852), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n853), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n854), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n855), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n856), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n857), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n858), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n859), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n860), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n861), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n862), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n863), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n864), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n865), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n866), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n867), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n868), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n869), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n870), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n871), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n872), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n873), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n874), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n875), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n876), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n877), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n878), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n879), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n880), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n881), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n882), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n883), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n884), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n885), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n886), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n887), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n888), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n889), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n890), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n891), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n892), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n893), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n894), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n895), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n896), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n897), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n898), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n899), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n900), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n901), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n902), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n903), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n904), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n905), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n906), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n907), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n908), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n909), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n910), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n911), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n912), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n913), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n914), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n915), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n2) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(N10), .Z(n621) );
  CLKBUF_X1 U4 ( .A(n621), .Z(n615) );
  CLKBUF_X1 U5 ( .A(n621), .Z(n616) );
  BUF_X1 U6 ( .A(n621), .Z(n614) );
  CLKBUF_X1 U7 ( .A(N11), .Z(n612) );
  INV_X2 U8 ( .A(n2), .ZN(data_out[3]) );
  BUF_X1 U9 ( .A(n622), .Z(n619) );
  BUF_X1 U10 ( .A(n622), .Z(n620) );
  BUF_X1 U11 ( .A(n621), .Z(n617) );
  BUF_X1 U12 ( .A(n621), .Z(n618) );
  BUF_X1 U13 ( .A(N11), .Z(n613) );
  BUF_X1 U14 ( .A(N10), .Z(n622) );
  NOR3_X1 U15 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1207) );
  NOR3_X1 U16 ( .A1(N11), .A2(N12), .A3(n623), .ZN(n1196) );
  NOR3_X1 U17 ( .A1(N10), .A2(N12), .A3(n624), .ZN(n1186) );
  NOR3_X1 U18 ( .A1(n623), .A2(N12), .A3(n624), .ZN(n1176) );
  INV_X1 U19 ( .A(n1133), .ZN(n848) );
  INV_X1 U20 ( .A(n1123), .ZN(n847) );
  INV_X1 U21 ( .A(n1114), .ZN(n846) );
  INV_X1 U22 ( .A(n1105), .ZN(n845) );
  INV_X1 U23 ( .A(n1060), .ZN(n840) );
  INV_X1 U24 ( .A(n1050), .ZN(n839) );
  INV_X1 U25 ( .A(n1041), .ZN(n838) );
  INV_X1 U26 ( .A(n1032), .ZN(n837) );
  INV_X1 U27 ( .A(n987), .ZN(n832) );
  INV_X1 U28 ( .A(n977), .ZN(n831) );
  INV_X1 U29 ( .A(n968), .ZN(n830) );
  INV_X1 U30 ( .A(n959), .ZN(n829) );
  INV_X1 U31 ( .A(n950), .ZN(n828) );
  INV_X1 U32 ( .A(n941), .ZN(n827) );
  INV_X1 U33 ( .A(n932), .ZN(n826) );
  INV_X1 U34 ( .A(n923), .ZN(n825) );
  INV_X1 U35 ( .A(n1096), .ZN(n844) );
  INV_X1 U36 ( .A(n1087), .ZN(n843) );
  INV_X1 U37 ( .A(n1078), .ZN(n842) );
  INV_X1 U38 ( .A(n1069), .ZN(n841) );
  INV_X1 U39 ( .A(n1023), .ZN(n836) );
  INV_X1 U40 ( .A(n1014), .ZN(n835) );
  INV_X1 U41 ( .A(n1005), .ZN(n834) );
  INV_X1 U42 ( .A(n996), .ZN(n833) );
  BUF_X1 U43 ( .A(N12), .Z(n609) );
  BUF_X1 U44 ( .A(N12), .Z(n610) );
  INV_X1 U45 ( .A(N13), .ZN(n850) );
  AND3_X1 U46 ( .A1(n623), .A2(n624), .A3(N12), .ZN(n1166) );
  AND3_X1 U47 ( .A1(N10), .A2(n624), .A3(N12), .ZN(n1156) );
  AND3_X1 U48 ( .A1(N11), .A2(n623), .A3(N12), .ZN(n1146) );
  AND3_X1 U49 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1136) );
  INV_X1 U50 ( .A(N14), .ZN(n851) );
  NAND2_X1 U51 ( .A1(n1196), .A2(n1206), .ZN(n1205) );
  NAND2_X1 U52 ( .A1(n1186), .A2(n1206), .ZN(n1195) );
  NAND2_X1 U53 ( .A1(n1176), .A2(n1206), .ZN(n1185) );
  NAND2_X1 U54 ( .A1(n1166), .A2(n1206), .ZN(n1175) );
  NAND2_X1 U55 ( .A1(n1156), .A2(n1206), .ZN(n1165) );
  NAND2_X1 U56 ( .A1(n1146), .A2(n1206), .ZN(n1155) );
  NAND2_X1 U57 ( .A1(n1136), .A2(n1206), .ZN(n1145) );
  NAND2_X1 U58 ( .A1(n1207), .A2(n1206), .ZN(n1216) );
  NAND2_X1 U59 ( .A1(n1125), .A2(n1207), .ZN(n1133) );
  NAND2_X1 U60 ( .A1(n1125), .A2(n1196), .ZN(n1123) );
  NAND2_X1 U61 ( .A1(n1125), .A2(n1186), .ZN(n1114) );
  NAND2_X1 U62 ( .A1(n1125), .A2(n1176), .ZN(n1105) );
  NAND2_X1 U63 ( .A1(n1052), .A2(n1207), .ZN(n1060) );
  NAND2_X1 U64 ( .A1(n1052), .A2(n1196), .ZN(n1050) );
  NAND2_X1 U65 ( .A1(n1052), .A2(n1186), .ZN(n1041) );
  NAND2_X1 U66 ( .A1(n1052), .A2(n1176), .ZN(n1032) );
  NAND2_X1 U67 ( .A1(n979), .A2(n1207), .ZN(n987) );
  NAND2_X1 U68 ( .A1(n979), .A2(n1196), .ZN(n977) );
  NAND2_X1 U69 ( .A1(n979), .A2(n1186), .ZN(n968) );
  NAND2_X1 U70 ( .A1(n979), .A2(n1176), .ZN(n959) );
  NAND2_X1 U71 ( .A1(n1125), .A2(n1166), .ZN(n1096) );
  NAND2_X1 U72 ( .A1(n1125), .A2(n1156), .ZN(n1087) );
  NAND2_X1 U73 ( .A1(n1125), .A2(n1146), .ZN(n1078) );
  NAND2_X1 U74 ( .A1(n1125), .A2(n1136), .ZN(n1069) );
  NAND2_X1 U75 ( .A1(n1052), .A2(n1166), .ZN(n1023) );
  NAND2_X1 U76 ( .A1(n1052), .A2(n1156), .ZN(n1014) );
  NAND2_X1 U77 ( .A1(n1052), .A2(n1146), .ZN(n1005) );
  NAND2_X1 U78 ( .A1(n1052), .A2(n1136), .ZN(n996) );
  NAND2_X1 U79 ( .A1(n979), .A2(n1166), .ZN(n950) );
  NAND2_X1 U80 ( .A1(n979), .A2(n1156), .ZN(n941) );
  NAND2_X1 U81 ( .A1(n979), .A2(n1146), .ZN(n932) );
  NAND2_X1 U82 ( .A1(n979), .A2(n1136), .ZN(n923) );
  AND3_X1 U83 ( .A1(n850), .A2(n851), .A3(n1135), .ZN(n1206) );
  AND3_X1 U84 ( .A1(N13), .A2(n1135), .A3(N14), .ZN(n979) );
  AND3_X1 U85 ( .A1(n1135), .A2(n851), .A3(N13), .ZN(n1125) );
  AND3_X1 U86 ( .A1(n1135), .A2(n850), .A3(N14), .ZN(n1052) );
  NOR2_X1 U87 ( .A1(n849), .A2(addr[5]), .ZN(n1135) );
  INV_X1 U88 ( .A(wr_en), .ZN(n849) );
  OAI21_X1 U89 ( .B1(n625), .B2(n1175), .A(n1174), .ZN(n883) );
  NAND2_X1 U90 ( .A1(\mem[4][0] ), .A2(n1175), .ZN(n1174) );
  OAI21_X1 U91 ( .B1(n626), .B2(n1175), .A(n1173), .ZN(n882) );
  NAND2_X1 U92 ( .A1(\mem[4][1] ), .A2(n1175), .ZN(n1173) );
  OAI21_X1 U93 ( .B1(n627), .B2(n1175), .A(n1172), .ZN(n881) );
  NAND2_X1 U94 ( .A1(\mem[4][2] ), .A2(n1175), .ZN(n1172) );
  OAI21_X1 U95 ( .B1(n628), .B2(n1175), .A(n1171), .ZN(n880) );
  NAND2_X1 U96 ( .A1(\mem[4][3] ), .A2(n1175), .ZN(n1171) );
  OAI21_X1 U97 ( .B1(n629), .B2(n1175), .A(n1170), .ZN(n879) );
  NAND2_X1 U98 ( .A1(\mem[4][4] ), .A2(n1175), .ZN(n1170) );
  OAI21_X1 U99 ( .B1(n630), .B2(n1175), .A(n1169), .ZN(n878) );
  NAND2_X1 U100 ( .A1(\mem[4][5] ), .A2(n1175), .ZN(n1169) );
  OAI21_X1 U101 ( .B1(n631), .B2(n1175), .A(n1168), .ZN(n877) );
  NAND2_X1 U102 ( .A1(\mem[4][6] ), .A2(n1175), .ZN(n1168) );
  OAI21_X1 U103 ( .B1(n632), .B2(n1175), .A(n1167), .ZN(n876) );
  NAND2_X1 U104 ( .A1(\mem[4][7] ), .A2(n1175), .ZN(n1167) );
  OAI21_X1 U105 ( .B1(n625), .B2(n1155), .A(n1154), .ZN(n867) );
  NAND2_X1 U106 ( .A1(\mem[6][0] ), .A2(n1155), .ZN(n1154) );
  OAI21_X1 U107 ( .B1(n626), .B2(n1155), .A(n1153), .ZN(n866) );
  NAND2_X1 U108 ( .A1(\mem[6][1] ), .A2(n1155), .ZN(n1153) );
  OAI21_X1 U109 ( .B1(n627), .B2(n1155), .A(n1152), .ZN(n865) );
  NAND2_X1 U110 ( .A1(\mem[6][2] ), .A2(n1155), .ZN(n1152) );
  OAI21_X1 U111 ( .B1(n628), .B2(n1155), .A(n1151), .ZN(n864) );
  NAND2_X1 U112 ( .A1(\mem[6][3] ), .A2(n1155), .ZN(n1151) );
  OAI21_X1 U113 ( .B1(n629), .B2(n1155), .A(n1150), .ZN(n863) );
  NAND2_X1 U114 ( .A1(\mem[6][4] ), .A2(n1155), .ZN(n1150) );
  OAI21_X1 U115 ( .B1(n630), .B2(n1155), .A(n1149), .ZN(n862) );
  NAND2_X1 U116 ( .A1(\mem[6][5] ), .A2(n1155), .ZN(n1149) );
  OAI21_X1 U117 ( .B1(n631), .B2(n1155), .A(n1148), .ZN(n861) );
  NAND2_X1 U118 ( .A1(\mem[6][6] ), .A2(n1155), .ZN(n1148) );
  OAI21_X1 U119 ( .B1(n632), .B2(n1155), .A(n1147), .ZN(n860) );
  NAND2_X1 U120 ( .A1(\mem[6][7] ), .A2(n1155), .ZN(n1147) );
  OAI21_X1 U121 ( .B1(n625), .B2(n1145), .A(n1144), .ZN(n859) );
  NAND2_X1 U122 ( .A1(\mem[7][0] ), .A2(n1145), .ZN(n1144) );
  OAI21_X1 U123 ( .B1(n626), .B2(n1145), .A(n1143), .ZN(n858) );
  NAND2_X1 U124 ( .A1(\mem[7][1] ), .A2(n1145), .ZN(n1143) );
  OAI21_X1 U125 ( .B1(n627), .B2(n1145), .A(n1142), .ZN(n857) );
  NAND2_X1 U126 ( .A1(\mem[7][2] ), .A2(n1145), .ZN(n1142) );
  OAI21_X1 U127 ( .B1(n628), .B2(n1145), .A(n1141), .ZN(n856) );
  NAND2_X1 U128 ( .A1(\mem[7][3] ), .A2(n1145), .ZN(n1141) );
  OAI21_X1 U129 ( .B1(n629), .B2(n1145), .A(n1140), .ZN(n855) );
  NAND2_X1 U130 ( .A1(\mem[7][4] ), .A2(n1145), .ZN(n1140) );
  OAI21_X1 U131 ( .B1(n630), .B2(n1145), .A(n1139), .ZN(n854) );
  NAND2_X1 U132 ( .A1(\mem[7][5] ), .A2(n1145), .ZN(n1139) );
  OAI21_X1 U133 ( .B1(n631), .B2(n1145), .A(n1138), .ZN(n853) );
  NAND2_X1 U134 ( .A1(\mem[7][6] ), .A2(n1145), .ZN(n1138) );
  OAI21_X1 U135 ( .B1(n632), .B2(n1145), .A(n1137), .ZN(n852) );
  NAND2_X1 U136 ( .A1(\mem[7][7] ), .A2(n1145), .ZN(n1137) );
  OAI21_X1 U137 ( .B1(n625), .B2(n1205), .A(n1204), .ZN(n907) );
  NAND2_X1 U138 ( .A1(\mem[1][0] ), .A2(n1205), .ZN(n1204) );
  OAI21_X1 U139 ( .B1(n626), .B2(n1205), .A(n1203), .ZN(n906) );
  NAND2_X1 U140 ( .A1(\mem[1][1] ), .A2(n1205), .ZN(n1203) );
  OAI21_X1 U141 ( .B1(n627), .B2(n1205), .A(n1202), .ZN(n905) );
  NAND2_X1 U142 ( .A1(\mem[1][2] ), .A2(n1205), .ZN(n1202) );
  OAI21_X1 U143 ( .B1(n628), .B2(n1205), .A(n1201), .ZN(n904) );
  NAND2_X1 U144 ( .A1(\mem[1][3] ), .A2(n1205), .ZN(n1201) );
  OAI21_X1 U145 ( .B1(n629), .B2(n1205), .A(n1200), .ZN(n903) );
  NAND2_X1 U146 ( .A1(\mem[1][4] ), .A2(n1205), .ZN(n1200) );
  OAI21_X1 U147 ( .B1(n630), .B2(n1205), .A(n1199), .ZN(n902) );
  NAND2_X1 U148 ( .A1(\mem[1][5] ), .A2(n1205), .ZN(n1199) );
  OAI21_X1 U149 ( .B1(n631), .B2(n1205), .A(n1198), .ZN(n901) );
  NAND2_X1 U150 ( .A1(\mem[1][6] ), .A2(n1205), .ZN(n1198) );
  OAI21_X1 U151 ( .B1(n632), .B2(n1205), .A(n1197), .ZN(n900) );
  NAND2_X1 U152 ( .A1(\mem[1][7] ), .A2(n1205), .ZN(n1197) );
  OAI21_X1 U153 ( .B1(n625), .B2(n1195), .A(n1194), .ZN(n899) );
  NAND2_X1 U154 ( .A1(\mem[2][0] ), .A2(n1195), .ZN(n1194) );
  OAI21_X1 U155 ( .B1(n626), .B2(n1195), .A(n1193), .ZN(n898) );
  NAND2_X1 U156 ( .A1(\mem[2][1] ), .A2(n1195), .ZN(n1193) );
  OAI21_X1 U157 ( .B1(n627), .B2(n1195), .A(n1192), .ZN(n897) );
  NAND2_X1 U158 ( .A1(\mem[2][2] ), .A2(n1195), .ZN(n1192) );
  OAI21_X1 U159 ( .B1(n628), .B2(n1195), .A(n1191), .ZN(n896) );
  NAND2_X1 U160 ( .A1(\mem[2][3] ), .A2(n1195), .ZN(n1191) );
  OAI21_X1 U161 ( .B1(n629), .B2(n1195), .A(n1190), .ZN(n895) );
  NAND2_X1 U162 ( .A1(\mem[2][4] ), .A2(n1195), .ZN(n1190) );
  OAI21_X1 U163 ( .B1(n630), .B2(n1195), .A(n1189), .ZN(n894) );
  NAND2_X1 U164 ( .A1(\mem[2][5] ), .A2(n1195), .ZN(n1189) );
  OAI21_X1 U165 ( .B1(n631), .B2(n1195), .A(n1188), .ZN(n893) );
  NAND2_X1 U166 ( .A1(\mem[2][6] ), .A2(n1195), .ZN(n1188) );
  OAI21_X1 U167 ( .B1(n632), .B2(n1195), .A(n1187), .ZN(n892) );
  NAND2_X1 U168 ( .A1(\mem[2][7] ), .A2(n1195), .ZN(n1187) );
  OAI21_X1 U169 ( .B1(n625), .B2(n1185), .A(n1184), .ZN(n891) );
  NAND2_X1 U170 ( .A1(\mem[3][0] ), .A2(n1185), .ZN(n1184) );
  OAI21_X1 U171 ( .B1(n626), .B2(n1185), .A(n1183), .ZN(n890) );
  NAND2_X1 U172 ( .A1(\mem[3][1] ), .A2(n1185), .ZN(n1183) );
  OAI21_X1 U173 ( .B1(n627), .B2(n1185), .A(n1182), .ZN(n889) );
  NAND2_X1 U174 ( .A1(\mem[3][2] ), .A2(n1185), .ZN(n1182) );
  OAI21_X1 U175 ( .B1(n628), .B2(n1185), .A(n1181), .ZN(n888) );
  NAND2_X1 U176 ( .A1(\mem[3][3] ), .A2(n1185), .ZN(n1181) );
  OAI21_X1 U177 ( .B1(n629), .B2(n1185), .A(n1180), .ZN(n887) );
  NAND2_X1 U178 ( .A1(\mem[3][4] ), .A2(n1185), .ZN(n1180) );
  OAI21_X1 U179 ( .B1(n630), .B2(n1185), .A(n1179), .ZN(n886) );
  NAND2_X1 U180 ( .A1(\mem[3][5] ), .A2(n1185), .ZN(n1179) );
  OAI21_X1 U181 ( .B1(n631), .B2(n1185), .A(n1178), .ZN(n885) );
  NAND2_X1 U182 ( .A1(\mem[3][6] ), .A2(n1185), .ZN(n1178) );
  OAI21_X1 U183 ( .B1(n632), .B2(n1185), .A(n1177), .ZN(n884) );
  NAND2_X1 U184 ( .A1(\mem[3][7] ), .A2(n1185), .ZN(n1177) );
  OAI21_X1 U185 ( .B1(n625), .B2(n1165), .A(n1164), .ZN(n875) );
  NAND2_X1 U186 ( .A1(\mem[5][0] ), .A2(n1165), .ZN(n1164) );
  OAI21_X1 U187 ( .B1(n626), .B2(n1165), .A(n1163), .ZN(n874) );
  NAND2_X1 U188 ( .A1(\mem[5][1] ), .A2(n1165), .ZN(n1163) );
  OAI21_X1 U189 ( .B1(n627), .B2(n1165), .A(n1162), .ZN(n873) );
  NAND2_X1 U190 ( .A1(\mem[5][2] ), .A2(n1165), .ZN(n1162) );
  OAI21_X1 U191 ( .B1(n628), .B2(n1165), .A(n1161), .ZN(n872) );
  NAND2_X1 U192 ( .A1(\mem[5][3] ), .A2(n1165), .ZN(n1161) );
  OAI21_X1 U193 ( .B1(n629), .B2(n1165), .A(n1160), .ZN(n871) );
  NAND2_X1 U194 ( .A1(\mem[5][4] ), .A2(n1165), .ZN(n1160) );
  OAI21_X1 U195 ( .B1(n630), .B2(n1165), .A(n1159), .ZN(n870) );
  NAND2_X1 U196 ( .A1(\mem[5][5] ), .A2(n1165), .ZN(n1159) );
  OAI21_X1 U197 ( .B1(n631), .B2(n1165), .A(n1158), .ZN(n869) );
  NAND2_X1 U198 ( .A1(\mem[5][6] ), .A2(n1165), .ZN(n1158) );
  OAI21_X1 U199 ( .B1(n632), .B2(n1165), .A(n1157), .ZN(n868) );
  NAND2_X1 U200 ( .A1(\mem[5][7] ), .A2(n1165), .ZN(n1157) );
  OAI21_X1 U201 ( .B1(n1216), .B2(n625), .A(n1215), .ZN(n915) );
  NAND2_X1 U202 ( .A1(\mem[0][0] ), .A2(n1216), .ZN(n1215) );
  OAI21_X1 U203 ( .B1(n1216), .B2(n626), .A(n1214), .ZN(n914) );
  NAND2_X1 U204 ( .A1(\mem[0][1] ), .A2(n1216), .ZN(n1214) );
  OAI21_X1 U205 ( .B1(n1216), .B2(n627), .A(n1213), .ZN(n913) );
  NAND2_X1 U206 ( .A1(\mem[0][2] ), .A2(n1216), .ZN(n1213) );
  OAI21_X1 U207 ( .B1(n1216), .B2(n628), .A(n1212), .ZN(n912) );
  NAND2_X1 U208 ( .A1(\mem[0][3] ), .A2(n1216), .ZN(n1212) );
  OAI21_X1 U209 ( .B1(n1216), .B2(n629), .A(n1211), .ZN(n911) );
  NAND2_X1 U210 ( .A1(\mem[0][4] ), .A2(n1216), .ZN(n1211) );
  OAI21_X1 U211 ( .B1(n1216), .B2(n630), .A(n1210), .ZN(n910) );
  NAND2_X1 U212 ( .A1(\mem[0][5] ), .A2(n1216), .ZN(n1210) );
  OAI21_X1 U213 ( .B1(n1216), .B2(n631), .A(n1209), .ZN(n909) );
  NAND2_X1 U214 ( .A1(\mem[0][6] ), .A2(n1216), .ZN(n1209) );
  OAI21_X1 U215 ( .B1(n1216), .B2(n632), .A(n1208), .ZN(n908) );
  NAND2_X1 U216 ( .A1(\mem[0][7] ), .A2(n1216), .ZN(n1208) );
  INV_X1 U217 ( .A(n1134), .ZN(n824) );
  AOI22_X1 U218 ( .A1(data_in[0]), .A2(n848), .B1(n1133), .B2(\mem[8][0] ), 
        .ZN(n1134) );
  INV_X1 U219 ( .A(n1132), .ZN(n823) );
  AOI22_X1 U220 ( .A1(data_in[1]), .A2(n848), .B1(n1133), .B2(\mem[8][1] ), 
        .ZN(n1132) );
  INV_X1 U221 ( .A(n1131), .ZN(n822) );
  AOI22_X1 U222 ( .A1(data_in[2]), .A2(n848), .B1(n1133), .B2(\mem[8][2] ), 
        .ZN(n1131) );
  INV_X1 U223 ( .A(n1130), .ZN(n821) );
  AOI22_X1 U224 ( .A1(data_in[3]), .A2(n848), .B1(n1133), .B2(\mem[8][3] ), 
        .ZN(n1130) );
  INV_X1 U225 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U226 ( .A1(data_in[4]), .A2(n848), .B1(n1133), .B2(\mem[8][4] ), 
        .ZN(n1129) );
  INV_X1 U227 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U228 ( .A1(data_in[5]), .A2(n848), .B1(n1133), .B2(\mem[8][5] ), 
        .ZN(n1128) );
  INV_X1 U229 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U230 ( .A1(data_in[6]), .A2(n848), .B1(n1133), .B2(\mem[8][6] ), 
        .ZN(n1127) );
  INV_X1 U231 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U232 ( .A1(data_in[7]), .A2(n848), .B1(n1133), .B2(\mem[8][7] ), 
        .ZN(n1126) );
  INV_X1 U233 ( .A(n1124), .ZN(n816) );
  AOI22_X1 U234 ( .A1(data_in[0]), .A2(n847), .B1(n1123), .B2(\mem[9][0] ), 
        .ZN(n1124) );
  INV_X1 U235 ( .A(n1122), .ZN(n815) );
  AOI22_X1 U236 ( .A1(data_in[1]), .A2(n847), .B1(n1123), .B2(\mem[9][1] ), 
        .ZN(n1122) );
  INV_X1 U237 ( .A(n1121), .ZN(n814) );
  AOI22_X1 U238 ( .A1(data_in[2]), .A2(n847), .B1(n1123), .B2(\mem[9][2] ), 
        .ZN(n1121) );
  INV_X1 U239 ( .A(n1120), .ZN(n813) );
  AOI22_X1 U240 ( .A1(data_in[3]), .A2(n847), .B1(n1123), .B2(\mem[9][3] ), 
        .ZN(n1120) );
  INV_X1 U241 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U242 ( .A1(data_in[4]), .A2(n847), .B1(n1123), .B2(\mem[9][4] ), 
        .ZN(n1119) );
  INV_X1 U243 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U244 ( .A1(data_in[5]), .A2(n847), .B1(n1123), .B2(\mem[9][5] ), 
        .ZN(n1118) );
  INV_X1 U245 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U246 ( .A1(data_in[6]), .A2(n847), .B1(n1123), .B2(\mem[9][6] ), 
        .ZN(n1117) );
  INV_X1 U247 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U248 ( .A1(data_in[7]), .A2(n847), .B1(n1123), .B2(\mem[9][7] ), 
        .ZN(n1116) );
  INV_X1 U249 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U250 ( .A1(data_in[0]), .A2(n846), .B1(n1114), .B2(\mem[10][0] ), 
        .ZN(n1115) );
  INV_X1 U251 ( .A(n1113), .ZN(n807) );
  AOI22_X1 U252 ( .A1(data_in[1]), .A2(n846), .B1(n1114), .B2(\mem[10][1] ), 
        .ZN(n1113) );
  INV_X1 U253 ( .A(n1112), .ZN(n806) );
  AOI22_X1 U254 ( .A1(data_in[2]), .A2(n846), .B1(n1114), .B2(\mem[10][2] ), 
        .ZN(n1112) );
  INV_X1 U255 ( .A(n1111), .ZN(n805) );
  AOI22_X1 U256 ( .A1(data_in[3]), .A2(n846), .B1(n1114), .B2(\mem[10][3] ), 
        .ZN(n1111) );
  INV_X1 U257 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U258 ( .A1(data_in[4]), .A2(n846), .B1(n1114), .B2(\mem[10][4] ), 
        .ZN(n1110) );
  INV_X1 U259 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U260 ( .A1(data_in[5]), .A2(n846), .B1(n1114), .B2(\mem[10][5] ), 
        .ZN(n1109) );
  INV_X1 U261 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U262 ( .A1(data_in[6]), .A2(n846), .B1(n1114), .B2(\mem[10][6] ), 
        .ZN(n1108) );
  INV_X1 U263 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U264 ( .A1(data_in[7]), .A2(n846), .B1(n1114), .B2(\mem[10][7] ), 
        .ZN(n1107) );
  INV_X1 U265 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U266 ( .A1(data_in[0]), .A2(n845), .B1(n1105), .B2(\mem[11][0] ), 
        .ZN(n1106) );
  INV_X1 U267 ( .A(n1104), .ZN(n799) );
  AOI22_X1 U268 ( .A1(data_in[1]), .A2(n845), .B1(n1105), .B2(\mem[11][1] ), 
        .ZN(n1104) );
  INV_X1 U269 ( .A(n1103), .ZN(n798) );
  AOI22_X1 U270 ( .A1(data_in[2]), .A2(n845), .B1(n1105), .B2(\mem[11][2] ), 
        .ZN(n1103) );
  INV_X1 U271 ( .A(n1102), .ZN(n797) );
  AOI22_X1 U272 ( .A1(data_in[3]), .A2(n845), .B1(n1105), .B2(\mem[11][3] ), 
        .ZN(n1102) );
  INV_X1 U273 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U274 ( .A1(data_in[4]), .A2(n845), .B1(n1105), .B2(\mem[11][4] ), 
        .ZN(n1101) );
  INV_X1 U275 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U276 ( .A1(data_in[5]), .A2(n845), .B1(n1105), .B2(\mem[11][5] ), 
        .ZN(n1100) );
  INV_X1 U277 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U278 ( .A1(data_in[6]), .A2(n845), .B1(n1105), .B2(\mem[11][6] ), 
        .ZN(n1099) );
  INV_X1 U279 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U280 ( .A1(data_in[7]), .A2(n845), .B1(n1105), .B2(\mem[11][7] ), 
        .ZN(n1098) );
  INV_X1 U281 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U282 ( .A1(data_in[0]), .A2(n844), .B1(n1096), .B2(\mem[12][0] ), 
        .ZN(n1097) );
  INV_X1 U283 ( .A(n1095), .ZN(n791) );
  AOI22_X1 U284 ( .A1(data_in[1]), .A2(n844), .B1(n1096), .B2(\mem[12][1] ), 
        .ZN(n1095) );
  INV_X1 U285 ( .A(n1094), .ZN(n790) );
  AOI22_X1 U286 ( .A1(data_in[2]), .A2(n844), .B1(n1096), .B2(\mem[12][2] ), 
        .ZN(n1094) );
  INV_X1 U287 ( .A(n1093), .ZN(n789) );
  AOI22_X1 U288 ( .A1(data_in[3]), .A2(n844), .B1(n1096), .B2(\mem[12][3] ), 
        .ZN(n1093) );
  INV_X1 U289 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U290 ( .A1(data_in[4]), .A2(n844), .B1(n1096), .B2(\mem[12][4] ), 
        .ZN(n1092) );
  INV_X1 U291 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U292 ( .A1(data_in[5]), .A2(n844), .B1(n1096), .B2(\mem[12][5] ), 
        .ZN(n1091) );
  INV_X1 U293 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U294 ( .A1(data_in[6]), .A2(n844), .B1(n1096), .B2(\mem[12][6] ), 
        .ZN(n1090) );
  INV_X1 U295 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U296 ( .A1(data_in[7]), .A2(n844), .B1(n1096), .B2(\mem[12][7] ), 
        .ZN(n1089) );
  INV_X1 U297 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U298 ( .A1(data_in[0]), .A2(n843), .B1(n1087), .B2(\mem[13][0] ), 
        .ZN(n1088) );
  INV_X1 U299 ( .A(n1086), .ZN(n783) );
  AOI22_X1 U300 ( .A1(data_in[1]), .A2(n843), .B1(n1087), .B2(\mem[13][1] ), 
        .ZN(n1086) );
  INV_X1 U301 ( .A(n1085), .ZN(n782) );
  AOI22_X1 U302 ( .A1(data_in[2]), .A2(n843), .B1(n1087), .B2(\mem[13][2] ), 
        .ZN(n1085) );
  INV_X1 U303 ( .A(n1084), .ZN(n781) );
  AOI22_X1 U304 ( .A1(data_in[3]), .A2(n843), .B1(n1087), .B2(\mem[13][3] ), 
        .ZN(n1084) );
  INV_X1 U305 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U306 ( .A1(data_in[4]), .A2(n843), .B1(n1087), .B2(\mem[13][4] ), 
        .ZN(n1083) );
  INV_X1 U307 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U308 ( .A1(data_in[5]), .A2(n843), .B1(n1087), .B2(\mem[13][5] ), 
        .ZN(n1082) );
  INV_X1 U309 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U310 ( .A1(data_in[6]), .A2(n843), .B1(n1087), .B2(\mem[13][6] ), 
        .ZN(n1081) );
  INV_X1 U311 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U312 ( .A1(data_in[7]), .A2(n843), .B1(n1087), .B2(\mem[13][7] ), 
        .ZN(n1080) );
  INV_X1 U313 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U314 ( .A1(data_in[0]), .A2(n842), .B1(n1078), .B2(\mem[14][0] ), 
        .ZN(n1079) );
  INV_X1 U315 ( .A(n1077), .ZN(n775) );
  AOI22_X1 U316 ( .A1(data_in[1]), .A2(n842), .B1(n1078), .B2(\mem[14][1] ), 
        .ZN(n1077) );
  INV_X1 U317 ( .A(n1076), .ZN(n774) );
  AOI22_X1 U318 ( .A1(data_in[2]), .A2(n842), .B1(n1078), .B2(\mem[14][2] ), 
        .ZN(n1076) );
  INV_X1 U319 ( .A(n1075), .ZN(n773) );
  AOI22_X1 U320 ( .A1(data_in[3]), .A2(n842), .B1(n1078), .B2(\mem[14][3] ), 
        .ZN(n1075) );
  INV_X1 U321 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U322 ( .A1(data_in[4]), .A2(n842), .B1(n1078), .B2(\mem[14][4] ), 
        .ZN(n1074) );
  INV_X1 U323 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U324 ( .A1(data_in[5]), .A2(n842), .B1(n1078), .B2(\mem[14][5] ), 
        .ZN(n1073) );
  INV_X1 U325 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U326 ( .A1(data_in[6]), .A2(n842), .B1(n1078), .B2(\mem[14][6] ), 
        .ZN(n1072) );
  INV_X1 U327 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U328 ( .A1(data_in[7]), .A2(n842), .B1(n1078), .B2(\mem[14][7] ), 
        .ZN(n1071) );
  INV_X1 U329 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U330 ( .A1(data_in[0]), .A2(n841), .B1(n1069), .B2(\mem[15][0] ), 
        .ZN(n1070) );
  INV_X1 U331 ( .A(n1068), .ZN(n767) );
  AOI22_X1 U332 ( .A1(data_in[1]), .A2(n841), .B1(n1069), .B2(\mem[15][1] ), 
        .ZN(n1068) );
  INV_X1 U333 ( .A(n1067), .ZN(n766) );
  AOI22_X1 U334 ( .A1(data_in[2]), .A2(n841), .B1(n1069), .B2(\mem[15][2] ), 
        .ZN(n1067) );
  INV_X1 U335 ( .A(n1066), .ZN(n765) );
  AOI22_X1 U336 ( .A1(data_in[3]), .A2(n841), .B1(n1069), .B2(\mem[15][3] ), 
        .ZN(n1066) );
  INV_X1 U337 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U338 ( .A1(data_in[4]), .A2(n841), .B1(n1069), .B2(\mem[15][4] ), 
        .ZN(n1065) );
  INV_X1 U339 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U340 ( .A1(data_in[5]), .A2(n841), .B1(n1069), .B2(\mem[15][5] ), 
        .ZN(n1064) );
  INV_X1 U341 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U342 ( .A1(data_in[6]), .A2(n841), .B1(n1069), .B2(\mem[15][6] ), 
        .ZN(n1063) );
  INV_X1 U343 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U344 ( .A1(data_in[7]), .A2(n841), .B1(n1069), .B2(\mem[15][7] ), 
        .ZN(n1062) );
  INV_X1 U345 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U346 ( .A1(data_in[0]), .A2(n840), .B1(n1060), .B2(\mem[16][0] ), 
        .ZN(n1061) );
  INV_X1 U347 ( .A(n1059), .ZN(n759) );
  AOI22_X1 U348 ( .A1(data_in[1]), .A2(n840), .B1(n1060), .B2(\mem[16][1] ), 
        .ZN(n1059) );
  INV_X1 U349 ( .A(n1058), .ZN(n758) );
  AOI22_X1 U350 ( .A1(data_in[2]), .A2(n840), .B1(n1060), .B2(\mem[16][2] ), 
        .ZN(n1058) );
  INV_X1 U351 ( .A(n1057), .ZN(n757) );
  AOI22_X1 U352 ( .A1(data_in[3]), .A2(n840), .B1(n1060), .B2(\mem[16][3] ), 
        .ZN(n1057) );
  INV_X1 U353 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U354 ( .A1(data_in[4]), .A2(n840), .B1(n1060), .B2(\mem[16][4] ), 
        .ZN(n1056) );
  INV_X1 U355 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U356 ( .A1(data_in[5]), .A2(n840), .B1(n1060), .B2(\mem[16][5] ), 
        .ZN(n1055) );
  INV_X1 U357 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U358 ( .A1(data_in[6]), .A2(n840), .B1(n1060), .B2(\mem[16][6] ), 
        .ZN(n1054) );
  INV_X1 U359 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U360 ( .A1(data_in[7]), .A2(n840), .B1(n1060), .B2(\mem[16][7] ), 
        .ZN(n1053) );
  INV_X1 U361 ( .A(n1051), .ZN(n752) );
  AOI22_X1 U362 ( .A1(data_in[0]), .A2(n839), .B1(n1050), .B2(\mem[17][0] ), 
        .ZN(n1051) );
  INV_X1 U363 ( .A(n1049), .ZN(n751) );
  AOI22_X1 U364 ( .A1(data_in[1]), .A2(n839), .B1(n1050), .B2(\mem[17][1] ), 
        .ZN(n1049) );
  INV_X1 U365 ( .A(n1048), .ZN(n750) );
  AOI22_X1 U366 ( .A1(data_in[2]), .A2(n839), .B1(n1050), .B2(\mem[17][2] ), 
        .ZN(n1048) );
  INV_X1 U367 ( .A(n1047), .ZN(n749) );
  AOI22_X1 U368 ( .A1(data_in[3]), .A2(n839), .B1(n1050), .B2(\mem[17][3] ), 
        .ZN(n1047) );
  INV_X1 U369 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U370 ( .A1(data_in[4]), .A2(n839), .B1(n1050), .B2(\mem[17][4] ), 
        .ZN(n1046) );
  INV_X1 U371 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U372 ( .A1(data_in[5]), .A2(n839), .B1(n1050), .B2(\mem[17][5] ), 
        .ZN(n1045) );
  INV_X1 U373 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U374 ( .A1(data_in[6]), .A2(n839), .B1(n1050), .B2(\mem[17][6] ), 
        .ZN(n1044) );
  INV_X1 U375 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U376 ( .A1(data_in[7]), .A2(n839), .B1(n1050), .B2(\mem[17][7] ), 
        .ZN(n1043) );
  INV_X1 U377 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U378 ( .A1(data_in[0]), .A2(n838), .B1(n1041), .B2(\mem[18][0] ), 
        .ZN(n1042) );
  INV_X1 U379 ( .A(n1040), .ZN(n743) );
  AOI22_X1 U380 ( .A1(data_in[1]), .A2(n838), .B1(n1041), .B2(\mem[18][1] ), 
        .ZN(n1040) );
  INV_X1 U381 ( .A(n1039), .ZN(n742) );
  AOI22_X1 U382 ( .A1(data_in[2]), .A2(n838), .B1(n1041), .B2(\mem[18][2] ), 
        .ZN(n1039) );
  INV_X1 U383 ( .A(n1038), .ZN(n741) );
  AOI22_X1 U384 ( .A1(data_in[3]), .A2(n838), .B1(n1041), .B2(\mem[18][3] ), 
        .ZN(n1038) );
  INV_X1 U385 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U386 ( .A1(data_in[4]), .A2(n838), .B1(n1041), .B2(\mem[18][4] ), 
        .ZN(n1037) );
  INV_X1 U387 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U388 ( .A1(data_in[5]), .A2(n838), .B1(n1041), .B2(\mem[18][5] ), 
        .ZN(n1036) );
  INV_X1 U389 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U390 ( .A1(data_in[6]), .A2(n838), .B1(n1041), .B2(\mem[18][6] ), 
        .ZN(n1035) );
  INV_X1 U391 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U392 ( .A1(data_in[7]), .A2(n838), .B1(n1041), .B2(\mem[18][7] ), 
        .ZN(n1034) );
  INV_X1 U393 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U394 ( .A1(data_in[0]), .A2(n837), .B1(n1032), .B2(\mem[19][0] ), 
        .ZN(n1033) );
  INV_X1 U395 ( .A(n1031), .ZN(n735) );
  AOI22_X1 U396 ( .A1(data_in[1]), .A2(n837), .B1(n1032), .B2(\mem[19][1] ), 
        .ZN(n1031) );
  INV_X1 U397 ( .A(n1030), .ZN(n734) );
  AOI22_X1 U398 ( .A1(data_in[2]), .A2(n837), .B1(n1032), .B2(\mem[19][2] ), 
        .ZN(n1030) );
  INV_X1 U399 ( .A(n1029), .ZN(n733) );
  AOI22_X1 U400 ( .A1(data_in[3]), .A2(n837), .B1(n1032), .B2(\mem[19][3] ), 
        .ZN(n1029) );
  INV_X1 U401 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U402 ( .A1(data_in[4]), .A2(n837), .B1(n1032), .B2(\mem[19][4] ), 
        .ZN(n1028) );
  INV_X1 U403 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U404 ( .A1(data_in[5]), .A2(n837), .B1(n1032), .B2(\mem[19][5] ), 
        .ZN(n1027) );
  INV_X1 U405 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U406 ( .A1(data_in[6]), .A2(n837), .B1(n1032), .B2(\mem[19][6] ), 
        .ZN(n1026) );
  INV_X1 U407 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U408 ( .A1(data_in[7]), .A2(n837), .B1(n1032), .B2(\mem[19][7] ), 
        .ZN(n1025) );
  INV_X1 U409 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U410 ( .A1(data_in[0]), .A2(n836), .B1(n1023), .B2(\mem[20][0] ), 
        .ZN(n1024) );
  INV_X1 U411 ( .A(n1022), .ZN(n727) );
  AOI22_X1 U412 ( .A1(data_in[1]), .A2(n836), .B1(n1023), .B2(\mem[20][1] ), 
        .ZN(n1022) );
  INV_X1 U413 ( .A(n1021), .ZN(n726) );
  AOI22_X1 U414 ( .A1(data_in[2]), .A2(n836), .B1(n1023), .B2(\mem[20][2] ), 
        .ZN(n1021) );
  INV_X1 U415 ( .A(n1020), .ZN(n725) );
  AOI22_X1 U416 ( .A1(data_in[3]), .A2(n836), .B1(n1023), .B2(\mem[20][3] ), 
        .ZN(n1020) );
  INV_X1 U417 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U418 ( .A1(data_in[4]), .A2(n836), .B1(n1023), .B2(\mem[20][4] ), 
        .ZN(n1019) );
  INV_X1 U419 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U420 ( .A1(data_in[5]), .A2(n836), .B1(n1023), .B2(\mem[20][5] ), 
        .ZN(n1018) );
  INV_X1 U421 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U422 ( .A1(data_in[6]), .A2(n836), .B1(n1023), .B2(\mem[20][6] ), 
        .ZN(n1017) );
  INV_X1 U423 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U424 ( .A1(data_in[7]), .A2(n836), .B1(n1023), .B2(\mem[20][7] ), 
        .ZN(n1016) );
  INV_X1 U425 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U426 ( .A1(data_in[0]), .A2(n835), .B1(n1014), .B2(\mem[21][0] ), 
        .ZN(n1015) );
  INV_X1 U427 ( .A(n1013), .ZN(n719) );
  AOI22_X1 U428 ( .A1(data_in[1]), .A2(n835), .B1(n1014), .B2(\mem[21][1] ), 
        .ZN(n1013) );
  INV_X1 U429 ( .A(n1012), .ZN(n718) );
  AOI22_X1 U430 ( .A1(data_in[2]), .A2(n835), .B1(n1014), .B2(\mem[21][2] ), 
        .ZN(n1012) );
  INV_X1 U431 ( .A(n1011), .ZN(n717) );
  AOI22_X1 U432 ( .A1(data_in[3]), .A2(n835), .B1(n1014), .B2(\mem[21][3] ), 
        .ZN(n1011) );
  INV_X1 U433 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U434 ( .A1(data_in[4]), .A2(n835), .B1(n1014), .B2(\mem[21][4] ), 
        .ZN(n1010) );
  INV_X1 U435 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U436 ( .A1(data_in[5]), .A2(n835), .B1(n1014), .B2(\mem[21][5] ), 
        .ZN(n1009) );
  INV_X1 U437 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U438 ( .A1(data_in[6]), .A2(n835), .B1(n1014), .B2(\mem[21][6] ), 
        .ZN(n1008) );
  INV_X1 U439 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U440 ( .A1(data_in[7]), .A2(n835), .B1(n1014), .B2(\mem[21][7] ), 
        .ZN(n1007) );
  INV_X1 U441 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U442 ( .A1(data_in[0]), .A2(n834), .B1(n1005), .B2(\mem[22][0] ), 
        .ZN(n1006) );
  INV_X1 U443 ( .A(n1004), .ZN(n711) );
  AOI22_X1 U444 ( .A1(data_in[1]), .A2(n834), .B1(n1005), .B2(\mem[22][1] ), 
        .ZN(n1004) );
  INV_X1 U445 ( .A(n1003), .ZN(n710) );
  AOI22_X1 U446 ( .A1(data_in[2]), .A2(n834), .B1(n1005), .B2(\mem[22][2] ), 
        .ZN(n1003) );
  INV_X1 U447 ( .A(n1002), .ZN(n709) );
  AOI22_X1 U448 ( .A1(data_in[3]), .A2(n834), .B1(n1005), .B2(\mem[22][3] ), 
        .ZN(n1002) );
  INV_X1 U449 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U450 ( .A1(data_in[4]), .A2(n834), .B1(n1005), .B2(\mem[22][4] ), 
        .ZN(n1001) );
  INV_X1 U451 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U452 ( .A1(data_in[5]), .A2(n834), .B1(n1005), .B2(\mem[22][5] ), 
        .ZN(n1000) );
  INV_X1 U453 ( .A(n999), .ZN(n706) );
  AOI22_X1 U454 ( .A1(data_in[6]), .A2(n834), .B1(n1005), .B2(\mem[22][6] ), 
        .ZN(n999) );
  INV_X1 U455 ( .A(n998), .ZN(n705) );
  AOI22_X1 U456 ( .A1(data_in[7]), .A2(n834), .B1(n1005), .B2(\mem[22][7] ), 
        .ZN(n998) );
  INV_X1 U457 ( .A(n997), .ZN(n704) );
  AOI22_X1 U458 ( .A1(data_in[0]), .A2(n833), .B1(n996), .B2(\mem[23][0] ), 
        .ZN(n997) );
  INV_X1 U459 ( .A(n995), .ZN(n703) );
  AOI22_X1 U460 ( .A1(data_in[1]), .A2(n833), .B1(n996), .B2(\mem[23][1] ), 
        .ZN(n995) );
  INV_X1 U461 ( .A(n994), .ZN(n702) );
  AOI22_X1 U462 ( .A1(data_in[2]), .A2(n833), .B1(n996), .B2(\mem[23][2] ), 
        .ZN(n994) );
  INV_X1 U463 ( .A(n993), .ZN(n701) );
  AOI22_X1 U464 ( .A1(data_in[3]), .A2(n833), .B1(n996), .B2(\mem[23][3] ), 
        .ZN(n993) );
  INV_X1 U465 ( .A(n992), .ZN(n700) );
  AOI22_X1 U466 ( .A1(data_in[4]), .A2(n833), .B1(n996), .B2(\mem[23][4] ), 
        .ZN(n992) );
  INV_X1 U467 ( .A(n991), .ZN(n699) );
  AOI22_X1 U468 ( .A1(data_in[5]), .A2(n833), .B1(n996), .B2(\mem[23][5] ), 
        .ZN(n991) );
  INV_X1 U469 ( .A(n990), .ZN(n698) );
  AOI22_X1 U470 ( .A1(data_in[6]), .A2(n833), .B1(n996), .B2(\mem[23][6] ), 
        .ZN(n990) );
  INV_X1 U471 ( .A(n989), .ZN(n697) );
  AOI22_X1 U472 ( .A1(data_in[7]), .A2(n833), .B1(n996), .B2(\mem[23][7] ), 
        .ZN(n989) );
  INV_X1 U473 ( .A(n988), .ZN(n696) );
  AOI22_X1 U474 ( .A1(data_in[0]), .A2(n832), .B1(n987), .B2(\mem[24][0] ), 
        .ZN(n988) );
  INV_X1 U475 ( .A(n986), .ZN(n695) );
  AOI22_X1 U476 ( .A1(data_in[1]), .A2(n832), .B1(n987), .B2(\mem[24][1] ), 
        .ZN(n986) );
  INV_X1 U477 ( .A(n985), .ZN(n694) );
  AOI22_X1 U478 ( .A1(data_in[2]), .A2(n832), .B1(n987), .B2(\mem[24][2] ), 
        .ZN(n985) );
  INV_X1 U479 ( .A(n984), .ZN(n693) );
  AOI22_X1 U480 ( .A1(data_in[3]), .A2(n832), .B1(n987), .B2(\mem[24][3] ), 
        .ZN(n984) );
  INV_X1 U481 ( .A(n983), .ZN(n692) );
  AOI22_X1 U482 ( .A1(data_in[4]), .A2(n832), .B1(n987), .B2(\mem[24][4] ), 
        .ZN(n983) );
  INV_X1 U483 ( .A(n982), .ZN(n691) );
  AOI22_X1 U484 ( .A1(data_in[5]), .A2(n832), .B1(n987), .B2(\mem[24][5] ), 
        .ZN(n982) );
  INV_X1 U485 ( .A(n981), .ZN(n690) );
  AOI22_X1 U486 ( .A1(data_in[6]), .A2(n832), .B1(n987), .B2(\mem[24][6] ), 
        .ZN(n981) );
  INV_X1 U487 ( .A(n980), .ZN(n689) );
  AOI22_X1 U488 ( .A1(data_in[7]), .A2(n832), .B1(n987), .B2(\mem[24][7] ), 
        .ZN(n980) );
  INV_X1 U489 ( .A(n978), .ZN(n688) );
  AOI22_X1 U490 ( .A1(data_in[0]), .A2(n831), .B1(n977), .B2(\mem[25][0] ), 
        .ZN(n978) );
  INV_X1 U491 ( .A(n976), .ZN(n687) );
  AOI22_X1 U492 ( .A1(data_in[1]), .A2(n831), .B1(n977), .B2(\mem[25][1] ), 
        .ZN(n976) );
  INV_X1 U493 ( .A(n975), .ZN(n686) );
  AOI22_X1 U494 ( .A1(data_in[2]), .A2(n831), .B1(n977), .B2(\mem[25][2] ), 
        .ZN(n975) );
  INV_X1 U495 ( .A(n974), .ZN(n685) );
  AOI22_X1 U496 ( .A1(data_in[3]), .A2(n831), .B1(n977), .B2(\mem[25][3] ), 
        .ZN(n974) );
  INV_X1 U497 ( .A(n973), .ZN(n684) );
  AOI22_X1 U498 ( .A1(data_in[4]), .A2(n831), .B1(n977), .B2(\mem[25][4] ), 
        .ZN(n973) );
  INV_X1 U499 ( .A(n972), .ZN(n683) );
  AOI22_X1 U500 ( .A1(data_in[5]), .A2(n831), .B1(n977), .B2(\mem[25][5] ), 
        .ZN(n972) );
  INV_X1 U501 ( .A(n971), .ZN(n682) );
  AOI22_X1 U502 ( .A1(data_in[6]), .A2(n831), .B1(n977), .B2(\mem[25][6] ), 
        .ZN(n971) );
  INV_X1 U503 ( .A(n970), .ZN(n681) );
  AOI22_X1 U504 ( .A1(data_in[7]), .A2(n831), .B1(n977), .B2(\mem[25][7] ), 
        .ZN(n970) );
  INV_X1 U505 ( .A(n969), .ZN(n680) );
  AOI22_X1 U506 ( .A1(data_in[0]), .A2(n830), .B1(n968), .B2(\mem[26][0] ), 
        .ZN(n969) );
  INV_X1 U507 ( .A(n967), .ZN(n679) );
  AOI22_X1 U508 ( .A1(data_in[1]), .A2(n830), .B1(n968), .B2(\mem[26][1] ), 
        .ZN(n967) );
  INV_X1 U509 ( .A(n966), .ZN(n678) );
  AOI22_X1 U510 ( .A1(data_in[2]), .A2(n830), .B1(n968), .B2(\mem[26][2] ), 
        .ZN(n966) );
  INV_X1 U511 ( .A(n965), .ZN(n677) );
  AOI22_X1 U512 ( .A1(data_in[3]), .A2(n830), .B1(n968), .B2(\mem[26][3] ), 
        .ZN(n965) );
  INV_X1 U513 ( .A(n964), .ZN(n676) );
  AOI22_X1 U514 ( .A1(data_in[4]), .A2(n830), .B1(n968), .B2(\mem[26][4] ), 
        .ZN(n964) );
  INV_X1 U515 ( .A(n963), .ZN(n675) );
  AOI22_X1 U516 ( .A1(data_in[5]), .A2(n830), .B1(n968), .B2(\mem[26][5] ), 
        .ZN(n963) );
  INV_X1 U517 ( .A(n962), .ZN(n674) );
  AOI22_X1 U518 ( .A1(data_in[6]), .A2(n830), .B1(n968), .B2(\mem[26][6] ), 
        .ZN(n962) );
  INV_X1 U519 ( .A(n961), .ZN(n673) );
  AOI22_X1 U520 ( .A1(data_in[7]), .A2(n830), .B1(n968), .B2(\mem[26][7] ), 
        .ZN(n961) );
  INV_X1 U521 ( .A(n960), .ZN(n672) );
  AOI22_X1 U522 ( .A1(data_in[0]), .A2(n829), .B1(n959), .B2(\mem[27][0] ), 
        .ZN(n960) );
  INV_X1 U523 ( .A(n958), .ZN(n671) );
  AOI22_X1 U524 ( .A1(data_in[1]), .A2(n829), .B1(n959), .B2(\mem[27][1] ), 
        .ZN(n958) );
  INV_X1 U525 ( .A(n957), .ZN(n670) );
  AOI22_X1 U526 ( .A1(data_in[2]), .A2(n829), .B1(n959), .B2(\mem[27][2] ), 
        .ZN(n957) );
  INV_X1 U527 ( .A(n956), .ZN(n669) );
  AOI22_X1 U528 ( .A1(data_in[3]), .A2(n829), .B1(n959), .B2(\mem[27][3] ), 
        .ZN(n956) );
  INV_X1 U529 ( .A(n955), .ZN(n668) );
  AOI22_X1 U530 ( .A1(data_in[4]), .A2(n829), .B1(n959), .B2(\mem[27][4] ), 
        .ZN(n955) );
  INV_X1 U531 ( .A(n954), .ZN(n667) );
  AOI22_X1 U532 ( .A1(data_in[5]), .A2(n829), .B1(n959), .B2(\mem[27][5] ), 
        .ZN(n954) );
  INV_X1 U533 ( .A(n953), .ZN(n666) );
  AOI22_X1 U534 ( .A1(data_in[6]), .A2(n829), .B1(n959), .B2(\mem[27][6] ), 
        .ZN(n953) );
  INV_X1 U535 ( .A(n952), .ZN(n665) );
  AOI22_X1 U536 ( .A1(data_in[7]), .A2(n829), .B1(n959), .B2(\mem[27][7] ), 
        .ZN(n952) );
  INV_X1 U537 ( .A(n951), .ZN(n664) );
  AOI22_X1 U538 ( .A1(data_in[0]), .A2(n828), .B1(n950), .B2(\mem[28][0] ), 
        .ZN(n951) );
  INV_X1 U539 ( .A(n949), .ZN(n663) );
  AOI22_X1 U540 ( .A1(data_in[1]), .A2(n828), .B1(n950), .B2(\mem[28][1] ), 
        .ZN(n949) );
  INV_X1 U541 ( .A(n948), .ZN(n662) );
  AOI22_X1 U542 ( .A1(data_in[2]), .A2(n828), .B1(n950), .B2(\mem[28][2] ), 
        .ZN(n948) );
  INV_X1 U543 ( .A(n947), .ZN(n661) );
  AOI22_X1 U544 ( .A1(data_in[3]), .A2(n828), .B1(n950), .B2(\mem[28][3] ), 
        .ZN(n947) );
  INV_X1 U545 ( .A(n946), .ZN(n660) );
  AOI22_X1 U546 ( .A1(data_in[4]), .A2(n828), .B1(n950), .B2(\mem[28][4] ), 
        .ZN(n946) );
  INV_X1 U547 ( .A(n945), .ZN(n659) );
  AOI22_X1 U548 ( .A1(data_in[5]), .A2(n828), .B1(n950), .B2(\mem[28][5] ), 
        .ZN(n945) );
  INV_X1 U549 ( .A(n944), .ZN(n658) );
  AOI22_X1 U550 ( .A1(data_in[6]), .A2(n828), .B1(n950), .B2(\mem[28][6] ), 
        .ZN(n944) );
  INV_X1 U551 ( .A(n943), .ZN(n657) );
  AOI22_X1 U552 ( .A1(data_in[7]), .A2(n828), .B1(n950), .B2(\mem[28][7] ), 
        .ZN(n943) );
  INV_X1 U553 ( .A(n942), .ZN(n656) );
  AOI22_X1 U554 ( .A1(data_in[0]), .A2(n827), .B1(n941), .B2(\mem[29][0] ), 
        .ZN(n942) );
  INV_X1 U555 ( .A(n940), .ZN(n655) );
  AOI22_X1 U556 ( .A1(data_in[1]), .A2(n827), .B1(n941), .B2(\mem[29][1] ), 
        .ZN(n940) );
  INV_X1 U557 ( .A(n939), .ZN(n654) );
  AOI22_X1 U558 ( .A1(data_in[2]), .A2(n827), .B1(n941), .B2(\mem[29][2] ), 
        .ZN(n939) );
  INV_X1 U559 ( .A(n938), .ZN(n653) );
  AOI22_X1 U560 ( .A1(data_in[3]), .A2(n827), .B1(n941), .B2(\mem[29][3] ), 
        .ZN(n938) );
  INV_X1 U561 ( .A(n937), .ZN(n652) );
  AOI22_X1 U562 ( .A1(data_in[4]), .A2(n827), .B1(n941), .B2(\mem[29][4] ), 
        .ZN(n937) );
  INV_X1 U563 ( .A(n936), .ZN(n651) );
  AOI22_X1 U564 ( .A1(data_in[5]), .A2(n827), .B1(n941), .B2(\mem[29][5] ), 
        .ZN(n936) );
  INV_X1 U565 ( .A(n935), .ZN(n650) );
  AOI22_X1 U566 ( .A1(data_in[6]), .A2(n827), .B1(n941), .B2(\mem[29][6] ), 
        .ZN(n935) );
  INV_X1 U567 ( .A(n934), .ZN(n649) );
  AOI22_X1 U568 ( .A1(data_in[7]), .A2(n827), .B1(n941), .B2(\mem[29][7] ), 
        .ZN(n934) );
  INV_X1 U569 ( .A(n933), .ZN(n648) );
  AOI22_X1 U570 ( .A1(data_in[0]), .A2(n826), .B1(n932), .B2(\mem[30][0] ), 
        .ZN(n933) );
  INV_X1 U571 ( .A(n931), .ZN(n647) );
  AOI22_X1 U572 ( .A1(data_in[1]), .A2(n826), .B1(n932), .B2(\mem[30][1] ), 
        .ZN(n931) );
  INV_X1 U573 ( .A(n930), .ZN(n646) );
  AOI22_X1 U574 ( .A1(data_in[2]), .A2(n826), .B1(n932), .B2(\mem[30][2] ), 
        .ZN(n930) );
  INV_X1 U575 ( .A(n929), .ZN(n645) );
  AOI22_X1 U576 ( .A1(data_in[3]), .A2(n826), .B1(n932), .B2(\mem[30][3] ), 
        .ZN(n929) );
  INV_X1 U577 ( .A(n928), .ZN(n644) );
  AOI22_X1 U578 ( .A1(data_in[4]), .A2(n826), .B1(n932), .B2(\mem[30][4] ), 
        .ZN(n928) );
  INV_X1 U579 ( .A(n927), .ZN(n643) );
  AOI22_X1 U580 ( .A1(data_in[5]), .A2(n826), .B1(n932), .B2(\mem[30][5] ), 
        .ZN(n927) );
  INV_X1 U581 ( .A(n926), .ZN(n642) );
  AOI22_X1 U582 ( .A1(data_in[6]), .A2(n826), .B1(n932), .B2(\mem[30][6] ), 
        .ZN(n926) );
  INV_X1 U583 ( .A(n925), .ZN(n641) );
  AOI22_X1 U584 ( .A1(data_in[7]), .A2(n826), .B1(n932), .B2(\mem[30][7] ), 
        .ZN(n925) );
  INV_X1 U585 ( .A(n924), .ZN(n640) );
  AOI22_X1 U586 ( .A1(data_in[0]), .A2(n825), .B1(n923), .B2(\mem[31][0] ), 
        .ZN(n924) );
  INV_X1 U587 ( .A(n922), .ZN(n639) );
  AOI22_X1 U588 ( .A1(data_in[1]), .A2(n825), .B1(n923), .B2(\mem[31][1] ), 
        .ZN(n922) );
  INV_X1 U589 ( .A(n921), .ZN(n638) );
  AOI22_X1 U590 ( .A1(data_in[2]), .A2(n825), .B1(n923), .B2(\mem[31][2] ), 
        .ZN(n921) );
  INV_X1 U591 ( .A(n920), .ZN(n637) );
  AOI22_X1 U592 ( .A1(data_in[3]), .A2(n825), .B1(n923), .B2(\mem[31][3] ), 
        .ZN(n920) );
  INV_X1 U593 ( .A(n919), .ZN(n636) );
  AOI22_X1 U594 ( .A1(data_in[4]), .A2(n825), .B1(n923), .B2(\mem[31][4] ), 
        .ZN(n919) );
  INV_X1 U595 ( .A(n918), .ZN(n635) );
  AOI22_X1 U596 ( .A1(data_in[5]), .A2(n825), .B1(n923), .B2(\mem[31][5] ), 
        .ZN(n918) );
  INV_X1 U597 ( .A(n917), .ZN(n634) );
  AOI22_X1 U598 ( .A1(data_in[6]), .A2(n825), .B1(n923), .B2(\mem[31][6] ), 
        .ZN(n917) );
  INV_X1 U599 ( .A(n916), .ZN(n633) );
  AOI22_X1 U600 ( .A1(data_in[7]), .A2(n825), .B1(n923), .B2(\mem[31][7] ), 
        .ZN(n916) );
  MUX2_X1 U601 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n614), .Z(n4) );
  MUX2_X1 U602 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n614), .Z(n5) );
  MUX2_X1 U603 ( .A(n5), .B(n4), .S(n611), .Z(n6) );
  MUX2_X1 U604 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n614), .Z(n7) );
  MUX2_X1 U605 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n614), .Z(n8) );
  MUX2_X1 U606 ( .A(n8), .B(n7), .S(n611), .Z(n9) );
  MUX2_X1 U607 ( .A(n9), .B(n6), .S(N12), .Z(n10) );
  MUX2_X1 U608 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n614), .Z(n11) );
  MUX2_X1 U609 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n614), .Z(n12) );
  MUX2_X1 U610 ( .A(n12), .B(n11), .S(n611), .Z(n13) );
  MUX2_X1 U611 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n614), .Z(n14) );
  MUX2_X1 U612 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n614), .Z(n15) );
  MUX2_X1 U613 ( .A(n15), .B(n14), .S(n611), .Z(n16) );
  MUX2_X1 U614 ( .A(n16), .B(n13), .S(n609), .Z(n17) );
  MUX2_X1 U615 ( .A(n17), .B(n10), .S(N13), .Z(n18) );
  MUX2_X1 U616 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n615), .Z(n19) );
  MUX2_X1 U617 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n615), .Z(n20) );
  MUX2_X1 U618 ( .A(n20), .B(n19), .S(n613), .Z(n21) );
  MUX2_X1 U619 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n615), .Z(n22) );
  MUX2_X1 U620 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n615), .Z(n23) );
  MUX2_X1 U621 ( .A(n23), .B(n22), .S(n611), .Z(n24) );
  MUX2_X1 U622 ( .A(n24), .B(n21), .S(n610), .Z(n25) );
  MUX2_X1 U623 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n615), .Z(n26) );
  MUX2_X1 U624 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n615), .Z(n27) );
  MUX2_X1 U625 ( .A(n27), .B(n26), .S(n611), .Z(n28) );
  MUX2_X1 U626 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n615), .Z(n29) );
  MUX2_X1 U627 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n615), .Z(n30) );
  MUX2_X1 U628 ( .A(n30), .B(n29), .S(n611), .Z(n31) );
  MUX2_X1 U629 ( .A(n31), .B(n28), .S(n610), .Z(n32) );
  MUX2_X1 U630 ( .A(n32), .B(n25), .S(N13), .Z(n33) );
  MUX2_X1 U631 ( .A(n33), .B(n18), .S(N14), .Z(N22) );
  MUX2_X1 U632 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n615), .Z(n34) );
  MUX2_X1 U633 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n615), .Z(n35) );
  MUX2_X1 U634 ( .A(n35), .B(n34), .S(n611), .Z(n36) );
  MUX2_X1 U635 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n615), .Z(n37) );
  MUX2_X1 U636 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n615), .Z(n38) );
  MUX2_X1 U637 ( .A(n38), .B(n37), .S(n611), .Z(n39) );
  MUX2_X1 U638 ( .A(n39), .B(n36), .S(N12), .Z(n40) );
  MUX2_X1 U639 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n616), .Z(n41) );
  MUX2_X1 U640 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n616), .Z(n42) );
  MUX2_X1 U641 ( .A(n42), .B(n41), .S(n611), .Z(n43) );
  MUX2_X1 U642 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n616), .Z(n44) );
  MUX2_X1 U643 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n616), .Z(n45) );
  MUX2_X1 U644 ( .A(n45), .B(n44), .S(n611), .Z(n46) );
  MUX2_X1 U645 ( .A(n46), .B(n43), .S(n610), .Z(n47) );
  MUX2_X1 U646 ( .A(n47), .B(n40), .S(N13), .Z(n48) );
  MUX2_X1 U647 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n616), .Z(n49) );
  MUX2_X1 U648 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n616), .Z(n50) );
  MUX2_X1 U649 ( .A(n50), .B(n49), .S(n611), .Z(n51) );
  MUX2_X1 U650 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n616), .Z(n52) );
  MUX2_X1 U651 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n616), .Z(n53) );
  MUX2_X1 U652 ( .A(n53), .B(n52), .S(n611), .Z(n54) );
  MUX2_X1 U653 ( .A(n54), .B(n51), .S(n609), .Z(n55) );
  MUX2_X1 U654 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n616), .Z(n56) );
  MUX2_X1 U655 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n616), .Z(n57) );
  MUX2_X1 U656 ( .A(n57), .B(n56), .S(n611), .Z(n58) );
  MUX2_X1 U657 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n616), .Z(n59) );
  MUX2_X1 U658 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n616), .Z(n60) );
  MUX2_X1 U659 ( .A(n60), .B(n59), .S(n612), .Z(n61) );
  MUX2_X1 U660 ( .A(n61), .B(n58), .S(N12), .Z(n62) );
  MUX2_X1 U661 ( .A(n62), .B(n55), .S(N13), .Z(n63) );
  MUX2_X1 U662 ( .A(n63), .B(n48), .S(N14), .Z(N21) );
  MUX2_X1 U663 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n617), .Z(n64) );
  MUX2_X1 U664 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n617), .Z(n65) );
  MUX2_X1 U665 ( .A(n65), .B(n64), .S(n612), .Z(n66) );
  MUX2_X1 U666 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n617), .Z(n67) );
  MUX2_X1 U667 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n617), .Z(n68) );
  MUX2_X1 U668 ( .A(n68), .B(n67), .S(n612), .Z(n69) );
  MUX2_X1 U669 ( .A(n69), .B(n66), .S(n609), .Z(n70) );
  MUX2_X1 U670 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n617), .Z(n71) );
  MUX2_X1 U671 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n617), .Z(n72) );
  MUX2_X1 U672 ( .A(n72), .B(n71), .S(n612), .Z(n73) );
  MUX2_X1 U673 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n617), .Z(n74) );
  MUX2_X1 U674 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n617), .Z(n75) );
  MUX2_X1 U675 ( .A(n75), .B(n74), .S(n612), .Z(n76) );
  MUX2_X1 U676 ( .A(n76), .B(n73), .S(n609), .Z(n77) );
  MUX2_X1 U677 ( .A(n77), .B(n70), .S(N13), .Z(n78) );
  MUX2_X1 U678 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n617), .Z(n79) );
  MUX2_X1 U679 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n617), .Z(n80) );
  MUX2_X1 U680 ( .A(n80), .B(n79), .S(n612), .Z(n81) );
  MUX2_X1 U681 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n617), .Z(n82) );
  MUX2_X1 U682 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n617), .Z(n83) );
  MUX2_X1 U683 ( .A(n83), .B(n82), .S(n612), .Z(n84) );
  MUX2_X1 U684 ( .A(n84), .B(n81), .S(n609), .Z(n85) );
  MUX2_X1 U685 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n618), .Z(n86) );
  MUX2_X1 U686 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n618), .Z(n87) );
  MUX2_X1 U687 ( .A(n87), .B(n86), .S(n612), .Z(n88) );
  MUX2_X1 U688 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n618), .Z(n89) );
  MUX2_X1 U689 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n618), .Z(n90) );
  MUX2_X1 U690 ( .A(n90), .B(n89), .S(n612), .Z(n91) );
  MUX2_X1 U691 ( .A(n91), .B(n88), .S(n609), .Z(n92) );
  MUX2_X1 U692 ( .A(n92), .B(n85), .S(N13), .Z(n93) );
  MUX2_X1 U693 ( .A(n93), .B(n78), .S(N14), .Z(N20) );
  MUX2_X1 U694 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n618), .Z(n94) );
  MUX2_X1 U695 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n618), .Z(n95) );
  MUX2_X1 U696 ( .A(n95), .B(n94), .S(n612), .Z(n96) );
  MUX2_X1 U697 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n618), .Z(n97) );
  MUX2_X1 U698 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n618), .Z(n98) );
  MUX2_X1 U699 ( .A(n98), .B(n97), .S(n612), .Z(n99) );
  MUX2_X1 U700 ( .A(n99), .B(n96), .S(n609), .Z(n100) );
  MUX2_X1 U701 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n618), .Z(n101) );
  MUX2_X1 U702 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n618), .Z(n102) );
  MUX2_X1 U703 ( .A(n102), .B(n101), .S(n612), .Z(n103) );
  MUX2_X1 U704 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n618), .Z(n104) );
  MUX2_X1 U705 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n618), .Z(n105) );
  MUX2_X1 U706 ( .A(n105), .B(n104), .S(n612), .Z(n106) );
  MUX2_X1 U707 ( .A(n106), .B(n103), .S(n609), .Z(n107) );
  MUX2_X1 U708 ( .A(n107), .B(n100), .S(N13), .Z(n108) );
  MUX2_X1 U709 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n619), .Z(n109) );
  MUX2_X1 U710 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n619), .Z(n110) );
  MUX2_X1 U711 ( .A(n110), .B(n109), .S(n613), .Z(n111) );
  MUX2_X1 U712 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n619), .Z(n112) );
  MUX2_X1 U713 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n619), .Z(n113) );
  MUX2_X1 U714 ( .A(n113), .B(n112), .S(n613), .Z(n114) );
  MUX2_X1 U715 ( .A(n114), .B(n111), .S(n609), .Z(n115) );
  MUX2_X1 U716 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n619), .Z(n116) );
  MUX2_X1 U717 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n619), .Z(n117) );
  MUX2_X1 U718 ( .A(n117), .B(n116), .S(n613), .Z(n118) );
  MUX2_X1 U719 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n619), .Z(n119) );
  MUX2_X1 U720 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n619), .Z(n120) );
  MUX2_X1 U721 ( .A(n120), .B(n119), .S(n613), .Z(n121) );
  MUX2_X1 U722 ( .A(n121), .B(n118), .S(n609), .Z(n122) );
  MUX2_X1 U723 ( .A(n122), .B(n115), .S(N13), .Z(n123) );
  MUX2_X1 U724 ( .A(n123), .B(n108), .S(N14), .Z(N19) );
  MUX2_X1 U725 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n619), .Z(n124) );
  MUX2_X1 U726 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n619), .Z(n125) );
  MUX2_X1 U727 ( .A(n125), .B(n124), .S(n613), .Z(n126) );
  MUX2_X1 U728 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n619), .Z(n127) );
  MUX2_X1 U729 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n619), .Z(n128) );
  MUX2_X1 U730 ( .A(n128), .B(n127), .S(n613), .Z(n129) );
  MUX2_X1 U731 ( .A(n129), .B(n126), .S(n609), .Z(n130) );
  MUX2_X1 U732 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n620), .Z(n131) );
  MUX2_X1 U733 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n620), .Z(n132) );
  MUX2_X1 U734 ( .A(n132), .B(n131), .S(n613), .Z(n133) );
  MUX2_X1 U735 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n620), .Z(n134) );
  MUX2_X1 U736 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n620), .Z(n135) );
  MUX2_X1 U737 ( .A(n135), .B(n134), .S(n613), .Z(n136) );
  MUX2_X1 U738 ( .A(n136), .B(n133), .S(n609), .Z(n137) );
  MUX2_X1 U739 ( .A(n137), .B(n130), .S(N13), .Z(n138) );
  MUX2_X1 U740 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n620), .Z(n139) );
  MUX2_X1 U741 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n620), .Z(n140) );
  MUX2_X1 U742 ( .A(n140), .B(n139), .S(n613), .Z(n141) );
  MUX2_X1 U743 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n620), .Z(n142) );
  MUX2_X1 U744 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n620), .Z(n143) );
  MUX2_X1 U745 ( .A(n143), .B(n142), .S(n613), .Z(n144) );
  MUX2_X1 U746 ( .A(n144), .B(n141), .S(n609), .Z(n145) );
  MUX2_X1 U747 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n620), .Z(n146) );
  MUX2_X1 U748 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n620), .Z(n147) );
  MUX2_X1 U749 ( .A(n147), .B(n146), .S(n613), .Z(n148) );
  MUX2_X1 U750 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n620), .Z(n149) );
  MUX2_X1 U751 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n620), .Z(n150) );
  MUX2_X1 U752 ( .A(n150), .B(n149), .S(n613), .Z(n151) );
  MUX2_X1 U753 ( .A(n151), .B(n148), .S(n609), .Z(n152) );
  MUX2_X1 U754 ( .A(n152), .B(n145), .S(N13), .Z(n153) );
  MUX2_X1 U755 ( .A(n153), .B(n138), .S(N14), .Z(N18) );
  MUX2_X1 U756 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n621), .Z(n154) );
  MUX2_X1 U757 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n621), .Z(n155) );
  MUX2_X1 U758 ( .A(n155), .B(n154), .S(n613), .Z(n156) );
  MUX2_X1 U759 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n616), .Z(n157) );
  MUX2_X1 U760 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n621), .Z(n158) );
  MUX2_X1 U761 ( .A(n158), .B(n157), .S(n611), .Z(n159) );
  MUX2_X1 U762 ( .A(n159), .B(n156), .S(n610), .Z(n160) );
  MUX2_X1 U763 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n622), .Z(n161) );
  MUX2_X1 U764 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n622), .Z(n162) );
  MUX2_X1 U765 ( .A(n162), .B(n161), .S(n613), .Z(n163) );
  MUX2_X1 U766 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n614), .Z(n164) );
  MUX2_X1 U767 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n622), .Z(n165) );
  MUX2_X1 U768 ( .A(n165), .B(n164), .S(n612), .Z(n166) );
  MUX2_X1 U769 ( .A(n166), .B(n163), .S(n610), .Z(n167) );
  MUX2_X1 U770 ( .A(n167), .B(n160), .S(N13), .Z(n168) );
  MUX2_X1 U771 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n615), .Z(n169) );
  MUX2_X1 U772 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n622), .Z(n170) );
  MUX2_X1 U773 ( .A(n170), .B(n169), .S(n612), .Z(n171) );
  MUX2_X1 U774 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n622), .Z(n172) );
  MUX2_X1 U775 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n621), .Z(n173) );
  MUX2_X1 U776 ( .A(n173), .B(n172), .S(n611), .Z(n174) );
  MUX2_X1 U777 ( .A(n174), .B(n171), .S(n610), .Z(n175) );
  MUX2_X1 U778 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n622), .Z(n176) );
  MUX2_X1 U779 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n622), .Z(n177) );
  MUX2_X1 U780 ( .A(n177), .B(n176), .S(n612), .Z(n178) );
  MUX2_X1 U781 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n622), .Z(n179) );
  MUX2_X1 U782 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n616), .Z(n180) );
  MUX2_X1 U783 ( .A(n180), .B(n179), .S(n612), .Z(n181) );
  MUX2_X1 U784 ( .A(n181), .B(n178), .S(n610), .Z(n182) );
  MUX2_X1 U785 ( .A(n182), .B(n175), .S(N13), .Z(n183) );
  MUX2_X1 U786 ( .A(n183), .B(n168), .S(N14), .Z(N17) );
  MUX2_X1 U787 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n614), .Z(n184) );
  MUX2_X1 U788 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n622), .Z(n185) );
  MUX2_X1 U789 ( .A(n185), .B(n184), .S(n611), .Z(n186) );
  MUX2_X1 U790 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n622), .Z(n187) );
  MUX2_X1 U791 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n622), .Z(n188) );
  MUX2_X1 U792 ( .A(n188), .B(n187), .S(n612), .Z(n189) );
  MUX2_X1 U793 ( .A(n189), .B(n186), .S(n610), .Z(n190) );
  MUX2_X1 U794 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n615), .Z(n191) );
  MUX2_X1 U795 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n618), .Z(n192) );
  MUX2_X1 U796 ( .A(n192), .B(n191), .S(N11), .Z(n193) );
  MUX2_X1 U797 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n622), .Z(n194) );
  MUX2_X1 U798 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n617), .Z(n195) );
  MUX2_X1 U799 ( .A(n195), .B(n194), .S(n613), .Z(n196) );
  MUX2_X1 U800 ( .A(n196), .B(n193), .S(n610), .Z(n197) );
  MUX2_X1 U801 ( .A(n197), .B(n190), .S(N13), .Z(n198) );
  MUX2_X1 U802 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n621), .Z(n199) );
  MUX2_X1 U803 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n619), .Z(n200) );
  MUX2_X1 U804 ( .A(n200), .B(n199), .S(n613), .Z(n201) );
  MUX2_X1 U805 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n618), .Z(n202) );
  MUX2_X1 U806 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n621), .Z(n203) );
  MUX2_X1 U807 ( .A(n203), .B(n202), .S(n612), .Z(n204) );
  MUX2_X1 U808 ( .A(n204), .B(n201), .S(n610), .Z(n205) );
  MUX2_X1 U809 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n620), .Z(n206) );
  MUX2_X1 U810 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n621), .Z(n207) );
  MUX2_X1 U811 ( .A(n207), .B(n206), .S(n613), .Z(n208) );
  MUX2_X1 U812 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n622), .Z(n209) );
  MUX2_X1 U813 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n210) );
  MUX2_X1 U814 ( .A(n210), .B(n209), .S(N11), .Z(n211) );
  MUX2_X1 U815 ( .A(n211), .B(n208), .S(n610), .Z(n212) );
  MUX2_X1 U816 ( .A(n212), .B(n205), .S(N13), .Z(n213) );
  MUX2_X1 U817 ( .A(n213), .B(n198), .S(N14), .Z(N16) );
  MUX2_X1 U818 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n614), .Z(n214) );
  MUX2_X1 U819 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n617), .Z(n215) );
  MUX2_X1 U820 ( .A(n215), .B(n214), .S(n611), .Z(n216) );
  MUX2_X1 U821 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n621), .Z(n217) );
  MUX2_X1 U822 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n622), .Z(n218) );
  MUX2_X1 U823 ( .A(n218), .B(n217), .S(n613), .Z(n219) );
  MUX2_X1 U824 ( .A(n219), .B(n216), .S(n610), .Z(n220) );
  MUX2_X1 U825 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n614), .Z(n221) );
  MUX2_X1 U826 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n622), .Z(n222) );
  MUX2_X1 U827 ( .A(n222), .B(n221), .S(n613), .Z(n223) );
  MUX2_X1 U828 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n622), .Z(n224) );
  MUX2_X1 U829 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n225) );
  MUX2_X1 U830 ( .A(n225), .B(n224), .S(N11), .Z(n226) );
  MUX2_X1 U831 ( .A(n226), .B(n223), .S(n610), .Z(n227) );
  MUX2_X1 U832 ( .A(n227), .B(n220), .S(N13), .Z(n228) );
  MUX2_X1 U833 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n614), .Z(n229) );
  MUX2_X1 U834 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n614), .Z(n595) );
  MUX2_X1 U835 ( .A(n595), .B(n229), .S(n611), .Z(n596) );
  MUX2_X1 U836 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n621), .Z(n597) );
  MUX2_X1 U837 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n598) );
  MUX2_X1 U838 ( .A(n598), .B(n597), .S(N11), .Z(n599) );
  MUX2_X1 U839 ( .A(n599), .B(n596), .S(n610), .Z(n600) );
  MUX2_X1 U840 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n614), .Z(n601) );
  MUX2_X1 U841 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n621), .Z(n602) );
  MUX2_X1 U842 ( .A(n602), .B(n601), .S(n613), .Z(n603) );
  MUX2_X1 U843 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n604) );
  MUX2_X1 U844 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n605) );
  MUX2_X1 U845 ( .A(n605), .B(n604), .S(N11), .Z(n606) );
  MUX2_X1 U846 ( .A(n606), .B(n603), .S(n610), .Z(n607) );
  MUX2_X1 U847 ( .A(n607), .B(n600), .S(N13), .Z(n608) );
  MUX2_X1 U848 ( .A(n608), .B(n228), .S(N14), .Z(N15) );
  CLKBUF_X1 U849 ( .A(N11), .Z(n611) );
  INV_X1 U850 ( .A(N10), .ZN(n623) );
  INV_X1 U851 ( .A(N11), .ZN(n624) );
  INV_X1 U852 ( .A(data_in[0]), .ZN(n625) );
  INV_X1 U853 ( .A(data_in[1]), .ZN(n626) );
  INV_X1 U854 ( .A(data_in[2]), .ZN(n627) );
  INV_X1 U855 ( .A(data_in[3]), .ZN(n628) );
  INV_X1 U856 ( .A(data_in[4]), .ZN(n629) );
  INV_X1 U857 ( .A(data_in[5]), .ZN(n630) );
  INV_X1 U858 ( .A(data_in[6]), .ZN(n631) );
  INV_X1 U859 ( .A(data_in[7]), .ZN(n632) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_9 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n634), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n635), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n636), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n637), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n638), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n639), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n640), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n641), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n642), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n643), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n644), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n645), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n646), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n647), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n648), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n649), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n650), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n651), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n652), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n653), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n654), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n655), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n656), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n657), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n658), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n659), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n660), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n661), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n662), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n663), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n664), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n665), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n666), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n667), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n668), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n669), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n670), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n671), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n672), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n673), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n674), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n675), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n676), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n677), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n678), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n679), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n680), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n681), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n682), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n683), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n684), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n685), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n686), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n687), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n688), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n689), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n690), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n691), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n692), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n693), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n694), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n695), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n696), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n697), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n698), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n699), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n700), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n701), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n702), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n703), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n704), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n705), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n706), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n707), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n708), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n709), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n710), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n711), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n712), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n713), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n714), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n715), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n716), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n717), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n718), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n719), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n720), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n721), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n722), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n723), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n724), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n725), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n726), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n727), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n728), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n729), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n730), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n731), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n732), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n733), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n734), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n735), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n736), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n737), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n738), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n739), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n740), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n741), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n742), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n743), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n744), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n745), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n746), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n747), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n748), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n749), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n750), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n751), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n752), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n753), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n754), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n755), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n756), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n757), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n758), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n759), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n760), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n761), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n762), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n763), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n764), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n765), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n766), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n767), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n768), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n769), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n770), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n771), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n772), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n773), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n774), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n775), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n776), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n777), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n778), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n779), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n780), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n781), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n782), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n783), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n784), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n785), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n786), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n787), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n788), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n789), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n790), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n791), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n792), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n793), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n794), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n795), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n796), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n797), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n798), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n799), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n800), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n801), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n802), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n803), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n804), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n805), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n806), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n807), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n808), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n809), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n810), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n811), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n812), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n813), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n814), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n815), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n816), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n817), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n818), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n819), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n820), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n821), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n822), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n823), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n824), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n825), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n853), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n854), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n855), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n856), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n857), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n858), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n859), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n860), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n861), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n862), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n863), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n864), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n865), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n866), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n867), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n868), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n869), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n870), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n871), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n872), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n873), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n874), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n875), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n876), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n877), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n878), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n879), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n880), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n881), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n882), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n883), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n884), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n885), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n886), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n887), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n888), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n889), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n890), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n891), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n892), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n893), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n894), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n895), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n896), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n897), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n898), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n899), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n900), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n901), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n902), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n903), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n904), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n905), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n906), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n907), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n908), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n909), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n910), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n911), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n912), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n913), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n914), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n915), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n916), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .QN(n2) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  CLKBUF_X1 U3 ( .A(N10), .Z(n623) );
  BUF_X1 U4 ( .A(n622), .Z(n614) );
  NOR2_X1 U5 ( .A1(n850), .A2(addr[5]), .ZN(n1136) );
  AND3_X1 U6 ( .A1(n851), .A2(n852), .A3(n1136), .ZN(n1207) );
  AND3_X1 U7 ( .A1(n1136), .A2(n852), .A3(N13), .ZN(n1126) );
  AND3_X1 U8 ( .A1(n1136), .A2(n851), .A3(N14), .ZN(n1053) );
  AND3_X1 U9 ( .A1(N13), .A2(n1136), .A3(N14), .ZN(n980) );
  INV_X2 U10 ( .A(n2), .ZN(data_out[1]) );
  BUF_X1 U11 ( .A(n623), .Z(n620) );
  BUF_X1 U12 ( .A(n623), .Z(n621) );
  BUF_X1 U13 ( .A(n623), .Z(n619) );
  BUF_X1 U14 ( .A(n622), .Z(n616) );
  BUF_X1 U15 ( .A(n622), .Z(n615) );
  BUF_X1 U16 ( .A(n622), .Z(n617) );
  BUF_X1 U17 ( .A(n622), .Z(n618) );
  BUF_X1 U18 ( .A(N11), .Z(n612) );
  BUF_X1 U19 ( .A(N11), .Z(n613) );
  BUF_X1 U20 ( .A(N10), .Z(n622) );
  NOR3_X1 U21 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1208) );
  NOR3_X1 U22 ( .A1(N11), .A2(N12), .A3(n624), .ZN(n1197) );
  NOR3_X1 U23 ( .A1(N10), .A2(N12), .A3(n625), .ZN(n1187) );
  NOR3_X1 U24 ( .A1(n624), .A2(N12), .A3(n625), .ZN(n1177) );
  INV_X1 U25 ( .A(n1134), .ZN(n849) );
  INV_X1 U26 ( .A(n1124), .ZN(n848) );
  INV_X1 U27 ( .A(n1115), .ZN(n847) );
  INV_X1 U28 ( .A(n1106), .ZN(n846) );
  INV_X1 U29 ( .A(n1061), .ZN(n841) );
  INV_X1 U30 ( .A(n1051), .ZN(n840) );
  INV_X1 U31 ( .A(n1042), .ZN(n839) );
  INV_X1 U32 ( .A(n1033), .ZN(n838) );
  INV_X1 U33 ( .A(n988), .ZN(n833) );
  INV_X1 U34 ( .A(n978), .ZN(n832) );
  INV_X1 U35 ( .A(n969), .ZN(n831) );
  INV_X1 U36 ( .A(n960), .ZN(n830) );
  INV_X1 U37 ( .A(n1097), .ZN(n845) );
  INV_X1 U38 ( .A(n1088), .ZN(n844) );
  INV_X1 U39 ( .A(n1079), .ZN(n843) );
  INV_X1 U40 ( .A(n1070), .ZN(n842) );
  INV_X1 U41 ( .A(n951), .ZN(n829) );
  INV_X1 U42 ( .A(n942), .ZN(n828) );
  INV_X1 U43 ( .A(n933), .ZN(n827) );
  INV_X1 U44 ( .A(n924), .ZN(n826) );
  INV_X1 U45 ( .A(n1024), .ZN(n837) );
  INV_X1 U46 ( .A(n1015), .ZN(n836) );
  INV_X1 U47 ( .A(n1006), .ZN(n835) );
  INV_X1 U48 ( .A(n997), .ZN(n834) );
  BUF_X1 U49 ( .A(N12), .Z(n609) );
  BUF_X1 U50 ( .A(N12), .Z(n610) );
  INV_X1 U51 ( .A(N13), .ZN(n851) );
  AND3_X1 U52 ( .A1(n624), .A2(n625), .A3(N12), .ZN(n1167) );
  AND3_X1 U53 ( .A1(N10), .A2(n625), .A3(N12), .ZN(n1157) );
  AND3_X1 U54 ( .A1(N11), .A2(n624), .A3(N12), .ZN(n1147) );
  AND3_X1 U55 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1137) );
  INV_X1 U56 ( .A(N14), .ZN(n852) );
  NAND2_X1 U57 ( .A1(n1197), .A2(n1207), .ZN(n1206) );
  NAND2_X1 U58 ( .A1(n1187), .A2(n1207), .ZN(n1196) );
  NAND2_X1 U59 ( .A1(n1177), .A2(n1207), .ZN(n1186) );
  NAND2_X1 U60 ( .A1(n1167), .A2(n1207), .ZN(n1176) );
  NAND2_X1 U61 ( .A1(n1157), .A2(n1207), .ZN(n1166) );
  NAND2_X1 U62 ( .A1(n1147), .A2(n1207), .ZN(n1156) );
  NAND2_X1 U63 ( .A1(n1137), .A2(n1207), .ZN(n1146) );
  NAND2_X1 U64 ( .A1(n1208), .A2(n1207), .ZN(n1217) );
  NAND2_X1 U65 ( .A1(n1126), .A2(n1208), .ZN(n1134) );
  NAND2_X1 U66 ( .A1(n1126), .A2(n1197), .ZN(n1124) );
  NAND2_X1 U67 ( .A1(n1126), .A2(n1187), .ZN(n1115) );
  NAND2_X1 U68 ( .A1(n1126), .A2(n1177), .ZN(n1106) );
  NAND2_X1 U69 ( .A1(n1053), .A2(n1208), .ZN(n1061) );
  NAND2_X1 U70 ( .A1(n1053), .A2(n1197), .ZN(n1051) );
  NAND2_X1 U71 ( .A1(n1053), .A2(n1187), .ZN(n1042) );
  NAND2_X1 U72 ( .A1(n1053), .A2(n1177), .ZN(n1033) );
  NAND2_X1 U73 ( .A1(n980), .A2(n1208), .ZN(n988) );
  NAND2_X1 U74 ( .A1(n980), .A2(n1197), .ZN(n978) );
  NAND2_X1 U75 ( .A1(n980), .A2(n1187), .ZN(n969) );
  NAND2_X1 U76 ( .A1(n980), .A2(n1177), .ZN(n960) );
  NAND2_X1 U77 ( .A1(n1126), .A2(n1167), .ZN(n1097) );
  NAND2_X1 U78 ( .A1(n1126), .A2(n1157), .ZN(n1088) );
  NAND2_X1 U79 ( .A1(n1126), .A2(n1147), .ZN(n1079) );
  NAND2_X1 U80 ( .A1(n1126), .A2(n1137), .ZN(n1070) );
  NAND2_X1 U81 ( .A1(n1053), .A2(n1167), .ZN(n1024) );
  NAND2_X1 U82 ( .A1(n1053), .A2(n1157), .ZN(n1015) );
  NAND2_X1 U83 ( .A1(n1053), .A2(n1147), .ZN(n1006) );
  NAND2_X1 U84 ( .A1(n1053), .A2(n1137), .ZN(n997) );
  NAND2_X1 U85 ( .A1(n980), .A2(n1167), .ZN(n951) );
  NAND2_X1 U86 ( .A1(n980), .A2(n1157), .ZN(n942) );
  NAND2_X1 U87 ( .A1(n980), .A2(n1147), .ZN(n933) );
  NAND2_X1 U88 ( .A1(n980), .A2(n1137), .ZN(n924) );
  INV_X1 U89 ( .A(wr_en), .ZN(n850) );
  OAI21_X1 U90 ( .B1(n626), .B2(n1176), .A(n1175), .ZN(n884) );
  NAND2_X1 U91 ( .A1(\mem[4][0] ), .A2(n1176), .ZN(n1175) );
  OAI21_X1 U92 ( .B1(n627), .B2(n1176), .A(n1174), .ZN(n883) );
  NAND2_X1 U93 ( .A1(\mem[4][1] ), .A2(n1176), .ZN(n1174) );
  OAI21_X1 U94 ( .B1(n628), .B2(n1176), .A(n1173), .ZN(n882) );
  NAND2_X1 U95 ( .A1(\mem[4][2] ), .A2(n1176), .ZN(n1173) );
  OAI21_X1 U96 ( .B1(n629), .B2(n1176), .A(n1172), .ZN(n881) );
  NAND2_X1 U97 ( .A1(\mem[4][3] ), .A2(n1176), .ZN(n1172) );
  OAI21_X1 U98 ( .B1(n630), .B2(n1176), .A(n1171), .ZN(n880) );
  NAND2_X1 U99 ( .A1(\mem[4][4] ), .A2(n1176), .ZN(n1171) );
  OAI21_X1 U100 ( .B1(n631), .B2(n1176), .A(n1170), .ZN(n879) );
  NAND2_X1 U101 ( .A1(\mem[4][5] ), .A2(n1176), .ZN(n1170) );
  OAI21_X1 U102 ( .B1(n632), .B2(n1176), .A(n1169), .ZN(n878) );
  NAND2_X1 U103 ( .A1(\mem[4][6] ), .A2(n1176), .ZN(n1169) );
  OAI21_X1 U104 ( .B1(n633), .B2(n1176), .A(n1168), .ZN(n877) );
  NAND2_X1 U105 ( .A1(\mem[4][7] ), .A2(n1176), .ZN(n1168) );
  OAI21_X1 U106 ( .B1(n626), .B2(n1156), .A(n1155), .ZN(n868) );
  NAND2_X1 U107 ( .A1(\mem[6][0] ), .A2(n1156), .ZN(n1155) );
  OAI21_X1 U108 ( .B1(n627), .B2(n1156), .A(n1154), .ZN(n867) );
  NAND2_X1 U109 ( .A1(\mem[6][1] ), .A2(n1156), .ZN(n1154) );
  OAI21_X1 U110 ( .B1(n628), .B2(n1156), .A(n1153), .ZN(n866) );
  NAND2_X1 U111 ( .A1(\mem[6][2] ), .A2(n1156), .ZN(n1153) );
  OAI21_X1 U112 ( .B1(n629), .B2(n1156), .A(n1152), .ZN(n865) );
  NAND2_X1 U113 ( .A1(\mem[6][3] ), .A2(n1156), .ZN(n1152) );
  OAI21_X1 U114 ( .B1(n630), .B2(n1156), .A(n1151), .ZN(n864) );
  NAND2_X1 U115 ( .A1(\mem[6][4] ), .A2(n1156), .ZN(n1151) );
  OAI21_X1 U116 ( .B1(n631), .B2(n1156), .A(n1150), .ZN(n863) );
  NAND2_X1 U117 ( .A1(\mem[6][5] ), .A2(n1156), .ZN(n1150) );
  OAI21_X1 U118 ( .B1(n632), .B2(n1156), .A(n1149), .ZN(n862) );
  NAND2_X1 U119 ( .A1(\mem[6][6] ), .A2(n1156), .ZN(n1149) );
  OAI21_X1 U120 ( .B1(n633), .B2(n1156), .A(n1148), .ZN(n861) );
  NAND2_X1 U121 ( .A1(\mem[6][7] ), .A2(n1156), .ZN(n1148) );
  OAI21_X1 U122 ( .B1(n626), .B2(n1146), .A(n1145), .ZN(n860) );
  NAND2_X1 U123 ( .A1(\mem[7][0] ), .A2(n1146), .ZN(n1145) );
  OAI21_X1 U124 ( .B1(n627), .B2(n1146), .A(n1144), .ZN(n859) );
  NAND2_X1 U125 ( .A1(\mem[7][1] ), .A2(n1146), .ZN(n1144) );
  OAI21_X1 U126 ( .B1(n628), .B2(n1146), .A(n1143), .ZN(n858) );
  NAND2_X1 U127 ( .A1(\mem[7][2] ), .A2(n1146), .ZN(n1143) );
  OAI21_X1 U128 ( .B1(n629), .B2(n1146), .A(n1142), .ZN(n857) );
  NAND2_X1 U129 ( .A1(\mem[7][3] ), .A2(n1146), .ZN(n1142) );
  OAI21_X1 U130 ( .B1(n630), .B2(n1146), .A(n1141), .ZN(n856) );
  NAND2_X1 U131 ( .A1(\mem[7][4] ), .A2(n1146), .ZN(n1141) );
  OAI21_X1 U132 ( .B1(n631), .B2(n1146), .A(n1140), .ZN(n855) );
  NAND2_X1 U133 ( .A1(\mem[7][5] ), .A2(n1146), .ZN(n1140) );
  OAI21_X1 U134 ( .B1(n632), .B2(n1146), .A(n1139), .ZN(n854) );
  NAND2_X1 U135 ( .A1(\mem[7][6] ), .A2(n1146), .ZN(n1139) );
  OAI21_X1 U136 ( .B1(n633), .B2(n1146), .A(n1138), .ZN(n853) );
  NAND2_X1 U137 ( .A1(\mem[7][7] ), .A2(n1146), .ZN(n1138) );
  OAI21_X1 U138 ( .B1(n626), .B2(n1206), .A(n1205), .ZN(n908) );
  NAND2_X1 U139 ( .A1(\mem[1][0] ), .A2(n1206), .ZN(n1205) );
  OAI21_X1 U140 ( .B1(n627), .B2(n1206), .A(n1204), .ZN(n907) );
  NAND2_X1 U141 ( .A1(\mem[1][1] ), .A2(n1206), .ZN(n1204) );
  OAI21_X1 U142 ( .B1(n628), .B2(n1206), .A(n1203), .ZN(n906) );
  NAND2_X1 U143 ( .A1(\mem[1][2] ), .A2(n1206), .ZN(n1203) );
  OAI21_X1 U144 ( .B1(n629), .B2(n1206), .A(n1202), .ZN(n905) );
  NAND2_X1 U145 ( .A1(\mem[1][3] ), .A2(n1206), .ZN(n1202) );
  OAI21_X1 U146 ( .B1(n630), .B2(n1206), .A(n1201), .ZN(n904) );
  NAND2_X1 U147 ( .A1(\mem[1][4] ), .A2(n1206), .ZN(n1201) );
  OAI21_X1 U148 ( .B1(n631), .B2(n1206), .A(n1200), .ZN(n903) );
  NAND2_X1 U149 ( .A1(\mem[1][5] ), .A2(n1206), .ZN(n1200) );
  OAI21_X1 U150 ( .B1(n632), .B2(n1206), .A(n1199), .ZN(n902) );
  NAND2_X1 U151 ( .A1(\mem[1][6] ), .A2(n1206), .ZN(n1199) );
  OAI21_X1 U152 ( .B1(n633), .B2(n1206), .A(n1198), .ZN(n901) );
  NAND2_X1 U153 ( .A1(\mem[1][7] ), .A2(n1206), .ZN(n1198) );
  OAI21_X1 U154 ( .B1(n626), .B2(n1196), .A(n1195), .ZN(n900) );
  NAND2_X1 U155 ( .A1(\mem[2][0] ), .A2(n1196), .ZN(n1195) );
  OAI21_X1 U156 ( .B1(n627), .B2(n1196), .A(n1194), .ZN(n899) );
  NAND2_X1 U157 ( .A1(\mem[2][1] ), .A2(n1196), .ZN(n1194) );
  OAI21_X1 U158 ( .B1(n628), .B2(n1196), .A(n1193), .ZN(n898) );
  NAND2_X1 U159 ( .A1(\mem[2][2] ), .A2(n1196), .ZN(n1193) );
  OAI21_X1 U160 ( .B1(n629), .B2(n1196), .A(n1192), .ZN(n897) );
  NAND2_X1 U161 ( .A1(\mem[2][3] ), .A2(n1196), .ZN(n1192) );
  OAI21_X1 U162 ( .B1(n630), .B2(n1196), .A(n1191), .ZN(n896) );
  NAND2_X1 U163 ( .A1(\mem[2][4] ), .A2(n1196), .ZN(n1191) );
  OAI21_X1 U164 ( .B1(n631), .B2(n1196), .A(n1190), .ZN(n895) );
  NAND2_X1 U165 ( .A1(\mem[2][5] ), .A2(n1196), .ZN(n1190) );
  OAI21_X1 U166 ( .B1(n632), .B2(n1196), .A(n1189), .ZN(n894) );
  NAND2_X1 U167 ( .A1(\mem[2][6] ), .A2(n1196), .ZN(n1189) );
  OAI21_X1 U168 ( .B1(n633), .B2(n1196), .A(n1188), .ZN(n893) );
  NAND2_X1 U169 ( .A1(\mem[2][7] ), .A2(n1196), .ZN(n1188) );
  OAI21_X1 U170 ( .B1(n626), .B2(n1186), .A(n1185), .ZN(n892) );
  NAND2_X1 U171 ( .A1(\mem[3][0] ), .A2(n1186), .ZN(n1185) );
  OAI21_X1 U172 ( .B1(n627), .B2(n1186), .A(n1184), .ZN(n891) );
  NAND2_X1 U173 ( .A1(\mem[3][1] ), .A2(n1186), .ZN(n1184) );
  OAI21_X1 U174 ( .B1(n628), .B2(n1186), .A(n1183), .ZN(n890) );
  NAND2_X1 U175 ( .A1(\mem[3][2] ), .A2(n1186), .ZN(n1183) );
  OAI21_X1 U176 ( .B1(n629), .B2(n1186), .A(n1182), .ZN(n889) );
  NAND2_X1 U177 ( .A1(\mem[3][3] ), .A2(n1186), .ZN(n1182) );
  OAI21_X1 U178 ( .B1(n630), .B2(n1186), .A(n1181), .ZN(n888) );
  NAND2_X1 U179 ( .A1(\mem[3][4] ), .A2(n1186), .ZN(n1181) );
  OAI21_X1 U180 ( .B1(n631), .B2(n1186), .A(n1180), .ZN(n887) );
  NAND2_X1 U181 ( .A1(\mem[3][5] ), .A2(n1186), .ZN(n1180) );
  OAI21_X1 U182 ( .B1(n632), .B2(n1186), .A(n1179), .ZN(n886) );
  NAND2_X1 U183 ( .A1(\mem[3][6] ), .A2(n1186), .ZN(n1179) );
  OAI21_X1 U184 ( .B1(n633), .B2(n1186), .A(n1178), .ZN(n885) );
  NAND2_X1 U185 ( .A1(\mem[3][7] ), .A2(n1186), .ZN(n1178) );
  OAI21_X1 U186 ( .B1(n626), .B2(n1166), .A(n1165), .ZN(n876) );
  NAND2_X1 U187 ( .A1(\mem[5][0] ), .A2(n1166), .ZN(n1165) );
  OAI21_X1 U188 ( .B1(n627), .B2(n1166), .A(n1164), .ZN(n875) );
  NAND2_X1 U189 ( .A1(\mem[5][1] ), .A2(n1166), .ZN(n1164) );
  OAI21_X1 U190 ( .B1(n628), .B2(n1166), .A(n1163), .ZN(n874) );
  NAND2_X1 U191 ( .A1(\mem[5][2] ), .A2(n1166), .ZN(n1163) );
  OAI21_X1 U192 ( .B1(n629), .B2(n1166), .A(n1162), .ZN(n873) );
  NAND2_X1 U193 ( .A1(\mem[5][3] ), .A2(n1166), .ZN(n1162) );
  OAI21_X1 U194 ( .B1(n630), .B2(n1166), .A(n1161), .ZN(n872) );
  NAND2_X1 U195 ( .A1(\mem[5][4] ), .A2(n1166), .ZN(n1161) );
  OAI21_X1 U196 ( .B1(n631), .B2(n1166), .A(n1160), .ZN(n871) );
  NAND2_X1 U197 ( .A1(\mem[5][5] ), .A2(n1166), .ZN(n1160) );
  OAI21_X1 U198 ( .B1(n632), .B2(n1166), .A(n1159), .ZN(n870) );
  NAND2_X1 U199 ( .A1(\mem[5][6] ), .A2(n1166), .ZN(n1159) );
  OAI21_X1 U200 ( .B1(n633), .B2(n1166), .A(n1158), .ZN(n869) );
  NAND2_X1 U201 ( .A1(\mem[5][7] ), .A2(n1166), .ZN(n1158) );
  OAI21_X1 U202 ( .B1(n1217), .B2(n626), .A(n1216), .ZN(n916) );
  NAND2_X1 U203 ( .A1(\mem[0][0] ), .A2(n1217), .ZN(n1216) );
  OAI21_X1 U204 ( .B1(n1217), .B2(n627), .A(n1215), .ZN(n915) );
  NAND2_X1 U205 ( .A1(\mem[0][1] ), .A2(n1217), .ZN(n1215) );
  OAI21_X1 U206 ( .B1(n1217), .B2(n628), .A(n1214), .ZN(n914) );
  NAND2_X1 U207 ( .A1(\mem[0][2] ), .A2(n1217), .ZN(n1214) );
  OAI21_X1 U208 ( .B1(n1217), .B2(n629), .A(n1213), .ZN(n913) );
  NAND2_X1 U209 ( .A1(\mem[0][3] ), .A2(n1217), .ZN(n1213) );
  OAI21_X1 U210 ( .B1(n1217), .B2(n630), .A(n1212), .ZN(n912) );
  NAND2_X1 U211 ( .A1(\mem[0][4] ), .A2(n1217), .ZN(n1212) );
  OAI21_X1 U212 ( .B1(n1217), .B2(n631), .A(n1211), .ZN(n911) );
  NAND2_X1 U213 ( .A1(\mem[0][5] ), .A2(n1217), .ZN(n1211) );
  OAI21_X1 U214 ( .B1(n1217), .B2(n632), .A(n1210), .ZN(n910) );
  NAND2_X1 U215 ( .A1(\mem[0][6] ), .A2(n1217), .ZN(n1210) );
  OAI21_X1 U216 ( .B1(n1217), .B2(n633), .A(n1209), .ZN(n909) );
  NAND2_X1 U217 ( .A1(\mem[0][7] ), .A2(n1217), .ZN(n1209) );
  INV_X1 U218 ( .A(n1135), .ZN(n825) );
  AOI22_X1 U219 ( .A1(data_in[0]), .A2(n849), .B1(n1134), .B2(\mem[8][0] ), 
        .ZN(n1135) );
  INV_X1 U220 ( .A(n1133), .ZN(n824) );
  AOI22_X1 U221 ( .A1(data_in[1]), .A2(n849), .B1(n1134), .B2(\mem[8][1] ), 
        .ZN(n1133) );
  INV_X1 U222 ( .A(n1132), .ZN(n823) );
  AOI22_X1 U223 ( .A1(data_in[2]), .A2(n849), .B1(n1134), .B2(\mem[8][2] ), 
        .ZN(n1132) );
  INV_X1 U224 ( .A(n1131), .ZN(n822) );
  AOI22_X1 U225 ( .A1(data_in[3]), .A2(n849), .B1(n1134), .B2(\mem[8][3] ), 
        .ZN(n1131) );
  INV_X1 U226 ( .A(n1130), .ZN(n821) );
  AOI22_X1 U227 ( .A1(data_in[4]), .A2(n849), .B1(n1134), .B2(\mem[8][4] ), 
        .ZN(n1130) );
  INV_X1 U228 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U229 ( .A1(data_in[5]), .A2(n849), .B1(n1134), .B2(\mem[8][5] ), 
        .ZN(n1129) );
  INV_X1 U230 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U231 ( .A1(data_in[6]), .A2(n849), .B1(n1134), .B2(\mem[8][6] ), 
        .ZN(n1128) );
  INV_X1 U232 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n849), .B1(n1134), .B2(\mem[8][7] ), 
        .ZN(n1127) );
  INV_X1 U234 ( .A(n1125), .ZN(n817) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n848), .B1(n1124), .B2(\mem[9][0] ), 
        .ZN(n1125) );
  INV_X1 U236 ( .A(n1123), .ZN(n816) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n848), .B1(n1124), .B2(\mem[9][1] ), 
        .ZN(n1123) );
  INV_X1 U238 ( .A(n1122), .ZN(n815) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n848), .B1(n1124), .B2(\mem[9][2] ), 
        .ZN(n1122) );
  INV_X1 U240 ( .A(n1121), .ZN(n814) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n848), .B1(n1124), .B2(\mem[9][3] ), 
        .ZN(n1121) );
  INV_X1 U242 ( .A(n1120), .ZN(n813) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n848), .B1(n1124), .B2(\mem[9][4] ), 
        .ZN(n1120) );
  INV_X1 U244 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n848), .B1(n1124), .B2(\mem[9][5] ), 
        .ZN(n1119) );
  INV_X1 U246 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n848), .B1(n1124), .B2(\mem[9][6] ), 
        .ZN(n1118) );
  INV_X1 U248 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n848), .B1(n1124), .B2(\mem[9][7] ), 
        .ZN(n1117) );
  INV_X1 U250 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n847), .B1(n1115), .B2(\mem[10][0] ), 
        .ZN(n1116) );
  INV_X1 U252 ( .A(n1114), .ZN(n808) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n847), .B1(n1115), .B2(\mem[10][1] ), 
        .ZN(n1114) );
  INV_X1 U254 ( .A(n1113), .ZN(n807) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n847), .B1(n1115), .B2(\mem[10][2] ), 
        .ZN(n1113) );
  INV_X1 U256 ( .A(n1112), .ZN(n806) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n847), .B1(n1115), .B2(\mem[10][3] ), 
        .ZN(n1112) );
  INV_X1 U258 ( .A(n1111), .ZN(n805) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n847), .B1(n1115), .B2(\mem[10][4] ), 
        .ZN(n1111) );
  INV_X1 U260 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n847), .B1(n1115), .B2(\mem[10][5] ), 
        .ZN(n1110) );
  INV_X1 U262 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n847), .B1(n1115), .B2(\mem[10][6] ), 
        .ZN(n1109) );
  INV_X1 U264 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n847), .B1(n1115), .B2(\mem[10][7] ), 
        .ZN(n1108) );
  INV_X1 U266 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n846), .B1(n1106), .B2(\mem[11][0] ), 
        .ZN(n1107) );
  INV_X1 U268 ( .A(n1105), .ZN(n800) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n846), .B1(n1106), .B2(\mem[11][1] ), 
        .ZN(n1105) );
  INV_X1 U270 ( .A(n1104), .ZN(n799) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n846), .B1(n1106), .B2(\mem[11][2] ), 
        .ZN(n1104) );
  INV_X1 U272 ( .A(n1103), .ZN(n798) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n846), .B1(n1106), .B2(\mem[11][3] ), 
        .ZN(n1103) );
  INV_X1 U274 ( .A(n1102), .ZN(n797) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n846), .B1(n1106), .B2(\mem[11][4] ), 
        .ZN(n1102) );
  INV_X1 U276 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n846), .B1(n1106), .B2(\mem[11][5] ), 
        .ZN(n1101) );
  INV_X1 U278 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n846), .B1(n1106), .B2(\mem[11][6] ), 
        .ZN(n1100) );
  INV_X1 U280 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n846), .B1(n1106), .B2(\mem[11][7] ), 
        .ZN(n1099) );
  INV_X1 U282 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n845), .B1(n1097), .B2(\mem[12][0] ), 
        .ZN(n1098) );
  INV_X1 U284 ( .A(n1096), .ZN(n792) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n845), .B1(n1097), .B2(\mem[12][1] ), 
        .ZN(n1096) );
  INV_X1 U286 ( .A(n1095), .ZN(n791) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n845), .B1(n1097), .B2(\mem[12][2] ), 
        .ZN(n1095) );
  INV_X1 U288 ( .A(n1094), .ZN(n790) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n845), .B1(n1097), .B2(\mem[12][3] ), 
        .ZN(n1094) );
  INV_X1 U290 ( .A(n1093), .ZN(n789) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n845), .B1(n1097), .B2(\mem[12][4] ), 
        .ZN(n1093) );
  INV_X1 U292 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n845), .B1(n1097), .B2(\mem[12][5] ), 
        .ZN(n1092) );
  INV_X1 U294 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n845), .B1(n1097), .B2(\mem[12][6] ), 
        .ZN(n1091) );
  INV_X1 U296 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n845), .B1(n1097), .B2(\mem[12][7] ), 
        .ZN(n1090) );
  INV_X1 U298 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n844), .B1(n1088), .B2(\mem[13][0] ), 
        .ZN(n1089) );
  INV_X1 U300 ( .A(n1087), .ZN(n784) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n844), .B1(n1088), .B2(\mem[13][1] ), 
        .ZN(n1087) );
  INV_X1 U302 ( .A(n1086), .ZN(n783) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n844), .B1(n1088), .B2(\mem[13][2] ), 
        .ZN(n1086) );
  INV_X1 U304 ( .A(n1085), .ZN(n782) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n844), .B1(n1088), .B2(\mem[13][3] ), 
        .ZN(n1085) );
  INV_X1 U306 ( .A(n1084), .ZN(n781) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n844), .B1(n1088), .B2(\mem[13][4] ), 
        .ZN(n1084) );
  INV_X1 U308 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n844), .B1(n1088), .B2(\mem[13][5] ), 
        .ZN(n1083) );
  INV_X1 U310 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n844), .B1(n1088), .B2(\mem[13][6] ), 
        .ZN(n1082) );
  INV_X1 U312 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n844), .B1(n1088), .B2(\mem[13][7] ), 
        .ZN(n1081) );
  INV_X1 U314 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n843), .B1(n1079), .B2(\mem[14][0] ), 
        .ZN(n1080) );
  INV_X1 U316 ( .A(n1078), .ZN(n776) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n843), .B1(n1079), .B2(\mem[14][1] ), 
        .ZN(n1078) );
  INV_X1 U318 ( .A(n1077), .ZN(n775) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n843), .B1(n1079), .B2(\mem[14][2] ), 
        .ZN(n1077) );
  INV_X1 U320 ( .A(n1076), .ZN(n774) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n843), .B1(n1079), .B2(\mem[14][3] ), 
        .ZN(n1076) );
  INV_X1 U322 ( .A(n1075), .ZN(n773) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n843), .B1(n1079), .B2(\mem[14][4] ), 
        .ZN(n1075) );
  INV_X1 U324 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n843), .B1(n1079), .B2(\mem[14][5] ), 
        .ZN(n1074) );
  INV_X1 U326 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n843), .B1(n1079), .B2(\mem[14][6] ), 
        .ZN(n1073) );
  INV_X1 U328 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n843), .B1(n1079), .B2(\mem[14][7] ), 
        .ZN(n1072) );
  INV_X1 U330 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U331 ( .A1(data_in[0]), .A2(n842), .B1(n1070), .B2(\mem[15][0] ), 
        .ZN(n1071) );
  INV_X1 U332 ( .A(n1069), .ZN(n768) );
  AOI22_X1 U333 ( .A1(data_in[1]), .A2(n842), .B1(n1070), .B2(\mem[15][1] ), 
        .ZN(n1069) );
  INV_X1 U334 ( .A(n1068), .ZN(n767) );
  AOI22_X1 U335 ( .A1(data_in[2]), .A2(n842), .B1(n1070), .B2(\mem[15][2] ), 
        .ZN(n1068) );
  INV_X1 U336 ( .A(n1067), .ZN(n766) );
  AOI22_X1 U337 ( .A1(data_in[3]), .A2(n842), .B1(n1070), .B2(\mem[15][3] ), 
        .ZN(n1067) );
  INV_X1 U338 ( .A(n1066), .ZN(n765) );
  AOI22_X1 U339 ( .A1(data_in[4]), .A2(n842), .B1(n1070), .B2(\mem[15][4] ), 
        .ZN(n1066) );
  INV_X1 U340 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U341 ( .A1(data_in[5]), .A2(n842), .B1(n1070), .B2(\mem[15][5] ), 
        .ZN(n1065) );
  INV_X1 U342 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U343 ( .A1(data_in[6]), .A2(n842), .B1(n1070), .B2(\mem[15][6] ), 
        .ZN(n1064) );
  INV_X1 U344 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U345 ( .A1(data_in[7]), .A2(n842), .B1(n1070), .B2(\mem[15][7] ), 
        .ZN(n1063) );
  INV_X1 U346 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U347 ( .A1(data_in[0]), .A2(n841), .B1(n1061), .B2(\mem[16][0] ), 
        .ZN(n1062) );
  INV_X1 U348 ( .A(n1060), .ZN(n760) );
  AOI22_X1 U349 ( .A1(data_in[1]), .A2(n841), .B1(n1061), .B2(\mem[16][1] ), 
        .ZN(n1060) );
  INV_X1 U350 ( .A(n1059), .ZN(n759) );
  AOI22_X1 U351 ( .A1(data_in[2]), .A2(n841), .B1(n1061), .B2(\mem[16][2] ), 
        .ZN(n1059) );
  INV_X1 U352 ( .A(n1058), .ZN(n758) );
  AOI22_X1 U353 ( .A1(data_in[3]), .A2(n841), .B1(n1061), .B2(\mem[16][3] ), 
        .ZN(n1058) );
  INV_X1 U354 ( .A(n1057), .ZN(n757) );
  AOI22_X1 U355 ( .A1(data_in[4]), .A2(n841), .B1(n1061), .B2(\mem[16][4] ), 
        .ZN(n1057) );
  INV_X1 U356 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U357 ( .A1(data_in[5]), .A2(n841), .B1(n1061), .B2(\mem[16][5] ), 
        .ZN(n1056) );
  INV_X1 U358 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U359 ( .A1(data_in[6]), .A2(n841), .B1(n1061), .B2(\mem[16][6] ), 
        .ZN(n1055) );
  INV_X1 U360 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U361 ( .A1(data_in[7]), .A2(n841), .B1(n1061), .B2(\mem[16][7] ), 
        .ZN(n1054) );
  INV_X1 U362 ( .A(n1052), .ZN(n753) );
  AOI22_X1 U363 ( .A1(data_in[0]), .A2(n840), .B1(n1051), .B2(\mem[17][0] ), 
        .ZN(n1052) );
  INV_X1 U364 ( .A(n1050), .ZN(n752) );
  AOI22_X1 U365 ( .A1(data_in[1]), .A2(n840), .B1(n1051), .B2(\mem[17][1] ), 
        .ZN(n1050) );
  INV_X1 U366 ( .A(n1049), .ZN(n751) );
  AOI22_X1 U367 ( .A1(data_in[2]), .A2(n840), .B1(n1051), .B2(\mem[17][2] ), 
        .ZN(n1049) );
  INV_X1 U368 ( .A(n1048), .ZN(n750) );
  AOI22_X1 U369 ( .A1(data_in[3]), .A2(n840), .B1(n1051), .B2(\mem[17][3] ), 
        .ZN(n1048) );
  INV_X1 U370 ( .A(n1047), .ZN(n749) );
  AOI22_X1 U371 ( .A1(data_in[4]), .A2(n840), .B1(n1051), .B2(\mem[17][4] ), 
        .ZN(n1047) );
  INV_X1 U372 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U373 ( .A1(data_in[5]), .A2(n840), .B1(n1051), .B2(\mem[17][5] ), 
        .ZN(n1046) );
  INV_X1 U374 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U375 ( .A1(data_in[6]), .A2(n840), .B1(n1051), .B2(\mem[17][6] ), 
        .ZN(n1045) );
  INV_X1 U376 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U377 ( .A1(data_in[7]), .A2(n840), .B1(n1051), .B2(\mem[17][7] ), 
        .ZN(n1044) );
  INV_X1 U378 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U379 ( .A1(data_in[0]), .A2(n839), .B1(n1042), .B2(\mem[18][0] ), 
        .ZN(n1043) );
  INV_X1 U380 ( .A(n1041), .ZN(n744) );
  AOI22_X1 U381 ( .A1(data_in[1]), .A2(n839), .B1(n1042), .B2(\mem[18][1] ), 
        .ZN(n1041) );
  INV_X1 U382 ( .A(n1040), .ZN(n743) );
  AOI22_X1 U383 ( .A1(data_in[2]), .A2(n839), .B1(n1042), .B2(\mem[18][2] ), 
        .ZN(n1040) );
  INV_X1 U384 ( .A(n1039), .ZN(n742) );
  AOI22_X1 U385 ( .A1(data_in[3]), .A2(n839), .B1(n1042), .B2(\mem[18][3] ), 
        .ZN(n1039) );
  INV_X1 U386 ( .A(n1038), .ZN(n741) );
  AOI22_X1 U387 ( .A1(data_in[4]), .A2(n839), .B1(n1042), .B2(\mem[18][4] ), 
        .ZN(n1038) );
  INV_X1 U388 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U389 ( .A1(data_in[5]), .A2(n839), .B1(n1042), .B2(\mem[18][5] ), 
        .ZN(n1037) );
  INV_X1 U390 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U391 ( .A1(data_in[6]), .A2(n839), .B1(n1042), .B2(\mem[18][6] ), 
        .ZN(n1036) );
  INV_X1 U392 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U393 ( .A1(data_in[7]), .A2(n839), .B1(n1042), .B2(\mem[18][7] ), 
        .ZN(n1035) );
  INV_X1 U394 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U395 ( .A1(data_in[0]), .A2(n838), .B1(n1033), .B2(\mem[19][0] ), 
        .ZN(n1034) );
  INV_X1 U396 ( .A(n1032), .ZN(n736) );
  AOI22_X1 U397 ( .A1(data_in[1]), .A2(n838), .B1(n1033), .B2(\mem[19][1] ), 
        .ZN(n1032) );
  INV_X1 U398 ( .A(n1031), .ZN(n735) );
  AOI22_X1 U399 ( .A1(data_in[2]), .A2(n838), .B1(n1033), .B2(\mem[19][2] ), 
        .ZN(n1031) );
  INV_X1 U400 ( .A(n1030), .ZN(n734) );
  AOI22_X1 U401 ( .A1(data_in[3]), .A2(n838), .B1(n1033), .B2(\mem[19][3] ), 
        .ZN(n1030) );
  INV_X1 U402 ( .A(n1029), .ZN(n733) );
  AOI22_X1 U403 ( .A1(data_in[4]), .A2(n838), .B1(n1033), .B2(\mem[19][4] ), 
        .ZN(n1029) );
  INV_X1 U404 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U405 ( .A1(data_in[5]), .A2(n838), .B1(n1033), .B2(\mem[19][5] ), 
        .ZN(n1028) );
  INV_X1 U406 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U407 ( .A1(data_in[6]), .A2(n838), .B1(n1033), .B2(\mem[19][6] ), 
        .ZN(n1027) );
  INV_X1 U408 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U409 ( .A1(data_in[7]), .A2(n838), .B1(n1033), .B2(\mem[19][7] ), 
        .ZN(n1026) );
  INV_X1 U410 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U411 ( .A1(data_in[0]), .A2(n837), .B1(n1024), .B2(\mem[20][0] ), 
        .ZN(n1025) );
  INV_X1 U412 ( .A(n1023), .ZN(n728) );
  AOI22_X1 U413 ( .A1(data_in[1]), .A2(n837), .B1(n1024), .B2(\mem[20][1] ), 
        .ZN(n1023) );
  INV_X1 U414 ( .A(n1022), .ZN(n727) );
  AOI22_X1 U415 ( .A1(data_in[2]), .A2(n837), .B1(n1024), .B2(\mem[20][2] ), 
        .ZN(n1022) );
  INV_X1 U416 ( .A(n1021), .ZN(n726) );
  AOI22_X1 U417 ( .A1(data_in[3]), .A2(n837), .B1(n1024), .B2(\mem[20][3] ), 
        .ZN(n1021) );
  INV_X1 U418 ( .A(n1020), .ZN(n725) );
  AOI22_X1 U419 ( .A1(data_in[4]), .A2(n837), .B1(n1024), .B2(\mem[20][4] ), 
        .ZN(n1020) );
  INV_X1 U420 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U421 ( .A1(data_in[5]), .A2(n837), .B1(n1024), .B2(\mem[20][5] ), 
        .ZN(n1019) );
  INV_X1 U422 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U423 ( .A1(data_in[6]), .A2(n837), .B1(n1024), .B2(\mem[20][6] ), 
        .ZN(n1018) );
  INV_X1 U424 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U425 ( .A1(data_in[7]), .A2(n837), .B1(n1024), .B2(\mem[20][7] ), 
        .ZN(n1017) );
  INV_X1 U426 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U427 ( .A1(data_in[0]), .A2(n836), .B1(n1015), .B2(\mem[21][0] ), 
        .ZN(n1016) );
  INV_X1 U428 ( .A(n1014), .ZN(n720) );
  AOI22_X1 U429 ( .A1(data_in[1]), .A2(n836), .B1(n1015), .B2(\mem[21][1] ), 
        .ZN(n1014) );
  INV_X1 U430 ( .A(n1013), .ZN(n719) );
  AOI22_X1 U431 ( .A1(data_in[2]), .A2(n836), .B1(n1015), .B2(\mem[21][2] ), 
        .ZN(n1013) );
  INV_X1 U432 ( .A(n1012), .ZN(n718) );
  AOI22_X1 U433 ( .A1(data_in[3]), .A2(n836), .B1(n1015), .B2(\mem[21][3] ), 
        .ZN(n1012) );
  INV_X1 U434 ( .A(n1011), .ZN(n717) );
  AOI22_X1 U435 ( .A1(data_in[4]), .A2(n836), .B1(n1015), .B2(\mem[21][4] ), 
        .ZN(n1011) );
  INV_X1 U436 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U437 ( .A1(data_in[5]), .A2(n836), .B1(n1015), .B2(\mem[21][5] ), 
        .ZN(n1010) );
  INV_X1 U438 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U439 ( .A1(data_in[6]), .A2(n836), .B1(n1015), .B2(\mem[21][6] ), 
        .ZN(n1009) );
  INV_X1 U440 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U441 ( .A1(data_in[7]), .A2(n836), .B1(n1015), .B2(\mem[21][7] ), 
        .ZN(n1008) );
  INV_X1 U442 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U443 ( .A1(data_in[0]), .A2(n835), .B1(n1006), .B2(\mem[22][0] ), 
        .ZN(n1007) );
  INV_X1 U444 ( .A(n1005), .ZN(n712) );
  AOI22_X1 U445 ( .A1(data_in[1]), .A2(n835), .B1(n1006), .B2(\mem[22][1] ), 
        .ZN(n1005) );
  INV_X1 U446 ( .A(n1004), .ZN(n711) );
  AOI22_X1 U447 ( .A1(data_in[2]), .A2(n835), .B1(n1006), .B2(\mem[22][2] ), 
        .ZN(n1004) );
  INV_X1 U448 ( .A(n1003), .ZN(n710) );
  AOI22_X1 U449 ( .A1(data_in[3]), .A2(n835), .B1(n1006), .B2(\mem[22][3] ), 
        .ZN(n1003) );
  INV_X1 U450 ( .A(n1002), .ZN(n709) );
  AOI22_X1 U451 ( .A1(data_in[4]), .A2(n835), .B1(n1006), .B2(\mem[22][4] ), 
        .ZN(n1002) );
  INV_X1 U452 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U453 ( .A1(data_in[5]), .A2(n835), .B1(n1006), .B2(\mem[22][5] ), 
        .ZN(n1001) );
  INV_X1 U454 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U455 ( .A1(data_in[6]), .A2(n835), .B1(n1006), .B2(\mem[22][6] ), 
        .ZN(n1000) );
  INV_X1 U456 ( .A(n999), .ZN(n706) );
  AOI22_X1 U457 ( .A1(data_in[7]), .A2(n835), .B1(n1006), .B2(\mem[22][7] ), 
        .ZN(n999) );
  INV_X1 U458 ( .A(n998), .ZN(n705) );
  AOI22_X1 U459 ( .A1(data_in[0]), .A2(n834), .B1(n997), .B2(\mem[23][0] ), 
        .ZN(n998) );
  INV_X1 U460 ( .A(n996), .ZN(n704) );
  AOI22_X1 U461 ( .A1(data_in[1]), .A2(n834), .B1(n997), .B2(\mem[23][1] ), 
        .ZN(n996) );
  INV_X1 U462 ( .A(n995), .ZN(n703) );
  AOI22_X1 U463 ( .A1(data_in[2]), .A2(n834), .B1(n997), .B2(\mem[23][2] ), 
        .ZN(n995) );
  INV_X1 U464 ( .A(n994), .ZN(n702) );
  AOI22_X1 U465 ( .A1(data_in[3]), .A2(n834), .B1(n997), .B2(\mem[23][3] ), 
        .ZN(n994) );
  INV_X1 U466 ( .A(n993), .ZN(n701) );
  AOI22_X1 U467 ( .A1(data_in[4]), .A2(n834), .B1(n997), .B2(\mem[23][4] ), 
        .ZN(n993) );
  INV_X1 U468 ( .A(n992), .ZN(n700) );
  AOI22_X1 U469 ( .A1(data_in[5]), .A2(n834), .B1(n997), .B2(\mem[23][5] ), 
        .ZN(n992) );
  INV_X1 U470 ( .A(n991), .ZN(n699) );
  AOI22_X1 U471 ( .A1(data_in[6]), .A2(n834), .B1(n997), .B2(\mem[23][6] ), 
        .ZN(n991) );
  INV_X1 U472 ( .A(n990), .ZN(n698) );
  AOI22_X1 U473 ( .A1(data_in[7]), .A2(n834), .B1(n997), .B2(\mem[23][7] ), 
        .ZN(n990) );
  INV_X1 U474 ( .A(n989), .ZN(n697) );
  AOI22_X1 U475 ( .A1(data_in[0]), .A2(n833), .B1(n988), .B2(\mem[24][0] ), 
        .ZN(n989) );
  INV_X1 U476 ( .A(n987), .ZN(n696) );
  AOI22_X1 U477 ( .A1(data_in[1]), .A2(n833), .B1(n988), .B2(\mem[24][1] ), 
        .ZN(n987) );
  INV_X1 U478 ( .A(n986), .ZN(n695) );
  AOI22_X1 U479 ( .A1(data_in[2]), .A2(n833), .B1(n988), .B2(\mem[24][2] ), 
        .ZN(n986) );
  INV_X1 U480 ( .A(n985), .ZN(n694) );
  AOI22_X1 U481 ( .A1(data_in[3]), .A2(n833), .B1(n988), .B2(\mem[24][3] ), 
        .ZN(n985) );
  INV_X1 U482 ( .A(n984), .ZN(n693) );
  AOI22_X1 U483 ( .A1(data_in[4]), .A2(n833), .B1(n988), .B2(\mem[24][4] ), 
        .ZN(n984) );
  INV_X1 U484 ( .A(n983), .ZN(n692) );
  AOI22_X1 U485 ( .A1(data_in[5]), .A2(n833), .B1(n988), .B2(\mem[24][5] ), 
        .ZN(n983) );
  INV_X1 U486 ( .A(n982), .ZN(n691) );
  AOI22_X1 U487 ( .A1(data_in[6]), .A2(n833), .B1(n988), .B2(\mem[24][6] ), 
        .ZN(n982) );
  INV_X1 U488 ( .A(n981), .ZN(n690) );
  AOI22_X1 U489 ( .A1(data_in[7]), .A2(n833), .B1(n988), .B2(\mem[24][7] ), 
        .ZN(n981) );
  INV_X1 U490 ( .A(n979), .ZN(n689) );
  AOI22_X1 U491 ( .A1(data_in[0]), .A2(n832), .B1(n978), .B2(\mem[25][0] ), 
        .ZN(n979) );
  INV_X1 U492 ( .A(n977), .ZN(n688) );
  AOI22_X1 U493 ( .A1(data_in[1]), .A2(n832), .B1(n978), .B2(\mem[25][1] ), 
        .ZN(n977) );
  INV_X1 U494 ( .A(n976), .ZN(n687) );
  AOI22_X1 U495 ( .A1(data_in[2]), .A2(n832), .B1(n978), .B2(\mem[25][2] ), 
        .ZN(n976) );
  INV_X1 U496 ( .A(n975), .ZN(n686) );
  AOI22_X1 U497 ( .A1(data_in[3]), .A2(n832), .B1(n978), .B2(\mem[25][3] ), 
        .ZN(n975) );
  INV_X1 U498 ( .A(n974), .ZN(n685) );
  AOI22_X1 U499 ( .A1(data_in[4]), .A2(n832), .B1(n978), .B2(\mem[25][4] ), 
        .ZN(n974) );
  INV_X1 U500 ( .A(n973), .ZN(n684) );
  AOI22_X1 U501 ( .A1(data_in[5]), .A2(n832), .B1(n978), .B2(\mem[25][5] ), 
        .ZN(n973) );
  INV_X1 U502 ( .A(n972), .ZN(n683) );
  AOI22_X1 U503 ( .A1(data_in[6]), .A2(n832), .B1(n978), .B2(\mem[25][6] ), 
        .ZN(n972) );
  INV_X1 U504 ( .A(n971), .ZN(n682) );
  AOI22_X1 U505 ( .A1(data_in[7]), .A2(n832), .B1(n978), .B2(\mem[25][7] ), 
        .ZN(n971) );
  INV_X1 U506 ( .A(n970), .ZN(n681) );
  AOI22_X1 U507 ( .A1(data_in[0]), .A2(n831), .B1(n969), .B2(\mem[26][0] ), 
        .ZN(n970) );
  INV_X1 U508 ( .A(n968), .ZN(n680) );
  AOI22_X1 U509 ( .A1(data_in[1]), .A2(n831), .B1(n969), .B2(\mem[26][1] ), 
        .ZN(n968) );
  INV_X1 U510 ( .A(n967), .ZN(n679) );
  AOI22_X1 U511 ( .A1(data_in[2]), .A2(n831), .B1(n969), .B2(\mem[26][2] ), 
        .ZN(n967) );
  INV_X1 U512 ( .A(n966), .ZN(n678) );
  AOI22_X1 U513 ( .A1(data_in[3]), .A2(n831), .B1(n969), .B2(\mem[26][3] ), 
        .ZN(n966) );
  INV_X1 U514 ( .A(n965), .ZN(n677) );
  AOI22_X1 U515 ( .A1(data_in[4]), .A2(n831), .B1(n969), .B2(\mem[26][4] ), 
        .ZN(n965) );
  INV_X1 U516 ( .A(n964), .ZN(n676) );
  AOI22_X1 U517 ( .A1(data_in[5]), .A2(n831), .B1(n969), .B2(\mem[26][5] ), 
        .ZN(n964) );
  INV_X1 U518 ( .A(n963), .ZN(n675) );
  AOI22_X1 U519 ( .A1(data_in[6]), .A2(n831), .B1(n969), .B2(\mem[26][6] ), 
        .ZN(n963) );
  INV_X1 U520 ( .A(n962), .ZN(n674) );
  AOI22_X1 U521 ( .A1(data_in[7]), .A2(n831), .B1(n969), .B2(\mem[26][7] ), 
        .ZN(n962) );
  INV_X1 U522 ( .A(n961), .ZN(n673) );
  AOI22_X1 U523 ( .A1(data_in[0]), .A2(n830), .B1(n960), .B2(\mem[27][0] ), 
        .ZN(n961) );
  INV_X1 U524 ( .A(n959), .ZN(n672) );
  AOI22_X1 U525 ( .A1(data_in[1]), .A2(n830), .B1(n960), .B2(\mem[27][1] ), 
        .ZN(n959) );
  INV_X1 U526 ( .A(n958), .ZN(n671) );
  AOI22_X1 U527 ( .A1(data_in[2]), .A2(n830), .B1(n960), .B2(\mem[27][2] ), 
        .ZN(n958) );
  INV_X1 U528 ( .A(n957), .ZN(n670) );
  AOI22_X1 U529 ( .A1(data_in[3]), .A2(n830), .B1(n960), .B2(\mem[27][3] ), 
        .ZN(n957) );
  INV_X1 U530 ( .A(n956), .ZN(n669) );
  AOI22_X1 U531 ( .A1(data_in[4]), .A2(n830), .B1(n960), .B2(\mem[27][4] ), 
        .ZN(n956) );
  INV_X1 U532 ( .A(n955), .ZN(n668) );
  AOI22_X1 U533 ( .A1(data_in[5]), .A2(n830), .B1(n960), .B2(\mem[27][5] ), 
        .ZN(n955) );
  INV_X1 U534 ( .A(n954), .ZN(n667) );
  AOI22_X1 U535 ( .A1(data_in[6]), .A2(n830), .B1(n960), .B2(\mem[27][6] ), 
        .ZN(n954) );
  INV_X1 U536 ( .A(n953), .ZN(n666) );
  AOI22_X1 U537 ( .A1(data_in[7]), .A2(n830), .B1(n960), .B2(\mem[27][7] ), 
        .ZN(n953) );
  INV_X1 U538 ( .A(n952), .ZN(n665) );
  AOI22_X1 U539 ( .A1(data_in[0]), .A2(n829), .B1(n951), .B2(\mem[28][0] ), 
        .ZN(n952) );
  INV_X1 U540 ( .A(n950), .ZN(n664) );
  AOI22_X1 U541 ( .A1(data_in[1]), .A2(n829), .B1(n951), .B2(\mem[28][1] ), 
        .ZN(n950) );
  INV_X1 U542 ( .A(n949), .ZN(n663) );
  AOI22_X1 U543 ( .A1(data_in[2]), .A2(n829), .B1(n951), .B2(\mem[28][2] ), 
        .ZN(n949) );
  INV_X1 U544 ( .A(n948), .ZN(n662) );
  AOI22_X1 U545 ( .A1(data_in[3]), .A2(n829), .B1(n951), .B2(\mem[28][3] ), 
        .ZN(n948) );
  INV_X1 U546 ( .A(n947), .ZN(n661) );
  AOI22_X1 U547 ( .A1(data_in[4]), .A2(n829), .B1(n951), .B2(\mem[28][4] ), 
        .ZN(n947) );
  INV_X1 U548 ( .A(n946), .ZN(n660) );
  AOI22_X1 U549 ( .A1(data_in[5]), .A2(n829), .B1(n951), .B2(\mem[28][5] ), 
        .ZN(n946) );
  INV_X1 U550 ( .A(n945), .ZN(n659) );
  AOI22_X1 U551 ( .A1(data_in[6]), .A2(n829), .B1(n951), .B2(\mem[28][6] ), 
        .ZN(n945) );
  INV_X1 U552 ( .A(n944), .ZN(n658) );
  AOI22_X1 U553 ( .A1(data_in[7]), .A2(n829), .B1(n951), .B2(\mem[28][7] ), 
        .ZN(n944) );
  INV_X1 U554 ( .A(n943), .ZN(n657) );
  AOI22_X1 U555 ( .A1(data_in[0]), .A2(n828), .B1(n942), .B2(\mem[29][0] ), 
        .ZN(n943) );
  INV_X1 U556 ( .A(n941), .ZN(n656) );
  AOI22_X1 U557 ( .A1(data_in[1]), .A2(n828), .B1(n942), .B2(\mem[29][1] ), 
        .ZN(n941) );
  INV_X1 U558 ( .A(n940), .ZN(n655) );
  AOI22_X1 U559 ( .A1(data_in[2]), .A2(n828), .B1(n942), .B2(\mem[29][2] ), 
        .ZN(n940) );
  INV_X1 U560 ( .A(n939), .ZN(n654) );
  AOI22_X1 U561 ( .A1(data_in[3]), .A2(n828), .B1(n942), .B2(\mem[29][3] ), 
        .ZN(n939) );
  INV_X1 U562 ( .A(n938), .ZN(n653) );
  AOI22_X1 U563 ( .A1(data_in[4]), .A2(n828), .B1(n942), .B2(\mem[29][4] ), 
        .ZN(n938) );
  INV_X1 U564 ( .A(n937), .ZN(n652) );
  AOI22_X1 U565 ( .A1(data_in[5]), .A2(n828), .B1(n942), .B2(\mem[29][5] ), 
        .ZN(n937) );
  INV_X1 U566 ( .A(n936), .ZN(n651) );
  AOI22_X1 U567 ( .A1(data_in[6]), .A2(n828), .B1(n942), .B2(\mem[29][6] ), 
        .ZN(n936) );
  INV_X1 U568 ( .A(n935), .ZN(n650) );
  AOI22_X1 U569 ( .A1(data_in[7]), .A2(n828), .B1(n942), .B2(\mem[29][7] ), 
        .ZN(n935) );
  INV_X1 U570 ( .A(n934), .ZN(n649) );
  AOI22_X1 U571 ( .A1(data_in[0]), .A2(n827), .B1(n933), .B2(\mem[30][0] ), 
        .ZN(n934) );
  INV_X1 U572 ( .A(n932), .ZN(n648) );
  AOI22_X1 U573 ( .A1(data_in[1]), .A2(n827), .B1(n933), .B2(\mem[30][1] ), 
        .ZN(n932) );
  INV_X1 U574 ( .A(n931), .ZN(n647) );
  AOI22_X1 U575 ( .A1(data_in[2]), .A2(n827), .B1(n933), .B2(\mem[30][2] ), 
        .ZN(n931) );
  INV_X1 U576 ( .A(n930), .ZN(n646) );
  AOI22_X1 U577 ( .A1(data_in[3]), .A2(n827), .B1(n933), .B2(\mem[30][3] ), 
        .ZN(n930) );
  INV_X1 U578 ( .A(n929), .ZN(n645) );
  AOI22_X1 U579 ( .A1(data_in[4]), .A2(n827), .B1(n933), .B2(\mem[30][4] ), 
        .ZN(n929) );
  INV_X1 U580 ( .A(n928), .ZN(n644) );
  AOI22_X1 U581 ( .A1(data_in[5]), .A2(n827), .B1(n933), .B2(\mem[30][5] ), 
        .ZN(n928) );
  INV_X1 U582 ( .A(n927), .ZN(n643) );
  AOI22_X1 U583 ( .A1(data_in[6]), .A2(n827), .B1(n933), .B2(\mem[30][6] ), 
        .ZN(n927) );
  INV_X1 U584 ( .A(n926), .ZN(n642) );
  AOI22_X1 U585 ( .A1(data_in[7]), .A2(n827), .B1(n933), .B2(\mem[30][7] ), 
        .ZN(n926) );
  INV_X1 U586 ( .A(n925), .ZN(n641) );
  AOI22_X1 U587 ( .A1(data_in[0]), .A2(n826), .B1(n924), .B2(\mem[31][0] ), 
        .ZN(n925) );
  INV_X1 U588 ( .A(n923), .ZN(n640) );
  AOI22_X1 U589 ( .A1(data_in[1]), .A2(n826), .B1(n924), .B2(\mem[31][1] ), 
        .ZN(n923) );
  INV_X1 U590 ( .A(n922), .ZN(n639) );
  AOI22_X1 U591 ( .A1(data_in[2]), .A2(n826), .B1(n924), .B2(\mem[31][2] ), 
        .ZN(n922) );
  INV_X1 U592 ( .A(n921), .ZN(n638) );
  AOI22_X1 U593 ( .A1(data_in[3]), .A2(n826), .B1(n924), .B2(\mem[31][3] ), 
        .ZN(n921) );
  INV_X1 U594 ( .A(n920), .ZN(n637) );
  AOI22_X1 U595 ( .A1(data_in[4]), .A2(n826), .B1(n924), .B2(\mem[31][4] ), 
        .ZN(n920) );
  INV_X1 U596 ( .A(n919), .ZN(n636) );
  AOI22_X1 U597 ( .A1(data_in[5]), .A2(n826), .B1(n924), .B2(\mem[31][5] ), 
        .ZN(n919) );
  INV_X1 U598 ( .A(n918), .ZN(n635) );
  AOI22_X1 U599 ( .A1(data_in[6]), .A2(n826), .B1(n924), .B2(\mem[31][6] ), 
        .ZN(n918) );
  INV_X1 U600 ( .A(n917), .ZN(n634) );
  AOI22_X1 U601 ( .A1(data_in[7]), .A2(n826), .B1(n924), .B2(\mem[31][7] ), 
        .ZN(n917) );
  MUX2_X1 U602 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n614), .Z(n4) );
  MUX2_X1 U603 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n614), .Z(n5) );
  MUX2_X1 U604 ( .A(n5), .B(n4), .S(n611), .Z(n6) );
  MUX2_X1 U605 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n614), .Z(n7) );
  MUX2_X1 U606 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n614), .Z(n8) );
  MUX2_X1 U607 ( .A(n8), .B(n7), .S(n611), .Z(n9) );
  MUX2_X1 U608 ( .A(n9), .B(n6), .S(n609), .Z(n10) );
  MUX2_X1 U609 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n614), .Z(n11) );
  MUX2_X1 U610 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n614), .Z(n12) );
  MUX2_X1 U611 ( .A(n12), .B(n11), .S(n611), .Z(n13) );
  MUX2_X1 U612 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n614), .Z(n14) );
  MUX2_X1 U613 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n614), .Z(n15) );
  MUX2_X1 U614 ( .A(n15), .B(n14), .S(n611), .Z(n16) );
  MUX2_X1 U615 ( .A(n16), .B(n13), .S(N12), .Z(n17) );
  MUX2_X1 U616 ( .A(n17), .B(n10), .S(N13), .Z(n18) );
  MUX2_X1 U617 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n615), .Z(n19) );
  MUX2_X1 U618 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n615), .Z(n20) );
  MUX2_X1 U619 ( .A(n20), .B(n19), .S(n611), .Z(n21) );
  MUX2_X1 U620 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n615), .Z(n22) );
  MUX2_X1 U621 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n615), .Z(n23) );
  MUX2_X1 U622 ( .A(n23), .B(n22), .S(n612), .Z(n24) );
  MUX2_X1 U623 ( .A(n24), .B(n21), .S(N12), .Z(n25) );
  MUX2_X1 U624 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n615), .Z(n26) );
  MUX2_X1 U625 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n615), .Z(n27) );
  MUX2_X1 U626 ( .A(n27), .B(n26), .S(n611), .Z(n28) );
  MUX2_X1 U627 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n615), .Z(n29) );
  MUX2_X1 U628 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n615), .Z(n30) );
  MUX2_X1 U629 ( .A(n30), .B(n29), .S(N11), .Z(n31) );
  MUX2_X1 U630 ( .A(n31), .B(n28), .S(n610), .Z(n32) );
  MUX2_X1 U631 ( .A(n32), .B(n25), .S(N13), .Z(n33) );
  MUX2_X1 U632 ( .A(n33), .B(n18), .S(N14), .Z(N22) );
  MUX2_X1 U633 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n615), .Z(n34) );
  MUX2_X1 U634 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n615), .Z(n35) );
  MUX2_X1 U635 ( .A(n35), .B(n34), .S(n611), .Z(n36) );
  MUX2_X1 U636 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n615), .Z(n37) );
  MUX2_X1 U637 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n615), .Z(n38) );
  MUX2_X1 U638 ( .A(n38), .B(n37), .S(n611), .Z(n39) );
  MUX2_X1 U639 ( .A(n39), .B(n36), .S(n610), .Z(n40) );
  MUX2_X1 U640 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n616), .Z(n41) );
  MUX2_X1 U641 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n616), .Z(n42) );
  MUX2_X1 U642 ( .A(n42), .B(n41), .S(n611), .Z(n43) );
  MUX2_X1 U643 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n616), .Z(n44) );
  MUX2_X1 U644 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n616), .Z(n45) );
  MUX2_X1 U645 ( .A(n45), .B(n44), .S(n612), .Z(n46) );
  MUX2_X1 U646 ( .A(n46), .B(n43), .S(n609), .Z(n47) );
  MUX2_X1 U647 ( .A(n47), .B(n40), .S(N13), .Z(n48) );
  MUX2_X1 U648 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n616), .Z(n49) );
  MUX2_X1 U649 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n616), .Z(n50) );
  MUX2_X1 U650 ( .A(n50), .B(n49), .S(n611), .Z(n51) );
  MUX2_X1 U651 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n616), .Z(n52) );
  MUX2_X1 U652 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n616), .Z(n53) );
  MUX2_X1 U653 ( .A(n53), .B(n52), .S(n613), .Z(n54) );
  MUX2_X1 U654 ( .A(n54), .B(n51), .S(N12), .Z(n55) );
  MUX2_X1 U655 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n616), .Z(n56) );
  MUX2_X1 U656 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n616), .Z(n57) );
  MUX2_X1 U657 ( .A(n57), .B(n56), .S(n611), .Z(n58) );
  MUX2_X1 U658 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n616), .Z(n59) );
  MUX2_X1 U659 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n616), .Z(n60) );
  MUX2_X1 U660 ( .A(n60), .B(n59), .S(n611), .Z(n61) );
  MUX2_X1 U661 ( .A(n61), .B(n58), .S(n609), .Z(n62) );
  MUX2_X1 U662 ( .A(n62), .B(n55), .S(N13), .Z(n63) );
  MUX2_X1 U663 ( .A(n63), .B(n48), .S(N14), .Z(N21) );
  MUX2_X1 U664 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n617), .Z(n64) );
  MUX2_X1 U665 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n617), .Z(n65) );
  MUX2_X1 U666 ( .A(n65), .B(n64), .S(n612), .Z(n66) );
  MUX2_X1 U667 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n617), .Z(n67) );
  MUX2_X1 U668 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n617), .Z(n68) );
  MUX2_X1 U669 ( .A(n68), .B(n67), .S(n612), .Z(n69) );
  MUX2_X1 U670 ( .A(n69), .B(n66), .S(n609), .Z(n70) );
  MUX2_X1 U671 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n617), .Z(n71) );
  MUX2_X1 U672 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n617), .Z(n72) );
  MUX2_X1 U673 ( .A(n72), .B(n71), .S(n612), .Z(n73) );
  MUX2_X1 U674 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n617), .Z(n74) );
  MUX2_X1 U675 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n617), .Z(n75) );
  MUX2_X1 U676 ( .A(n75), .B(n74), .S(n612), .Z(n76) );
  MUX2_X1 U677 ( .A(n76), .B(n73), .S(n609), .Z(n77) );
  MUX2_X1 U678 ( .A(n77), .B(n70), .S(N13), .Z(n78) );
  MUX2_X1 U679 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n617), .Z(n79) );
  MUX2_X1 U680 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n617), .Z(n80) );
  MUX2_X1 U681 ( .A(n80), .B(n79), .S(n612), .Z(n81) );
  MUX2_X1 U682 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n617), .Z(n82) );
  MUX2_X1 U683 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n617), .Z(n83) );
  MUX2_X1 U684 ( .A(n83), .B(n82), .S(n612), .Z(n84) );
  MUX2_X1 U685 ( .A(n84), .B(n81), .S(n609), .Z(n85) );
  MUX2_X1 U686 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n618), .Z(n86) );
  MUX2_X1 U687 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n618), .Z(n87) );
  MUX2_X1 U688 ( .A(n87), .B(n86), .S(n612), .Z(n88) );
  MUX2_X1 U689 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n618), .Z(n89) );
  MUX2_X1 U690 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n618), .Z(n90) );
  MUX2_X1 U691 ( .A(n90), .B(n89), .S(n612), .Z(n91) );
  MUX2_X1 U692 ( .A(n91), .B(n88), .S(n609), .Z(n92) );
  MUX2_X1 U693 ( .A(n92), .B(n85), .S(N13), .Z(n93) );
  MUX2_X1 U694 ( .A(n93), .B(n78), .S(N14), .Z(N20) );
  MUX2_X1 U695 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n618), .Z(n94) );
  MUX2_X1 U696 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n618), .Z(n95) );
  MUX2_X1 U697 ( .A(n95), .B(n94), .S(n612), .Z(n96) );
  MUX2_X1 U698 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n618), .Z(n97) );
  MUX2_X1 U699 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n618), .Z(n98) );
  MUX2_X1 U700 ( .A(n98), .B(n97), .S(n612), .Z(n99) );
  MUX2_X1 U701 ( .A(n99), .B(n96), .S(n609), .Z(n100) );
  MUX2_X1 U702 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n618), .Z(n101) );
  MUX2_X1 U703 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n618), .Z(n102) );
  MUX2_X1 U704 ( .A(n102), .B(n101), .S(n612), .Z(n103) );
  MUX2_X1 U705 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n618), .Z(n104) );
  MUX2_X1 U706 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n618), .Z(n105) );
  MUX2_X1 U707 ( .A(n105), .B(n104), .S(n612), .Z(n106) );
  MUX2_X1 U708 ( .A(n106), .B(n103), .S(n609), .Z(n107) );
  MUX2_X1 U709 ( .A(n107), .B(n100), .S(N13), .Z(n108) );
  MUX2_X1 U710 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n622), .Z(n109) );
  MUX2_X1 U711 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n622), .Z(n110) );
  MUX2_X1 U712 ( .A(n110), .B(n109), .S(n613), .Z(n111) );
  MUX2_X1 U713 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n623), .Z(n112) );
  MUX2_X1 U714 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n622), .Z(n113) );
  MUX2_X1 U715 ( .A(n113), .B(n112), .S(n613), .Z(n114) );
  MUX2_X1 U716 ( .A(n114), .B(n111), .S(n609), .Z(n115) );
  MUX2_X1 U717 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n623), .Z(n116) );
  MUX2_X1 U718 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n623), .Z(n117) );
  MUX2_X1 U719 ( .A(n117), .B(n116), .S(n613), .Z(n118) );
  MUX2_X1 U720 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n623), .Z(n119) );
  MUX2_X1 U721 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n623), .Z(n120) );
  MUX2_X1 U722 ( .A(n120), .B(n119), .S(n613), .Z(n121) );
  MUX2_X1 U723 ( .A(n121), .B(n118), .S(n609), .Z(n122) );
  MUX2_X1 U724 ( .A(n122), .B(n115), .S(N13), .Z(n123) );
  MUX2_X1 U725 ( .A(n123), .B(n108), .S(N14), .Z(N19) );
  MUX2_X1 U726 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n622), .Z(n124) );
  MUX2_X1 U727 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n622), .Z(n125) );
  MUX2_X1 U728 ( .A(n125), .B(n124), .S(n613), .Z(n126) );
  MUX2_X1 U729 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n622), .Z(n127) );
  MUX2_X1 U730 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n128) );
  MUX2_X1 U731 ( .A(n128), .B(n127), .S(n613), .Z(n129) );
  MUX2_X1 U732 ( .A(n129), .B(n126), .S(n609), .Z(n130) );
  MUX2_X1 U733 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n614), .Z(n131) );
  MUX2_X1 U734 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n622), .Z(n132) );
  MUX2_X1 U735 ( .A(n132), .B(n131), .S(n613), .Z(n133) );
  MUX2_X1 U736 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n622), .Z(n134) );
  MUX2_X1 U737 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(N10), .Z(n135) );
  MUX2_X1 U738 ( .A(n135), .B(n134), .S(n613), .Z(n136) );
  MUX2_X1 U739 ( .A(n136), .B(n133), .S(n609), .Z(n137) );
  MUX2_X1 U740 ( .A(n137), .B(n130), .S(N13), .Z(n138) );
  MUX2_X1 U741 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n614), .Z(n139) );
  MUX2_X1 U742 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n623), .Z(n140) );
  MUX2_X1 U743 ( .A(n140), .B(n139), .S(n613), .Z(n141) );
  MUX2_X1 U744 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n614), .Z(n142) );
  MUX2_X1 U745 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n143) );
  MUX2_X1 U746 ( .A(n143), .B(n142), .S(n613), .Z(n144) );
  MUX2_X1 U747 ( .A(n144), .B(n141), .S(n609), .Z(n145) );
  MUX2_X1 U748 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n614), .Z(n146) );
  MUX2_X1 U749 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n147) );
  MUX2_X1 U750 ( .A(n147), .B(n146), .S(n613), .Z(n148) );
  MUX2_X1 U751 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n623), .Z(n149) );
  MUX2_X1 U752 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n150) );
  MUX2_X1 U753 ( .A(n150), .B(n149), .S(n613), .Z(n151) );
  MUX2_X1 U754 ( .A(n151), .B(n148), .S(n609), .Z(n152) );
  MUX2_X1 U755 ( .A(n152), .B(n145), .S(N13), .Z(n153) );
  MUX2_X1 U756 ( .A(n153), .B(n138), .S(N14), .Z(N18) );
  MUX2_X1 U757 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n619), .Z(n154) );
  MUX2_X1 U758 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n619), .Z(n155) );
  MUX2_X1 U759 ( .A(n155), .B(n154), .S(n611), .Z(n156) );
  MUX2_X1 U760 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n619), .Z(n157) );
  MUX2_X1 U761 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n619), .Z(n158) );
  MUX2_X1 U762 ( .A(n158), .B(n157), .S(n613), .Z(n159) );
  MUX2_X1 U763 ( .A(n159), .B(n156), .S(n610), .Z(n160) );
  MUX2_X1 U764 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n619), .Z(n161) );
  MUX2_X1 U765 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n619), .Z(n162) );
  MUX2_X1 U766 ( .A(n162), .B(n161), .S(N11), .Z(n163) );
  MUX2_X1 U767 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n619), .Z(n164) );
  MUX2_X1 U768 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n619), .Z(n165) );
  MUX2_X1 U769 ( .A(n165), .B(n164), .S(n613), .Z(n166) );
  MUX2_X1 U770 ( .A(n166), .B(n163), .S(n610), .Z(n167) );
  MUX2_X1 U771 ( .A(n167), .B(n160), .S(N13), .Z(n168) );
  MUX2_X1 U772 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n619), .Z(n169) );
  MUX2_X1 U773 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n619), .Z(n170) );
  MUX2_X1 U774 ( .A(n170), .B(n169), .S(n613), .Z(n171) );
  MUX2_X1 U775 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n619), .Z(n172) );
  MUX2_X1 U776 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n619), .Z(n173) );
  MUX2_X1 U777 ( .A(n173), .B(n172), .S(n611), .Z(n174) );
  MUX2_X1 U778 ( .A(n174), .B(n171), .S(n610), .Z(n175) );
  MUX2_X1 U779 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n620), .Z(n176) );
  MUX2_X1 U780 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n620), .Z(n177) );
  MUX2_X1 U781 ( .A(n177), .B(n176), .S(n612), .Z(n178) );
  MUX2_X1 U782 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n620), .Z(n179) );
  MUX2_X1 U783 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n620), .Z(n180) );
  MUX2_X1 U784 ( .A(n180), .B(n179), .S(n612), .Z(n181) );
  MUX2_X1 U785 ( .A(n181), .B(n178), .S(n610), .Z(n182) );
  MUX2_X1 U786 ( .A(n182), .B(n175), .S(N13), .Z(n183) );
  MUX2_X1 U787 ( .A(n183), .B(n168), .S(N14), .Z(N17) );
  MUX2_X1 U788 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n620), .Z(n184) );
  MUX2_X1 U789 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n620), .Z(n185) );
  MUX2_X1 U790 ( .A(n185), .B(n184), .S(n612), .Z(n186) );
  MUX2_X1 U791 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n620), .Z(n187) );
  MUX2_X1 U792 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n620), .Z(n188) );
  MUX2_X1 U793 ( .A(n188), .B(n187), .S(n611), .Z(n189) );
  MUX2_X1 U794 ( .A(n189), .B(n186), .S(n610), .Z(n190) );
  MUX2_X1 U795 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n620), .Z(n191) );
  MUX2_X1 U796 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n620), .Z(n192) );
  MUX2_X1 U797 ( .A(n192), .B(n191), .S(n612), .Z(n193) );
  MUX2_X1 U798 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n620), .Z(n194) );
  MUX2_X1 U799 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n620), .Z(n195) );
  MUX2_X1 U800 ( .A(n195), .B(n194), .S(n611), .Z(n196) );
  MUX2_X1 U801 ( .A(n196), .B(n193), .S(n610), .Z(n197) );
  MUX2_X1 U802 ( .A(n197), .B(n190), .S(N13), .Z(n198) );
  MUX2_X1 U803 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n621), .Z(n199) );
  MUX2_X1 U804 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n621), .Z(n200) );
  MUX2_X1 U805 ( .A(n200), .B(n199), .S(n613), .Z(n201) );
  MUX2_X1 U806 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n621), .Z(n202) );
  MUX2_X1 U807 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n621), .Z(n203) );
  MUX2_X1 U808 ( .A(n203), .B(n202), .S(N11), .Z(n204) );
  MUX2_X1 U809 ( .A(n204), .B(n201), .S(n610), .Z(n205) );
  MUX2_X1 U810 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n621), .Z(n206) );
  MUX2_X1 U811 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n621), .Z(n207) );
  MUX2_X1 U812 ( .A(n207), .B(n206), .S(n613), .Z(n208) );
  MUX2_X1 U813 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n621), .Z(n209) );
  MUX2_X1 U814 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n621), .Z(n210) );
  MUX2_X1 U815 ( .A(n210), .B(n209), .S(n612), .Z(n211) );
  MUX2_X1 U816 ( .A(n211), .B(n208), .S(n610), .Z(n212) );
  MUX2_X1 U817 ( .A(n212), .B(n205), .S(N13), .Z(n213) );
  MUX2_X1 U818 ( .A(n213), .B(n198), .S(N14), .Z(N16) );
  MUX2_X1 U819 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n621), .Z(n214) );
  MUX2_X1 U820 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n621), .Z(n215) );
  MUX2_X1 U821 ( .A(n215), .B(n214), .S(n612), .Z(n216) );
  MUX2_X1 U822 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n621), .Z(n217) );
  MUX2_X1 U823 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n621), .Z(n218) );
  MUX2_X1 U824 ( .A(n218), .B(n217), .S(n612), .Z(n219) );
  MUX2_X1 U825 ( .A(n219), .B(n216), .S(n610), .Z(n220) );
  MUX2_X1 U826 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n622), .Z(n221) );
  MUX2_X1 U827 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n623), .Z(n222) );
  MUX2_X1 U828 ( .A(n222), .B(n221), .S(n611), .Z(n223) );
  MUX2_X1 U829 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n622), .Z(n224) );
  MUX2_X1 U830 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n622), .Z(n225) );
  MUX2_X1 U831 ( .A(n225), .B(n224), .S(N11), .Z(n226) );
  MUX2_X1 U832 ( .A(n226), .B(n223), .S(n610), .Z(n227) );
  MUX2_X1 U833 ( .A(n227), .B(n220), .S(N13), .Z(n228) );
  MUX2_X1 U834 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n623), .Z(n229) );
  MUX2_X1 U835 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n622), .Z(n595) );
  MUX2_X1 U836 ( .A(n595), .B(n229), .S(n611), .Z(n596) );
  MUX2_X1 U837 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n623), .Z(n597) );
  MUX2_X1 U838 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n623), .Z(n598) );
  MUX2_X1 U839 ( .A(n598), .B(n597), .S(N11), .Z(n599) );
  MUX2_X1 U840 ( .A(n599), .B(n596), .S(n610), .Z(n600) );
  MUX2_X1 U841 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n622), .Z(n601) );
  MUX2_X1 U842 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n622), .Z(n602) );
  MUX2_X1 U843 ( .A(n602), .B(n601), .S(n613), .Z(n603) );
  MUX2_X1 U844 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n623), .Z(n604) );
  MUX2_X1 U845 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n623), .Z(n605) );
  MUX2_X1 U846 ( .A(n605), .B(n604), .S(n613), .Z(n606) );
  MUX2_X1 U847 ( .A(n606), .B(n603), .S(n610), .Z(n607) );
  MUX2_X1 U848 ( .A(n607), .B(n600), .S(N13), .Z(n608) );
  MUX2_X1 U849 ( .A(n608), .B(n228), .S(N14), .Z(N15) );
  CLKBUF_X1 U850 ( .A(N11), .Z(n611) );
  INV_X1 U851 ( .A(N10), .ZN(n624) );
  INV_X1 U852 ( .A(N11), .ZN(n625) );
  INV_X1 U853 ( .A(data_in[0]), .ZN(n626) );
  INV_X1 U854 ( .A(data_in[1]), .ZN(n627) );
  INV_X1 U855 ( .A(data_in[2]), .ZN(n628) );
  INV_X1 U856 ( .A(data_in[3]), .ZN(n629) );
  INV_X1 U857 ( .A(data_in[4]), .ZN(n630) );
  INV_X1 U858 ( .A(data_in[5]), .ZN(n631) );
  INV_X1 U859 ( .A(data_in[6]), .ZN(n632) );
  INV_X1 U860 ( .A(data_in[7]), .ZN(n633) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_8 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n631), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n632), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n633), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n634), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n635), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n636), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n637), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n638), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n639), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n640), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n641), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n642), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n643), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n644), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n645), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n646), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n647), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n648), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n649), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n650), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n651), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n652), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n653), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n654), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n655), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n656), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n657), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n658), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n659), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n660), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n661), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n662), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n663), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n664), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n665), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n666), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n667), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n668), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n669), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n670), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n671), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n672), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n673), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n674), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n675), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n676), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n677), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n678), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n679), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n680), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n681), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n682), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n683), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n684), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n685), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n686), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n687), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n688), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n689), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n690), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n691), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n692), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n693), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n694), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n695), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n696), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n697), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n698), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n699), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n700), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n701), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n702), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n703), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n704), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n705), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n706), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n707), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n708), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n709), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n710), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n711), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n712), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n713), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n714), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n715), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n716), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n717), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n718), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n719), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n720), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n721), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n722), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n723), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n724), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n725), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n726), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n727), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n728), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n729), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n730), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n731), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n732), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n733), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n734), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n735), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n736), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n737), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n738), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n739), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n740), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n741), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n742), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n743), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n744), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n745), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n746), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n747), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n748), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n749), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n750), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n751), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n752), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n753), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n754), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n755), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n756), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n757), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n758), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n759), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n760), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n761), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n762), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n763), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n764), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n765), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n766), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n767), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n768), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n769), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n770), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n771), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n772), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n773), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n774), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n775), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n776), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n777), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n778), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n779), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n780), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n781), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n782), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n783), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n784), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n785), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n786), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n787), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n788), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n789), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n790), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n791), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n792), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n793), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n794), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n795), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n796), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n797), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n798), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n799), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n800), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n801), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n802), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n803), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n804), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n805), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n806), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n807), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n808), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n809), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n810), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n811), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n812), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n813), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n814), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n815), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n816), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n817), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n818), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n819), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n820), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n821), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n822), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n850), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n851), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n852), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n853), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n854), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n855), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n856), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n857), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n858), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n859), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n860), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n861), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n862), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n863), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n864), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n865), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n866), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n867), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n868), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n869), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n870), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n871), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n872), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n873), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n874), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n875), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n876), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n877), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n878), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n879), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n880), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n881), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n882), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n883), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n884), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n885), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n886), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n887), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n888), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n889), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n890), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n891), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n892), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n893), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n894), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n895), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n896), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n897), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n898), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n899), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n900), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n901), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n902), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n903), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n904), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n905), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n906), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n907), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n908), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n909), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n910), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n911), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n912), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n913), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  BUF_X1 U3 ( .A(n619), .Z(n612) );
  BUF_X1 U4 ( .A(n620), .Z(n617) );
  BUF_X1 U5 ( .A(n620), .Z(n618) );
  BUF_X1 U6 ( .A(n620), .Z(n616) );
  BUF_X1 U7 ( .A(n619), .Z(n613) );
  BUF_X1 U8 ( .A(n619), .Z(n614) );
  BUF_X1 U9 ( .A(n619), .Z(n615) );
  BUF_X1 U10 ( .A(N11), .Z(n610) );
  BUF_X1 U11 ( .A(N11), .Z(n611) );
  BUF_X1 U12 ( .A(N10), .Z(n620) );
  BUF_X1 U13 ( .A(N10), .Z(n619) );
  NOR3_X1 U14 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1205) );
  NOR3_X1 U15 ( .A1(N11), .A2(N12), .A3(n621), .ZN(n1194) );
  NOR3_X1 U16 ( .A1(N10), .A2(N12), .A3(n622), .ZN(n1184) );
  NOR3_X1 U17 ( .A1(n621), .A2(N12), .A3(n622), .ZN(n1174) );
  INV_X1 U18 ( .A(n1131), .ZN(n846) );
  INV_X1 U19 ( .A(n1121), .ZN(n845) );
  INV_X1 U20 ( .A(n1112), .ZN(n844) );
  INV_X1 U21 ( .A(n1103), .ZN(n843) );
  INV_X1 U22 ( .A(n1058), .ZN(n838) );
  INV_X1 U23 ( .A(n1048), .ZN(n837) );
  INV_X1 U24 ( .A(n1039), .ZN(n836) );
  INV_X1 U25 ( .A(n1030), .ZN(n835) );
  INV_X1 U26 ( .A(n985), .ZN(n830) );
  INV_X1 U27 ( .A(n975), .ZN(n829) );
  INV_X1 U28 ( .A(n966), .ZN(n828) );
  INV_X1 U29 ( .A(n957), .ZN(n827) );
  INV_X1 U30 ( .A(n948), .ZN(n826) );
  INV_X1 U31 ( .A(n939), .ZN(n825) );
  INV_X1 U32 ( .A(n930), .ZN(n824) );
  INV_X1 U33 ( .A(n921), .ZN(n823) );
  INV_X1 U34 ( .A(n1094), .ZN(n842) );
  INV_X1 U35 ( .A(n1085), .ZN(n841) );
  INV_X1 U36 ( .A(n1076), .ZN(n840) );
  INV_X1 U37 ( .A(n1067), .ZN(n839) );
  INV_X1 U38 ( .A(n1021), .ZN(n834) );
  INV_X1 U39 ( .A(n1012), .ZN(n833) );
  INV_X1 U40 ( .A(n1003), .ZN(n832) );
  INV_X1 U41 ( .A(n994), .ZN(n831) );
  BUF_X1 U42 ( .A(N12), .Z(n607) );
  BUF_X1 U43 ( .A(N12), .Z(n608) );
  INV_X1 U44 ( .A(N13), .ZN(n848) );
  AND3_X1 U45 ( .A1(n621), .A2(n622), .A3(N12), .ZN(n1164) );
  AND3_X1 U46 ( .A1(N10), .A2(n622), .A3(N12), .ZN(n1154) );
  AND3_X1 U47 ( .A1(N11), .A2(n621), .A3(N12), .ZN(n1144) );
  AND3_X1 U48 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1134) );
  INV_X1 U49 ( .A(N14), .ZN(n849) );
  NAND2_X1 U50 ( .A1(n1194), .A2(n1204), .ZN(n1203) );
  NAND2_X1 U51 ( .A1(n1184), .A2(n1204), .ZN(n1193) );
  NAND2_X1 U52 ( .A1(n1174), .A2(n1204), .ZN(n1183) );
  NAND2_X1 U53 ( .A1(n1164), .A2(n1204), .ZN(n1173) );
  NAND2_X1 U54 ( .A1(n1154), .A2(n1204), .ZN(n1163) );
  NAND2_X1 U55 ( .A1(n1144), .A2(n1204), .ZN(n1153) );
  NAND2_X1 U56 ( .A1(n1134), .A2(n1204), .ZN(n1143) );
  NAND2_X1 U57 ( .A1(n1205), .A2(n1204), .ZN(n1214) );
  NAND2_X1 U58 ( .A1(n1123), .A2(n1205), .ZN(n1131) );
  NAND2_X1 U59 ( .A1(n1123), .A2(n1194), .ZN(n1121) );
  NAND2_X1 U60 ( .A1(n1123), .A2(n1184), .ZN(n1112) );
  NAND2_X1 U61 ( .A1(n1123), .A2(n1174), .ZN(n1103) );
  NAND2_X1 U62 ( .A1(n1050), .A2(n1205), .ZN(n1058) );
  NAND2_X1 U63 ( .A1(n1050), .A2(n1194), .ZN(n1048) );
  NAND2_X1 U64 ( .A1(n1050), .A2(n1184), .ZN(n1039) );
  NAND2_X1 U65 ( .A1(n1050), .A2(n1174), .ZN(n1030) );
  NAND2_X1 U66 ( .A1(n977), .A2(n1205), .ZN(n985) );
  NAND2_X1 U67 ( .A1(n977), .A2(n1194), .ZN(n975) );
  NAND2_X1 U68 ( .A1(n977), .A2(n1184), .ZN(n966) );
  NAND2_X1 U69 ( .A1(n977), .A2(n1174), .ZN(n957) );
  NAND2_X1 U70 ( .A1(n1123), .A2(n1164), .ZN(n1094) );
  NAND2_X1 U71 ( .A1(n1123), .A2(n1154), .ZN(n1085) );
  NAND2_X1 U72 ( .A1(n1123), .A2(n1144), .ZN(n1076) );
  NAND2_X1 U73 ( .A1(n1123), .A2(n1134), .ZN(n1067) );
  NAND2_X1 U74 ( .A1(n1050), .A2(n1164), .ZN(n1021) );
  NAND2_X1 U75 ( .A1(n1050), .A2(n1154), .ZN(n1012) );
  NAND2_X1 U76 ( .A1(n1050), .A2(n1144), .ZN(n1003) );
  NAND2_X1 U77 ( .A1(n1050), .A2(n1134), .ZN(n994) );
  NAND2_X1 U78 ( .A1(n977), .A2(n1164), .ZN(n948) );
  NAND2_X1 U79 ( .A1(n977), .A2(n1154), .ZN(n939) );
  NAND2_X1 U80 ( .A1(n977), .A2(n1144), .ZN(n930) );
  NAND2_X1 U81 ( .A1(n977), .A2(n1134), .ZN(n921) );
  AND3_X1 U82 ( .A1(n848), .A2(n849), .A3(n1133), .ZN(n1204) );
  AND3_X1 U83 ( .A1(N13), .A2(n1133), .A3(N14), .ZN(n977) );
  AND3_X1 U84 ( .A1(n1133), .A2(n849), .A3(N13), .ZN(n1123) );
  AND3_X1 U85 ( .A1(n1133), .A2(n848), .A3(N14), .ZN(n1050) );
  NOR2_X1 U86 ( .A1(n847), .A2(addr[5]), .ZN(n1133) );
  INV_X1 U87 ( .A(wr_en), .ZN(n847) );
  OAI21_X1 U88 ( .B1(n623), .B2(n1173), .A(n1172), .ZN(n881) );
  NAND2_X1 U89 ( .A1(\mem[4][0] ), .A2(n1173), .ZN(n1172) );
  OAI21_X1 U90 ( .B1(n624), .B2(n1173), .A(n1171), .ZN(n880) );
  NAND2_X1 U91 ( .A1(\mem[4][1] ), .A2(n1173), .ZN(n1171) );
  OAI21_X1 U92 ( .B1(n625), .B2(n1173), .A(n1170), .ZN(n879) );
  NAND2_X1 U93 ( .A1(\mem[4][2] ), .A2(n1173), .ZN(n1170) );
  OAI21_X1 U94 ( .B1(n626), .B2(n1173), .A(n1169), .ZN(n878) );
  NAND2_X1 U95 ( .A1(\mem[4][3] ), .A2(n1173), .ZN(n1169) );
  OAI21_X1 U96 ( .B1(n627), .B2(n1173), .A(n1168), .ZN(n877) );
  NAND2_X1 U97 ( .A1(\mem[4][4] ), .A2(n1173), .ZN(n1168) );
  OAI21_X1 U98 ( .B1(n628), .B2(n1173), .A(n1167), .ZN(n876) );
  NAND2_X1 U99 ( .A1(\mem[4][5] ), .A2(n1173), .ZN(n1167) );
  OAI21_X1 U100 ( .B1(n629), .B2(n1173), .A(n1166), .ZN(n875) );
  NAND2_X1 U101 ( .A1(\mem[4][6] ), .A2(n1173), .ZN(n1166) );
  OAI21_X1 U102 ( .B1(n630), .B2(n1173), .A(n1165), .ZN(n874) );
  NAND2_X1 U103 ( .A1(\mem[4][7] ), .A2(n1173), .ZN(n1165) );
  OAI21_X1 U104 ( .B1(n623), .B2(n1153), .A(n1152), .ZN(n865) );
  NAND2_X1 U105 ( .A1(\mem[6][0] ), .A2(n1153), .ZN(n1152) );
  OAI21_X1 U106 ( .B1(n624), .B2(n1153), .A(n1151), .ZN(n864) );
  NAND2_X1 U107 ( .A1(\mem[6][1] ), .A2(n1153), .ZN(n1151) );
  OAI21_X1 U108 ( .B1(n625), .B2(n1153), .A(n1150), .ZN(n863) );
  NAND2_X1 U109 ( .A1(\mem[6][2] ), .A2(n1153), .ZN(n1150) );
  OAI21_X1 U110 ( .B1(n626), .B2(n1153), .A(n1149), .ZN(n862) );
  NAND2_X1 U111 ( .A1(\mem[6][3] ), .A2(n1153), .ZN(n1149) );
  OAI21_X1 U112 ( .B1(n627), .B2(n1153), .A(n1148), .ZN(n861) );
  NAND2_X1 U113 ( .A1(\mem[6][4] ), .A2(n1153), .ZN(n1148) );
  OAI21_X1 U114 ( .B1(n628), .B2(n1153), .A(n1147), .ZN(n860) );
  NAND2_X1 U115 ( .A1(\mem[6][5] ), .A2(n1153), .ZN(n1147) );
  OAI21_X1 U116 ( .B1(n629), .B2(n1153), .A(n1146), .ZN(n859) );
  NAND2_X1 U117 ( .A1(\mem[6][6] ), .A2(n1153), .ZN(n1146) );
  OAI21_X1 U118 ( .B1(n630), .B2(n1153), .A(n1145), .ZN(n858) );
  NAND2_X1 U119 ( .A1(\mem[6][7] ), .A2(n1153), .ZN(n1145) );
  OAI21_X1 U120 ( .B1(n623), .B2(n1143), .A(n1142), .ZN(n857) );
  NAND2_X1 U121 ( .A1(\mem[7][0] ), .A2(n1143), .ZN(n1142) );
  OAI21_X1 U122 ( .B1(n624), .B2(n1143), .A(n1141), .ZN(n856) );
  NAND2_X1 U123 ( .A1(\mem[7][1] ), .A2(n1143), .ZN(n1141) );
  OAI21_X1 U124 ( .B1(n625), .B2(n1143), .A(n1140), .ZN(n855) );
  NAND2_X1 U125 ( .A1(\mem[7][2] ), .A2(n1143), .ZN(n1140) );
  OAI21_X1 U126 ( .B1(n626), .B2(n1143), .A(n1139), .ZN(n854) );
  NAND2_X1 U127 ( .A1(\mem[7][3] ), .A2(n1143), .ZN(n1139) );
  OAI21_X1 U128 ( .B1(n627), .B2(n1143), .A(n1138), .ZN(n853) );
  NAND2_X1 U129 ( .A1(\mem[7][4] ), .A2(n1143), .ZN(n1138) );
  OAI21_X1 U130 ( .B1(n628), .B2(n1143), .A(n1137), .ZN(n852) );
  NAND2_X1 U131 ( .A1(\mem[7][5] ), .A2(n1143), .ZN(n1137) );
  OAI21_X1 U132 ( .B1(n629), .B2(n1143), .A(n1136), .ZN(n851) );
  NAND2_X1 U133 ( .A1(\mem[7][6] ), .A2(n1143), .ZN(n1136) );
  OAI21_X1 U134 ( .B1(n630), .B2(n1143), .A(n1135), .ZN(n850) );
  NAND2_X1 U135 ( .A1(\mem[7][7] ), .A2(n1143), .ZN(n1135) );
  OAI21_X1 U136 ( .B1(n623), .B2(n1203), .A(n1202), .ZN(n905) );
  NAND2_X1 U137 ( .A1(\mem[1][0] ), .A2(n1203), .ZN(n1202) );
  OAI21_X1 U138 ( .B1(n624), .B2(n1203), .A(n1201), .ZN(n904) );
  NAND2_X1 U139 ( .A1(\mem[1][1] ), .A2(n1203), .ZN(n1201) );
  OAI21_X1 U140 ( .B1(n625), .B2(n1203), .A(n1200), .ZN(n903) );
  NAND2_X1 U141 ( .A1(\mem[1][2] ), .A2(n1203), .ZN(n1200) );
  OAI21_X1 U142 ( .B1(n626), .B2(n1203), .A(n1199), .ZN(n902) );
  NAND2_X1 U143 ( .A1(\mem[1][3] ), .A2(n1203), .ZN(n1199) );
  OAI21_X1 U144 ( .B1(n627), .B2(n1203), .A(n1198), .ZN(n901) );
  NAND2_X1 U145 ( .A1(\mem[1][4] ), .A2(n1203), .ZN(n1198) );
  OAI21_X1 U146 ( .B1(n628), .B2(n1203), .A(n1197), .ZN(n900) );
  NAND2_X1 U147 ( .A1(\mem[1][5] ), .A2(n1203), .ZN(n1197) );
  OAI21_X1 U148 ( .B1(n629), .B2(n1203), .A(n1196), .ZN(n899) );
  NAND2_X1 U149 ( .A1(\mem[1][6] ), .A2(n1203), .ZN(n1196) );
  OAI21_X1 U150 ( .B1(n630), .B2(n1203), .A(n1195), .ZN(n898) );
  NAND2_X1 U151 ( .A1(\mem[1][7] ), .A2(n1203), .ZN(n1195) );
  OAI21_X1 U152 ( .B1(n623), .B2(n1193), .A(n1192), .ZN(n897) );
  NAND2_X1 U153 ( .A1(\mem[2][0] ), .A2(n1193), .ZN(n1192) );
  OAI21_X1 U154 ( .B1(n624), .B2(n1193), .A(n1191), .ZN(n896) );
  NAND2_X1 U155 ( .A1(\mem[2][1] ), .A2(n1193), .ZN(n1191) );
  OAI21_X1 U156 ( .B1(n625), .B2(n1193), .A(n1190), .ZN(n895) );
  NAND2_X1 U157 ( .A1(\mem[2][2] ), .A2(n1193), .ZN(n1190) );
  OAI21_X1 U158 ( .B1(n626), .B2(n1193), .A(n1189), .ZN(n894) );
  NAND2_X1 U159 ( .A1(\mem[2][3] ), .A2(n1193), .ZN(n1189) );
  OAI21_X1 U160 ( .B1(n627), .B2(n1193), .A(n1188), .ZN(n893) );
  NAND2_X1 U161 ( .A1(\mem[2][4] ), .A2(n1193), .ZN(n1188) );
  OAI21_X1 U162 ( .B1(n628), .B2(n1193), .A(n1187), .ZN(n892) );
  NAND2_X1 U163 ( .A1(\mem[2][5] ), .A2(n1193), .ZN(n1187) );
  OAI21_X1 U164 ( .B1(n629), .B2(n1193), .A(n1186), .ZN(n891) );
  NAND2_X1 U165 ( .A1(\mem[2][6] ), .A2(n1193), .ZN(n1186) );
  OAI21_X1 U166 ( .B1(n630), .B2(n1193), .A(n1185), .ZN(n890) );
  NAND2_X1 U167 ( .A1(\mem[2][7] ), .A2(n1193), .ZN(n1185) );
  OAI21_X1 U168 ( .B1(n623), .B2(n1183), .A(n1182), .ZN(n889) );
  NAND2_X1 U169 ( .A1(\mem[3][0] ), .A2(n1183), .ZN(n1182) );
  OAI21_X1 U170 ( .B1(n624), .B2(n1183), .A(n1181), .ZN(n888) );
  NAND2_X1 U171 ( .A1(\mem[3][1] ), .A2(n1183), .ZN(n1181) );
  OAI21_X1 U172 ( .B1(n625), .B2(n1183), .A(n1180), .ZN(n887) );
  NAND2_X1 U173 ( .A1(\mem[3][2] ), .A2(n1183), .ZN(n1180) );
  OAI21_X1 U174 ( .B1(n626), .B2(n1183), .A(n1179), .ZN(n886) );
  NAND2_X1 U175 ( .A1(\mem[3][3] ), .A2(n1183), .ZN(n1179) );
  OAI21_X1 U176 ( .B1(n627), .B2(n1183), .A(n1178), .ZN(n885) );
  NAND2_X1 U177 ( .A1(\mem[3][4] ), .A2(n1183), .ZN(n1178) );
  OAI21_X1 U178 ( .B1(n628), .B2(n1183), .A(n1177), .ZN(n884) );
  NAND2_X1 U179 ( .A1(\mem[3][5] ), .A2(n1183), .ZN(n1177) );
  OAI21_X1 U180 ( .B1(n629), .B2(n1183), .A(n1176), .ZN(n883) );
  NAND2_X1 U181 ( .A1(\mem[3][6] ), .A2(n1183), .ZN(n1176) );
  OAI21_X1 U182 ( .B1(n630), .B2(n1183), .A(n1175), .ZN(n882) );
  NAND2_X1 U183 ( .A1(\mem[3][7] ), .A2(n1183), .ZN(n1175) );
  OAI21_X1 U184 ( .B1(n623), .B2(n1163), .A(n1162), .ZN(n873) );
  NAND2_X1 U185 ( .A1(\mem[5][0] ), .A2(n1163), .ZN(n1162) );
  OAI21_X1 U186 ( .B1(n624), .B2(n1163), .A(n1161), .ZN(n872) );
  NAND2_X1 U187 ( .A1(\mem[5][1] ), .A2(n1163), .ZN(n1161) );
  OAI21_X1 U188 ( .B1(n625), .B2(n1163), .A(n1160), .ZN(n871) );
  NAND2_X1 U189 ( .A1(\mem[5][2] ), .A2(n1163), .ZN(n1160) );
  OAI21_X1 U190 ( .B1(n626), .B2(n1163), .A(n1159), .ZN(n870) );
  NAND2_X1 U191 ( .A1(\mem[5][3] ), .A2(n1163), .ZN(n1159) );
  OAI21_X1 U192 ( .B1(n627), .B2(n1163), .A(n1158), .ZN(n869) );
  NAND2_X1 U193 ( .A1(\mem[5][4] ), .A2(n1163), .ZN(n1158) );
  OAI21_X1 U194 ( .B1(n628), .B2(n1163), .A(n1157), .ZN(n868) );
  NAND2_X1 U195 ( .A1(\mem[5][5] ), .A2(n1163), .ZN(n1157) );
  OAI21_X1 U196 ( .B1(n629), .B2(n1163), .A(n1156), .ZN(n867) );
  NAND2_X1 U197 ( .A1(\mem[5][6] ), .A2(n1163), .ZN(n1156) );
  OAI21_X1 U198 ( .B1(n630), .B2(n1163), .A(n1155), .ZN(n866) );
  NAND2_X1 U199 ( .A1(\mem[5][7] ), .A2(n1163), .ZN(n1155) );
  OAI21_X1 U200 ( .B1(n1214), .B2(n623), .A(n1213), .ZN(n913) );
  NAND2_X1 U201 ( .A1(\mem[0][0] ), .A2(n1214), .ZN(n1213) );
  OAI21_X1 U202 ( .B1(n1214), .B2(n624), .A(n1212), .ZN(n912) );
  NAND2_X1 U203 ( .A1(\mem[0][1] ), .A2(n1214), .ZN(n1212) );
  OAI21_X1 U204 ( .B1(n1214), .B2(n625), .A(n1211), .ZN(n911) );
  NAND2_X1 U205 ( .A1(\mem[0][2] ), .A2(n1214), .ZN(n1211) );
  OAI21_X1 U206 ( .B1(n1214), .B2(n626), .A(n1210), .ZN(n910) );
  NAND2_X1 U207 ( .A1(\mem[0][3] ), .A2(n1214), .ZN(n1210) );
  OAI21_X1 U208 ( .B1(n1214), .B2(n627), .A(n1209), .ZN(n909) );
  NAND2_X1 U209 ( .A1(\mem[0][4] ), .A2(n1214), .ZN(n1209) );
  OAI21_X1 U210 ( .B1(n1214), .B2(n628), .A(n1208), .ZN(n908) );
  NAND2_X1 U211 ( .A1(\mem[0][5] ), .A2(n1214), .ZN(n1208) );
  OAI21_X1 U212 ( .B1(n1214), .B2(n629), .A(n1207), .ZN(n907) );
  NAND2_X1 U213 ( .A1(\mem[0][6] ), .A2(n1214), .ZN(n1207) );
  OAI21_X1 U214 ( .B1(n1214), .B2(n630), .A(n1206), .ZN(n906) );
  NAND2_X1 U215 ( .A1(\mem[0][7] ), .A2(n1214), .ZN(n1206) );
  INV_X1 U216 ( .A(n1132), .ZN(n822) );
  AOI22_X1 U217 ( .A1(data_in[0]), .A2(n846), .B1(n1131), .B2(\mem[8][0] ), 
        .ZN(n1132) );
  INV_X1 U218 ( .A(n1130), .ZN(n821) );
  AOI22_X1 U219 ( .A1(data_in[1]), .A2(n846), .B1(n1131), .B2(\mem[8][1] ), 
        .ZN(n1130) );
  INV_X1 U220 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U221 ( .A1(data_in[2]), .A2(n846), .B1(n1131), .B2(\mem[8][2] ), 
        .ZN(n1129) );
  INV_X1 U222 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U223 ( .A1(data_in[3]), .A2(n846), .B1(n1131), .B2(\mem[8][3] ), 
        .ZN(n1128) );
  INV_X1 U224 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U225 ( .A1(data_in[4]), .A2(n846), .B1(n1131), .B2(\mem[8][4] ), 
        .ZN(n1127) );
  INV_X1 U226 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U227 ( .A1(data_in[5]), .A2(n846), .B1(n1131), .B2(\mem[8][5] ), 
        .ZN(n1126) );
  INV_X1 U228 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U229 ( .A1(data_in[6]), .A2(n846), .B1(n1131), .B2(\mem[8][6] ), 
        .ZN(n1125) );
  INV_X1 U230 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U231 ( .A1(data_in[7]), .A2(n846), .B1(n1131), .B2(\mem[8][7] ), 
        .ZN(n1124) );
  INV_X1 U232 ( .A(n1122), .ZN(n814) );
  AOI22_X1 U233 ( .A1(data_in[0]), .A2(n845), .B1(n1121), .B2(\mem[9][0] ), 
        .ZN(n1122) );
  INV_X1 U234 ( .A(n1120), .ZN(n813) );
  AOI22_X1 U235 ( .A1(data_in[1]), .A2(n845), .B1(n1121), .B2(\mem[9][1] ), 
        .ZN(n1120) );
  INV_X1 U236 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U237 ( .A1(data_in[2]), .A2(n845), .B1(n1121), .B2(\mem[9][2] ), 
        .ZN(n1119) );
  INV_X1 U238 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U239 ( .A1(data_in[3]), .A2(n845), .B1(n1121), .B2(\mem[9][3] ), 
        .ZN(n1118) );
  INV_X1 U240 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U241 ( .A1(data_in[4]), .A2(n845), .B1(n1121), .B2(\mem[9][4] ), 
        .ZN(n1117) );
  INV_X1 U242 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U243 ( .A1(data_in[5]), .A2(n845), .B1(n1121), .B2(\mem[9][5] ), 
        .ZN(n1116) );
  INV_X1 U244 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U245 ( .A1(data_in[6]), .A2(n845), .B1(n1121), .B2(\mem[9][6] ), 
        .ZN(n1115) );
  INV_X1 U246 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U247 ( .A1(data_in[7]), .A2(n845), .B1(n1121), .B2(\mem[9][7] ), 
        .ZN(n1114) );
  INV_X1 U248 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U249 ( .A1(data_in[0]), .A2(n844), .B1(n1112), .B2(\mem[10][0] ), 
        .ZN(n1113) );
  INV_X1 U250 ( .A(n1111), .ZN(n805) );
  AOI22_X1 U251 ( .A1(data_in[1]), .A2(n844), .B1(n1112), .B2(\mem[10][1] ), 
        .ZN(n1111) );
  INV_X1 U252 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U253 ( .A1(data_in[2]), .A2(n844), .B1(n1112), .B2(\mem[10][2] ), 
        .ZN(n1110) );
  INV_X1 U254 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U255 ( .A1(data_in[3]), .A2(n844), .B1(n1112), .B2(\mem[10][3] ), 
        .ZN(n1109) );
  INV_X1 U256 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U257 ( .A1(data_in[4]), .A2(n844), .B1(n1112), .B2(\mem[10][4] ), 
        .ZN(n1108) );
  INV_X1 U258 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U259 ( .A1(data_in[5]), .A2(n844), .B1(n1112), .B2(\mem[10][5] ), 
        .ZN(n1107) );
  INV_X1 U260 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U261 ( .A1(data_in[6]), .A2(n844), .B1(n1112), .B2(\mem[10][6] ), 
        .ZN(n1106) );
  INV_X1 U262 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U263 ( .A1(data_in[7]), .A2(n844), .B1(n1112), .B2(\mem[10][7] ), 
        .ZN(n1105) );
  INV_X1 U264 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U265 ( .A1(data_in[0]), .A2(n843), .B1(n1103), .B2(\mem[11][0] ), 
        .ZN(n1104) );
  INV_X1 U266 ( .A(n1102), .ZN(n797) );
  AOI22_X1 U267 ( .A1(data_in[1]), .A2(n843), .B1(n1103), .B2(\mem[11][1] ), 
        .ZN(n1102) );
  INV_X1 U268 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U269 ( .A1(data_in[2]), .A2(n843), .B1(n1103), .B2(\mem[11][2] ), 
        .ZN(n1101) );
  INV_X1 U270 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U271 ( .A1(data_in[3]), .A2(n843), .B1(n1103), .B2(\mem[11][3] ), 
        .ZN(n1100) );
  INV_X1 U272 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U273 ( .A1(data_in[4]), .A2(n843), .B1(n1103), .B2(\mem[11][4] ), 
        .ZN(n1099) );
  INV_X1 U274 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U275 ( .A1(data_in[5]), .A2(n843), .B1(n1103), .B2(\mem[11][5] ), 
        .ZN(n1098) );
  INV_X1 U276 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U277 ( .A1(data_in[6]), .A2(n843), .B1(n1103), .B2(\mem[11][6] ), 
        .ZN(n1097) );
  INV_X1 U278 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U279 ( .A1(data_in[7]), .A2(n843), .B1(n1103), .B2(\mem[11][7] ), 
        .ZN(n1096) );
  INV_X1 U280 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U281 ( .A1(data_in[0]), .A2(n842), .B1(n1094), .B2(\mem[12][0] ), 
        .ZN(n1095) );
  INV_X1 U282 ( .A(n1093), .ZN(n789) );
  AOI22_X1 U283 ( .A1(data_in[1]), .A2(n842), .B1(n1094), .B2(\mem[12][1] ), 
        .ZN(n1093) );
  INV_X1 U284 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U285 ( .A1(data_in[2]), .A2(n842), .B1(n1094), .B2(\mem[12][2] ), 
        .ZN(n1092) );
  INV_X1 U286 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U287 ( .A1(data_in[3]), .A2(n842), .B1(n1094), .B2(\mem[12][3] ), 
        .ZN(n1091) );
  INV_X1 U288 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U289 ( .A1(data_in[4]), .A2(n842), .B1(n1094), .B2(\mem[12][4] ), 
        .ZN(n1090) );
  INV_X1 U290 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U291 ( .A1(data_in[5]), .A2(n842), .B1(n1094), .B2(\mem[12][5] ), 
        .ZN(n1089) );
  INV_X1 U292 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U293 ( .A1(data_in[6]), .A2(n842), .B1(n1094), .B2(\mem[12][6] ), 
        .ZN(n1088) );
  INV_X1 U294 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U295 ( .A1(data_in[7]), .A2(n842), .B1(n1094), .B2(\mem[12][7] ), 
        .ZN(n1087) );
  INV_X1 U296 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U297 ( .A1(data_in[0]), .A2(n841), .B1(n1085), .B2(\mem[13][0] ), 
        .ZN(n1086) );
  INV_X1 U298 ( .A(n1084), .ZN(n781) );
  AOI22_X1 U299 ( .A1(data_in[1]), .A2(n841), .B1(n1085), .B2(\mem[13][1] ), 
        .ZN(n1084) );
  INV_X1 U300 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U301 ( .A1(data_in[2]), .A2(n841), .B1(n1085), .B2(\mem[13][2] ), 
        .ZN(n1083) );
  INV_X1 U302 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U303 ( .A1(data_in[3]), .A2(n841), .B1(n1085), .B2(\mem[13][3] ), 
        .ZN(n1082) );
  INV_X1 U304 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U305 ( .A1(data_in[4]), .A2(n841), .B1(n1085), .B2(\mem[13][4] ), 
        .ZN(n1081) );
  INV_X1 U306 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U307 ( .A1(data_in[5]), .A2(n841), .B1(n1085), .B2(\mem[13][5] ), 
        .ZN(n1080) );
  INV_X1 U308 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U309 ( .A1(data_in[6]), .A2(n841), .B1(n1085), .B2(\mem[13][6] ), 
        .ZN(n1079) );
  INV_X1 U310 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U311 ( .A1(data_in[7]), .A2(n841), .B1(n1085), .B2(\mem[13][7] ), 
        .ZN(n1078) );
  INV_X1 U312 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U313 ( .A1(data_in[0]), .A2(n840), .B1(n1076), .B2(\mem[14][0] ), 
        .ZN(n1077) );
  INV_X1 U314 ( .A(n1075), .ZN(n773) );
  AOI22_X1 U315 ( .A1(data_in[1]), .A2(n840), .B1(n1076), .B2(\mem[14][1] ), 
        .ZN(n1075) );
  INV_X1 U316 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U317 ( .A1(data_in[2]), .A2(n840), .B1(n1076), .B2(\mem[14][2] ), 
        .ZN(n1074) );
  INV_X1 U318 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U319 ( .A1(data_in[3]), .A2(n840), .B1(n1076), .B2(\mem[14][3] ), 
        .ZN(n1073) );
  INV_X1 U320 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U321 ( .A1(data_in[4]), .A2(n840), .B1(n1076), .B2(\mem[14][4] ), 
        .ZN(n1072) );
  INV_X1 U322 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U323 ( .A1(data_in[5]), .A2(n840), .B1(n1076), .B2(\mem[14][5] ), 
        .ZN(n1071) );
  INV_X1 U324 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U325 ( .A1(data_in[6]), .A2(n840), .B1(n1076), .B2(\mem[14][6] ), 
        .ZN(n1070) );
  INV_X1 U326 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U327 ( .A1(data_in[7]), .A2(n840), .B1(n1076), .B2(\mem[14][7] ), 
        .ZN(n1069) );
  INV_X1 U328 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U329 ( .A1(data_in[0]), .A2(n839), .B1(n1067), .B2(\mem[15][0] ), 
        .ZN(n1068) );
  INV_X1 U330 ( .A(n1066), .ZN(n765) );
  AOI22_X1 U331 ( .A1(data_in[1]), .A2(n839), .B1(n1067), .B2(\mem[15][1] ), 
        .ZN(n1066) );
  INV_X1 U332 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U333 ( .A1(data_in[2]), .A2(n839), .B1(n1067), .B2(\mem[15][2] ), 
        .ZN(n1065) );
  INV_X1 U334 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U335 ( .A1(data_in[3]), .A2(n839), .B1(n1067), .B2(\mem[15][3] ), 
        .ZN(n1064) );
  INV_X1 U336 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U337 ( .A1(data_in[4]), .A2(n839), .B1(n1067), .B2(\mem[15][4] ), 
        .ZN(n1063) );
  INV_X1 U338 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U339 ( .A1(data_in[5]), .A2(n839), .B1(n1067), .B2(\mem[15][5] ), 
        .ZN(n1062) );
  INV_X1 U340 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U341 ( .A1(data_in[6]), .A2(n839), .B1(n1067), .B2(\mem[15][6] ), 
        .ZN(n1061) );
  INV_X1 U342 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U343 ( .A1(data_in[7]), .A2(n839), .B1(n1067), .B2(\mem[15][7] ), 
        .ZN(n1060) );
  INV_X1 U344 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U345 ( .A1(data_in[0]), .A2(n838), .B1(n1058), .B2(\mem[16][0] ), 
        .ZN(n1059) );
  INV_X1 U346 ( .A(n1057), .ZN(n757) );
  AOI22_X1 U347 ( .A1(data_in[1]), .A2(n838), .B1(n1058), .B2(\mem[16][1] ), 
        .ZN(n1057) );
  INV_X1 U348 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U349 ( .A1(data_in[2]), .A2(n838), .B1(n1058), .B2(\mem[16][2] ), 
        .ZN(n1056) );
  INV_X1 U350 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U351 ( .A1(data_in[3]), .A2(n838), .B1(n1058), .B2(\mem[16][3] ), 
        .ZN(n1055) );
  INV_X1 U352 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U353 ( .A1(data_in[4]), .A2(n838), .B1(n1058), .B2(\mem[16][4] ), 
        .ZN(n1054) );
  INV_X1 U354 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U355 ( .A1(data_in[5]), .A2(n838), .B1(n1058), .B2(\mem[16][5] ), 
        .ZN(n1053) );
  INV_X1 U356 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U357 ( .A1(data_in[6]), .A2(n838), .B1(n1058), .B2(\mem[16][6] ), 
        .ZN(n1052) );
  INV_X1 U358 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U359 ( .A1(data_in[7]), .A2(n838), .B1(n1058), .B2(\mem[16][7] ), 
        .ZN(n1051) );
  INV_X1 U360 ( .A(n1049), .ZN(n750) );
  AOI22_X1 U361 ( .A1(data_in[0]), .A2(n837), .B1(n1048), .B2(\mem[17][0] ), 
        .ZN(n1049) );
  INV_X1 U362 ( .A(n1047), .ZN(n749) );
  AOI22_X1 U363 ( .A1(data_in[1]), .A2(n837), .B1(n1048), .B2(\mem[17][1] ), 
        .ZN(n1047) );
  INV_X1 U364 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U365 ( .A1(data_in[2]), .A2(n837), .B1(n1048), .B2(\mem[17][2] ), 
        .ZN(n1046) );
  INV_X1 U366 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U367 ( .A1(data_in[3]), .A2(n837), .B1(n1048), .B2(\mem[17][3] ), 
        .ZN(n1045) );
  INV_X1 U368 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U369 ( .A1(data_in[4]), .A2(n837), .B1(n1048), .B2(\mem[17][4] ), 
        .ZN(n1044) );
  INV_X1 U370 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U371 ( .A1(data_in[5]), .A2(n837), .B1(n1048), .B2(\mem[17][5] ), 
        .ZN(n1043) );
  INV_X1 U372 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U373 ( .A1(data_in[6]), .A2(n837), .B1(n1048), .B2(\mem[17][6] ), 
        .ZN(n1042) );
  INV_X1 U374 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U375 ( .A1(data_in[7]), .A2(n837), .B1(n1048), .B2(\mem[17][7] ), 
        .ZN(n1041) );
  INV_X1 U376 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U377 ( .A1(data_in[0]), .A2(n836), .B1(n1039), .B2(\mem[18][0] ), 
        .ZN(n1040) );
  INV_X1 U378 ( .A(n1038), .ZN(n741) );
  AOI22_X1 U379 ( .A1(data_in[1]), .A2(n836), .B1(n1039), .B2(\mem[18][1] ), 
        .ZN(n1038) );
  INV_X1 U380 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U381 ( .A1(data_in[2]), .A2(n836), .B1(n1039), .B2(\mem[18][2] ), 
        .ZN(n1037) );
  INV_X1 U382 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U383 ( .A1(data_in[3]), .A2(n836), .B1(n1039), .B2(\mem[18][3] ), 
        .ZN(n1036) );
  INV_X1 U384 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U385 ( .A1(data_in[4]), .A2(n836), .B1(n1039), .B2(\mem[18][4] ), 
        .ZN(n1035) );
  INV_X1 U386 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U387 ( .A1(data_in[5]), .A2(n836), .B1(n1039), .B2(\mem[18][5] ), 
        .ZN(n1034) );
  INV_X1 U388 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U389 ( .A1(data_in[6]), .A2(n836), .B1(n1039), .B2(\mem[18][6] ), 
        .ZN(n1033) );
  INV_X1 U390 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U391 ( .A1(data_in[7]), .A2(n836), .B1(n1039), .B2(\mem[18][7] ), 
        .ZN(n1032) );
  INV_X1 U392 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U393 ( .A1(data_in[0]), .A2(n835), .B1(n1030), .B2(\mem[19][0] ), 
        .ZN(n1031) );
  INV_X1 U394 ( .A(n1029), .ZN(n733) );
  AOI22_X1 U395 ( .A1(data_in[1]), .A2(n835), .B1(n1030), .B2(\mem[19][1] ), 
        .ZN(n1029) );
  INV_X1 U396 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U397 ( .A1(data_in[2]), .A2(n835), .B1(n1030), .B2(\mem[19][2] ), 
        .ZN(n1028) );
  INV_X1 U398 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U399 ( .A1(data_in[3]), .A2(n835), .B1(n1030), .B2(\mem[19][3] ), 
        .ZN(n1027) );
  INV_X1 U400 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U401 ( .A1(data_in[4]), .A2(n835), .B1(n1030), .B2(\mem[19][4] ), 
        .ZN(n1026) );
  INV_X1 U402 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U403 ( .A1(data_in[5]), .A2(n835), .B1(n1030), .B2(\mem[19][5] ), 
        .ZN(n1025) );
  INV_X1 U404 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U405 ( .A1(data_in[6]), .A2(n835), .B1(n1030), .B2(\mem[19][6] ), 
        .ZN(n1024) );
  INV_X1 U406 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U407 ( .A1(data_in[7]), .A2(n835), .B1(n1030), .B2(\mem[19][7] ), 
        .ZN(n1023) );
  INV_X1 U408 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U409 ( .A1(data_in[0]), .A2(n834), .B1(n1021), .B2(\mem[20][0] ), 
        .ZN(n1022) );
  INV_X1 U410 ( .A(n1020), .ZN(n725) );
  AOI22_X1 U411 ( .A1(data_in[1]), .A2(n834), .B1(n1021), .B2(\mem[20][1] ), 
        .ZN(n1020) );
  INV_X1 U412 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U413 ( .A1(data_in[2]), .A2(n834), .B1(n1021), .B2(\mem[20][2] ), 
        .ZN(n1019) );
  INV_X1 U414 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U415 ( .A1(data_in[3]), .A2(n834), .B1(n1021), .B2(\mem[20][3] ), 
        .ZN(n1018) );
  INV_X1 U416 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U417 ( .A1(data_in[4]), .A2(n834), .B1(n1021), .B2(\mem[20][4] ), 
        .ZN(n1017) );
  INV_X1 U418 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U419 ( .A1(data_in[5]), .A2(n834), .B1(n1021), .B2(\mem[20][5] ), 
        .ZN(n1016) );
  INV_X1 U420 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U421 ( .A1(data_in[6]), .A2(n834), .B1(n1021), .B2(\mem[20][6] ), 
        .ZN(n1015) );
  INV_X1 U422 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U423 ( .A1(data_in[7]), .A2(n834), .B1(n1021), .B2(\mem[20][7] ), 
        .ZN(n1014) );
  INV_X1 U424 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U425 ( .A1(data_in[0]), .A2(n833), .B1(n1012), .B2(\mem[21][0] ), 
        .ZN(n1013) );
  INV_X1 U426 ( .A(n1011), .ZN(n717) );
  AOI22_X1 U427 ( .A1(data_in[1]), .A2(n833), .B1(n1012), .B2(\mem[21][1] ), 
        .ZN(n1011) );
  INV_X1 U428 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U429 ( .A1(data_in[2]), .A2(n833), .B1(n1012), .B2(\mem[21][2] ), 
        .ZN(n1010) );
  INV_X1 U430 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U431 ( .A1(data_in[3]), .A2(n833), .B1(n1012), .B2(\mem[21][3] ), 
        .ZN(n1009) );
  INV_X1 U432 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U433 ( .A1(data_in[4]), .A2(n833), .B1(n1012), .B2(\mem[21][4] ), 
        .ZN(n1008) );
  INV_X1 U434 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U435 ( .A1(data_in[5]), .A2(n833), .B1(n1012), .B2(\mem[21][5] ), 
        .ZN(n1007) );
  INV_X1 U436 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U437 ( .A1(data_in[6]), .A2(n833), .B1(n1012), .B2(\mem[21][6] ), 
        .ZN(n1006) );
  INV_X1 U438 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U439 ( .A1(data_in[7]), .A2(n833), .B1(n1012), .B2(\mem[21][7] ), 
        .ZN(n1005) );
  INV_X1 U440 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U441 ( .A1(data_in[0]), .A2(n832), .B1(n1003), .B2(\mem[22][0] ), 
        .ZN(n1004) );
  INV_X1 U442 ( .A(n1002), .ZN(n709) );
  AOI22_X1 U443 ( .A1(data_in[1]), .A2(n832), .B1(n1003), .B2(\mem[22][1] ), 
        .ZN(n1002) );
  INV_X1 U444 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U445 ( .A1(data_in[2]), .A2(n832), .B1(n1003), .B2(\mem[22][2] ), 
        .ZN(n1001) );
  INV_X1 U446 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U447 ( .A1(data_in[3]), .A2(n832), .B1(n1003), .B2(\mem[22][3] ), 
        .ZN(n1000) );
  INV_X1 U448 ( .A(n999), .ZN(n706) );
  AOI22_X1 U449 ( .A1(data_in[4]), .A2(n832), .B1(n1003), .B2(\mem[22][4] ), 
        .ZN(n999) );
  INV_X1 U450 ( .A(n998), .ZN(n705) );
  AOI22_X1 U451 ( .A1(data_in[5]), .A2(n832), .B1(n1003), .B2(\mem[22][5] ), 
        .ZN(n998) );
  INV_X1 U452 ( .A(n997), .ZN(n704) );
  AOI22_X1 U453 ( .A1(data_in[6]), .A2(n832), .B1(n1003), .B2(\mem[22][6] ), 
        .ZN(n997) );
  INV_X1 U454 ( .A(n996), .ZN(n703) );
  AOI22_X1 U455 ( .A1(data_in[7]), .A2(n832), .B1(n1003), .B2(\mem[22][7] ), 
        .ZN(n996) );
  INV_X1 U456 ( .A(n995), .ZN(n702) );
  AOI22_X1 U457 ( .A1(data_in[0]), .A2(n831), .B1(n994), .B2(\mem[23][0] ), 
        .ZN(n995) );
  INV_X1 U458 ( .A(n993), .ZN(n701) );
  AOI22_X1 U459 ( .A1(data_in[1]), .A2(n831), .B1(n994), .B2(\mem[23][1] ), 
        .ZN(n993) );
  INV_X1 U460 ( .A(n992), .ZN(n700) );
  AOI22_X1 U461 ( .A1(data_in[2]), .A2(n831), .B1(n994), .B2(\mem[23][2] ), 
        .ZN(n992) );
  INV_X1 U462 ( .A(n991), .ZN(n699) );
  AOI22_X1 U463 ( .A1(data_in[3]), .A2(n831), .B1(n994), .B2(\mem[23][3] ), 
        .ZN(n991) );
  INV_X1 U464 ( .A(n990), .ZN(n698) );
  AOI22_X1 U465 ( .A1(data_in[4]), .A2(n831), .B1(n994), .B2(\mem[23][4] ), 
        .ZN(n990) );
  INV_X1 U466 ( .A(n989), .ZN(n697) );
  AOI22_X1 U467 ( .A1(data_in[5]), .A2(n831), .B1(n994), .B2(\mem[23][5] ), 
        .ZN(n989) );
  INV_X1 U468 ( .A(n988), .ZN(n696) );
  AOI22_X1 U469 ( .A1(data_in[6]), .A2(n831), .B1(n994), .B2(\mem[23][6] ), 
        .ZN(n988) );
  INV_X1 U470 ( .A(n987), .ZN(n695) );
  AOI22_X1 U471 ( .A1(data_in[7]), .A2(n831), .B1(n994), .B2(\mem[23][7] ), 
        .ZN(n987) );
  INV_X1 U472 ( .A(n986), .ZN(n694) );
  AOI22_X1 U473 ( .A1(data_in[0]), .A2(n830), .B1(n985), .B2(\mem[24][0] ), 
        .ZN(n986) );
  INV_X1 U474 ( .A(n984), .ZN(n693) );
  AOI22_X1 U475 ( .A1(data_in[1]), .A2(n830), .B1(n985), .B2(\mem[24][1] ), 
        .ZN(n984) );
  INV_X1 U476 ( .A(n983), .ZN(n692) );
  AOI22_X1 U477 ( .A1(data_in[2]), .A2(n830), .B1(n985), .B2(\mem[24][2] ), 
        .ZN(n983) );
  INV_X1 U478 ( .A(n982), .ZN(n691) );
  AOI22_X1 U479 ( .A1(data_in[3]), .A2(n830), .B1(n985), .B2(\mem[24][3] ), 
        .ZN(n982) );
  INV_X1 U480 ( .A(n981), .ZN(n690) );
  AOI22_X1 U481 ( .A1(data_in[4]), .A2(n830), .B1(n985), .B2(\mem[24][4] ), 
        .ZN(n981) );
  INV_X1 U482 ( .A(n980), .ZN(n689) );
  AOI22_X1 U483 ( .A1(data_in[5]), .A2(n830), .B1(n985), .B2(\mem[24][5] ), 
        .ZN(n980) );
  INV_X1 U484 ( .A(n979), .ZN(n688) );
  AOI22_X1 U485 ( .A1(data_in[6]), .A2(n830), .B1(n985), .B2(\mem[24][6] ), 
        .ZN(n979) );
  INV_X1 U486 ( .A(n978), .ZN(n687) );
  AOI22_X1 U487 ( .A1(data_in[7]), .A2(n830), .B1(n985), .B2(\mem[24][7] ), 
        .ZN(n978) );
  INV_X1 U488 ( .A(n976), .ZN(n686) );
  AOI22_X1 U489 ( .A1(data_in[0]), .A2(n829), .B1(n975), .B2(\mem[25][0] ), 
        .ZN(n976) );
  INV_X1 U490 ( .A(n974), .ZN(n685) );
  AOI22_X1 U491 ( .A1(data_in[1]), .A2(n829), .B1(n975), .B2(\mem[25][1] ), 
        .ZN(n974) );
  INV_X1 U492 ( .A(n973), .ZN(n684) );
  AOI22_X1 U493 ( .A1(data_in[2]), .A2(n829), .B1(n975), .B2(\mem[25][2] ), 
        .ZN(n973) );
  INV_X1 U494 ( .A(n972), .ZN(n683) );
  AOI22_X1 U495 ( .A1(data_in[3]), .A2(n829), .B1(n975), .B2(\mem[25][3] ), 
        .ZN(n972) );
  INV_X1 U496 ( .A(n971), .ZN(n682) );
  AOI22_X1 U497 ( .A1(data_in[4]), .A2(n829), .B1(n975), .B2(\mem[25][4] ), 
        .ZN(n971) );
  INV_X1 U498 ( .A(n970), .ZN(n681) );
  AOI22_X1 U499 ( .A1(data_in[5]), .A2(n829), .B1(n975), .B2(\mem[25][5] ), 
        .ZN(n970) );
  INV_X1 U500 ( .A(n969), .ZN(n680) );
  AOI22_X1 U501 ( .A1(data_in[6]), .A2(n829), .B1(n975), .B2(\mem[25][6] ), 
        .ZN(n969) );
  INV_X1 U502 ( .A(n968), .ZN(n679) );
  AOI22_X1 U503 ( .A1(data_in[7]), .A2(n829), .B1(n975), .B2(\mem[25][7] ), 
        .ZN(n968) );
  INV_X1 U504 ( .A(n967), .ZN(n678) );
  AOI22_X1 U505 ( .A1(data_in[0]), .A2(n828), .B1(n966), .B2(\mem[26][0] ), 
        .ZN(n967) );
  INV_X1 U506 ( .A(n965), .ZN(n677) );
  AOI22_X1 U507 ( .A1(data_in[1]), .A2(n828), .B1(n966), .B2(\mem[26][1] ), 
        .ZN(n965) );
  INV_X1 U508 ( .A(n964), .ZN(n676) );
  AOI22_X1 U509 ( .A1(data_in[2]), .A2(n828), .B1(n966), .B2(\mem[26][2] ), 
        .ZN(n964) );
  INV_X1 U510 ( .A(n963), .ZN(n675) );
  AOI22_X1 U511 ( .A1(data_in[3]), .A2(n828), .B1(n966), .B2(\mem[26][3] ), 
        .ZN(n963) );
  INV_X1 U512 ( .A(n962), .ZN(n674) );
  AOI22_X1 U513 ( .A1(data_in[4]), .A2(n828), .B1(n966), .B2(\mem[26][4] ), 
        .ZN(n962) );
  INV_X1 U514 ( .A(n961), .ZN(n673) );
  AOI22_X1 U515 ( .A1(data_in[5]), .A2(n828), .B1(n966), .B2(\mem[26][5] ), 
        .ZN(n961) );
  INV_X1 U516 ( .A(n960), .ZN(n672) );
  AOI22_X1 U517 ( .A1(data_in[6]), .A2(n828), .B1(n966), .B2(\mem[26][6] ), 
        .ZN(n960) );
  INV_X1 U518 ( .A(n959), .ZN(n671) );
  AOI22_X1 U519 ( .A1(data_in[7]), .A2(n828), .B1(n966), .B2(\mem[26][7] ), 
        .ZN(n959) );
  INV_X1 U520 ( .A(n958), .ZN(n670) );
  AOI22_X1 U521 ( .A1(data_in[0]), .A2(n827), .B1(n957), .B2(\mem[27][0] ), 
        .ZN(n958) );
  INV_X1 U522 ( .A(n956), .ZN(n669) );
  AOI22_X1 U523 ( .A1(data_in[1]), .A2(n827), .B1(n957), .B2(\mem[27][1] ), 
        .ZN(n956) );
  INV_X1 U524 ( .A(n955), .ZN(n668) );
  AOI22_X1 U525 ( .A1(data_in[2]), .A2(n827), .B1(n957), .B2(\mem[27][2] ), 
        .ZN(n955) );
  INV_X1 U526 ( .A(n954), .ZN(n667) );
  AOI22_X1 U527 ( .A1(data_in[3]), .A2(n827), .B1(n957), .B2(\mem[27][3] ), 
        .ZN(n954) );
  INV_X1 U528 ( .A(n953), .ZN(n666) );
  AOI22_X1 U529 ( .A1(data_in[4]), .A2(n827), .B1(n957), .B2(\mem[27][4] ), 
        .ZN(n953) );
  INV_X1 U530 ( .A(n952), .ZN(n665) );
  AOI22_X1 U531 ( .A1(data_in[5]), .A2(n827), .B1(n957), .B2(\mem[27][5] ), 
        .ZN(n952) );
  INV_X1 U532 ( .A(n951), .ZN(n664) );
  AOI22_X1 U533 ( .A1(data_in[6]), .A2(n827), .B1(n957), .B2(\mem[27][6] ), 
        .ZN(n951) );
  INV_X1 U534 ( .A(n950), .ZN(n663) );
  AOI22_X1 U535 ( .A1(data_in[7]), .A2(n827), .B1(n957), .B2(\mem[27][7] ), 
        .ZN(n950) );
  INV_X1 U536 ( .A(n949), .ZN(n662) );
  AOI22_X1 U537 ( .A1(data_in[0]), .A2(n826), .B1(n948), .B2(\mem[28][0] ), 
        .ZN(n949) );
  INV_X1 U538 ( .A(n947), .ZN(n661) );
  AOI22_X1 U539 ( .A1(data_in[1]), .A2(n826), .B1(n948), .B2(\mem[28][1] ), 
        .ZN(n947) );
  INV_X1 U540 ( .A(n946), .ZN(n660) );
  AOI22_X1 U541 ( .A1(data_in[2]), .A2(n826), .B1(n948), .B2(\mem[28][2] ), 
        .ZN(n946) );
  INV_X1 U542 ( .A(n945), .ZN(n659) );
  AOI22_X1 U543 ( .A1(data_in[3]), .A2(n826), .B1(n948), .B2(\mem[28][3] ), 
        .ZN(n945) );
  INV_X1 U544 ( .A(n944), .ZN(n658) );
  AOI22_X1 U545 ( .A1(data_in[4]), .A2(n826), .B1(n948), .B2(\mem[28][4] ), 
        .ZN(n944) );
  INV_X1 U546 ( .A(n943), .ZN(n657) );
  AOI22_X1 U547 ( .A1(data_in[5]), .A2(n826), .B1(n948), .B2(\mem[28][5] ), 
        .ZN(n943) );
  INV_X1 U548 ( .A(n942), .ZN(n656) );
  AOI22_X1 U549 ( .A1(data_in[6]), .A2(n826), .B1(n948), .B2(\mem[28][6] ), 
        .ZN(n942) );
  INV_X1 U550 ( .A(n941), .ZN(n655) );
  AOI22_X1 U551 ( .A1(data_in[7]), .A2(n826), .B1(n948), .B2(\mem[28][7] ), 
        .ZN(n941) );
  INV_X1 U552 ( .A(n940), .ZN(n654) );
  AOI22_X1 U553 ( .A1(data_in[0]), .A2(n825), .B1(n939), .B2(\mem[29][0] ), 
        .ZN(n940) );
  INV_X1 U554 ( .A(n938), .ZN(n653) );
  AOI22_X1 U555 ( .A1(data_in[1]), .A2(n825), .B1(n939), .B2(\mem[29][1] ), 
        .ZN(n938) );
  INV_X1 U556 ( .A(n937), .ZN(n652) );
  AOI22_X1 U557 ( .A1(data_in[2]), .A2(n825), .B1(n939), .B2(\mem[29][2] ), 
        .ZN(n937) );
  INV_X1 U558 ( .A(n936), .ZN(n651) );
  AOI22_X1 U559 ( .A1(data_in[3]), .A2(n825), .B1(n939), .B2(\mem[29][3] ), 
        .ZN(n936) );
  INV_X1 U560 ( .A(n935), .ZN(n650) );
  AOI22_X1 U561 ( .A1(data_in[4]), .A2(n825), .B1(n939), .B2(\mem[29][4] ), 
        .ZN(n935) );
  INV_X1 U562 ( .A(n934), .ZN(n649) );
  AOI22_X1 U563 ( .A1(data_in[5]), .A2(n825), .B1(n939), .B2(\mem[29][5] ), 
        .ZN(n934) );
  INV_X1 U564 ( .A(n933), .ZN(n648) );
  AOI22_X1 U565 ( .A1(data_in[6]), .A2(n825), .B1(n939), .B2(\mem[29][6] ), 
        .ZN(n933) );
  INV_X1 U566 ( .A(n932), .ZN(n647) );
  AOI22_X1 U567 ( .A1(data_in[7]), .A2(n825), .B1(n939), .B2(\mem[29][7] ), 
        .ZN(n932) );
  INV_X1 U568 ( .A(n931), .ZN(n646) );
  AOI22_X1 U569 ( .A1(data_in[0]), .A2(n824), .B1(n930), .B2(\mem[30][0] ), 
        .ZN(n931) );
  INV_X1 U570 ( .A(n929), .ZN(n645) );
  AOI22_X1 U571 ( .A1(data_in[1]), .A2(n824), .B1(n930), .B2(\mem[30][1] ), 
        .ZN(n929) );
  INV_X1 U572 ( .A(n928), .ZN(n644) );
  AOI22_X1 U573 ( .A1(data_in[2]), .A2(n824), .B1(n930), .B2(\mem[30][2] ), 
        .ZN(n928) );
  INV_X1 U574 ( .A(n927), .ZN(n643) );
  AOI22_X1 U575 ( .A1(data_in[3]), .A2(n824), .B1(n930), .B2(\mem[30][3] ), 
        .ZN(n927) );
  INV_X1 U576 ( .A(n926), .ZN(n642) );
  AOI22_X1 U577 ( .A1(data_in[4]), .A2(n824), .B1(n930), .B2(\mem[30][4] ), 
        .ZN(n926) );
  INV_X1 U578 ( .A(n925), .ZN(n641) );
  AOI22_X1 U579 ( .A1(data_in[5]), .A2(n824), .B1(n930), .B2(\mem[30][5] ), 
        .ZN(n925) );
  INV_X1 U580 ( .A(n924), .ZN(n640) );
  AOI22_X1 U581 ( .A1(data_in[6]), .A2(n824), .B1(n930), .B2(\mem[30][6] ), 
        .ZN(n924) );
  INV_X1 U582 ( .A(n923), .ZN(n639) );
  AOI22_X1 U583 ( .A1(data_in[7]), .A2(n824), .B1(n930), .B2(\mem[30][7] ), 
        .ZN(n923) );
  INV_X1 U584 ( .A(n922), .ZN(n638) );
  AOI22_X1 U585 ( .A1(data_in[0]), .A2(n823), .B1(n921), .B2(\mem[31][0] ), 
        .ZN(n922) );
  INV_X1 U586 ( .A(n920), .ZN(n637) );
  AOI22_X1 U587 ( .A1(data_in[1]), .A2(n823), .B1(n921), .B2(\mem[31][1] ), 
        .ZN(n920) );
  INV_X1 U588 ( .A(n919), .ZN(n636) );
  AOI22_X1 U589 ( .A1(data_in[2]), .A2(n823), .B1(n921), .B2(\mem[31][2] ), 
        .ZN(n919) );
  INV_X1 U590 ( .A(n918), .ZN(n635) );
  AOI22_X1 U591 ( .A1(data_in[3]), .A2(n823), .B1(n921), .B2(\mem[31][3] ), 
        .ZN(n918) );
  INV_X1 U592 ( .A(n917), .ZN(n634) );
  AOI22_X1 U593 ( .A1(data_in[4]), .A2(n823), .B1(n921), .B2(\mem[31][4] ), 
        .ZN(n917) );
  INV_X1 U594 ( .A(n916), .ZN(n633) );
  AOI22_X1 U595 ( .A1(data_in[5]), .A2(n823), .B1(n921), .B2(\mem[31][5] ), 
        .ZN(n916) );
  INV_X1 U596 ( .A(n915), .ZN(n632) );
  AOI22_X1 U597 ( .A1(data_in[6]), .A2(n823), .B1(n921), .B2(\mem[31][6] ), 
        .ZN(n915) );
  INV_X1 U598 ( .A(n914), .ZN(n631) );
  AOI22_X1 U599 ( .A1(data_in[7]), .A2(n823), .B1(n921), .B2(\mem[31][7] ), 
        .ZN(n914) );
  MUX2_X1 U600 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n612), .Z(n2) );
  MUX2_X1 U601 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n612), .Z(n3) );
  MUX2_X1 U602 ( .A(n3), .B(n2), .S(n609), .Z(n4) );
  MUX2_X1 U603 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n612), .Z(n5) );
  MUX2_X1 U604 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n612), .Z(n6) );
  MUX2_X1 U605 ( .A(n6), .B(n5), .S(n609), .Z(n7) );
  MUX2_X1 U606 ( .A(n7), .B(n4), .S(n608), .Z(n8) );
  MUX2_X1 U607 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n612), .Z(n9) );
  MUX2_X1 U608 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n612), .Z(n10) );
  MUX2_X1 U609 ( .A(n10), .B(n9), .S(n609), .Z(n11) );
  MUX2_X1 U610 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n612), .Z(n12) );
  MUX2_X1 U611 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n612), .Z(n13) );
  MUX2_X1 U612 ( .A(n13), .B(n12), .S(n609), .Z(n14) );
  MUX2_X1 U613 ( .A(n14), .B(n11), .S(N12), .Z(n15) );
  MUX2_X1 U614 ( .A(n15), .B(n8), .S(N13), .Z(n16) );
  MUX2_X1 U615 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n613), .Z(n17) );
  MUX2_X1 U616 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n613), .Z(n18) );
  MUX2_X1 U617 ( .A(n18), .B(n17), .S(n610), .Z(n19) );
  MUX2_X1 U618 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n613), .Z(n20) );
  MUX2_X1 U619 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n613), .Z(n21) );
  MUX2_X1 U620 ( .A(n21), .B(n20), .S(n610), .Z(n22) );
  MUX2_X1 U621 ( .A(n22), .B(n19), .S(N12), .Z(n23) );
  MUX2_X1 U622 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n613), .Z(n24) );
  MUX2_X1 U623 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n613), .Z(n25) );
  MUX2_X1 U624 ( .A(n25), .B(n24), .S(n610), .Z(n26) );
  MUX2_X1 U625 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n613), .Z(n27) );
  MUX2_X1 U626 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n613), .Z(n28) );
  MUX2_X1 U627 ( .A(n28), .B(n27), .S(n610), .Z(n29) );
  MUX2_X1 U628 ( .A(n29), .B(n26), .S(n607), .Z(n30) );
  MUX2_X1 U629 ( .A(n30), .B(n23), .S(N13), .Z(n31) );
  MUX2_X1 U630 ( .A(n31), .B(n16), .S(N14), .Z(N22) );
  MUX2_X1 U631 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n613), .Z(n32) );
  MUX2_X1 U632 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n613), .Z(n33) );
  MUX2_X1 U633 ( .A(n33), .B(n32), .S(n610), .Z(n34) );
  MUX2_X1 U634 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n613), .Z(n35) );
  MUX2_X1 U635 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n613), .Z(n36) );
  MUX2_X1 U636 ( .A(n36), .B(n35), .S(n610), .Z(n37) );
  MUX2_X1 U637 ( .A(n37), .B(n34), .S(n607), .Z(n38) );
  MUX2_X1 U638 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n614), .Z(n39) );
  MUX2_X1 U639 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n614), .Z(n40) );
  MUX2_X1 U640 ( .A(n40), .B(n39), .S(n610), .Z(n41) );
  MUX2_X1 U641 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n614), .Z(n42) );
  MUX2_X1 U642 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n614), .Z(n43) );
  MUX2_X1 U643 ( .A(n43), .B(n42), .S(n610), .Z(n44) );
  MUX2_X1 U644 ( .A(n44), .B(n41), .S(N12), .Z(n45) );
  MUX2_X1 U645 ( .A(n45), .B(n38), .S(N13), .Z(n46) );
  MUX2_X1 U646 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n614), .Z(n47) );
  MUX2_X1 U647 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n614), .Z(n48) );
  MUX2_X1 U648 ( .A(n48), .B(n47), .S(n610), .Z(n49) );
  MUX2_X1 U649 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n614), .Z(n50) );
  MUX2_X1 U650 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n614), .Z(n51) );
  MUX2_X1 U651 ( .A(n51), .B(n50), .S(n610), .Z(n52) );
  MUX2_X1 U652 ( .A(n52), .B(n49), .S(n608), .Z(n53) );
  MUX2_X1 U653 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n614), .Z(n54) );
  MUX2_X1 U654 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n614), .Z(n55) );
  MUX2_X1 U655 ( .A(n55), .B(n54), .S(n610), .Z(n56) );
  MUX2_X1 U656 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n614), .Z(n57) );
  MUX2_X1 U657 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n614), .Z(n58) );
  MUX2_X1 U658 ( .A(n58), .B(n57), .S(n610), .Z(n59) );
  MUX2_X1 U659 ( .A(n59), .B(n56), .S(n608), .Z(n60) );
  MUX2_X1 U660 ( .A(n60), .B(n53), .S(N13), .Z(n61) );
  MUX2_X1 U661 ( .A(n61), .B(n46), .S(N14), .Z(N21) );
  MUX2_X1 U662 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n614), .Z(n62) );
  MUX2_X1 U663 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n619), .Z(n63) );
  MUX2_X1 U664 ( .A(n63), .B(n62), .S(n611), .Z(n64) );
  MUX2_X1 U665 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n612), .Z(n65) );
  MUX2_X1 U666 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n620), .Z(n66) );
  MUX2_X1 U667 ( .A(n66), .B(n65), .S(n611), .Z(n67) );
  MUX2_X1 U668 ( .A(n67), .B(n64), .S(n607), .Z(n68) );
  MUX2_X1 U669 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n619), .Z(n69) );
  MUX2_X1 U670 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n619), .Z(n70) );
  MUX2_X1 U671 ( .A(n70), .B(n69), .S(n611), .Z(n71) );
  MUX2_X1 U672 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n618), .Z(n72) );
  MUX2_X1 U673 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n619), .Z(n73) );
  MUX2_X1 U674 ( .A(n73), .B(n72), .S(n611), .Z(n74) );
  MUX2_X1 U675 ( .A(n74), .B(n71), .S(n607), .Z(n75) );
  MUX2_X1 U676 ( .A(n75), .B(n68), .S(N13), .Z(n76) );
  MUX2_X1 U677 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n613), .Z(n77) );
  MUX2_X1 U678 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n619), .Z(n78) );
  MUX2_X1 U679 ( .A(n78), .B(n77), .S(n611), .Z(n79) );
  MUX2_X1 U680 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n616), .Z(n80) );
  MUX2_X1 U681 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n620), .Z(n81) );
  MUX2_X1 U682 ( .A(n81), .B(n80), .S(n611), .Z(n82) );
  MUX2_X1 U683 ( .A(n82), .B(n79), .S(n607), .Z(n83) );
  MUX2_X1 U684 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n615), .Z(n84) );
  MUX2_X1 U685 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n615), .Z(n85) );
  MUX2_X1 U686 ( .A(n85), .B(n84), .S(n611), .Z(n86) );
  MUX2_X1 U687 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n615), .Z(n87) );
  MUX2_X1 U688 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n615), .Z(n88) );
  MUX2_X1 U689 ( .A(n88), .B(n87), .S(n611), .Z(n89) );
  MUX2_X1 U690 ( .A(n89), .B(n86), .S(n607), .Z(n90) );
  MUX2_X1 U691 ( .A(n90), .B(n83), .S(N13), .Z(n91) );
  MUX2_X1 U692 ( .A(n91), .B(n76), .S(N14), .Z(N20) );
  MUX2_X1 U693 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n615), .Z(n92) );
  MUX2_X1 U694 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n615), .Z(n93) );
  MUX2_X1 U695 ( .A(n93), .B(n92), .S(n611), .Z(n94) );
  MUX2_X1 U696 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n615), .Z(n95) );
  MUX2_X1 U697 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n615), .Z(n96) );
  MUX2_X1 U698 ( .A(n96), .B(n95), .S(n611), .Z(n97) );
  MUX2_X1 U699 ( .A(n97), .B(n94), .S(n607), .Z(n98) );
  MUX2_X1 U700 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n615), .Z(n99) );
  MUX2_X1 U701 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n615), .Z(n100) );
  MUX2_X1 U702 ( .A(n100), .B(n99), .S(n611), .Z(n101) );
  MUX2_X1 U703 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n615), .Z(n102) );
  MUX2_X1 U704 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n615), .Z(n103) );
  MUX2_X1 U705 ( .A(n103), .B(n102), .S(n611), .Z(n104) );
  MUX2_X1 U706 ( .A(n104), .B(n101), .S(n607), .Z(n105) );
  MUX2_X1 U707 ( .A(n105), .B(n98), .S(N13), .Z(n106) );
  MUX2_X1 U708 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n616), .Z(n107) );
  MUX2_X1 U709 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n620), .Z(n108) );
  MUX2_X1 U710 ( .A(n108), .B(n107), .S(n611), .Z(n109) );
  MUX2_X1 U711 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n619), .Z(n110) );
  MUX2_X1 U712 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n111) );
  MUX2_X1 U713 ( .A(n111), .B(n110), .S(n610), .Z(n112) );
  MUX2_X1 U714 ( .A(n112), .B(n109), .S(n607), .Z(n113) );
  MUX2_X1 U715 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n618), .Z(n114) );
  MUX2_X1 U716 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n620), .Z(n115) );
  MUX2_X1 U717 ( .A(n115), .B(n114), .S(n609), .Z(n116) );
  MUX2_X1 U718 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n619), .Z(n117) );
  MUX2_X1 U719 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n619), .Z(n118) );
  MUX2_X1 U720 ( .A(n118), .B(n117), .S(n611), .Z(n119) );
  MUX2_X1 U721 ( .A(n119), .B(n116), .S(n607), .Z(n120) );
  MUX2_X1 U722 ( .A(n120), .B(n113), .S(N13), .Z(n121) );
  MUX2_X1 U723 ( .A(n121), .B(n106), .S(N14), .Z(N19) );
  MUX2_X1 U724 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n620), .Z(n122) );
  MUX2_X1 U725 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n619), .Z(n123) );
  MUX2_X1 U726 ( .A(n123), .B(n122), .S(n609), .Z(n124) );
  MUX2_X1 U727 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(N10), .Z(n125) );
  MUX2_X1 U728 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n620), .Z(n126) );
  MUX2_X1 U729 ( .A(n126), .B(n125), .S(n609), .Z(n127) );
  MUX2_X1 U730 ( .A(n127), .B(n124), .S(n607), .Z(n128) );
  MUX2_X1 U731 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n617), .Z(n129) );
  MUX2_X1 U732 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(N10), .Z(n130) );
  MUX2_X1 U733 ( .A(n130), .B(n129), .S(n611), .Z(n131) );
  MUX2_X1 U734 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n619), .Z(n132) );
  MUX2_X1 U735 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(N10), .Z(n133) );
  MUX2_X1 U736 ( .A(n133), .B(n132), .S(n610), .Z(n134) );
  MUX2_X1 U737 ( .A(n134), .B(n131), .S(n607), .Z(n135) );
  MUX2_X1 U738 ( .A(n135), .B(n128), .S(N13), .Z(n136) );
  MUX2_X1 U739 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n619), .Z(n137) );
  MUX2_X1 U740 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n620), .Z(n138) );
  MUX2_X1 U741 ( .A(n138), .B(n137), .S(n610), .Z(n139) );
  MUX2_X1 U742 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n612), .Z(n140) );
  MUX2_X1 U743 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n612), .Z(n141) );
  MUX2_X1 U744 ( .A(n141), .B(n140), .S(n609), .Z(n142) );
  MUX2_X1 U745 ( .A(n142), .B(n139), .S(n607), .Z(n143) );
  MUX2_X1 U746 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n620), .Z(n144) );
  MUX2_X1 U747 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n145) );
  MUX2_X1 U748 ( .A(n145), .B(n144), .S(n610), .Z(n146) );
  MUX2_X1 U749 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n612), .Z(n147) );
  MUX2_X1 U750 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n612), .Z(n148) );
  MUX2_X1 U751 ( .A(n148), .B(n147), .S(n609), .Z(n149) );
  MUX2_X1 U752 ( .A(n149), .B(n146), .S(n607), .Z(n150) );
  MUX2_X1 U753 ( .A(n150), .B(n143), .S(N13), .Z(n151) );
  MUX2_X1 U754 ( .A(n151), .B(n136), .S(N14), .Z(N18) );
  MUX2_X1 U755 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n616), .Z(n152) );
  MUX2_X1 U756 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n616), .Z(n153) );
  MUX2_X1 U757 ( .A(n153), .B(n152), .S(n610), .Z(n154) );
  MUX2_X1 U758 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n616), .Z(n155) );
  MUX2_X1 U759 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n616), .Z(n156) );
  MUX2_X1 U760 ( .A(n156), .B(n155), .S(N11), .Z(n157) );
  MUX2_X1 U761 ( .A(n157), .B(n154), .S(n608), .Z(n158) );
  MUX2_X1 U762 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n616), .Z(n159) );
  MUX2_X1 U763 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n616), .Z(n160) );
  MUX2_X1 U764 ( .A(n160), .B(n159), .S(n609), .Z(n161) );
  MUX2_X1 U765 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n616), .Z(n162) );
  MUX2_X1 U766 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n616), .Z(n163) );
  MUX2_X1 U767 ( .A(n163), .B(n162), .S(N11), .Z(n164) );
  MUX2_X1 U768 ( .A(n164), .B(n161), .S(n608), .Z(n165) );
  MUX2_X1 U769 ( .A(n165), .B(n158), .S(N13), .Z(n166) );
  MUX2_X1 U770 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n616), .Z(n167) );
  MUX2_X1 U771 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n616), .Z(n168) );
  MUX2_X1 U772 ( .A(n168), .B(n167), .S(n611), .Z(n169) );
  MUX2_X1 U773 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n616), .Z(n170) );
  MUX2_X1 U774 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n616), .Z(n171) );
  MUX2_X1 U775 ( .A(n171), .B(n170), .S(n611), .Z(n172) );
  MUX2_X1 U776 ( .A(n172), .B(n169), .S(n608), .Z(n173) );
  MUX2_X1 U777 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n617), .Z(n174) );
  MUX2_X1 U778 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n617), .Z(n175) );
  MUX2_X1 U779 ( .A(n175), .B(n174), .S(n611), .Z(n176) );
  MUX2_X1 U780 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n617), .Z(n177) );
  MUX2_X1 U781 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n617), .Z(n178) );
  MUX2_X1 U782 ( .A(n178), .B(n177), .S(n610), .Z(n179) );
  MUX2_X1 U783 ( .A(n179), .B(n176), .S(n608), .Z(n180) );
  MUX2_X1 U784 ( .A(n180), .B(n173), .S(N13), .Z(n181) );
  MUX2_X1 U785 ( .A(n181), .B(n166), .S(N14), .Z(N17) );
  MUX2_X1 U786 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n617), .Z(n182) );
  MUX2_X1 U787 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n617), .Z(n183) );
  MUX2_X1 U788 ( .A(n183), .B(n182), .S(N11), .Z(n184) );
  MUX2_X1 U789 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n617), .Z(n185) );
  MUX2_X1 U790 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n617), .Z(n186) );
  MUX2_X1 U791 ( .A(n186), .B(n185), .S(n610), .Z(n187) );
  MUX2_X1 U792 ( .A(n187), .B(n184), .S(n608), .Z(n188) );
  MUX2_X1 U793 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n617), .Z(n189) );
  MUX2_X1 U794 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n617), .Z(n190) );
  MUX2_X1 U795 ( .A(n190), .B(n189), .S(N11), .Z(n191) );
  MUX2_X1 U796 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n617), .Z(n192) );
  MUX2_X1 U797 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n617), .Z(n193) );
  MUX2_X1 U798 ( .A(n193), .B(n192), .S(n610), .Z(n194) );
  MUX2_X1 U799 ( .A(n194), .B(n191), .S(n608), .Z(n195) );
  MUX2_X1 U800 ( .A(n195), .B(n188), .S(N13), .Z(n196) );
  MUX2_X1 U801 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n618), .Z(n197) );
  MUX2_X1 U802 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n618), .Z(n198) );
  MUX2_X1 U803 ( .A(n198), .B(n197), .S(n609), .Z(n199) );
  MUX2_X1 U804 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n618), .Z(n200) );
  MUX2_X1 U805 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n618), .Z(n201) );
  MUX2_X1 U806 ( .A(n201), .B(n200), .S(n610), .Z(n202) );
  MUX2_X1 U807 ( .A(n202), .B(n199), .S(n608), .Z(n203) );
  MUX2_X1 U808 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n618), .Z(n204) );
  MUX2_X1 U809 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n618), .Z(n205) );
  MUX2_X1 U810 ( .A(n205), .B(n204), .S(n609), .Z(n206) );
  MUX2_X1 U811 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n618), .Z(n207) );
  MUX2_X1 U812 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n618), .Z(n208) );
  MUX2_X1 U813 ( .A(n208), .B(n207), .S(n611), .Z(n209) );
  MUX2_X1 U814 ( .A(n209), .B(n206), .S(n608), .Z(n210) );
  MUX2_X1 U815 ( .A(n210), .B(n203), .S(N13), .Z(n211) );
  MUX2_X1 U816 ( .A(n211), .B(n196), .S(N14), .Z(N16) );
  MUX2_X1 U817 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n618), .Z(n212) );
  MUX2_X1 U818 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n618), .Z(n213) );
  MUX2_X1 U819 ( .A(n213), .B(n212), .S(n609), .Z(n214) );
  MUX2_X1 U820 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n618), .Z(n215) );
  MUX2_X1 U821 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n618), .Z(n216) );
  MUX2_X1 U822 ( .A(n216), .B(n215), .S(n609), .Z(n217) );
  MUX2_X1 U823 ( .A(n217), .B(n214), .S(n608), .Z(n218) );
  MUX2_X1 U824 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n620), .Z(n219) );
  MUX2_X1 U825 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n617), .Z(n220) );
  MUX2_X1 U826 ( .A(n220), .B(n219), .S(n609), .Z(n221) );
  MUX2_X1 U827 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n619), .Z(n222) );
  MUX2_X1 U828 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n619), .Z(n223) );
  MUX2_X1 U829 ( .A(n223), .B(n222), .S(n611), .Z(n224) );
  MUX2_X1 U830 ( .A(n224), .B(n221), .S(n608), .Z(n225) );
  MUX2_X1 U831 ( .A(n225), .B(n218), .S(N13), .Z(n226) );
  MUX2_X1 U832 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n619), .Z(n227) );
  MUX2_X1 U833 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n619), .Z(n228) );
  MUX2_X1 U834 ( .A(n228), .B(n227), .S(n609), .Z(n229) );
  MUX2_X1 U835 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n620), .Z(n595) );
  MUX2_X1 U836 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n620), .Z(n596) );
  MUX2_X1 U837 ( .A(n596), .B(n595), .S(N11), .Z(n597) );
  MUX2_X1 U838 ( .A(n597), .B(n229), .S(n608), .Z(n598) );
  MUX2_X1 U839 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n620), .Z(n599) );
  MUX2_X1 U840 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n619), .Z(n600) );
  MUX2_X1 U841 ( .A(n600), .B(n599), .S(n609), .Z(n601) );
  MUX2_X1 U842 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n620), .Z(n602) );
  MUX2_X1 U843 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n620), .Z(n603) );
  MUX2_X1 U844 ( .A(n603), .B(n602), .S(n609), .Z(n604) );
  MUX2_X1 U845 ( .A(n604), .B(n601), .S(n608), .Z(n605) );
  MUX2_X1 U846 ( .A(n605), .B(n598), .S(N13), .Z(n606) );
  MUX2_X1 U847 ( .A(n606), .B(n226), .S(N14), .Z(N15) );
  CLKBUF_X1 U848 ( .A(N11), .Z(n609) );
  INV_X1 U849 ( .A(N10), .ZN(n621) );
  INV_X1 U850 ( .A(N11), .ZN(n622) );
  INV_X1 U851 ( .A(data_in[0]), .ZN(n623) );
  INV_X1 U852 ( .A(data_in[1]), .ZN(n624) );
  INV_X1 U853 ( .A(data_in[2]), .ZN(n625) );
  INV_X1 U854 ( .A(data_in[3]), .ZN(n626) );
  INV_X1 U855 ( .A(data_in[4]), .ZN(n627) );
  INV_X1 U856 ( .A(data_in[5]), .ZN(n628) );
  INV_X1 U857 ( .A(data_in[6]), .ZN(n629) );
  INV_X1 U858 ( .A(data_in[7]), .ZN(n630) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_7 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n632), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n633), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n634), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n635), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n636), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n637), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n638), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n639), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n640), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n641), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n642), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n643), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n644), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n645), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n646), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n647), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n648), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n649), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n650), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n651), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n652), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n653), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n654), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n655), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n656), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n657), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n658), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n659), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n660), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n661), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n662), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n663), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n664), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n665), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n666), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n667), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n668), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n669), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n670), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n671), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n672), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n673), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n674), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n675), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n676), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n677), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n678), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n679), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n680), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n681), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n682), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n683), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n684), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n685), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n686), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n687), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n688), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n689), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n690), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n691), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n692), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n693), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n694), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n695), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n696), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n697), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n698), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n699), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n700), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n701), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n702), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n703), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n704), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n705), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n706), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n707), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n708), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n709), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n710), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n711), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n712), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n713), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n714), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n715), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n716), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n717), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n718), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n719), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n720), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n721), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n722), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n723), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n724), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n725), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n726), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n727), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n728), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n729), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n730), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n731), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n732), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n733), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n734), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n735), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n736), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n737), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n738), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n739), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n740), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n741), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n742), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n743), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n744), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n745), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n746), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n747), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n748), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n749), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n750), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n751), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n752), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n753), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n754), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n755), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n756), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n757), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n758), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n759), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n760), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n761), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n762), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n763), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n764), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n765), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n766), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n767), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n768), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n769), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n770), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n771), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n772), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n773), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n774), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n775), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n776), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n777), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n778), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n779), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n780), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n781), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n782), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n783), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n784), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n785), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n786), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n787), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n788), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n789), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n790), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n791), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n792), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n793), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n794), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n795), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n796), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n797), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n798), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n799), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n800), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n801), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n802), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n803), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n804), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n805), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n806), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n807), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n808), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n809), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n810), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n811), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n812), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n813), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n814), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n815), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n816), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n817), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n818), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n819), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n820), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n821), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n822), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n823), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n851), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n852), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n853), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n854), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n855), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n856), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n857), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n858), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n859), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n860), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n861), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n862), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n863), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n864), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n865), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n866), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n867), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n868), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n869), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n870), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n871), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n872), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n873), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n874), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n875), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n876), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n877), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n878), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n879), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n880), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n881), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n882), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n883), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n884), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n885), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n886), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n887), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n888), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n889), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n890), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n891), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n892), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n893), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n894), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n895), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n896), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n897), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n898), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n899), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n900), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n901), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n902), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n903), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n904), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n905), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n906), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n907), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n908), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n909), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n910), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n911), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n912), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n913), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n914), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n2) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  BUF_X1 U3 ( .A(n621), .Z(n614) );
  INV_X2 U4 ( .A(n2), .ZN(data_out[3]) );
  BUF_X1 U5 ( .A(n621), .Z(n618) );
  BUF_X1 U6 ( .A(n621), .Z(n619) );
  BUF_X1 U7 ( .A(n621), .Z(n620) );
  BUF_X1 U8 ( .A(n621), .Z(n617) );
  BUF_X1 U9 ( .A(N10), .Z(n615) );
  BUF_X1 U10 ( .A(N10), .Z(n616) );
  BUF_X1 U11 ( .A(N11), .Z(n612) );
  BUF_X1 U12 ( .A(N11), .Z(n613) );
  BUF_X1 U13 ( .A(N10), .Z(n621) );
  NOR3_X1 U14 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1206) );
  NOR3_X1 U15 ( .A1(N11), .A2(N12), .A3(n622), .ZN(n1195) );
  NOR3_X1 U16 ( .A1(N10), .A2(N12), .A3(n623), .ZN(n1185) );
  NOR3_X1 U17 ( .A1(n622), .A2(N12), .A3(n623), .ZN(n1175) );
  INV_X1 U18 ( .A(n1132), .ZN(n847) );
  INV_X1 U19 ( .A(n1122), .ZN(n846) );
  INV_X1 U20 ( .A(n1113), .ZN(n845) );
  INV_X1 U21 ( .A(n1104), .ZN(n844) );
  INV_X1 U22 ( .A(n1059), .ZN(n839) );
  INV_X1 U23 ( .A(n1049), .ZN(n838) );
  INV_X1 U24 ( .A(n1040), .ZN(n837) );
  INV_X1 U25 ( .A(n1031), .ZN(n836) );
  INV_X1 U26 ( .A(n986), .ZN(n831) );
  INV_X1 U27 ( .A(n976), .ZN(n830) );
  INV_X1 U28 ( .A(n967), .ZN(n829) );
  INV_X1 U29 ( .A(n958), .ZN(n828) );
  INV_X1 U30 ( .A(n1095), .ZN(n843) );
  INV_X1 U31 ( .A(n1086), .ZN(n842) );
  INV_X1 U32 ( .A(n1077), .ZN(n841) );
  INV_X1 U33 ( .A(n1068), .ZN(n840) );
  INV_X1 U34 ( .A(n949), .ZN(n827) );
  INV_X1 U35 ( .A(n940), .ZN(n826) );
  INV_X1 U36 ( .A(n931), .ZN(n825) );
  INV_X1 U37 ( .A(n922), .ZN(n824) );
  INV_X1 U38 ( .A(n1022), .ZN(n835) );
  INV_X1 U39 ( .A(n1013), .ZN(n834) );
  INV_X1 U40 ( .A(n1004), .ZN(n833) );
  INV_X1 U41 ( .A(n995), .ZN(n832) );
  BUF_X1 U42 ( .A(N12), .Z(n609) );
  BUF_X1 U43 ( .A(N12), .Z(n610) );
  INV_X1 U44 ( .A(N13), .ZN(n849) );
  AND3_X1 U45 ( .A1(n622), .A2(n623), .A3(N12), .ZN(n1165) );
  AND3_X1 U46 ( .A1(N10), .A2(n623), .A3(N12), .ZN(n1155) );
  AND3_X1 U47 ( .A1(N11), .A2(n622), .A3(N12), .ZN(n1145) );
  AND3_X1 U48 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1135) );
  INV_X1 U49 ( .A(N14), .ZN(n850) );
  NAND2_X1 U50 ( .A1(n1195), .A2(n1205), .ZN(n1204) );
  NAND2_X1 U51 ( .A1(n1185), .A2(n1205), .ZN(n1194) );
  NAND2_X1 U52 ( .A1(n1175), .A2(n1205), .ZN(n1184) );
  NAND2_X1 U53 ( .A1(n1165), .A2(n1205), .ZN(n1174) );
  NAND2_X1 U54 ( .A1(n1155), .A2(n1205), .ZN(n1164) );
  NAND2_X1 U55 ( .A1(n1145), .A2(n1205), .ZN(n1154) );
  NAND2_X1 U56 ( .A1(n1135), .A2(n1205), .ZN(n1144) );
  NAND2_X1 U57 ( .A1(n1206), .A2(n1205), .ZN(n1215) );
  NAND2_X1 U58 ( .A1(n1124), .A2(n1206), .ZN(n1132) );
  NAND2_X1 U59 ( .A1(n1124), .A2(n1195), .ZN(n1122) );
  NAND2_X1 U60 ( .A1(n1124), .A2(n1185), .ZN(n1113) );
  NAND2_X1 U61 ( .A1(n1124), .A2(n1175), .ZN(n1104) );
  NAND2_X1 U62 ( .A1(n1051), .A2(n1206), .ZN(n1059) );
  NAND2_X1 U63 ( .A1(n1051), .A2(n1195), .ZN(n1049) );
  NAND2_X1 U64 ( .A1(n1051), .A2(n1185), .ZN(n1040) );
  NAND2_X1 U65 ( .A1(n1051), .A2(n1175), .ZN(n1031) );
  NAND2_X1 U66 ( .A1(n978), .A2(n1206), .ZN(n986) );
  NAND2_X1 U67 ( .A1(n978), .A2(n1195), .ZN(n976) );
  NAND2_X1 U68 ( .A1(n978), .A2(n1185), .ZN(n967) );
  NAND2_X1 U69 ( .A1(n978), .A2(n1175), .ZN(n958) );
  NAND2_X1 U70 ( .A1(n1124), .A2(n1165), .ZN(n1095) );
  NAND2_X1 U71 ( .A1(n1124), .A2(n1155), .ZN(n1086) );
  NAND2_X1 U72 ( .A1(n1124), .A2(n1145), .ZN(n1077) );
  NAND2_X1 U73 ( .A1(n1124), .A2(n1135), .ZN(n1068) );
  NAND2_X1 U74 ( .A1(n1051), .A2(n1165), .ZN(n1022) );
  NAND2_X1 U75 ( .A1(n1051), .A2(n1155), .ZN(n1013) );
  NAND2_X1 U76 ( .A1(n1051), .A2(n1145), .ZN(n1004) );
  NAND2_X1 U77 ( .A1(n1051), .A2(n1135), .ZN(n995) );
  NAND2_X1 U78 ( .A1(n978), .A2(n1165), .ZN(n949) );
  NAND2_X1 U79 ( .A1(n978), .A2(n1155), .ZN(n940) );
  NAND2_X1 U80 ( .A1(n978), .A2(n1145), .ZN(n931) );
  NAND2_X1 U81 ( .A1(n978), .A2(n1135), .ZN(n922) );
  AND3_X1 U82 ( .A1(n849), .A2(n850), .A3(n1134), .ZN(n1205) );
  AND3_X1 U83 ( .A1(N13), .A2(n1134), .A3(N14), .ZN(n978) );
  AND3_X1 U84 ( .A1(n1134), .A2(n850), .A3(N13), .ZN(n1124) );
  AND3_X1 U85 ( .A1(n1134), .A2(n849), .A3(N14), .ZN(n1051) );
  NOR2_X1 U86 ( .A1(n848), .A2(addr[5]), .ZN(n1134) );
  INV_X1 U87 ( .A(wr_en), .ZN(n848) );
  OAI21_X1 U88 ( .B1(n624), .B2(n1174), .A(n1173), .ZN(n882) );
  NAND2_X1 U89 ( .A1(\mem[4][0] ), .A2(n1174), .ZN(n1173) );
  OAI21_X1 U90 ( .B1(n625), .B2(n1174), .A(n1172), .ZN(n881) );
  NAND2_X1 U91 ( .A1(\mem[4][1] ), .A2(n1174), .ZN(n1172) );
  OAI21_X1 U92 ( .B1(n626), .B2(n1174), .A(n1171), .ZN(n880) );
  NAND2_X1 U93 ( .A1(\mem[4][2] ), .A2(n1174), .ZN(n1171) );
  OAI21_X1 U94 ( .B1(n627), .B2(n1174), .A(n1170), .ZN(n879) );
  NAND2_X1 U95 ( .A1(\mem[4][3] ), .A2(n1174), .ZN(n1170) );
  OAI21_X1 U96 ( .B1(n628), .B2(n1174), .A(n1169), .ZN(n878) );
  NAND2_X1 U97 ( .A1(\mem[4][4] ), .A2(n1174), .ZN(n1169) );
  OAI21_X1 U98 ( .B1(n629), .B2(n1174), .A(n1168), .ZN(n877) );
  NAND2_X1 U99 ( .A1(\mem[4][5] ), .A2(n1174), .ZN(n1168) );
  OAI21_X1 U100 ( .B1(n630), .B2(n1174), .A(n1167), .ZN(n876) );
  NAND2_X1 U101 ( .A1(\mem[4][6] ), .A2(n1174), .ZN(n1167) );
  OAI21_X1 U102 ( .B1(n631), .B2(n1174), .A(n1166), .ZN(n875) );
  NAND2_X1 U103 ( .A1(\mem[4][7] ), .A2(n1174), .ZN(n1166) );
  OAI21_X1 U104 ( .B1(n624), .B2(n1154), .A(n1153), .ZN(n866) );
  NAND2_X1 U105 ( .A1(\mem[6][0] ), .A2(n1154), .ZN(n1153) );
  OAI21_X1 U106 ( .B1(n625), .B2(n1154), .A(n1152), .ZN(n865) );
  NAND2_X1 U107 ( .A1(\mem[6][1] ), .A2(n1154), .ZN(n1152) );
  OAI21_X1 U108 ( .B1(n626), .B2(n1154), .A(n1151), .ZN(n864) );
  NAND2_X1 U109 ( .A1(\mem[6][2] ), .A2(n1154), .ZN(n1151) );
  OAI21_X1 U110 ( .B1(n627), .B2(n1154), .A(n1150), .ZN(n863) );
  NAND2_X1 U111 ( .A1(\mem[6][3] ), .A2(n1154), .ZN(n1150) );
  OAI21_X1 U112 ( .B1(n628), .B2(n1154), .A(n1149), .ZN(n862) );
  NAND2_X1 U113 ( .A1(\mem[6][4] ), .A2(n1154), .ZN(n1149) );
  OAI21_X1 U114 ( .B1(n629), .B2(n1154), .A(n1148), .ZN(n861) );
  NAND2_X1 U115 ( .A1(\mem[6][5] ), .A2(n1154), .ZN(n1148) );
  OAI21_X1 U116 ( .B1(n630), .B2(n1154), .A(n1147), .ZN(n860) );
  NAND2_X1 U117 ( .A1(\mem[6][6] ), .A2(n1154), .ZN(n1147) );
  OAI21_X1 U118 ( .B1(n631), .B2(n1154), .A(n1146), .ZN(n859) );
  NAND2_X1 U119 ( .A1(\mem[6][7] ), .A2(n1154), .ZN(n1146) );
  OAI21_X1 U120 ( .B1(n624), .B2(n1144), .A(n1143), .ZN(n858) );
  NAND2_X1 U121 ( .A1(\mem[7][0] ), .A2(n1144), .ZN(n1143) );
  OAI21_X1 U122 ( .B1(n625), .B2(n1144), .A(n1142), .ZN(n857) );
  NAND2_X1 U123 ( .A1(\mem[7][1] ), .A2(n1144), .ZN(n1142) );
  OAI21_X1 U124 ( .B1(n626), .B2(n1144), .A(n1141), .ZN(n856) );
  NAND2_X1 U125 ( .A1(\mem[7][2] ), .A2(n1144), .ZN(n1141) );
  OAI21_X1 U126 ( .B1(n627), .B2(n1144), .A(n1140), .ZN(n855) );
  NAND2_X1 U127 ( .A1(\mem[7][3] ), .A2(n1144), .ZN(n1140) );
  OAI21_X1 U128 ( .B1(n628), .B2(n1144), .A(n1139), .ZN(n854) );
  NAND2_X1 U129 ( .A1(\mem[7][4] ), .A2(n1144), .ZN(n1139) );
  OAI21_X1 U130 ( .B1(n629), .B2(n1144), .A(n1138), .ZN(n853) );
  NAND2_X1 U131 ( .A1(\mem[7][5] ), .A2(n1144), .ZN(n1138) );
  OAI21_X1 U132 ( .B1(n630), .B2(n1144), .A(n1137), .ZN(n852) );
  NAND2_X1 U133 ( .A1(\mem[7][6] ), .A2(n1144), .ZN(n1137) );
  OAI21_X1 U134 ( .B1(n631), .B2(n1144), .A(n1136), .ZN(n851) );
  NAND2_X1 U135 ( .A1(\mem[7][7] ), .A2(n1144), .ZN(n1136) );
  OAI21_X1 U136 ( .B1(n624), .B2(n1204), .A(n1203), .ZN(n906) );
  NAND2_X1 U137 ( .A1(\mem[1][0] ), .A2(n1204), .ZN(n1203) );
  OAI21_X1 U138 ( .B1(n625), .B2(n1204), .A(n1202), .ZN(n905) );
  NAND2_X1 U139 ( .A1(\mem[1][1] ), .A2(n1204), .ZN(n1202) );
  OAI21_X1 U140 ( .B1(n626), .B2(n1204), .A(n1201), .ZN(n904) );
  NAND2_X1 U141 ( .A1(\mem[1][2] ), .A2(n1204), .ZN(n1201) );
  OAI21_X1 U142 ( .B1(n627), .B2(n1204), .A(n1200), .ZN(n903) );
  NAND2_X1 U143 ( .A1(\mem[1][3] ), .A2(n1204), .ZN(n1200) );
  OAI21_X1 U144 ( .B1(n628), .B2(n1204), .A(n1199), .ZN(n902) );
  NAND2_X1 U145 ( .A1(\mem[1][4] ), .A2(n1204), .ZN(n1199) );
  OAI21_X1 U146 ( .B1(n629), .B2(n1204), .A(n1198), .ZN(n901) );
  NAND2_X1 U147 ( .A1(\mem[1][5] ), .A2(n1204), .ZN(n1198) );
  OAI21_X1 U148 ( .B1(n630), .B2(n1204), .A(n1197), .ZN(n900) );
  NAND2_X1 U149 ( .A1(\mem[1][6] ), .A2(n1204), .ZN(n1197) );
  OAI21_X1 U150 ( .B1(n631), .B2(n1204), .A(n1196), .ZN(n899) );
  NAND2_X1 U151 ( .A1(\mem[1][7] ), .A2(n1204), .ZN(n1196) );
  OAI21_X1 U152 ( .B1(n624), .B2(n1194), .A(n1193), .ZN(n898) );
  NAND2_X1 U153 ( .A1(\mem[2][0] ), .A2(n1194), .ZN(n1193) );
  OAI21_X1 U154 ( .B1(n625), .B2(n1194), .A(n1192), .ZN(n897) );
  NAND2_X1 U155 ( .A1(\mem[2][1] ), .A2(n1194), .ZN(n1192) );
  OAI21_X1 U156 ( .B1(n626), .B2(n1194), .A(n1191), .ZN(n896) );
  NAND2_X1 U157 ( .A1(\mem[2][2] ), .A2(n1194), .ZN(n1191) );
  OAI21_X1 U158 ( .B1(n627), .B2(n1194), .A(n1190), .ZN(n895) );
  NAND2_X1 U159 ( .A1(\mem[2][3] ), .A2(n1194), .ZN(n1190) );
  OAI21_X1 U160 ( .B1(n628), .B2(n1194), .A(n1189), .ZN(n894) );
  NAND2_X1 U161 ( .A1(\mem[2][4] ), .A2(n1194), .ZN(n1189) );
  OAI21_X1 U162 ( .B1(n629), .B2(n1194), .A(n1188), .ZN(n893) );
  NAND2_X1 U163 ( .A1(\mem[2][5] ), .A2(n1194), .ZN(n1188) );
  OAI21_X1 U164 ( .B1(n630), .B2(n1194), .A(n1187), .ZN(n892) );
  NAND2_X1 U165 ( .A1(\mem[2][6] ), .A2(n1194), .ZN(n1187) );
  OAI21_X1 U166 ( .B1(n631), .B2(n1194), .A(n1186), .ZN(n891) );
  NAND2_X1 U167 ( .A1(\mem[2][7] ), .A2(n1194), .ZN(n1186) );
  OAI21_X1 U168 ( .B1(n624), .B2(n1184), .A(n1183), .ZN(n890) );
  NAND2_X1 U169 ( .A1(\mem[3][0] ), .A2(n1184), .ZN(n1183) );
  OAI21_X1 U170 ( .B1(n625), .B2(n1184), .A(n1182), .ZN(n889) );
  NAND2_X1 U171 ( .A1(\mem[3][1] ), .A2(n1184), .ZN(n1182) );
  OAI21_X1 U172 ( .B1(n626), .B2(n1184), .A(n1181), .ZN(n888) );
  NAND2_X1 U173 ( .A1(\mem[3][2] ), .A2(n1184), .ZN(n1181) );
  OAI21_X1 U174 ( .B1(n627), .B2(n1184), .A(n1180), .ZN(n887) );
  NAND2_X1 U175 ( .A1(\mem[3][3] ), .A2(n1184), .ZN(n1180) );
  OAI21_X1 U176 ( .B1(n628), .B2(n1184), .A(n1179), .ZN(n886) );
  NAND2_X1 U177 ( .A1(\mem[3][4] ), .A2(n1184), .ZN(n1179) );
  OAI21_X1 U178 ( .B1(n629), .B2(n1184), .A(n1178), .ZN(n885) );
  NAND2_X1 U179 ( .A1(\mem[3][5] ), .A2(n1184), .ZN(n1178) );
  OAI21_X1 U180 ( .B1(n630), .B2(n1184), .A(n1177), .ZN(n884) );
  NAND2_X1 U181 ( .A1(\mem[3][6] ), .A2(n1184), .ZN(n1177) );
  OAI21_X1 U182 ( .B1(n631), .B2(n1184), .A(n1176), .ZN(n883) );
  NAND2_X1 U183 ( .A1(\mem[3][7] ), .A2(n1184), .ZN(n1176) );
  OAI21_X1 U184 ( .B1(n624), .B2(n1164), .A(n1163), .ZN(n874) );
  NAND2_X1 U185 ( .A1(\mem[5][0] ), .A2(n1164), .ZN(n1163) );
  OAI21_X1 U186 ( .B1(n625), .B2(n1164), .A(n1162), .ZN(n873) );
  NAND2_X1 U187 ( .A1(\mem[5][1] ), .A2(n1164), .ZN(n1162) );
  OAI21_X1 U188 ( .B1(n626), .B2(n1164), .A(n1161), .ZN(n872) );
  NAND2_X1 U189 ( .A1(\mem[5][2] ), .A2(n1164), .ZN(n1161) );
  OAI21_X1 U190 ( .B1(n627), .B2(n1164), .A(n1160), .ZN(n871) );
  NAND2_X1 U191 ( .A1(\mem[5][3] ), .A2(n1164), .ZN(n1160) );
  OAI21_X1 U192 ( .B1(n628), .B2(n1164), .A(n1159), .ZN(n870) );
  NAND2_X1 U193 ( .A1(\mem[5][4] ), .A2(n1164), .ZN(n1159) );
  OAI21_X1 U194 ( .B1(n629), .B2(n1164), .A(n1158), .ZN(n869) );
  NAND2_X1 U195 ( .A1(\mem[5][5] ), .A2(n1164), .ZN(n1158) );
  OAI21_X1 U196 ( .B1(n630), .B2(n1164), .A(n1157), .ZN(n868) );
  NAND2_X1 U197 ( .A1(\mem[5][6] ), .A2(n1164), .ZN(n1157) );
  OAI21_X1 U198 ( .B1(n631), .B2(n1164), .A(n1156), .ZN(n867) );
  NAND2_X1 U199 ( .A1(\mem[5][7] ), .A2(n1164), .ZN(n1156) );
  OAI21_X1 U200 ( .B1(n1215), .B2(n624), .A(n1214), .ZN(n914) );
  NAND2_X1 U201 ( .A1(\mem[0][0] ), .A2(n1215), .ZN(n1214) );
  OAI21_X1 U202 ( .B1(n1215), .B2(n625), .A(n1213), .ZN(n913) );
  NAND2_X1 U203 ( .A1(\mem[0][1] ), .A2(n1215), .ZN(n1213) );
  OAI21_X1 U204 ( .B1(n1215), .B2(n626), .A(n1212), .ZN(n912) );
  NAND2_X1 U205 ( .A1(\mem[0][2] ), .A2(n1215), .ZN(n1212) );
  OAI21_X1 U206 ( .B1(n1215), .B2(n627), .A(n1211), .ZN(n911) );
  NAND2_X1 U207 ( .A1(\mem[0][3] ), .A2(n1215), .ZN(n1211) );
  OAI21_X1 U208 ( .B1(n1215), .B2(n628), .A(n1210), .ZN(n910) );
  NAND2_X1 U209 ( .A1(\mem[0][4] ), .A2(n1215), .ZN(n1210) );
  OAI21_X1 U210 ( .B1(n1215), .B2(n629), .A(n1209), .ZN(n909) );
  NAND2_X1 U211 ( .A1(\mem[0][5] ), .A2(n1215), .ZN(n1209) );
  OAI21_X1 U212 ( .B1(n1215), .B2(n630), .A(n1208), .ZN(n908) );
  NAND2_X1 U213 ( .A1(\mem[0][6] ), .A2(n1215), .ZN(n1208) );
  OAI21_X1 U214 ( .B1(n1215), .B2(n631), .A(n1207), .ZN(n907) );
  NAND2_X1 U215 ( .A1(\mem[0][7] ), .A2(n1215), .ZN(n1207) );
  INV_X1 U216 ( .A(n1133), .ZN(n823) );
  AOI22_X1 U217 ( .A1(data_in[0]), .A2(n847), .B1(n1132), .B2(\mem[8][0] ), 
        .ZN(n1133) );
  INV_X1 U218 ( .A(n1131), .ZN(n822) );
  AOI22_X1 U219 ( .A1(data_in[1]), .A2(n847), .B1(n1132), .B2(\mem[8][1] ), 
        .ZN(n1131) );
  INV_X1 U220 ( .A(n1130), .ZN(n821) );
  AOI22_X1 U221 ( .A1(data_in[2]), .A2(n847), .B1(n1132), .B2(\mem[8][2] ), 
        .ZN(n1130) );
  INV_X1 U222 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U223 ( .A1(data_in[3]), .A2(n847), .B1(n1132), .B2(\mem[8][3] ), 
        .ZN(n1129) );
  INV_X1 U224 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U225 ( .A1(data_in[4]), .A2(n847), .B1(n1132), .B2(\mem[8][4] ), 
        .ZN(n1128) );
  INV_X1 U226 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U227 ( .A1(data_in[5]), .A2(n847), .B1(n1132), .B2(\mem[8][5] ), 
        .ZN(n1127) );
  INV_X1 U228 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U229 ( .A1(data_in[6]), .A2(n847), .B1(n1132), .B2(\mem[8][6] ), 
        .ZN(n1126) );
  INV_X1 U230 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U231 ( .A1(data_in[7]), .A2(n847), .B1(n1132), .B2(\mem[8][7] ), 
        .ZN(n1125) );
  INV_X1 U232 ( .A(n1123), .ZN(n815) );
  AOI22_X1 U233 ( .A1(data_in[0]), .A2(n846), .B1(n1122), .B2(\mem[9][0] ), 
        .ZN(n1123) );
  INV_X1 U234 ( .A(n1121), .ZN(n814) );
  AOI22_X1 U235 ( .A1(data_in[1]), .A2(n846), .B1(n1122), .B2(\mem[9][1] ), 
        .ZN(n1121) );
  INV_X1 U236 ( .A(n1120), .ZN(n813) );
  AOI22_X1 U237 ( .A1(data_in[2]), .A2(n846), .B1(n1122), .B2(\mem[9][2] ), 
        .ZN(n1120) );
  INV_X1 U238 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U239 ( .A1(data_in[3]), .A2(n846), .B1(n1122), .B2(\mem[9][3] ), 
        .ZN(n1119) );
  INV_X1 U240 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U241 ( .A1(data_in[4]), .A2(n846), .B1(n1122), .B2(\mem[9][4] ), 
        .ZN(n1118) );
  INV_X1 U242 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U243 ( .A1(data_in[5]), .A2(n846), .B1(n1122), .B2(\mem[9][5] ), 
        .ZN(n1117) );
  INV_X1 U244 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U245 ( .A1(data_in[6]), .A2(n846), .B1(n1122), .B2(\mem[9][6] ), 
        .ZN(n1116) );
  INV_X1 U246 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U247 ( .A1(data_in[7]), .A2(n846), .B1(n1122), .B2(\mem[9][7] ), 
        .ZN(n1115) );
  INV_X1 U248 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U249 ( .A1(data_in[0]), .A2(n845), .B1(n1113), .B2(\mem[10][0] ), 
        .ZN(n1114) );
  INV_X1 U250 ( .A(n1112), .ZN(n806) );
  AOI22_X1 U251 ( .A1(data_in[1]), .A2(n845), .B1(n1113), .B2(\mem[10][1] ), 
        .ZN(n1112) );
  INV_X1 U252 ( .A(n1111), .ZN(n805) );
  AOI22_X1 U253 ( .A1(data_in[2]), .A2(n845), .B1(n1113), .B2(\mem[10][2] ), 
        .ZN(n1111) );
  INV_X1 U254 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U255 ( .A1(data_in[3]), .A2(n845), .B1(n1113), .B2(\mem[10][3] ), 
        .ZN(n1110) );
  INV_X1 U256 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U257 ( .A1(data_in[4]), .A2(n845), .B1(n1113), .B2(\mem[10][4] ), 
        .ZN(n1109) );
  INV_X1 U258 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U259 ( .A1(data_in[5]), .A2(n845), .B1(n1113), .B2(\mem[10][5] ), 
        .ZN(n1108) );
  INV_X1 U260 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U261 ( .A1(data_in[6]), .A2(n845), .B1(n1113), .B2(\mem[10][6] ), 
        .ZN(n1107) );
  INV_X1 U262 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U263 ( .A1(data_in[7]), .A2(n845), .B1(n1113), .B2(\mem[10][7] ), 
        .ZN(n1106) );
  INV_X1 U264 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U265 ( .A1(data_in[0]), .A2(n844), .B1(n1104), .B2(\mem[11][0] ), 
        .ZN(n1105) );
  INV_X1 U266 ( .A(n1103), .ZN(n798) );
  AOI22_X1 U267 ( .A1(data_in[1]), .A2(n844), .B1(n1104), .B2(\mem[11][1] ), 
        .ZN(n1103) );
  INV_X1 U268 ( .A(n1102), .ZN(n797) );
  AOI22_X1 U269 ( .A1(data_in[2]), .A2(n844), .B1(n1104), .B2(\mem[11][2] ), 
        .ZN(n1102) );
  INV_X1 U270 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U271 ( .A1(data_in[3]), .A2(n844), .B1(n1104), .B2(\mem[11][3] ), 
        .ZN(n1101) );
  INV_X1 U272 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U273 ( .A1(data_in[4]), .A2(n844), .B1(n1104), .B2(\mem[11][4] ), 
        .ZN(n1100) );
  INV_X1 U274 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U275 ( .A1(data_in[5]), .A2(n844), .B1(n1104), .B2(\mem[11][5] ), 
        .ZN(n1099) );
  INV_X1 U276 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U277 ( .A1(data_in[6]), .A2(n844), .B1(n1104), .B2(\mem[11][6] ), 
        .ZN(n1098) );
  INV_X1 U278 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U279 ( .A1(data_in[7]), .A2(n844), .B1(n1104), .B2(\mem[11][7] ), 
        .ZN(n1097) );
  INV_X1 U280 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U281 ( .A1(data_in[0]), .A2(n843), .B1(n1095), .B2(\mem[12][0] ), 
        .ZN(n1096) );
  INV_X1 U282 ( .A(n1094), .ZN(n790) );
  AOI22_X1 U283 ( .A1(data_in[1]), .A2(n843), .B1(n1095), .B2(\mem[12][1] ), 
        .ZN(n1094) );
  INV_X1 U284 ( .A(n1093), .ZN(n789) );
  AOI22_X1 U285 ( .A1(data_in[2]), .A2(n843), .B1(n1095), .B2(\mem[12][2] ), 
        .ZN(n1093) );
  INV_X1 U286 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U287 ( .A1(data_in[3]), .A2(n843), .B1(n1095), .B2(\mem[12][3] ), 
        .ZN(n1092) );
  INV_X1 U288 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U289 ( .A1(data_in[4]), .A2(n843), .B1(n1095), .B2(\mem[12][4] ), 
        .ZN(n1091) );
  INV_X1 U290 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U291 ( .A1(data_in[5]), .A2(n843), .B1(n1095), .B2(\mem[12][5] ), 
        .ZN(n1090) );
  INV_X1 U292 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U293 ( .A1(data_in[6]), .A2(n843), .B1(n1095), .B2(\mem[12][6] ), 
        .ZN(n1089) );
  INV_X1 U294 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U295 ( .A1(data_in[7]), .A2(n843), .B1(n1095), .B2(\mem[12][7] ), 
        .ZN(n1088) );
  INV_X1 U296 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U297 ( .A1(data_in[0]), .A2(n842), .B1(n1086), .B2(\mem[13][0] ), 
        .ZN(n1087) );
  INV_X1 U298 ( .A(n1085), .ZN(n782) );
  AOI22_X1 U299 ( .A1(data_in[1]), .A2(n842), .B1(n1086), .B2(\mem[13][1] ), 
        .ZN(n1085) );
  INV_X1 U300 ( .A(n1084), .ZN(n781) );
  AOI22_X1 U301 ( .A1(data_in[2]), .A2(n842), .B1(n1086), .B2(\mem[13][2] ), 
        .ZN(n1084) );
  INV_X1 U302 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U303 ( .A1(data_in[3]), .A2(n842), .B1(n1086), .B2(\mem[13][3] ), 
        .ZN(n1083) );
  INV_X1 U304 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U305 ( .A1(data_in[4]), .A2(n842), .B1(n1086), .B2(\mem[13][4] ), 
        .ZN(n1082) );
  INV_X1 U306 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U307 ( .A1(data_in[5]), .A2(n842), .B1(n1086), .B2(\mem[13][5] ), 
        .ZN(n1081) );
  INV_X1 U308 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U309 ( .A1(data_in[6]), .A2(n842), .B1(n1086), .B2(\mem[13][6] ), 
        .ZN(n1080) );
  INV_X1 U310 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U311 ( .A1(data_in[7]), .A2(n842), .B1(n1086), .B2(\mem[13][7] ), 
        .ZN(n1079) );
  INV_X1 U312 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U313 ( .A1(data_in[0]), .A2(n841), .B1(n1077), .B2(\mem[14][0] ), 
        .ZN(n1078) );
  INV_X1 U314 ( .A(n1076), .ZN(n774) );
  AOI22_X1 U315 ( .A1(data_in[1]), .A2(n841), .B1(n1077), .B2(\mem[14][1] ), 
        .ZN(n1076) );
  INV_X1 U316 ( .A(n1075), .ZN(n773) );
  AOI22_X1 U317 ( .A1(data_in[2]), .A2(n841), .B1(n1077), .B2(\mem[14][2] ), 
        .ZN(n1075) );
  INV_X1 U318 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U319 ( .A1(data_in[3]), .A2(n841), .B1(n1077), .B2(\mem[14][3] ), 
        .ZN(n1074) );
  INV_X1 U320 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U321 ( .A1(data_in[4]), .A2(n841), .B1(n1077), .B2(\mem[14][4] ), 
        .ZN(n1073) );
  INV_X1 U322 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U323 ( .A1(data_in[5]), .A2(n841), .B1(n1077), .B2(\mem[14][5] ), 
        .ZN(n1072) );
  INV_X1 U324 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U325 ( .A1(data_in[6]), .A2(n841), .B1(n1077), .B2(\mem[14][6] ), 
        .ZN(n1071) );
  INV_X1 U326 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U327 ( .A1(data_in[7]), .A2(n841), .B1(n1077), .B2(\mem[14][7] ), 
        .ZN(n1070) );
  INV_X1 U328 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U329 ( .A1(data_in[0]), .A2(n840), .B1(n1068), .B2(\mem[15][0] ), 
        .ZN(n1069) );
  INV_X1 U330 ( .A(n1067), .ZN(n766) );
  AOI22_X1 U331 ( .A1(data_in[1]), .A2(n840), .B1(n1068), .B2(\mem[15][1] ), 
        .ZN(n1067) );
  INV_X1 U332 ( .A(n1066), .ZN(n765) );
  AOI22_X1 U333 ( .A1(data_in[2]), .A2(n840), .B1(n1068), .B2(\mem[15][2] ), 
        .ZN(n1066) );
  INV_X1 U334 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U335 ( .A1(data_in[3]), .A2(n840), .B1(n1068), .B2(\mem[15][3] ), 
        .ZN(n1065) );
  INV_X1 U336 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U337 ( .A1(data_in[4]), .A2(n840), .B1(n1068), .B2(\mem[15][4] ), 
        .ZN(n1064) );
  INV_X1 U338 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U339 ( .A1(data_in[5]), .A2(n840), .B1(n1068), .B2(\mem[15][5] ), 
        .ZN(n1063) );
  INV_X1 U340 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U341 ( .A1(data_in[6]), .A2(n840), .B1(n1068), .B2(\mem[15][6] ), 
        .ZN(n1062) );
  INV_X1 U342 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U343 ( .A1(data_in[7]), .A2(n840), .B1(n1068), .B2(\mem[15][7] ), 
        .ZN(n1061) );
  INV_X1 U344 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U345 ( .A1(data_in[0]), .A2(n839), .B1(n1059), .B2(\mem[16][0] ), 
        .ZN(n1060) );
  INV_X1 U346 ( .A(n1058), .ZN(n758) );
  AOI22_X1 U347 ( .A1(data_in[1]), .A2(n839), .B1(n1059), .B2(\mem[16][1] ), 
        .ZN(n1058) );
  INV_X1 U348 ( .A(n1057), .ZN(n757) );
  AOI22_X1 U349 ( .A1(data_in[2]), .A2(n839), .B1(n1059), .B2(\mem[16][2] ), 
        .ZN(n1057) );
  INV_X1 U350 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U351 ( .A1(data_in[3]), .A2(n839), .B1(n1059), .B2(\mem[16][3] ), 
        .ZN(n1056) );
  INV_X1 U352 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U353 ( .A1(data_in[4]), .A2(n839), .B1(n1059), .B2(\mem[16][4] ), 
        .ZN(n1055) );
  INV_X1 U354 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U355 ( .A1(data_in[5]), .A2(n839), .B1(n1059), .B2(\mem[16][5] ), 
        .ZN(n1054) );
  INV_X1 U356 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U357 ( .A1(data_in[6]), .A2(n839), .B1(n1059), .B2(\mem[16][6] ), 
        .ZN(n1053) );
  INV_X1 U358 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U359 ( .A1(data_in[7]), .A2(n839), .B1(n1059), .B2(\mem[16][7] ), 
        .ZN(n1052) );
  INV_X1 U360 ( .A(n1050), .ZN(n751) );
  AOI22_X1 U361 ( .A1(data_in[0]), .A2(n838), .B1(n1049), .B2(\mem[17][0] ), 
        .ZN(n1050) );
  INV_X1 U362 ( .A(n1048), .ZN(n750) );
  AOI22_X1 U363 ( .A1(data_in[1]), .A2(n838), .B1(n1049), .B2(\mem[17][1] ), 
        .ZN(n1048) );
  INV_X1 U364 ( .A(n1047), .ZN(n749) );
  AOI22_X1 U365 ( .A1(data_in[2]), .A2(n838), .B1(n1049), .B2(\mem[17][2] ), 
        .ZN(n1047) );
  INV_X1 U366 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U367 ( .A1(data_in[3]), .A2(n838), .B1(n1049), .B2(\mem[17][3] ), 
        .ZN(n1046) );
  INV_X1 U368 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U369 ( .A1(data_in[4]), .A2(n838), .B1(n1049), .B2(\mem[17][4] ), 
        .ZN(n1045) );
  INV_X1 U370 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U371 ( .A1(data_in[5]), .A2(n838), .B1(n1049), .B2(\mem[17][5] ), 
        .ZN(n1044) );
  INV_X1 U372 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U373 ( .A1(data_in[6]), .A2(n838), .B1(n1049), .B2(\mem[17][6] ), 
        .ZN(n1043) );
  INV_X1 U374 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U375 ( .A1(data_in[7]), .A2(n838), .B1(n1049), .B2(\mem[17][7] ), 
        .ZN(n1042) );
  INV_X1 U376 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U377 ( .A1(data_in[0]), .A2(n837), .B1(n1040), .B2(\mem[18][0] ), 
        .ZN(n1041) );
  INV_X1 U378 ( .A(n1039), .ZN(n742) );
  AOI22_X1 U379 ( .A1(data_in[1]), .A2(n837), .B1(n1040), .B2(\mem[18][1] ), 
        .ZN(n1039) );
  INV_X1 U380 ( .A(n1038), .ZN(n741) );
  AOI22_X1 U381 ( .A1(data_in[2]), .A2(n837), .B1(n1040), .B2(\mem[18][2] ), 
        .ZN(n1038) );
  INV_X1 U382 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U383 ( .A1(data_in[3]), .A2(n837), .B1(n1040), .B2(\mem[18][3] ), 
        .ZN(n1037) );
  INV_X1 U384 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U385 ( .A1(data_in[4]), .A2(n837), .B1(n1040), .B2(\mem[18][4] ), 
        .ZN(n1036) );
  INV_X1 U386 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U387 ( .A1(data_in[5]), .A2(n837), .B1(n1040), .B2(\mem[18][5] ), 
        .ZN(n1035) );
  INV_X1 U388 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U389 ( .A1(data_in[6]), .A2(n837), .B1(n1040), .B2(\mem[18][6] ), 
        .ZN(n1034) );
  INV_X1 U390 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U391 ( .A1(data_in[7]), .A2(n837), .B1(n1040), .B2(\mem[18][7] ), 
        .ZN(n1033) );
  INV_X1 U392 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U393 ( .A1(data_in[0]), .A2(n836), .B1(n1031), .B2(\mem[19][0] ), 
        .ZN(n1032) );
  INV_X1 U394 ( .A(n1030), .ZN(n734) );
  AOI22_X1 U395 ( .A1(data_in[1]), .A2(n836), .B1(n1031), .B2(\mem[19][1] ), 
        .ZN(n1030) );
  INV_X1 U396 ( .A(n1029), .ZN(n733) );
  AOI22_X1 U397 ( .A1(data_in[2]), .A2(n836), .B1(n1031), .B2(\mem[19][2] ), 
        .ZN(n1029) );
  INV_X1 U398 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U399 ( .A1(data_in[3]), .A2(n836), .B1(n1031), .B2(\mem[19][3] ), 
        .ZN(n1028) );
  INV_X1 U400 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U401 ( .A1(data_in[4]), .A2(n836), .B1(n1031), .B2(\mem[19][4] ), 
        .ZN(n1027) );
  INV_X1 U402 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U403 ( .A1(data_in[5]), .A2(n836), .B1(n1031), .B2(\mem[19][5] ), 
        .ZN(n1026) );
  INV_X1 U404 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U405 ( .A1(data_in[6]), .A2(n836), .B1(n1031), .B2(\mem[19][6] ), 
        .ZN(n1025) );
  INV_X1 U406 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U407 ( .A1(data_in[7]), .A2(n836), .B1(n1031), .B2(\mem[19][7] ), 
        .ZN(n1024) );
  INV_X1 U408 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U409 ( .A1(data_in[0]), .A2(n835), .B1(n1022), .B2(\mem[20][0] ), 
        .ZN(n1023) );
  INV_X1 U410 ( .A(n1021), .ZN(n726) );
  AOI22_X1 U411 ( .A1(data_in[1]), .A2(n835), .B1(n1022), .B2(\mem[20][1] ), 
        .ZN(n1021) );
  INV_X1 U412 ( .A(n1020), .ZN(n725) );
  AOI22_X1 U413 ( .A1(data_in[2]), .A2(n835), .B1(n1022), .B2(\mem[20][2] ), 
        .ZN(n1020) );
  INV_X1 U414 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U415 ( .A1(data_in[3]), .A2(n835), .B1(n1022), .B2(\mem[20][3] ), 
        .ZN(n1019) );
  INV_X1 U416 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U417 ( .A1(data_in[4]), .A2(n835), .B1(n1022), .B2(\mem[20][4] ), 
        .ZN(n1018) );
  INV_X1 U418 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U419 ( .A1(data_in[5]), .A2(n835), .B1(n1022), .B2(\mem[20][5] ), 
        .ZN(n1017) );
  INV_X1 U420 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U421 ( .A1(data_in[6]), .A2(n835), .B1(n1022), .B2(\mem[20][6] ), 
        .ZN(n1016) );
  INV_X1 U422 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U423 ( .A1(data_in[7]), .A2(n835), .B1(n1022), .B2(\mem[20][7] ), 
        .ZN(n1015) );
  INV_X1 U424 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U425 ( .A1(data_in[0]), .A2(n834), .B1(n1013), .B2(\mem[21][0] ), 
        .ZN(n1014) );
  INV_X1 U426 ( .A(n1012), .ZN(n718) );
  AOI22_X1 U427 ( .A1(data_in[1]), .A2(n834), .B1(n1013), .B2(\mem[21][1] ), 
        .ZN(n1012) );
  INV_X1 U428 ( .A(n1011), .ZN(n717) );
  AOI22_X1 U429 ( .A1(data_in[2]), .A2(n834), .B1(n1013), .B2(\mem[21][2] ), 
        .ZN(n1011) );
  INV_X1 U430 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U431 ( .A1(data_in[3]), .A2(n834), .B1(n1013), .B2(\mem[21][3] ), 
        .ZN(n1010) );
  INV_X1 U432 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U433 ( .A1(data_in[4]), .A2(n834), .B1(n1013), .B2(\mem[21][4] ), 
        .ZN(n1009) );
  INV_X1 U434 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U435 ( .A1(data_in[5]), .A2(n834), .B1(n1013), .B2(\mem[21][5] ), 
        .ZN(n1008) );
  INV_X1 U436 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U437 ( .A1(data_in[6]), .A2(n834), .B1(n1013), .B2(\mem[21][6] ), 
        .ZN(n1007) );
  INV_X1 U438 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U439 ( .A1(data_in[7]), .A2(n834), .B1(n1013), .B2(\mem[21][7] ), 
        .ZN(n1006) );
  INV_X1 U440 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U441 ( .A1(data_in[0]), .A2(n833), .B1(n1004), .B2(\mem[22][0] ), 
        .ZN(n1005) );
  INV_X1 U442 ( .A(n1003), .ZN(n710) );
  AOI22_X1 U443 ( .A1(data_in[1]), .A2(n833), .B1(n1004), .B2(\mem[22][1] ), 
        .ZN(n1003) );
  INV_X1 U444 ( .A(n1002), .ZN(n709) );
  AOI22_X1 U445 ( .A1(data_in[2]), .A2(n833), .B1(n1004), .B2(\mem[22][2] ), 
        .ZN(n1002) );
  INV_X1 U446 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U447 ( .A1(data_in[3]), .A2(n833), .B1(n1004), .B2(\mem[22][3] ), 
        .ZN(n1001) );
  INV_X1 U448 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U449 ( .A1(data_in[4]), .A2(n833), .B1(n1004), .B2(\mem[22][4] ), 
        .ZN(n1000) );
  INV_X1 U450 ( .A(n999), .ZN(n706) );
  AOI22_X1 U451 ( .A1(data_in[5]), .A2(n833), .B1(n1004), .B2(\mem[22][5] ), 
        .ZN(n999) );
  INV_X1 U452 ( .A(n998), .ZN(n705) );
  AOI22_X1 U453 ( .A1(data_in[6]), .A2(n833), .B1(n1004), .B2(\mem[22][6] ), 
        .ZN(n998) );
  INV_X1 U454 ( .A(n997), .ZN(n704) );
  AOI22_X1 U455 ( .A1(data_in[7]), .A2(n833), .B1(n1004), .B2(\mem[22][7] ), 
        .ZN(n997) );
  INV_X1 U456 ( .A(n996), .ZN(n703) );
  AOI22_X1 U457 ( .A1(data_in[0]), .A2(n832), .B1(n995), .B2(\mem[23][0] ), 
        .ZN(n996) );
  INV_X1 U458 ( .A(n994), .ZN(n702) );
  AOI22_X1 U459 ( .A1(data_in[1]), .A2(n832), .B1(n995), .B2(\mem[23][1] ), 
        .ZN(n994) );
  INV_X1 U460 ( .A(n993), .ZN(n701) );
  AOI22_X1 U461 ( .A1(data_in[2]), .A2(n832), .B1(n995), .B2(\mem[23][2] ), 
        .ZN(n993) );
  INV_X1 U462 ( .A(n992), .ZN(n700) );
  AOI22_X1 U463 ( .A1(data_in[3]), .A2(n832), .B1(n995), .B2(\mem[23][3] ), 
        .ZN(n992) );
  INV_X1 U464 ( .A(n991), .ZN(n699) );
  AOI22_X1 U465 ( .A1(data_in[4]), .A2(n832), .B1(n995), .B2(\mem[23][4] ), 
        .ZN(n991) );
  INV_X1 U466 ( .A(n990), .ZN(n698) );
  AOI22_X1 U467 ( .A1(data_in[5]), .A2(n832), .B1(n995), .B2(\mem[23][5] ), 
        .ZN(n990) );
  INV_X1 U468 ( .A(n989), .ZN(n697) );
  AOI22_X1 U469 ( .A1(data_in[6]), .A2(n832), .B1(n995), .B2(\mem[23][6] ), 
        .ZN(n989) );
  INV_X1 U470 ( .A(n988), .ZN(n696) );
  AOI22_X1 U471 ( .A1(data_in[7]), .A2(n832), .B1(n995), .B2(\mem[23][7] ), 
        .ZN(n988) );
  INV_X1 U472 ( .A(n987), .ZN(n695) );
  AOI22_X1 U473 ( .A1(data_in[0]), .A2(n831), .B1(n986), .B2(\mem[24][0] ), 
        .ZN(n987) );
  INV_X1 U474 ( .A(n985), .ZN(n694) );
  AOI22_X1 U475 ( .A1(data_in[1]), .A2(n831), .B1(n986), .B2(\mem[24][1] ), 
        .ZN(n985) );
  INV_X1 U476 ( .A(n984), .ZN(n693) );
  AOI22_X1 U477 ( .A1(data_in[2]), .A2(n831), .B1(n986), .B2(\mem[24][2] ), 
        .ZN(n984) );
  INV_X1 U478 ( .A(n983), .ZN(n692) );
  AOI22_X1 U479 ( .A1(data_in[3]), .A2(n831), .B1(n986), .B2(\mem[24][3] ), 
        .ZN(n983) );
  INV_X1 U480 ( .A(n982), .ZN(n691) );
  AOI22_X1 U481 ( .A1(data_in[4]), .A2(n831), .B1(n986), .B2(\mem[24][4] ), 
        .ZN(n982) );
  INV_X1 U482 ( .A(n981), .ZN(n690) );
  AOI22_X1 U483 ( .A1(data_in[5]), .A2(n831), .B1(n986), .B2(\mem[24][5] ), 
        .ZN(n981) );
  INV_X1 U484 ( .A(n980), .ZN(n689) );
  AOI22_X1 U485 ( .A1(data_in[6]), .A2(n831), .B1(n986), .B2(\mem[24][6] ), 
        .ZN(n980) );
  INV_X1 U486 ( .A(n979), .ZN(n688) );
  AOI22_X1 U487 ( .A1(data_in[7]), .A2(n831), .B1(n986), .B2(\mem[24][7] ), 
        .ZN(n979) );
  INV_X1 U488 ( .A(n977), .ZN(n687) );
  AOI22_X1 U489 ( .A1(data_in[0]), .A2(n830), .B1(n976), .B2(\mem[25][0] ), 
        .ZN(n977) );
  INV_X1 U490 ( .A(n975), .ZN(n686) );
  AOI22_X1 U491 ( .A1(data_in[1]), .A2(n830), .B1(n976), .B2(\mem[25][1] ), 
        .ZN(n975) );
  INV_X1 U492 ( .A(n974), .ZN(n685) );
  AOI22_X1 U493 ( .A1(data_in[2]), .A2(n830), .B1(n976), .B2(\mem[25][2] ), 
        .ZN(n974) );
  INV_X1 U494 ( .A(n973), .ZN(n684) );
  AOI22_X1 U495 ( .A1(data_in[3]), .A2(n830), .B1(n976), .B2(\mem[25][3] ), 
        .ZN(n973) );
  INV_X1 U496 ( .A(n972), .ZN(n683) );
  AOI22_X1 U497 ( .A1(data_in[4]), .A2(n830), .B1(n976), .B2(\mem[25][4] ), 
        .ZN(n972) );
  INV_X1 U498 ( .A(n971), .ZN(n682) );
  AOI22_X1 U499 ( .A1(data_in[5]), .A2(n830), .B1(n976), .B2(\mem[25][5] ), 
        .ZN(n971) );
  INV_X1 U500 ( .A(n970), .ZN(n681) );
  AOI22_X1 U501 ( .A1(data_in[6]), .A2(n830), .B1(n976), .B2(\mem[25][6] ), 
        .ZN(n970) );
  INV_X1 U502 ( .A(n969), .ZN(n680) );
  AOI22_X1 U503 ( .A1(data_in[7]), .A2(n830), .B1(n976), .B2(\mem[25][7] ), 
        .ZN(n969) );
  INV_X1 U504 ( .A(n968), .ZN(n679) );
  AOI22_X1 U505 ( .A1(data_in[0]), .A2(n829), .B1(n967), .B2(\mem[26][0] ), 
        .ZN(n968) );
  INV_X1 U506 ( .A(n966), .ZN(n678) );
  AOI22_X1 U507 ( .A1(data_in[1]), .A2(n829), .B1(n967), .B2(\mem[26][1] ), 
        .ZN(n966) );
  INV_X1 U508 ( .A(n965), .ZN(n677) );
  AOI22_X1 U509 ( .A1(data_in[2]), .A2(n829), .B1(n967), .B2(\mem[26][2] ), 
        .ZN(n965) );
  INV_X1 U510 ( .A(n964), .ZN(n676) );
  AOI22_X1 U511 ( .A1(data_in[3]), .A2(n829), .B1(n967), .B2(\mem[26][3] ), 
        .ZN(n964) );
  INV_X1 U512 ( .A(n963), .ZN(n675) );
  AOI22_X1 U513 ( .A1(data_in[4]), .A2(n829), .B1(n967), .B2(\mem[26][4] ), 
        .ZN(n963) );
  INV_X1 U514 ( .A(n962), .ZN(n674) );
  AOI22_X1 U515 ( .A1(data_in[5]), .A2(n829), .B1(n967), .B2(\mem[26][5] ), 
        .ZN(n962) );
  INV_X1 U516 ( .A(n961), .ZN(n673) );
  AOI22_X1 U517 ( .A1(data_in[6]), .A2(n829), .B1(n967), .B2(\mem[26][6] ), 
        .ZN(n961) );
  INV_X1 U518 ( .A(n960), .ZN(n672) );
  AOI22_X1 U519 ( .A1(data_in[7]), .A2(n829), .B1(n967), .B2(\mem[26][7] ), 
        .ZN(n960) );
  INV_X1 U520 ( .A(n959), .ZN(n671) );
  AOI22_X1 U521 ( .A1(data_in[0]), .A2(n828), .B1(n958), .B2(\mem[27][0] ), 
        .ZN(n959) );
  INV_X1 U522 ( .A(n957), .ZN(n670) );
  AOI22_X1 U523 ( .A1(data_in[1]), .A2(n828), .B1(n958), .B2(\mem[27][1] ), 
        .ZN(n957) );
  INV_X1 U524 ( .A(n956), .ZN(n669) );
  AOI22_X1 U525 ( .A1(data_in[2]), .A2(n828), .B1(n958), .B2(\mem[27][2] ), 
        .ZN(n956) );
  INV_X1 U526 ( .A(n955), .ZN(n668) );
  AOI22_X1 U527 ( .A1(data_in[3]), .A2(n828), .B1(n958), .B2(\mem[27][3] ), 
        .ZN(n955) );
  INV_X1 U528 ( .A(n954), .ZN(n667) );
  AOI22_X1 U529 ( .A1(data_in[4]), .A2(n828), .B1(n958), .B2(\mem[27][4] ), 
        .ZN(n954) );
  INV_X1 U530 ( .A(n953), .ZN(n666) );
  AOI22_X1 U531 ( .A1(data_in[5]), .A2(n828), .B1(n958), .B2(\mem[27][5] ), 
        .ZN(n953) );
  INV_X1 U532 ( .A(n952), .ZN(n665) );
  AOI22_X1 U533 ( .A1(data_in[6]), .A2(n828), .B1(n958), .B2(\mem[27][6] ), 
        .ZN(n952) );
  INV_X1 U534 ( .A(n951), .ZN(n664) );
  AOI22_X1 U535 ( .A1(data_in[7]), .A2(n828), .B1(n958), .B2(\mem[27][7] ), 
        .ZN(n951) );
  INV_X1 U536 ( .A(n950), .ZN(n663) );
  AOI22_X1 U537 ( .A1(data_in[0]), .A2(n827), .B1(n949), .B2(\mem[28][0] ), 
        .ZN(n950) );
  INV_X1 U538 ( .A(n948), .ZN(n662) );
  AOI22_X1 U539 ( .A1(data_in[1]), .A2(n827), .B1(n949), .B2(\mem[28][1] ), 
        .ZN(n948) );
  INV_X1 U540 ( .A(n947), .ZN(n661) );
  AOI22_X1 U541 ( .A1(data_in[2]), .A2(n827), .B1(n949), .B2(\mem[28][2] ), 
        .ZN(n947) );
  INV_X1 U542 ( .A(n946), .ZN(n660) );
  AOI22_X1 U543 ( .A1(data_in[3]), .A2(n827), .B1(n949), .B2(\mem[28][3] ), 
        .ZN(n946) );
  INV_X1 U544 ( .A(n945), .ZN(n659) );
  AOI22_X1 U545 ( .A1(data_in[4]), .A2(n827), .B1(n949), .B2(\mem[28][4] ), 
        .ZN(n945) );
  INV_X1 U546 ( .A(n944), .ZN(n658) );
  AOI22_X1 U547 ( .A1(data_in[5]), .A2(n827), .B1(n949), .B2(\mem[28][5] ), 
        .ZN(n944) );
  INV_X1 U548 ( .A(n943), .ZN(n657) );
  AOI22_X1 U549 ( .A1(data_in[6]), .A2(n827), .B1(n949), .B2(\mem[28][6] ), 
        .ZN(n943) );
  INV_X1 U550 ( .A(n942), .ZN(n656) );
  AOI22_X1 U551 ( .A1(data_in[7]), .A2(n827), .B1(n949), .B2(\mem[28][7] ), 
        .ZN(n942) );
  INV_X1 U552 ( .A(n941), .ZN(n655) );
  AOI22_X1 U553 ( .A1(data_in[0]), .A2(n826), .B1(n940), .B2(\mem[29][0] ), 
        .ZN(n941) );
  INV_X1 U554 ( .A(n939), .ZN(n654) );
  AOI22_X1 U555 ( .A1(data_in[1]), .A2(n826), .B1(n940), .B2(\mem[29][1] ), 
        .ZN(n939) );
  INV_X1 U556 ( .A(n938), .ZN(n653) );
  AOI22_X1 U557 ( .A1(data_in[2]), .A2(n826), .B1(n940), .B2(\mem[29][2] ), 
        .ZN(n938) );
  INV_X1 U558 ( .A(n937), .ZN(n652) );
  AOI22_X1 U559 ( .A1(data_in[3]), .A2(n826), .B1(n940), .B2(\mem[29][3] ), 
        .ZN(n937) );
  INV_X1 U560 ( .A(n936), .ZN(n651) );
  AOI22_X1 U561 ( .A1(data_in[4]), .A2(n826), .B1(n940), .B2(\mem[29][4] ), 
        .ZN(n936) );
  INV_X1 U562 ( .A(n935), .ZN(n650) );
  AOI22_X1 U563 ( .A1(data_in[5]), .A2(n826), .B1(n940), .B2(\mem[29][5] ), 
        .ZN(n935) );
  INV_X1 U564 ( .A(n934), .ZN(n649) );
  AOI22_X1 U565 ( .A1(data_in[6]), .A2(n826), .B1(n940), .B2(\mem[29][6] ), 
        .ZN(n934) );
  INV_X1 U566 ( .A(n933), .ZN(n648) );
  AOI22_X1 U567 ( .A1(data_in[7]), .A2(n826), .B1(n940), .B2(\mem[29][7] ), 
        .ZN(n933) );
  INV_X1 U568 ( .A(n932), .ZN(n647) );
  AOI22_X1 U569 ( .A1(data_in[0]), .A2(n825), .B1(n931), .B2(\mem[30][0] ), 
        .ZN(n932) );
  INV_X1 U570 ( .A(n930), .ZN(n646) );
  AOI22_X1 U571 ( .A1(data_in[1]), .A2(n825), .B1(n931), .B2(\mem[30][1] ), 
        .ZN(n930) );
  INV_X1 U572 ( .A(n929), .ZN(n645) );
  AOI22_X1 U573 ( .A1(data_in[2]), .A2(n825), .B1(n931), .B2(\mem[30][2] ), 
        .ZN(n929) );
  INV_X1 U574 ( .A(n928), .ZN(n644) );
  AOI22_X1 U575 ( .A1(data_in[3]), .A2(n825), .B1(n931), .B2(\mem[30][3] ), 
        .ZN(n928) );
  INV_X1 U576 ( .A(n927), .ZN(n643) );
  AOI22_X1 U577 ( .A1(data_in[4]), .A2(n825), .B1(n931), .B2(\mem[30][4] ), 
        .ZN(n927) );
  INV_X1 U578 ( .A(n926), .ZN(n642) );
  AOI22_X1 U579 ( .A1(data_in[5]), .A2(n825), .B1(n931), .B2(\mem[30][5] ), 
        .ZN(n926) );
  INV_X1 U580 ( .A(n925), .ZN(n641) );
  AOI22_X1 U581 ( .A1(data_in[6]), .A2(n825), .B1(n931), .B2(\mem[30][6] ), 
        .ZN(n925) );
  INV_X1 U582 ( .A(n924), .ZN(n640) );
  AOI22_X1 U583 ( .A1(data_in[7]), .A2(n825), .B1(n931), .B2(\mem[30][7] ), 
        .ZN(n924) );
  INV_X1 U584 ( .A(n923), .ZN(n639) );
  AOI22_X1 U585 ( .A1(data_in[0]), .A2(n824), .B1(n922), .B2(\mem[31][0] ), 
        .ZN(n923) );
  INV_X1 U586 ( .A(n921), .ZN(n638) );
  AOI22_X1 U587 ( .A1(data_in[1]), .A2(n824), .B1(n922), .B2(\mem[31][1] ), 
        .ZN(n921) );
  INV_X1 U588 ( .A(n920), .ZN(n637) );
  AOI22_X1 U589 ( .A1(data_in[2]), .A2(n824), .B1(n922), .B2(\mem[31][2] ), 
        .ZN(n920) );
  INV_X1 U590 ( .A(n919), .ZN(n636) );
  AOI22_X1 U591 ( .A1(data_in[3]), .A2(n824), .B1(n922), .B2(\mem[31][3] ), 
        .ZN(n919) );
  INV_X1 U592 ( .A(n918), .ZN(n635) );
  AOI22_X1 U593 ( .A1(data_in[4]), .A2(n824), .B1(n922), .B2(\mem[31][4] ), 
        .ZN(n918) );
  INV_X1 U594 ( .A(n917), .ZN(n634) );
  AOI22_X1 U595 ( .A1(data_in[5]), .A2(n824), .B1(n922), .B2(\mem[31][5] ), 
        .ZN(n917) );
  INV_X1 U596 ( .A(n916), .ZN(n633) );
  AOI22_X1 U597 ( .A1(data_in[6]), .A2(n824), .B1(n922), .B2(\mem[31][6] ), 
        .ZN(n916) );
  INV_X1 U598 ( .A(n915), .ZN(n632) );
  AOI22_X1 U599 ( .A1(data_in[7]), .A2(n824), .B1(n922), .B2(\mem[31][7] ), 
        .ZN(n915) );
  MUX2_X1 U600 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n614), .Z(n4) );
  MUX2_X1 U601 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n614), .Z(n5) );
  MUX2_X1 U602 ( .A(n5), .B(n4), .S(n611), .Z(n6) );
  MUX2_X1 U603 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n614), .Z(n7) );
  MUX2_X1 U604 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n614), .Z(n8) );
  MUX2_X1 U605 ( .A(n8), .B(n7), .S(n611), .Z(n9) );
  MUX2_X1 U606 ( .A(n9), .B(n6), .S(N12), .Z(n10) );
  MUX2_X1 U607 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n614), .Z(n11) );
  MUX2_X1 U608 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n614), .Z(n12) );
  MUX2_X1 U609 ( .A(n12), .B(n11), .S(n611), .Z(n13) );
  MUX2_X1 U610 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n614), .Z(n14) );
  MUX2_X1 U611 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n614), .Z(n15) );
  MUX2_X1 U612 ( .A(n15), .B(n14), .S(n611), .Z(n16) );
  MUX2_X1 U613 ( .A(n16), .B(n13), .S(n609), .Z(n17) );
  MUX2_X1 U614 ( .A(n17), .B(n10), .S(N13), .Z(n18) );
  MUX2_X1 U615 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n621), .Z(n19) );
  MUX2_X1 U616 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n621), .Z(n20) );
  MUX2_X1 U617 ( .A(n20), .B(n19), .S(n611), .Z(n21) );
  MUX2_X1 U618 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n621), .Z(n22) );
  MUX2_X1 U619 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n23) );
  MUX2_X1 U620 ( .A(n23), .B(n22), .S(N11), .Z(n24) );
  MUX2_X1 U621 ( .A(n24), .B(n21), .S(n610), .Z(n25) );
  MUX2_X1 U622 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n621), .Z(n26) );
  MUX2_X1 U623 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n27) );
  MUX2_X1 U624 ( .A(n27), .B(n26), .S(N11), .Z(n28) );
  MUX2_X1 U625 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n29) );
  MUX2_X1 U626 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n30) );
  MUX2_X1 U627 ( .A(n30), .B(n29), .S(n613), .Z(n31) );
  MUX2_X1 U628 ( .A(n31), .B(n28), .S(n610), .Z(n32) );
  MUX2_X1 U629 ( .A(n32), .B(n25), .S(N13), .Z(n33) );
  MUX2_X1 U630 ( .A(n33), .B(n18), .S(N14), .Z(N22) );
  MUX2_X1 U631 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n614), .Z(n34) );
  MUX2_X1 U632 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n614), .Z(n35) );
  MUX2_X1 U633 ( .A(n35), .B(n34), .S(n612), .Z(n36) );
  MUX2_X1 U634 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n614), .Z(n37) );
  MUX2_X1 U635 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n614), .Z(n38) );
  MUX2_X1 U636 ( .A(n38), .B(n37), .S(N11), .Z(n39) );
  MUX2_X1 U637 ( .A(n39), .B(n36), .S(N12), .Z(n40) );
  MUX2_X1 U638 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n615), .Z(n41) );
  MUX2_X1 U639 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(N10), .Z(n42) );
  MUX2_X1 U640 ( .A(n42), .B(n41), .S(n612), .Z(n43) );
  MUX2_X1 U641 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n621), .Z(n44) );
  MUX2_X1 U642 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n615), .Z(n45) );
  MUX2_X1 U643 ( .A(n45), .B(n44), .S(n613), .Z(n46) );
  MUX2_X1 U644 ( .A(n46), .B(n43), .S(n610), .Z(n47) );
  MUX2_X1 U645 ( .A(n47), .B(n40), .S(N13), .Z(n48) );
  MUX2_X1 U646 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n618), .Z(n49) );
  MUX2_X1 U647 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n617), .Z(n50) );
  MUX2_X1 U648 ( .A(n50), .B(n49), .S(n613), .Z(n51) );
  MUX2_X1 U649 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n620), .Z(n52) );
  MUX2_X1 U650 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n619), .Z(n53) );
  MUX2_X1 U651 ( .A(n53), .B(n52), .S(n611), .Z(n54) );
  MUX2_X1 U652 ( .A(n54), .B(n51), .S(n609), .Z(n55) );
  MUX2_X1 U653 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n621), .Z(n56) );
  MUX2_X1 U654 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n621), .Z(n57) );
  MUX2_X1 U655 ( .A(n57), .B(n56), .S(N11), .Z(n58) );
  MUX2_X1 U656 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n621), .Z(n59) );
  MUX2_X1 U657 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n621), .Z(n60) );
  MUX2_X1 U658 ( .A(n60), .B(n59), .S(n612), .Z(n61) );
  MUX2_X1 U659 ( .A(n61), .B(n58), .S(N12), .Z(n62) );
  MUX2_X1 U660 ( .A(n62), .B(n55), .S(N13), .Z(n63) );
  MUX2_X1 U661 ( .A(n63), .B(n48), .S(N14), .Z(N21) );
  MUX2_X1 U662 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n615), .Z(n64) );
  MUX2_X1 U663 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n615), .Z(n65) );
  MUX2_X1 U664 ( .A(n65), .B(n64), .S(n611), .Z(n66) );
  MUX2_X1 U665 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n615), .Z(n67) );
  MUX2_X1 U666 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n615), .Z(n68) );
  MUX2_X1 U667 ( .A(n68), .B(n67), .S(n611), .Z(n69) );
  MUX2_X1 U668 ( .A(n69), .B(n66), .S(n609), .Z(n70) );
  MUX2_X1 U669 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n615), .Z(n71) );
  MUX2_X1 U670 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n615), .Z(n72) );
  MUX2_X1 U671 ( .A(n72), .B(n71), .S(n611), .Z(n73) );
  MUX2_X1 U672 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n615), .Z(n74) );
  MUX2_X1 U673 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n615), .Z(n75) );
  MUX2_X1 U674 ( .A(n75), .B(n74), .S(n611), .Z(n76) );
  MUX2_X1 U675 ( .A(n76), .B(n73), .S(n609), .Z(n77) );
  MUX2_X1 U676 ( .A(n77), .B(n70), .S(N13), .Z(n78) );
  MUX2_X1 U677 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n615), .Z(n79) );
  MUX2_X1 U678 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n615), .Z(n80) );
  MUX2_X1 U679 ( .A(n80), .B(n79), .S(n611), .Z(n81) );
  MUX2_X1 U680 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n615), .Z(n82) );
  MUX2_X1 U681 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n615), .Z(n83) );
  MUX2_X1 U682 ( .A(n83), .B(n82), .S(n613), .Z(n84) );
  MUX2_X1 U683 ( .A(n84), .B(n81), .S(n609), .Z(n85) );
  MUX2_X1 U684 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n616), .Z(n86) );
  MUX2_X1 U685 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n616), .Z(n87) );
  MUX2_X1 U686 ( .A(n87), .B(n86), .S(n612), .Z(n88) );
  MUX2_X1 U687 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n616), .Z(n89) );
  MUX2_X1 U688 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n616), .Z(n90) );
  MUX2_X1 U689 ( .A(n90), .B(n89), .S(n611), .Z(n91) );
  MUX2_X1 U690 ( .A(n91), .B(n88), .S(n609), .Z(n92) );
  MUX2_X1 U691 ( .A(n92), .B(n85), .S(N13), .Z(n93) );
  MUX2_X1 U692 ( .A(n93), .B(n78), .S(N14), .Z(N20) );
  MUX2_X1 U693 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n616), .Z(n94) );
  MUX2_X1 U694 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n616), .Z(n95) );
  MUX2_X1 U695 ( .A(n95), .B(n94), .S(n611), .Z(n96) );
  MUX2_X1 U696 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n616), .Z(n97) );
  MUX2_X1 U697 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n616), .Z(n98) );
  MUX2_X1 U698 ( .A(n98), .B(n97), .S(n611), .Z(n99) );
  MUX2_X1 U699 ( .A(n99), .B(n96), .S(n609), .Z(n100) );
  MUX2_X1 U700 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n616), .Z(n101) );
  MUX2_X1 U701 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n616), .Z(n102) );
  MUX2_X1 U702 ( .A(n102), .B(n101), .S(n611), .Z(n103) );
  MUX2_X1 U703 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n616), .Z(n104) );
  MUX2_X1 U704 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n616), .Z(n105) );
  MUX2_X1 U705 ( .A(n105), .B(n104), .S(n613), .Z(n106) );
  MUX2_X1 U706 ( .A(n106), .B(n103), .S(n609), .Z(n107) );
  MUX2_X1 U707 ( .A(n107), .B(n100), .S(N13), .Z(n108) );
  MUX2_X1 U708 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n617), .Z(n109) );
  MUX2_X1 U709 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n617), .Z(n110) );
  MUX2_X1 U710 ( .A(n110), .B(n109), .S(n612), .Z(n111) );
  MUX2_X1 U711 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n617), .Z(n112) );
  MUX2_X1 U712 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n617), .Z(n113) );
  MUX2_X1 U713 ( .A(n113), .B(n112), .S(n612), .Z(n114) );
  MUX2_X1 U714 ( .A(n114), .B(n111), .S(n609), .Z(n115) );
  MUX2_X1 U715 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n617), .Z(n116) );
  MUX2_X1 U716 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n617), .Z(n117) );
  MUX2_X1 U717 ( .A(n117), .B(n116), .S(n612), .Z(n118) );
  MUX2_X1 U718 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n617), .Z(n119) );
  MUX2_X1 U719 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n617), .Z(n120) );
  MUX2_X1 U720 ( .A(n120), .B(n119), .S(n612), .Z(n121) );
  MUX2_X1 U721 ( .A(n121), .B(n118), .S(n609), .Z(n122) );
  MUX2_X1 U722 ( .A(n122), .B(n115), .S(N13), .Z(n123) );
  MUX2_X1 U723 ( .A(n123), .B(n108), .S(N14), .Z(N19) );
  MUX2_X1 U724 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n617), .Z(n124) );
  MUX2_X1 U725 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n617), .Z(n125) );
  MUX2_X1 U726 ( .A(n125), .B(n124), .S(n612), .Z(n126) );
  MUX2_X1 U727 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n617), .Z(n127) );
  MUX2_X1 U728 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n617), .Z(n128) );
  MUX2_X1 U729 ( .A(n128), .B(n127), .S(n612), .Z(n129) );
  MUX2_X1 U730 ( .A(n129), .B(n126), .S(n609), .Z(n130) );
  MUX2_X1 U731 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n615), .Z(n131) );
  MUX2_X1 U732 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n616), .Z(n132) );
  MUX2_X1 U733 ( .A(n132), .B(n131), .S(n612), .Z(n133) );
  MUX2_X1 U734 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n616), .Z(n134) );
  MUX2_X1 U735 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n614), .Z(n135) );
  MUX2_X1 U736 ( .A(n135), .B(n134), .S(n612), .Z(n136) );
  MUX2_X1 U737 ( .A(n136), .B(n133), .S(n609), .Z(n137) );
  MUX2_X1 U738 ( .A(n137), .B(n130), .S(N13), .Z(n138) );
  MUX2_X1 U739 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n616), .Z(n139) );
  MUX2_X1 U740 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n615), .Z(n140) );
  MUX2_X1 U741 ( .A(n140), .B(n139), .S(n612), .Z(n141) );
  MUX2_X1 U742 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n616), .Z(n142) );
  MUX2_X1 U743 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n614), .Z(n143) );
  MUX2_X1 U744 ( .A(n143), .B(n142), .S(n612), .Z(n144) );
  MUX2_X1 U745 ( .A(n144), .B(n141), .S(n609), .Z(n145) );
  MUX2_X1 U746 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n615), .Z(n146) );
  MUX2_X1 U747 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n617), .Z(n147) );
  MUX2_X1 U748 ( .A(n147), .B(n146), .S(n612), .Z(n148) );
  MUX2_X1 U749 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n615), .Z(n149) );
  MUX2_X1 U750 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n618), .Z(n150) );
  MUX2_X1 U751 ( .A(n150), .B(n149), .S(n612), .Z(n151) );
  MUX2_X1 U752 ( .A(n151), .B(n148), .S(n609), .Z(n152) );
  MUX2_X1 U753 ( .A(n152), .B(n145), .S(N13), .Z(n153) );
  MUX2_X1 U754 ( .A(n153), .B(n138), .S(N14), .Z(N18) );
  MUX2_X1 U755 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n616), .Z(n154) );
  MUX2_X1 U756 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n615), .Z(n155) );
  MUX2_X1 U757 ( .A(n155), .B(n154), .S(n613), .Z(n156) );
  MUX2_X1 U758 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n615), .Z(n157) );
  MUX2_X1 U759 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n615), .Z(n158) );
  MUX2_X1 U760 ( .A(n158), .B(n157), .S(n613), .Z(n159) );
  MUX2_X1 U761 ( .A(n159), .B(n156), .S(n610), .Z(n160) );
  MUX2_X1 U762 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n616), .Z(n161) );
  MUX2_X1 U763 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n616), .Z(n162) );
  MUX2_X1 U764 ( .A(n162), .B(n161), .S(n613), .Z(n163) );
  MUX2_X1 U765 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n615), .Z(n164) );
  MUX2_X1 U766 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n616), .Z(n165) );
  MUX2_X1 U767 ( .A(n165), .B(n164), .S(n613), .Z(n166) );
  MUX2_X1 U768 ( .A(n166), .B(n163), .S(n610), .Z(n167) );
  MUX2_X1 U769 ( .A(n167), .B(n160), .S(N13), .Z(n168) );
  MUX2_X1 U770 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n616), .Z(n169) );
  MUX2_X1 U771 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n616), .Z(n170) );
  MUX2_X1 U772 ( .A(n170), .B(n169), .S(n613), .Z(n171) );
  MUX2_X1 U773 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n616), .Z(n172) );
  MUX2_X1 U774 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n615), .Z(n173) );
  MUX2_X1 U775 ( .A(n173), .B(n172), .S(n613), .Z(n174) );
  MUX2_X1 U776 ( .A(n174), .B(n171), .S(n610), .Z(n175) );
  MUX2_X1 U777 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n618), .Z(n176) );
  MUX2_X1 U778 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n618), .Z(n177) );
  MUX2_X1 U779 ( .A(n177), .B(n176), .S(n613), .Z(n178) );
  MUX2_X1 U780 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n618), .Z(n179) );
  MUX2_X1 U781 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n618), .Z(n180) );
  MUX2_X1 U782 ( .A(n180), .B(n179), .S(n613), .Z(n181) );
  MUX2_X1 U783 ( .A(n181), .B(n178), .S(n610), .Z(n182) );
  MUX2_X1 U784 ( .A(n182), .B(n175), .S(N13), .Z(n183) );
  MUX2_X1 U785 ( .A(n183), .B(n168), .S(N14), .Z(N17) );
  MUX2_X1 U786 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n618), .Z(n184) );
  MUX2_X1 U787 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n618), .Z(n185) );
  MUX2_X1 U788 ( .A(n185), .B(n184), .S(n613), .Z(n186) );
  MUX2_X1 U789 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n618), .Z(n187) );
  MUX2_X1 U790 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n618), .Z(n188) );
  MUX2_X1 U791 ( .A(n188), .B(n187), .S(n613), .Z(n189) );
  MUX2_X1 U792 ( .A(n189), .B(n186), .S(n610), .Z(n190) );
  MUX2_X1 U793 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n618), .Z(n191) );
  MUX2_X1 U794 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n618), .Z(n192) );
  MUX2_X1 U795 ( .A(n192), .B(n191), .S(n613), .Z(n193) );
  MUX2_X1 U796 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n618), .Z(n194) );
  MUX2_X1 U797 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n618), .Z(n195) );
  MUX2_X1 U798 ( .A(n195), .B(n194), .S(n613), .Z(n196) );
  MUX2_X1 U799 ( .A(n196), .B(n193), .S(n610), .Z(n197) );
  MUX2_X1 U800 ( .A(n197), .B(n190), .S(N13), .Z(n198) );
  MUX2_X1 U801 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n619), .Z(n199) );
  MUX2_X1 U802 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n619), .Z(n200) );
  MUX2_X1 U803 ( .A(n200), .B(n199), .S(n612), .Z(n201) );
  MUX2_X1 U804 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n619), .Z(n202) );
  MUX2_X1 U805 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n619), .Z(n203) );
  MUX2_X1 U806 ( .A(n203), .B(n202), .S(n613), .Z(n204) );
  MUX2_X1 U807 ( .A(n204), .B(n201), .S(n610), .Z(n205) );
  MUX2_X1 U808 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n619), .Z(n206) );
  MUX2_X1 U809 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n619), .Z(n207) );
  MUX2_X1 U810 ( .A(n207), .B(n206), .S(n612), .Z(n208) );
  MUX2_X1 U811 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n619), .Z(n209) );
  MUX2_X1 U812 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n619), .Z(n210) );
  MUX2_X1 U813 ( .A(n210), .B(n209), .S(n611), .Z(n211) );
  MUX2_X1 U814 ( .A(n211), .B(n208), .S(n610), .Z(n212) );
  MUX2_X1 U815 ( .A(n212), .B(n205), .S(N13), .Z(n213) );
  MUX2_X1 U816 ( .A(n213), .B(n198), .S(N14), .Z(N16) );
  MUX2_X1 U817 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n619), .Z(n214) );
  MUX2_X1 U818 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n619), .Z(n215) );
  MUX2_X1 U819 ( .A(n215), .B(n214), .S(n613), .Z(n216) );
  MUX2_X1 U820 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n619), .Z(n217) );
  MUX2_X1 U821 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n619), .Z(n218) );
  MUX2_X1 U822 ( .A(n218), .B(n217), .S(n613), .Z(n219) );
  MUX2_X1 U823 ( .A(n219), .B(n216), .S(n610), .Z(n220) );
  MUX2_X1 U824 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n620), .Z(n221) );
  MUX2_X1 U825 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n620), .Z(n222) );
  MUX2_X1 U826 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U827 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n620), .Z(n224) );
  MUX2_X1 U828 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n620), .Z(n225) );
  MUX2_X1 U829 ( .A(n225), .B(n224), .S(n612), .Z(n226) );
  MUX2_X1 U830 ( .A(n226), .B(n223), .S(n610), .Z(n227) );
  MUX2_X1 U831 ( .A(n227), .B(n220), .S(N13), .Z(n228) );
  MUX2_X1 U832 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n620), .Z(n229) );
  MUX2_X1 U833 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n620), .Z(n595) );
  MUX2_X1 U834 ( .A(n595), .B(n229), .S(n611), .Z(n596) );
  MUX2_X1 U835 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n620), .Z(n597) );
  MUX2_X1 U836 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n620), .Z(n598) );
  MUX2_X1 U837 ( .A(n598), .B(n597), .S(n612), .Z(n599) );
  MUX2_X1 U838 ( .A(n599), .B(n596), .S(n610), .Z(n600) );
  MUX2_X1 U839 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n620), .Z(n601) );
  MUX2_X1 U840 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n620), .Z(n602) );
  MUX2_X1 U841 ( .A(n602), .B(n601), .S(n611), .Z(n603) );
  MUX2_X1 U842 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n620), .Z(n604) );
  MUX2_X1 U843 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n620), .Z(n605) );
  MUX2_X1 U844 ( .A(n605), .B(n604), .S(n613), .Z(n606) );
  MUX2_X1 U845 ( .A(n606), .B(n603), .S(n610), .Z(n607) );
  MUX2_X1 U846 ( .A(n607), .B(n600), .S(N13), .Z(n608) );
  MUX2_X1 U847 ( .A(n608), .B(n228), .S(N14), .Z(N15) );
  CLKBUF_X1 U848 ( .A(N11), .Z(n611) );
  INV_X1 U849 ( .A(N10), .ZN(n622) );
  INV_X1 U850 ( .A(N11), .ZN(n623) );
  INV_X1 U851 ( .A(data_in[0]), .ZN(n624) );
  INV_X1 U852 ( .A(data_in[1]), .ZN(n625) );
  INV_X1 U853 ( .A(data_in[2]), .ZN(n626) );
  INV_X1 U854 ( .A(data_in[3]), .ZN(n627) );
  INV_X1 U855 ( .A(data_in[4]), .ZN(n628) );
  INV_X1 U856 ( .A(data_in[5]), .ZN(n629) );
  INV_X1 U857 ( .A(data_in[6]), .ZN(n630) );
  INV_X1 U858 ( .A(data_in[7]), .ZN(n631) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_6 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n632), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n633), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n634), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n635), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n636), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n637), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n638), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n639), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n640), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n641), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n642), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n643), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n644), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n645), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n646), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n647), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n648), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n649), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n650), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n651), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n652), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n653), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n654), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n655), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n656), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n657), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n658), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n659), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n660), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n661), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n662), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n663), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n664), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n665), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n666), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n667), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n668), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n669), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n670), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n671), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n672), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n673), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n674), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n675), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n676), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n677), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n678), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n679), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n680), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n681), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n682), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n683), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n684), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n685), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n686), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n687), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n688), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n689), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n690), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n691), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n692), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n693), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n694), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n695), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n696), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n697), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n698), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n699), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n700), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n701), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n702), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n703), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n704), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n705), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n706), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n707), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n708), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n709), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n710), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n711), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n712), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n713), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n714), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n715), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n716), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n717), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n718), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n719), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n720), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n721), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n722), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n723), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n724), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n725), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n726), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n727), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n728), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n729), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n730), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n731), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n732), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n733), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n734), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n735), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n736), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n737), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n738), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n739), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n740), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n741), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n742), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n743), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n744), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n745), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n746), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n747), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n748), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n749), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n750), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n751), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n752), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n753), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n754), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n755), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n756), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n757), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n758), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n759), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n760), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n761), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n762), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n763), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n764), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n765), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n766), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n767), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n768), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n769), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n770), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n771), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n772), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n773), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n774), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n775), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n776), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n777), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n778), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n779), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n780), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n781), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n782), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n783), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n784), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n785), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n786), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n787), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n788), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n789), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n790), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n791), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n792), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n793), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n794), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n795), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n796), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n797), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n798), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n799), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n800), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n801), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n802), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n803), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n804), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n805), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n806), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n807), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n808), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n809), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n810), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n811), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n812), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n813), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n814), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n815), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n816), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n817), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n818), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n819), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n820), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n821), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n822), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n823), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n851), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n852), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n853), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n854), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n855), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n856), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n857), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n858), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n859), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n860), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n861), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n862), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n863), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n864), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n865), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n866), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n867), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n868), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n869), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n870), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n871), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n872), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n873), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n874), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n875), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n876), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n877), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n878), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n879), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n880), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n881), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n882), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n883), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n884), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n885), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n886), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n887), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n888), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n889), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n890), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n891), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n892), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n893), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n894), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n895), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n896), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n897), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n898), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n899), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n900), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n901), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n902), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n903), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n904), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n905), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n906), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n907), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n908), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n909), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n910), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n911), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n912), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n913), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n914), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n2) );
  BUF_X1 U3 ( .A(n621), .Z(n614) );
  INV_X2 U4 ( .A(n2), .ZN(data_out[3]) );
  BUF_X1 U5 ( .A(N10), .Z(n620) );
  BUF_X1 U6 ( .A(N10), .Z(n617) );
  BUF_X1 U7 ( .A(n621), .Z(n618) );
  BUF_X1 U8 ( .A(n621), .Z(n619) );
  BUF_X1 U9 ( .A(n621), .Z(n615) );
  BUF_X1 U10 ( .A(n621), .Z(n616) );
  BUF_X1 U11 ( .A(N11), .Z(n612) );
  BUF_X1 U12 ( .A(N11), .Z(n613) );
  BUF_X1 U13 ( .A(N10), .Z(n621) );
  NOR3_X1 U14 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1206) );
  NOR3_X1 U15 ( .A1(N11), .A2(N12), .A3(n622), .ZN(n1195) );
  NOR3_X1 U16 ( .A1(N10), .A2(N12), .A3(n623), .ZN(n1185) );
  NOR3_X1 U17 ( .A1(n622), .A2(N12), .A3(n623), .ZN(n1175) );
  INV_X1 U18 ( .A(n1132), .ZN(n847) );
  INV_X1 U19 ( .A(n1122), .ZN(n846) );
  INV_X1 U20 ( .A(n1113), .ZN(n845) );
  INV_X1 U21 ( .A(n1104), .ZN(n844) );
  INV_X1 U22 ( .A(n1059), .ZN(n839) );
  INV_X1 U23 ( .A(n1049), .ZN(n838) );
  INV_X1 U24 ( .A(n1040), .ZN(n837) );
  INV_X1 U25 ( .A(n1031), .ZN(n836) );
  INV_X1 U26 ( .A(n986), .ZN(n831) );
  INV_X1 U27 ( .A(n976), .ZN(n830) );
  INV_X1 U28 ( .A(n967), .ZN(n829) );
  INV_X1 U29 ( .A(n958), .ZN(n828) );
  INV_X1 U30 ( .A(n1095), .ZN(n843) );
  INV_X1 U31 ( .A(n1086), .ZN(n842) );
  INV_X1 U32 ( .A(n1077), .ZN(n841) );
  INV_X1 U33 ( .A(n1068), .ZN(n840) );
  INV_X1 U34 ( .A(n949), .ZN(n827) );
  INV_X1 U35 ( .A(n940), .ZN(n826) );
  INV_X1 U36 ( .A(n931), .ZN(n825) );
  INV_X1 U37 ( .A(n922), .ZN(n824) );
  INV_X1 U38 ( .A(n1022), .ZN(n835) );
  INV_X1 U39 ( .A(n1013), .ZN(n834) );
  INV_X1 U40 ( .A(n1004), .ZN(n833) );
  INV_X1 U41 ( .A(n995), .ZN(n832) );
  BUF_X1 U42 ( .A(N12), .Z(n610) );
  INV_X1 U43 ( .A(N13), .ZN(n849) );
  AND3_X1 U44 ( .A1(n622), .A2(n623), .A3(N12), .ZN(n1165) );
  AND3_X1 U45 ( .A1(N10), .A2(n623), .A3(N12), .ZN(n1155) );
  AND3_X1 U46 ( .A1(N11), .A2(n622), .A3(N12), .ZN(n1145) );
  AND3_X1 U47 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1135) );
  BUF_X1 U48 ( .A(N12), .Z(n609) );
  INV_X1 U49 ( .A(N14), .ZN(n850) );
  NAND2_X1 U50 ( .A1(n1195), .A2(n1205), .ZN(n1204) );
  NAND2_X1 U51 ( .A1(n1185), .A2(n1205), .ZN(n1194) );
  NAND2_X1 U52 ( .A1(n1175), .A2(n1205), .ZN(n1184) );
  NAND2_X1 U53 ( .A1(n1165), .A2(n1205), .ZN(n1174) );
  NAND2_X1 U54 ( .A1(n1155), .A2(n1205), .ZN(n1164) );
  NAND2_X1 U55 ( .A1(n1145), .A2(n1205), .ZN(n1154) );
  NAND2_X1 U56 ( .A1(n1135), .A2(n1205), .ZN(n1144) );
  NAND2_X1 U57 ( .A1(n1206), .A2(n1205), .ZN(n1215) );
  NAND2_X1 U58 ( .A1(n1124), .A2(n1206), .ZN(n1132) );
  NAND2_X1 U59 ( .A1(n1124), .A2(n1195), .ZN(n1122) );
  NAND2_X1 U60 ( .A1(n1124), .A2(n1185), .ZN(n1113) );
  NAND2_X1 U61 ( .A1(n1124), .A2(n1175), .ZN(n1104) );
  NAND2_X1 U62 ( .A1(n1051), .A2(n1206), .ZN(n1059) );
  NAND2_X1 U63 ( .A1(n1051), .A2(n1195), .ZN(n1049) );
  NAND2_X1 U64 ( .A1(n1051), .A2(n1185), .ZN(n1040) );
  NAND2_X1 U65 ( .A1(n1051), .A2(n1175), .ZN(n1031) );
  NAND2_X1 U66 ( .A1(n978), .A2(n1206), .ZN(n986) );
  NAND2_X1 U67 ( .A1(n978), .A2(n1195), .ZN(n976) );
  NAND2_X1 U68 ( .A1(n978), .A2(n1185), .ZN(n967) );
  NAND2_X1 U69 ( .A1(n978), .A2(n1175), .ZN(n958) );
  NAND2_X1 U70 ( .A1(n1124), .A2(n1165), .ZN(n1095) );
  NAND2_X1 U71 ( .A1(n1124), .A2(n1155), .ZN(n1086) );
  NAND2_X1 U72 ( .A1(n1124), .A2(n1145), .ZN(n1077) );
  NAND2_X1 U73 ( .A1(n1124), .A2(n1135), .ZN(n1068) );
  NAND2_X1 U74 ( .A1(n1051), .A2(n1165), .ZN(n1022) );
  NAND2_X1 U75 ( .A1(n1051), .A2(n1155), .ZN(n1013) );
  NAND2_X1 U76 ( .A1(n1051), .A2(n1145), .ZN(n1004) );
  NAND2_X1 U77 ( .A1(n1051), .A2(n1135), .ZN(n995) );
  NAND2_X1 U78 ( .A1(n978), .A2(n1165), .ZN(n949) );
  NAND2_X1 U79 ( .A1(n978), .A2(n1155), .ZN(n940) );
  NAND2_X1 U80 ( .A1(n978), .A2(n1145), .ZN(n931) );
  NAND2_X1 U81 ( .A1(n978), .A2(n1135), .ZN(n922) );
  AND3_X1 U82 ( .A1(n849), .A2(n850), .A3(n1134), .ZN(n1205) );
  AND3_X1 U83 ( .A1(N13), .A2(n1134), .A3(N14), .ZN(n978) );
  AND3_X1 U84 ( .A1(n1134), .A2(n850), .A3(N13), .ZN(n1124) );
  AND3_X1 U85 ( .A1(n1134), .A2(n849), .A3(N14), .ZN(n1051) );
  NOR2_X1 U86 ( .A1(n848), .A2(addr[5]), .ZN(n1134) );
  INV_X1 U87 ( .A(wr_en), .ZN(n848) );
  OAI21_X1 U88 ( .B1(n624), .B2(n1174), .A(n1173), .ZN(n882) );
  NAND2_X1 U89 ( .A1(\mem[4][0] ), .A2(n1174), .ZN(n1173) );
  OAI21_X1 U90 ( .B1(n625), .B2(n1174), .A(n1172), .ZN(n881) );
  NAND2_X1 U91 ( .A1(\mem[4][1] ), .A2(n1174), .ZN(n1172) );
  OAI21_X1 U92 ( .B1(n626), .B2(n1174), .A(n1171), .ZN(n880) );
  NAND2_X1 U93 ( .A1(\mem[4][2] ), .A2(n1174), .ZN(n1171) );
  OAI21_X1 U94 ( .B1(n627), .B2(n1174), .A(n1170), .ZN(n879) );
  NAND2_X1 U95 ( .A1(\mem[4][3] ), .A2(n1174), .ZN(n1170) );
  OAI21_X1 U96 ( .B1(n628), .B2(n1174), .A(n1169), .ZN(n878) );
  NAND2_X1 U97 ( .A1(\mem[4][4] ), .A2(n1174), .ZN(n1169) );
  OAI21_X1 U98 ( .B1(n629), .B2(n1174), .A(n1168), .ZN(n877) );
  NAND2_X1 U99 ( .A1(\mem[4][5] ), .A2(n1174), .ZN(n1168) );
  OAI21_X1 U100 ( .B1(n630), .B2(n1174), .A(n1167), .ZN(n876) );
  NAND2_X1 U101 ( .A1(\mem[4][6] ), .A2(n1174), .ZN(n1167) );
  OAI21_X1 U102 ( .B1(n631), .B2(n1174), .A(n1166), .ZN(n875) );
  NAND2_X1 U103 ( .A1(\mem[4][7] ), .A2(n1174), .ZN(n1166) );
  OAI21_X1 U104 ( .B1(n624), .B2(n1154), .A(n1153), .ZN(n866) );
  NAND2_X1 U105 ( .A1(\mem[6][0] ), .A2(n1154), .ZN(n1153) );
  OAI21_X1 U106 ( .B1(n625), .B2(n1154), .A(n1152), .ZN(n865) );
  NAND2_X1 U107 ( .A1(\mem[6][1] ), .A2(n1154), .ZN(n1152) );
  OAI21_X1 U108 ( .B1(n626), .B2(n1154), .A(n1151), .ZN(n864) );
  NAND2_X1 U109 ( .A1(\mem[6][2] ), .A2(n1154), .ZN(n1151) );
  OAI21_X1 U110 ( .B1(n627), .B2(n1154), .A(n1150), .ZN(n863) );
  NAND2_X1 U111 ( .A1(\mem[6][3] ), .A2(n1154), .ZN(n1150) );
  OAI21_X1 U112 ( .B1(n628), .B2(n1154), .A(n1149), .ZN(n862) );
  NAND2_X1 U113 ( .A1(\mem[6][4] ), .A2(n1154), .ZN(n1149) );
  OAI21_X1 U114 ( .B1(n629), .B2(n1154), .A(n1148), .ZN(n861) );
  NAND2_X1 U115 ( .A1(\mem[6][5] ), .A2(n1154), .ZN(n1148) );
  OAI21_X1 U116 ( .B1(n630), .B2(n1154), .A(n1147), .ZN(n860) );
  NAND2_X1 U117 ( .A1(\mem[6][6] ), .A2(n1154), .ZN(n1147) );
  OAI21_X1 U118 ( .B1(n631), .B2(n1154), .A(n1146), .ZN(n859) );
  NAND2_X1 U119 ( .A1(\mem[6][7] ), .A2(n1154), .ZN(n1146) );
  OAI21_X1 U120 ( .B1(n624), .B2(n1144), .A(n1143), .ZN(n858) );
  NAND2_X1 U121 ( .A1(\mem[7][0] ), .A2(n1144), .ZN(n1143) );
  OAI21_X1 U122 ( .B1(n625), .B2(n1144), .A(n1142), .ZN(n857) );
  NAND2_X1 U123 ( .A1(\mem[7][1] ), .A2(n1144), .ZN(n1142) );
  OAI21_X1 U124 ( .B1(n626), .B2(n1144), .A(n1141), .ZN(n856) );
  NAND2_X1 U125 ( .A1(\mem[7][2] ), .A2(n1144), .ZN(n1141) );
  OAI21_X1 U126 ( .B1(n627), .B2(n1144), .A(n1140), .ZN(n855) );
  NAND2_X1 U127 ( .A1(\mem[7][3] ), .A2(n1144), .ZN(n1140) );
  OAI21_X1 U128 ( .B1(n628), .B2(n1144), .A(n1139), .ZN(n854) );
  NAND2_X1 U129 ( .A1(\mem[7][4] ), .A2(n1144), .ZN(n1139) );
  OAI21_X1 U130 ( .B1(n629), .B2(n1144), .A(n1138), .ZN(n853) );
  NAND2_X1 U131 ( .A1(\mem[7][5] ), .A2(n1144), .ZN(n1138) );
  OAI21_X1 U132 ( .B1(n630), .B2(n1144), .A(n1137), .ZN(n852) );
  NAND2_X1 U133 ( .A1(\mem[7][6] ), .A2(n1144), .ZN(n1137) );
  OAI21_X1 U134 ( .B1(n631), .B2(n1144), .A(n1136), .ZN(n851) );
  NAND2_X1 U135 ( .A1(\mem[7][7] ), .A2(n1144), .ZN(n1136) );
  OAI21_X1 U136 ( .B1(n624), .B2(n1204), .A(n1203), .ZN(n906) );
  NAND2_X1 U137 ( .A1(\mem[1][0] ), .A2(n1204), .ZN(n1203) );
  OAI21_X1 U138 ( .B1(n625), .B2(n1204), .A(n1202), .ZN(n905) );
  NAND2_X1 U139 ( .A1(\mem[1][1] ), .A2(n1204), .ZN(n1202) );
  OAI21_X1 U140 ( .B1(n626), .B2(n1204), .A(n1201), .ZN(n904) );
  NAND2_X1 U141 ( .A1(\mem[1][2] ), .A2(n1204), .ZN(n1201) );
  OAI21_X1 U142 ( .B1(n627), .B2(n1204), .A(n1200), .ZN(n903) );
  NAND2_X1 U143 ( .A1(\mem[1][3] ), .A2(n1204), .ZN(n1200) );
  OAI21_X1 U144 ( .B1(n628), .B2(n1204), .A(n1199), .ZN(n902) );
  NAND2_X1 U145 ( .A1(\mem[1][4] ), .A2(n1204), .ZN(n1199) );
  OAI21_X1 U146 ( .B1(n629), .B2(n1204), .A(n1198), .ZN(n901) );
  NAND2_X1 U147 ( .A1(\mem[1][5] ), .A2(n1204), .ZN(n1198) );
  OAI21_X1 U148 ( .B1(n630), .B2(n1204), .A(n1197), .ZN(n900) );
  NAND2_X1 U149 ( .A1(\mem[1][6] ), .A2(n1204), .ZN(n1197) );
  OAI21_X1 U150 ( .B1(n631), .B2(n1204), .A(n1196), .ZN(n899) );
  NAND2_X1 U151 ( .A1(\mem[1][7] ), .A2(n1204), .ZN(n1196) );
  OAI21_X1 U152 ( .B1(n624), .B2(n1194), .A(n1193), .ZN(n898) );
  NAND2_X1 U153 ( .A1(\mem[2][0] ), .A2(n1194), .ZN(n1193) );
  OAI21_X1 U154 ( .B1(n625), .B2(n1194), .A(n1192), .ZN(n897) );
  NAND2_X1 U155 ( .A1(\mem[2][1] ), .A2(n1194), .ZN(n1192) );
  OAI21_X1 U156 ( .B1(n626), .B2(n1194), .A(n1191), .ZN(n896) );
  NAND2_X1 U157 ( .A1(\mem[2][2] ), .A2(n1194), .ZN(n1191) );
  OAI21_X1 U158 ( .B1(n627), .B2(n1194), .A(n1190), .ZN(n895) );
  NAND2_X1 U159 ( .A1(\mem[2][3] ), .A2(n1194), .ZN(n1190) );
  OAI21_X1 U160 ( .B1(n628), .B2(n1194), .A(n1189), .ZN(n894) );
  NAND2_X1 U161 ( .A1(\mem[2][4] ), .A2(n1194), .ZN(n1189) );
  OAI21_X1 U162 ( .B1(n629), .B2(n1194), .A(n1188), .ZN(n893) );
  NAND2_X1 U163 ( .A1(\mem[2][5] ), .A2(n1194), .ZN(n1188) );
  OAI21_X1 U164 ( .B1(n630), .B2(n1194), .A(n1187), .ZN(n892) );
  NAND2_X1 U165 ( .A1(\mem[2][6] ), .A2(n1194), .ZN(n1187) );
  OAI21_X1 U166 ( .B1(n631), .B2(n1194), .A(n1186), .ZN(n891) );
  NAND2_X1 U167 ( .A1(\mem[2][7] ), .A2(n1194), .ZN(n1186) );
  OAI21_X1 U168 ( .B1(n624), .B2(n1184), .A(n1183), .ZN(n890) );
  NAND2_X1 U169 ( .A1(\mem[3][0] ), .A2(n1184), .ZN(n1183) );
  OAI21_X1 U170 ( .B1(n625), .B2(n1184), .A(n1182), .ZN(n889) );
  NAND2_X1 U171 ( .A1(\mem[3][1] ), .A2(n1184), .ZN(n1182) );
  OAI21_X1 U172 ( .B1(n626), .B2(n1184), .A(n1181), .ZN(n888) );
  NAND2_X1 U173 ( .A1(\mem[3][2] ), .A2(n1184), .ZN(n1181) );
  OAI21_X1 U174 ( .B1(n627), .B2(n1184), .A(n1180), .ZN(n887) );
  NAND2_X1 U175 ( .A1(\mem[3][3] ), .A2(n1184), .ZN(n1180) );
  OAI21_X1 U176 ( .B1(n628), .B2(n1184), .A(n1179), .ZN(n886) );
  NAND2_X1 U177 ( .A1(\mem[3][4] ), .A2(n1184), .ZN(n1179) );
  OAI21_X1 U178 ( .B1(n629), .B2(n1184), .A(n1178), .ZN(n885) );
  NAND2_X1 U179 ( .A1(\mem[3][5] ), .A2(n1184), .ZN(n1178) );
  OAI21_X1 U180 ( .B1(n630), .B2(n1184), .A(n1177), .ZN(n884) );
  NAND2_X1 U181 ( .A1(\mem[3][6] ), .A2(n1184), .ZN(n1177) );
  OAI21_X1 U182 ( .B1(n631), .B2(n1184), .A(n1176), .ZN(n883) );
  NAND2_X1 U183 ( .A1(\mem[3][7] ), .A2(n1184), .ZN(n1176) );
  OAI21_X1 U184 ( .B1(n624), .B2(n1164), .A(n1163), .ZN(n874) );
  NAND2_X1 U185 ( .A1(\mem[5][0] ), .A2(n1164), .ZN(n1163) );
  OAI21_X1 U186 ( .B1(n625), .B2(n1164), .A(n1162), .ZN(n873) );
  NAND2_X1 U187 ( .A1(\mem[5][1] ), .A2(n1164), .ZN(n1162) );
  OAI21_X1 U188 ( .B1(n626), .B2(n1164), .A(n1161), .ZN(n872) );
  NAND2_X1 U189 ( .A1(\mem[5][2] ), .A2(n1164), .ZN(n1161) );
  OAI21_X1 U190 ( .B1(n627), .B2(n1164), .A(n1160), .ZN(n871) );
  NAND2_X1 U191 ( .A1(\mem[5][3] ), .A2(n1164), .ZN(n1160) );
  OAI21_X1 U192 ( .B1(n628), .B2(n1164), .A(n1159), .ZN(n870) );
  NAND2_X1 U193 ( .A1(\mem[5][4] ), .A2(n1164), .ZN(n1159) );
  OAI21_X1 U194 ( .B1(n629), .B2(n1164), .A(n1158), .ZN(n869) );
  NAND2_X1 U195 ( .A1(\mem[5][5] ), .A2(n1164), .ZN(n1158) );
  OAI21_X1 U196 ( .B1(n630), .B2(n1164), .A(n1157), .ZN(n868) );
  NAND2_X1 U197 ( .A1(\mem[5][6] ), .A2(n1164), .ZN(n1157) );
  OAI21_X1 U198 ( .B1(n631), .B2(n1164), .A(n1156), .ZN(n867) );
  NAND2_X1 U199 ( .A1(\mem[5][7] ), .A2(n1164), .ZN(n1156) );
  OAI21_X1 U200 ( .B1(n1215), .B2(n624), .A(n1214), .ZN(n914) );
  NAND2_X1 U201 ( .A1(\mem[0][0] ), .A2(n1215), .ZN(n1214) );
  OAI21_X1 U202 ( .B1(n1215), .B2(n625), .A(n1213), .ZN(n913) );
  NAND2_X1 U203 ( .A1(\mem[0][1] ), .A2(n1215), .ZN(n1213) );
  OAI21_X1 U204 ( .B1(n1215), .B2(n626), .A(n1212), .ZN(n912) );
  NAND2_X1 U205 ( .A1(\mem[0][2] ), .A2(n1215), .ZN(n1212) );
  OAI21_X1 U206 ( .B1(n1215), .B2(n627), .A(n1211), .ZN(n911) );
  NAND2_X1 U207 ( .A1(\mem[0][3] ), .A2(n1215), .ZN(n1211) );
  OAI21_X1 U208 ( .B1(n1215), .B2(n628), .A(n1210), .ZN(n910) );
  NAND2_X1 U209 ( .A1(\mem[0][4] ), .A2(n1215), .ZN(n1210) );
  OAI21_X1 U210 ( .B1(n1215), .B2(n629), .A(n1209), .ZN(n909) );
  NAND2_X1 U211 ( .A1(\mem[0][5] ), .A2(n1215), .ZN(n1209) );
  OAI21_X1 U212 ( .B1(n1215), .B2(n630), .A(n1208), .ZN(n908) );
  NAND2_X1 U213 ( .A1(\mem[0][6] ), .A2(n1215), .ZN(n1208) );
  OAI21_X1 U214 ( .B1(n1215), .B2(n631), .A(n1207), .ZN(n907) );
  NAND2_X1 U215 ( .A1(\mem[0][7] ), .A2(n1215), .ZN(n1207) );
  INV_X1 U216 ( .A(n1133), .ZN(n823) );
  AOI22_X1 U217 ( .A1(data_in[0]), .A2(n847), .B1(n1132), .B2(\mem[8][0] ), 
        .ZN(n1133) );
  INV_X1 U218 ( .A(n1131), .ZN(n822) );
  AOI22_X1 U219 ( .A1(data_in[1]), .A2(n847), .B1(n1132), .B2(\mem[8][1] ), 
        .ZN(n1131) );
  INV_X1 U220 ( .A(n1130), .ZN(n821) );
  AOI22_X1 U221 ( .A1(data_in[2]), .A2(n847), .B1(n1132), .B2(\mem[8][2] ), 
        .ZN(n1130) );
  INV_X1 U222 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U223 ( .A1(data_in[3]), .A2(n847), .B1(n1132), .B2(\mem[8][3] ), 
        .ZN(n1129) );
  INV_X1 U224 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U225 ( .A1(data_in[4]), .A2(n847), .B1(n1132), .B2(\mem[8][4] ), 
        .ZN(n1128) );
  INV_X1 U226 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U227 ( .A1(data_in[5]), .A2(n847), .B1(n1132), .B2(\mem[8][5] ), 
        .ZN(n1127) );
  INV_X1 U228 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U229 ( .A1(data_in[6]), .A2(n847), .B1(n1132), .B2(\mem[8][6] ), 
        .ZN(n1126) );
  INV_X1 U230 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U231 ( .A1(data_in[7]), .A2(n847), .B1(n1132), .B2(\mem[8][7] ), 
        .ZN(n1125) );
  INV_X1 U232 ( .A(n1123), .ZN(n815) );
  AOI22_X1 U233 ( .A1(data_in[0]), .A2(n846), .B1(n1122), .B2(\mem[9][0] ), 
        .ZN(n1123) );
  INV_X1 U234 ( .A(n1121), .ZN(n814) );
  AOI22_X1 U235 ( .A1(data_in[1]), .A2(n846), .B1(n1122), .B2(\mem[9][1] ), 
        .ZN(n1121) );
  INV_X1 U236 ( .A(n1120), .ZN(n813) );
  AOI22_X1 U237 ( .A1(data_in[2]), .A2(n846), .B1(n1122), .B2(\mem[9][2] ), 
        .ZN(n1120) );
  INV_X1 U238 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U239 ( .A1(data_in[3]), .A2(n846), .B1(n1122), .B2(\mem[9][3] ), 
        .ZN(n1119) );
  INV_X1 U240 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U241 ( .A1(data_in[4]), .A2(n846), .B1(n1122), .B2(\mem[9][4] ), 
        .ZN(n1118) );
  INV_X1 U242 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U243 ( .A1(data_in[5]), .A2(n846), .B1(n1122), .B2(\mem[9][5] ), 
        .ZN(n1117) );
  INV_X1 U244 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U245 ( .A1(data_in[6]), .A2(n846), .B1(n1122), .B2(\mem[9][6] ), 
        .ZN(n1116) );
  INV_X1 U246 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U247 ( .A1(data_in[7]), .A2(n846), .B1(n1122), .B2(\mem[9][7] ), 
        .ZN(n1115) );
  INV_X1 U248 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U249 ( .A1(data_in[0]), .A2(n845), .B1(n1113), .B2(\mem[10][0] ), 
        .ZN(n1114) );
  INV_X1 U250 ( .A(n1112), .ZN(n806) );
  AOI22_X1 U251 ( .A1(data_in[1]), .A2(n845), .B1(n1113), .B2(\mem[10][1] ), 
        .ZN(n1112) );
  INV_X1 U252 ( .A(n1111), .ZN(n805) );
  AOI22_X1 U253 ( .A1(data_in[2]), .A2(n845), .B1(n1113), .B2(\mem[10][2] ), 
        .ZN(n1111) );
  INV_X1 U254 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U255 ( .A1(data_in[3]), .A2(n845), .B1(n1113), .B2(\mem[10][3] ), 
        .ZN(n1110) );
  INV_X1 U256 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U257 ( .A1(data_in[4]), .A2(n845), .B1(n1113), .B2(\mem[10][4] ), 
        .ZN(n1109) );
  INV_X1 U258 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U259 ( .A1(data_in[5]), .A2(n845), .B1(n1113), .B2(\mem[10][5] ), 
        .ZN(n1108) );
  INV_X1 U260 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U261 ( .A1(data_in[6]), .A2(n845), .B1(n1113), .B2(\mem[10][6] ), 
        .ZN(n1107) );
  INV_X1 U262 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U263 ( .A1(data_in[7]), .A2(n845), .B1(n1113), .B2(\mem[10][7] ), 
        .ZN(n1106) );
  INV_X1 U264 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U265 ( .A1(data_in[0]), .A2(n844), .B1(n1104), .B2(\mem[11][0] ), 
        .ZN(n1105) );
  INV_X1 U266 ( .A(n1103), .ZN(n798) );
  AOI22_X1 U267 ( .A1(data_in[1]), .A2(n844), .B1(n1104), .B2(\mem[11][1] ), 
        .ZN(n1103) );
  INV_X1 U268 ( .A(n1102), .ZN(n797) );
  AOI22_X1 U269 ( .A1(data_in[2]), .A2(n844), .B1(n1104), .B2(\mem[11][2] ), 
        .ZN(n1102) );
  INV_X1 U270 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U271 ( .A1(data_in[3]), .A2(n844), .B1(n1104), .B2(\mem[11][3] ), 
        .ZN(n1101) );
  INV_X1 U272 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U273 ( .A1(data_in[4]), .A2(n844), .B1(n1104), .B2(\mem[11][4] ), 
        .ZN(n1100) );
  INV_X1 U274 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U275 ( .A1(data_in[5]), .A2(n844), .B1(n1104), .B2(\mem[11][5] ), 
        .ZN(n1099) );
  INV_X1 U276 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U277 ( .A1(data_in[6]), .A2(n844), .B1(n1104), .B2(\mem[11][6] ), 
        .ZN(n1098) );
  INV_X1 U278 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U279 ( .A1(data_in[7]), .A2(n844), .B1(n1104), .B2(\mem[11][7] ), 
        .ZN(n1097) );
  INV_X1 U280 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U281 ( .A1(data_in[0]), .A2(n843), .B1(n1095), .B2(\mem[12][0] ), 
        .ZN(n1096) );
  INV_X1 U282 ( .A(n1094), .ZN(n790) );
  AOI22_X1 U283 ( .A1(data_in[1]), .A2(n843), .B1(n1095), .B2(\mem[12][1] ), 
        .ZN(n1094) );
  INV_X1 U284 ( .A(n1093), .ZN(n789) );
  AOI22_X1 U285 ( .A1(data_in[2]), .A2(n843), .B1(n1095), .B2(\mem[12][2] ), 
        .ZN(n1093) );
  INV_X1 U286 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U287 ( .A1(data_in[3]), .A2(n843), .B1(n1095), .B2(\mem[12][3] ), 
        .ZN(n1092) );
  INV_X1 U288 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U289 ( .A1(data_in[4]), .A2(n843), .B1(n1095), .B2(\mem[12][4] ), 
        .ZN(n1091) );
  INV_X1 U290 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U291 ( .A1(data_in[5]), .A2(n843), .B1(n1095), .B2(\mem[12][5] ), 
        .ZN(n1090) );
  INV_X1 U292 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U293 ( .A1(data_in[6]), .A2(n843), .B1(n1095), .B2(\mem[12][6] ), 
        .ZN(n1089) );
  INV_X1 U294 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U295 ( .A1(data_in[7]), .A2(n843), .B1(n1095), .B2(\mem[12][7] ), 
        .ZN(n1088) );
  INV_X1 U296 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U297 ( .A1(data_in[0]), .A2(n842), .B1(n1086), .B2(\mem[13][0] ), 
        .ZN(n1087) );
  INV_X1 U298 ( .A(n1085), .ZN(n782) );
  AOI22_X1 U299 ( .A1(data_in[1]), .A2(n842), .B1(n1086), .B2(\mem[13][1] ), 
        .ZN(n1085) );
  INV_X1 U300 ( .A(n1084), .ZN(n781) );
  AOI22_X1 U301 ( .A1(data_in[2]), .A2(n842), .B1(n1086), .B2(\mem[13][2] ), 
        .ZN(n1084) );
  INV_X1 U302 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U303 ( .A1(data_in[3]), .A2(n842), .B1(n1086), .B2(\mem[13][3] ), 
        .ZN(n1083) );
  INV_X1 U304 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U305 ( .A1(data_in[4]), .A2(n842), .B1(n1086), .B2(\mem[13][4] ), 
        .ZN(n1082) );
  INV_X1 U306 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U307 ( .A1(data_in[5]), .A2(n842), .B1(n1086), .B2(\mem[13][5] ), 
        .ZN(n1081) );
  INV_X1 U308 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U309 ( .A1(data_in[6]), .A2(n842), .B1(n1086), .B2(\mem[13][6] ), 
        .ZN(n1080) );
  INV_X1 U310 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U311 ( .A1(data_in[7]), .A2(n842), .B1(n1086), .B2(\mem[13][7] ), 
        .ZN(n1079) );
  INV_X1 U312 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U313 ( .A1(data_in[0]), .A2(n841), .B1(n1077), .B2(\mem[14][0] ), 
        .ZN(n1078) );
  INV_X1 U314 ( .A(n1076), .ZN(n774) );
  AOI22_X1 U315 ( .A1(data_in[1]), .A2(n841), .B1(n1077), .B2(\mem[14][1] ), 
        .ZN(n1076) );
  INV_X1 U316 ( .A(n1075), .ZN(n773) );
  AOI22_X1 U317 ( .A1(data_in[2]), .A2(n841), .B1(n1077), .B2(\mem[14][2] ), 
        .ZN(n1075) );
  INV_X1 U318 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U319 ( .A1(data_in[3]), .A2(n841), .B1(n1077), .B2(\mem[14][3] ), 
        .ZN(n1074) );
  INV_X1 U320 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U321 ( .A1(data_in[4]), .A2(n841), .B1(n1077), .B2(\mem[14][4] ), 
        .ZN(n1073) );
  INV_X1 U322 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U323 ( .A1(data_in[5]), .A2(n841), .B1(n1077), .B2(\mem[14][5] ), 
        .ZN(n1072) );
  INV_X1 U324 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U325 ( .A1(data_in[6]), .A2(n841), .B1(n1077), .B2(\mem[14][6] ), 
        .ZN(n1071) );
  INV_X1 U326 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U327 ( .A1(data_in[7]), .A2(n841), .B1(n1077), .B2(\mem[14][7] ), 
        .ZN(n1070) );
  INV_X1 U328 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U329 ( .A1(data_in[0]), .A2(n840), .B1(n1068), .B2(\mem[15][0] ), 
        .ZN(n1069) );
  INV_X1 U330 ( .A(n1067), .ZN(n766) );
  AOI22_X1 U331 ( .A1(data_in[1]), .A2(n840), .B1(n1068), .B2(\mem[15][1] ), 
        .ZN(n1067) );
  INV_X1 U332 ( .A(n1066), .ZN(n765) );
  AOI22_X1 U333 ( .A1(data_in[2]), .A2(n840), .B1(n1068), .B2(\mem[15][2] ), 
        .ZN(n1066) );
  INV_X1 U334 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U335 ( .A1(data_in[3]), .A2(n840), .B1(n1068), .B2(\mem[15][3] ), 
        .ZN(n1065) );
  INV_X1 U336 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U337 ( .A1(data_in[4]), .A2(n840), .B1(n1068), .B2(\mem[15][4] ), 
        .ZN(n1064) );
  INV_X1 U338 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U339 ( .A1(data_in[5]), .A2(n840), .B1(n1068), .B2(\mem[15][5] ), 
        .ZN(n1063) );
  INV_X1 U340 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U341 ( .A1(data_in[6]), .A2(n840), .B1(n1068), .B2(\mem[15][6] ), 
        .ZN(n1062) );
  INV_X1 U342 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U343 ( .A1(data_in[7]), .A2(n840), .B1(n1068), .B2(\mem[15][7] ), 
        .ZN(n1061) );
  INV_X1 U344 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U345 ( .A1(data_in[0]), .A2(n839), .B1(n1059), .B2(\mem[16][0] ), 
        .ZN(n1060) );
  INV_X1 U346 ( .A(n1058), .ZN(n758) );
  AOI22_X1 U347 ( .A1(data_in[1]), .A2(n839), .B1(n1059), .B2(\mem[16][1] ), 
        .ZN(n1058) );
  INV_X1 U348 ( .A(n1057), .ZN(n757) );
  AOI22_X1 U349 ( .A1(data_in[2]), .A2(n839), .B1(n1059), .B2(\mem[16][2] ), 
        .ZN(n1057) );
  INV_X1 U350 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U351 ( .A1(data_in[3]), .A2(n839), .B1(n1059), .B2(\mem[16][3] ), 
        .ZN(n1056) );
  INV_X1 U352 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U353 ( .A1(data_in[4]), .A2(n839), .B1(n1059), .B2(\mem[16][4] ), 
        .ZN(n1055) );
  INV_X1 U354 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U355 ( .A1(data_in[5]), .A2(n839), .B1(n1059), .B2(\mem[16][5] ), 
        .ZN(n1054) );
  INV_X1 U356 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U357 ( .A1(data_in[6]), .A2(n839), .B1(n1059), .B2(\mem[16][6] ), 
        .ZN(n1053) );
  INV_X1 U358 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U359 ( .A1(data_in[7]), .A2(n839), .B1(n1059), .B2(\mem[16][7] ), 
        .ZN(n1052) );
  INV_X1 U360 ( .A(n1050), .ZN(n751) );
  AOI22_X1 U361 ( .A1(data_in[0]), .A2(n838), .B1(n1049), .B2(\mem[17][0] ), 
        .ZN(n1050) );
  INV_X1 U362 ( .A(n1048), .ZN(n750) );
  AOI22_X1 U363 ( .A1(data_in[1]), .A2(n838), .B1(n1049), .B2(\mem[17][1] ), 
        .ZN(n1048) );
  INV_X1 U364 ( .A(n1047), .ZN(n749) );
  AOI22_X1 U365 ( .A1(data_in[2]), .A2(n838), .B1(n1049), .B2(\mem[17][2] ), 
        .ZN(n1047) );
  INV_X1 U366 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U367 ( .A1(data_in[3]), .A2(n838), .B1(n1049), .B2(\mem[17][3] ), 
        .ZN(n1046) );
  INV_X1 U368 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U369 ( .A1(data_in[4]), .A2(n838), .B1(n1049), .B2(\mem[17][4] ), 
        .ZN(n1045) );
  INV_X1 U370 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U371 ( .A1(data_in[5]), .A2(n838), .B1(n1049), .B2(\mem[17][5] ), 
        .ZN(n1044) );
  INV_X1 U372 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U373 ( .A1(data_in[6]), .A2(n838), .B1(n1049), .B2(\mem[17][6] ), 
        .ZN(n1043) );
  INV_X1 U374 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U375 ( .A1(data_in[7]), .A2(n838), .B1(n1049), .B2(\mem[17][7] ), 
        .ZN(n1042) );
  INV_X1 U376 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U377 ( .A1(data_in[0]), .A2(n837), .B1(n1040), .B2(\mem[18][0] ), 
        .ZN(n1041) );
  INV_X1 U378 ( .A(n1039), .ZN(n742) );
  AOI22_X1 U379 ( .A1(data_in[1]), .A2(n837), .B1(n1040), .B2(\mem[18][1] ), 
        .ZN(n1039) );
  INV_X1 U380 ( .A(n1038), .ZN(n741) );
  AOI22_X1 U381 ( .A1(data_in[2]), .A2(n837), .B1(n1040), .B2(\mem[18][2] ), 
        .ZN(n1038) );
  INV_X1 U382 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U383 ( .A1(data_in[3]), .A2(n837), .B1(n1040), .B2(\mem[18][3] ), 
        .ZN(n1037) );
  INV_X1 U384 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U385 ( .A1(data_in[4]), .A2(n837), .B1(n1040), .B2(\mem[18][4] ), 
        .ZN(n1036) );
  INV_X1 U386 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U387 ( .A1(data_in[5]), .A2(n837), .B1(n1040), .B2(\mem[18][5] ), 
        .ZN(n1035) );
  INV_X1 U388 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U389 ( .A1(data_in[6]), .A2(n837), .B1(n1040), .B2(\mem[18][6] ), 
        .ZN(n1034) );
  INV_X1 U390 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U391 ( .A1(data_in[7]), .A2(n837), .B1(n1040), .B2(\mem[18][7] ), 
        .ZN(n1033) );
  INV_X1 U392 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U393 ( .A1(data_in[0]), .A2(n836), .B1(n1031), .B2(\mem[19][0] ), 
        .ZN(n1032) );
  INV_X1 U394 ( .A(n1030), .ZN(n734) );
  AOI22_X1 U395 ( .A1(data_in[1]), .A2(n836), .B1(n1031), .B2(\mem[19][1] ), 
        .ZN(n1030) );
  INV_X1 U396 ( .A(n1029), .ZN(n733) );
  AOI22_X1 U397 ( .A1(data_in[2]), .A2(n836), .B1(n1031), .B2(\mem[19][2] ), 
        .ZN(n1029) );
  INV_X1 U398 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U399 ( .A1(data_in[3]), .A2(n836), .B1(n1031), .B2(\mem[19][3] ), 
        .ZN(n1028) );
  INV_X1 U400 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U401 ( .A1(data_in[4]), .A2(n836), .B1(n1031), .B2(\mem[19][4] ), 
        .ZN(n1027) );
  INV_X1 U402 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U403 ( .A1(data_in[5]), .A2(n836), .B1(n1031), .B2(\mem[19][5] ), 
        .ZN(n1026) );
  INV_X1 U404 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U405 ( .A1(data_in[6]), .A2(n836), .B1(n1031), .B2(\mem[19][6] ), 
        .ZN(n1025) );
  INV_X1 U406 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U407 ( .A1(data_in[7]), .A2(n836), .B1(n1031), .B2(\mem[19][7] ), 
        .ZN(n1024) );
  INV_X1 U408 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U409 ( .A1(data_in[0]), .A2(n835), .B1(n1022), .B2(\mem[20][0] ), 
        .ZN(n1023) );
  INV_X1 U410 ( .A(n1021), .ZN(n726) );
  AOI22_X1 U411 ( .A1(data_in[1]), .A2(n835), .B1(n1022), .B2(\mem[20][1] ), 
        .ZN(n1021) );
  INV_X1 U412 ( .A(n1020), .ZN(n725) );
  AOI22_X1 U413 ( .A1(data_in[2]), .A2(n835), .B1(n1022), .B2(\mem[20][2] ), 
        .ZN(n1020) );
  INV_X1 U414 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U415 ( .A1(data_in[3]), .A2(n835), .B1(n1022), .B2(\mem[20][3] ), 
        .ZN(n1019) );
  INV_X1 U416 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U417 ( .A1(data_in[4]), .A2(n835), .B1(n1022), .B2(\mem[20][4] ), 
        .ZN(n1018) );
  INV_X1 U418 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U419 ( .A1(data_in[5]), .A2(n835), .B1(n1022), .B2(\mem[20][5] ), 
        .ZN(n1017) );
  INV_X1 U420 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U421 ( .A1(data_in[6]), .A2(n835), .B1(n1022), .B2(\mem[20][6] ), 
        .ZN(n1016) );
  INV_X1 U422 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U423 ( .A1(data_in[7]), .A2(n835), .B1(n1022), .B2(\mem[20][7] ), 
        .ZN(n1015) );
  INV_X1 U424 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U425 ( .A1(data_in[0]), .A2(n834), .B1(n1013), .B2(\mem[21][0] ), 
        .ZN(n1014) );
  INV_X1 U426 ( .A(n1012), .ZN(n718) );
  AOI22_X1 U427 ( .A1(data_in[1]), .A2(n834), .B1(n1013), .B2(\mem[21][1] ), 
        .ZN(n1012) );
  INV_X1 U428 ( .A(n1011), .ZN(n717) );
  AOI22_X1 U429 ( .A1(data_in[2]), .A2(n834), .B1(n1013), .B2(\mem[21][2] ), 
        .ZN(n1011) );
  INV_X1 U430 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U431 ( .A1(data_in[3]), .A2(n834), .B1(n1013), .B2(\mem[21][3] ), 
        .ZN(n1010) );
  INV_X1 U432 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U433 ( .A1(data_in[4]), .A2(n834), .B1(n1013), .B2(\mem[21][4] ), 
        .ZN(n1009) );
  INV_X1 U434 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U435 ( .A1(data_in[5]), .A2(n834), .B1(n1013), .B2(\mem[21][5] ), 
        .ZN(n1008) );
  INV_X1 U436 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U437 ( .A1(data_in[6]), .A2(n834), .B1(n1013), .B2(\mem[21][6] ), 
        .ZN(n1007) );
  INV_X1 U438 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U439 ( .A1(data_in[7]), .A2(n834), .B1(n1013), .B2(\mem[21][7] ), 
        .ZN(n1006) );
  INV_X1 U440 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U441 ( .A1(data_in[0]), .A2(n833), .B1(n1004), .B2(\mem[22][0] ), 
        .ZN(n1005) );
  INV_X1 U442 ( .A(n1003), .ZN(n710) );
  AOI22_X1 U443 ( .A1(data_in[1]), .A2(n833), .B1(n1004), .B2(\mem[22][1] ), 
        .ZN(n1003) );
  INV_X1 U444 ( .A(n1002), .ZN(n709) );
  AOI22_X1 U445 ( .A1(data_in[2]), .A2(n833), .B1(n1004), .B2(\mem[22][2] ), 
        .ZN(n1002) );
  INV_X1 U446 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U447 ( .A1(data_in[3]), .A2(n833), .B1(n1004), .B2(\mem[22][3] ), 
        .ZN(n1001) );
  INV_X1 U448 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U449 ( .A1(data_in[4]), .A2(n833), .B1(n1004), .B2(\mem[22][4] ), 
        .ZN(n1000) );
  INV_X1 U450 ( .A(n999), .ZN(n706) );
  AOI22_X1 U451 ( .A1(data_in[5]), .A2(n833), .B1(n1004), .B2(\mem[22][5] ), 
        .ZN(n999) );
  INV_X1 U452 ( .A(n998), .ZN(n705) );
  AOI22_X1 U453 ( .A1(data_in[6]), .A2(n833), .B1(n1004), .B2(\mem[22][6] ), 
        .ZN(n998) );
  INV_X1 U454 ( .A(n997), .ZN(n704) );
  AOI22_X1 U455 ( .A1(data_in[7]), .A2(n833), .B1(n1004), .B2(\mem[22][7] ), 
        .ZN(n997) );
  INV_X1 U456 ( .A(n996), .ZN(n703) );
  AOI22_X1 U457 ( .A1(data_in[0]), .A2(n832), .B1(n995), .B2(\mem[23][0] ), 
        .ZN(n996) );
  INV_X1 U458 ( .A(n994), .ZN(n702) );
  AOI22_X1 U459 ( .A1(data_in[1]), .A2(n832), .B1(n995), .B2(\mem[23][1] ), 
        .ZN(n994) );
  INV_X1 U460 ( .A(n993), .ZN(n701) );
  AOI22_X1 U461 ( .A1(data_in[2]), .A2(n832), .B1(n995), .B2(\mem[23][2] ), 
        .ZN(n993) );
  INV_X1 U462 ( .A(n992), .ZN(n700) );
  AOI22_X1 U463 ( .A1(data_in[3]), .A2(n832), .B1(n995), .B2(\mem[23][3] ), 
        .ZN(n992) );
  INV_X1 U464 ( .A(n991), .ZN(n699) );
  AOI22_X1 U465 ( .A1(data_in[4]), .A2(n832), .B1(n995), .B2(\mem[23][4] ), 
        .ZN(n991) );
  INV_X1 U466 ( .A(n990), .ZN(n698) );
  AOI22_X1 U467 ( .A1(data_in[5]), .A2(n832), .B1(n995), .B2(\mem[23][5] ), 
        .ZN(n990) );
  INV_X1 U468 ( .A(n989), .ZN(n697) );
  AOI22_X1 U469 ( .A1(data_in[6]), .A2(n832), .B1(n995), .B2(\mem[23][6] ), 
        .ZN(n989) );
  INV_X1 U470 ( .A(n988), .ZN(n696) );
  AOI22_X1 U471 ( .A1(data_in[7]), .A2(n832), .B1(n995), .B2(\mem[23][7] ), 
        .ZN(n988) );
  INV_X1 U472 ( .A(n987), .ZN(n695) );
  AOI22_X1 U473 ( .A1(data_in[0]), .A2(n831), .B1(n986), .B2(\mem[24][0] ), 
        .ZN(n987) );
  INV_X1 U474 ( .A(n985), .ZN(n694) );
  AOI22_X1 U475 ( .A1(data_in[1]), .A2(n831), .B1(n986), .B2(\mem[24][1] ), 
        .ZN(n985) );
  INV_X1 U476 ( .A(n984), .ZN(n693) );
  AOI22_X1 U477 ( .A1(data_in[2]), .A2(n831), .B1(n986), .B2(\mem[24][2] ), 
        .ZN(n984) );
  INV_X1 U478 ( .A(n983), .ZN(n692) );
  AOI22_X1 U479 ( .A1(data_in[3]), .A2(n831), .B1(n986), .B2(\mem[24][3] ), 
        .ZN(n983) );
  INV_X1 U480 ( .A(n982), .ZN(n691) );
  AOI22_X1 U481 ( .A1(data_in[4]), .A2(n831), .B1(n986), .B2(\mem[24][4] ), 
        .ZN(n982) );
  INV_X1 U482 ( .A(n981), .ZN(n690) );
  AOI22_X1 U483 ( .A1(data_in[5]), .A2(n831), .B1(n986), .B2(\mem[24][5] ), 
        .ZN(n981) );
  INV_X1 U484 ( .A(n980), .ZN(n689) );
  AOI22_X1 U485 ( .A1(data_in[6]), .A2(n831), .B1(n986), .B2(\mem[24][6] ), 
        .ZN(n980) );
  INV_X1 U486 ( .A(n979), .ZN(n688) );
  AOI22_X1 U487 ( .A1(data_in[7]), .A2(n831), .B1(n986), .B2(\mem[24][7] ), 
        .ZN(n979) );
  INV_X1 U488 ( .A(n977), .ZN(n687) );
  AOI22_X1 U489 ( .A1(data_in[0]), .A2(n830), .B1(n976), .B2(\mem[25][0] ), 
        .ZN(n977) );
  INV_X1 U490 ( .A(n975), .ZN(n686) );
  AOI22_X1 U491 ( .A1(data_in[1]), .A2(n830), .B1(n976), .B2(\mem[25][1] ), 
        .ZN(n975) );
  INV_X1 U492 ( .A(n974), .ZN(n685) );
  AOI22_X1 U493 ( .A1(data_in[2]), .A2(n830), .B1(n976), .B2(\mem[25][2] ), 
        .ZN(n974) );
  INV_X1 U494 ( .A(n973), .ZN(n684) );
  AOI22_X1 U495 ( .A1(data_in[3]), .A2(n830), .B1(n976), .B2(\mem[25][3] ), 
        .ZN(n973) );
  INV_X1 U496 ( .A(n972), .ZN(n683) );
  AOI22_X1 U497 ( .A1(data_in[4]), .A2(n830), .B1(n976), .B2(\mem[25][4] ), 
        .ZN(n972) );
  INV_X1 U498 ( .A(n971), .ZN(n682) );
  AOI22_X1 U499 ( .A1(data_in[5]), .A2(n830), .B1(n976), .B2(\mem[25][5] ), 
        .ZN(n971) );
  INV_X1 U500 ( .A(n970), .ZN(n681) );
  AOI22_X1 U501 ( .A1(data_in[6]), .A2(n830), .B1(n976), .B2(\mem[25][6] ), 
        .ZN(n970) );
  INV_X1 U502 ( .A(n969), .ZN(n680) );
  AOI22_X1 U503 ( .A1(data_in[7]), .A2(n830), .B1(n976), .B2(\mem[25][7] ), 
        .ZN(n969) );
  INV_X1 U504 ( .A(n968), .ZN(n679) );
  AOI22_X1 U505 ( .A1(data_in[0]), .A2(n829), .B1(n967), .B2(\mem[26][0] ), 
        .ZN(n968) );
  INV_X1 U506 ( .A(n966), .ZN(n678) );
  AOI22_X1 U507 ( .A1(data_in[1]), .A2(n829), .B1(n967), .B2(\mem[26][1] ), 
        .ZN(n966) );
  INV_X1 U508 ( .A(n965), .ZN(n677) );
  AOI22_X1 U509 ( .A1(data_in[2]), .A2(n829), .B1(n967), .B2(\mem[26][2] ), 
        .ZN(n965) );
  INV_X1 U510 ( .A(n964), .ZN(n676) );
  AOI22_X1 U511 ( .A1(data_in[3]), .A2(n829), .B1(n967), .B2(\mem[26][3] ), 
        .ZN(n964) );
  INV_X1 U512 ( .A(n963), .ZN(n675) );
  AOI22_X1 U513 ( .A1(data_in[4]), .A2(n829), .B1(n967), .B2(\mem[26][4] ), 
        .ZN(n963) );
  INV_X1 U514 ( .A(n962), .ZN(n674) );
  AOI22_X1 U515 ( .A1(data_in[5]), .A2(n829), .B1(n967), .B2(\mem[26][5] ), 
        .ZN(n962) );
  INV_X1 U516 ( .A(n961), .ZN(n673) );
  AOI22_X1 U517 ( .A1(data_in[6]), .A2(n829), .B1(n967), .B2(\mem[26][6] ), 
        .ZN(n961) );
  INV_X1 U518 ( .A(n960), .ZN(n672) );
  AOI22_X1 U519 ( .A1(data_in[7]), .A2(n829), .B1(n967), .B2(\mem[26][7] ), 
        .ZN(n960) );
  INV_X1 U520 ( .A(n959), .ZN(n671) );
  AOI22_X1 U521 ( .A1(data_in[0]), .A2(n828), .B1(n958), .B2(\mem[27][0] ), 
        .ZN(n959) );
  INV_X1 U522 ( .A(n957), .ZN(n670) );
  AOI22_X1 U523 ( .A1(data_in[1]), .A2(n828), .B1(n958), .B2(\mem[27][1] ), 
        .ZN(n957) );
  INV_X1 U524 ( .A(n956), .ZN(n669) );
  AOI22_X1 U525 ( .A1(data_in[2]), .A2(n828), .B1(n958), .B2(\mem[27][2] ), 
        .ZN(n956) );
  INV_X1 U526 ( .A(n955), .ZN(n668) );
  AOI22_X1 U527 ( .A1(data_in[3]), .A2(n828), .B1(n958), .B2(\mem[27][3] ), 
        .ZN(n955) );
  INV_X1 U528 ( .A(n954), .ZN(n667) );
  AOI22_X1 U529 ( .A1(data_in[4]), .A2(n828), .B1(n958), .B2(\mem[27][4] ), 
        .ZN(n954) );
  INV_X1 U530 ( .A(n953), .ZN(n666) );
  AOI22_X1 U531 ( .A1(data_in[5]), .A2(n828), .B1(n958), .B2(\mem[27][5] ), 
        .ZN(n953) );
  INV_X1 U532 ( .A(n952), .ZN(n665) );
  AOI22_X1 U533 ( .A1(data_in[6]), .A2(n828), .B1(n958), .B2(\mem[27][6] ), 
        .ZN(n952) );
  INV_X1 U534 ( .A(n951), .ZN(n664) );
  AOI22_X1 U535 ( .A1(data_in[7]), .A2(n828), .B1(n958), .B2(\mem[27][7] ), 
        .ZN(n951) );
  INV_X1 U536 ( .A(n950), .ZN(n663) );
  AOI22_X1 U537 ( .A1(data_in[0]), .A2(n827), .B1(n949), .B2(\mem[28][0] ), 
        .ZN(n950) );
  INV_X1 U538 ( .A(n948), .ZN(n662) );
  AOI22_X1 U539 ( .A1(data_in[1]), .A2(n827), .B1(n949), .B2(\mem[28][1] ), 
        .ZN(n948) );
  INV_X1 U540 ( .A(n947), .ZN(n661) );
  AOI22_X1 U541 ( .A1(data_in[2]), .A2(n827), .B1(n949), .B2(\mem[28][2] ), 
        .ZN(n947) );
  INV_X1 U542 ( .A(n946), .ZN(n660) );
  AOI22_X1 U543 ( .A1(data_in[3]), .A2(n827), .B1(n949), .B2(\mem[28][3] ), 
        .ZN(n946) );
  INV_X1 U544 ( .A(n945), .ZN(n659) );
  AOI22_X1 U545 ( .A1(data_in[4]), .A2(n827), .B1(n949), .B2(\mem[28][4] ), 
        .ZN(n945) );
  INV_X1 U546 ( .A(n944), .ZN(n658) );
  AOI22_X1 U547 ( .A1(data_in[5]), .A2(n827), .B1(n949), .B2(\mem[28][5] ), 
        .ZN(n944) );
  INV_X1 U548 ( .A(n943), .ZN(n657) );
  AOI22_X1 U549 ( .A1(data_in[6]), .A2(n827), .B1(n949), .B2(\mem[28][6] ), 
        .ZN(n943) );
  INV_X1 U550 ( .A(n942), .ZN(n656) );
  AOI22_X1 U551 ( .A1(data_in[7]), .A2(n827), .B1(n949), .B2(\mem[28][7] ), 
        .ZN(n942) );
  INV_X1 U552 ( .A(n941), .ZN(n655) );
  AOI22_X1 U553 ( .A1(data_in[0]), .A2(n826), .B1(n940), .B2(\mem[29][0] ), 
        .ZN(n941) );
  INV_X1 U554 ( .A(n939), .ZN(n654) );
  AOI22_X1 U555 ( .A1(data_in[1]), .A2(n826), .B1(n940), .B2(\mem[29][1] ), 
        .ZN(n939) );
  INV_X1 U556 ( .A(n938), .ZN(n653) );
  AOI22_X1 U557 ( .A1(data_in[2]), .A2(n826), .B1(n940), .B2(\mem[29][2] ), 
        .ZN(n938) );
  INV_X1 U558 ( .A(n937), .ZN(n652) );
  AOI22_X1 U559 ( .A1(data_in[3]), .A2(n826), .B1(n940), .B2(\mem[29][3] ), 
        .ZN(n937) );
  INV_X1 U560 ( .A(n936), .ZN(n651) );
  AOI22_X1 U561 ( .A1(data_in[4]), .A2(n826), .B1(n940), .B2(\mem[29][4] ), 
        .ZN(n936) );
  INV_X1 U562 ( .A(n935), .ZN(n650) );
  AOI22_X1 U563 ( .A1(data_in[5]), .A2(n826), .B1(n940), .B2(\mem[29][5] ), 
        .ZN(n935) );
  INV_X1 U564 ( .A(n934), .ZN(n649) );
  AOI22_X1 U565 ( .A1(data_in[6]), .A2(n826), .B1(n940), .B2(\mem[29][6] ), 
        .ZN(n934) );
  INV_X1 U566 ( .A(n933), .ZN(n648) );
  AOI22_X1 U567 ( .A1(data_in[7]), .A2(n826), .B1(n940), .B2(\mem[29][7] ), 
        .ZN(n933) );
  INV_X1 U568 ( .A(n932), .ZN(n647) );
  AOI22_X1 U569 ( .A1(data_in[0]), .A2(n825), .B1(n931), .B2(\mem[30][0] ), 
        .ZN(n932) );
  INV_X1 U570 ( .A(n930), .ZN(n646) );
  AOI22_X1 U571 ( .A1(data_in[1]), .A2(n825), .B1(n931), .B2(\mem[30][1] ), 
        .ZN(n930) );
  INV_X1 U572 ( .A(n929), .ZN(n645) );
  AOI22_X1 U573 ( .A1(data_in[2]), .A2(n825), .B1(n931), .B2(\mem[30][2] ), 
        .ZN(n929) );
  INV_X1 U574 ( .A(n928), .ZN(n644) );
  AOI22_X1 U575 ( .A1(data_in[3]), .A2(n825), .B1(n931), .B2(\mem[30][3] ), 
        .ZN(n928) );
  INV_X1 U576 ( .A(n927), .ZN(n643) );
  AOI22_X1 U577 ( .A1(data_in[4]), .A2(n825), .B1(n931), .B2(\mem[30][4] ), 
        .ZN(n927) );
  INV_X1 U578 ( .A(n926), .ZN(n642) );
  AOI22_X1 U579 ( .A1(data_in[5]), .A2(n825), .B1(n931), .B2(\mem[30][5] ), 
        .ZN(n926) );
  INV_X1 U580 ( .A(n925), .ZN(n641) );
  AOI22_X1 U581 ( .A1(data_in[6]), .A2(n825), .B1(n931), .B2(\mem[30][6] ), 
        .ZN(n925) );
  INV_X1 U582 ( .A(n924), .ZN(n640) );
  AOI22_X1 U583 ( .A1(data_in[7]), .A2(n825), .B1(n931), .B2(\mem[30][7] ), 
        .ZN(n924) );
  INV_X1 U584 ( .A(n923), .ZN(n639) );
  AOI22_X1 U585 ( .A1(data_in[0]), .A2(n824), .B1(n922), .B2(\mem[31][0] ), 
        .ZN(n923) );
  INV_X1 U586 ( .A(n921), .ZN(n638) );
  AOI22_X1 U587 ( .A1(data_in[1]), .A2(n824), .B1(n922), .B2(\mem[31][1] ), 
        .ZN(n921) );
  INV_X1 U588 ( .A(n920), .ZN(n637) );
  AOI22_X1 U589 ( .A1(data_in[2]), .A2(n824), .B1(n922), .B2(\mem[31][2] ), 
        .ZN(n920) );
  INV_X1 U590 ( .A(n919), .ZN(n636) );
  AOI22_X1 U591 ( .A1(data_in[3]), .A2(n824), .B1(n922), .B2(\mem[31][3] ), 
        .ZN(n919) );
  INV_X1 U592 ( .A(n918), .ZN(n635) );
  AOI22_X1 U593 ( .A1(data_in[4]), .A2(n824), .B1(n922), .B2(\mem[31][4] ), 
        .ZN(n918) );
  INV_X1 U594 ( .A(n917), .ZN(n634) );
  AOI22_X1 U595 ( .A1(data_in[5]), .A2(n824), .B1(n922), .B2(\mem[31][5] ), 
        .ZN(n917) );
  INV_X1 U596 ( .A(n916), .ZN(n633) );
  AOI22_X1 U597 ( .A1(data_in[6]), .A2(n824), .B1(n922), .B2(\mem[31][6] ), 
        .ZN(n916) );
  INV_X1 U598 ( .A(n915), .ZN(n632) );
  AOI22_X1 U599 ( .A1(data_in[7]), .A2(n824), .B1(n922), .B2(\mem[31][7] ), 
        .ZN(n915) );
  MUX2_X1 U600 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n614), .Z(n4) );
  MUX2_X1 U601 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n614), .Z(n5) );
  MUX2_X1 U602 ( .A(n5), .B(n4), .S(n611), .Z(n6) );
  MUX2_X1 U603 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n614), .Z(n7) );
  MUX2_X1 U604 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n614), .Z(n8) );
  MUX2_X1 U605 ( .A(n8), .B(n7), .S(n611), .Z(n9) );
  MUX2_X1 U606 ( .A(n9), .B(n6), .S(n609), .Z(n10) );
  MUX2_X1 U607 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n614), .Z(n11) );
  MUX2_X1 U608 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n614), .Z(n12) );
  MUX2_X1 U609 ( .A(n12), .B(n11), .S(n611), .Z(n13) );
  MUX2_X1 U610 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n614), .Z(n14) );
  MUX2_X1 U611 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n614), .Z(n15) );
  MUX2_X1 U612 ( .A(n15), .B(n14), .S(n611), .Z(n16) );
  MUX2_X1 U613 ( .A(n16), .B(n13), .S(n609), .Z(n17) );
  MUX2_X1 U614 ( .A(n17), .B(n10), .S(N13), .Z(n18) );
  MUX2_X1 U615 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n615), .Z(n19) );
  MUX2_X1 U616 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n615), .Z(n20) );
  MUX2_X1 U617 ( .A(n20), .B(n19), .S(n611), .Z(n21) );
  MUX2_X1 U618 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n615), .Z(n22) );
  MUX2_X1 U619 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n615), .Z(n23) );
  MUX2_X1 U620 ( .A(n23), .B(n22), .S(n612), .Z(n24) );
  MUX2_X1 U621 ( .A(n24), .B(n21), .S(n609), .Z(n25) );
  MUX2_X1 U622 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n615), .Z(n26) );
  MUX2_X1 U623 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n615), .Z(n27) );
  MUX2_X1 U624 ( .A(n27), .B(n26), .S(N11), .Z(n28) );
  MUX2_X1 U625 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n615), .Z(n29) );
  MUX2_X1 U626 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n615), .Z(n30) );
  MUX2_X1 U627 ( .A(n30), .B(n29), .S(n613), .Z(n31) );
  MUX2_X1 U628 ( .A(n31), .B(n28), .S(n609), .Z(n32) );
  MUX2_X1 U629 ( .A(n32), .B(n25), .S(N13), .Z(n33) );
  MUX2_X1 U630 ( .A(n33), .B(n18), .S(N14), .Z(N22) );
  MUX2_X1 U631 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n615), .Z(n34) );
  MUX2_X1 U632 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n615), .Z(n35) );
  MUX2_X1 U633 ( .A(n35), .B(n34), .S(n612), .Z(n36) );
  MUX2_X1 U634 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n615), .Z(n37) );
  MUX2_X1 U635 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n615), .Z(n38) );
  MUX2_X1 U636 ( .A(n38), .B(n37), .S(N11), .Z(n39) );
  MUX2_X1 U637 ( .A(n39), .B(n36), .S(n609), .Z(n40) );
  MUX2_X1 U638 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n616), .Z(n41) );
  MUX2_X1 U639 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n616), .Z(n42) );
  MUX2_X1 U640 ( .A(n42), .B(n41), .S(n611), .Z(n43) );
  MUX2_X1 U641 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n616), .Z(n44) );
  MUX2_X1 U642 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n616), .Z(n45) );
  MUX2_X1 U643 ( .A(n45), .B(n44), .S(N11), .Z(n46) );
  MUX2_X1 U644 ( .A(n46), .B(n43), .S(n609), .Z(n47) );
  MUX2_X1 U645 ( .A(n47), .B(n40), .S(N13), .Z(n48) );
  MUX2_X1 U646 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n616), .Z(n49) );
  MUX2_X1 U647 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n616), .Z(n50) );
  MUX2_X1 U648 ( .A(n50), .B(n49), .S(n613), .Z(n51) );
  MUX2_X1 U649 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n616), .Z(n52) );
  MUX2_X1 U650 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n616), .Z(n53) );
  MUX2_X1 U651 ( .A(n53), .B(n52), .S(n613), .Z(n54) );
  MUX2_X1 U652 ( .A(n54), .B(n51), .S(n609), .Z(n55) );
  MUX2_X1 U653 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n616), .Z(n56) );
  MUX2_X1 U654 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n616), .Z(n57) );
  MUX2_X1 U655 ( .A(n57), .B(n56), .S(n612), .Z(n58) );
  MUX2_X1 U656 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n616), .Z(n59) );
  MUX2_X1 U657 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n616), .Z(n60) );
  MUX2_X1 U658 ( .A(n60), .B(n59), .S(n612), .Z(n61) );
  MUX2_X1 U659 ( .A(n61), .B(n58), .S(n609), .Z(n62) );
  MUX2_X1 U660 ( .A(n62), .B(n55), .S(N13), .Z(n63) );
  MUX2_X1 U661 ( .A(n63), .B(n48), .S(N14), .Z(N21) );
  MUX2_X1 U662 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n620), .Z(n64) );
  MUX2_X1 U663 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n620), .Z(n65) );
  MUX2_X1 U664 ( .A(n65), .B(n64), .S(n611), .Z(n66) );
  MUX2_X1 U665 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n617), .Z(n67) );
  MUX2_X1 U666 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n617), .Z(n68) );
  MUX2_X1 U667 ( .A(n68), .B(n67), .S(n611), .Z(n69) );
  MUX2_X1 U668 ( .A(n69), .B(n66), .S(n609), .Z(n70) );
  MUX2_X1 U669 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n617), .Z(n71) );
  MUX2_X1 U670 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n619), .Z(n72) );
  MUX2_X1 U671 ( .A(n72), .B(n71), .S(n611), .Z(n73) );
  MUX2_X1 U672 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n621), .Z(n74) );
  MUX2_X1 U673 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n621), .Z(n75) );
  MUX2_X1 U674 ( .A(n75), .B(n74), .S(N11), .Z(n76) );
  MUX2_X1 U675 ( .A(n76), .B(n73), .S(N12), .Z(n77) );
  MUX2_X1 U676 ( .A(n77), .B(n70), .S(N13), .Z(n78) );
  MUX2_X1 U677 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n620), .Z(n79) );
  MUX2_X1 U678 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n620), .Z(n80) );
  MUX2_X1 U679 ( .A(n80), .B(n79), .S(n611), .Z(n81) );
  MUX2_X1 U680 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n618), .Z(n82) );
  MUX2_X1 U681 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n621), .Z(n83) );
  MUX2_X1 U682 ( .A(n83), .B(n82), .S(n612), .Z(n84) );
  MUX2_X1 U683 ( .A(n84), .B(n81), .S(n609), .Z(n85) );
  MUX2_X1 U684 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n617), .Z(n86) );
  MUX2_X1 U685 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n617), .Z(n87) );
  MUX2_X1 U686 ( .A(n87), .B(n86), .S(n612), .Z(n88) );
  MUX2_X1 U687 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n617), .Z(n89) );
  MUX2_X1 U688 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n620), .Z(n90) );
  MUX2_X1 U689 ( .A(n90), .B(n89), .S(n611), .Z(n91) );
  MUX2_X1 U690 ( .A(n91), .B(n88), .S(n609), .Z(n92) );
  MUX2_X1 U691 ( .A(n92), .B(n85), .S(N13), .Z(n93) );
  MUX2_X1 U692 ( .A(n93), .B(n78), .S(N14), .Z(N20) );
  MUX2_X1 U693 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n620), .Z(n94) );
  MUX2_X1 U694 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n620), .Z(n95) );
  MUX2_X1 U695 ( .A(n95), .B(n94), .S(n611), .Z(n96) );
  MUX2_X1 U696 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n617), .Z(n97) );
  MUX2_X1 U697 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n617), .Z(n98) );
  MUX2_X1 U698 ( .A(n98), .B(n97), .S(n611), .Z(n99) );
  MUX2_X1 U699 ( .A(n99), .B(n96), .S(n609), .Z(n100) );
  MUX2_X1 U700 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n617), .Z(n101) );
  MUX2_X1 U701 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n620), .Z(n102) );
  MUX2_X1 U702 ( .A(n102), .B(n101), .S(n611), .Z(n103) );
  MUX2_X1 U703 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n620), .Z(n104) );
  MUX2_X1 U704 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n617), .Z(n105) );
  MUX2_X1 U705 ( .A(n105), .B(n104), .S(n613), .Z(n106) );
  MUX2_X1 U706 ( .A(n106), .B(n103), .S(N12), .Z(n107) );
  MUX2_X1 U707 ( .A(n107), .B(n100), .S(N13), .Z(n108) );
  MUX2_X1 U708 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n617), .Z(n109) );
  MUX2_X1 U709 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n617), .Z(n110) );
  MUX2_X1 U710 ( .A(n110), .B(n109), .S(n612), .Z(n111) );
  MUX2_X1 U711 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n617), .Z(n112) );
  MUX2_X1 U712 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n617), .Z(n113) );
  MUX2_X1 U713 ( .A(n113), .B(n112), .S(n612), .Z(n114) );
  MUX2_X1 U714 ( .A(n114), .B(n111), .S(n609), .Z(n115) );
  MUX2_X1 U715 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n617), .Z(n116) );
  MUX2_X1 U716 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n617), .Z(n117) );
  MUX2_X1 U717 ( .A(n117), .B(n116), .S(n612), .Z(n118) );
  MUX2_X1 U718 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n617), .Z(n119) );
  MUX2_X1 U719 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n617), .Z(n120) );
  MUX2_X1 U720 ( .A(n120), .B(n119), .S(n612), .Z(n121) );
  MUX2_X1 U721 ( .A(n121), .B(n118), .S(n610), .Z(n122) );
  MUX2_X1 U722 ( .A(n122), .B(n115), .S(N13), .Z(n123) );
  MUX2_X1 U723 ( .A(n123), .B(n108), .S(N14), .Z(N19) );
  MUX2_X1 U724 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n617), .Z(n124) );
  MUX2_X1 U725 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n617), .Z(n125) );
  MUX2_X1 U726 ( .A(n125), .B(n124), .S(n612), .Z(n126) );
  MUX2_X1 U727 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n617), .Z(n127) );
  MUX2_X1 U728 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n617), .Z(n128) );
  MUX2_X1 U729 ( .A(n128), .B(n127), .S(n612), .Z(n129) );
  MUX2_X1 U730 ( .A(n129), .B(n126), .S(n609), .Z(n130) );
  MUX2_X1 U731 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n618), .Z(n131) );
  MUX2_X1 U732 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n618), .Z(n132) );
  MUX2_X1 U733 ( .A(n132), .B(n131), .S(n612), .Z(n133) );
  MUX2_X1 U734 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n618), .Z(n134) );
  MUX2_X1 U735 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n618), .Z(n135) );
  MUX2_X1 U736 ( .A(n135), .B(n134), .S(n612), .Z(n136) );
  MUX2_X1 U737 ( .A(n136), .B(n133), .S(N12), .Z(n137) );
  MUX2_X1 U738 ( .A(n137), .B(n130), .S(N13), .Z(n138) );
  MUX2_X1 U739 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n618), .Z(n139) );
  MUX2_X1 U740 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n618), .Z(n140) );
  MUX2_X1 U741 ( .A(n140), .B(n139), .S(n612), .Z(n141) );
  MUX2_X1 U742 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n618), .Z(n142) );
  MUX2_X1 U743 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n618), .Z(n143) );
  MUX2_X1 U744 ( .A(n143), .B(n142), .S(n612), .Z(n144) );
  MUX2_X1 U745 ( .A(n144), .B(n141), .S(n610), .Z(n145) );
  MUX2_X1 U746 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n618), .Z(n146) );
  MUX2_X1 U747 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n618), .Z(n147) );
  MUX2_X1 U748 ( .A(n147), .B(n146), .S(n612), .Z(n148) );
  MUX2_X1 U749 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n618), .Z(n149) );
  MUX2_X1 U750 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n618), .Z(n150) );
  MUX2_X1 U751 ( .A(n150), .B(n149), .S(n612), .Z(n151) );
  MUX2_X1 U752 ( .A(n151), .B(n148), .S(n609), .Z(n152) );
  MUX2_X1 U753 ( .A(n152), .B(n145), .S(N13), .Z(n153) );
  MUX2_X1 U754 ( .A(n153), .B(n138), .S(N14), .Z(N18) );
  MUX2_X1 U755 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n619), .Z(n154) );
  MUX2_X1 U756 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n619), .Z(n155) );
  MUX2_X1 U757 ( .A(n155), .B(n154), .S(n613), .Z(n156) );
  MUX2_X1 U758 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n619), .Z(n157) );
  MUX2_X1 U759 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n619), .Z(n158) );
  MUX2_X1 U760 ( .A(n158), .B(n157), .S(n613), .Z(n159) );
  MUX2_X1 U761 ( .A(n159), .B(n156), .S(n610), .Z(n160) );
  MUX2_X1 U762 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n619), .Z(n161) );
  MUX2_X1 U763 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n619), .Z(n162) );
  MUX2_X1 U764 ( .A(n162), .B(n161), .S(n613), .Z(n163) );
  MUX2_X1 U765 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n619), .Z(n164) );
  MUX2_X1 U766 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n619), .Z(n165) );
  MUX2_X1 U767 ( .A(n165), .B(n164), .S(n613), .Z(n166) );
  MUX2_X1 U768 ( .A(n166), .B(n163), .S(n610), .Z(n167) );
  MUX2_X1 U769 ( .A(n167), .B(n160), .S(N13), .Z(n168) );
  MUX2_X1 U770 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n619), .Z(n169) );
  MUX2_X1 U771 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n619), .Z(n170) );
  MUX2_X1 U772 ( .A(n170), .B(n169), .S(n613), .Z(n171) );
  MUX2_X1 U773 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n619), .Z(n172) );
  MUX2_X1 U774 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n619), .Z(n173) );
  MUX2_X1 U775 ( .A(n173), .B(n172), .S(n613), .Z(n174) );
  MUX2_X1 U776 ( .A(n174), .B(n171), .S(n610), .Z(n175) );
  MUX2_X1 U777 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n621), .Z(n176) );
  MUX2_X1 U778 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n621), .Z(n177) );
  MUX2_X1 U779 ( .A(n177), .B(n176), .S(n613), .Z(n178) );
  MUX2_X1 U780 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n621), .Z(n179) );
  MUX2_X1 U781 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n621), .Z(n180) );
  MUX2_X1 U782 ( .A(n180), .B(n179), .S(n613), .Z(n181) );
  MUX2_X1 U783 ( .A(n181), .B(n178), .S(n610), .Z(n182) );
  MUX2_X1 U784 ( .A(n182), .B(n175), .S(N13), .Z(n183) );
  MUX2_X1 U785 ( .A(n183), .B(n168), .S(N14), .Z(N17) );
  MUX2_X1 U786 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n617), .Z(n184) );
  MUX2_X1 U787 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n614), .Z(n185) );
  MUX2_X1 U788 ( .A(n185), .B(n184), .S(n613), .Z(n186) );
  MUX2_X1 U789 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n618), .Z(n187) );
  MUX2_X1 U790 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n621), .Z(n188) );
  MUX2_X1 U791 ( .A(n188), .B(n187), .S(n613), .Z(n189) );
  MUX2_X1 U792 ( .A(n189), .B(n186), .S(n610), .Z(n190) );
  MUX2_X1 U793 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n620), .Z(n191) );
  MUX2_X1 U794 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(N10), .Z(n192) );
  MUX2_X1 U795 ( .A(n192), .B(n191), .S(n613), .Z(n193) );
  MUX2_X1 U796 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n621), .Z(n194) );
  MUX2_X1 U797 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n620), .Z(n195) );
  MUX2_X1 U798 ( .A(n195), .B(n194), .S(n613), .Z(n196) );
  MUX2_X1 U799 ( .A(n196), .B(n193), .S(n610), .Z(n197) );
  MUX2_X1 U800 ( .A(n197), .B(n190), .S(N13), .Z(n198) );
  MUX2_X1 U801 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n614), .Z(n199) );
  MUX2_X1 U802 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n621), .Z(n200) );
  MUX2_X1 U803 ( .A(n200), .B(n199), .S(n612), .Z(n201) );
  MUX2_X1 U804 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n615), .Z(n202) );
  MUX2_X1 U805 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n203) );
  MUX2_X1 U806 ( .A(n203), .B(n202), .S(n613), .Z(n204) );
  MUX2_X1 U807 ( .A(n204), .B(n201), .S(n610), .Z(n205) );
  MUX2_X1 U808 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n206) );
  MUX2_X1 U809 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n207) );
  MUX2_X1 U810 ( .A(n207), .B(n206), .S(n613), .Z(n208) );
  MUX2_X1 U811 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n614), .Z(n209) );
  MUX2_X1 U812 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n614), .Z(n210) );
  MUX2_X1 U813 ( .A(n210), .B(n209), .S(n611), .Z(n211) );
  MUX2_X1 U814 ( .A(n211), .B(n208), .S(n610), .Z(n212) );
  MUX2_X1 U815 ( .A(n212), .B(n205), .S(N13), .Z(n213) );
  MUX2_X1 U816 ( .A(n213), .B(n198), .S(N14), .Z(N16) );
  MUX2_X1 U817 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n614), .Z(n214) );
  MUX2_X1 U818 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n616), .Z(n215) );
  MUX2_X1 U819 ( .A(n215), .B(n214), .S(n613), .Z(n216) );
  MUX2_X1 U820 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n621), .Z(n217) );
  MUX2_X1 U821 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n218) );
  MUX2_X1 U822 ( .A(n218), .B(n217), .S(N11), .Z(n219) );
  MUX2_X1 U823 ( .A(n219), .B(n216), .S(n610), .Z(n220) );
  MUX2_X1 U824 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n620), .Z(n221) );
  MUX2_X1 U825 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n620), .Z(n222) );
  MUX2_X1 U826 ( .A(n222), .B(n221), .S(n611), .Z(n223) );
  MUX2_X1 U827 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n620), .Z(n224) );
  MUX2_X1 U828 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n620), .Z(n225) );
  MUX2_X1 U829 ( .A(n225), .B(n224), .S(n612), .Z(n226) );
  MUX2_X1 U830 ( .A(n226), .B(n223), .S(n610), .Z(n227) );
  MUX2_X1 U831 ( .A(n227), .B(n220), .S(N13), .Z(n228) );
  MUX2_X1 U832 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n620), .Z(n229) );
  MUX2_X1 U833 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n620), .Z(n595) );
  MUX2_X1 U834 ( .A(n595), .B(n229), .S(n613), .Z(n596) );
  MUX2_X1 U835 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n620), .Z(n597) );
  MUX2_X1 U836 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n620), .Z(n598) );
  MUX2_X1 U837 ( .A(n598), .B(n597), .S(n611), .Z(n599) );
  MUX2_X1 U838 ( .A(n599), .B(n596), .S(n610), .Z(n600) );
  MUX2_X1 U839 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n620), .Z(n601) );
  MUX2_X1 U840 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n620), .Z(n602) );
  MUX2_X1 U841 ( .A(n602), .B(n601), .S(n611), .Z(n603) );
  MUX2_X1 U842 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n620), .Z(n604) );
  MUX2_X1 U843 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n620), .Z(n605) );
  MUX2_X1 U844 ( .A(n605), .B(n604), .S(n612), .Z(n606) );
  MUX2_X1 U845 ( .A(n606), .B(n603), .S(n610), .Z(n607) );
  MUX2_X1 U846 ( .A(n607), .B(n600), .S(N13), .Z(n608) );
  MUX2_X1 U847 ( .A(n608), .B(n228), .S(N14), .Z(N15) );
  CLKBUF_X1 U848 ( .A(N11), .Z(n611) );
  INV_X1 U849 ( .A(N10), .ZN(n622) );
  INV_X1 U850 ( .A(N11), .ZN(n623) );
  INV_X1 U851 ( .A(data_in[0]), .ZN(n624) );
  INV_X1 U852 ( .A(data_in[1]), .ZN(n625) );
  INV_X1 U853 ( .A(data_in[2]), .ZN(n626) );
  INV_X1 U854 ( .A(data_in[3]), .ZN(n627) );
  INV_X1 U855 ( .A(data_in[4]), .ZN(n628) );
  INV_X1 U856 ( .A(data_in[5]), .ZN(n629) );
  INV_X1 U857 ( .A(data_in[6]), .ZN(n630) );
  INV_X1 U858 ( .A(data_in[7]), .ZN(n631) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_5 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n630), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n631), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n632), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n633), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n634), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n635), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n636), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n637), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n638), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n639), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n640), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n641), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n642), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n643), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n644), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n645), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n646), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n647), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n648), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n649), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n650), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n651), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n652), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n653), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n654), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n655), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n656), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n657), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n658), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n659), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n660), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n661), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n662), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n663), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n664), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n665), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n666), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n667), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n668), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n669), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n670), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n671), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n672), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n673), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n674), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n675), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n676), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n677), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n678), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n679), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n680), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n681), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n682), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n683), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n684), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n685), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n686), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n687), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n688), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n689), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n690), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n691), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n692), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n693), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n694), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n695), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n696), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n697), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n698), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n699), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n700), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n701), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n702), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n703), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n704), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n705), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n706), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n707), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n708), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n709), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n710), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n711), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n712), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n713), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n714), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n715), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n716), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n717), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n718), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n719), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n720), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n721), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n722), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n723), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n724), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n725), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n726), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n727), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n728), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n729), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n730), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n731), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n732), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n733), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n734), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n735), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n736), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n737), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n738), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n739), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n740), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n741), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n742), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n743), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n744), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n745), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n746), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n747), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n748), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n749), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n750), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n751), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n752), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n753), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n754), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n755), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n756), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n757), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n758), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n759), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n760), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n761), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n762), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n763), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n764), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n765), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n766), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n767), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n768), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n769), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n770), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n771), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n772), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n773), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n774), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n775), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n776), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n777), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n778), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n779), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n780), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n781), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n782), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n783), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n784), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n785), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n786), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n787), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n788), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n789), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n790), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n791), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n792), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n793), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n794), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n795), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n796), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n797), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n798), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n799), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n800), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n801), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n802), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n803), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n804), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n805), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n806), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n807), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n808), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n809), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n810), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n811), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n812), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n813), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n814), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n815), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n816), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n817), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n818), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n819), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n820), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n821), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n849), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n850), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n851), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n852), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n853), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n854), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n855), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n856), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n857), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n858), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n859), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n860), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n861), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n862), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n863), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n864), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n865), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n866), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n867), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n868), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n869), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n870), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n871), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n872), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n873), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n874), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n875), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n876), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n877), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n878), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n879), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n880), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n881), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n882), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n883), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n884), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n885), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n886), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n887), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n888), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n889), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n890), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n891), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n892), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n893), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n894), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n895), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n896), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n897), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n898), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n899), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n900), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n901), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n902), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n903), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n904), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n905), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n906), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n907), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n908), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n909), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n910), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n911), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n912), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  CLKBUF_X1 U3 ( .A(N10), .Z(n619) );
  BUF_X1 U4 ( .A(N10), .Z(n613) );
  INV_X2 U5 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U6 ( .A(n619), .Z(n618) );
  BUF_X1 U7 ( .A(N10), .Z(n615) );
  BUF_X1 U8 ( .A(N10), .Z(n614) );
  BUF_X1 U9 ( .A(n619), .Z(n616) );
  BUF_X1 U10 ( .A(N10), .Z(n617) );
  BUF_X1 U11 ( .A(N11), .Z(n611) );
  BUF_X1 U12 ( .A(N11), .Z(n612) );
  NOR3_X1 U13 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1204) );
  NOR3_X1 U14 ( .A1(N11), .A2(N12), .A3(n620), .ZN(n1193) );
  NOR3_X1 U15 ( .A1(N10), .A2(N12), .A3(n621), .ZN(n1183) );
  NOR3_X1 U16 ( .A1(n620), .A2(N12), .A3(n621), .ZN(n1173) );
  INV_X1 U17 ( .A(n1130), .ZN(n845) );
  INV_X1 U18 ( .A(n1120), .ZN(n844) );
  INV_X1 U19 ( .A(n1111), .ZN(n843) );
  INV_X1 U20 ( .A(n1102), .ZN(n842) );
  INV_X1 U21 ( .A(n1057), .ZN(n837) );
  INV_X1 U22 ( .A(n1047), .ZN(n836) );
  INV_X1 U23 ( .A(n1038), .ZN(n835) );
  INV_X1 U24 ( .A(n1029), .ZN(n834) );
  INV_X1 U25 ( .A(n984), .ZN(n829) );
  INV_X1 U26 ( .A(n974), .ZN(n828) );
  INV_X1 U27 ( .A(n965), .ZN(n827) );
  INV_X1 U28 ( .A(n956), .ZN(n826) );
  INV_X1 U29 ( .A(n1093), .ZN(n841) );
  INV_X1 U30 ( .A(n1084), .ZN(n840) );
  INV_X1 U31 ( .A(n1075), .ZN(n839) );
  INV_X1 U32 ( .A(n1066), .ZN(n838) );
  INV_X1 U33 ( .A(n947), .ZN(n825) );
  INV_X1 U34 ( .A(n938), .ZN(n824) );
  INV_X1 U35 ( .A(n929), .ZN(n823) );
  INV_X1 U36 ( .A(n920), .ZN(n822) );
  INV_X1 U37 ( .A(n1020), .ZN(n833) );
  INV_X1 U38 ( .A(n1011), .ZN(n832) );
  INV_X1 U39 ( .A(n1002), .ZN(n831) );
  INV_X1 U40 ( .A(n993), .ZN(n830) );
  BUF_X1 U41 ( .A(N12), .Z(n608) );
  BUF_X1 U42 ( .A(N12), .Z(n609) );
  INV_X1 U43 ( .A(N13), .ZN(n847) );
  AND3_X1 U44 ( .A1(n620), .A2(n621), .A3(N12), .ZN(n1163) );
  AND3_X1 U45 ( .A1(N10), .A2(n621), .A3(N12), .ZN(n1153) );
  AND3_X1 U46 ( .A1(N11), .A2(n620), .A3(N12), .ZN(n1143) );
  AND3_X1 U47 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1133) );
  INV_X1 U48 ( .A(N14), .ZN(n848) );
  NAND2_X1 U49 ( .A1(n1193), .A2(n1203), .ZN(n1202) );
  NAND2_X1 U50 ( .A1(n1183), .A2(n1203), .ZN(n1192) );
  NAND2_X1 U51 ( .A1(n1173), .A2(n1203), .ZN(n1182) );
  NAND2_X1 U52 ( .A1(n1163), .A2(n1203), .ZN(n1172) );
  NAND2_X1 U53 ( .A1(n1153), .A2(n1203), .ZN(n1162) );
  NAND2_X1 U54 ( .A1(n1143), .A2(n1203), .ZN(n1152) );
  NAND2_X1 U55 ( .A1(n1133), .A2(n1203), .ZN(n1142) );
  NAND2_X1 U56 ( .A1(n1204), .A2(n1203), .ZN(n1213) );
  NAND2_X1 U57 ( .A1(n1122), .A2(n1204), .ZN(n1130) );
  NAND2_X1 U58 ( .A1(n1122), .A2(n1193), .ZN(n1120) );
  NAND2_X1 U59 ( .A1(n1122), .A2(n1183), .ZN(n1111) );
  NAND2_X1 U60 ( .A1(n1122), .A2(n1173), .ZN(n1102) );
  NAND2_X1 U61 ( .A1(n1049), .A2(n1204), .ZN(n1057) );
  NAND2_X1 U62 ( .A1(n1049), .A2(n1193), .ZN(n1047) );
  NAND2_X1 U63 ( .A1(n1049), .A2(n1183), .ZN(n1038) );
  NAND2_X1 U64 ( .A1(n1049), .A2(n1173), .ZN(n1029) );
  NAND2_X1 U65 ( .A1(n976), .A2(n1204), .ZN(n984) );
  NAND2_X1 U66 ( .A1(n976), .A2(n1193), .ZN(n974) );
  NAND2_X1 U67 ( .A1(n976), .A2(n1183), .ZN(n965) );
  NAND2_X1 U68 ( .A1(n976), .A2(n1173), .ZN(n956) );
  NAND2_X1 U69 ( .A1(n1122), .A2(n1163), .ZN(n1093) );
  NAND2_X1 U70 ( .A1(n1122), .A2(n1153), .ZN(n1084) );
  NAND2_X1 U71 ( .A1(n1122), .A2(n1143), .ZN(n1075) );
  NAND2_X1 U72 ( .A1(n1122), .A2(n1133), .ZN(n1066) );
  NAND2_X1 U73 ( .A1(n1049), .A2(n1163), .ZN(n1020) );
  NAND2_X1 U74 ( .A1(n1049), .A2(n1153), .ZN(n1011) );
  NAND2_X1 U75 ( .A1(n1049), .A2(n1143), .ZN(n1002) );
  NAND2_X1 U76 ( .A1(n1049), .A2(n1133), .ZN(n993) );
  NAND2_X1 U77 ( .A1(n976), .A2(n1163), .ZN(n947) );
  NAND2_X1 U78 ( .A1(n976), .A2(n1153), .ZN(n938) );
  NAND2_X1 U79 ( .A1(n976), .A2(n1143), .ZN(n929) );
  NAND2_X1 U80 ( .A1(n976), .A2(n1133), .ZN(n920) );
  AND3_X1 U81 ( .A1(n847), .A2(n848), .A3(n1132), .ZN(n1203) );
  AND3_X1 U82 ( .A1(N13), .A2(n1132), .A3(N14), .ZN(n976) );
  AND3_X1 U83 ( .A1(n1132), .A2(n848), .A3(N13), .ZN(n1122) );
  AND3_X1 U84 ( .A1(n1132), .A2(n847), .A3(N14), .ZN(n1049) );
  NOR2_X1 U85 ( .A1(n846), .A2(addr[5]), .ZN(n1132) );
  INV_X1 U86 ( .A(wr_en), .ZN(n846) );
  OAI21_X1 U87 ( .B1(n622), .B2(n1172), .A(n1171), .ZN(n880) );
  NAND2_X1 U88 ( .A1(\mem[4][0] ), .A2(n1172), .ZN(n1171) );
  OAI21_X1 U89 ( .B1(n623), .B2(n1172), .A(n1170), .ZN(n879) );
  NAND2_X1 U90 ( .A1(\mem[4][1] ), .A2(n1172), .ZN(n1170) );
  OAI21_X1 U91 ( .B1(n624), .B2(n1172), .A(n1169), .ZN(n878) );
  NAND2_X1 U92 ( .A1(\mem[4][2] ), .A2(n1172), .ZN(n1169) );
  OAI21_X1 U93 ( .B1(n625), .B2(n1172), .A(n1168), .ZN(n877) );
  NAND2_X1 U94 ( .A1(\mem[4][3] ), .A2(n1172), .ZN(n1168) );
  OAI21_X1 U95 ( .B1(n626), .B2(n1172), .A(n1167), .ZN(n876) );
  NAND2_X1 U96 ( .A1(\mem[4][4] ), .A2(n1172), .ZN(n1167) );
  OAI21_X1 U97 ( .B1(n627), .B2(n1172), .A(n1166), .ZN(n875) );
  NAND2_X1 U98 ( .A1(\mem[4][5] ), .A2(n1172), .ZN(n1166) );
  OAI21_X1 U99 ( .B1(n628), .B2(n1172), .A(n1165), .ZN(n874) );
  NAND2_X1 U100 ( .A1(\mem[4][6] ), .A2(n1172), .ZN(n1165) );
  OAI21_X1 U101 ( .B1(n629), .B2(n1172), .A(n1164), .ZN(n873) );
  NAND2_X1 U102 ( .A1(\mem[4][7] ), .A2(n1172), .ZN(n1164) );
  OAI21_X1 U103 ( .B1(n622), .B2(n1152), .A(n1151), .ZN(n864) );
  NAND2_X1 U104 ( .A1(\mem[6][0] ), .A2(n1152), .ZN(n1151) );
  OAI21_X1 U105 ( .B1(n623), .B2(n1152), .A(n1150), .ZN(n863) );
  NAND2_X1 U106 ( .A1(\mem[6][1] ), .A2(n1152), .ZN(n1150) );
  OAI21_X1 U107 ( .B1(n624), .B2(n1152), .A(n1149), .ZN(n862) );
  NAND2_X1 U108 ( .A1(\mem[6][2] ), .A2(n1152), .ZN(n1149) );
  OAI21_X1 U109 ( .B1(n625), .B2(n1152), .A(n1148), .ZN(n861) );
  NAND2_X1 U110 ( .A1(\mem[6][3] ), .A2(n1152), .ZN(n1148) );
  OAI21_X1 U111 ( .B1(n626), .B2(n1152), .A(n1147), .ZN(n860) );
  NAND2_X1 U112 ( .A1(\mem[6][4] ), .A2(n1152), .ZN(n1147) );
  OAI21_X1 U113 ( .B1(n627), .B2(n1152), .A(n1146), .ZN(n859) );
  NAND2_X1 U114 ( .A1(\mem[6][5] ), .A2(n1152), .ZN(n1146) );
  OAI21_X1 U115 ( .B1(n628), .B2(n1152), .A(n1145), .ZN(n858) );
  NAND2_X1 U116 ( .A1(\mem[6][6] ), .A2(n1152), .ZN(n1145) );
  OAI21_X1 U117 ( .B1(n629), .B2(n1152), .A(n1144), .ZN(n857) );
  NAND2_X1 U118 ( .A1(\mem[6][7] ), .A2(n1152), .ZN(n1144) );
  OAI21_X1 U119 ( .B1(n622), .B2(n1142), .A(n1141), .ZN(n856) );
  NAND2_X1 U120 ( .A1(\mem[7][0] ), .A2(n1142), .ZN(n1141) );
  OAI21_X1 U121 ( .B1(n623), .B2(n1142), .A(n1140), .ZN(n855) );
  NAND2_X1 U122 ( .A1(\mem[7][1] ), .A2(n1142), .ZN(n1140) );
  OAI21_X1 U123 ( .B1(n624), .B2(n1142), .A(n1139), .ZN(n854) );
  NAND2_X1 U124 ( .A1(\mem[7][2] ), .A2(n1142), .ZN(n1139) );
  OAI21_X1 U125 ( .B1(n625), .B2(n1142), .A(n1138), .ZN(n853) );
  NAND2_X1 U126 ( .A1(\mem[7][3] ), .A2(n1142), .ZN(n1138) );
  OAI21_X1 U127 ( .B1(n626), .B2(n1142), .A(n1137), .ZN(n852) );
  NAND2_X1 U128 ( .A1(\mem[7][4] ), .A2(n1142), .ZN(n1137) );
  OAI21_X1 U129 ( .B1(n627), .B2(n1142), .A(n1136), .ZN(n851) );
  NAND2_X1 U130 ( .A1(\mem[7][5] ), .A2(n1142), .ZN(n1136) );
  OAI21_X1 U131 ( .B1(n628), .B2(n1142), .A(n1135), .ZN(n850) );
  NAND2_X1 U132 ( .A1(\mem[7][6] ), .A2(n1142), .ZN(n1135) );
  OAI21_X1 U133 ( .B1(n629), .B2(n1142), .A(n1134), .ZN(n849) );
  NAND2_X1 U134 ( .A1(\mem[7][7] ), .A2(n1142), .ZN(n1134) );
  OAI21_X1 U135 ( .B1(n622), .B2(n1202), .A(n1201), .ZN(n904) );
  NAND2_X1 U136 ( .A1(\mem[1][0] ), .A2(n1202), .ZN(n1201) );
  OAI21_X1 U137 ( .B1(n623), .B2(n1202), .A(n1200), .ZN(n903) );
  NAND2_X1 U138 ( .A1(\mem[1][1] ), .A2(n1202), .ZN(n1200) );
  OAI21_X1 U139 ( .B1(n624), .B2(n1202), .A(n1199), .ZN(n902) );
  NAND2_X1 U140 ( .A1(\mem[1][2] ), .A2(n1202), .ZN(n1199) );
  OAI21_X1 U141 ( .B1(n625), .B2(n1202), .A(n1198), .ZN(n901) );
  NAND2_X1 U142 ( .A1(\mem[1][3] ), .A2(n1202), .ZN(n1198) );
  OAI21_X1 U143 ( .B1(n626), .B2(n1202), .A(n1197), .ZN(n900) );
  NAND2_X1 U144 ( .A1(\mem[1][4] ), .A2(n1202), .ZN(n1197) );
  OAI21_X1 U145 ( .B1(n627), .B2(n1202), .A(n1196), .ZN(n899) );
  NAND2_X1 U146 ( .A1(\mem[1][5] ), .A2(n1202), .ZN(n1196) );
  OAI21_X1 U147 ( .B1(n628), .B2(n1202), .A(n1195), .ZN(n898) );
  NAND2_X1 U148 ( .A1(\mem[1][6] ), .A2(n1202), .ZN(n1195) );
  OAI21_X1 U149 ( .B1(n629), .B2(n1202), .A(n1194), .ZN(n897) );
  NAND2_X1 U150 ( .A1(\mem[1][7] ), .A2(n1202), .ZN(n1194) );
  OAI21_X1 U151 ( .B1(n622), .B2(n1192), .A(n1191), .ZN(n896) );
  NAND2_X1 U152 ( .A1(\mem[2][0] ), .A2(n1192), .ZN(n1191) );
  OAI21_X1 U153 ( .B1(n623), .B2(n1192), .A(n1190), .ZN(n895) );
  NAND2_X1 U154 ( .A1(\mem[2][1] ), .A2(n1192), .ZN(n1190) );
  OAI21_X1 U155 ( .B1(n624), .B2(n1192), .A(n1189), .ZN(n894) );
  NAND2_X1 U156 ( .A1(\mem[2][2] ), .A2(n1192), .ZN(n1189) );
  OAI21_X1 U157 ( .B1(n625), .B2(n1192), .A(n1188), .ZN(n893) );
  NAND2_X1 U158 ( .A1(\mem[2][3] ), .A2(n1192), .ZN(n1188) );
  OAI21_X1 U159 ( .B1(n626), .B2(n1192), .A(n1187), .ZN(n892) );
  NAND2_X1 U160 ( .A1(\mem[2][4] ), .A2(n1192), .ZN(n1187) );
  OAI21_X1 U161 ( .B1(n627), .B2(n1192), .A(n1186), .ZN(n891) );
  NAND2_X1 U162 ( .A1(\mem[2][5] ), .A2(n1192), .ZN(n1186) );
  OAI21_X1 U163 ( .B1(n628), .B2(n1192), .A(n1185), .ZN(n890) );
  NAND2_X1 U164 ( .A1(\mem[2][6] ), .A2(n1192), .ZN(n1185) );
  OAI21_X1 U165 ( .B1(n629), .B2(n1192), .A(n1184), .ZN(n889) );
  NAND2_X1 U166 ( .A1(\mem[2][7] ), .A2(n1192), .ZN(n1184) );
  OAI21_X1 U167 ( .B1(n622), .B2(n1182), .A(n1181), .ZN(n888) );
  NAND2_X1 U168 ( .A1(\mem[3][0] ), .A2(n1182), .ZN(n1181) );
  OAI21_X1 U169 ( .B1(n623), .B2(n1182), .A(n1180), .ZN(n887) );
  NAND2_X1 U170 ( .A1(\mem[3][1] ), .A2(n1182), .ZN(n1180) );
  OAI21_X1 U171 ( .B1(n624), .B2(n1182), .A(n1179), .ZN(n886) );
  NAND2_X1 U172 ( .A1(\mem[3][2] ), .A2(n1182), .ZN(n1179) );
  OAI21_X1 U173 ( .B1(n625), .B2(n1182), .A(n1178), .ZN(n885) );
  NAND2_X1 U174 ( .A1(\mem[3][3] ), .A2(n1182), .ZN(n1178) );
  OAI21_X1 U175 ( .B1(n626), .B2(n1182), .A(n1177), .ZN(n884) );
  NAND2_X1 U176 ( .A1(\mem[3][4] ), .A2(n1182), .ZN(n1177) );
  OAI21_X1 U177 ( .B1(n627), .B2(n1182), .A(n1176), .ZN(n883) );
  NAND2_X1 U178 ( .A1(\mem[3][5] ), .A2(n1182), .ZN(n1176) );
  OAI21_X1 U179 ( .B1(n628), .B2(n1182), .A(n1175), .ZN(n882) );
  NAND2_X1 U180 ( .A1(\mem[3][6] ), .A2(n1182), .ZN(n1175) );
  OAI21_X1 U181 ( .B1(n629), .B2(n1182), .A(n1174), .ZN(n881) );
  NAND2_X1 U182 ( .A1(\mem[3][7] ), .A2(n1182), .ZN(n1174) );
  OAI21_X1 U183 ( .B1(n622), .B2(n1162), .A(n1161), .ZN(n872) );
  NAND2_X1 U184 ( .A1(\mem[5][0] ), .A2(n1162), .ZN(n1161) );
  OAI21_X1 U185 ( .B1(n623), .B2(n1162), .A(n1160), .ZN(n871) );
  NAND2_X1 U186 ( .A1(\mem[5][1] ), .A2(n1162), .ZN(n1160) );
  OAI21_X1 U187 ( .B1(n624), .B2(n1162), .A(n1159), .ZN(n870) );
  NAND2_X1 U188 ( .A1(\mem[5][2] ), .A2(n1162), .ZN(n1159) );
  OAI21_X1 U189 ( .B1(n625), .B2(n1162), .A(n1158), .ZN(n869) );
  NAND2_X1 U190 ( .A1(\mem[5][3] ), .A2(n1162), .ZN(n1158) );
  OAI21_X1 U191 ( .B1(n626), .B2(n1162), .A(n1157), .ZN(n868) );
  NAND2_X1 U192 ( .A1(\mem[5][4] ), .A2(n1162), .ZN(n1157) );
  OAI21_X1 U193 ( .B1(n627), .B2(n1162), .A(n1156), .ZN(n867) );
  NAND2_X1 U194 ( .A1(\mem[5][5] ), .A2(n1162), .ZN(n1156) );
  OAI21_X1 U195 ( .B1(n628), .B2(n1162), .A(n1155), .ZN(n866) );
  NAND2_X1 U196 ( .A1(\mem[5][6] ), .A2(n1162), .ZN(n1155) );
  OAI21_X1 U197 ( .B1(n629), .B2(n1162), .A(n1154), .ZN(n865) );
  NAND2_X1 U198 ( .A1(\mem[5][7] ), .A2(n1162), .ZN(n1154) );
  OAI21_X1 U199 ( .B1(n1213), .B2(n622), .A(n1212), .ZN(n912) );
  NAND2_X1 U200 ( .A1(\mem[0][0] ), .A2(n1213), .ZN(n1212) );
  OAI21_X1 U201 ( .B1(n1213), .B2(n623), .A(n1211), .ZN(n911) );
  NAND2_X1 U202 ( .A1(\mem[0][1] ), .A2(n1213), .ZN(n1211) );
  OAI21_X1 U203 ( .B1(n1213), .B2(n624), .A(n1210), .ZN(n910) );
  NAND2_X1 U204 ( .A1(\mem[0][2] ), .A2(n1213), .ZN(n1210) );
  OAI21_X1 U205 ( .B1(n1213), .B2(n625), .A(n1209), .ZN(n909) );
  NAND2_X1 U206 ( .A1(\mem[0][3] ), .A2(n1213), .ZN(n1209) );
  OAI21_X1 U207 ( .B1(n1213), .B2(n626), .A(n1208), .ZN(n908) );
  NAND2_X1 U208 ( .A1(\mem[0][4] ), .A2(n1213), .ZN(n1208) );
  OAI21_X1 U209 ( .B1(n1213), .B2(n627), .A(n1207), .ZN(n907) );
  NAND2_X1 U210 ( .A1(\mem[0][5] ), .A2(n1213), .ZN(n1207) );
  OAI21_X1 U211 ( .B1(n1213), .B2(n628), .A(n1206), .ZN(n906) );
  NAND2_X1 U212 ( .A1(\mem[0][6] ), .A2(n1213), .ZN(n1206) );
  OAI21_X1 U213 ( .B1(n1213), .B2(n629), .A(n1205), .ZN(n905) );
  NAND2_X1 U214 ( .A1(\mem[0][7] ), .A2(n1213), .ZN(n1205) );
  INV_X1 U215 ( .A(n1131), .ZN(n821) );
  AOI22_X1 U216 ( .A1(data_in[0]), .A2(n845), .B1(n1130), .B2(\mem[8][0] ), 
        .ZN(n1131) );
  INV_X1 U217 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U218 ( .A1(data_in[1]), .A2(n845), .B1(n1130), .B2(\mem[8][1] ), 
        .ZN(n1129) );
  INV_X1 U219 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U220 ( .A1(data_in[2]), .A2(n845), .B1(n1130), .B2(\mem[8][2] ), 
        .ZN(n1128) );
  INV_X1 U221 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U222 ( .A1(data_in[3]), .A2(n845), .B1(n1130), .B2(\mem[8][3] ), 
        .ZN(n1127) );
  INV_X1 U223 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U224 ( .A1(data_in[4]), .A2(n845), .B1(n1130), .B2(\mem[8][4] ), 
        .ZN(n1126) );
  INV_X1 U225 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U226 ( .A1(data_in[5]), .A2(n845), .B1(n1130), .B2(\mem[8][5] ), 
        .ZN(n1125) );
  INV_X1 U227 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U228 ( .A1(data_in[6]), .A2(n845), .B1(n1130), .B2(\mem[8][6] ), 
        .ZN(n1124) );
  INV_X1 U229 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U230 ( .A1(data_in[7]), .A2(n845), .B1(n1130), .B2(\mem[8][7] ), 
        .ZN(n1123) );
  INV_X1 U231 ( .A(n1121), .ZN(n813) );
  AOI22_X1 U232 ( .A1(data_in[0]), .A2(n844), .B1(n1120), .B2(\mem[9][0] ), 
        .ZN(n1121) );
  INV_X1 U233 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U234 ( .A1(data_in[1]), .A2(n844), .B1(n1120), .B2(\mem[9][1] ), 
        .ZN(n1119) );
  INV_X1 U235 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U236 ( .A1(data_in[2]), .A2(n844), .B1(n1120), .B2(\mem[9][2] ), 
        .ZN(n1118) );
  INV_X1 U237 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U238 ( .A1(data_in[3]), .A2(n844), .B1(n1120), .B2(\mem[9][3] ), 
        .ZN(n1117) );
  INV_X1 U239 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U240 ( .A1(data_in[4]), .A2(n844), .B1(n1120), .B2(\mem[9][4] ), 
        .ZN(n1116) );
  INV_X1 U241 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U242 ( .A1(data_in[5]), .A2(n844), .B1(n1120), .B2(\mem[9][5] ), 
        .ZN(n1115) );
  INV_X1 U243 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U244 ( .A1(data_in[6]), .A2(n844), .B1(n1120), .B2(\mem[9][6] ), 
        .ZN(n1114) );
  INV_X1 U245 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U246 ( .A1(data_in[7]), .A2(n844), .B1(n1120), .B2(\mem[9][7] ), 
        .ZN(n1113) );
  INV_X1 U247 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U248 ( .A1(data_in[0]), .A2(n843), .B1(n1111), .B2(\mem[10][0] ), 
        .ZN(n1112) );
  INV_X1 U249 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U250 ( .A1(data_in[1]), .A2(n843), .B1(n1111), .B2(\mem[10][1] ), 
        .ZN(n1110) );
  INV_X1 U251 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U252 ( .A1(data_in[2]), .A2(n843), .B1(n1111), .B2(\mem[10][2] ), 
        .ZN(n1109) );
  INV_X1 U253 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U254 ( .A1(data_in[3]), .A2(n843), .B1(n1111), .B2(\mem[10][3] ), 
        .ZN(n1108) );
  INV_X1 U255 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U256 ( .A1(data_in[4]), .A2(n843), .B1(n1111), .B2(\mem[10][4] ), 
        .ZN(n1107) );
  INV_X1 U257 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U258 ( .A1(data_in[5]), .A2(n843), .B1(n1111), .B2(\mem[10][5] ), 
        .ZN(n1106) );
  INV_X1 U259 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U260 ( .A1(data_in[6]), .A2(n843), .B1(n1111), .B2(\mem[10][6] ), 
        .ZN(n1105) );
  INV_X1 U261 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U262 ( .A1(data_in[7]), .A2(n843), .B1(n1111), .B2(\mem[10][7] ), 
        .ZN(n1104) );
  INV_X1 U263 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U264 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[11][0] ), 
        .ZN(n1103) );
  INV_X1 U265 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U266 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[11][1] ), 
        .ZN(n1101) );
  INV_X1 U267 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U268 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[11][2] ), 
        .ZN(n1100) );
  INV_X1 U269 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U270 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[11][3] ), 
        .ZN(n1099) );
  INV_X1 U271 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U272 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[11][4] ), 
        .ZN(n1098) );
  INV_X1 U273 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U274 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[11][5] ), 
        .ZN(n1097) );
  INV_X1 U275 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U276 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[11][6] ), 
        .ZN(n1096) );
  INV_X1 U277 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U278 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[11][7] ), 
        .ZN(n1095) );
  INV_X1 U279 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U280 ( .A1(data_in[0]), .A2(n841), .B1(n1093), .B2(\mem[12][0] ), 
        .ZN(n1094) );
  INV_X1 U281 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U282 ( .A1(data_in[1]), .A2(n841), .B1(n1093), .B2(\mem[12][1] ), 
        .ZN(n1092) );
  INV_X1 U283 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U284 ( .A1(data_in[2]), .A2(n841), .B1(n1093), .B2(\mem[12][2] ), 
        .ZN(n1091) );
  INV_X1 U285 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U286 ( .A1(data_in[3]), .A2(n841), .B1(n1093), .B2(\mem[12][3] ), 
        .ZN(n1090) );
  INV_X1 U287 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U288 ( .A1(data_in[4]), .A2(n841), .B1(n1093), .B2(\mem[12][4] ), 
        .ZN(n1089) );
  INV_X1 U289 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U290 ( .A1(data_in[5]), .A2(n841), .B1(n1093), .B2(\mem[12][5] ), 
        .ZN(n1088) );
  INV_X1 U291 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U292 ( .A1(data_in[6]), .A2(n841), .B1(n1093), .B2(\mem[12][6] ), 
        .ZN(n1087) );
  INV_X1 U293 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U294 ( .A1(data_in[7]), .A2(n841), .B1(n1093), .B2(\mem[12][7] ), 
        .ZN(n1086) );
  INV_X1 U295 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U296 ( .A1(data_in[0]), .A2(n840), .B1(n1084), .B2(\mem[13][0] ), 
        .ZN(n1085) );
  INV_X1 U297 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U298 ( .A1(data_in[1]), .A2(n840), .B1(n1084), .B2(\mem[13][1] ), 
        .ZN(n1083) );
  INV_X1 U299 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U300 ( .A1(data_in[2]), .A2(n840), .B1(n1084), .B2(\mem[13][2] ), 
        .ZN(n1082) );
  INV_X1 U301 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U302 ( .A1(data_in[3]), .A2(n840), .B1(n1084), .B2(\mem[13][3] ), 
        .ZN(n1081) );
  INV_X1 U303 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U304 ( .A1(data_in[4]), .A2(n840), .B1(n1084), .B2(\mem[13][4] ), 
        .ZN(n1080) );
  INV_X1 U305 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U306 ( .A1(data_in[5]), .A2(n840), .B1(n1084), .B2(\mem[13][5] ), 
        .ZN(n1079) );
  INV_X1 U307 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U308 ( .A1(data_in[6]), .A2(n840), .B1(n1084), .B2(\mem[13][6] ), 
        .ZN(n1078) );
  INV_X1 U309 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U310 ( .A1(data_in[7]), .A2(n840), .B1(n1084), .B2(\mem[13][7] ), 
        .ZN(n1077) );
  INV_X1 U311 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U312 ( .A1(data_in[0]), .A2(n839), .B1(n1075), .B2(\mem[14][0] ), 
        .ZN(n1076) );
  INV_X1 U313 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U314 ( .A1(data_in[1]), .A2(n839), .B1(n1075), .B2(\mem[14][1] ), 
        .ZN(n1074) );
  INV_X1 U315 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U316 ( .A1(data_in[2]), .A2(n839), .B1(n1075), .B2(\mem[14][2] ), 
        .ZN(n1073) );
  INV_X1 U317 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U318 ( .A1(data_in[3]), .A2(n839), .B1(n1075), .B2(\mem[14][3] ), 
        .ZN(n1072) );
  INV_X1 U319 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U320 ( .A1(data_in[4]), .A2(n839), .B1(n1075), .B2(\mem[14][4] ), 
        .ZN(n1071) );
  INV_X1 U321 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U322 ( .A1(data_in[5]), .A2(n839), .B1(n1075), .B2(\mem[14][5] ), 
        .ZN(n1070) );
  INV_X1 U323 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U324 ( .A1(data_in[6]), .A2(n839), .B1(n1075), .B2(\mem[14][6] ), 
        .ZN(n1069) );
  INV_X1 U325 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U326 ( .A1(data_in[7]), .A2(n839), .B1(n1075), .B2(\mem[14][7] ), 
        .ZN(n1068) );
  INV_X1 U327 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U328 ( .A1(data_in[0]), .A2(n838), .B1(n1066), .B2(\mem[15][0] ), 
        .ZN(n1067) );
  INV_X1 U329 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U330 ( .A1(data_in[1]), .A2(n838), .B1(n1066), .B2(\mem[15][1] ), 
        .ZN(n1065) );
  INV_X1 U331 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U332 ( .A1(data_in[2]), .A2(n838), .B1(n1066), .B2(\mem[15][2] ), 
        .ZN(n1064) );
  INV_X1 U333 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U334 ( .A1(data_in[3]), .A2(n838), .B1(n1066), .B2(\mem[15][3] ), 
        .ZN(n1063) );
  INV_X1 U335 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U336 ( .A1(data_in[4]), .A2(n838), .B1(n1066), .B2(\mem[15][4] ), 
        .ZN(n1062) );
  INV_X1 U337 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U338 ( .A1(data_in[5]), .A2(n838), .B1(n1066), .B2(\mem[15][5] ), 
        .ZN(n1061) );
  INV_X1 U339 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U340 ( .A1(data_in[6]), .A2(n838), .B1(n1066), .B2(\mem[15][6] ), 
        .ZN(n1060) );
  INV_X1 U341 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U342 ( .A1(data_in[7]), .A2(n838), .B1(n1066), .B2(\mem[15][7] ), 
        .ZN(n1059) );
  INV_X1 U343 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U344 ( .A1(data_in[0]), .A2(n837), .B1(n1057), .B2(\mem[16][0] ), 
        .ZN(n1058) );
  INV_X1 U345 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U346 ( .A1(data_in[1]), .A2(n837), .B1(n1057), .B2(\mem[16][1] ), 
        .ZN(n1056) );
  INV_X1 U347 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U348 ( .A1(data_in[2]), .A2(n837), .B1(n1057), .B2(\mem[16][2] ), 
        .ZN(n1055) );
  INV_X1 U349 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U350 ( .A1(data_in[3]), .A2(n837), .B1(n1057), .B2(\mem[16][3] ), 
        .ZN(n1054) );
  INV_X1 U351 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U352 ( .A1(data_in[4]), .A2(n837), .B1(n1057), .B2(\mem[16][4] ), 
        .ZN(n1053) );
  INV_X1 U353 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U354 ( .A1(data_in[5]), .A2(n837), .B1(n1057), .B2(\mem[16][5] ), 
        .ZN(n1052) );
  INV_X1 U355 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U356 ( .A1(data_in[6]), .A2(n837), .B1(n1057), .B2(\mem[16][6] ), 
        .ZN(n1051) );
  INV_X1 U357 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U358 ( .A1(data_in[7]), .A2(n837), .B1(n1057), .B2(\mem[16][7] ), 
        .ZN(n1050) );
  INV_X1 U359 ( .A(n1048), .ZN(n749) );
  AOI22_X1 U360 ( .A1(data_in[0]), .A2(n836), .B1(n1047), .B2(\mem[17][0] ), 
        .ZN(n1048) );
  INV_X1 U361 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U362 ( .A1(data_in[1]), .A2(n836), .B1(n1047), .B2(\mem[17][1] ), 
        .ZN(n1046) );
  INV_X1 U363 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U364 ( .A1(data_in[2]), .A2(n836), .B1(n1047), .B2(\mem[17][2] ), 
        .ZN(n1045) );
  INV_X1 U365 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U366 ( .A1(data_in[3]), .A2(n836), .B1(n1047), .B2(\mem[17][3] ), 
        .ZN(n1044) );
  INV_X1 U367 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U368 ( .A1(data_in[4]), .A2(n836), .B1(n1047), .B2(\mem[17][4] ), 
        .ZN(n1043) );
  INV_X1 U369 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U370 ( .A1(data_in[5]), .A2(n836), .B1(n1047), .B2(\mem[17][5] ), 
        .ZN(n1042) );
  INV_X1 U371 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U372 ( .A1(data_in[6]), .A2(n836), .B1(n1047), .B2(\mem[17][6] ), 
        .ZN(n1041) );
  INV_X1 U373 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U374 ( .A1(data_in[7]), .A2(n836), .B1(n1047), .B2(\mem[17][7] ), 
        .ZN(n1040) );
  INV_X1 U375 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U376 ( .A1(data_in[0]), .A2(n835), .B1(n1038), .B2(\mem[18][0] ), 
        .ZN(n1039) );
  INV_X1 U377 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U378 ( .A1(data_in[1]), .A2(n835), .B1(n1038), .B2(\mem[18][1] ), 
        .ZN(n1037) );
  INV_X1 U379 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U380 ( .A1(data_in[2]), .A2(n835), .B1(n1038), .B2(\mem[18][2] ), 
        .ZN(n1036) );
  INV_X1 U381 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U382 ( .A1(data_in[3]), .A2(n835), .B1(n1038), .B2(\mem[18][3] ), 
        .ZN(n1035) );
  INV_X1 U383 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U384 ( .A1(data_in[4]), .A2(n835), .B1(n1038), .B2(\mem[18][4] ), 
        .ZN(n1034) );
  INV_X1 U385 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U386 ( .A1(data_in[5]), .A2(n835), .B1(n1038), .B2(\mem[18][5] ), 
        .ZN(n1033) );
  INV_X1 U387 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U388 ( .A1(data_in[6]), .A2(n835), .B1(n1038), .B2(\mem[18][6] ), 
        .ZN(n1032) );
  INV_X1 U389 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U390 ( .A1(data_in[7]), .A2(n835), .B1(n1038), .B2(\mem[18][7] ), 
        .ZN(n1031) );
  INV_X1 U391 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U392 ( .A1(data_in[0]), .A2(n834), .B1(n1029), .B2(\mem[19][0] ), 
        .ZN(n1030) );
  INV_X1 U393 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U394 ( .A1(data_in[1]), .A2(n834), .B1(n1029), .B2(\mem[19][1] ), 
        .ZN(n1028) );
  INV_X1 U395 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U396 ( .A1(data_in[2]), .A2(n834), .B1(n1029), .B2(\mem[19][2] ), 
        .ZN(n1027) );
  INV_X1 U397 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U398 ( .A1(data_in[3]), .A2(n834), .B1(n1029), .B2(\mem[19][3] ), 
        .ZN(n1026) );
  INV_X1 U399 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U400 ( .A1(data_in[4]), .A2(n834), .B1(n1029), .B2(\mem[19][4] ), 
        .ZN(n1025) );
  INV_X1 U401 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U402 ( .A1(data_in[5]), .A2(n834), .B1(n1029), .B2(\mem[19][5] ), 
        .ZN(n1024) );
  INV_X1 U403 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U404 ( .A1(data_in[6]), .A2(n834), .B1(n1029), .B2(\mem[19][6] ), 
        .ZN(n1023) );
  INV_X1 U405 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U406 ( .A1(data_in[7]), .A2(n834), .B1(n1029), .B2(\mem[19][7] ), 
        .ZN(n1022) );
  INV_X1 U407 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U408 ( .A1(data_in[0]), .A2(n833), .B1(n1020), .B2(\mem[20][0] ), 
        .ZN(n1021) );
  INV_X1 U409 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U410 ( .A1(data_in[1]), .A2(n833), .B1(n1020), .B2(\mem[20][1] ), 
        .ZN(n1019) );
  INV_X1 U411 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U412 ( .A1(data_in[2]), .A2(n833), .B1(n1020), .B2(\mem[20][2] ), 
        .ZN(n1018) );
  INV_X1 U413 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U414 ( .A1(data_in[3]), .A2(n833), .B1(n1020), .B2(\mem[20][3] ), 
        .ZN(n1017) );
  INV_X1 U415 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U416 ( .A1(data_in[4]), .A2(n833), .B1(n1020), .B2(\mem[20][4] ), 
        .ZN(n1016) );
  INV_X1 U417 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U418 ( .A1(data_in[5]), .A2(n833), .B1(n1020), .B2(\mem[20][5] ), 
        .ZN(n1015) );
  INV_X1 U419 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U420 ( .A1(data_in[6]), .A2(n833), .B1(n1020), .B2(\mem[20][6] ), 
        .ZN(n1014) );
  INV_X1 U421 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U422 ( .A1(data_in[7]), .A2(n833), .B1(n1020), .B2(\mem[20][7] ), 
        .ZN(n1013) );
  INV_X1 U423 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U424 ( .A1(data_in[0]), .A2(n832), .B1(n1011), .B2(\mem[21][0] ), 
        .ZN(n1012) );
  INV_X1 U425 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U426 ( .A1(data_in[1]), .A2(n832), .B1(n1011), .B2(\mem[21][1] ), 
        .ZN(n1010) );
  INV_X1 U427 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U428 ( .A1(data_in[2]), .A2(n832), .B1(n1011), .B2(\mem[21][2] ), 
        .ZN(n1009) );
  INV_X1 U429 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U430 ( .A1(data_in[3]), .A2(n832), .B1(n1011), .B2(\mem[21][3] ), 
        .ZN(n1008) );
  INV_X1 U431 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U432 ( .A1(data_in[4]), .A2(n832), .B1(n1011), .B2(\mem[21][4] ), 
        .ZN(n1007) );
  INV_X1 U433 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U434 ( .A1(data_in[5]), .A2(n832), .B1(n1011), .B2(\mem[21][5] ), 
        .ZN(n1006) );
  INV_X1 U435 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U436 ( .A1(data_in[6]), .A2(n832), .B1(n1011), .B2(\mem[21][6] ), 
        .ZN(n1005) );
  INV_X1 U437 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U438 ( .A1(data_in[7]), .A2(n832), .B1(n1011), .B2(\mem[21][7] ), 
        .ZN(n1004) );
  INV_X1 U439 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U440 ( .A1(data_in[0]), .A2(n831), .B1(n1002), .B2(\mem[22][0] ), 
        .ZN(n1003) );
  INV_X1 U441 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U442 ( .A1(data_in[1]), .A2(n831), .B1(n1002), .B2(\mem[22][1] ), 
        .ZN(n1001) );
  INV_X1 U443 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U444 ( .A1(data_in[2]), .A2(n831), .B1(n1002), .B2(\mem[22][2] ), 
        .ZN(n1000) );
  INV_X1 U445 ( .A(n999), .ZN(n706) );
  AOI22_X1 U446 ( .A1(data_in[3]), .A2(n831), .B1(n1002), .B2(\mem[22][3] ), 
        .ZN(n999) );
  INV_X1 U447 ( .A(n998), .ZN(n705) );
  AOI22_X1 U448 ( .A1(data_in[4]), .A2(n831), .B1(n1002), .B2(\mem[22][4] ), 
        .ZN(n998) );
  INV_X1 U449 ( .A(n997), .ZN(n704) );
  AOI22_X1 U450 ( .A1(data_in[5]), .A2(n831), .B1(n1002), .B2(\mem[22][5] ), 
        .ZN(n997) );
  INV_X1 U451 ( .A(n996), .ZN(n703) );
  AOI22_X1 U452 ( .A1(data_in[6]), .A2(n831), .B1(n1002), .B2(\mem[22][6] ), 
        .ZN(n996) );
  INV_X1 U453 ( .A(n995), .ZN(n702) );
  AOI22_X1 U454 ( .A1(data_in[7]), .A2(n831), .B1(n1002), .B2(\mem[22][7] ), 
        .ZN(n995) );
  INV_X1 U455 ( .A(n994), .ZN(n701) );
  AOI22_X1 U456 ( .A1(data_in[0]), .A2(n830), .B1(n993), .B2(\mem[23][0] ), 
        .ZN(n994) );
  INV_X1 U457 ( .A(n992), .ZN(n700) );
  AOI22_X1 U458 ( .A1(data_in[1]), .A2(n830), .B1(n993), .B2(\mem[23][1] ), 
        .ZN(n992) );
  INV_X1 U459 ( .A(n991), .ZN(n699) );
  AOI22_X1 U460 ( .A1(data_in[2]), .A2(n830), .B1(n993), .B2(\mem[23][2] ), 
        .ZN(n991) );
  INV_X1 U461 ( .A(n990), .ZN(n698) );
  AOI22_X1 U462 ( .A1(data_in[3]), .A2(n830), .B1(n993), .B2(\mem[23][3] ), 
        .ZN(n990) );
  INV_X1 U463 ( .A(n989), .ZN(n697) );
  AOI22_X1 U464 ( .A1(data_in[4]), .A2(n830), .B1(n993), .B2(\mem[23][4] ), 
        .ZN(n989) );
  INV_X1 U465 ( .A(n988), .ZN(n696) );
  AOI22_X1 U466 ( .A1(data_in[5]), .A2(n830), .B1(n993), .B2(\mem[23][5] ), 
        .ZN(n988) );
  INV_X1 U467 ( .A(n987), .ZN(n695) );
  AOI22_X1 U468 ( .A1(data_in[6]), .A2(n830), .B1(n993), .B2(\mem[23][6] ), 
        .ZN(n987) );
  INV_X1 U469 ( .A(n986), .ZN(n694) );
  AOI22_X1 U470 ( .A1(data_in[7]), .A2(n830), .B1(n993), .B2(\mem[23][7] ), 
        .ZN(n986) );
  INV_X1 U471 ( .A(n985), .ZN(n693) );
  AOI22_X1 U472 ( .A1(data_in[0]), .A2(n829), .B1(n984), .B2(\mem[24][0] ), 
        .ZN(n985) );
  INV_X1 U473 ( .A(n983), .ZN(n692) );
  AOI22_X1 U474 ( .A1(data_in[1]), .A2(n829), .B1(n984), .B2(\mem[24][1] ), 
        .ZN(n983) );
  INV_X1 U475 ( .A(n982), .ZN(n691) );
  AOI22_X1 U476 ( .A1(data_in[2]), .A2(n829), .B1(n984), .B2(\mem[24][2] ), 
        .ZN(n982) );
  INV_X1 U477 ( .A(n981), .ZN(n690) );
  AOI22_X1 U478 ( .A1(data_in[3]), .A2(n829), .B1(n984), .B2(\mem[24][3] ), 
        .ZN(n981) );
  INV_X1 U479 ( .A(n980), .ZN(n689) );
  AOI22_X1 U480 ( .A1(data_in[4]), .A2(n829), .B1(n984), .B2(\mem[24][4] ), 
        .ZN(n980) );
  INV_X1 U481 ( .A(n979), .ZN(n688) );
  AOI22_X1 U482 ( .A1(data_in[5]), .A2(n829), .B1(n984), .B2(\mem[24][5] ), 
        .ZN(n979) );
  INV_X1 U483 ( .A(n978), .ZN(n687) );
  AOI22_X1 U484 ( .A1(data_in[6]), .A2(n829), .B1(n984), .B2(\mem[24][6] ), 
        .ZN(n978) );
  INV_X1 U485 ( .A(n977), .ZN(n686) );
  AOI22_X1 U486 ( .A1(data_in[7]), .A2(n829), .B1(n984), .B2(\mem[24][7] ), 
        .ZN(n977) );
  INV_X1 U487 ( .A(n975), .ZN(n685) );
  AOI22_X1 U488 ( .A1(data_in[0]), .A2(n828), .B1(n974), .B2(\mem[25][0] ), 
        .ZN(n975) );
  INV_X1 U489 ( .A(n973), .ZN(n684) );
  AOI22_X1 U490 ( .A1(data_in[1]), .A2(n828), .B1(n974), .B2(\mem[25][1] ), 
        .ZN(n973) );
  INV_X1 U491 ( .A(n972), .ZN(n683) );
  AOI22_X1 U492 ( .A1(data_in[2]), .A2(n828), .B1(n974), .B2(\mem[25][2] ), 
        .ZN(n972) );
  INV_X1 U493 ( .A(n971), .ZN(n682) );
  AOI22_X1 U494 ( .A1(data_in[3]), .A2(n828), .B1(n974), .B2(\mem[25][3] ), 
        .ZN(n971) );
  INV_X1 U495 ( .A(n970), .ZN(n681) );
  AOI22_X1 U496 ( .A1(data_in[4]), .A2(n828), .B1(n974), .B2(\mem[25][4] ), 
        .ZN(n970) );
  INV_X1 U497 ( .A(n969), .ZN(n680) );
  AOI22_X1 U498 ( .A1(data_in[5]), .A2(n828), .B1(n974), .B2(\mem[25][5] ), 
        .ZN(n969) );
  INV_X1 U499 ( .A(n968), .ZN(n679) );
  AOI22_X1 U500 ( .A1(data_in[6]), .A2(n828), .B1(n974), .B2(\mem[25][6] ), 
        .ZN(n968) );
  INV_X1 U501 ( .A(n967), .ZN(n678) );
  AOI22_X1 U502 ( .A1(data_in[7]), .A2(n828), .B1(n974), .B2(\mem[25][7] ), 
        .ZN(n967) );
  INV_X1 U503 ( .A(n966), .ZN(n677) );
  AOI22_X1 U504 ( .A1(data_in[0]), .A2(n827), .B1(n965), .B2(\mem[26][0] ), 
        .ZN(n966) );
  INV_X1 U505 ( .A(n964), .ZN(n676) );
  AOI22_X1 U506 ( .A1(data_in[1]), .A2(n827), .B1(n965), .B2(\mem[26][1] ), 
        .ZN(n964) );
  INV_X1 U507 ( .A(n963), .ZN(n675) );
  AOI22_X1 U508 ( .A1(data_in[2]), .A2(n827), .B1(n965), .B2(\mem[26][2] ), 
        .ZN(n963) );
  INV_X1 U509 ( .A(n962), .ZN(n674) );
  AOI22_X1 U510 ( .A1(data_in[3]), .A2(n827), .B1(n965), .B2(\mem[26][3] ), 
        .ZN(n962) );
  INV_X1 U511 ( .A(n961), .ZN(n673) );
  AOI22_X1 U512 ( .A1(data_in[4]), .A2(n827), .B1(n965), .B2(\mem[26][4] ), 
        .ZN(n961) );
  INV_X1 U513 ( .A(n960), .ZN(n672) );
  AOI22_X1 U514 ( .A1(data_in[5]), .A2(n827), .B1(n965), .B2(\mem[26][5] ), 
        .ZN(n960) );
  INV_X1 U515 ( .A(n959), .ZN(n671) );
  AOI22_X1 U516 ( .A1(data_in[6]), .A2(n827), .B1(n965), .B2(\mem[26][6] ), 
        .ZN(n959) );
  INV_X1 U517 ( .A(n958), .ZN(n670) );
  AOI22_X1 U518 ( .A1(data_in[7]), .A2(n827), .B1(n965), .B2(\mem[26][7] ), 
        .ZN(n958) );
  INV_X1 U519 ( .A(n957), .ZN(n669) );
  AOI22_X1 U520 ( .A1(data_in[0]), .A2(n826), .B1(n956), .B2(\mem[27][0] ), 
        .ZN(n957) );
  INV_X1 U521 ( .A(n955), .ZN(n668) );
  AOI22_X1 U522 ( .A1(data_in[1]), .A2(n826), .B1(n956), .B2(\mem[27][1] ), 
        .ZN(n955) );
  INV_X1 U523 ( .A(n954), .ZN(n667) );
  AOI22_X1 U524 ( .A1(data_in[2]), .A2(n826), .B1(n956), .B2(\mem[27][2] ), 
        .ZN(n954) );
  INV_X1 U525 ( .A(n953), .ZN(n666) );
  AOI22_X1 U526 ( .A1(data_in[3]), .A2(n826), .B1(n956), .B2(\mem[27][3] ), 
        .ZN(n953) );
  INV_X1 U527 ( .A(n952), .ZN(n665) );
  AOI22_X1 U528 ( .A1(data_in[4]), .A2(n826), .B1(n956), .B2(\mem[27][4] ), 
        .ZN(n952) );
  INV_X1 U529 ( .A(n951), .ZN(n664) );
  AOI22_X1 U530 ( .A1(data_in[5]), .A2(n826), .B1(n956), .B2(\mem[27][5] ), 
        .ZN(n951) );
  INV_X1 U531 ( .A(n950), .ZN(n663) );
  AOI22_X1 U532 ( .A1(data_in[6]), .A2(n826), .B1(n956), .B2(\mem[27][6] ), 
        .ZN(n950) );
  INV_X1 U533 ( .A(n949), .ZN(n662) );
  AOI22_X1 U534 ( .A1(data_in[7]), .A2(n826), .B1(n956), .B2(\mem[27][7] ), 
        .ZN(n949) );
  INV_X1 U535 ( .A(n948), .ZN(n661) );
  AOI22_X1 U536 ( .A1(data_in[0]), .A2(n825), .B1(n947), .B2(\mem[28][0] ), 
        .ZN(n948) );
  INV_X1 U537 ( .A(n946), .ZN(n660) );
  AOI22_X1 U538 ( .A1(data_in[1]), .A2(n825), .B1(n947), .B2(\mem[28][1] ), 
        .ZN(n946) );
  INV_X1 U539 ( .A(n945), .ZN(n659) );
  AOI22_X1 U540 ( .A1(data_in[2]), .A2(n825), .B1(n947), .B2(\mem[28][2] ), 
        .ZN(n945) );
  INV_X1 U541 ( .A(n944), .ZN(n658) );
  AOI22_X1 U542 ( .A1(data_in[3]), .A2(n825), .B1(n947), .B2(\mem[28][3] ), 
        .ZN(n944) );
  INV_X1 U543 ( .A(n943), .ZN(n657) );
  AOI22_X1 U544 ( .A1(data_in[4]), .A2(n825), .B1(n947), .B2(\mem[28][4] ), 
        .ZN(n943) );
  INV_X1 U545 ( .A(n942), .ZN(n656) );
  AOI22_X1 U546 ( .A1(data_in[5]), .A2(n825), .B1(n947), .B2(\mem[28][5] ), 
        .ZN(n942) );
  INV_X1 U547 ( .A(n941), .ZN(n655) );
  AOI22_X1 U548 ( .A1(data_in[6]), .A2(n825), .B1(n947), .B2(\mem[28][6] ), 
        .ZN(n941) );
  INV_X1 U549 ( .A(n940), .ZN(n654) );
  AOI22_X1 U550 ( .A1(data_in[7]), .A2(n825), .B1(n947), .B2(\mem[28][7] ), 
        .ZN(n940) );
  INV_X1 U551 ( .A(n939), .ZN(n653) );
  AOI22_X1 U552 ( .A1(data_in[0]), .A2(n824), .B1(n938), .B2(\mem[29][0] ), 
        .ZN(n939) );
  INV_X1 U553 ( .A(n937), .ZN(n652) );
  AOI22_X1 U554 ( .A1(data_in[1]), .A2(n824), .B1(n938), .B2(\mem[29][1] ), 
        .ZN(n937) );
  INV_X1 U555 ( .A(n936), .ZN(n651) );
  AOI22_X1 U556 ( .A1(data_in[2]), .A2(n824), .B1(n938), .B2(\mem[29][2] ), 
        .ZN(n936) );
  INV_X1 U557 ( .A(n935), .ZN(n650) );
  AOI22_X1 U558 ( .A1(data_in[3]), .A2(n824), .B1(n938), .B2(\mem[29][3] ), 
        .ZN(n935) );
  INV_X1 U559 ( .A(n934), .ZN(n649) );
  AOI22_X1 U560 ( .A1(data_in[4]), .A2(n824), .B1(n938), .B2(\mem[29][4] ), 
        .ZN(n934) );
  INV_X1 U561 ( .A(n933), .ZN(n648) );
  AOI22_X1 U562 ( .A1(data_in[5]), .A2(n824), .B1(n938), .B2(\mem[29][5] ), 
        .ZN(n933) );
  INV_X1 U563 ( .A(n932), .ZN(n647) );
  AOI22_X1 U564 ( .A1(data_in[6]), .A2(n824), .B1(n938), .B2(\mem[29][6] ), 
        .ZN(n932) );
  INV_X1 U565 ( .A(n931), .ZN(n646) );
  AOI22_X1 U566 ( .A1(data_in[7]), .A2(n824), .B1(n938), .B2(\mem[29][7] ), 
        .ZN(n931) );
  INV_X1 U567 ( .A(n930), .ZN(n645) );
  AOI22_X1 U568 ( .A1(data_in[0]), .A2(n823), .B1(n929), .B2(\mem[30][0] ), 
        .ZN(n930) );
  INV_X1 U569 ( .A(n928), .ZN(n644) );
  AOI22_X1 U570 ( .A1(data_in[1]), .A2(n823), .B1(n929), .B2(\mem[30][1] ), 
        .ZN(n928) );
  INV_X1 U571 ( .A(n927), .ZN(n643) );
  AOI22_X1 U572 ( .A1(data_in[2]), .A2(n823), .B1(n929), .B2(\mem[30][2] ), 
        .ZN(n927) );
  INV_X1 U573 ( .A(n926), .ZN(n642) );
  AOI22_X1 U574 ( .A1(data_in[3]), .A2(n823), .B1(n929), .B2(\mem[30][3] ), 
        .ZN(n926) );
  INV_X1 U575 ( .A(n925), .ZN(n641) );
  AOI22_X1 U576 ( .A1(data_in[4]), .A2(n823), .B1(n929), .B2(\mem[30][4] ), 
        .ZN(n925) );
  INV_X1 U577 ( .A(n924), .ZN(n640) );
  AOI22_X1 U578 ( .A1(data_in[5]), .A2(n823), .B1(n929), .B2(\mem[30][5] ), 
        .ZN(n924) );
  INV_X1 U579 ( .A(n923), .ZN(n639) );
  AOI22_X1 U580 ( .A1(data_in[6]), .A2(n823), .B1(n929), .B2(\mem[30][6] ), 
        .ZN(n923) );
  INV_X1 U581 ( .A(n922), .ZN(n638) );
  AOI22_X1 U582 ( .A1(data_in[7]), .A2(n823), .B1(n929), .B2(\mem[30][7] ), 
        .ZN(n922) );
  INV_X1 U583 ( .A(n921), .ZN(n637) );
  AOI22_X1 U584 ( .A1(data_in[0]), .A2(n822), .B1(n920), .B2(\mem[31][0] ), 
        .ZN(n921) );
  INV_X1 U585 ( .A(n919), .ZN(n636) );
  AOI22_X1 U586 ( .A1(data_in[1]), .A2(n822), .B1(n920), .B2(\mem[31][1] ), 
        .ZN(n919) );
  INV_X1 U587 ( .A(n918), .ZN(n635) );
  AOI22_X1 U588 ( .A1(data_in[2]), .A2(n822), .B1(n920), .B2(\mem[31][2] ), 
        .ZN(n918) );
  INV_X1 U589 ( .A(n917), .ZN(n634) );
  AOI22_X1 U590 ( .A1(data_in[3]), .A2(n822), .B1(n920), .B2(\mem[31][3] ), 
        .ZN(n917) );
  INV_X1 U591 ( .A(n916), .ZN(n633) );
  AOI22_X1 U592 ( .A1(data_in[4]), .A2(n822), .B1(n920), .B2(\mem[31][4] ), 
        .ZN(n916) );
  INV_X1 U593 ( .A(n915), .ZN(n632) );
  AOI22_X1 U594 ( .A1(data_in[5]), .A2(n822), .B1(n920), .B2(\mem[31][5] ), 
        .ZN(n915) );
  INV_X1 U595 ( .A(n914), .ZN(n631) );
  AOI22_X1 U596 ( .A1(data_in[6]), .A2(n822), .B1(n920), .B2(\mem[31][6] ), 
        .ZN(n914) );
  INV_X1 U597 ( .A(n913), .ZN(n630) );
  AOI22_X1 U598 ( .A1(data_in[7]), .A2(n822), .B1(n920), .B2(\mem[31][7] ), 
        .ZN(n913) );
  MUX2_X1 U599 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n613), .Z(n3) );
  MUX2_X1 U600 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n613), .Z(n4) );
  MUX2_X1 U601 ( .A(n4), .B(n3), .S(n610), .Z(n5) );
  MUX2_X1 U602 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n613), .Z(n6) );
  MUX2_X1 U603 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n613), .Z(n7) );
  MUX2_X1 U604 ( .A(n7), .B(n6), .S(n610), .Z(n8) );
  MUX2_X1 U605 ( .A(n8), .B(n5), .S(n608), .Z(n9) );
  MUX2_X1 U606 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n613), .Z(n10) );
  MUX2_X1 U607 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n613), .Z(n11) );
  MUX2_X1 U608 ( .A(n11), .B(n10), .S(n610), .Z(n12) );
  MUX2_X1 U609 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n613), .Z(n13) );
  MUX2_X1 U610 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n613), .Z(n14) );
  MUX2_X1 U611 ( .A(n14), .B(n13), .S(n610), .Z(n15) );
  MUX2_X1 U612 ( .A(n15), .B(n12), .S(N12), .Z(n16) );
  MUX2_X1 U613 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U614 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n614), .Z(n18) );
  MUX2_X1 U615 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n614), .Z(n19) );
  MUX2_X1 U616 ( .A(n19), .B(n18), .S(n612), .Z(n20) );
  MUX2_X1 U617 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n614), .Z(n21) );
  MUX2_X1 U618 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n614), .Z(n22) );
  MUX2_X1 U619 ( .A(n22), .B(n21), .S(n612), .Z(n23) );
  MUX2_X1 U620 ( .A(n23), .B(n20), .S(N12), .Z(n24) );
  MUX2_X1 U621 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n614), .Z(n25) );
  MUX2_X1 U622 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n614), .Z(n26) );
  MUX2_X1 U623 ( .A(n26), .B(n25), .S(n611), .Z(n27) );
  MUX2_X1 U624 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n614), .Z(n28) );
  MUX2_X1 U625 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n614), .Z(n29) );
  MUX2_X1 U626 ( .A(n29), .B(n28), .S(n610), .Z(n30) );
  MUX2_X1 U627 ( .A(n30), .B(n27), .S(n609), .Z(n31) );
  MUX2_X1 U628 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U629 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U630 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n614), .Z(n33) );
  MUX2_X1 U631 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n614), .Z(n34) );
  MUX2_X1 U632 ( .A(n34), .B(n33), .S(n611), .Z(n35) );
  MUX2_X1 U633 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n614), .Z(n36) );
  MUX2_X1 U634 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n614), .Z(n37) );
  MUX2_X1 U635 ( .A(n37), .B(n36), .S(N11), .Z(n38) );
  MUX2_X1 U636 ( .A(n38), .B(n35), .S(n609), .Z(n39) );
  MUX2_X1 U637 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n615), .Z(n40) );
  MUX2_X1 U638 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n615), .Z(n41) );
  MUX2_X1 U639 ( .A(n41), .B(n40), .S(n610), .Z(n42) );
  MUX2_X1 U640 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n615), .Z(n43) );
  MUX2_X1 U641 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n615), .Z(n44) );
  MUX2_X1 U642 ( .A(n44), .B(n43), .S(n612), .Z(n45) );
  MUX2_X1 U643 ( .A(n45), .B(n42), .S(N12), .Z(n46) );
  MUX2_X1 U644 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U645 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n615), .Z(n48) );
  MUX2_X1 U646 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n615), .Z(n49) );
  MUX2_X1 U647 ( .A(n49), .B(n48), .S(n611), .Z(n50) );
  MUX2_X1 U648 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n615), .Z(n51) );
  MUX2_X1 U649 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n615), .Z(n52) );
  MUX2_X1 U650 ( .A(n52), .B(n51), .S(n611), .Z(n53) );
  MUX2_X1 U651 ( .A(n53), .B(n50), .S(n608), .Z(n54) );
  MUX2_X1 U652 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n615), .Z(n55) );
  MUX2_X1 U653 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n615), .Z(n56) );
  MUX2_X1 U654 ( .A(n56), .B(n55), .S(n610), .Z(n57) );
  MUX2_X1 U655 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n615), .Z(n58) );
  MUX2_X1 U656 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n615), .Z(n59) );
  MUX2_X1 U657 ( .A(n59), .B(n58), .S(n612), .Z(n60) );
  MUX2_X1 U658 ( .A(n60), .B(n57), .S(n608), .Z(n61) );
  MUX2_X1 U659 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U660 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U661 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n616), .Z(n63) );
  MUX2_X1 U662 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n616), .Z(n64) );
  MUX2_X1 U663 ( .A(n64), .B(n63), .S(n610), .Z(n65) );
  MUX2_X1 U664 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n616), .Z(n66) );
  MUX2_X1 U665 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n616), .Z(n67) );
  MUX2_X1 U666 ( .A(n67), .B(n66), .S(N11), .Z(n68) );
  MUX2_X1 U667 ( .A(n68), .B(n65), .S(n608), .Z(n69) );
  MUX2_X1 U668 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n616), .Z(n70) );
  MUX2_X1 U669 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n616), .Z(n71) );
  MUX2_X1 U670 ( .A(n71), .B(n70), .S(n610), .Z(n72) );
  MUX2_X1 U671 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n616), .Z(n73) );
  MUX2_X1 U672 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n616), .Z(n74) );
  MUX2_X1 U673 ( .A(n74), .B(n73), .S(N11), .Z(n75) );
  MUX2_X1 U674 ( .A(n75), .B(n72), .S(n608), .Z(n76) );
  MUX2_X1 U675 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U676 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n616), .Z(n78) );
  MUX2_X1 U677 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n616), .Z(n79) );
  MUX2_X1 U678 ( .A(n79), .B(n78), .S(n611), .Z(n80) );
  MUX2_X1 U679 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n616), .Z(n81) );
  MUX2_X1 U680 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n616), .Z(n82) );
  MUX2_X1 U681 ( .A(n82), .B(n81), .S(n611), .Z(n83) );
  MUX2_X1 U682 ( .A(n83), .B(n80), .S(n608), .Z(n84) );
  MUX2_X1 U683 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n617), .Z(n85) );
  MUX2_X1 U684 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n617), .Z(n86) );
  MUX2_X1 U685 ( .A(n86), .B(n85), .S(n612), .Z(n87) );
  MUX2_X1 U686 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n617), .Z(n88) );
  MUX2_X1 U687 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n617), .Z(n89) );
  MUX2_X1 U688 ( .A(n89), .B(n88), .S(n612), .Z(n90) );
  MUX2_X1 U689 ( .A(n90), .B(n87), .S(n608), .Z(n91) );
  MUX2_X1 U690 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U691 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U692 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n617), .Z(n93) );
  MUX2_X1 U693 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n617), .Z(n94) );
  MUX2_X1 U694 ( .A(n94), .B(n93), .S(n612), .Z(n95) );
  MUX2_X1 U695 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n617), .Z(n96) );
  MUX2_X1 U696 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n617), .Z(n97) );
  MUX2_X1 U697 ( .A(n97), .B(n96), .S(n612), .Z(n98) );
  MUX2_X1 U698 ( .A(n98), .B(n95), .S(n608), .Z(n99) );
  MUX2_X1 U699 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n617), .Z(n100) );
  MUX2_X1 U700 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n617), .Z(n101) );
  MUX2_X1 U701 ( .A(n101), .B(n100), .S(N11), .Z(n102) );
  MUX2_X1 U702 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n617), .Z(n103) );
  MUX2_X1 U703 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n617), .Z(n104) );
  MUX2_X1 U704 ( .A(n104), .B(n103), .S(N11), .Z(n105) );
  MUX2_X1 U705 ( .A(n105), .B(n102), .S(n608), .Z(n106) );
  MUX2_X1 U706 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U707 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n617), .Z(n108) );
  MUX2_X1 U708 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n617), .Z(n109) );
  MUX2_X1 U709 ( .A(n109), .B(n108), .S(n610), .Z(n110) );
  MUX2_X1 U710 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n615), .Z(n111) );
  MUX2_X1 U711 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n613), .Z(n112) );
  MUX2_X1 U712 ( .A(n112), .B(n111), .S(n612), .Z(n113) );
  MUX2_X1 U713 ( .A(n113), .B(n110), .S(n608), .Z(n114) );
  MUX2_X1 U714 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n615), .Z(n115) );
  MUX2_X1 U715 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n614), .Z(n116) );
  MUX2_X1 U716 ( .A(n116), .B(n115), .S(n610), .Z(n117) );
  MUX2_X1 U717 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n619), .Z(n118) );
  MUX2_X1 U718 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n119) );
  MUX2_X1 U719 ( .A(n119), .B(n118), .S(n611), .Z(n120) );
  MUX2_X1 U720 ( .A(n120), .B(n117), .S(n608), .Z(n121) );
  MUX2_X1 U721 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U722 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U723 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n615), .Z(n123) );
  MUX2_X1 U724 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n614), .Z(n124) );
  MUX2_X1 U725 ( .A(n124), .B(n123), .S(n610), .Z(n125) );
  MUX2_X1 U726 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n613), .Z(n126) );
  MUX2_X1 U727 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n613), .Z(n127) );
  MUX2_X1 U728 ( .A(n127), .B(n126), .S(n610), .Z(n128) );
  MUX2_X1 U729 ( .A(n128), .B(n125), .S(n608), .Z(n129) );
  MUX2_X1 U730 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n615), .Z(n130) );
  MUX2_X1 U731 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n615), .Z(n131) );
  MUX2_X1 U732 ( .A(n131), .B(n130), .S(n610), .Z(n132) );
  MUX2_X1 U733 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n617), .Z(n133) );
  MUX2_X1 U734 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n614), .Z(n134) );
  MUX2_X1 U735 ( .A(n134), .B(n133), .S(n611), .Z(n135) );
  MUX2_X1 U736 ( .A(n135), .B(n132), .S(n608), .Z(n136) );
  MUX2_X1 U737 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U738 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n614), .Z(n138) );
  MUX2_X1 U739 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n614), .Z(n139) );
  MUX2_X1 U740 ( .A(n139), .B(n138), .S(n610), .Z(n140) );
  MUX2_X1 U741 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n613), .Z(n141) );
  MUX2_X1 U742 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n614), .Z(n142) );
  MUX2_X1 U743 ( .A(n142), .B(n141), .S(n610), .Z(n143) );
  MUX2_X1 U744 ( .A(n143), .B(n140), .S(n608), .Z(n144) );
  MUX2_X1 U745 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n617), .Z(n145) );
  MUX2_X1 U746 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n615), .Z(n146) );
  MUX2_X1 U747 ( .A(n146), .B(n145), .S(n610), .Z(n147) );
  MUX2_X1 U748 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n617), .Z(n148) );
  MUX2_X1 U749 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n613), .Z(n149) );
  MUX2_X1 U750 ( .A(n149), .B(n148), .S(n610), .Z(n150) );
  MUX2_X1 U751 ( .A(n150), .B(n147), .S(n608), .Z(n151) );
  MUX2_X1 U752 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U753 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U754 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n613), .Z(n153) );
  MUX2_X1 U755 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n614), .Z(n154) );
  MUX2_X1 U756 ( .A(n154), .B(n153), .S(n611), .Z(n155) );
  MUX2_X1 U757 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n613), .Z(n156) );
  MUX2_X1 U758 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n614), .Z(n157) );
  MUX2_X1 U759 ( .A(n157), .B(n156), .S(n611), .Z(n158) );
  MUX2_X1 U760 ( .A(n158), .B(n155), .S(n609), .Z(n159) );
  MUX2_X1 U761 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n615), .Z(n160) );
  MUX2_X1 U762 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n615), .Z(n161) );
  MUX2_X1 U763 ( .A(n161), .B(n160), .S(n611), .Z(n162) );
  MUX2_X1 U764 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n613), .Z(n163) );
  MUX2_X1 U765 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n617), .Z(n164) );
  MUX2_X1 U766 ( .A(n164), .B(n163), .S(n611), .Z(n165) );
  MUX2_X1 U767 ( .A(n165), .B(n162), .S(n609), .Z(n166) );
  MUX2_X1 U768 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U769 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n613), .Z(n168) );
  MUX2_X1 U770 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n617), .Z(n169) );
  MUX2_X1 U771 ( .A(n169), .B(n168), .S(n611), .Z(n170) );
  MUX2_X1 U772 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n617), .Z(n171) );
  MUX2_X1 U773 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n613), .Z(n172) );
  MUX2_X1 U774 ( .A(n172), .B(n171), .S(n611), .Z(n173) );
  MUX2_X1 U775 ( .A(n173), .B(n170), .S(n609), .Z(n174) );
  MUX2_X1 U776 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n618), .Z(n175) );
  MUX2_X1 U777 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n618), .Z(n176) );
  MUX2_X1 U778 ( .A(n176), .B(n175), .S(n611), .Z(n177) );
  MUX2_X1 U779 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n618), .Z(n178) );
  MUX2_X1 U780 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n618), .Z(n179) );
  MUX2_X1 U781 ( .A(n179), .B(n178), .S(n611), .Z(n180) );
  MUX2_X1 U782 ( .A(n180), .B(n177), .S(n609), .Z(n181) );
  MUX2_X1 U783 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U784 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U785 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n618), .Z(n183) );
  MUX2_X1 U786 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n618), .Z(n184) );
  MUX2_X1 U787 ( .A(n184), .B(n183), .S(n611), .Z(n185) );
  MUX2_X1 U788 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n618), .Z(n186) );
  MUX2_X1 U789 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n618), .Z(n187) );
  MUX2_X1 U790 ( .A(n187), .B(n186), .S(n611), .Z(n188) );
  MUX2_X1 U791 ( .A(n188), .B(n185), .S(n609), .Z(n189) );
  MUX2_X1 U792 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n618), .Z(n190) );
  MUX2_X1 U793 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n618), .Z(n191) );
  MUX2_X1 U794 ( .A(n191), .B(n190), .S(n611), .Z(n192) );
  MUX2_X1 U795 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n618), .Z(n193) );
  MUX2_X1 U796 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n618), .Z(n194) );
  MUX2_X1 U797 ( .A(n194), .B(n193), .S(n611), .Z(n195) );
  MUX2_X1 U798 ( .A(n195), .B(n192), .S(n609), .Z(n196) );
  MUX2_X1 U799 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U800 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n617), .Z(n198) );
  MUX2_X1 U801 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n613), .Z(n199) );
  MUX2_X1 U802 ( .A(n199), .B(n198), .S(n612), .Z(n200) );
  MUX2_X1 U803 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n613), .Z(n201) );
  MUX2_X1 U804 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n613), .Z(n202) );
  MUX2_X1 U805 ( .A(n202), .B(n201), .S(n612), .Z(n203) );
  MUX2_X1 U806 ( .A(n203), .B(n200), .S(n609), .Z(n204) );
  MUX2_X1 U807 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n619), .Z(n205) );
  MUX2_X1 U808 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n619), .Z(n206) );
  MUX2_X1 U809 ( .A(n206), .B(n205), .S(n612), .Z(n207) );
  MUX2_X1 U810 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n619), .Z(n208) );
  MUX2_X1 U811 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n619), .Z(n209) );
  MUX2_X1 U812 ( .A(n209), .B(n208), .S(n612), .Z(n210) );
  MUX2_X1 U813 ( .A(n210), .B(n207), .S(n609), .Z(n211) );
  MUX2_X1 U814 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U815 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U816 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n619), .Z(n213) );
  MUX2_X1 U817 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n615), .Z(n214) );
  MUX2_X1 U818 ( .A(n214), .B(n213), .S(n612), .Z(n215) );
  MUX2_X1 U819 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n614), .Z(n216) );
  MUX2_X1 U820 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n619), .Z(n217) );
  MUX2_X1 U821 ( .A(n217), .B(n216), .S(n612), .Z(n218) );
  MUX2_X1 U822 ( .A(n218), .B(n215), .S(n609), .Z(n219) );
  MUX2_X1 U823 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n614), .Z(n220) );
  MUX2_X1 U824 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n617), .Z(n221) );
  MUX2_X1 U825 ( .A(n221), .B(n220), .S(n612), .Z(n222) );
  MUX2_X1 U826 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n613), .Z(n223) );
  MUX2_X1 U827 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n224) );
  MUX2_X1 U828 ( .A(n224), .B(n223), .S(n612), .Z(n225) );
  MUX2_X1 U829 ( .A(n225), .B(n222), .S(n609), .Z(n226) );
  MUX2_X1 U830 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U831 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n617), .Z(n228) );
  MUX2_X1 U832 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n619), .Z(n229) );
  MUX2_X1 U833 ( .A(n229), .B(n228), .S(n612), .Z(n595) );
  MUX2_X1 U834 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n615), .Z(n596) );
  MUX2_X1 U835 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n615), .Z(n597) );
  MUX2_X1 U836 ( .A(n597), .B(n596), .S(n612), .Z(n598) );
  MUX2_X1 U837 ( .A(n598), .B(n595), .S(n609), .Z(n599) );
  MUX2_X1 U838 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n619), .Z(n600) );
  MUX2_X1 U839 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n613), .Z(n601) );
  MUX2_X1 U840 ( .A(n601), .B(n600), .S(n612), .Z(n602) );
  MUX2_X1 U841 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n614), .Z(n603) );
  MUX2_X1 U842 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n604) );
  MUX2_X1 U843 ( .A(n604), .B(n603), .S(n612), .Z(n605) );
  MUX2_X1 U844 ( .A(n605), .B(n602), .S(n609), .Z(n606) );
  MUX2_X1 U845 ( .A(n606), .B(n599), .S(N13), .Z(n607) );
  MUX2_X1 U846 ( .A(n607), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U847 ( .A(N11), .Z(n610) );
  INV_X1 U848 ( .A(N10), .ZN(n620) );
  INV_X1 U849 ( .A(N11), .ZN(n621) );
  INV_X1 U850 ( .A(data_in[0]), .ZN(n622) );
  INV_X1 U851 ( .A(data_in[1]), .ZN(n623) );
  INV_X1 U852 ( .A(data_in[2]), .ZN(n624) );
  INV_X1 U853 ( .A(data_in[3]), .ZN(n625) );
  INV_X1 U854 ( .A(data_in[4]), .ZN(n626) );
  INV_X1 U855 ( .A(data_in[5]), .ZN(n627) );
  INV_X1 U856 ( .A(data_in[6]), .ZN(n628) );
  INV_X1 U857 ( .A(data_in[7]), .ZN(n629) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_4 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n630), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n631), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n632), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n633), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n634), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n635), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n636), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n637), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n638), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n639), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n640), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n641), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n642), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n643), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n644), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n645), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n646), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n647), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n648), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n649), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n650), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n651), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n652), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n653), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n654), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n655), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n656), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n657), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n658), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n659), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n660), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n661), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n662), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n663), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n664), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n665), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n666), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n667), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n668), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n669), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n670), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n671), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n672), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n673), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n674), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n675), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n676), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n677), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n678), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n679), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n680), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n681), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n682), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n683), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n684), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n685), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n686), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n687), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n688), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n689), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n690), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n691), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n692), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n693), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n694), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n695), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n696), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n697), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n698), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n699), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n700), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n701), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n702), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n703), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n704), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n705), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n706), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n707), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n708), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n709), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n710), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n711), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n712), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n713), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n714), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n715), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n716), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n717), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n718), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n719), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n720), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n721), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n722), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n723), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n724), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n725), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n726), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n727), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n728), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n729), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n730), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n731), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n732), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n733), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n734), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n735), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n736), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n737), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n738), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n739), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n740), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n741), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n742), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n743), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n744), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n745), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n746), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n747), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n748), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n749), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n750), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n751), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n752), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n753), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n754), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n755), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n756), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n757), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n758), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n759), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n760), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n761), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n762), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n763), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n764), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n765), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n766), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n767), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n768), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n769), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n770), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n771), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n772), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n773), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n774), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n775), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n776), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n777), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n778), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n779), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n780), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n781), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n782), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n783), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n784), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n785), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n786), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n787), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n788), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n789), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n790), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n791), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n792), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n793), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n794), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n795), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n796), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n797), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n798), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n799), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n800), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n801), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n802), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n803), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n804), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n805), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n806), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n807), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n808), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n809), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n810), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n811), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n812), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n813), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n814), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n815), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n816), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n817), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n818), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n819), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n820), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n821), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n849), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n850), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n851), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n852), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n853), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n854), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n855), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n856), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n857), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n858), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n859), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n860), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n861), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n862), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n863), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n864), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n865), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n866), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n867), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n868), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n869), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n870), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n871), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n872), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n873), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n874), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n875), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n876), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n877), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n878), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n879), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n880), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n881), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n882), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n883), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n884), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n885), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n886), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n887), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n888), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n889), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n890), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n891), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n892), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n893), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n894), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n895), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n896), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n897), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n898), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n899), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n900), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n901), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n902), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n903), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n904), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n905), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n906), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n907), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n908), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n909), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n910), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n911), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n912), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  BUF_X1 U3 ( .A(n619), .Z(n616) );
  BUF_X1 U4 ( .A(n619), .Z(n617) );
  BUF_X1 U5 ( .A(n619), .Z(n618) );
  BUF_X1 U6 ( .A(n619), .Z(n615) );
  BUF_X1 U7 ( .A(n619), .Z(n612) );
  BUF_X1 U8 ( .A(N10), .Z(n613) );
  BUF_X1 U9 ( .A(n619), .Z(n614) );
  BUF_X1 U10 ( .A(N11), .Z(n609) );
  BUF_X1 U11 ( .A(N11), .Z(n610) );
  BUF_X1 U12 ( .A(N10), .Z(n619) );
  NOR3_X1 U13 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1204) );
  NOR3_X1 U14 ( .A1(N11), .A2(N12), .A3(n620), .ZN(n1193) );
  NOR3_X1 U15 ( .A1(N10), .A2(N12), .A3(n621), .ZN(n1183) );
  NOR3_X1 U16 ( .A1(n620), .A2(N12), .A3(n621), .ZN(n1173) );
  INV_X1 U17 ( .A(n1130), .ZN(n845) );
  INV_X1 U18 ( .A(n1120), .ZN(n844) );
  INV_X1 U19 ( .A(n1111), .ZN(n843) );
  INV_X1 U20 ( .A(n1102), .ZN(n842) );
  INV_X1 U21 ( .A(n1057), .ZN(n837) );
  INV_X1 U22 ( .A(n1047), .ZN(n836) );
  INV_X1 U23 ( .A(n1038), .ZN(n835) );
  INV_X1 U24 ( .A(n1029), .ZN(n834) );
  INV_X1 U25 ( .A(n984), .ZN(n829) );
  INV_X1 U26 ( .A(n974), .ZN(n828) );
  INV_X1 U27 ( .A(n965), .ZN(n827) );
  INV_X1 U28 ( .A(n956), .ZN(n826) );
  INV_X1 U29 ( .A(n1093), .ZN(n841) );
  INV_X1 U30 ( .A(n1084), .ZN(n840) );
  INV_X1 U31 ( .A(n1075), .ZN(n839) );
  INV_X1 U32 ( .A(n1066), .ZN(n838) );
  INV_X1 U33 ( .A(n947), .ZN(n825) );
  INV_X1 U34 ( .A(n938), .ZN(n824) );
  INV_X1 U35 ( .A(n929), .ZN(n823) );
  INV_X1 U36 ( .A(n920), .ZN(n822) );
  INV_X1 U37 ( .A(n1020), .ZN(n833) );
  INV_X1 U38 ( .A(n1011), .ZN(n832) );
  INV_X1 U39 ( .A(n1002), .ZN(n831) );
  INV_X1 U40 ( .A(n993), .ZN(n830) );
  BUF_X1 U41 ( .A(N12), .Z(n607) );
  INV_X1 U42 ( .A(N13), .ZN(n847) );
  AND3_X1 U43 ( .A1(n620), .A2(n621), .A3(N12), .ZN(n1163) );
  AND3_X1 U44 ( .A1(N10), .A2(n621), .A3(N12), .ZN(n1153) );
  AND3_X1 U45 ( .A1(N11), .A2(n620), .A3(N12), .ZN(n1143) );
  AND3_X1 U46 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1133) );
  BUF_X1 U47 ( .A(N12), .Z(n606) );
  INV_X1 U48 ( .A(N14), .ZN(n848) );
  NAND2_X1 U49 ( .A1(n1193), .A2(n1203), .ZN(n1202) );
  NAND2_X1 U50 ( .A1(n1183), .A2(n1203), .ZN(n1192) );
  NAND2_X1 U51 ( .A1(n1173), .A2(n1203), .ZN(n1182) );
  NAND2_X1 U52 ( .A1(n1163), .A2(n1203), .ZN(n1172) );
  NAND2_X1 U53 ( .A1(n1153), .A2(n1203), .ZN(n1162) );
  NAND2_X1 U54 ( .A1(n1143), .A2(n1203), .ZN(n1152) );
  NAND2_X1 U55 ( .A1(n1133), .A2(n1203), .ZN(n1142) );
  NAND2_X1 U56 ( .A1(n1204), .A2(n1203), .ZN(n1213) );
  NAND2_X1 U57 ( .A1(n1122), .A2(n1204), .ZN(n1130) );
  NAND2_X1 U58 ( .A1(n1122), .A2(n1193), .ZN(n1120) );
  NAND2_X1 U59 ( .A1(n1122), .A2(n1183), .ZN(n1111) );
  NAND2_X1 U60 ( .A1(n1122), .A2(n1173), .ZN(n1102) );
  NAND2_X1 U61 ( .A1(n1049), .A2(n1204), .ZN(n1057) );
  NAND2_X1 U62 ( .A1(n1049), .A2(n1193), .ZN(n1047) );
  NAND2_X1 U63 ( .A1(n1049), .A2(n1183), .ZN(n1038) );
  NAND2_X1 U64 ( .A1(n1049), .A2(n1173), .ZN(n1029) );
  NAND2_X1 U65 ( .A1(n976), .A2(n1204), .ZN(n984) );
  NAND2_X1 U66 ( .A1(n976), .A2(n1193), .ZN(n974) );
  NAND2_X1 U67 ( .A1(n976), .A2(n1183), .ZN(n965) );
  NAND2_X1 U68 ( .A1(n976), .A2(n1173), .ZN(n956) );
  NAND2_X1 U69 ( .A1(n1122), .A2(n1163), .ZN(n1093) );
  NAND2_X1 U70 ( .A1(n1122), .A2(n1153), .ZN(n1084) );
  NAND2_X1 U71 ( .A1(n1122), .A2(n1143), .ZN(n1075) );
  NAND2_X1 U72 ( .A1(n1122), .A2(n1133), .ZN(n1066) );
  NAND2_X1 U73 ( .A1(n1049), .A2(n1163), .ZN(n1020) );
  NAND2_X1 U74 ( .A1(n1049), .A2(n1153), .ZN(n1011) );
  NAND2_X1 U75 ( .A1(n1049), .A2(n1143), .ZN(n1002) );
  NAND2_X1 U76 ( .A1(n1049), .A2(n1133), .ZN(n993) );
  NAND2_X1 U77 ( .A1(n976), .A2(n1163), .ZN(n947) );
  NAND2_X1 U78 ( .A1(n976), .A2(n1153), .ZN(n938) );
  NAND2_X1 U79 ( .A1(n976), .A2(n1143), .ZN(n929) );
  NAND2_X1 U80 ( .A1(n976), .A2(n1133), .ZN(n920) );
  AND3_X1 U81 ( .A1(n847), .A2(n848), .A3(n1132), .ZN(n1203) );
  AND3_X1 U82 ( .A1(N13), .A2(n1132), .A3(N14), .ZN(n976) );
  AND3_X1 U83 ( .A1(n1132), .A2(n848), .A3(N13), .ZN(n1122) );
  AND3_X1 U84 ( .A1(n1132), .A2(n847), .A3(N14), .ZN(n1049) );
  NOR2_X1 U85 ( .A1(n846), .A2(addr[5]), .ZN(n1132) );
  INV_X1 U86 ( .A(wr_en), .ZN(n846) );
  OAI21_X1 U87 ( .B1(n622), .B2(n1172), .A(n1171), .ZN(n880) );
  NAND2_X1 U88 ( .A1(\mem[4][0] ), .A2(n1172), .ZN(n1171) );
  OAI21_X1 U89 ( .B1(n623), .B2(n1172), .A(n1170), .ZN(n879) );
  NAND2_X1 U90 ( .A1(\mem[4][1] ), .A2(n1172), .ZN(n1170) );
  OAI21_X1 U91 ( .B1(n624), .B2(n1172), .A(n1169), .ZN(n878) );
  NAND2_X1 U92 ( .A1(\mem[4][2] ), .A2(n1172), .ZN(n1169) );
  OAI21_X1 U93 ( .B1(n625), .B2(n1172), .A(n1168), .ZN(n877) );
  NAND2_X1 U94 ( .A1(\mem[4][3] ), .A2(n1172), .ZN(n1168) );
  OAI21_X1 U95 ( .B1(n626), .B2(n1172), .A(n1167), .ZN(n876) );
  NAND2_X1 U96 ( .A1(\mem[4][4] ), .A2(n1172), .ZN(n1167) );
  OAI21_X1 U97 ( .B1(n627), .B2(n1172), .A(n1166), .ZN(n875) );
  NAND2_X1 U98 ( .A1(\mem[4][5] ), .A2(n1172), .ZN(n1166) );
  OAI21_X1 U99 ( .B1(n628), .B2(n1172), .A(n1165), .ZN(n874) );
  NAND2_X1 U100 ( .A1(\mem[4][6] ), .A2(n1172), .ZN(n1165) );
  OAI21_X1 U101 ( .B1(n629), .B2(n1172), .A(n1164), .ZN(n873) );
  NAND2_X1 U102 ( .A1(\mem[4][7] ), .A2(n1172), .ZN(n1164) );
  OAI21_X1 U103 ( .B1(n622), .B2(n1152), .A(n1151), .ZN(n864) );
  NAND2_X1 U104 ( .A1(\mem[6][0] ), .A2(n1152), .ZN(n1151) );
  OAI21_X1 U105 ( .B1(n623), .B2(n1152), .A(n1150), .ZN(n863) );
  NAND2_X1 U106 ( .A1(\mem[6][1] ), .A2(n1152), .ZN(n1150) );
  OAI21_X1 U107 ( .B1(n624), .B2(n1152), .A(n1149), .ZN(n862) );
  NAND2_X1 U108 ( .A1(\mem[6][2] ), .A2(n1152), .ZN(n1149) );
  OAI21_X1 U109 ( .B1(n625), .B2(n1152), .A(n1148), .ZN(n861) );
  NAND2_X1 U110 ( .A1(\mem[6][3] ), .A2(n1152), .ZN(n1148) );
  OAI21_X1 U111 ( .B1(n626), .B2(n1152), .A(n1147), .ZN(n860) );
  NAND2_X1 U112 ( .A1(\mem[6][4] ), .A2(n1152), .ZN(n1147) );
  OAI21_X1 U113 ( .B1(n627), .B2(n1152), .A(n1146), .ZN(n859) );
  NAND2_X1 U114 ( .A1(\mem[6][5] ), .A2(n1152), .ZN(n1146) );
  OAI21_X1 U115 ( .B1(n628), .B2(n1152), .A(n1145), .ZN(n858) );
  NAND2_X1 U116 ( .A1(\mem[6][6] ), .A2(n1152), .ZN(n1145) );
  OAI21_X1 U117 ( .B1(n629), .B2(n1152), .A(n1144), .ZN(n857) );
  NAND2_X1 U118 ( .A1(\mem[6][7] ), .A2(n1152), .ZN(n1144) );
  OAI21_X1 U119 ( .B1(n622), .B2(n1142), .A(n1141), .ZN(n856) );
  NAND2_X1 U120 ( .A1(\mem[7][0] ), .A2(n1142), .ZN(n1141) );
  OAI21_X1 U121 ( .B1(n623), .B2(n1142), .A(n1140), .ZN(n855) );
  NAND2_X1 U122 ( .A1(\mem[7][1] ), .A2(n1142), .ZN(n1140) );
  OAI21_X1 U123 ( .B1(n624), .B2(n1142), .A(n1139), .ZN(n854) );
  NAND2_X1 U124 ( .A1(\mem[7][2] ), .A2(n1142), .ZN(n1139) );
  OAI21_X1 U125 ( .B1(n625), .B2(n1142), .A(n1138), .ZN(n853) );
  NAND2_X1 U126 ( .A1(\mem[7][3] ), .A2(n1142), .ZN(n1138) );
  OAI21_X1 U127 ( .B1(n626), .B2(n1142), .A(n1137), .ZN(n852) );
  NAND2_X1 U128 ( .A1(\mem[7][4] ), .A2(n1142), .ZN(n1137) );
  OAI21_X1 U129 ( .B1(n627), .B2(n1142), .A(n1136), .ZN(n851) );
  NAND2_X1 U130 ( .A1(\mem[7][5] ), .A2(n1142), .ZN(n1136) );
  OAI21_X1 U131 ( .B1(n628), .B2(n1142), .A(n1135), .ZN(n850) );
  NAND2_X1 U132 ( .A1(\mem[7][6] ), .A2(n1142), .ZN(n1135) );
  OAI21_X1 U133 ( .B1(n629), .B2(n1142), .A(n1134), .ZN(n849) );
  NAND2_X1 U134 ( .A1(\mem[7][7] ), .A2(n1142), .ZN(n1134) );
  OAI21_X1 U135 ( .B1(n622), .B2(n1202), .A(n1201), .ZN(n904) );
  NAND2_X1 U136 ( .A1(\mem[1][0] ), .A2(n1202), .ZN(n1201) );
  OAI21_X1 U137 ( .B1(n623), .B2(n1202), .A(n1200), .ZN(n903) );
  NAND2_X1 U138 ( .A1(\mem[1][1] ), .A2(n1202), .ZN(n1200) );
  OAI21_X1 U139 ( .B1(n624), .B2(n1202), .A(n1199), .ZN(n902) );
  NAND2_X1 U140 ( .A1(\mem[1][2] ), .A2(n1202), .ZN(n1199) );
  OAI21_X1 U141 ( .B1(n625), .B2(n1202), .A(n1198), .ZN(n901) );
  NAND2_X1 U142 ( .A1(\mem[1][3] ), .A2(n1202), .ZN(n1198) );
  OAI21_X1 U143 ( .B1(n626), .B2(n1202), .A(n1197), .ZN(n900) );
  NAND2_X1 U144 ( .A1(\mem[1][4] ), .A2(n1202), .ZN(n1197) );
  OAI21_X1 U145 ( .B1(n627), .B2(n1202), .A(n1196), .ZN(n899) );
  NAND2_X1 U146 ( .A1(\mem[1][5] ), .A2(n1202), .ZN(n1196) );
  OAI21_X1 U147 ( .B1(n628), .B2(n1202), .A(n1195), .ZN(n898) );
  NAND2_X1 U148 ( .A1(\mem[1][6] ), .A2(n1202), .ZN(n1195) );
  OAI21_X1 U149 ( .B1(n629), .B2(n1202), .A(n1194), .ZN(n897) );
  NAND2_X1 U150 ( .A1(\mem[1][7] ), .A2(n1202), .ZN(n1194) );
  OAI21_X1 U151 ( .B1(n622), .B2(n1192), .A(n1191), .ZN(n896) );
  NAND2_X1 U152 ( .A1(\mem[2][0] ), .A2(n1192), .ZN(n1191) );
  OAI21_X1 U153 ( .B1(n623), .B2(n1192), .A(n1190), .ZN(n895) );
  NAND2_X1 U154 ( .A1(\mem[2][1] ), .A2(n1192), .ZN(n1190) );
  OAI21_X1 U155 ( .B1(n624), .B2(n1192), .A(n1189), .ZN(n894) );
  NAND2_X1 U156 ( .A1(\mem[2][2] ), .A2(n1192), .ZN(n1189) );
  OAI21_X1 U157 ( .B1(n625), .B2(n1192), .A(n1188), .ZN(n893) );
  NAND2_X1 U158 ( .A1(\mem[2][3] ), .A2(n1192), .ZN(n1188) );
  OAI21_X1 U159 ( .B1(n626), .B2(n1192), .A(n1187), .ZN(n892) );
  NAND2_X1 U160 ( .A1(\mem[2][4] ), .A2(n1192), .ZN(n1187) );
  OAI21_X1 U161 ( .B1(n627), .B2(n1192), .A(n1186), .ZN(n891) );
  NAND2_X1 U162 ( .A1(\mem[2][5] ), .A2(n1192), .ZN(n1186) );
  OAI21_X1 U163 ( .B1(n628), .B2(n1192), .A(n1185), .ZN(n890) );
  NAND2_X1 U164 ( .A1(\mem[2][6] ), .A2(n1192), .ZN(n1185) );
  OAI21_X1 U165 ( .B1(n629), .B2(n1192), .A(n1184), .ZN(n889) );
  NAND2_X1 U166 ( .A1(\mem[2][7] ), .A2(n1192), .ZN(n1184) );
  OAI21_X1 U167 ( .B1(n622), .B2(n1182), .A(n1181), .ZN(n888) );
  NAND2_X1 U168 ( .A1(\mem[3][0] ), .A2(n1182), .ZN(n1181) );
  OAI21_X1 U169 ( .B1(n623), .B2(n1182), .A(n1180), .ZN(n887) );
  NAND2_X1 U170 ( .A1(\mem[3][1] ), .A2(n1182), .ZN(n1180) );
  OAI21_X1 U171 ( .B1(n624), .B2(n1182), .A(n1179), .ZN(n886) );
  NAND2_X1 U172 ( .A1(\mem[3][2] ), .A2(n1182), .ZN(n1179) );
  OAI21_X1 U173 ( .B1(n625), .B2(n1182), .A(n1178), .ZN(n885) );
  NAND2_X1 U174 ( .A1(\mem[3][3] ), .A2(n1182), .ZN(n1178) );
  OAI21_X1 U175 ( .B1(n626), .B2(n1182), .A(n1177), .ZN(n884) );
  NAND2_X1 U176 ( .A1(\mem[3][4] ), .A2(n1182), .ZN(n1177) );
  OAI21_X1 U177 ( .B1(n627), .B2(n1182), .A(n1176), .ZN(n883) );
  NAND2_X1 U178 ( .A1(\mem[3][5] ), .A2(n1182), .ZN(n1176) );
  OAI21_X1 U179 ( .B1(n628), .B2(n1182), .A(n1175), .ZN(n882) );
  NAND2_X1 U180 ( .A1(\mem[3][6] ), .A2(n1182), .ZN(n1175) );
  OAI21_X1 U181 ( .B1(n629), .B2(n1182), .A(n1174), .ZN(n881) );
  NAND2_X1 U182 ( .A1(\mem[3][7] ), .A2(n1182), .ZN(n1174) );
  OAI21_X1 U183 ( .B1(n622), .B2(n1162), .A(n1161), .ZN(n872) );
  NAND2_X1 U184 ( .A1(\mem[5][0] ), .A2(n1162), .ZN(n1161) );
  OAI21_X1 U185 ( .B1(n623), .B2(n1162), .A(n1160), .ZN(n871) );
  NAND2_X1 U186 ( .A1(\mem[5][1] ), .A2(n1162), .ZN(n1160) );
  OAI21_X1 U187 ( .B1(n624), .B2(n1162), .A(n1159), .ZN(n870) );
  NAND2_X1 U188 ( .A1(\mem[5][2] ), .A2(n1162), .ZN(n1159) );
  OAI21_X1 U189 ( .B1(n625), .B2(n1162), .A(n1158), .ZN(n869) );
  NAND2_X1 U190 ( .A1(\mem[5][3] ), .A2(n1162), .ZN(n1158) );
  OAI21_X1 U191 ( .B1(n626), .B2(n1162), .A(n1157), .ZN(n868) );
  NAND2_X1 U192 ( .A1(\mem[5][4] ), .A2(n1162), .ZN(n1157) );
  OAI21_X1 U193 ( .B1(n627), .B2(n1162), .A(n1156), .ZN(n867) );
  NAND2_X1 U194 ( .A1(\mem[5][5] ), .A2(n1162), .ZN(n1156) );
  OAI21_X1 U195 ( .B1(n628), .B2(n1162), .A(n1155), .ZN(n866) );
  NAND2_X1 U196 ( .A1(\mem[5][6] ), .A2(n1162), .ZN(n1155) );
  OAI21_X1 U197 ( .B1(n629), .B2(n1162), .A(n1154), .ZN(n865) );
  NAND2_X1 U198 ( .A1(\mem[5][7] ), .A2(n1162), .ZN(n1154) );
  OAI21_X1 U199 ( .B1(n1213), .B2(n622), .A(n1212), .ZN(n912) );
  NAND2_X1 U200 ( .A1(\mem[0][0] ), .A2(n1213), .ZN(n1212) );
  OAI21_X1 U201 ( .B1(n1213), .B2(n623), .A(n1211), .ZN(n911) );
  NAND2_X1 U202 ( .A1(\mem[0][1] ), .A2(n1213), .ZN(n1211) );
  OAI21_X1 U203 ( .B1(n1213), .B2(n624), .A(n1210), .ZN(n910) );
  NAND2_X1 U204 ( .A1(\mem[0][2] ), .A2(n1213), .ZN(n1210) );
  OAI21_X1 U205 ( .B1(n1213), .B2(n625), .A(n1209), .ZN(n909) );
  NAND2_X1 U206 ( .A1(\mem[0][3] ), .A2(n1213), .ZN(n1209) );
  OAI21_X1 U207 ( .B1(n1213), .B2(n626), .A(n1208), .ZN(n908) );
  NAND2_X1 U208 ( .A1(\mem[0][4] ), .A2(n1213), .ZN(n1208) );
  OAI21_X1 U209 ( .B1(n1213), .B2(n627), .A(n1207), .ZN(n907) );
  NAND2_X1 U210 ( .A1(\mem[0][5] ), .A2(n1213), .ZN(n1207) );
  OAI21_X1 U211 ( .B1(n1213), .B2(n628), .A(n1206), .ZN(n906) );
  NAND2_X1 U212 ( .A1(\mem[0][6] ), .A2(n1213), .ZN(n1206) );
  OAI21_X1 U213 ( .B1(n1213), .B2(n629), .A(n1205), .ZN(n905) );
  NAND2_X1 U214 ( .A1(\mem[0][7] ), .A2(n1213), .ZN(n1205) );
  INV_X1 U215 ( .A(n1131), .ZN(n821) );
  AOI22_X1 U216 ( .A1(data_in[0]), .A2(n845), .B1(n1130), .B2(\mem[8][0] ), 
        .ZN(n1131) );
  INV_X1 U217 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U218 ( .A1(data_in[1]), .A2(n845), .B1(n1130), .B2(\mem[8][1] ), 
        .ZN(n1129) );
  INV_X1 U219 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U220 ( .A1(data_in[2]), .A2(n845), .B1(n1130), .B2(\mem[8][2] ), 
        .ZN(n1128) );
  INV_X1 U221 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U222 ( .A1(data_in[3]), .A2(n845), .B1(n1130), .B2(\mem[8][3] ), 
        .ZN(n1127) );
  INV_X1 U223 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U224 ( .A1(data_in[4]), .A2(n845), .B1(n1130), .B2(\mem[8][4] ), 
        .ZN(n1126) );
  INV_X1 U225 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U226 ( .A1(data_in[5]), .A2(n845), .B1(n1130), .B2(\mem[8][5] ), 
        .ZN(n1125) );
  INV_X1 U227 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U228 ( .A1(data_in[6]), .A2(n845), .B1(n1130), .B2(\mem[8][6] ), 
        .ZN(n1124) );
  INV_X1 U229 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U230 ( .A1(data_in[7]), .A2(n845), .B1(n1130), .B2(\mem[8][7] ), 
        .ZN(n1123) );
  INV_X1 U231 ( .A(n1121), .ZN(n813) );
  AOI22_X1 U232 ( .A1(data_in[0]), .A2(n844), .B1(n1120), .B2(\mem[9][0] ), 
        .ZN(n1121) );
  INV_X1 U233 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U234 ( .A1(data_in[1]), .A2(n844), .B1(n1120), .B2(\mem[9][1] ), 
        .ZN(n1119) );
  INV_X1 U235 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U236 ( .A1(data_in[2]), .A2(n844), .B1(n1120), .B2(\mem[9][2] ), 
        .ZN(n1118) );
  INV_X1 U237 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U238 ( .A1(data_in[3]), .A2(n844), .B1(n1120), .B2(\mem[9][3] ), 
        .ZN(n1117) );
  INV_X1 U239 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U240 ( .A1(data_in[4]), .A2(n844), .B1(n1120), .B2(\mem[9][4] ), 
        .ZN(n1116) );
  INV_X1 U241 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U242 ( .A1(data_in[5]), .A2(n844), .B1(n1120), .B2(\mem[9][5] ), 
        .ZN(n1115) );
  INV_X1 U243 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U244 ( .A1(data_in[6]), .A2(n844), .B1(n1120), .B2(\mem[9][6] ), 
        .ZN(n1114) );
  INV_X1 U245 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U246 ( .A1(data_in[7]), .A2(n844), .B1(n1120), .B2(\mem[9][7] ), 
        .ZN(n1113) );
  INV_X1 U247 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U248 ( .A1(data_in[0]), .A2(n843), .B1(n1111), .B2(\mem[10][0] ), 
        .ZN(n1112) );
  INV_X1 U249 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U250 ( .A1(data_in[1]), .A2(n843), .B1(n1111), .B2(\mem[10][1] ), 
        .ZN(n1110) );
  INV_X1 U251 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U252 ( .A1(data_in[2]), .A2(n843), .B1(n1111), .B2(\mem[10][2] ), 
        .ZN(n1109) );
  INV_X1 U253 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U254 ( .A1(data_in[3]), .A2(n843), .B1(n1111), .B2(\mem[10][3] ), 
        .ZN(n1108) );
  INV_X1 U255 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U256 ( .A1(data_in[4]), .A2(n843), .B1(n1111), .B2(\mem[10][4] ), 
        .ZN(n1107) );
  INV_X1 U257 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U258 ( .A1(data_in[5]), .A2(n843), .B1(n1111), .B2(\mem[10][5] ), 
        .ZN(n1106) );
  INV_X1 U259 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U260 ( .A1(data_in[6]), .A2(n843), .B1(n1111), .B2(\mem[10][6] ), 
        .ZN(n1105) );
  INV_X1 U261 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U262 ( .A1(data_in[7]), .A2(n843), .B1(n1111), .B2(\mem[10][7] ), 
        .ZN(n1104) );
  INV_X1 U263 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U264 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[11][0] ), 
        .ZN(n1103) );
  INV_X1 U265 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U266 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[11][1] ), 
        .ZN(n1101) );
  INV_X1 U267 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U268 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[11][2] ), 
        .ZN(n1100) );
  INV_X1 U269 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U270 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[11][3] ), 
        .ZN(n1099) );
  INV_X1 U271 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U272 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[11][4] ), 
        .ZN(n1098) );
  INV_X1 U273 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U274 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[11][5] ), 
        .ZN(n1097) );
  INV_X1 U275 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U276 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[11][6] ), 
        .ZN(n1096) );
  INV_X1 U277 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U278 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[11][7] ), 
        .ZN(n1095) );
  INV_X1 U279 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U280 ( .A1(data_in[0]), .A2(n841), .B1(n1093), .B2(\mem[12][0] ), 
        .ZN(n1094) );
  INV_X1 U281 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U282 ( .A1(data_in[1]), .A2(n841), .B1(n1093), .B2(\mem[12][1] ), 
        .ZN(n1092) );
  INV_X1 U283 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U284 ( .A1(data_in[2]), .A2(n841), .B1(n1093), .B2(\mem[12][2] ), 
        .ZN(n1091) );
  INV_X1 U285 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U286 ( .A1(data_in[3]), .A2(n841), .B1(n1093), .B2(\mem[12][3] ), 
        .ZN(n1090) );
  INV_X1 U287 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U288 ( .A1(data_in[4]), .A2(n841), .B1(n1093), .B2(\mem[12][4] ), 
        .ZN(n1089) );
  INV_X1 U289 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U290 ( .A1(data_in[5]), .A2(n841), .B1(n1093), .B2(\mem[12][5] ), 
        .ZN(n1088) );
  INV_X1 U291 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U292 ( .A1(data_in[6]), .A2(n841), .B1(n1093), .B2(\mem[12][6] ), 
        .ZN(n1087) );
  INV_X1 U293 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U294 ( .A1(data_in[7]), .A2(n841), .B1(n1093), .B2(\mem[12][7] ), 
        .ZN(n1086) );
  INV_X1 U295 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U296 ( .A1(data_in[0]), .A2(n840), .B1(n1084), .B2(\mem[13][0] ), 
        .ZN(n1085) );
  INV_X1 U297 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U298 ( .A1(data_in[1]), .A2(n840), .B1(n1084), .B2(\mem[13][1] ), 
        .ZN(n1083) );
  INV_X1 U299 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U300 ( .A1(data_in[2]), .A2(n840), .B1(n1084), .B2(\mem[13][2] ), 
        .ZN(n1082) );
  INV_X1 U301 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U302 ( .A1(data_in[3]), .A2(n840), .B1(n1084), .B2(\mem[13][3] ), 
        .ZN(n1081) );
  INV_X1 U303 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U304 ( .A1(data_in[4]), .A2(n840), .B1(n1084), .B2(\mem[13][4] ), 
        .ZN(n1080) );
  INV_X1 U305 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U306 ( .A1(data_in[5]), .A2(n840), .B1(n1084), .B2(\mem[13][5] ), 
        .ZN(n1079) );
  INV_X1 U307 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U308 ( .A1(data_in[6]), .A2(n840), .B1(n1084), .B2(\mem[13][6] ), 
        .ZN(n1078) );
  INV_X1 U309 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U310 ( .A1(data_in[7]), .A2(n840), .B1(n1084), .B2(\mem[13][7] ), 
        .ZN(n1077) );
  INV_X1 U311 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U312 ( .A1(data_in[0]), .A2(n839), .B1(n1075), .B2(\mem[14][0] ), 
        .ZN(n1076) );
  INV_X1 U313 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U314 ( .A1(data_in[1]), .A2(n839), .B1(n1075), .B2(\mem[14][1] ), 
        .ZN(n1074) );
  INV_X1 U315 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U316 ( .A1(data_in[2]), .A2(n839), .B1(n1075), .B2(\mem[14][2] ), 
        .ZN(n1073) );
  INV_X1 U317 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U318 ( .A1(data_in[3]), .A2(n839), .B1(n1075), .B2(\mem[14][3] ), 
        .ZN(n1072) );
  INV_X1 U319 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U320 ( .A1(data_in[4]), .A2(n839), .B1(n1075), .B2(\mem[14][4] ), 
        .ZN(n1071) );
  INV_X1 U321 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U322 ( .A1(data_in[5]), .A2(n839), .B1(n1075), .B2(\mem[14][5] ), 
        .ZN(n1070) );
  INV_X1 U323 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U324 ( .A1(data_in[6]), .A2(n839), .B1(n1075), .B2(\mem[14][6] ), 
        .ZN(n1069) );
  INV_X1 U325 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U326 ( .A1(data_in[7]), .A2(n839), .B1(n1075), .B2(\mem[14][7] ), 
        .ZN(n1068) );
  INV_X1 U327 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U328 ( .A1(data_in[0]), .A2(n838), .B1(n1066), .B2(\mem[15][0] ), 
        .ZN(n1067) );
  INV_X1 U329 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U330 ( .A1(data_in[1]), .A2(n838), .B1(n1066), .B2(\mem[15][1] ), 
        .ZN(n1065) );
  INV_X1 U331 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U332 ( .A1(data_in[2]), .A2(n838), .B1(n1066), .B2(\mem[15][2] ), 
        .ZN(n1064) );
  INV_X1 U333 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U334 ( .A1(data_in[3]), .A2(n838), .B1(n1066), .B2(\mem[15][3] ), 
        .ZN(n1063) );
  INV_X1 U335 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U336 ( .A1(data_in[4]), .A2(n838), .B1(n1066), .B2(\mem[15][4] ), 
        .ZN(n1062) );
  INV_X1 U337 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U338 ( .A1(data_in[5]), .A2(n838), .B1(n1066), .B2(\mem[15][5] ), 
        .ZN(n1061) );
  INV_X1 U339 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U340 ( .A1(data_in[6]), .A2(n838), .B1(n1066), .B2(\mem[15][6] ), 
        .ZN(n1060) );
  INV_X1 U341 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U342 ( .A1(data_in[7]), .A2(n838), .B1(n1066), .B2(\mem[15][7] ), 
        .ZN(n1059) );
  INV_X1 U343 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U344 ( .A1(data_in[0]), .A2(n837), .B1(n1057), .B2(\mem[16][0] ), 
        .ZN(n1058) );
  INV_X1 U345 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U346 ( .A1(data_in[1]), .A2(n837), .B1(n1057), .B2(\mem[16][1] ), 
        .ZN(n1056) );
  INV_X1 U347 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U348 ( .A1(data_in[2]), .A2(n837), .B1(n1057), .B2(\mem[16][2] ), 
        .ZN(n1055) );
  INV_X1 U349 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U350 ( .A1(data_in[3]), .A2(n837), .B1(n1057), .B2(\mem[16][3] ), 
        .ZN(n1054) );
  INV_X1 U351 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U352 ( .A1(data_in[4]), .A2(n837), .B1(n1057), .B2(\mem[16][4] ), 
        .ZN(n1053) );
  INV_X1 U353 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U354 ( .A1(data_in[5]), .A2(n837), .B1(n1057), .B2(\mem[16][5] ), 
        .ZN(n1052) );
  INV_X1 U355 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U356 ( .A1(data_in[6]), .A2(n837), .B1(n1057), .B2(\mem[16][6] ), 
        .ZN(n1051) );
  INV_X1 U357 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U358 ( .A1(data_in[7]), .A2(n837), .B1(n1057), .B2(\mem[16][7] ), 
        .ZN(n1050) );
  INV_X1 U359 ( .A(n1048), .ZN(n749) );
  AOI22_X1 U360 ( .A1(data_in[0]), .A2(n836), .B1(n1047), .B2(\mem[17][0] ), 
        .ZN(n1048) );
  INV_X1 U361 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U362 ( .A1(data_in[1]), .A2(n836), .B1(n1047), .B2(\mem[17][1] ), 
        .ZN(n1046) );
  INV_X1 U363 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U364 ( .A1(data_in[2]), .A2(n836), .B1(n1047), .B2(\mem[17][2] ), 
        .ZN(n1045) );
  INV_X1 U365 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U366 ( .A1(data_in[3]), .A2(n836), .B1(n1047), .B2(\mem[17][3] ), 
        .ZN(n1044) );
  INV_X1 U367 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U368 ( .A1(data_in[4]), .A2(n836), .B1(n1047), .B2(\mem[17][4] ), 
        .ZN(n1043) );
  INV_X1 U369 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U370 ( .A1(data_in[5]), .A2(n836), .B1(n1047), .B2(\mem[17][5] ), 
        .ZN(n1042) );
  INV_X1 U371 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U372 ( .A1(data_in[6]), .A2(n836), .B1(n1047), .B2(\mem[17][6] ), 
        .ZN(n1041) );
  INV_X1 U373 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U374 ( .A1(data_in[7]), .A2(n836), .B1(n1047), .B2(\mem[17][7] ), 
        .ZN(n1040) );
  INV_X1 U375 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U376 ( .A1(data_in[0]), .A2(n835), .B1(n1038), .B2(\mem[18][0] ), 
        .ZN(n1039) );
  INV_X1 U377 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U378 ( .A1(data_in[1]), .A2(n835), .B1(n1038), .B2(\mem[18][1] ), 
        .ZN(n1037) );
  INV_X1 U379 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U380 ( .A1(data_in[2]), .A2(n835), .B1(n1038), .B2(\mem[18][2] ), 
        .ZN(n1036) );
  INV_X1 U381 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U382 ( .A1(data_in[3]), .A2(n835), .B1(n1038), .B2(\mem[18][3] ), 
        .ZN(n1035) );
  INV_X1 U383 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U384 ( .A1(data_in[4]), .A2(n835), .B1(n1038), .B2(\mem[18][4] ), 
        .ZN(n1034) );
  INV_X1 U385 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U386 ( .A1(data_in[5]), .A2(n835), .B1(n1038), .B2(\mem[18][5] ), 
        .ZN(n1033) );
  INV_X1 U387 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U388 ( .A1(data_in[6]), .A2(n835), .B1(n1038), .B2(\mem[18][6] ), 
        .ZN(n1032) );
  INV_X1 U389 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U390 ( .A1(data_in[7]), .A2(n835), .B1(n1038), .B2(\mem[18][7] ), 
        .ZN(n1031) );
  INV_X1 U391 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U392 ( .A1(data_in[0]), .A2(n834), .B1(n1029), .B2(\mem[19][0] ), 
        .ZN(n1030) );
  INV_X1 U393 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U394 ( .A1(data_in[1]), .A2(n834), .B1(n1029), .B2(\mem[19][1] ), 
        .ZN(n1028) );
  INV_X1 U395 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U396 ( .A1(data_in[2]), .A2(n834), .B1(n1029), .B2(\mem[19][2] ), 
        .ZN(n1027) );
  INV_X1 U397 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U398 ( .A1(data_in[3]), .A2(n834), .B1(n1029), .B2(\mem[19][3] ), 
        .ZN(n1026) );
  INV_X1 U399 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U400 ( .A1(data_in[4]), .A2(n834), .B1(n1029), .B2(\mem[19][4] ), 
        .ZN(n1025) );
  INV_X1 U401 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U402 ( .A1(data_in[5]), .A2(n834), .B1(n1029), .B2(\mem[19][5] ), 
        .ZN(n1024) );
  INV_X1 U403 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U404 ( .A1(data_in[6]), .A2(n834), .B1(n1029), .B2(\mem[19][6] ), 
        .ZN(n1023) );
  INV_X1 U405 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U406 ( .A1(data_in[7]), .A2(n834), .B1(n1029), .B2(\mem[19][7] ), 
        .ZN(n1022) );
  INV_X1 U407 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U408 ( .A1(data_in[0]), .A2(n833), .B1(n1020), .B2(\mem[20][0] ), 
        .ZN(n1021) );
  INV_X1 U409 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U410 ( .A1(data_in[1]), .A2(n833), .B1(n1020), .B2(\mem[20][1] ), 
        .ZN(n1019) );
  INV_X1 U411 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U412 ( .A1(data_in[2]), .A2(n833), .B1(n1020), .B2(\mem[20][2] ), 
        .ZN(n1018) );
  INV_X1 U413 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U414 ( .A1(data_in[3]), .A2(n833), .B1(n1020), .B2(\mem[20][3] ), 
        .ZN(n1017) );
  INV_X1 U415 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U416 ( .A1(data_in[4]), .A2(n833), .B1(n1020), .B2(\mem[20][4] ), 
        .ZN(n1016) );
  INV_X1 U417 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U418 ( .A1(data_in[5]), .A2(n833), .B1(n1020), .B2(\mem[20][5] ), 
        .ZN(n1015) );
  INV_X1 U419 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U420 ( .A1(data_in[6]), .A2(n833), .B1(n1020), .B2(\mem[20][6] ), 
        .ZN(n1014) );
  INV_X1 U421 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U422 ( .A1(data_in[7]), .A2(n833), .B1(n1020), .B2(\mem[20][7] ), 
        .ZN(n1013) );
  INV_X1 U423 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U424 ( .A1(data_in[0]), .A2(n832), .B1(n1011), .B2(\mem[21][0] ), 
        .ZN(n1012) );
  INV_X1 U425 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U426 ( .A1(data_in[1]), .A2(n832), .B1(n1011), .B2(\mem[21][1] ), 
        .ZN(n1010) );
  INV_X1 U427 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U428 ( .A1(data_in[2]), .A2(n832), .B1(n1011), .B2(\mem[21][2] ), 
        .ZN(n1009) );
  INV_X1 U429 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U430 ( .A1(data_in[3]), .A2(n832), .B1(n1011), .B2(\mem[21][3] ), 
        .ZN(n1008) );
  INV_X1 U431 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U432 ( .A1(data_in[4]), .A2(n832), .B1(n1011), .B2(\mem[21][4] ), 
        .ZN(n1007) );
  INV_X1 U433 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U434 ( .A1(data_in[5]), .A2(n832), .B1(n1011), .B2(\mem[21][5] ), 
        .ZN(n1006) );
  INV_X1 U435 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U436 ( .A1(data_in[6]), .A2(n832), .B1(n1011), .B2(\mem[21][6] ), 
        .ZN(n1005) );
  INV_X1 U437 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U438 ( .A1(data_in[7]), .A2(n832), .B1(n1011), .B2(\mem[21][7] ), 
        .ZN(n1004) );
  INV_X1 U439 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U440 ( .A1(data_in[0]), .A2(n831), .B1(n1002), .B2(\mem[22][0] ), 
        .ZN(n1003) );
  INV_X1 U441 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U442 ( .A1(data_in[1]), .A2(n831), .B1(n1002), .B2(\mem[22][1] ), 
        .ZN(n1001) );
  INV_X1 U443 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U444 ( .A1(data_in[2]), .A2(n831), .B1(n1002), .B2(\mem[22][2] ), 
        .ZN(n1000) );
  INV_X1 U445 ( .A(n999), .ZN(n706) );
  AOI22_X1 U446 ( .A1(data_in[3]), .A2(n831), .B1(n1002), .B2(\mem[22][3] ), 
        .ZN(n999) );
  INV_X1 U447 ( .A(n998), .ZN(n705) );
  AOI22_X1 U448 ( .A1(data_in[4]), .A2(n831), .B1(n1002), .B2(\mem[22][4] ), 
        .ZN(n998) );
  INV_X1 U449 ( .A(n997), .ZN(n704) );
  AOI22_X1 U450 ( .A1(data_in[5]), .A2(n831), .B1(n1002), .B2(\mem[22][5] ), 
        .ZN(n997) );
  INV_X1 U451 ( .A(n996), .ZN(n703) );
  AOI22_X1 U452 ( .A1(data_in[6]), .A2(n831), .B1(n1002), .B2(\mem[22][6] ), 
        .ZN(n996) );
  INV_X1 U453 ( .A(n995), .ZN(n702) );
  AOI22_X1 U454 ( .A1(data_in[7]), .A2(n831), .B1(n1002), .B2(\mem[22][7] ), 
        .ZN(n995) );
  INV_X1 U455 ( .A(n994), .ZN(n701) );
  AOI22_X1 U456 ( .A1(data_in[0]), .A2(n830), .B1(n993), .B2(\mem[23][0] ), 
        .ZN(n994) );
  INV_X1 U457 ( .A(n992), .ZN(n700) );
  AOI22_X1 U458 ( .A1(data_in[1]), .A2(n830), .B1(n993), .B2(\mem[23][1] ), 
        .ZN(n992) );
  INV_X1 U459 ( .A(n991), .ZN(n699) );
  AOI22_X1 U460 ( .A1(data_in[2]), .A2(n830), .B1(n993), .B2(\mem[23][2] ), 
        .ZN(n991) );
  INV_X1 U461 ( .A(n990), .ZN(n698) );
  AOI22_X1 U462 ( .A1(data_in[3]), .A2(n830), .B1(n993), .B2(\mem[23][3] ), 
        .ZN(n990) );
  INV_X1 U463 ( .A(n989), .ZN(n697) );
  AOI22_X1 U464 ( .A1(data_in[4]), .A2(n830), .B1(n993), .B2(\mem[23][4] ), 
        .ZN(n989) );
  INV_X1 U465 ( .A(n988), .ZN(n696) );
  AOI22_X1 U466 ( .A1(data_in[5]), .A2(n830), .B1(n993), .B2(\mem[23][5] ), 
        .ZN(n988) );
  INV_X1 U467 ( .A(n987), .ZN(n695) );
  AOI22_X1 U468 ( .A1(data_in[6]), .A2(n830), .B1(n993), .B2(\mem[23][6] ), 
        .ZN(n987) );
  INV_X1 U469 ( .A(n986), .ZN(n694) );
  AOI22_X1 U470 ( .A1(data_in[7]), .A2(n830), .B1(n993), .B2(\mem[23][7] ), 
        .ZN(n986) );
  INV_X1 U471 ( .A(n985), .ZN(n693) );
  AOI22_X1 U472 ( .A1(data_in[0]), .A2(n829), .B1(n984), .B2(\mem[24][0] ), 
        .ZN(n985) );
  INV_X1 U473 ( .A(n983), .ZN(n692) );
  AOI22_X1 U474 ( .A1(data_in[1]), .A2(n829), .B1(n984), .B2(\mem[24][1] ), 
        .ZN(n983) );
  INV_X1 U475 ( .A(n982), .ZN(n691) );
  AOI22_X1 U476 ( .A1(data_in[2]), .A2(n829), .B1(n984), .B2(\mem[24][2] ), 
        .ZN(n982) );
  INV_X1 U477 ( .A(n981), .ZN(n690) );
  AOI22_X1 U478 ( .A1(data_in[3]), .A2(n829), .B1(n984), .B2(\mem[24][3] ), 
        .ZN(n981) );
  INV_X1 U479 ( .A(n980), .ZN(n689) );
  AOI22_X1 U480 ( .A1(data_in[4]), .A2(n829), .B1(n984), .B2(\mem[24][4] ), 
        .ZN(n980) );
  INV_X1 U481 ( .A(n979), .ZN(n688) );
  AOI22_X1 U482 ( .A1(data_in[5]), .A2(n829), .B1(n984), .B2(\mem[24][5] ), 
        .ZN(n979) );
  INV_X1 U483 ( .A(n978), .ZN(n687) );
  AOI22_X1 U484 ( .A1(data_in[6]), .A2(n829), .B1(n984), .B2(\mem[24][6] ), 
        .ZN(n978) );
  INV_X1 U485 ( .A(n977), .ZN(n686) );
  AOI22_X1 U486 ( .A1(data_in[7]), .A2(n829), .B1(n984), .B2(\mem[24][7] ), 
        .ZN(n977) );
  INV_X1 U487 ( .A(n975), .ZN(n685) );
  AOI22_X1 U488 ( .A1(data_in[0]), .A2(n828), .B1(n974), .B2(\mem[25][0] ), 
        .ZN(n975) );
  INV_X1 U489 ( .A(n973), .ZN(n684) );
  AOI22_X1 U490 ( .A1(data_in[1]), .A2(n828), .B1(n974), .B2(\mem[25][1] ), 
        .ZN(n973) );
  INV_X1 U491 ( .A(n972), .ZN(n683) );
  AOI22_X1 U492 ( .A1(data_in[2]), .A2(n828), .B1(n974), .B2(\mem[25][2] ), 
        .ZN(n972) );
  INV_X1 U493 ( .A(n971), .ZN(n682) );
  AOI22_X1 U494 ( .A1(data_in[3]), .A2(n828), .B1(n974), .B2(\mem[25][3] ), 
        .ZN(n971) );
  INV_X1 U495 ( .A(n970), .ZN(n681) );
  AOI22_X1 U496 ( .A1(data_in[4]), .A2(n828), .B1(n974), .B2(\mem[25][4] ), 
        .ZN(n970) );
  INV_X1 U497 ( .A(n969), .ZN(n680) );
  AOI22_X1 U498 ( .A1(data_in[5]), .A2(n828), .B1(n974), .B2(\mem[25][5] ), 
        .ZN(n969) );
  INV_X1 U499 ( .A(n968), .ZN(n679) );
  AOI22_X1 U500 ( .A1(data_in[6]), .A2(n828), .B1(n974), .B2(\mem[25][6] ), 
        .ZN(n968) );
  INV_X1 U501 ( .A(n967), .ZN(n678) );
  AOI22_X1 U502 ( .A1(data_in[7]), .A2(n828), .B1(n974), .B2(\mem[25][7] ), 
        .ZN(n967) );
  INV_X1 U503 ( .A(n966), .ZN(n677) );
  AOI22_X1 U504 ( .A1(data_in[0]), .A2(n827), .B1(n965), .B2(\mem[26][0] ), 
        .ZN(n966) );
  INV_X1 U505 ( .A(n964), .ZN(n676) );
  AOI22_X1 U506 ( .A1(data_in[1]), .A2(n827), .B1(n965), .B2(\mem[26][1] ), 
        .ZN(n964) );
  INV_X1 U507 ( .A(n963), .ZN(n675) );
  AOI22_X1 U508 ( .A1(data_in[2]), .A2(n827), .B1(n965), .B2(\mem[26][2] ), 
        .ZN(n963) );
  INV_X1 U509 ( .A(n962), .ZN(n674) );
  AOI22_X1 U510 ( .A1(data_in[3]), .A2(n827), .B1(n965), .B2(\mem[26][3] ), 
        .ZN(n962) );
  INV_X1 U511 ( .A(n961), .ZN(n673) );
  AOI22_X1 U512 ( .A1(data_in[4]), .A2(n827), .B1(n965), .B2(\mem[26][4] ), 
        .ZN(n961) );
  INV_X1 U513 ( .A(n960), .ZN(n672) );
  AOI22_X1 U514 ( .A1(data_in[5]), .A2(n827), .B1(n965), .B2(\mem[26][5] ), 
        .ZN(n960) );
  INV_X1 U515 ( .A(n959), .ZN(n671) );
  AOI22_X1 U516 ( .A1(data_in[6]), .A2(n827), .B1(n965), .B2(\mem[26][6] ), 
        .ZN(n959) );
  INV_X1 U517 ( .A(n958), .ZN(n670) );
  AOI22_X1 U518 ( .A1(data_in[7]), .A2(n827), .B1(n965), .B2(\mem[26][7] ), 
        .ZN(n958) );
  INV_X1 U519 ( .A(n957), .ZN(n669) );
  AOI22_X1 U520 ( .A1(data_in[0]), .A2(n826), .B1(n956), .B2(\mem[27][0] ), 
        .ZN(n957) );
  INV_X1 U521 ( .A(n955), .ZN(n668) );
  AOI22_X1 U522 ( .A1(data_in[1]), .A2(n826), .B1(n956), .B2(\mem[27][1] ), 
        .ZN(n955) );
  INV_X1 U523 ( .A(n954), .ZN(n667) );
  AOI22_X1 U524 ( .A1(data_in[2]), .A2(n826), .B1(n956), .B2(\mem[27][2] ), 
        .ZN(n954) );
  INV_X1 U525 ( .A(n953), .ZN(n666) );
  AOI22_X1 U526 ( .A1(data_in[3]), .A2(n826), .B1(n956), .B2(\mem[27][3] ), 
        .ZN(n953) );
  INV_X1 U527 ( .A(n952), .ZN(n665) );
  AOI22_X1 U528 ( .A1(data_in[4]), .A2(n826), .B1(n956), .B2(\mem[27][4] ), 
        .ZN(n952) );
  INV_X1 U529 ( .A(n951), .ZN(n664) );
  AOI22_X1 U530 ( .A1(data_in[5]), .A2(n826), .B1(n956), .B2(\mem[27][5] ), 
        .ZN(n951) );
  INV_X1 U531 ( .A(n950), .ZN(n663) );
  AOI22_X1 U532 ( .A1(data_in[6]), .A2(n826), .B1(n956), .B2(\mem[27][6] ), 
        .ZN(n950) );
  INV_X1 U533 ( .A(n949), .ZN(n662) );
  AOI22_X1 U534 ( .A1(data_in[7]), .A2(n826), .B1(n956), .B2(\mem[27][7] ), 
        .ZN(n949) );
  INV_X1 U535 ( .A(n948), .ZN(n661) );
  AOI22_X1 U536 ( .A1(data_in[0]), .A2(n825), .B1(n947), .B2(\mem[28][0] ), 
        .ZN(n948) );
  INV_X1 U537 ( .A(n946), .ZN(n660) );
  AOI22_X1 U538 ( .A1(data_in[1]), .A2(n825), .B1(n947), .B2(\mem[28][1] ), 
        .ZN(n946) );
  INV_X1 U539 ( .A(n945), .ZN(n659) );
  AOI22_X1 U540 ( .A1(data_in[2]), .A2(n825), .B1(n947), .B2(\mem[28][2] ), 
        .ZN(n945) );
  INV_X1 U541 ( .A(n944), .ZN(n658) );
  AOI22_X1 U542 ( .A1(data_in[3]), .A2(n825), .B1(n947), .B2(\mem[28][3] ), 
        .ZN(n944) );
  INV_X1 U543 ( .A(n943), .ZN(n657) );
  AOI22_X1 U544 ( .A1(data_in[4]), .A2(n825), .B1(n947), .B2(\mem[28][4] ), 
        .ZN(n943) );
  INV_X1 U545 ( .A(n942), .ZN(n656) );
  AOI22_X1 U546 ( .A1(data_in[5]), .A2(n825), .B1(n947), .B2(\mem[28][5] ), 
        .ZN(n942) );
  INV_X1 U547 ( .A(n941), .ZN(n655) );
  AOI22_X1 U548 ( .A1(data_in[6]), .A2(n825), .B1(n947), .B2(\mem[28][6] ), 
        .ZN(n941) );
  INV_X1 U549 ( .A(n940), .ZN(n654) );
  AOI22_X1 U550 ( .A1(data_in[7]), .A2(n825), .B1(n947), .B2(\mem[28][7] ), 
        .ZN(n940) );
  INV_X1 U551 ( .A(n939), .ZN(n653) );
  AOI22_X1 U552 ( .A1(data_in[0]), .A2(n824), .B1(n938), .B2(\mem[29][0] ), 
        .ZN(n939) );
  INV_X1 U553 ( .A(n937), .ZN(n652) );
  AOI22_X1 U554 ( .A1(data_in[1]), .A2(n824), .B1(n938), .B2(\mem[29][1] ), 
        .ZN(n937) );
  INV_X1 U555 ( .A(n936), .ZN(n651) );
  AOI22_X1 U556 ( .A1(data_in[2]), .A2(n824), .B1(n938), .B2(\mem[29][2] ), 
        .ZN(n936) );
  INV_X1 U557 ( .A(n935), .ZN(n650) );
  AOI22_X1 U558 ( .A1(data_in[3]), .A2(n824), .B1(n938), .B2(\mem[29][3] ), 
        .ZN(n935) );
  INV_X1 U559 ( .A(n934), .ZN(n649) );
  AOI22_X1 U560 ( .A1(data_in[4]), .A2(n824), .B1(n938), .B2(\mem[29][4] ), 
        .ZN(n934) );
  INV_X1 U561 ( .A(n933), .ZN(n648) );
  AOI22_X1 U562 ( .A1(data_in[5]), .A2(n824), .B1(n938), .B2(\mem[29][5] ), 
        .ZN(n933) );
  INV_X1 U563 ( .A(n932), .ZN(n647) );
  AOI22_X1 U564 ( .A1(data_in[6]), .A2(n824), .B1(n938), .B2(\mem[29][6] ), 
        .ZN(n932) );
  INV_X1 U565 ( .A(n931), .ZN(n646) );
  AOI22_X1 U566 ( .A1(data_in[7]), .A2(n824), .B1(n938), .B2(\mem[29][7] ), 
        .ZN(n931) );
  INV_X1 U567 ( .A(n930), .ZN(n645) );
  AOI22_X1 U568 ( .A1(data_in[0]), .A2(n823), .B1(n929), .B2(\mem[30][0] ), 
        .ZN(n930) );
  INV_X1 U569 ( .A(n928), .ZN(n644) );
  AOI22_X1 U570 ( .A1(data_in[1]), .A2(n823), .B1(n929), .B2(\mem[30][1] ), 
        .ZN(n928) );
  INV_X1 U571 ( .A(n927), .ZN(n643) );
  AOI22_X1 U572 ( .A1(data_in[2]), .A2(n823), .B1(n929), .B2(\mem[30][2] ), 
        .ZN(n927) );
  INV_X1 U573 ( .A(n926), .ZN(n642) );
  AOI22_X1 U574 ( .A1(data_in[3]), .A2(n823), .B1(n929), .B2(\mem[30][3] ), 
        .ZN(n926) );
  INV_X1 U575 ( .A(n925), .ZN(n641) );
  AOI22_X1 U576 ( .A1(data_in[4]), .A2(n823), .B1(n929), .B2(\mem[30][4] ), 
        .ZN(n925) );
  INV_X1 U577 ( .A(n924), .ZN(n640) );
  AOI22_X1 U578 ( .A1(data_in[5]), .A2(n823), .B1(n929), .B2(\mem[30][5] ), 
        .ZN(n924) );
  INV_X1 U579 ( .A(n923), .ZN(n639) );
  AOI22_X1 U580 ( .A1(data_in[6]), .A2(n823), .B1(n929), .B2(\mem[30][6] ), 
        .ZN(n923) );
  INV_X1 U581 ( .A(n922), .ZN(n638) );
  AOI22_X1 U582 ( .A1(data_in[7]), .A2(n823), .B1(n929), .B2(\mem[30][7] ), 
        .ZN(n922) );
  INV_X1 U583 ( .A(n921), .ZN(n637) );
  AOI22_X1 U584 ( .A1(data_in[0]), .A2(n822), .B1(n920), .B2(\mem[31][0] ), 
        .ZN(n921) );
  INV_X1 U585 ( .A(n919), .ZN(n636) );
  AOI22_X1 U586 ( .A1(data_in[1]), .A2(n822), .B1(n920), .B2(\mem[31][1] ), 
        .ZN(n919) );
  INV_X1 U587 ( .A(n918), .ZN(n635) );
  AOI22_X1 U588 ( .A1(data_in[2]), .A2(n822), .B1(n920), .B2(\mem[31][2] ), 
        .ZN(n918) );
  INV_X1 U589 ( .A(n917), .ZN(n634) );
  AOI22_X1 U590 ( .A1(data_in[3]), .A2(n822), .B1(n920), .B2(\mem[31][3] ), 
        .ZN(n917) );
  INV_X1 U591 ( .A(n916), .ZN(n633) );
  AOI22_X1 U592 ( .A1(data_in[4]), .A2(n822), .B1(n920), .B2(\mem[31][4] ), 
        .ZN(n916) );
  INV_X1 U593 ( .A(n915), .ZN(n632) );
  AOI22_X1 U594 ( .A1(data_in[5]), .A2(n822), .B1(n920), .B2(\mem[31][5] ), 
        .ZN(n915) );
  INV_X1 U595 ( .A(n914), .ZN(n631) );
  AOI22_X1 U596 ( .A1(data_in[6]), .A2(n822), .B1(n920), .B2(\mem[31][6] ), 
        .ZN(n914) );
  INV_X1 U597 ( .A(n913), .ZN(n630) );
  AOI22_X1 U598 ( .A1(data_in[7]), .A2(n822), .B1(n920), .B2(\mem[31][7] ), 
        .ZN(n913) );
  MUX2_X1 U599 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n611), .Z(n1) );
  MUX2_X1 U600 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n611), .Z(n2) );
  MUX2_X1 U601 ( .A(n2), .B(n1), .S(n608), .Z(n3) );
  MUX2_X1 U602 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n611), .Z(n4) );
  MUX2_X1 U603 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n611), .Z(n5) );
  MUX2_X1 U604 ( .A(n5), .B(n4), .S(n608), .Z(n6) );
  MUX2_X1 U605 ( .A(n6), .B(n3), .S(n606), .Z(n7) );
  MUX2_X1 U606 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n611), .Z(n8) );
  MUX2_X1 U607 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n611), .Z(n9) );
  MUX2_X1 U608 ( .A(n9), .B(n8), .S(n608), .Z(n10) );
  MUX2_X1 U609 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n611), .Z(n11) );
  MUX2_X1 U610 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n611), .Z(n12) );
  MUX2_X1 U611 ( .A(n12), .B(n11), .S(n608), .Z(n13) );
  MUX2_X1 U612 ( .A(n13), .B(n10), .S(n606), .Z(n14) );
  MUX2_X1 U613 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U614 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n612), .Z(n16) );
  MUX2_X1 U615 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n612), .Z(n17) );
  MUX2_X1 U616 ( .A(n17), .B(n16), .S(n609), .Z(n18) );
  MUX2_X1 U617 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n612), .Z(n19) );
  MUX2_X1 U618 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n612), .Z(n20) );
  MUX2_X1 U619 ( .A(n20), .B(n19), .S(n609), .Z(n21) );
  MUX2_X1 U620 ( .A(n21), .B(n18), .S(n606), .Z(n22) );
  MUX2_X1 U621 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n612), .Z(n23) );
  MUX2_X1 U622 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n612), .Z(n24) );
  MUX2_X1 U623 ( .A(n24), .B(n23), .S(n609), .Z(n25) );
  MUX2_X1 U624 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n612), .Z(n26) );
  MUX2_X1 U625 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n612), .Z(n27) );
  MUX2_X1 U626 ( .A(n27), .B(n26), .S(n609), .Z(n28) );
  MUX2_X1 U627 ( .A(n28), .B(n25), .S(n606), .Z(n29) );
  MUX2_X1 U628 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U629 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U630 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n612), .Z(n31) );
  MUX2_X1 U631 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n612), .Z(n32) );
  MUX2_X1 U632 ( .A(n32), .B(n31), .S(n609), .Z(n33) );
  MUX2_X1 U633 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n612), .Z(n34) );
  MUX2_X1 U634 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n612), .Z(n35) );
  MUX2_X1 U635 ( .A(n35), .B(n34), .S(n609), .Z(n36) );
  MUX2_X1 U636 ( .A(n36), .B(n33), .S(n606), .Z(n37) );
  MUX2_X1 U637 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n611), .Z(n38) );
  MUX2_X1 U638 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n616), .Z(n39) );
  MUX2_X1 U639 ( .A(n39), .B(n38), .S(n609), .Z(n40) );
  MUX2_X1 U640 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n615), .Z(n41) );
  MUX2_X1 U641 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n617), .Z(n42) );
  MUX2_X1 U642 ( .A(n42), .B(n41), .S(n609), .Z(n43) );
  MUX2_X1 U643 ( .A(n43), .B(n40), .S(n606), .Z(n44) );
  MUX2_X1 U644 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U645 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n611), .Z(n46) );
  MUX2_X1 U646 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n619), .Z(n47) );
  MUX2_X1 U647 ( .A(n47), .B(n46), .S(n609), .Z(n48) );
  MUX2_X1 U648 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n611), .Z(n49) );
  MUX2_X1 U649 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n612), .Z(n50) );
  MUX2_X1 U650 ( .A(n50), .B(n49), .S(n609), .Z(n51) );
  MUX2_X1 U651 ( .A(n51), .B(n48), .S(n606), .Z(n52) );
  MUX2_X1 U652 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n611), .Z(n53) );
  MUX2_X1 U653 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n618), .Z(n54) );
  MUX2_X1 U654 ( .A(n54), .B(n53), .S(n609), .Z(n55) );
  MUX2_X1 U655 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n619), .Z(n56) );
  MUX2_X1 U656 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n619), .Z(n57) );
  MUX2_X1 U657 ( .A(n57), .B(n56), .S(n609), .Z(n58) );
  MUX2_X1 U658 ( .A(n58), .B(n55), .S(n606), .Z(n59) );
  MUX2_X1 U659 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U660 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U661 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n613), .Z(n61) );
  MUX2_X1 U662 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n613), .Z(n62) );
  MUX2_X1 U663 ( .A(n62), .B(n61), .S(n610), .Z(n63) );
  MUX2_X1 U664 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n613), .Z(n64) );
  MUX2_X1 U665 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n613), .Z(n65) );
  MUX2_X1 U666 ( .A(n65), .B(n64), .S(n610), .Z(n66) );
  MUX2_X1 U667 ( .A(n66), .B(n63), .S(n607), .Z(n67) );
  MUX2_X1 U668 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n613), .Z(n68) );
  MUX2_X1 U669 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n613), .Z(n69) );
  MUX2_X1 U670 ( .A(n69), .B(n68), .S(n610), .Z(n70) );
  MUX2_X1 U671 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n613), .Z(n71) );
  MUX2_X1 U672 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n613), .Z(n72) );
  MUX2_X1 U673 ( .A(n72), .B(n71), .S(n610), .Z(n73) );
  MUX2_X1 U674 ( .A(n73), .B(n70), .S(N12), .Z(n74) );
  MUX2_X1 U675 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U676 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n613), .Z(n76) );
  MUX2_X1 U677 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n613), .Z(n77) );
  MUX2_X1 U678 ( .A(n77), .B(n76), .S(n610), .Z(n78) );
  MUX2_X1 U679 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n613), .Z(n79) );
  MUX2_X1 U680 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n613), .Z(n80) );
  MUX2_X1 U681 ( .A(n80), .B(n79), .S(n610), .Z(n81) );
  MUX2_X1 U682 ( .A(n81), .B(n78), .S(n606), .Z(n82) );
  MUX2_X1 U683 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n614), .Z(n83) );
  MUX2_X1 U684 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n614), .Z(n84) );
  MUX2_X1 U685 ( .A(n84), .B(n83), .S(n610), .Z(n85) );
  MUX2_X1 U686 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n614), .Z(n86) );
  MUX2_X1 U687 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n614), .Z(n87) );
  MUX2_X1 U688 ( .A(n87), .B(n86), .S(n610), .Z(n88) );
  MUX2_X1 U689 ( .A(n88), .B(n85), .S(n606), .Z(n89) );
  MUX2_X1 U690 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U691 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U692 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n614), .Z(n91) );
  MUX2_X1 U693 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n614), .Z(n92) );
  MUX2_X1 U694 ( .A(n92), .B(n91), .S(n610), .Z(n93) );
  MUX2_X1 U695 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n614), .Z(n94) );
  MUX2_X1 U696 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n614), .Z(n95) );
  MUX2_X1 U697 ( .A(n95), .B(n94), .S(n610), .Z(n96) );
  MUX2_X1 U698 ( .A(n96), .B(n93), .S(n606), .Z(n97) );
  MUX2_X1 U699 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n614), .Z(n98) );
  MUX2_X1 U700 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n614), .Z(n99) );
  MUX2_X1 U701 ( .A(n99), .B(n98), .S(n610), .Z(n100) );
  MUX2_X1 U702 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n614), .Z(n101) );
  MUX2_X1 U703 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n614), .Z(n102) );
  MUX2_X1 U704 ( .A(n102), .B(n101), .S(n610), .Z(n103) );
  MUX2_X1 U705 ( .A(n103), .B(n100), .S(n606), .Z(n104) );
  MUX2_X1 U706 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U707 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n615), .Z(n106) );
  MUX2_X1 U708 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n615), .Z(n107) );
  MUX2_X1 U709 ( .A(n107), .B(n106), .S(n610), .Z(n108) );
  MUX2_X1 U710 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n615), .Z(n109) );
  MUX2_X1 U711 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n615), .Z(n110) );
  MUX2_X1 U712 ( .A(n110), .B(n109), .S(n609), .Z(n111) );
  MUX2_X1 U713 ( .A(n111), .B(n108), .S(n606), .Z(n112) );
  MUX2_X1 U714 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n615), .Z(n113) );
  MUX2_X1 U715 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n615), .Z(n114) );
  MUX2_X1 U716 ( .A(n114), .B(n113), .S(n608), .Z(n115) );
  MUX2_X1 U717 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n615), .Z(n116) );
  MUX2_X1 U718 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n615), .Z(n117) );
  MUX2_X1 U719 ( .A(n117), .B(n116), .S(n610), .Z(n118) );
  MUX2_X1 U720 ( .A(n118), .B(n115), .S(n606), .Z(n119) );
  MUX2_X1 U721 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U722 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U723 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n615), .Z(n121) );
  MUX2_X1 U724 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n615), .Z(n122) );
  MUX2_X1 U725 ( .A(n122), .B(n121), .S(n608), .Z(n123) );
  MUX2_X1 U726 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n615), .Z(n124) );
  MUX2_X1 U727 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n615), .Z(n125) );
  MUX2_X1 U728 ( .A(n125), .B(n124), .S(n608), .Z(n126) );
  MUX2_X1 U729 ( .A(n126), .B(n123), .S(N12), .Z(n127) );
  MUX2_X1 U730 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(N10), .Z(n128) );
  MUX2_X1 U731 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n618), .Z(n129) );
  MUX2_X1 U732 ( .A(n129), .B(n128), .S(n610), .Z(n130) );
  MUX2_X1 U733 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n612), .Z(n131) );
  MUX2_X1 U734 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n619), .Z(n132) );
  MUX2_X1 U735 ( .A(n132), .B(n131), .S(n609), .Z(n133) );
  MUX2_X1 U736 ( .A(n133), .B(n130), .S(n607), .Z(n134) );
  MUX2_X1 U737 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U738 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(N10), .Z(n136) );
  MUX2_X1 U739 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n616), .Z(n137) );
  MUX2_X1 U740 ( .A(n137), .B(n136), .S(n609), .Z(n138) );
  MUX2_X1 U741 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n619), .Z(n139) );
  MUX2_X1 U742 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n140) );
  MUX2_X1 U743 ( .A(n140), .B(n139), .S(n608), .Z(n141) );
  MUX2_X1 U744 ( .A(n141), .B(n138), .S(N12), .Z(n142) );
  MUX2_X1 U745 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(N10), .Z(n143) );
  MUX2_X1 U746 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n619), .Z(n144) );
  MUX2_X1 U747 ( .A(n144), .B(n143), .S(n609), .Z(n145) );
  MUX2_X1 U748 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n619), .Z(n146) );
  MUX2_X1 U749 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n147) );
  MUX2_X1 U750 ( .A(n147), .B(n146), .S(n608), .Z(n148) );
  MUX2_X1 U751 ( .A(n148), .B(n145), .S(n607), .Z(n149) );
  MUX2_X1 U752 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U753 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U754 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n613), .Z(n151) );
  MUX2_X1 U755 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n613), .Z(n152) );
  MUX2_X1 U756 ( .A(n152), .B(n151), .S(n609), .Z(n153) );
  MUX2_X1 U757 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n613), .Z(n154) );
  MUX2_X1 U758 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n613), .Z(n155) );
  MUX2_X1 U759 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U760 ( .A(n156), .B(n153), .S(n607), .Z(n157) );
  MUX2_X1 U761 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n613), .Z(n158) );
  MUX2_X1 U762 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n613), .Z(n159) );
  MUX2_X1 U763 ( .A(n159), .B(n158), .S(n608), .Z(n160) );
  MUX2_X1 U764 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n613), .Z(n161) );
  MUX2_X1 U765 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n614), .Z(n162) );
  MUX2_X1 U766 ( .A(n162), .B(n161), .S(N11), .Z(n163) );
  MUX2_X1 U767 ( .A(n163), .B(n160), .S(n607), .Z(n164) );
  MUX2_X1 U768 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U769 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n613), .Z(n166) );
  MUX2_X1 U770 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n613), .Z(n167) );
  MUX2_X1 U771 ( .A(n167), .B(n166), .S(n610), .Z(n168) );
  MUX2_X1 U772 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n613), .Z(n169) );
  MUX2_X1 U773 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n613), .Z(n170) );
  MUX2_X1 U774 ( .A(n170), .B(n169), .S(n610), .Z(n171) );
  MUX2_X1 U775 ( .A(n171), .B(n168), .S(n607), .Z(n172) );
  MUX2_X1 U776 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n616), .Z(n173) );
  MUX2_X1 U777 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n616), .Z(n174) );
  MUX2_X1 U778 ( .A(n174), .B(n173), .S(n610), .Z(n175) );
  MUX2_X1 U779 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n616), .Z(n176) );
  MUX2_X1 U780 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n616), .Z(n177) );
  MUX2_X1 U781 ( .A(n177), .B(n176), .S(n609), .Z(n178) );
  MUX2_X1 U782 ( .A(n178), .B(n175), .S(n607), .Z(n179) );
  MUX2_X1 U783 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U784 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U785 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n616), .Z(n181) );
  MUX2_X1 U786 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n616), .Z(n182) );
  MUX2_X1 U787 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U788 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n616), .Z(n184) );
  MUX2_X1 U789 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n616), .Z(n185) );
  MUX2_X1 U790 ( .A(n185), .B(n184), .S(n609), .Z(n186) );
  MUX2_X1 U791 ( .A(n186), .B(n183), .S(n607), .Z(n187) );
  MUX2_X1 U792 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n616), .Z(n188) );
  MUX2_X1 U793 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n616), .Z(n189) );
  MUX2_X1 U794 ( .A(n189), .B(n188), .S(N11), .Z(n190) );
  MUX2_X1 U795 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n616), .Z(n191) );
  MUX2_X1 U796 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n616), .Z(n192) );
  MUX2_X1 U797 ( .A(n192), .B(n191), .S(n609), .Z(n193) );
  MUX2_X1 U798 ( .A(n193), .B(n190), .S(n607), .Z(n194) );
  MUX2_X1 U799 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U800 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n617), .Z(n196) );
  MUX2_X1 U801 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n617), .Z(n197) );
  MUX2_X1 U802 ( .A(n197), .B(n196), .S(n608), .Z(n198) );
  MUX2_X1 U803 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n617), .Z(n199) );
  MUX2_X1 U804 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n617), .Z(n200) );
  MUX2_X1 U805 ( .A(n200), .B(n199), .S(n609), .Z(n201) );
  MUX2_X1 U806 ( .A(n201), .B(n198), .S(n607), .Z(n202) );
  MUX2_X1 U807 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n617), .Z(n203) );
  MUX2_X1 U808 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n617), .Z(n204) );
  MUX2_X1 U809 ( .A(n204), .B(n203), .S(n608), .Z(n205) );
  MUX2_X1 U810 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n617), .Z(n206) );
  MUX2_X1 U811 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n617), .Z(n207) );
  MUX2_X1 U812 ( .A(n207), .B(n206), .S(n610), .Z(n208) );
  MUX2_X1 U813 ( .A(n208), .B(n205), .S(n607), .Z(n209) );
  MUX2_X1 U814 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U815 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U816 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n617), .Z(n211) );
  MUX2_X1 U817 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n617), .Z(n212) );
  MUX2_X1 U818 ( .A(n212), .B(n211), .S(n608), .Z(n213) );
  MUX2_X1 U819 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n617), .Z(n214) );
  MUX2_X1 U820 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n617), .Z(n215) );
  MUX2_X1 U821 ( .A(n215), .B(n214), .S(n608), .Z(n216) );
  MUX2_X1 U822 ( .A(n216), .B(n213), .S(n607), .Z(n217) );
  MUX2_X1 U823 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n618), .Z(n218) );
  MUX2_X1 U824 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n618), .Z(n219) );
  MUX2_X1 U825 ( .A(n219), .B(n218), .S(n608), .Z(n220) );
  MUX2_X1 U826 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n618), .Z(n221) );
  MUX2_X1 U827 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n618), .Z(n222) );
  MUX2_X1 U828 ( .A(n222), .B(n221), .S(n610), .Z(n223) );
  MUX2_X1 U829 ( .A(n223), .B(n220), .S(n607), .Z(n224) );
  MUX2_X1 U830 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U831 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n618), .Z(n226) );
  MUX2_X1 U832 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n618), .Z(n227) );
  MUX2_X1 U833 ( .A(n227), .B(n226), .S(n608), .Z(n228) );
  MUX2_X1 U834 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n618), .Z(n229) );
  MUX2_X1 U835 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n618), .Z(n595) );
  MUX2_X1 U836 ( .A(n595), .B(n229), .S(N11), .Z(n596) );
  MUX2_X1 U837 ( .A(n596), .B(n228), .S(n607), .Z(n597) );
  MUX2_X1 U838 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n618), .Z(n598) );
  MUX2_X1 U839 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n618), .Z(n599) );
  MUX2_X1 U840 ( .A(n599), .B(n598), .S(n608), .Z(n600) );
  MUX2_X1 U841 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n618), .Z(n601) );
  MUX2_X1 U842 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n618), .Z(n602) );
  MUX2_X1 U843 ( .A(n602), .B(n601), .S(n608), .Z(n603) );
  MUX2_X1 U844 ( .A(n603), .B(n600), .S(n607), .Z(n604) );
  MUX2_X1 U845 ( .A(n604), .B(n597), .S(N13), .Z(n605) );
  MUX2_X1 U846 ( .A(n605), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U847 ( .A(N11), .Z(n608) );
  CLKBUF_X1 U848 ( .A(n619), .Z(n611) );
  INV_X1 U849 ( .A(N10), .ZN(n620) );
  INV_X1 U850 ( .A(N11), .ZN(n621) );
  INV_X1 U851 ( .A(data_in[0]), .ZN(n622) );
  INV_X1 U852 ( .A(data_in[1]), .ZN(n623) );
  INV_X1 U853 ( .A(data_in[2]), .ZN(n624) );
  INV_X1 U854 ( .A(data_in[3]), .ZN(n625) );
  INV_X1 U855 ( .A(data_in[4]), .ZN(n626) );
  INV_X1 U856 ( .A(data_in[5]), .ZN(n627) );
  INV_X1 U857 ( .A(data_in[6]), .ZN(n628) );
  INV_X1 U858 ( .A(data_in[7]), .ZN(n629) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_3 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n633), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n634), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n635), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n636), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n637), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n638), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n639), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n640), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n641), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n642), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n643), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n644), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n645), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n646), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n647), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n648), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n649), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n650), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n651), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n652), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n653), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n654), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n655), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n656), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n657), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n658), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n659), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n660), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n661), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n662), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n663), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n664), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n665), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n666), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n667), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n668), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n669), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n670), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n671), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n672), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n673), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n674), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n675), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n676), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n677), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n678), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n679), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n680), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n681), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n682), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n683), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n684), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n685), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n686), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n687), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n688), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n689), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n690), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n691), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n692), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n693), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n694), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n695), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n696), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n697), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n698), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n699), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n700), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n701), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n702), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n703), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n704), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n705), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n706), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n707), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n708), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n709), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n710), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n711), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n712), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n713), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n714), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n715), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n716), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n717), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n718), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n719), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n720), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n721), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n722), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n723), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n724), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n725), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n726), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n727), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n728), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n729), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n730), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n731), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n732), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n733), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n734), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n735), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n736), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n737), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n738), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n739), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n740), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n741), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n742), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n743), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n744), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n745), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n746), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n747), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n748), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n749), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n750), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n751), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n752), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n753), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n754), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n755), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n756), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n757), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n758), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n759), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n760), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n761), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n762), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n763), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n764), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n765), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n766), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n767), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n768), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n769), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n770), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n771), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n772), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n773), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n774), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n775), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n776), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n777), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n778), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n779), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n780), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n781), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n782), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n783), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n784), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n785), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n786), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n787), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n788), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n789), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n790), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n791), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n792), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n793), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n794), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n795), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n796), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n797), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n798), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n799), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n800), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n801), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n802), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n803), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n804), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n805), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n806), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n807), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n808), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n809), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n810), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n811), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n812), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n813), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n814), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n815), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n816), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n817), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n818), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n819), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n820), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n821), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n822), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n823), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n824), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n852), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n853), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n854), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n855), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n856), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n857), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n858), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n859), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n860), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n861), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n862), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n863), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n864), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n865), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n866), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n867), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n868), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n869), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n870), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n871), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n872), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n873), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n874), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n875), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n876), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n877), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n878), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n879), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n880), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n881), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n882), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n883), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n884), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n885), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n886), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n887), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n888), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n889), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n890), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n891), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n892), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n893), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n894), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n895), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n896), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n897), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n898), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n899), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n900), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n901), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n902), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n903), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n904), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n905), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n906), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n907), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n908), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n909), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n910), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n911), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n912), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n913), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n914), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n915), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  CLKBUF_X1 U3 ( .A(N10), .Z(n622) );
  BUF_X1 U4 ( .A(n621), .Z(n613) );
  INV_X2 U5 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U6 ( .A(n622), .Z(n618) );
  BUF_X1 U7 ( .A(n622), .Z(n619) );
  BUF_X1 U8 ( .A(n622), .Z(n620) );
  BUF_X1 U9 ( .A(n621), .Z(n615) );
  BUF_X1 U10 ( .A(n621), .Z(n614) );
  BUF_X1 U11 ( .A(n621), .Z(n616) );
  BUF_X1 U12 ( .A(n621), .Z(n617) );
  BUF_X1 U13 ( .A(N11), .Z(n611) );
  BUF_X1 U14 ( .A(N11), .Z(n612) );
  BUF_X1 U15 ( .A(N10), .Z(n621) );
  NOR3_X1 U16 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1207) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(n623), .ZN(n1196) );
  NOR3_X1 U18 ( .A1(N10), .A2(N12), .A3(n624), .ZN(n1186) );
  NOR3_X1 U19 ( .A1(n623), .A2(N12), .A3(n624), .ZN(n1176) );
  INV_X1 U20 ( .A(n1133), .ZN(n848) );
  INV_X1 U21 ( .A(n1123), .ZN(n847) );
  INV_X1 U22 ( .A(n1114), .ZN(n846) );
  INV_X1 U23 ( .A(n1105), .ZN(n845) );
  INV_X1 U24 ( .A(n1060), .ZN(n840) );
  INV_X1 U25 ( .A(n1050), .ZN(n839) );
  INV_X1 U26 ( .A(n1041), .ZN(n838) );
  INV_X1 U27 ( .A(n1032), .ZN(n837) );
  INV_X1 U28 ( .A(n987), .ZN(n832) );
  INV_X1 U29 ( .A(n977), .ZN(n831) );
  INV_X1 U30 ( .A(n968), .ZN(n830) );
  INV_X1 U31 ( .A(n959), .ZN(n829) );
  INV_X1 U32 ( .A(n1096), .ZN(n844) );
  INV_X1 U33 ( .A(n1087), .ZN(n843) );
  INV_X1 U34 ( .A(n1078), .ZN(n842) );
  INV_X1 U35 ( .A(n1069), .ZN(n841) );
  INV_X1 U36 ( .A(n950), .ZN(n828) );
  INV_X1 U37 ( .A(n941), .ZN(n827) );
  INV_X1 U38 ( .A(n932), .ZN(n826) );
  INV_X1 U39 ( .A(n923), .ZN(n825) );
  INV_X1 U40 ( .A(n1023), .ZN(n836) );
  INV_X1 U41 ( .A(n1014), .ZN(n835) );
  INV_X1 U42 ( .A(n1005), .ZN(n834) );
  INV_X1 U43 ( .A(n996), .ZN(n833) );
  BUF_X1 U44 ( .A(N12), .Z(n608) );
  BUF_X1 U45 ( .A(N12), .Z(n609) );
  INV_X1 U46 ( .A(N13), .ZN(n850) );
  AND3_X1 U47 ( .A1(n623), .A2(n624), .A3(N12), .ZN(n1166) );
  AND3_X1 U48 ( .A1(N10), .A2(n624), .A3(N12), .ZN(n1156) );
  AND3_X1 U49 ( .A1(N11), .A2(n623), .A3(N12), .ZN(n1146) );
  AND3_X1 U50 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1136) );
  INV_X1 U51 ( .A(N14), .ZN(n851) );
  NAND2_X1 U52 ( .A1(n1196), .A2(n1206), .ZN(n1205) );
  NAND2_X1 U53 ( .A1(n1186), .A2(n1206), .ZN(n1195) );
  NAND2_X1 U54 ( .A1(n1176), .A2(n1206), .ZN(n1185) );
  NAND2_X1 U55 ( .A1(n1166), .A2(n1206), .ZN(n1175) );
  NAND2_X1 U56 ( .A1(n1156), .A2(n1206), .ZN(n1165) );
  NAND2_X1 U57 ( .A1(n1146), .A2(n1206), .ZN(n1155) );
  NAND2_X1 U58 ( .A1(n1136), .A2(n1206), .ZN(n1145) );
  NAND2_X1 U59 ( .A1(n1207), .A2(n1206), .ZN(n1216) );
  NAND2_X1 U60 ( .A1(n1125), .A2(n1207), .ZN(n1133) );
  NAND2_X1 U61 ( .A1(n1125), .A2(n1196), .ZN(n1123) );
  NAND2_X1 U62 ( .A1(n1125), .A2(n1186), .ZN(n1114) );
  NAND2_X1 U63 ( .A1(n1125), .A2(n1176), .ZN(n1105) );
  NAND2_X1 U64 ( .A1(n1052), .A2(n1207), .ZN(n1060) );
  NAND2_X1 U65 ( .A1(n1052), .A2(n1196), .ZN(n1050) );
  NAND2_X1 U66 ( .A1(n1052), .A2(n1186), .ZN(n1041) );
  NAND2_X1 U67 ( .A1(n1052), .A2(n1176), .ZN(n1032) );
  NAND2_X1 U68 ( .A1(n979), .A2(n1207), .ZN(n987) );
  NAND2_X1 U69 ( .A1(n979), .A2(n1196), .ZN(n977) );
  NAND2_X1 U70 ( .A1(n979), .A2(n1186), .ZN(n968) );
  NAND2_X1 U71 ( .A1(n979), .A2(n1176), .ZN(n959) );
  NAND2_X1 U72 ( .A1(n1125), .A2(n1166), .ZN(n1096) );
  NAND2_X1 U73 ( .A1(n1125), .A2(n1156), .ZN(n1087) );
  NAND2_X1 U74 ( .A1(n1125), .A2(n1146), .ZN(n1078) );
  NAND2_X1 U75 ( .A1(n1125), .A2(n1136), .ZN(n1069) );
  NAND2_X1 U76 ( .A1(n1052), .A2(n1166), .ZN(n1023) );
  NAND2_X1 U77 ( .A1(n1052), .A2(n1156), .ZN(n1014) );
  NAND2_X1 U78 ( .A1(n1052), .A2(n1146), .ZN(n1005) );
  NAND2_X1 U79 ( .A1(n1052), .A2(n1136), .ZN(n996) );
  NAND2_X1 U80 ( .A1(n979), .A2(n1166), .ZN(n950) );
  NAND2_X1 U81 ( .A1(n979), .A2(n1156), .ZN(n941) );
  NAND2_X1 U82 ( .A1(n979), .A2(n1146), .ZN(n932) );
  NAND2_X1 U83 ( .A1(n979), .A2(n1136), .ZN(n923) );
  AND3_X1 U84 ( .A1(n850), .A2(n851), .A3(n1135), .ZN(n1206) );
  AND3_X1 U85 ( .A1(N13), .A2(n1135), .A3(N14), .ZN(n979) );
  AND3_X1 U86 ( .A1(n1135), .A2(n851), .A3(N13), .ZN(n1125) );
  AND3_X1 U87 ( .A1(n1135), .A2(n850), .A3(N14), .ZN(n1052) );
  NOR2_X1 U88 ( .A1(n849), .A2(addr[5]), .ZN(n1135) );
  INV_X1 U89 ( .A(wr_en), .ZN(n849) );
  OAI21_X1 U90 ( .B1(n625), .B2(n1175), .A(n1174), .ZN(n883) );
  NAND2_X1 U91 ( .A1(\mem[4][0] ), .A2(n1175), .ZN(n1174) );
  OAI21_X1 U92 ( .B1(n626), .B2(n1175), .A(n1173), .ZN(n882) );
  NAND2_X1 U93 ( .A1(\mem[4][1] ), .A2(n1175), .ZN(n1173) );
  OAI21_X1 U94 ( .B1(n627), .B2(n1175), .A(n1172), .ZN(n881) );
  NAND2_X1 U95 ( .A1(\mem[4][2] ), .A2(n1175), .ZN(n1172) );
  OAI21_X1 U96 ( .B1(n628), .B2(n1175), .A(n1171), .ZN(n880) );
  NAND2_X1 U97 ( .A1(\mem[4][3] ), .A2(n1175), .ZN(n1171) );
  OAI21_X1 U98 ( .B1(n629), .B2(n1175), .A(n1170), .ZN(n879) );
  NAND2_X1 U99 ( .A1(\mem[4][4] ), .A2(n1175), .ZN(n1170) );
  OAI21_X1 U100 ( .B1(n630), .B2(n1175), .A(n1169), .ZN(n878) );
  NAND2_X1 U101 ( .A1(\mem[4][5] ), .A2(n1175), .ZN(n1169) );
  OAI21_X1 U102 ( .B1(n631), .B2(n1175), .A(n1168), .ZN(n877) );
  NAND2_X1 U103 ( .A1(\mem[4][6] ), .A2(n1175), .ZN(n1168) );
  OAI21_X1 U104 ( .B1(n632), .B2(n1175), .A(n1167), .ZN(n876) );
  NAND2_X1 U105 ( .A1(\mem[4][7] ), .A2(n1175), .ZN(n1167) );
  OAI21_X1 U106 ( .B1(n625), .B2(n1155), .A(n1154), .ZN(n867) );
  NAND2_X1 U107 ( .A1(\mem[6][0] ), .A2(n1155), .ZN(n1154) );
  OAI21_X1 U108 ( .B1(n626), .B2(n1155), .A(n1153), .ZN(n866) );
  NAND2_X1 U109 ( .A1(\mem[6][1] ), .A2(n1155), .ZN(n1153) );
  OAI21_X1 U110 ( .B1(n627), .B2(n1155), .A(n1152), .ZN(n865) );
  NAND2_X1 U111 ( .A1(\mem[6][2] ), .A2(n1155), .ZN(n1152) );
  OAI21_X1 U112 ( .B1(n628), .B2(n1155), .A(n1151), .ZN(n864) );
  NAND2_X1 U113 ( .A1(\mem[6][3] ), .A2(n1155), .ZN(n1151) );
  OAI21_X1 U114 ( .B1(n629), .B2(n1155), .A(n1150), .ZN(n863) );
  NAND2_X1 U115 ( .A1(\mem[6][4] ), .A2(n1155), .ZN(n1150) );
  OAI21_X1 U116 ( .B1(n630), .B2(n1155), .A(n1149), .ZN(n862) );
  NAND2_X1 U117 ( .A1(\mem[6][5] ), .A2(n1155), .ZN(n1149) );
  OAI21_X1 U118 ( .B1(n631), .B2(n1155), .A(n1148), .ZN(n861) );
  NAND2_X1 U119 ( .A1(\mem[6][6] ), .A2(n1155), .ZN(n1148) );
  OAI21_X1 U120 ( .B1(n632), .B2(n1155), .A(n1147), .ZN(n860) );
  NAND2_X1 U121 ( .A1(\mem[6][7] ), .A2(n1155), .ZN(n1147) );
  OAI21_X1 U122 ( .B1(n625), .B2(n1145), .A(n1144), .ZN(n859) );
  NAND2_X1 U123 ( .A1(\mem[7][0] ), .A2(n1145), .ZN(n1144) );
  OAI21_X1 U124 ( .B1(n626), .B2(n1145), .A(n1143), .ZN(n858) );
  NAND2_X1 U125 ( .A1(\mem[7][1] ), .A2(n1145), .ZN(n1143) );
  OAI21_X1 U126 ( .B1(n627), .B2(n1145), .A(n1142), .ZN(n857) );
  NAND2_X1 U127 ( .A1(\mem[7][2] ), .A2(n1145), .ZN(n1142) );
  OAI21_X1 U128 ( .B1(n628), .B2(n1145), .A(n1141), .ZN(n856) );
  NAND2_X1 U129 ( .A1(\mem[7][3] ), .A2(n1145), .ZN(n1141) );
  OAI21_X1 U130 ( .B1(n629), .B2(n1145), .A(n1140), .ZN(n855) );
  NAND2_X1 U131 ( .A1(\mem[7][4] ), .A2(n1145), .ZN(n1140) );
  OAI21_X1 U132 ( .B1(n630), .B2(n1145), .A(n1139), .ZN(n854) );
  NAND2_X1 U133 ( .A1(\mem[7][5] ), .A2(n1145), .ZN(n1139) );
  OAI21_X1 U134 ( .B1(n631), .B2(n1145), .A(n1138), .ZN(n853) );
  NAND2_X1 U135 ( .A1(\mem[7][6] ), .A2(n1145), .ZN(n1138) );
  OAI21_X1 U136 ( .B1(n632), .B2(n1145), .A(n1137), .ZN(n852) );
  NAND2_X1 U137 ( .A1(\mem[7][7] ), .A2(n1145), .ZN(n1137) );
  OAI21_X1 U138 ( .B1(n625), .B2(n1205), .A(n1204), .ZN(n907) );
  NAND2_X1 U139 ( .A1(\mem[1][0] ), .A2(n1205), .ZN(n1204) );
  OAI21_X1 U140 ( .B1(n626), .B2(n1205), .A(n1203), .ZN(n906) );
  NAND2_X1 U141 ( .A1(\mem[1][1] ), .A2(n1205), .ZN(n1203) );
  OAI21_X1 U142 ( .B1(n627), .B2(n1205), .A(n1202), .ZN(n905) );
  NAND2_X1 U143 ( .A1(\mem[1][2] ), .A2(n1205), .ZN(n1202) );
  OAI21_X1 U144 ( .B1(n628), .B2(n1205), .A(n1201), .ZN(n904) );
  NAND2_X1 U145 ( .A1(\mem[1][3] ), .A2(n1205), .ZN(n1201) );
  OAI21_X1 U146 ( .B1(n629), .B2(n1205), .A(n1200), .ZN(n903) );
  NAND2_X1 U147 ( .A1(\mem[1][4] ), .A2(n1205), .ZN(n1200) );
  OAI21_X1 U148 ( .B1(n630), .B2(n1205), .A(n1199), .ZN(n902) );
  NAND2_X1 U149 ( .A1(\mem[1][5] ), .A2(n1205), .ZN(n1199) );
  OAI21_X1 U150 ( .B1(n631), .B2(n1205), .A(n1198), .ZN(n901) );
  NAND2_X1 U151 ( .A1(\mem[1][6] ), .A2(n1205), .ZN(n1198) );
  OAI21_X1 U152 ( .B1(n632), .B2(n1205), .A(n1197), .ZN(n900) );
  NAND2_X1 U153 ( .A1(\mem[1][7] ), .A2(n1205), .ZN(n1197) );
  OAI21_X1 U154 ( .B1(n625), .B2(n1195), .A(n1194), .ZN(n899) );
  NAND2_X1 U155 ( .A1(\mem[2][0] ), .A2(n1195), .ZN(n1194) );
  OAI21_X1 U156 ( .B1(n626), .B2(n1195), .A(n1193), .ZN(n898) );
  NAND2_X1 U157 ( .A1(\mem[2][1] ), .A2(n1195), .ZN(n1193) );
  OAI21_X1 U158 ( .B1(n627), .B2(n1195), .A(n1192), .ZN(n897) );
  NAND2_X1 U159 ( .A1(\mem[2][2] ), .A2(n1195), .ZN(n1192) );
  OAI21_X1 U160 ( .B1(n628), .B2(n1195), .A(n1191), .ZN(n896) );
  NAND2_X1 U161 ( .A1(\mem[2][3] ), .A2(n1195), .ZN(n1191) );
  OAI21_X1 U162 ( .B1(n629), .B2(n1195), .A(n1190), .ZN(n895) );
  NAND2_X1 U163 ( .A1(\mem[2][4] ), .A2(n1195), .ZN(n1190) );
  OAI21_X1 U164 ( .B1(n630), .B2(n1195), .A(n1189), .ZN(n894) );
  NAND2_X1 U165 ( .A1(\mem[2][5] ), .A2(n1195), .ZN(n1189) );
  OAI21_X1 U166 ( .B1(n631), .B2(n1195), .A(n1188), .ZN(n893) );
  NAND2_X1 U167 ( .A1(\mem[2][6] ), .A2(n1195), .ZN(n1188) );
  OAI21_X1 U168 ( .B1(n632), .B2(n1195), .A(n1187), .ZN(n892) );
  NAND2_X1 U169 ( .A1(\mem[2][7] ), .A2(n1195), .ZN(n1187) );
  OAI21_X1 U170 ( .B1(n625), .B2(n1185), .A(n1184), .ZN(n891) );
  NAND2_X1 U171 ( .A1(\mem[3][0] ), .A2(n1185), .ZN(n1184) );
  OAI21_X1 U172 ( .B1(n626), .B2(n1185), .A(n1183), .ZN(n890) );
  NAND2_X1 U173 ( .A1(\mem[3][1] ), .A2(n1185), .ZN(n1183) );
  OAI21_X1 U174 ( .B1(n627), .B2(n1185), .A(n1182), .ZN(n889) );
  NAND2_X1 U175 ( .A1(\mem[3][2] ), .A2(n1185), .ZN(n1182) );
  OAI21_X1 U176 ( .B1(n628), .B2(n1185), .A(n1181), .ZN(n888) );
  NAND2_X1 U177 ( .A1(\mem[3][3] ), .A2(n1185), .ZN(n1181) );
  OAI21_X1 U178 ( .B1(n629), .B2(n1185), .A(n1180), .ZN(n887) );
  NAND2_X1 U179 ( .A1(\mem[3][4] ), .A2(n1185), .ZN(n1180) );
  OAI21_X1 U180 ( .B1(n630), .B2(n1185), .A(n1179), .ZN(n886) );
  NAND2_X1 U181 ( .A1(\mem[3][5] ), .A2(n1185), .ZN(n1179) );
  OAI21_X1 U182 ( .B1(n631), .B2(n1185), .A(n1178), .ZN(n885) );
  NAND2_X1 U183 ( .A1(\mem[3][6] ), .A2(n1185), .ZN(n1178) );
  OAI21_X1 U184 ( .B1(n632), .B2(n1185), .A(n1177), .ZN(n884) );
  NAND2_X1 U185 ( .A1(\mem[3][7] ), .A2(n1185), .ZN(n1177) );
  OAI21_X1 U186 ( .B1(n625), .B2(n1165), .A(n1164), .ZN(n875) );
  NAND2_X1 U187 ( .A1(\mem[5][0] ), .A2(n1165), .ZN(n1164) );
  OAI21_X1 U188 ( .B1(n626), .B2(n1165), .A(n1163), .ZN(n874) );
  NAND2_X1 U189 ( .A1(\mem[5][1] ), .A2(n1165), .ZN(n1163) );
  OAI21_X1 U190 ( .B1(n627), .B2(n1165), .A(n1162), .ZN(n873) );
  NAND2_X1 U191 ( .A1(\mem[5][2] ), .A2(n1165), .ZN(n1162) );
  OAI21_X1 U192 ( .B1(n628), .B2(n1165), .A(n1161), .ZN(n872) );
  NAND2_X1 U193 ( .A1(\mem[5][3] ), .A2(n1165), .ZN(n1161) );
  OAI21_X1 U194 ( .B1(n629), .B2(n1165), .A(n1160), .ZN(n871) );
  NAND2_X1 U195 ( .A1(\mem[5][4] ), .A2(n1165), .ZN(n1160) );
  OAI21_X1 U196 ( .B1(n630), .B2(n1165), .A(n1159), .ZN(n870) );
  NAND2_X1 U197 ( .A1(\mem[5][5] ), .A2(n1165), .ZN(n1159) );
  OAI21_X1 U198 ( .B1(n631), .B2(n1165), .A(n1158), .ZN(n869) );
  NAND2_X1 U199 ( .A1(\mem[5][6] ), .A2(n1165), .ZN(n1158) );
  OAI21_X1 U200 ( .B1(n632), .B2(n1165), .A(n1157), .ZN(n868) );
  NAND2_X1 U201 ( .A1(\mem[5][7] ), .A2(n1165), .ZN(n1157) );
  OAI21_X1 U202 ( .B1(n1216), .B2(n625), .A(n1215), .ZN(n915) );
  NAND2_X1 U203 ( .A1(\mem[0][0] ), .A2(n1216), .ZN(n1215) );
  OAI21_X1 U204 ( .B1(n1216), .B2(n626), .A(n1214), .ZN(n914) );
  NAND2_X1 U205 ( .A1(\mem[0][1] ), .A2(n1216), .ZN(n1214) );
  OAI21_X1 U206 ( .B1(n1216), .B2(n627), .A(n1213), .ZN(n913) );
  NAND2_X1 U207 ( .A1(\mem[0][2] ), .A2(n1216), .ZN(n1213) );
  OAI21_X1 U208 ( .B1(n1216), .B2(n628), .A(n1212), .ZN(n912) );
  NAND2_X1 U209 ( .A1(\mem[0][3] ), .A2(n1216), .ZN(n1212) );
  OAI21_X1 U210 ( .B1(n1216), .B2(n629), .A(n1211), .ZN(n911) );
  NAND2_X1 U211 ( .A1(\mem[0][4] ), .A2(n1216), .ZN(n1211) );
  OAI21_X1 U212 ( .B1(n1216), .B2(n630), .A(n1210), .ZN(n910) );
  NAND2_X1 U213 ( .A1(\mem[0][5] ), .A2(n1216), .ZN(n1210) );
  OAI21_X1 U214 ( .B1(n1216), .B2(n631), .A(n1209), .ZN(n909) );
  NAND2_X1 U215 ( .A1(\mem[0][6] ), .A2(n1216), .ZN(n1209) );
  OAI21_X1 U216 ( .B1(n1216), .B2(n632), .A(n1208), .ZN(n908) );
  NAND2_X1 U217 ( .A1(\mem[0][7] ), .A2(n1216), .ZN(n1208) );
  INV_X1 U218 ( .A(n1134), .ZN(n824) );
  AOI22_X1 U219 ( .A1(data_in[0]), .A2(n848), .B1(n1133), .B2(\mem[8][0] ), 
        .ZN(n1134) );
  INV_X1 U220 ( .A(n1132), .ZN(n823) );
  AOI22_X1 U221 ( .A1(data_in[1]), .A2(n848), .B1(n1133), .B2(\mem[8][1] ), 
        .ZN(n1132) );
  INV_X1 U222 ( .A(n1131), .ZN(n822) );
  AOI22_X1 U223 ( .A1(data_in[2]), .A2(n848), .B1(n1133), .B2(\mem[8][2] ), 
        .ZN(n1131) );
  INV_X1 U224 ( .A(n1130), .ZN(n821) );
  AOI22_X1 U225 ( .A1(data_in[3]), .A2(n848), .B1(n1133), .B2(\mem[8][3] ), 
        .ZN(n1130) );
  INV_X1 U226 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U227 ( .A1(data_in[4]), .A2(n848), .B1(n1133), .B2(\mem[8][4] ), 
        .ZN(n1129) );
  INV_X1 U228 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U229 ( .A1(data_in[5]), .A2(n848), .B1(n1133), .B2(\mem[8][5] ), 
        .ZN(n1128) );
  INV_X1 U230 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U231 ( .A1(data_in[6]), .A2(n848), .B1(n1133), .B2(\mem[8][6] ), 
        .ZN(n1127) );
  INV_X1 U232 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n848), .B1(n1133), .B2(\mem[8][7] ), 
        .ZN(n1126) );
  INV_X1 U234 ( .A(n1124), .ZN(n816) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n847), .B1(n1123), .B2(\mem[9][0] ), 
        .ZN(n1124) );
  INV_X1 U236 ( .A(n1122), .ZN(n815) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n847), .B1(n1123), .B2(\mem[9][1] ), 
        .ZN(n1122) );
  INV_X1 U238 ( .A(n1121), .ZN(n814) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n847), .B1(n1123), .B2(\mem[9][2] ), 
        .ZN(n1121) );
  INV_X1 U240 ( .A(n1120), .ZN(n813) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n847), .B1(n1123), .B2(\mem[9][3] ), 
        .ZN(n1120) );
  INV_X1 U242 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n847), .B1(n1123), .B2(\mem[9][4] ), 
        .ZN(n1119) );
  INV_X1 U244 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n847), .B1(n1123), .B2(\mem[9][5] ), 
        .ZN(n1118) );
  INV_X1 U246 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n847), .B1(n1123), .B2(\mem[9][6] ), 
        .ZN(n1117) );
  INV_X1 U248 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n847), .B1(n1123), .B2(\mem[9][7] ), 
        .ZN(n1116) );
  INV_X1 U250 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n846), .B1(n1114), .B2(\mem[10][0] ), 
        .ZN(n1115) );
  INV_X1 U252 ( .A(n1113), .ZN(n807) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n846), .B1(n1114), .B2(\mem[10][1] ), 
        .ZN(n1113) );
  INV_X1 U254 ( .A(n1112), .ZN(n806) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n846), .B1(n1114), .B2(\mem[10][2] ), 
        .ZN(n1112) );
  INV_X1 U256 ( .A(n1111), .ZN(n805) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n846), .B1(n1114), .B2(\mem[10][3] ), 
        .ZN(n1111) );
  INV_X1 U258 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n846), .B1(n1114), .B2(\mem[10][4] ), 
        .ZN(n1110) );
  INV_X1 U260 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n846), .B1(n1114), .B2(\mem[10][5] ), 
        .ZN(n1109) );
  INV_X1 U262 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n846), .B1(n1114), .B2(\mem[10][6] ), 
        .ZN(n1108) );
  INV_X1 U264 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n846), .B1(n1114), .B2(\mem[10][7] ), 
        .ZN(n1107) );
  INV_X1 U266 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n845), .B1(n1105), .B2(\mem[11][0] ), 
        .ZN(n1106) );
  INV_X1 U268 ( .A(n1104), .ZN(n799) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n845), .B1(n1105), .B2(\mem[11][1] ), 
        .ZN(n1104) );
  INV_X1 U270 ( .A(n1103), .ZN(n798) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n845), .B1(n1105), .B2(\mem[11][2] ), 
        .ZN(n1103) );
  INV_X1 U272 ( .A(n1102), .ZN(n797) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n845), .B1(n1105), .B2(\mem[11][3] ), 
        .ZN(n1102) );
  INV_X1 U274 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n845), .B1(n1105), .B2(\mem[11][4] ), 
        .ZN(n1101) );
  INV_X1 U276 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n845), .B1(n1105), .B2(\mem[11][5] ), 
        .ZN(n1100) );
  INV_X1 U278 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n845), .B1(n1105), .B2(\mem[11][6] ), 
        .ZN(n1099) );
  INV_X1 U280 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n845), .B1(n1105), .B2(\mem[11][7] ), 
        .ZN(n1098) );
  INV_X1 U282 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n844), .B1(n1096), .B2(\mem[12][0] ), 
        .ZN(n1097) );
  INV_X1 U284 ( .A(n1095), .ZN(n791) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n844), .B1(n1096), .B2(\mem[12][1] ), 
        .ZN(n1095) );
  INV_X1 U286 ( .A(n1094), .ZN(n790) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n844), .B1(n1096), .B2(\mem[12][2] ), 
        .ZN(n1094) );
  INV_X1 U288 ( .A(n1093), .ZN(n789) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n844), .B1(n1096), .B2(\mem[12][3] ), 
        .ZN(n1093) );
  INV_X1 U290 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n844), .B1(n1096), .B2(\mem[12][4] ), 
        .ZN(n1092) );
  INV_X1 U292 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n844), .B1(n1096), .B2(\mem[12][5] ), 
        .ZN(n1091) );
  INV_X1 U294 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n844), .B1(n1096), .B2(\mem[12][6] ), 
        .ZN(n1090) );
  INV_X1 U296 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n844), .B1(n1096), .B2(\mem[12][7] ), 
        .ZN(n1089) );
  INV_X1 U298 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n843), .B1(n1087), .B2(\mem[13][0] ), 
        .ZN(n1088) );
  INV_X1 U300 ( .A(n1086), .ZN(n783) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n843), .B1(n1087), .B2(\mem[13][1] ), 
        .ZN(n1086) );
  INV_X1 U302 ( .A(n1085), .ZN(n782) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n843), .B1(n1087), .B2(\mem[13][2] ), 
        .ZN(n1085) );
  INV_X1 U304 ( .A(n1084), .ZN(n781) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n843), .B1(n1087), .B2(\mem[13][3] ), 
        .ZN(n1084) );
  INV_X1 U306 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n843), .B1(n1087), .B2(\mem[13][4] ), 
        .ZN(n1083) );
  INV_X1 U308 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n843), .B1(n1087), .B2(\mem[13][5] ), 
        .ZN(n1082) );
  INV_X1 U310 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n843), .B1(n1087), .B2(\mem[13][6] ), 
        .ZN(n1081) );
  INV_X1 U312 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n843), .B1(n1087), .B2(\mem[13][7] ), 
        .ZN(n1080) );
  INV_X1 U314 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n842), .B1(n1078), .B2(\mem[14][0] ), 
        .ZN(n1079) );
  INV_X1 U316 ( .A(n1077), .ZN(n775) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n842), .B1(n1078), .B2(\mem[14][1] ), 
        .ZN(n1077) );
  INV_X1 U318 ( .A(n1076), .ZN(n774) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n842), .B1(n1078), .B2(\mem[14][2] ), 
        .ZN(n1076) );
  INV_X1 U320 ( .A(n1075), .ZN(n773) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n842), .B1(n1078), .B2(\mem[14][3] ), 
        .ZN(n1075) );
  INV_X1 U322 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n842), .B1(n1078), .B2(\mem[14][4] ), 
        .ZN(n1074) );
  INV_X1 U324 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n842), .B1(n1078), .B2(\mem[14][5] ), 
        .ZN(n1073) );
  INV_X1 U326 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n842), .B1(n1078), .B2(\mem[14][6] ), 
        .ZN(n1072) );
  INV_X1 U328 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n842), .B1(n1078), .B2(\mem[14][7] ), 
        .ZN(n1071) );
  INV_X1 U330 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U331 ( .A1(data_in[0]), .A2(n841), .B1(n1069), .B2(\mem[15][0] ), 
        .ZN(n1070) );
  INV_X1 U332 ( .A(n1068), .ZN(n767) );
  AOI22_X1 U333 ( .A1(data_in[1]), .A2(n841), .B1(n1069), .B2(\mem[15][1] ), 
        .ZN(n1068) );
  INV_X1 U334 ( .A(n1067), .ZN(n766) );
  AOI22_X1 U335 ( .A1(data_in[2]), .A2(n841), .B1(n1069), .B2(\mem[15][2] ), 
        .ZN(n1067) );
  INV_X1 U336 ( .A(n1066), .ZN(n765) );
  AOI22_X1 U337 ( .A1(data_in[3]), .A2(n841), .B1(n1069), .B2(\mem[15][3] ), 
        .ZN(n1066) );
  INV_X1 U338 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U339 ( .A1(data_in[4]), .A2(n841), .B1(n1069), .B2(\mem[15][4] ), 
        .ZN(n1065) );
  INV_X1 U340 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U341 ( .A1(data_in[5]), .A2(n841), .B1(n1069), .B2(\mem[15][5] ), 
        .ZN(n1064) );
  INV_X1 U342 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U343 ( .A1(data_in[6]), .A2(n841), .B1(n1069), .B2(\mem[15][6] ), 
        .ZN(n1063) );
  INV_X1 U344 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U345 ( .A1(data_in[7]), .A2(n841), .B1(n1069), .B2(\mem[15][7] ), 
        .ZN(n1062) );
  INV_X1 U346 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U347 ( .A1(data_in[0]), .A2(n840), .B1(n1060), .B2(\mem[16][0] ), 
        .ZN(n1061) );
  INV_X1 U348 ( .A(n1059), .ZN(n759) );
  AOI22_X1 U349 ( .A1(data_in[1]), .A2(n840), .B1(n1060), .B2(\mem[16][1] ), 
        .ZN(n1059) );
  INV_X1 U350 ( .A(n1058), .ZN(n758) );
  AOI22_X1 U351 ( .A1(data_in[2]), .A2(n840), .B1(n1060), .B2(\mem[16][2] ), 
        .ZN(n1058) );
  INV_X1 U352 ( .A(n1057), .ZN(n757) );
  AOI22_X1 U353 ( .A1(data_in[3]), .A2(n840), .B1(n1060), .B2(\mem[16][3] ), 
        .ZN(n1057) );
  INV_X1 U354 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U355 ( .A1(data_in[4]), .A2(n840), .B1(n1060), .B2(\mem[16][4] ), 
        .ZN(n1056) );
  INV_X1 U356 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U357 ( .A1(data_in[5]), .A2(n840), .B1(n1060), .B2(\mem[16][5] ), 
        .ZN(n1055) );
  INV_X1 U358 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U359 ( .A1(data_in[6]), .A2(n840), .B1(n1060), .B2(\mem[16][6] ), 
        .ZN(n1054) );
  INV_X1 U360 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U361 ( .A1(data_in[7]), .A2(n840), .B1(n1060), .B2(\mem[16][7] ), 
        .ZN(n1053) );
  INV_X1 U362 ( .A(n1051), .ZN(n752) );
  AOI22_X1 U363 ( .A1(data_in[0]), .A2(n839), .B1(n1050), .B2(\mem[17][0] ), 
        .ZN(n1051) );
  INV_X1 U364 ( .A(n1049), .ZN(n751) );
  AOI22_X1 U365 ( .A1(data_in[1]), .A2(n839), .B1(n1050), .B2(\mem[17][1] ), 
        .ZN(n1049) );
  INV_X1 U366 ( .A(n1048), .ZN(n750) );
  AOI22_X1 U367 ( .A1(data_in[2]), .A2(n839), .B1(n1050), .B2(\mem[17][2] ), 
        .ZN(n1048) );
  INV_X1 U368 ( .A(n1047), .ZN(n749) );
  AOI22_X1 U369 ( .A1(data_in[3]), .A2(n839), .B1(n1050), .B2(\mem[17][3] ), 
        .ZN(n1047) );
  INV_X1 U370 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U371 ( .A1(data_in[4]), .A2(n839), .B1(n1050), .B2(\mem[17][4] ), 
        .ZN(n1046) );
  INV_X1 U372 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U373 ( .A1(data_in[5]), .A2(n839), .B1(n1050), .B2(\mem[17][5] ), 
        .ZN(n1045) );
  INV_X1 U374 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U375 ( .A1(data_in[6]), .A2(n839), .B1(n1050), .B2(\mem[17][6] ), 
        .ZN(n1044) );
  INV_X1 U376 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U377 ( .A1(data_in[7]), .A2(n839), .B1(n1050), .B2(\mem[17][7] ), 
        .ZN(n1043) );
  INV_X1 U378 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U379 ( .A1(data_in[0]), .A2(n838), .B1(n1041), .B2(\mem[18][0] ), 
        .ZN(n1042) );
  INV_X1 U380 ( .A(n1040), .ZN(n743) );
  AOI22_X1 U381 ( .A1(data_in[1]), .A2(n838), .B1(n1041), .B2(\mem[18][1] ), 
        .ZN(n1040) );
  INV_X1 U382 ( .A(n1039), .ZN(n742) );
  AOI22_X1 U383 ( .A1(data_in[2]), .A2(n838), .B1(n1041), .B2(\mem[18][2] ), 
        .ZN(n1039) );
  INV_X1 U384 ( .A(n1038), .ZN(n741) );
  AOI22_X1 U385 ( .A1(data_in[3]), .A2(n838), .B1(n1041), .B2(\mem[18][3] ), 
        .ZN(n1038) );
  INV_X1 U386 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U387 ( .A1(data_in[4]), .A2(n838), .B1(n1041), .B2(\mem[18][4] ), 
        .ZN(n1037) );
  INV_X1 U388 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U389 ( .A1(data_in[5]), .A2(n838), .B1(n1041), .B2(\mem[18][5] ), 
        .ZN(n1036) );
  INV_X1 U390 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U391 ( .A1(data_in[6]), .A2(n838), .B1(n1041), .B2(\mem[18][6] ), 
        .ZN(n1035) );
  INV_X1 U392 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U393 ( .A1(data_in[7]), .A2(n838), .B1(n1041), .B2(\mem[18][7] ), 
        .ZN(n1034) );
  INV_X1 U394 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U395 ( .A1(data_in[0]), .A2(n837), .B1(n1032), .B2(\mem[19][0] ), 
        .ZN(n1033) );
  INV_X1 U396 ( .A(n1031), .ZN(n735) );
  AOI22_X1 U397 ( .A1(data_in[1]), .A2(n837), .B1(n1032), .B2(\mem[19][1] ), 
        .ZN(n1031) );
  INV_X1 U398 ( .A(n1030), .ZN(n734) );
  AOI22_X1 U399 ( .A1(data_in[2]), .A2(n837), .B1(n1032), .B2(\mem[19][2] ), 
        .ZN(n1030) );
  INV_X1 U400 ( .A(n1029), .ZN(n733) );
  AOI22_X1 U401 ( .A1(data_in[3]), .A2(n837), .B1(n1032), .B2(\mem[19][3] ), 
        .ZN(n1029) );
  INV_X1 U402 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U403 ( .A1(data_in[4]), .A2(n837), .B1(n1032), .B2(\mem[19][4] ), 
        .ZN(n1028) );
  INV_X1 U404 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U405 ( .A1(data_in[5]), .A2(n837), .B1(n1032), .B2(\mem[19][5] ), 
        .ZN(n1027) );
  INV_X1 U406 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U407 ( .A1(data_in[6]), .A2(n837), .B1(n1032), .B2(\mem[19][6] ), 
        .ZN(n1026) );
  INV_X1 U408 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U409 ( .A1(data_in[7]), .A2(n837), .B1(n1032), .B2(\mem[19][7] ), 
        .ZN(n1025) );
  INV_X1 U410 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U411 ( .A1(data_in[0]), .A2(n836), .B1(n1023), .B2(\mem[20][0] ), 
        .ZN(n1024) );
  INV_X1 U412 ( .A(n1022), .ZN(n727) );
  AOI22_X1 U413 ( .A1(data_in[1]), .A2(n836), .B1(n1023), .B2(\mem[20][1] ), 
        .ZN(n1022) );
  INV_X1 U414 ( .A(n1021), .ZN(n726) );
  AOI22_X1 U415 ( .A1(data_in[2]), .A2(n836), .B1(n1023), .B2(\mem[20][2] ), 
        .ZN(n1021) );
  INV_X1 U416 ( .A(n1020), .ZN(n725) );
  AOI22_X1 U417 ( .A1(data_in[3]), .A2(n836), .B1(n1023), .B2(\mem[20][3] ), 
        .ZN(n1020) );
  INV_X1 U418 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U419 ( .A1(data_in[4]), .A2(n836), .B1(n1023), .B2(\mem[20][4] ), 
        .ZN(n1019) );
  INV_X1 U420 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U421 ( .A1(data_in[5]), .A2(n836), .B1(n1023), .B2(\mem[20][5] ), 
        .ZN(n1018) );
  INV_X1 U422 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U423 ( .A1(data_in[6]), .A2(n836), .B1(n1023), .B2(\mem[20][6] ), 
        .ZN(n1017) );
  INV_X1 U424 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U425 ( .A1(data_in[7]), .A2(n836), .B1(n1023), .B2(\mem[20][7] ), 
        .ZN(n1016) );
  INV_X1 U426 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U427 ( .A1(data_in[0]), .A2(n835), .B1(n1014), .B2(\mem[21][0] ), 
        .ZN(n1015) );
  INV_X1 U428 ( .A(n1013), .ZN(n719) );
  AOI22_X1 U429 ( .A1(data_in[1]), .A2(n835), .B1(n1014), .B2(\mem[21][1] ), 
        .ZN(n1013) );
  INV_X1 U430 ( .A(n1012), .ZN(n718) );
  AOI22_X1 U431 ( .A1(data_in[2]), .A2(n835), .B1(n1014), .B2(\mem[21][2] ), 
        .ZN(n1012) );
  INV_X1 U432 ( .A(n1011), .ZN(n717) );
  AOI22_X1 U433 ( .A1(data_in[3]), .A2(n835), .B1(n1014), .B2(\mem[21][3] ), 
        .ZN(n1011) );
  INV_X1 U434 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U435 ( .A1(data_in[4]), .A2(n835), .B1(n1014), .B2(\mem[21][4] ), 
        .ZN(n1010) );
  INV_X1 U436 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U437 ( .A1(data_in[5]), .A2(n835), .B1(n1014), .B2(\mem[21][5] ), 
        .ZN(n1009) );
  INV_X1 U438 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U439 ( .A1(data_in[6]), .A2(n835), .B1(n1014), .B2(\mem[21][6] ), 
        .ZN(n1008) );
  INV_X1 U440 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U441 ( .A1(data_in[7]), .A2(n835), .B1(n1014), .B2(\mem[21][7] ), 
        .ZN(n1007) );
  INV_X1 U442 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U443 ( .A1(data_in[0]), .A2(n834), .B1(n1005), .B2(\mem[22][0] ), 
        .ZN(n1006) );
  INV_X1 U444 ( .A(n1004), .ZN(n711) );
  AOI22_X1 U445 ( .A1(data_in[1]), .A2(n834), .B1(n1005), .B2(\mem[22][1] ), 
        .ZN(n1004) );
  INV_X1 U446 ( .A(n1003), .ZN(n710) );
  AOI22_X1 U447 ( .A1(data_in[2]), .A2(n834), .B1(n1005), .B2(\mem[22][2] ), 
        .ZN(n1003) );
  INV_X1 U448 ( .A(n1002), .ZN(n709) );
  AOI22_X1 U449 ( .A1(data_in[3]), .A2(n834), .B1(n1005), .B2(\mem[22][3] ), 
        .ZN(n1002) );
  INV_X1 U450 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U451 ( .A1(data_in[4]), .A2(n834), .B1(n1005), .B2(\mem[22][4] ), 
        .ZN(n1001) );
  INV_X1 U452 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U453 ( .A1(data_in[5]), .A2(n834), .B1(n1005), .B2(\mem[22][5] ), 
        .ZN(n1000) );
  INV_X1 U454 ( .A(n999), .ZN(n706) );
  AOI22_X1 U455 ( .A1(data_in[6]), .A2(n834), .B1(n1005), .B2(\mem[22][6] ), 
        .ZN(n999) );
  INV_X1 U456 ( .A(n998), .ZN(n705) );
  AOI22_X1 U457 ( .A1(data_in[7]), .A2(n834), .B1(n1005), .B2(\mem[22][7] ), 
        .ZN(n998) );
  INV_X1 U458 ( .A(n997), .ZN(n704) );
  AOI22_X1 U459 ( .A1(data_in[0]), .A2(n833), .B1(n996), .B2(\mem[23][0] ), 
        .ZN(n997) );
  INV_X1 U460 ( .A(n995), .ZN(n703) );
  AOI22_X1 U461 ( .A1(data_in[1]), .A2(n833), .B1(n996), .B2(\mem[23][1] ), 
        .ZN(n995) );
  INV_X1 U462 ( .A(n994), .ZN(n702) );
  AOI22_X1 U463 ( .A1(data_in[2]), .A2(n833), .B1(n996), .B2(\mem[23][2] ), 
        .ZN(n994) );
  INV_X1 U464 ( .A(n993), .ZN(n701) );
  AOI22_X1 U465 ( .A1(data_in[3]), .A2(n833), .B1(n996), .B2(\mem[23][3] ), 
        .ZN(n993) );
  INV_X1 U466 ( .A(n992), .ZN(n700) );
  AOI22_X1 U467 ( .A1(data_in[4]), .A2(n833), .B1(n996), .B2(\mem[23][4] ), 
        .ZN(n992) );
  INV_X1 U468 ( .A(n991), .ZN(n699) );
  AOI22_X1 U469 ( .A1(data_in[5]), .A2(n833), .B1(n996), .B2(\mem[23][5] ), 
        .ZN(n991) );
  INV_X1 U470 ( .A(n990), .ZN(n698) );
  AOI22_X1 U471 ( .A1(data_in[6]), .A2(n833), .B1(n996), .B2(\mem[23][6] ), 
        .ZN(n990) );
  INV_X1 U472 ( .A(n989), .ZN(n697) );
  AOI22_X1 U473 ( .A1(data_in[7]), .A2(n833), .B1(n996), .B2(\mem[23][7] ), 
        .ZN(n989) );
  INV_X1 U474 ( .A(n988), .ZN(n696) );
  AOI22_X1 U475 ( .A1(data_in[0]), .A2(n832), .B1(n987), .B2(\mem[24][0] ), 
        .ZN(n988) );
  INV_X1 U476 ( .A(n986), .ZN(n695) );
  AOI22_X1 U477 ( .A1(data_in[1]), .A2(n832), .B1(n987), .B2(\mem[24][1] ), 
        .ZN(n986) );
  INV_X1 U478 ( .A(n985), .ZN(n694) );
  AOI22_X1 U479 ( .A1(data_in[2]), .A2(n832), .B1(n987), .B2(\mem[24][2] ), 
        .ZN(n985) );
  INV_X1 U480 ( .A(n984), .ZN(n693) );
  AOI22_X1 U481 ( .A1(data_in[3]), .A2(n832), .B1(n987), .B2(\mem[24][3] ), 
        .ZN(n984) );
  INV_X1 U482 ( .A(n983), .ZN(n692) );
  AOI22_X1 U483 ( .A1(data_in[4]), .A2(n832), .B1(n987), .B2(\mem[24][4] ), 
        .ZN(n983) );
  INV_X1 U484 ( .A(n982), .ZN(n691) );
  AOI22_X1 U485 ( .A1(data_in[5]), .A2(n832), .B1(n987), .B2(\mem[24][5] ), 
        .ZN(n982) );
  INV_X1 U486 ( .A(n981), .ZN(n690) );
  AOI22_X1 U487 ( .A1(data_in[6]), .A2(n832), .B1(n987), .B2(\mem[24][6] ), 
        .ZN(n981) );
  INV_X1 U488 ( .A(n980), .ZN(n689) );
  AOI22_X1 U489 ( .A1(data_in[7]), .A2(n832), .B1(n987), .B2(\mem[24][7] ), 
        .ZN(n980) );
  INV_X1 U490 ( .A(n978), .ZN(n688) );
  AOI22_X1 U491 ( .A1(data_in[0]), .A2(n831), .B1(n977), .B2(\mem[25][0] ), 
        .ZN(n978) );
  INV_X1 U492 ( .A(n976), .ZN(n687) );
  AOI22_X1 U493 ( .A1(data_in[1]), .A2(n831), .B1(n977), .B2(\mem[25][1] ), 
        .ZN(n976) );
  INV_X1 U494 ( .A(n975), .ZN(n686) );
  AOI22_X1 U495 ( .A1(data_in[2]), .A2(n831), .B1(n977), .B2(\mem[25][2] ), 
        .ZN(n975) );
  INV_X1 U496 ( .A(n974), .ZN(n685) );
  AOI22_X1 U497 ( .A1(data_in[3]), .A2(n831), .B1(n977), .B2(\mem[25][3] ), 
        .ZN(n974) );
  INV_X1 U498 ( .A(n973), .ZN(n684) );
  AOI22_X1 U499 ( .A1(data_in[4]), .A2(n831), .B1(n977), .B2(\mem[25][4] ), 
        .ZN(n973) );
  INV_X1 U500 ( .A(n972), .ZN(n683) );
  AOI22_X1 U501 ( .A1(data_in[5]), .A2(n831), .B1(n977), .B2(\mem[25][5] ), 
        .ZN(n972) );
  INV_X1 U502 ( .A(n971), .ZN(n682) );
  AOI22_X1 U503 ( .A1(data_in[6]), .A2(n831), .B1(n977), .B2(\mem[25][6] ), 
        .ZN(n971) );
  INV_X1 U504 ( .A(n970), .ZN(n681) );
  AOI22_X1 U505 ( .A1(data_in[7]), .A2(n831), .B1(n977), .B2(\mem[25][7] ), 
        .ZN(n970) );
  INV_X1 U506 ( .A(n969), .ZN(n680) );
  AOI22_X1 U507 ( .A1(data_in[0]), .A2(n830), .B1(n968), .B2(\mem[26][0] ), 
        .ZN(n969) );
  INV_X1 U508 ( .A(n967), .ZN(n679) );
  AOI22_X1 U509 ( .A1(data_in[1]), .A2(n830), .B1(n968), .B2(\mem[26][1] ), 
        .ZN(n967) );
  INV_X1 U510 ( .A(n966), .ZN(n678) );
  AOI22_X1 U511 ( .A1(data_in[2]), .A2(n830), .B1(n968), .B2(\mem[26][2] ), 
        .ZN(n966) );
  INV_X1 U512 ( .A(n965), .ZN(n677) );
  AOI22_X1 U513 ( .A1(data_in[3]), .A2(n830), .B1(n968), .B2(\mem[26][3] ), 
        .ZN(n965) );
  INV_X1 U514 ( .A(n964), .ZN(n676) );
  AOI22_X1 U515 ( .A1(data_in[4]), .A2(n830), .B1(n968), .B2(\mem[26][4] ), 
        .ZN(n964) );
  INV_X1 U516 ( .A(n963), .ZN(n675) );
  AOI22_X1 U517 ( .A1(data_in[5]), .A2(n830), .B1(n968), .B2(\mem[26][5] ), 
        .ZN(n963) );
  INV_X1 U518 ( .A(n962), .ZN(n674) );
  AOI22_X1 U519 ( .A1(data_in[6]), .A2(n830), .B1(n968), .B2(\mem[26][6] ), 
        .ZN(n962) );
  INV_X1 U520 ( .A(n961), .ZN(n673) );
  AOI22_X1 U521 ( .A1(data_in[7]), .A2(n830), .B1(n968), .B2(\mem[26][7] ), 
        .ZN(n961) );
  INV_X1 U522 ( .A(n960), .ZN(n672) );
  AOI22_X1 U523 ( .A1(data_in[0]), .A2(n829), .B1(n959), .B2(\mem[27][0] ), 
        .ZN(n960) );
  INV_X1 U524 ( .A(n958), .ZN(n671) );
  AOI22_X1 U525 ( .A1(data_in[1]), .A2(n829), .B1(n959), .B2(\mem[27][1] ), 
        .ZN(n958) );
  INV_X1 U526 ( .A(n957), .ZN(n670) );
  AOI22_X1 U527 ( .A1(data_in[2]), .A2(n829), .B1(n959), .B2(\mem[27][2] ), 
        .ZN(n957) );
  INV_X1 U528 ( .A(n956), .ZN(n669) );
  AOI22_X1 U529 ( .A1(data_in[3]), .A2(n829), .B1(n959), .B2(\mem[27][3] ), 
        .ZN(n956) );
  INV_X1 U530 ( .A(n955), .ZN(n668) );
  AOI22_X1 U531 ( .A1(data_in[4]), .A2(n829), .B1(n959), .B2(\mem[27][4] ), 
        .ZN(n955) );
  INV_X1 U532 ( .A(n954), .ZN(n667) );
  AOI22_X1 U533 ( .A1(data_in[5]), .A2(n829), .B1(n959), .B2(\mem[27][5] ), 
        .ZN(n954) );
  INV_X1 U534 ( .A(n953), .ZN(n666) );
  AOI22_X1 U535 ( .A1(data_in[6]), .A2(n829), .B1(n959), .B2(\mem[27][6] ), 
        .ZN(n953) );
  INV_X1 U536 ( .A(n952), .ZN(n665) );
  AOI22_X1 U537 ( .A1(data_in[7]), .A2(n829), .B1(n959), .B2(\mem[27][7] ), 
        .ZN(n952) );
  INV_X1 U538 ( .A(n951), .ZN(n664) );
  AOI22_X1 U539 ( .A1(data_in[0]), .A2(n828), .B1(n950), .B2(\mem[28][0] ), 
        .ZN(n951) );
  INV_X1 U540 ( .A(n949), .ZN(n663) );
  AOI22_X1 U541 ( .A1(data_in[1]), .A2(n828), .B1(n950), .B2(\mem[28][1] ), 
        .ZN(n949) );
  INV_X1 U542 ( .A(n948), .ZN(n662) );
  AOI22_X1 U543 ( .A1(data_in[2]), .A2(n828), .B1(n950), .B2(\mem[28][2] ), 
        .ZN(n948) );
  INV_X1 U544 ( .A(n947), .ZN(n661) );
  AOI22_X1 U545 ( .A1(data_in[3]), .A2(n828), .B1(n950), .B2(\mem[28][3] ), 
        .ZN(n947) );
  INV_X1 U546 ( .A(n946), .ZN(n660) );
  AOI22_X1 U547 ( .A1(data_in[4]), .A2(n828), .B1(n950), .B2(\mem[28][4] ), 
        .ZN(n946) );
  INV_X1 U548 ( .A(n945), .ZN(n659) );
  AOI22_X1 U549 ( .A1(data_in[5]), .A2(n828), .B1(n950), .B2(\mem[28][5] ), 
        .ZN(n945) );
  INV_X1 U550 ( .A(n944), .ZN(n658) );
  AOI22_X1 U551 ( .A1(data_in[6]), .A2(n828), .B1(n950), .B2(\mem[28][6] ), 
        .ZN(n944) );
  INV_X1 U552 ( .A(n943), .ZN(n657) );
  AOI22_X1 U553 ( .A1(data_in[7]), .A2(n828), .B1(n950), .B2(\mem[28][7] ), 
        .ZN(n943) );
  INV_X1 U554 ( .A(n942), .ZN(n656) );
  AOI22_X1 U555 ( .A1(data_in[0]), .A2(n827), .B1(n941), .B2(\mem[29][0] ), 
        .ZN(n942) );
  INV_X1 U556 ( .A(n940), .ZN(n655) );
  AOI22_X1 U557 ( .A1(data_in[1]), .A2(n827), .B1(n941), .B2(\mem[29][1] ), 
        .ZN(n940) );
  INV_X1 U558 ( .A(n939), .ZN(n654) );
  AOI22_X1 U559 ( .A1(data_in[2]), .A2(n827), .B1(n941), .B2(\mem[29][2] ), 
        .ZN(n939) );
  INV_X1 U560 ( .A(n938), .ZN(n653) );
  AOI22_X1 U561 ( .A1(data_in[3]), .A2(n827), .B1(n941), .B2(\mem[29][3] ), 
        .ZN(n938) );
  INV_X1 U562 ( .A(n937), .ZN(n652) );
  AOI22_X1 U563 ( .A1(data_in[4]), .A2(n827), .B1(n941), .B2(\mem[29][4] ), 
        .ZN(n937) );
  INV_X1 U564 ( .A(n936), .ZN(n651) );
  AOI22_X1 U565 ( .A1(data_in[5]), .A2(n827), .B1(n941), .B2(\mem[29][5] ), 
        .ZN(n936) );
  INV_X1 U566 ( .A(n935), .ZN(n650) );
  AOI22_X1 U567 ( .A1(data_in[6]), .A2(n827), .B1(n941), .B2(\mem[29][6] ), 
        .ZN(n935) );
  INV_X1 U568 ( .A(n934), .ZN(n649) );
  AOI22_X1 U569 ( .A1(data_in[7]), .A2(n827), .B1(n941), .B2(\mem[29][7] ), 
        .ZN(n934) );
  INV_X1 U570 ( .A(n933), .ZN(n648) );
  AOI22_X1 U571 ( .A1(data_in[0]), .A2(n826), .B1(n932), .B2(\mem[30][0] ), 
        .ZN(n933) );
  INV_X1 U572 ( .A(n931), .ZN(n647) );
  AOI22_X1 U573 ( .A1(data_in[1]), .A2(n826), .B1(n932), .B2(\mem[30][1] ), 
        .ZN(n931) );
  INV_X1 U574 ( .A(n930), .ZN(n646) );
  AOI22_X1 U575 ( .A1(data_in[2]), .A2(n826), .B1(n932), .B2(\mem[30][2] ), 
        .ZN(n930) );
  INV_X1 U576 ( .A(n929), .ZN(n645) );
  AOI22_X1 U577 ( .A1(data_in[3]), .A2(n826), .B1(n932), .B2(\mem[30][3] ), 
        .ZN(n929) );
  INV_X1 U578 ( .A(n928), .ZN(n644) );
  AOI22_X1 U579 ( .A1(data_in[4]), .A2(n826), .B1(n932), .B2(\mem[30][4] ), 
        .ZN(n928) );
  INV_X1 U580 ( .A(n927), .ZN(n643) );
  AOI22_X1 U581 ( .A1(data_in[5]), .A2(n826), .B1(n932), .B2(\mem[30][5] ), 
        .ZN(n927) );
  INV_X1 U582 ( .A(n926), .ZN(n642) );
  AOI22_X1 U583 ( .A1(data_in[6]), .A2(n826), .B1(n932), .B2(\mem[30][6] ), 
        .ZN(n926) );
  INV_X1 U584 ( .A(n925), .ZN(n641) );
  AOI22_X1 U585 ( .A1(data_in[7]), .A2(n826), .B1(n932), .B2(\mem[30][7] ), 
        .ZN(n925) );
  INV_X1 U586 ( .A(n924), .ZN(n640) );
  AOI22_X1 U587 ( .A1(data_in[0]), .A2(n825), .B1(n923), .B2(\mem[31][0] ), 
        .ZN(n924) );
  INV_X1 U588 ( .A(n922), .ZN(n639) );
  AOI22_X1 U589 ( .A1(data_in[1]), .A2(n825), .B1(n923), .B2(\mem[31][1] ), 
        .ZN(n922) );
  INV_X1 U590 ( .A(n921), .ZN(n638) );
  AOI22_X1 U591 ( .A1(data_in[2]), .A2(n825), .B1(n923), .B2(\mem[31][2] ), 
        .ZN(n921) );
  INV_X1 U592 ( .A(n920), .ZN(n637) );
  AOI22_X1 U593 ( .A1(data_in[3]), .A2(n825), .B1(n923), .B2(\mem[31][3] ), 
        .ZN(n920) );
  INV_X1 U594 ( .A(n919), .ZN(n636) );
  AOI22_X1 U595 ( .A1(data_in[4]), .A2(n825), .B1(n923), .B2(\mem[31][4] ), 
        .ZN(n919) );
  INV_X1 U596 ( .A(n918), .ZN(n635) );
  AOI22_X1 U597 ( .A1(data_in[5]), .A2(n825), .B1(n923), .B2(\mem[31][5] ), 
        .ZN(n918) );
  INV_X1 U598 ( .A(n917), .ZN(n634) );
  AOI22_X1 U599 ( .A1(data_in[6]), .A2(n825), .B1(n923), .B2(\mem[31][6] ), 
        .ZN(n917) );
  INV_X1 U600 ( .A(n916), .ZN(n633) );
  AOI22_X1 U601 ( .A1(data_in[7]), .A2(n825), .B1(n923), .B2(\mem[31][7] ), 
        .ZN(n916) );
  MUX2_X1 U602 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n613), .Z(n3) );
  MUX2_X1 U603 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n613), .Z(n4) );
  MUX2_X1 U604 ( .A(n4), .B(n3), .S(n610), .Z(n5) );
  MUX2_X1 U605 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n613), .Z(n6) );
  MUX2_X1 U606 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n613), .Z(n7) );
  MUX2_X1 U607 ( .A(n7), .B(n6), .S(n610), .Z(n8) );
  MUX2_X1 U608 ( .A(n8), .B(n5), .S(n608), .Z(n9) );
  MUX2_X1 U609 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n613), .Z(n10) );
  MUX2_X1 U610 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n613), .Z(n11) );
  MUX2_X1 U611 ( .A(n11), .B(n10), .S(n610), .Z(n12) );
  MUX2_X1 U612 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n613), .Z(n13) );
  MUX2_X1 U613 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n613), .Z(n14) );
  MUX2_X1 U614 ( .A(n14), .B(n13), .S(n610), .Z(n15) );
  MUX2_X1 U615 ( .A(n15), .B(n12), .S(N12), .Z(n16) );
  MUX2_X1 U616 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U617 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n614), .Z(n18) );
  MUX2_X1 U618 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n614), .Z(n19) );
  MUX2_X1 U619 ( .A(n19), .B(n18), .S(n610), .Z(n20) );
  MUX2_X1 U620 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n614), .Z(n21) );
  MUX2_X1 U621 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n614), .Z(n22) );
  MUX2_X1 U622 ( .A(n22), .B(n21), .S(n611), .Z(n23) );
  MUX2_X1 U623 ( .A(n23), .B(n20), .S(N12), .Z(n24) );
  MUX2_X1 U624 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n614), .Z(n25) );
  MUX2_X1 U625 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n614), .Z(n26) );
  MUX2_X1 U626 ( .A(n26), .B(n25), .S(n610), .Z(n27) );
  MUX2_X1 U627 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n614), .Z(n28) );
  MUX2_X1 U628 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n614), .Z(n29) );
  MUX2_X1 U629 ( .A(n29), .B(n28), .S(N11), .Z(n30) );
  MUX2_X1 U630 ( .A(n30), .B(n27), .S(n609), .Z(n31) );
  MUX2_X1 U631 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U632 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U633 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n614), .Z(n33) );
  MUX2_X1 U634 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n614), .Z(n34) );
  MUX2_X1 U635 ( .A(n34), .B(n33), .S(n610), .Z(n35) );
  MUX2_X1 U636 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n614), .Z(n36) );
  MUX2_X1 U637 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n614), .Z(n37) );
  MUX2_X1 U638 ( .A(n37), .B(n36), .S(n610), .Z(n38) );
  MUX2_X1 U639 ( .A(n38), .B(n35), .S(n609), .Z(n39) );
  MUX2_X1 U640 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n615), .Z(n40) );
  MUX2_X1 U641 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n615), .Z(n41) );
  MUX2_X1 U642 ( .A(n41), .B(n40), .S(n610), .Z(n42) );
  MUX2_X1 U643 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n615), .Z(n43) );
  MUX2_X1 U644 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n615), .Z(n44) );
  MUX2_X1 U645 ( .A(n44), .B(n43), .S(n611), .Z(n45) );
  MUX2_X1 U646 ( .A(n45), .B(n42), .S(n608), .Z(n46) );
  MUX2_X1 U647 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U648 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n615), .Z(n48) );
  MUX2_X1 U649 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n615), .Z(n49) );
  MUX2_X1 U650 ( .A(n49), .B(n48), .S(n610), .Z(n50) );
  MUX2_X1 U651 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n615), .Z(n51) );
  MUX2_X1 U652 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n615), .Z(n52) );
  MUX2_X1 U653 ( .A(n52), .B(n51), .S(n612), .Z(n53) );
  MUX2_X1 U654 ( .A(n53), .B(n50), .S(N12), .Z(n54) );
  MUX2_X1 U655 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n615), .Z(n55) );
  MUX2_X1 U656 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n615), .Z(n56) );
  MUX2_X1 U657 ( .A(n56), .B(n55), .S(n610), .Z(n57) );
  MUX2_X1 U658 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n615), .Z(n58) );
  MUX2_X1 U659 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n615), .Z(n59) );
  MUX2_X1 U660 ( .A(n59), .B(n58), .S(n610), .Z(n60) );
  MUX2_X1 U661 ( .A(n60), .B(n57), .S(n608), .Z(n61) );
  MUX2_X1 U662 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U663 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U664 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n616), .Z(n63) );
  MUX2_X1 U665 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n616), .Z(n64) );
  MUX2_X1 U666 ( .A(n64), .B(n63), .S(n611), .Z(n65) );
  MUX2_X1 U667 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n616), .Z(n66) );
  MUX2_X1 U668 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n616), .Z(n67) );
  MUX2_X1 U669 ( .A(n67), .B(n66), .S(n611), .Z(n68) );
  MUX2_X1 U670 ( .A(n68), .B(n65), .S(n608), .Z(n69) );
  MUX2_X1 U671 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n616), .Z(n70) );
  MUX2_X1 U672 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n616), .Z(n71) );
  MUX2_X1 U673 ( .A(n71), .B(n70), .S(n611), .Z(n72) );
  MUX2_X1 U674 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n616), .Z(n73) );
  MUX2_X1 U675 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n616), .Z(n74) );
  MUX2_X1 U676 ( .A(n74), .B(n73), .S(n611), .Z(n75) );
  MUX2_X1 U677 ( .A(n75), .B(n72), .S(n608), .Z(n76) );
  MUX2_X1 U678 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U679 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n616), .Z(n78) );
  MUX2_X1 U680 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n616), .Z(n79) );
  MUX2_X1 U681 ( .A(n79), .B(n78), .S(n611), .Z(n80) );
  MUX2_X1 U682 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n616), .Z(n81) );
  MUX2_X1 U683 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n616), .Z(n82) );
  MUX2_X1 U684 ( .A(n82), .B(n81), .S(n611), .Z(n83) );
  MUX2_X1 U685 ( .A(n83), .B(n80), .S(n608), .Z(n84) );
  MUX2_X1 U686 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n617), .Z(n85) );
  MUX2_X1 U687 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n617), .Z(n86) );
  MUX2_X1 U688 ( .A(n86), .B(n85), .S(n611), .Z(n87) );
  MUX2_X1 U689 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n617), .Z(n88) );
  MUX2_X1 U690 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n617), .Z(n89) );
  MUX2_X1 U691 ( .A(n89), .B(n88), .S(n611), .Z(n90) );
  MUX2_X1 U692 ( .A(n90), .B(n87), .S(n608), .Z(n91) );
  MUX2_X1 U693 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U694 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U695 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n617), .Z(n93) );
  MUX2_X1 U696 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n617), .Z(n94) );
  MUX2_X1 U697 ( .A(n94), .B(n93), .S(n611), .Z(n95) );
  MUX2_X1 U698 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n617), .Z(n96) );
  MUX2_X1 U699 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n617), .Z(n97) );
  MUX2_X1 U700 ( .A(n97), .B(n96), .S(n611), .Z(n98) );
  MUX2_X1 U701 ( .A(n98), .B(n95), .S(n608), .Z(n99) );
  MUX2_X1 U702 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n617), .Z(n100) );
  MUX2_X1 U703 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n617), .Z(n101) );
  MUX2_X1 U704 ( .A(n101), .B(n100), .S(n611), .Z(n102) );
  MUX2_X1 U705 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n617), .Z(n103) );
  MUX2_X1 U706 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n617), .Z(n104) );
  MUX2_X1 U707 ( .A(n104), .B(n103), .S(n611), .Z(n105) );
  MUX2_X1 U708 ( .A(n105), .B(n102), .S(n608), .Z(n106) );
  MUX2_X1 U709 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U710 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n616), .Z(n108) );
  MUX2_X1 U711 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n621), .Z(n109) );
  MUX2_X1 U712 ( .A(n109), .B(n108), .S(n612), .Z(n110) );
  MUX2_X1 U713 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n622), .Z(n111) );
  MUX2_X1 U714 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n622), .Z(n112) );
  MUX2_X1 U715 ( .A(n112), .B(n111), .S(n612), .Z(n113) );
  MUX2_X1 U716 ( .A(n113), .B(n110), .S(n608), .Z(n114) );
  MUX2_X1 U717 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n621), .Z(n115) );
  MUX2_X1 U718 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n621), .Z(n116) );
  MUX2_X1 U719 ( .A(n116), .B(n115), .S(n612), .Z(n117) );
  MUX2_X1 U720 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n621), .Z(n118) );
  MUX2_X1 U721 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n622), .Z(n119) );
  MUX2_X1 U722 ( .A(n119), .B(n118), .S(n612), .Z(n120) );
  MUX2_X1 U723 ( .A(n120), .B(n117), .S(n608), .Z(n121) );
  MUX2_X1 U724 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U725 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U726 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n622), .Z(n123) );
  MUX2_X1 U727 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n621), .Z(n124) );
  MUX2_X1 U728 ( .A(n124), .B(n123), .S(n612), .Z(n125) );
  MUX2_X1 U729 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n617), .Z(n126) );
  MUX2_X1 U730 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n622), .Z(n127) );
  MUX2_X1 U731 ( .A(n127), .B(n126), .S(n612), .Z(n128) );
  MUX2_X1 U732 ( .A(n128), .B(n125), .S(n608), .Z(n129) );
  MUX2_X1 U733 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n621), .Z(n130) );
  MUX2_X1 U734 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n621), .Z(n131) );
  MUX2_X1 U735 ( .A(n131), .B(n130), .S(n612), .Z(n132) );
  MUX2_X1 U736 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n621), .Z(n133) );
  MUX2_X1 U737 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n622), .Z(n134) );
  MUX2_X1 U738 ( .A(n134), .B(n133), .S(n612), .Z(n135) );
  MUX2_X1 U739 ( .A(n135), .B(n132), .S(n608), .Z(n136) );
  MUX2_X1 U740 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U741 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n613), .Z(n138) );
  MUX2_X1 U742 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n622), .Z(n139) );
  MUX2_X1 U743 ( .A(n139), .B(n138), .S(n612), .Z(n140) );
  MUX2_X1 U744 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n621), .Z(n141) );
  MUX2_X1 U745 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n622), .Z(n142) );
  MUX2_X1 U746 ( .A(n142), .B(n141), .S(n612), .Z(n143) );
  MUX2_X1 U747 ( .A(n143), .B(n140), .S(n608), .Z(n144) );
  MUX2_X1 U748 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n621), .Z(n145) );
  MUX2_X1 U749 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n621), .Z(n146) );
  MUX2_X1 U750 ( .A(n146), .B(n145), .S(n612), .Z(n147) );
  MUX2_X1 U751 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n622), .Z(n148) );
  MUX2_X1 U752 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n622), .Z(n149) );
  MUX2_X1 U753 ( .A(n149), .B(n148), .S(n612), .Z(n150) );
  MUX2_X1 U754 ( .A(n150), .B(n147), .S(n608), .Z(n151) );
  MUX2_X1 U755 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U756 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U757 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n613), .Z(n153) );
  MUX2_X1 U758 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n613), .Z(n154) );
  MUX2_X1 U759 ( .A(n154), .B(n153), .S(n610), .Z(n155) );
  MUX2_X1 U760 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n621), .Z(n156) );
  MUX2_X1 U761 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(N10), .Z(n157) );
  MUX2_X1 U762 ( .A(n157), .B(n156), .S(n612), .Z(n158) );
  MUX2_X1 U763 ( .A(n158), .B(n155), .S(n609), .Z(n159) );
  MUX2_X1 U764 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n622), .Z(n160) );
  MUX2_X1 U765 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(N10), .Z(n161) );
  MUX2_X1 U766 ( .A(n161), .B(n160), .S(N11), .Z(n162) );
  MUX2_X1 U767 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n622), .Z(n163) );
  MUX2_X1 U768 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(N10), .Z(n164) );
  MUX2_X1 U769 ( .A(n164), .B(n163), .S(n612), .Z(n165) );
  MUX2_X1 U770 ( .A(n165), .B(n162), .S(n609), .Z(n166) );
  MUX2_X1 U771 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U772 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n613), .Z(n168) );
  MUX2_X1 U773 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(N10), .Z(n169) );
  MUX2_X1 U774 ( .A(n169), .B(n168), .S(n612), .Z(n170) );
  MUX2_X1 U775 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n621), .Z(n171) );
  MUX2_X1 U776 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(N10), .Z(n172) );
  MUX2_X1 U777 ( .A(n172), .B(n171), .S(n612), .Z(n173) );
  MUX2_X1 U778 ( .A(n173), .B(n170), .S(n609), .Z(n174) );
  MUX2_X1 U779 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n618), .Z(n175) );
  MUX2_X1 U780 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n618), .Z(n176) );
  MUX2_X1 U781 ( .A(n176), .B(n175), .S(n611), .Z(n177) );
  MUX2_X1 U782 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n618), .Z(n178) );
  MUX2_X1 U783 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n618), .Z(n179) );
  MUX2_X1 U784 ( .A(n179), .B(n178), .S(n611), .Z(n180) );
  MUX2_X1 U785 ( .A(n180), .B(n177), .S(n609), .Z(n181) );
  MUX2_X1 U786 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U787 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U788 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n618), .Z(n183) );
  MUX2_X1 U789 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n618), .Z(n184) );
  MUX2_X1 U790 ( .A(n184), .B(n183), .S(n611), .Z(n185) );
  MUX2_X1 U791 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n618), .Z(n186) );
  MUX2_X1 U792 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n618), .Z(n187) );
  MUX2_X1 U793 ( .A(n187), .B(n186), .S(n610), .Z(n188) );
  MUX2_X1 U794 ( .A(n188), .B(n185), .S(n609), .Z(n189) );
  MUX2_X1 U795 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n618), .Z(n190) );
  MUX2_X1 U796 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n618), .Z(n191) );
  MUX2_X1 U797 ( .A(n191), .B(n190), .S(n611), .Z(n192) );
  MUX2_X1 U798 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n618), .Z(n193) );
  MUX2_X1 U799 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n618), .Z(n194) );
  MUX2_X1 U800 ( .A(n194), .B(n193), .S(n610), .Z(n195) );
  MUX2_X1 U801 ( .A(n195), .B(n192), .S(n609), .Z(n196) );
  MUX2_X1 U802 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U803 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n619), .Z(n198) );
  MUX2_X1 U804 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n619), .Z(n199) );
  MUX2_X1 U805 ( .A(n199), .B(n198), .S(n612), .Z(n200) );
  MUX2_X1 U806 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n619), .Z(n201) );
  MUX2_X1 U807 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n619), .Z(n202) );
  MUX2_X1 U808 ( .A(n202), .B(n201), .S(n612), .Z(n203) );
  MUX2_X1 U809 ( .A(n203), .B(n200), .S(n609), .Z(n204) );
  MUX2_X1 U810 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n619), .Z(n205) );
  MUX2_X1 U811 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n619), .Z(n206) );
  MUX2_X1 U812 ( .A(n206), .B(n205), .S(N11), .Z(n207) );
  MUX2_X1 U813 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n619), .Z(n208) );
  MUX2_X1 U814 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n619), .Z(n209) );
  MUX2_X1 U815 ( .A(n209), .B(n208), .S(n611), .Z(n210) );
  MUX2_X1 U816 ( .A(n210), .B(n207), .S(n609), .Z(n211) );
  MUX2_X1 U817 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U818 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U819 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n619), .Z(n213) );
  MUX2_X1 U820 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n619), .Z(n214) );
  MUX2_X1 U821 ( .A(n214), .B(n213), .S(n611), .Z(n215) );
  MUX2_X1 U822 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n619), .Z(n216) );
  MUX2_X1 U823 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n619), .Z(n217) );
  MUX2_X1 U824 ( .A(n217), .B(n216), .S(N11), .Z(n218) );
  MUX2_X1 U825 ( .A(n218), .B(n215), .S(n609), .Z(n219) );
  MUX2_X1 U826 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n620), .Z(n220) );
  MUX2_X1 U827 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n620), .Z(n221) );
  MUX2_X1 U828 ( .A(n221), .B(n220), .S(n610), .Z(n222) );
  MUX2_X1 U829 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n620), .Z(n223) );
  MUX2_X1 U830 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n620), .Z(n224) );
  MUX2_X1 U831 ( .A(n224), .B(n223), .S(N11), .Z(n225) );
  MUX2_X1 U832 ( .A(n225), .B(n222), .S(n609), .Z(n226) );
  MUX2_X1 U833 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U834 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n620), .Z(n228) );
  MUX2_X1 U835 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n620), .Z(n229) );
  MUX2_X1 U836 ( .A(n229), .B(n228), .S(n610), .Z(n595) );
  MUX2_X1 U837 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n620), .Z(n596) );
  MUX2_X1 U838 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n620), .Z(n597) );
  MUX2_X1 U839 ( .A(n597), .B(n596), .S(n610), .Z(n598) );
  MUX2_X1 U840 ( .A(n598), .B(n595), .S(n609), .Z(n599) );
  MUX2_X1 U841 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n620), .Z(n600) );
  MUX2_X1 U842 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n620), .Z(n601) );
  MUX2_X1 U843 ( .A(n601), .B(n600), .S(n611), .Z(n602) );
  MUX2_X1 U844 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n620), .Z(n603) );
  MUX2_X1 U845 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n620), .Z(n604) );
  MUX2_X1 U846 ( .A(n604), .B(n603), .S(n612), .Z(n605) );
  MUX2_X1 U847 ( .A(n605), .B(n602), .S(n609), .Z(n606) );
  MUX2_X1 U848 ( .A(n606), .B(n599), .S(N13), .Z(n607) );
  MUX2_X1 U849 ( .A(n607), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U850 ( .A(N11), .Z(n610) );
  INV_X1 U851 ( .A(N10), .ZN(n623) );
  INV_X1 U852 ( .A(N11), .ZN(n624) );
  INV_X1 U853 ( .A(data_in[0]), .ZN(n625) );
  INV_X1 U854 ( .A(data_in[1]), .ZN(n626) );
  INV_X1 U855 ( .A(data_in[2]), .ZN(n627) );
  INV_X1 U856 ( .A(data_in[3]), .ZN(n628) );
  INV_X1 U857 ( .A(data_in[4]), .ZN(n629) );
  INV_X1 U858 ( .A(data_in[5]), .ZN(n630) );
  INV_X1 U859 ( .A(data_in[6]), .ZN(n631) );
  INV_X1 U860 ( .A(data_in[7]), .ZN(n632) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_2 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n630), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n631), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n632), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n633), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n634), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n635), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n636), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n637), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n638), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n639), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n640), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n641), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n642), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n643), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n644), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n645), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n646), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n647), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n648), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n649), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n650), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n651), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n652), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n653), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n654), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n655), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n656), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n657), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n658), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n659), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n660), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n661), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n662), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n663), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n664), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n665), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n666), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n667), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n668), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n669), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n670), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n671), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n672), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n673), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n674), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n675), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n676), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n677), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n678), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n679), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n680), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n681), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n682), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n683), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n684), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n685), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n686), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n687), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n688), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n689), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n690), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n691), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n692), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n693), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n694), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n695), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n696), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n697), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n698), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n699), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n700), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n701), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n702), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n703), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n704), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n705), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n706), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n707), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n708), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n709), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n710), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n711), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n712), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n713), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n714), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n715), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n716), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n717), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n718), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n719), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n720), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n721), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n722), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n723), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n724), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n725), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n726), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n727), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n728), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n729), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n730), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n731), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n732), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n733), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n734), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n735), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n736), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n737), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n738), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n739), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n740), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n741), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n742), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n743), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n744), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n745), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n746), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n747), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n748), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n749), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n750), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n751), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n752), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n753), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n754), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n755), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n756), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n757), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n758), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n759), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n760), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n761), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n762), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n763), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n764), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n765), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n766), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n767), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n768), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n769), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n770), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n771), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n772), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n773), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n774), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n775), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n776), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n777), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n778), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n779), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n780), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n781), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n782), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n783), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n784), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n785), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n786), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n787), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n788), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n789), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n790), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n791), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n792), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n793), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n794), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n795), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n796), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n797), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n798), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n799), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n800), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n801), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n802), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n803), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n804), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n805), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n806), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n807), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n808), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n809), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n810), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n811), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n812), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n813), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n814), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n815), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n816), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n817), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n818), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n819), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n820), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n821), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n849), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n850), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n851), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n852), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n853), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n854), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n855), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n856), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n857), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n858), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n859), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n860), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n861), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n862), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n863), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n864), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n865), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n866), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n867), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n868), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n869), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n870), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n871), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n872), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n873), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n874), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n875), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n876), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n877), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n878), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n879), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n880), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n881), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n882), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n883), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n884), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n885), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n886), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n887), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n888), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n889), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n890), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n891), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n892), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n893), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n894), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n895), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n896), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n897), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n898), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n899), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n900), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n901), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n902), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n903), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n904), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n905), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n906), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n907), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n908), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n909), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n910), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n911), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n912), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n618), .Z(n611) );
  BUF_X1 U4 ( .A(N11), .Z(n610) );
  BUF_X1 U5 ( .A(N11), .Z(n608) );
  CLKBUF_X1 U6 ( .A(N11), .Z(n609) );
  NOR2_X1 U7 ( .A1(n846), .A2(addr[5]), .ZN(n1132) );
  AND3_X1 U8 ( .A1(n847), .A2(n848), .A3(n1132), .ZN(n1203) );
  AND3_X1 U9 ( .A1(n1132), .A2(n848), .A3(N13), .ZN(n1122) );
  AND3_X1 U10 ( .A1(n1132), .A2(n847), .A3(N14), .ZN(n1049) );
  AND3_X1 U11 ( .A1(N13), .A2(n1132), .A3(N14), .ZN(n976) );
  BUF_X1 U12 ( .A(n619), .Z(n617) );
  BUF_X1 U13 ( .A(n619), .Z(n616) );
  BUF_X1 U14 ( .A(n618), .Z(n612) );
  BUF_X1 U15 ( .A(n618), .Z(n613) );
  BUF_X1 U16 ( .A(n618), .Z(n614) );
  BUF_X1 U17 ( .A(n618), .Z(n615) );
  BUF_X1 U18 ( .A(N10), .Z(n619) );
  BUF_X1 U19 ( .A(N10), .Z(n618) );
  NOR3_X1 U20 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1204) );
  NOR3_X1 U21 ( .A1(N11), .A2(N12), .A3(n620), .ZN(n1193) );
  NOR3_X1 U22 ( .A1(N10), .A2(N12), .A3(n621), .ZN(n1183) );
  NOR3_X1 U23 ( .A1(n620), .A2(N12), .A3(n621), .ZN(n1173) );
  INV_X1 U24 ( .A(n1130), .ZN(n845) );
  INV_X1 U25 ( .A(n1120), .ZN(n844) );
  INV_X1 U26 ( .A(n1111), .ZN(n843) );
  INV_X1 U27 ( .A(n1102), .ZN(n842) );
  INV_X1 U28 ( .A(n1057), .ZN(n837) );
  INV_X1 U29 ( .A(n1047), .ZN(n836) );
  INV_X1 U30 ( .A(n1038), .ZN(n835) );
  INV_X1 U31 ( .A(n1029), .ZN(n834) );
  INV_X1 U32 ( .A(n984), .ZN(n829) );
  INV_X1 U33 ( .A(n974), .ZN(n828) );
  INV_X1 U34 ( .A(n965), .ZN(n827) );
  INV_X1 U35 ( .A(n956), .ZN(n826) );
  INV_X1 U36 ( .A(n1093), .ZN(n841) );
  INV_X1 U37 ( .A(n1084), .ZN(n840) );
  INV_X1 U38 ( .A(n1075), .ZN(n839) );
  INV_X1 U39 ( .A(n1066), .ZN(n838) );
  INV_X1 U40 ( .A(n947), .ZN(n825) );
  INV_X1 U41 ( .A(n938), .ZN(n824) );
  INV_X1 U42 ( .A(n929), .ZN(n823) );
  INV_X1 U43 ( .A(n920), .ZN(n822) );
  INV_X1 U44 ( .A(n1020), .ZN(n833) );
  INV_X1 U45 ( .A(n1011), .ZN(n832) );
  INV_X1 U46 ( .A(n1002), .ZN(n831) );
  INV_X1 U47 ( .A(n993), .ZN(n830) );
  BUF_X1 U48 ( .A(N12), .Z(n607) );
  INV_X1 U49 ( .A(N13), .ZN(n847) );
  AND3_X1 U50 ( .A1(n620), .A2(n621), .A3(N12), .ZN(n1163) );
  AND3_X1 U51 ( .A1(N10), .A2(n621), .A3(N12), .ZN(n1153) );
  AND3_X1 U52 ( .A1(N11), .A2(n620), .A3(N12), .ZN(n1143) );
  AND3_X1 U53 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1133) );
  BUF_X1 U54 ( .A(N12), .Z(n606) );
  INV_X1 U55 ( .A(N14), .ZN(n848) );
  NAND2_X1 U56 ( .A1(n1193), .A2(n1203), .ZN(n1202) );
  NAND2_X1 U57 ( .A1(n1183), .A2(n1203), .ZN(n1192) );
  NAND2_X1 U58 ( .A1(n1173), .A2(n1203), .ZN(n1182) );
  NAND2_X1 U59 ( .A1(n1163), .A2(n1203), .ZN(n1172) );
  NAND2_X1 U60 ( .A1(n1153), .A2(n1203), .ZN(n1162) );
  NAND2_X1 U61 ( .A1(n1143), .A2(n1203), .ZN(n1152) );
  NAND2_X1 U62 ( .A1(n1133), .A2(n1203), .ZN(n1142) );
  NAND2_X1 U63 ( .A1(n1204), .A2(n1203), .ZN(n1213) );
  NAND2_X1 U64 ( .A1(n1122), .A2(n1204), .ZN(n1130) );
  NAND2_X1 U65 ( .A1(n1122), .A2(n1193), .ZN(n1120) );
  NAND2_X1 U66 ( .A1(n1122), .A2(n1183), .ZN(n1111) );
  NAND2_X1 U67 ( .A1(n1122), .A2(n1173), .ZN(n1102) );
  NAND2_X1 U68 ( .A1(n1049), .A2(n1204), .ZN(n1057) );
  NAND2_X1 U69 ( .A1(n1049), .A2(n1193), .ZN(n1047) );
  NAND2_X1 U70 ( .A1(n1049), .A2(n1183), .ZN(n1038) );
  NAND2_X1 U71 ( .A1(n1049), .A2(n1173), .ZN(n1029) );
  NAND2_X1 U72 ( .A1(n976), .A2(n1204), .ZN(n984) );
  NAND2_X1 U73 ( .A1(n976), .A2(n1193), .ZN(n974) );
  NAND2_X1 U74 ( .A1(n976), .A2(n1183), .ZN(n965) );
  NAND2_X1 U75 ( .A1(n976), .A2(n1173), .ZN(n956) );
  NAND2_X1 U76 ( .A1(n1122), .A2(n1163), .ZN(n1093) );
  NAND2_X1 U77 ( .A1(n1122), .A2(n1153), .ZN(n1084) );
  NAND2_X1 U78 ( .A1(n1122), .A2(n1143), .ZN(n1075) );
  NAND2_X1 U79 ( .A1(n1122), .A2(n1133), .ZN(n1066) );
  NAND2_X1 U80 ( .A1(n1049), .A2(n1163), .ZN(n1020) );
  NAND2_X1 U81 ( .A1(n1049), .A2(n1153), .ZN(n1011) );
  NAND2_X1 U82 ( .A1(n1049), .A2(n1143), .ZN(n1002) );
  NAND2_X1 U83 ( .A1(n1049), .A2(n1133), .ZN(n993) );
  NAND2_X1 U84 ( .A1(n976), .A2(n1163), .ZN(n947) );
  NAND2_X1 U85 ( .A1(n976), .A2(n1153), .ZN(n938) );
  NAND2_X1 U86 ( .A1(n976), .A2(n1143), .ZN(n929) );
  NAND2_X1 U87 ( .A1(n976), .A2(n1133), .ZN(n920) );
  INV_X1 U88 ( .A(wr_en), .ZN(n846) );
  OAI21_X1 U89 ( .B1(n622), .B2(n1172), .A(n1171), .ZN(n880) );
  NAND2_X1 U90 ( .A1(\mem[4][0] ), .A2(n1172), .ZN(n1171) );
  OAI21_X1 U91 ( .B1(n623), .B2(n1172), .A(n1170), .ZN(n879) );
  NAND2_X1 U92 ( .A1(\mem[4][1] ), .A2(n1172), .ZN(n1170) );
  OAI21_X1 U93 ( .B1(n624), .B2(n1172), .A(n1169), .ZN(n878) );
  NAND2_X1 U94 ( .A1(\mem[4][2] ), .A2(n1172), .ZN(n1169) );
  OAI21_X1 U95 ( .B1(n625), .B2(n1172), .A(n1168), .ZN(n877) );
  NAND2_X1 U96 ( .A1(\mem[4][3] ), .A2(n1172), .ZN(n1168) );
  OAI21_X1 U97 ( .B1(n626), .B2(n1172), .A(n1167), .ZN(n876) );
  NAND2_X1 U98 ( .A1(\mem[4][4] ), .A2(n1172), .ZN(n1167) );
  OAI21_X1 U99 ( .B1(n627), .B2(n1172), .A(n1166), .ZN(n875) );
  NAND2_X1 U100 ( .A1(\mem[4][5] ), .A2(n1172), .ZN(n1166) );
  OAI21_X1 U101 ( .B1(n628), .B2(n1172), .A(n1165), .ZN(n874) );
  NAND2_X1 U102 ( .A1(\mem[4][6] ), .A2(n1172), .ZN(n1165) );
  OAI21_X1 U103 ( .B1(n629), .B2(n1172), .A(n1164), .ZN(n873) );
  NAND2_X1 U104 ( .A1(\mem[4][7] ), .A2(n1172), .ZN(n1164) );
  OAI21_X1 U105 ( .B1(n622), .B2(n1152), .A(n1151), .ZN(n864) );
  NAND2_X1 U106 ( .A1(\mem[6][0] ), .A2(n1152), .ZN(n1151) );
  OAI21_X1 U107 ( .B1(n623), .B2(n1152), .A(n1150), .ZN(n863) );
  NAND2_X1 U108 ( .A1(\mem[6][1] ), .A2(n1152), .ZN(n1150) );
  OAI21_X1 U109 ( .B1(n624), .B2(n1152), .A(n1149), .ZN(n862) );
  NAND2_X1 U110 ( .A1(\mem[6][2] ), .A2(n1152), .ZN(n1149) );
  OAI21_X1 U111 ( .B1(n625), .B2(n1152), .A(n1148), .ZN(n861) );
  NAND2_X1 U112 ( .A1(\mem[6][3] ), .A2(n1152), .ZN(n1148) );
  OAI21_X1 U113 ( .B1(n626), .B2(n1152), .A(n1147), .ZN(n860) );
  NAND2_X1 U114 ( .A1(\mem[6][4] ), .A2(n1152), .ZN(n1147) );
  OAI21_X1 U115 ( .B1(n627), .B2(n1152), .A(n1146), .ZN(n859) );
  NAND2_X1 U116 ( .A1(\mem[6][5] ), .A2(n1152), .ZN(n1146) );
  OAI21_X1 U117 ( .B1(n628), .B2(n1152), .A(n1145), .ZN(n858) );
  NAND2_X1 U118 ( .A1(\mem[6][6] ), .A2(n1152), .ZN(n1145) );
  OAI21_X1 U119 ( .B1(n629), .B2(n1152), .A(n1144), .ZN(n857) );
  NAND2_X1 U120 ( .A1(\mem[6][7] ), .A2(n1152), .ZN(n1144) );
  OAI21_X1 U121 ( .B1(n622), .B2(n1142), .A(n1141), .ZN(n856) );
  NAND2_X1 U122 ( .A1(\mem[7][0] ), .A2(n1142), .ZN(n1141) );
  OAI21_X1 U123 ( .B1(n623), .B2(n1142), .A(n1140), .ZN(n855) );
  NAND2_X1 U124 ( .A1(\mem[7][1] ), .A2(n1142), .ZN(n1140) );
  OAI21_X1 U125 ( .B1(n624), .B2(n1142), .A(n1139), .ZN(n854) );
  NAND2_X1 U126 ( .A1(\mem[7][2] ), .A2(n1142), .ZN(n1139) );
  OAI21_X1 U127 ( .B1(n625), .B2(n1142), .A(n1138), .ZN(n853) );
  NAND2_X1 U128 ( .A1(\mem[7][3] ), .A2(n1142), .ZN(n1138) );
  OAI21_X1 U129 ( .B1(n626), .B2(n1142), .A(n1137), .ZN(n852) );
  NAND2_X1 U130 ( .A1(\mem[7][4] ), .A2(n1142), .ZN(n1137) );
  OAI21_X1 U131 ( .B1(n627), .B2(n1142), .A(n1136), .ZN(n851) );
  NAND2_X1 U132 ( .A1(\mem[7][5] ), .A2(n1142), .ZN(n1136) );
  OAI21_X1 U133 ( .B1(n628), .B2(n1142), .A(n1135), .ZN(n850) );
  NAND2_X1 U134 ( .A1(\mem[7][6] ), .A2(n1142), .ZN(n1135) );
  OAI21_X1 U135 ( .B1(n629), .B2(n1142), .A(n1134), .ZN(n849) );
  NAND2_X1 U136 ( .A1(\mem[7][7] ), .A2(n1142), .ZN(n1134) );
  OAI21_X1 U137 ( .B1(n622), .B2(n1202), .A(n1201), .ZN(n904) );
  NAND2_X1 U138 ( .A1(\mem[1][0] ), .A2(n1202), .ZN(n1201) );
  OAI21_X1 U139 ( .B1(n623), .B2(n1202), .A(n1200), .ZN(n903) );
  NAND2_X1 U140 ( .A1(\mem[1][1] ), .A2(n1202), .ZN(n1200) );
  OAI21_X1 U141 ( .B1(n624), .B2(n1202), .A(n1199), .ZN(n902) );
  NAND2_X1 U142 ( .A1(\mem[1][2] ), .A2(n1202), .ZN(n1199) );
  OAI21_X1 U143 ( .B1(n625), .B2(n1202), .A(n1198), .ZN(n901) );
  NAND2_X1 U144 ( .A1(\mem[1][3] ), .A2(n1202), .ZN(n1198) );
  OAI21_X1 U145 ( .B1(n626), .B2(n1202), .A(n1197), .ZN(n900) );
  NAND2_X1 U146 ( .A1(\mem[1][4] ), .A2(n1202), .ZN(n1197) );
  OAI21_X1 U147 ( .B1(n627), .B2(n1202), .A(n1196), .ZN(n899) );
  NAND2_X1 U148 ( .A1(\mem[1][5] ), .A2(n1202), .ZN(n1196) );
  OAI21_X1 U149 ( .B1(n628), .B2(n1202), .A(n1195), .ZN(n898) );
  NAND2_X1 U150 ( .A1(\mem[1][6] ), .A2(n1202), .ZN(n1195) );
  OAI21_X1 U151 ( .B1(n629), .B2(n1202), .A(n1194), .ZN(n897) );
  NAND2_X1 U152 ( .A1(\mem[1][7] ), .A2(n1202), .ZN(n1194) );
  OAI21_X1 U153 ( .B1(n622), .B2(n1192), .A(n1191), .ZN(n896) );
  NAND2_X1 U154 ( .A1(\mem[2][0] ), .A2(n1192), .ZN(n1191) );
  OAI21_X1 U155 ( .B1(n623), .B2(n1192), .A(n1190), .ZN(n895) );
  NAND2_X1 U156 ( .A1(\mem[2][1] ), .A2(n1192), .ZN(n1190) );
  OAI21_X1 U157 ( .B1(n624), .B2(n1192), .A(n1189), .ZN(n894) );
  NAND2_X1 U158 ( .A1(\mem[2][2] ), .A2(n1192), .ZN(n1189) );
  OAI21_X1 U159 ( .B1(n625), .B2(n1192), .A(n1188), .ZN(n893) );
  NAND2_X1 U160 ( .A1(\mem[2][3] ), .A2(n1192), .ZN(n1188) );
  OAI21_X1 U161 ( .B1(n626), .B2(n1192), .A(n1187), .ZN(n892) );
  NAND2_X1 U162 ( .A1(\mem[2][4] ), .A2(n1192), .ZN(n1187) );
  OAI21_X1 U163 ( .B1(n627), .B2(n1192), .A(n1186), .ZN(n891) );
  NAND2_X1 U164 ( .A1(\mem[2][5] ), .A2(n1192), .ZN(n1186) );
  OAI21_X1 U165 ( .B1(n628), .B2(n1192), .A(n1185), .ZN(n890) );
  NAND2_X1 U166 ( .A1(\mem[2][6] ), .A2(n1192), .ZN(n1185) );
  OAI21_X1 U167 ( .B1(n629), .B2(n1192), .A(n1184), .ZN(n889) );
  NAND2_X1 U168 ( .A1(\mem[2][7] ), .A2(n1192), .ZN(n1184) );
  OAI21_X1 U169 ( .B1(n622), .B2(n1182), .A(n1181), .ZN(n888) );
  NAND2_X1 U170 ( .A1(\mem[3][0] ), .A2(n1182), .ZN(n1181) );
  OAI21_X1 U171 ( .B1(n623), .B2(n1182), .A(n1180), .ZN(n887) );
  NAND2_X1 U172 ( .A1(\mem[3][1] ), .A2(n1182), .ZN(n1180) );
  OAI21_X1 U173 ( .B1(n624), .B2(n1182), .A(n1179), .ZN(n886) );
  NAND2_X1 U174 ( .A1(\mem[3][2] ), .A2(n1182), .ZN(n1179) );
  OAI21_X1 U175 ( .B1(n625), .B2(n1182), .A(n1178), .ZN(n885) );
  NAND2_X1 U176 ( .A1(\mem[3][3] ), .A2(n1182), .ZN(n1178) );
  OAI21_X1 U177 ( .B1(n626), .B2(n1182), .A(n1177), .ZN(n884) );
  NAND2_X1 U178 ( .A1(\mem[3][4] ), .A2(n1182), .ZN(n1177) );
  OAI21_X1 U179 ( .B1(n627), .B2(n1182), .A(n1176), .ZN(n883) );
  NAND2_X1 U180 ( .A1(\mem[3][5] ), .A2(n1182), .ZN(n1176) );
  OAI21_X1 U181 ( .B1(n628), .B2(n1182), .A(n1175), .ZN(n882) );
  NAND2_X1 U182 ( .A1(\mem[3][6] ), .A2(n1182), .ZN(n1175) );
  OAI21_X1 U183 ( .B1(n629), .B2(n1182), .A(n1174), .ZN(n881) );
  NAND2_X1 U184 ( .A1(\mem[3][7] ), .A2(n1182), .ZN(n1174) );
  OAI21_X1 U185 ( .B1(n622), .B2(n1162), .A(n1161), .ZN(n872) );
  NAND2_X1 U186 ( .A1(\mem[5][0] ), .A2(n1162), .ZN(n1161) );
  OAI21_X1 U187 ( .B1(n623), .B2(n1162), .A(n1160), .ZN(n871) );
  NAND2_X1 U188 ( .A1(\mem[5][1] ), .A2(n1162), .ZN(n1160) );
  OAI21_X1 U189 ( .B1(n624), .B2(n1162), .A(n1159), .ZN(n870) );
  NAND2_X1 U190 ( .A1(\mem[5][2] ), .A2(n1162), .ZN(n1159) );
  OAI21_X1 U191 ( .B1(n625), .B2(n1162), .A(n1158), .ZN(n869) );
  NAND2_X1 U192 ( .A1(\mem[5][3] ), .A2(n1162), .ZN(n1158) );
  OAI21_X1 U193 ( .B1(n626), .B2(n1162), .A(n1157), .ZN(n868) );
  NAND2_X1 U194 ( .A1(\mem[5][4] ), .A2(n1162), .ZN(n1157) );
  OAI21_X1 U195 ( .B1(n627), .B2(n1162), .A(n1156), .ZN(n867) );
  NAND2_X1 U196 ( .A1(\mem[5][5] ), .A2(n1162), .ZN(n1156) );
  OAI21_X1 U197 ( .B1(n628), .B2(n1162), .A(n1155), .ZN(n866) );
  NAND2_X1 U198 ( .A1(\mem[5][6] ), .A2(n1162), .ZN(n1155) );
  OAI21_X1 U199 ( .B1(n629), .B2(n1162), .A(n1154), .ZN(n865) );
  NAND2_X1 U200 ( .A1(\mem[5][7] ), .A2(n1162), .ZN(n1154) );
  OAI21_X1 U201 ( .B1(n1213), .B2(n622), .A(n1212), .ZN(n912) );
  NAND2_X1 U202 ( .A1(\mem[0][0] ), .A2(n1213), .ZN(n1212) );
  OAI21_X1 U203 ( .B1(n1213), .B2(n623), .A(n1211), .ZN(n911) );
  NAND2_X1 U204 ( .A1(\mem[0][1] ), .A2(n1213), .ZN(n1211) );
  OAI21_X1 U205 ( .B1(n1213), .B2(n624), .A(n1210), .ZN(n910) );
  NAND2_X1 U206 ( .A1(\mem[0][2] ), .A2(n1213), .ZN(n1210) );
  OAI21_X1 U207 ( .B1(n1213), .B2(n625), .A(n1209), .ZN(n909) );
  NAND2_X1 U208 ( .A1(\mem[0][3] ), .A2(n1213), .ZN(n1209) );
  OAI21_X1 U209 ( .B1(n1213), .B2(n626), .A(n1208), .ZN(n908) );
  NAND2_X1 U210 ( .A1(\mem[0][4] ), .A2(n1213), .ZN(n1208) );
  OAI21_X1 U211 ( .B1(n1213), .B2(n627), .A(n1207), .ZN(n907) );
  NAND2_X1 U212 ( .A1(\mem[0][5] ), .A2(n1213), .ZN(n1207) );
  OAI21_X1 U213 ( .B1(n1213), .B2(n628), .A(n1206), .ZN(n906) );
  NAND2_X1 U214 ( .A1(\mem[0][6] ), .A2(n1213), .ZN(n1206) );
  OAI21_X1 U215 ( .B1(n1213), .B2(n629), .A(n1205), .ZN(n905) );
  NAND2_X1 U216 ( .A1(\mem[0][7] ), .A2(n1213), .ZN(n1205) );
  INV_X1 U217 ( .A(n1131), .ZN(n821) );
  AOI22_X1 U218 ( .A1(data_in[0]), .A2(n845), .B1(n1130), .B2(\mem[8][0] ), 
        .ZN(n1131) );
  INV_X1 U219 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U220 ( .A1(data_in[1]), .A2(n845), .B1(n1130), .B2(\mem[8][1] ), 
        .ZN(n1129) );
  INV_X1 U221 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U222 ( .A1(data_in[2]), .A2(n845), .B1(n1130), .B2(\mem[8][2] ), 
        .ZN(n1128) );
  INV_X1 U223 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U224 ( .A1(data_in[3]), .A2(n845), .B1(n1130), .B2(\mem[8][3] ), 
        .ZN(n1127) );
  INV_X1 U225 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U226 ( .A1(data_in[4]), .A2(n845), .B1(n1130), .B2(\mem[8][4] ), 
        .ZN(n1126) );
  INV_X1 U227 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U228 ( .A1(data_in[5]), .A2(n845), .B1(n1130), .B2(\mem[8][5] ), 
        .ZN(n1125) );
  INV_X1 U229 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U230 ( .A1(data_in[6]), .A2(n845), .B1(n1130), .B2(\mem[8][6] ), 
        .ZN(n1124) );
  INV_X1 U231 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U232 ( .A1(data_in[7]), .A2(n845), .B1(n1130), .B2(\mem[8][7] ), 
        .ZN(n1123) );
  INV_X1 U233 ( .A(n1121), .ZN(n813) );
  AOI22_X1 U234 ( .A1(data_in[0]), .A2(n844), .B1(n1120), .B2(\mem[9][0] ), 
        .ZN(n1121) );
  INV_X1 U235 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U236 ( .A1(data_in[1]), .A2(n844), .B1(n1120), .B2(\mem[9][1] ), 
        .ZN(n1119) );
  INV_X1 U237 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U238 ( .A1(data_in[2]), .A2(n844), .B1(n1120), .B2(\mem[9][2] ), 
        .ZN(n1118) );
  INV_X1 U239 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U240 ( .A1(data_in[3]), .A2(n844), .B1(n1120), .B2(\mem[9][3] ), 
        .ZN(n1117) );
  INV_X1 U241 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U242 ( .A1(data_in[4]), .A2(n844), .B1(n1120), .B2(\mem[9][4] ), 
        .ZN(n1116) );
  INV_X1 U243 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U244 ( .A1(data_in[5]), .A2(n844), .B1(n1120), .B2(\mem[9][5] ), 
        .ZN(n1115) );
  INV_X1 U245 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U246 ( .A1(data_in[6]), .A2(n844), .B1(n1120), .B2(\mem[9][6] ), 
        .ZN(n1114) );
  INV_X1 U247 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U248 ( .A1(data_in[7]), .A2(n844), .B1(n1120), .B2(\mem[9][7] ), 
        .ZN(n1113) );
  INV_X1 U249 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U250 ( .A1(data_in[0]), .A2(n843), .B1(n1111), .B2(\mem[10][0] ), 
        .ZN(n1112) );
  INV_X1 U251 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U252 ( .A1(data_in[1]), .A2(n843), .B1(n1111), .B2(\mem[10][1] ), 
        .ZN(n1110) );
  INV_X1 U253 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U254 ( .A1(data_in[2]), .A2(n843), .B1(n1111), .B2(\mem[10][2] ), 
        .ZN(n1109) );
  INV_X1 U255 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U256 ( .A1(data_in[3]), .A2(n843), .B1(n1111), .B2(\mem[10][3] ), 
        .ZN(n1108) );
  INV_X1 U257 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U258 ( .A1(data_in[4]), .A2(n843), .B1(n1111), .B2(\mem[10][4] ), 
        .ZN(n1107) );
  INV_X1 U259 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U260 ( .A1(data_in[5]), .A2(n843), .B1(n1111), .B2(\mem[10][5] ), 
        .ZN(n1106) );
  INV_X1 U261 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U262 ( .A1(data_in[6]), .A2(n843), .B1(n1111), .B2(\mem[10][6] ), 
        .ZN(n1105) );
  INV_X1 U263 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U264 ( .A1(data_in[7]), .A2(n843), .B1(n1111), .B2(\mem[10][7] ), 
        .ZN(n1104) );
  INV_X1 U265 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U266 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[11][0] ), 
        .ZN(n1103) );
  INV_X1 U267 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U268 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[11][1] ), 
        .ZN(n1101) );
  INV_X1 U269 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U270 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[11][2] ), 
        .ZN(n1100) );
  INV_X1 U271 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U272 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[11][3] ), 
        .ZN(n1099) );
  INV_X1 U273 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U274 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[11][4] ), 
        .ZN(n1098) );
  INV_X1 U275 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U276 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[11][5] ), 
        .ZN(n1097) );
  INV_X1 U277 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U278 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[11][6] ), 
        .ZN(n1096) );
  INV_X1 U279 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U280 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[11][7] ), 
        .ZN(n1095) );
  INV_X1 U281 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U282 ( .A1(data_in[0]), .A2(n841), .B1(n1093), .B2(\mem[12][0] ), 
        .ZN(n1094) );
  INV_X1 U283 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U284 ( .A1(data_in[1]), .A2(n841), .B1(n1093), .B2(\mem[12][1] ), 
        .ZN(n1092) );
  INV_X1 U285 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U286 ( .A1(data_in[2]), .A2(n841), .B1(n1093), .B2(\mem[12][2] ), 
        .ZN(n1091) );
  INV_X1 U287 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U288 ( .A1(data_in[3]), .A2(n841), .B1(n1093), .B2(\mem[12][3] ), 
        .ZN(n1090) );
  INV_X1 U289 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U290 ( .A1(data_in[4]), .A2(n841), .B1(n1093), .B2(\mem[12][4] ), 
        .ZN(n1089) );
  INV_X1 U291 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U292 ( .A1(data_in[5]), .A2(n841), .B1(n1093), .B2(\mem[12][5] ), 
        .ZN(n1088) );
  INV_X1 U293 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U294 ( .A1(data_in[6]), .A2(n841), .B1(n1093), .B2(\mem[12][6] ), 
        .ZN(n1087) );
  INV_X1 U295 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U296 ( .A1(data_in[7]), .A2(n841), .B1(n1093), .B2(\mem[12][7] ), 
        .ZN(n1086) );
  INV_X1 U297 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U298 ( .A1(data_in[0]), .A2(n840), .B1(n1084), .B2(\mem[13][0] ), 
        .ZN(n1085) );
  INV_X1 U299 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U300 ( .A1(data_in[1]), .A2(n840), .B1(n1084), .B2(\mem[13][1] ), 
        .ZN(n1083) );
  INV_X1 U301 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U302 ( .A1(data_in[2]), .A2(n840), .B1(n1084), .B2(\mem[13][2] ), 
        .ZN(n1082) );
  INV_X1 U303 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U304 ( .A1(data_in[3]), .A2(n840), .B1(n1084), .B2(\mem[13][3] ), 
        .ZN(n1081) );
  INV_X1 U305 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U306 ( .A1(data_in[4]), .A2(n840), .B1(n1084), .B2(\mem[13][4] ), 
        .ZN(n1080) );
  INV_X1 U307 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U308 ( .A1(data_in[5]), .A2(n840), .B1(n1084), .B2(\mem[13][5] ), 
        .ZN(n1079) );
  INV_X1 U309 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U310 ( .A1(data_in[6]), .A2(n840), .B1(n1084), .B2(\mem[13][6] ), 
        .ZN(n1078) );
  INV_X1 U311 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U312 ( .A1(data_in[7]), .A2(n840), .B1(n1084), .B2(\mem[13][7] ), 
        .ZN(n1077) );
  INV_X1 U313 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U314 ( .A1(data_in[0]), .A2(n839), .B1(n1075), .B2(\mem[14][0] ), 
        .ZN(n1076) );
  INV_X1 U315 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U316 ( .A1(data_in[1]), .A2(n839), .B1(n1075), .B2(\mem[14][1] ), 
        .ZN(n1074) );
  INV_X1 U317 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U318 ( .A1(data_in[2]), .A2(n839), .B1(n1075), .B2(\mem[14][2] ), 
        .ZN(n1073) );
  INV_X1 U319 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U320 ( .A1(data_in[3]), .A2(n839), .B1(n1075), .B2(\mem[14][3] ), 
        .ZN(n1072) );
  INV_X1 U321 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U322 ( .A1(data_in[4]), .A2(n839), .B1(n1075), .B2(\mem[14][4] ), 
        .ZN(n1071) );
  INV_X1 U323 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U324 ( .A1(data_in[5]), .A2(n839), .B1(n1075), .B2(\mem[14][5] ), 
        .ZN(n1070) );
  INV_X1 U325 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U326 ( .A1(data_in[6]), .A2(n839), .B1(n1075), .B2(\mem[14][6] ), 
        .ZN(n1069) );
  INV_X1 U327 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U328 ( .A1(data_in[7]), .A2(n839), .B1(n1075), .B2(\mem[14][7] ), 
        .ZN(n1068) );
  INV_X1 U329 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U330 ( .A1(data_in[0]), .A2(n838), .B1(n1066), .B2(\mem[15][0] ), 
        .ZN(n1067) );
  INV_X1 U331 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U332 ( .A1(data_in[1]), .A2(n838), .B1(n1066), .B2(\mem[15][1] ), 
        .ZN(n1065) );
  INV_X1 U333 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U334 ( .A1(data_in[2]), .A2(n838), .B1(n1066), .B2(\mem[15][2] ), 
        .ZN(n1064) );
  INV_X1 U335 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U336 ( .A1(data_in[3]), .A2(n838), .B1(n1066), .B2(\mem[15][3] ), 
        .ZN(n1063) );
  INV_X1 U337 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U338 ( .A1(data_in[4]), .A2(n838), .B1(n1066), .B2(\mem[15][4] ), 
        .ZN(n1062) );
  INV_X1 U339 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U340 ( .A1(data_in[5]), .A2(n838), .B1(n1066), .B2(\mem[15][5] ), 
        .ZN(n1061) );
  INV_X1 U341 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U342 ( .A1(data_in[6]), .A2(n838), .B1(n1066), .B2(\mem[15][6] ), 
        .ZN(n1060) );
  INV_X1 U343 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U344 ( .A1(data_in[7]), .A2(n838), .B1(n1066), .B2(\mem[15][7] ), 
        .ZN(n1059) );
  INV_X1 U345 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U346 ( .A1(data_in[0]), .A2(n837), .B1(n1057), .B2(\mem[16][0] ), 
        .ZN(n1058) );
  INV_X1 U347 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U348 ( .A1(data_in[1]), .A2(n837), .B1(n1057), .B2(\mem[16][1] ), 
        .ZN(n1056) );
  INV_X1 U349 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U350 ( .A1(data_in[2]), .A2(n837), .B1(n1057), .B2(\mem[16][2] ), 
        .ZN(n1055) );
  INV_X1 U351 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U352 ( .A1(data_in[3]), .A2(n837), .B1(n1057), .B2(\mem[16][3] ), 
        .ZN(n1054) );
  INV_X1 U353 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U354 ( .A1(data_in[4]), .A2(n837), .B1(n1057), .B2(\mem[16][4] ), 
        .ZN(n1053) );
  INV_X1 U355 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U356 ( .A1(data_in[5]), .A2(n837), .B1(n1057), .B2(\mem[16][5] ), 
        .ZN(n1052) );
  INV_X1 U357 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U358 ( .A1(data_in[6]), .A2(n837), .B1(n1057), .B2(\mem[16][6] ), 
        .ZN(n1051) );
  INV_X1 U359 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U360 ( .A1(data_in[7]), .A2(n837), .B1(n1057), .B2(\mem[16][7] ), 
        .ZN(n1050) );
  INV_X1 U361 ( .A(n1048), .ZN(n749) );
  AOI22_X1 U362 ( .A1(data_in[0]), .A2(n836), .B1(n1047), .B2(\mem[17][0] ), 
        .ZN(n1048) );
  INV_X1 U363 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U364 ( .A1(data_in[1]), .A2(n836), .B1(n1047), .B2(\mem[17][1] ), 
        .ZN(n1046) );
  INV_X1 U365 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U366 ( .A1(data_in[2]), .A2(n836), .B1(n1047), .B2(\mem[17][2] ), 
        .ZN(n1045) );
  INV_X1 U367 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U368 ( .A1(data_in[3]), .A2(n836), .B1(n1047), .B2(\mem[17][3] ), 
        .ZN(n1044) );
  INV_X1 U369 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U370 ( .A1(data_in[4]), .A2(n836), .B1(n1047), .B2(\mem[17][4] ), 
        .ZN(n1043) );
  INV_X1 U371 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U372 ( .A1(data_in[5]), .A2(n836), .B1(n1047), .B2(\mem[17][5] ), 
        .ZN(n1042) );
  INV_X1 U373 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U374 ( .A1(data_in[6]), .A2(n836), .B1(n1047), .B2(\mem[17][6] ), 
        .ZN(n1041) );
  INV_X1 U375 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U376 ( .A1(data_in[7]), .A2(n836), .B1(n1047), .B2(\mem[17][7] ), 
        .ZN(n1040) );
  INV_X1 U377 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U378 ( .A1(data_in[0]), .A2(n835), .B1(n1038), .B2(\mem[18][0] ), 
        .ZN(n1039) );
  INV_X1 U379 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U380 ( .A1(data_in[1]), .A2(n835), .B1(n1038), .B2(\mem[18][1] ), 
        .ZN(n1037) );
  INV_X1 U381 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U382 ( .A1(data_in[2]), .A2(n835), .B1(n1038), .B2(\mem[18][2] ), 
        .ZN(n1036) );
  INV_X1 U383 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U384 ( .A1(data_in[3]), .A2(n835), .B1(n1038), .B2(\mem[18][3] ), 
        .ZN(n1035) );
  INV_X1 U385 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U386 ( .A1(data_in[4]), .A2(n835), .B1(n1038), .B2(\mem[18][4] ), 
        .ZN(n1034) );
  INV_X1 U387 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U388 ( .A1(data_in[5]), .A2(n835), .B1(n1038), .B2(\mem[18][5] ), 
        .ZN(n1033) );
  INV_X1 U389 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U390 ( .A1(data_in[6]), .A2(n835), .B1(n1038), .B2(\mem[18][6] ), 
        .ZN(n1032) );
  INV_X1 U391 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U392 ( .A1(data_in[7]), .A2(n835), .B1(n1038), .B2(\mem[18][7] ), 
        .ZN(n1031) );
  INV_X1 U393 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U394 ( .A1(data_in[0]), .A2(n834), .B1(n1029), .B2(\mem[19][0] ), 
        .ZN(n1030) );
  INV_X1 U395 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U396 ( .A1(data_in[1]), .A2(n834), .B1(n1029), .B2(\mem[19][1] ), 
        .ZN(n1028) );
  INV_X1 U397 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U398 ( .A1(data_in[2]), .A2(n834), .B1(n1029), .B2(\mem[19][2] ), 
        .ZN(n1027) );
  INV_X1 U399 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U400 ( .A1(data_in[3]), .A2(n834), .B1(n1029), .B2(\mem[19][3] ), 
        .ZN(n1026) );
  INV_X1 U401 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U402 ( .A1(data_in[4]), .A2(n834), .B1(n1029), .B2(\mem[19][4] ), 
        .ZN(n1025) );
  INV_X1 U403 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U404 ( .A1(data_in[5]), .A2(n834), .B1(n1029), .B2(\mem[19][5] ), 
        .ZN(n1024) );
  INV_X1 U405 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U406 ( .A1(data_in[6]), .A2(n834), .B1(n1029), .B2(\mem[19][6] ), 
        .ZN(n1023) );
  INV_X1 U407 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U408 ( .A1(data_in[7]), .A2(n834), .B1(n1029), .B2(\mem[19][7] ), 
        .ZN(n1022) );
  INV_X1 U409 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U410 ( .A1(data_in[0]), .A2(n833), .B1(n1020), .B2(\mem[20][0] ), 
        .ZN(n1021) );
  INV_X1 U411 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U412 ( .A1(data_in[1]), .A2(n833), .B1(n1020), .B2(\mem[20][1] ), 
        .ZN(n1019) );
  INV_X1 U413 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U414 ( .A1(data_in[2]), .A2(n833), .B1(n1020), .B2(\mem[20][2] ), 
        .ZN(n1018) );
  INV_X1 U415 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U416 ( .A1(data_in[3]), .A2(n833), .B1(n1020), .B2(\mem[20][3] ), 
        .ZN(n1017) );
  INV_X1 U417 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U418 ( .A1(data_in[4]), .A2(n833), .B1(n1020), .B2(\mem[20][4] ), 
        .ZN(n1016) );
  INV_X1 U419 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U420 ( .A1(data_in[5]), .A2(n833), .B1(n1020), .B2(\mem[20][5] ), 
        .ZN(n1015) );
  INV_X1 U421 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U422 ( .A1(data_in[6]), .A2(n833), .B1(n1020), .B2(\mem[20][6] ), 
        .ZN(n1014) );
  INV_X1 U423 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U424 ( .A1(data_in[7]), .A2(n833), .B1(n1020), .B2(\mem[20][7] ), 
        .ZN(n1013) );
  INV_X1 U425 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U426 ( .A1(data_in[0]), .A2(n832), .B1(n1011), .B2(\mem[21][0] ), 
        .ZN(n1012) );
  INV_X1 U427 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U428 ( .A1(data_in[1]), .A2(n832), .B1(n1011), .B2(\mem[21][1] ), 
        .ZN(n1010) );
  INV_X1 U429 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U430 ( .A1(data_in[2]), .A2(n832), .B1(n1011), .B2(\mem[21][2] ), 
        .ZN(n1009) );
  INV_X1 U431 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U432 ( .A1(data_in[3]), .A2(n832), .B1(n1011), .B2(\mem[21][3] ), 
        .ZN(n1008) );
  INV_X1 U433 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U434 ( .A1(data_in[4]), .A2(n832), .B1(n1011), .B2(\mem[21][4] ), 
        .ZN(n1007) );
  INV_X1 U435 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U436 ( .A1(data_in[5]), .A2(n832), .B1(n1011), .B2(\mem[21][5] ), 
        .ZN(n1006) );
  INV_X1 U437 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U438 ( .A1(data_in[6]), .A2(n832), .B1(n1011), .B2(\mem[21][6] ), 
        .ZN(n1005) );
  INV_X1 U439 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U440 ( .A1(data_in[7]), .A2(n832), .B1(n1011), .B2(\mem[21][7] ), 
        .ZN(n1004) );
  INV_X1 U441 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U442 ( .A1(data_in[0]), .A2(n831), .B1(n1002), .B2(\mem[22][0] ), 
        .ZN(n1003) );
  INV_X1 U443 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U444 ( .A1(data_in[1]), .A2(n831), .B1(n1002), .B2(\mem[22][1] ), 
        .ZN(n1001) );
  INV_X1 U445 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U446 ( .A1(data_in[2]), .A2(n831), .B1(n1002), .B2(\mem[22][2] ), 
        .ZN(n1000) );
  INV_X1 U447 ( .A(n999), .ZN(n706) );
  AOI22_X1 U448 ( .A1(data_in[3]), .A2(n831), .B1(n1002), .B2(\mem[22][3] ), 
        .ZN(n999) );
  INV_X1 U449 ( .A(n998), .ZN(n705) );
  AOI22_X1 U450 ( .A1(data_in[4]), .A2(n831), .B1(n1002), .B2(\mem[22][4] ), 
        .ZN(n998) );
  INV_X1 U451 ( .A(n997), .ZN(n704) );
  AOI22_X1 U452 ( .A1(data_in[5]), .A2(n831), .B1(n1002), .B2(\mem[22][5] ), 
        .ZN(n997) );
  INV_X1 U453 ( .A(n996), .ZN(n703) );
  AOI22_X1 U454 ( .A1(data_in[6]), .A2(n831), .B1(n1002), .B2(\mem[22][6] ), 
        .ZN(n996) );
  INV_X1 U455 ( .A(n995), .ZN(n702) );
  AOI22_X1 U456 ( .A1(data_in[7]), .A2(n831), .B1(n1002), .B2(\mem[22][7] ), 
        .ZN(n995) );
  INV_X1 U457 ( .A(n994), .ZN(n701) );
  AOI22_X1 U458 ( .A1(data_in[0]), .A2(n830), .B1(n993), .B2(\mem[23][0] ), 
        .ZN(n994) );
  INV_X1 U459 ( .A(n992), .ZN(n700) );
  AOI22_X1 U460 ( .A1(data_in[1]), .A2(n830), .B1(n993), .B2(\mem[23][1] ), 
        .ZN(n992) );
  INV_X1 U461 ( .A(n991), .ZN(n699) );
  AOI22_X1 U462 ( .A1(data_in[2]), .A2(n830), .B1(n993), .B2(\mem[23][2] ), 
        .ZN(n991) );
  INV_X1 U463 ( .A(n990), .ZN(n698) );
  AOI22_X1 U464 ( .A1(data_in[3]), .A2(n830), .B1(n993), .B2(\mem[23][3] ), 
        .ZN(n990) );
  INV_X1 U465 ( .A(n989), .ZN(n697) );
  AOI22_X1 U466 ( .A1(data_in[4]), .A2(n830), .B1(n993), .B2(\mem[23][4] ), 
        .ZN(n989) );
  INV_X1 U467 ( .A(n988), .ZN(n696) );
  AOI22_X1 U468 ( .A1(data_in[5]), .A2(n830), .B1(n993), .B2(\mem[23][5] ), 
        .ZN(n988) );
  INV_X1 U469 ( .A(n987), .ZN(n695) );
  AOI22_X1 U470 ( .A1(data_in[6]), .A2(n830), .B1(n993), .B2(\mem[23][6] ), 
        .ZN(n987) );
  INV_X1 U471 ( .A(n986), .ZN(n694) );
  AOI22_X1 U472 ( .A1(data_in[7]), .A2(n830), .B1(n993), .B2(\mem[23][7] ), 
        .ZN(n986) );
  INV_X1 U473 ( .A(n985), .ZN(n693) );
  AOI22_X1 U474 ( .A1(data_in[0]), .A2(n829), .B1(n984), .B2(\mem[24][0] ), 
        .ZN(n985) );
  INV_X1 U475 ( .A(n983), .ZN(n692) );
  AOI22_X1 U476 ( .A1(data_in[1]), .A2(n829), .B1(n984), .B2(\mem[24][1] ), 
        .ZN(n983) );
  INV_X1 U477 ( .A(n982), .ZN(n691) );
  AOI22_X1 U478 ( .A1(data_in[2]), .A2(n829), .B1(n984), .B2(\mem[24][2] ), 
        .ZN(n982) );
  INV_X1 U479 ( .A(n981), .ZN(n690) );
  AOI22_X1 U480 ( .A1(data_in[3]), .A2(n829), .B1(n984), .B2(\mem[24][3] ), 
        .ZN(n981) );
  INV_X1 U481 ( .A(n980), .ZN(n689) );
  AOI22_X1 U482 ( .A1(data_in[4]), .A2(n829), .B1(n984), .B2(\mem[24][4] ), 
        .ZN(n980) );
  INV_X1 U483 ( .A(n979), .ZN(n688) );
  AOI22_X1 U484 ( .A1(data_in[5]), .A2(n829), .B1(n984), .B2(\mem[24][5] ), 
        .ZN(n979) );
  INV_X1 U485 ( .A(n978), .ZN(n687) );
  AOI22_X1 U486 ( .A1(data_in[6]), .A2(n829), .B1(n984), .B2(\mem[24][6] ), 
        .ZN(n978) );
  INV_X1 U487 ( .A(n977), .ZN(n686) );
  AOI22_X1 U488 ( .A1(data_in[7]), .A2(n829), .B1(n984), .B2(\mem[24][7] ), 
        .ZN(n977) );
  INV_X1 U489 ( .A(n975), .ZN(n685) );
  AOI22_X1 U490 ( .A1(data_in[0]), .A2(n828), .B1(n974), .B2(\mem[25][0] ), 
        .ZN(n975) );
  INV_X1 U491 ( .A(n973), .ZN(n684) );
  AOI22_X1 U492 ( .A1(data_in[1]), .A2(n828), .B1(n974), .B2(\mem[25][1] ), 
        .ZN(n973) );
  INV_X1 U493 ( .A(n972), .ZN(n683) );
  AOI22_X1 U494 ( .A1(data_in[2]), .A2(n828), .B1(n974), .B2(\mem[25][2] ), 
        .ZN(n972) );
  INV_X1 U495 ( .A(n971), .ZN(n682) );
  AOI22_X1 U496 ( .A1(data_in[3]), .A2(n828), .B1(n974), .B2(\mem[25][3] ), 
        .ZN(n971) );
  INV_X1 U497 ( .A(n970), .ZN(n681) );
  AOI22_X1 U498 ( .A1(data_in[4]), .A2(n828), .B1(n974), .B2(\mem[25][4] ), 
        .ZN(n970) );
  INV_X1 U499 ( .A(n969), .ZN(n680) );
  AOI22_X1 U500 ( .A1(data_in[5]), .A2(n828), .B1(n974), .B2(\mem[25][5] ), 
        .ZN(n969) );
  INV_X1 U501 ( .A(n968), .ZN(n679) );
  AOI22_X1 U502 ( .A1(data_in[6]), .A2(n828), .B1(n974), .B2(\mem[25][6] ), 
        .ZN(n968) );
  INV_X1 U503 ( .A(n967), .ZN(n678) );
  AOI22_X1 U504 ( .A1(data_in[7]), .A2(n828), .B1(n974), .B2(\mem[25][7] ), 
        .ZN(n967) );
  INV_X1 U505 ( .A(n966), .ZN(n677) );
  AOI22_X1 U506 ( .A1(data_in[0]), .A2(n827), .B1(n965), .B2(\mem[26][0] ), 
        .ZN(n966) );
  INV_X1 U507 ( .A(n964), .ZN(n676) );
  AOI22_X1 U508 ( .A1(data_in[1]), .A2(n827), .B1(n965), .B2(\mem[26][1] ), 
        .ZN(n964) );
  INV_X1 U509 ( .A(n963), .ZN(n675) );
  AOI22_X1 U510 ( .A1(data_in[2]), .A2(n827), .B1(n965), .B2(\mem[26][2] ), 
        .ZN(n963) );
  INV_X1 U511 ( .A(n962), .ZN(n674) );
  AOI22_X1 U512 ( .A1(data_in[3]), .A2(n827), .B1(n965), .B2(\mem[26][3] ), 
        .ZN(n962) );
  INV_X1 U513 ( .A(n961), .ZN(n673) );
  AOI22_X1 U514 ( .A1(data_in[4]), .A2(n827), .B1(n965), .B2(\mem[26][4] ), 
        .ZN(n961) );
  INV_X1 U515 ( .A(n960), .ZN(n672) );
  AOI22_X1 U516 ( .A1(data_in[5]), .A2(n827), .B1(n965), .B2(\mem[26][5] ), 
        .ZN(n960) );
  INV_X1 U517 ( .A(n959), .ZN(n671) );
  AOI22_X1 U518 ( .A1(data_in[6]), .A2(n827), .B1(n965), .B2(\mem[26][6] ), 
        .ZN(n959) );
  INV_X1 U519 ( .A(n958), .ZN(n670) );
  AOI22_X1 U520 ( .A1(data_in[7]), .A2(n827), .B1(n965), .B2(\mem[26][7] ), 
        .ZN(n958) );
  INV_X1 U521 ( .A(n957), .ZN(n669) );
  AOI22_X1 U522 ( .A1(data_in[0]), .A2(n826), .B1(n956), .B2(\mem[27][0] ), 
        .ZN(n957) );
  INV_X1 U523 ( .A(n955), .ZN(n668) );
  AOI22_X1 U524 ( .A1(data_in[1]), .A2(n826), .B1(n956), .B2(\mem[27][1] ), 
        .ZN(n955) );
  INV_X1 U525 ( .A(n954), .ZN(n667) );
  AOI22_X1 U526 ( .A1(data_in[2]), .A2(n826), .B1(n956), .B2(\mem[27][2] ), 
        .ZN(n954) );
  INV_X1 U527 ( .A(n953), .ZN(n666) );
  AOI22_X1 U528 ( .A1(data_in[3]), .A2(n826), .B1(n956), .B2(\mem[27][3] ), 
        .ZN(n953) );
  INV_X1 U529 ( .A(n952), .ZN(n665) );
  AOI22_X1 U530 ( .A1(data_in[4]), .A2(n826), .B1(n956), .B2(\mem[27][4] ), 
        .ZN(n952) );
  INV_X1 U531 ( .A(n951), .ZN(n664) );
  AOI22_X1 U532 ( .A1(data_in[5]), .A2(n826), .B1(n956), .B2(\mem[27][5] ), 
        .ZN(n951) );
  INV_X1 U533 ( .A(n950), .ZN(n663) );
  AOI22_X1 U534 ( .A1(data_in[6]), .A2(n826), .B1(n956), .B2(\mem[27][6] ), 
        .ZN(n950) );
  INV_X1 U535 ( .A(n949), .ZN(n662) );
  AOI22_X1 U536 ( .A1(data_in[7]), .A2(n826), .B1(n956), .B2(\mem[27][7] ), 
        .ZN(n949) );
  INV_X1 U537 ( .A(n948), .ZN(n661) );
  AOI22_X1 U538 ( .A1(data_in[0]), .A2(n825), .B1(n947), .B2(\mem[28][0] ), 
        .ZN(n948) );
  INV_X1 U539 ( .A(n946), .ZN(n660) );
  AOI22_X1 U540 ( .A1(data_in[1]), .A2(n825), .B1(n947), .B2(\mem[28][1] ), 
        .ZN(n946) );
  INV_X1 U541 ( .A(n945), .ZN(n659) );
  AOI22_X1 U542 ( .A1(data_in[2]), .A2(n825), .B1(n947), .B2(\mem[28][2] ), 
        .ZN(n945) );
  INV_X1 U543 ( .A(n944), .ZN(n658) );
  AOI22_X1 U544 ( .A1(data_in[3]), .A2(n825), .B1(n947), .B2(\mem[28][3] ), 
        .ZN(n944) );
  INV_X1 U545 ( .A(n943), .ZN(n657) );
  AOI22_X1 U546 ( .A1(data_in[4]), .A2(n825), .B1(n947), .B2(\mem[28][4] ), 
        .ZN(n943) );
  INV_X1 U547 ( .A(n942), .ZN(n656) );
  AOI22_X1 U548 ( .A1(data_in[5]), .A2(n825), .B1(n947), .B2(\mem[28][5] ), 
        .ZN(n942) );
  INV_X1 U549 ( .A(n941), .ZN(n655) );
  AOI22_X1 U550 ( .A1(data_in[6]), .A2(n825), .B1(n947), .B2(\mem[28][6] ), 
        .ZN(n941) );
  INV_X1 U551 ( .A(n940), .ZN(n654) );
  AOI22_X1 U552 ( .A1(data_in[7]), .A2(n825), .B1(n947), .B2(\mem[28][7] ), 
        .ZN(n940) );
  INV_X1 U553 ( .A(n939), .ZN(n653) );
  AOI22_X1 U554 ( .A1(data_in[0]), .A2(n824), .B1(n938), .B2(\mem[29][0] ), 
        .ZN(n939) );
  INV_X1 U555 ( .A(n937), .ZN(n652) );
  AOI22_X1 U556 ( .A1(data_in[1]), .A2(n824), .B1(n938), .B2(\mem[29][1] ), 
        .ZN(n937) );
  INV_X1 U557 ( .A(n936), .ZN(n651) );
  AOI22_X1 U558 ( .A1(data_in[2]), .A2(n824), .B1(n938), .B2(\mem[29][2] ), 
        .ZN(n936) );
  INV_X1 U559 ( .A(n935), .ZN(n650) );
  AOI22_X1 U560 ( .A1(data_in[3]), .A2(n824), .B1(n938), .B2(\mem[29][3] ), 
        .ZN(n935) );
  INV_X1 U561 ( .A(n934), .ZN(n649) );
  AOI22_X1 U562 ( .A1(data_in[4]), .A2(n824), .B1(n938), .B2(\mem[29][4] ), 
        .ZN(n934) );
  INV_X1 U563 ( .A(n933), .ZN(n648) );
  AOI22_X1 U564 ( .A1(data_in[5]), .A2(n824), .B1(n938), .B2(\mem[29][5] ), 
        .ZN(n933) );
  INV_X1 U565 ( .A(n932), .ZN(n647) );
  AOI22_X1 U566 ( .A1(data_in[6]), .A2(n824), .B1(n938), .B2(\mem[29][6] ), 
        .ZN(n932) );
  INV_X1 U567 ( .A(n931), .ZN(n646) );
  AOI22_X1 U568 ( .A1(data_in[7]), .A2(n824), .B1(n938), .B2(\mem[29][7] ), 
        .ZN(n931) );
  INV_X1 U569 ( .A(n930), .ZN(n645) );
  AOI22_X1 U570 ( .A1(data_in[0]), .A2(n823), .B1(n929), .B2(\mem[30][0] ), 
        .ZN(n930) );
  INV_X1 U571 ( .A(n928), .ZN(n644) );
  AOI22_X1 U572 ( .A1(data_in[1]), .A2(n823), .B1(n929), .B2(\mem[30][1] ), 
        .ZN(n928) );
  INV_X1 U573 ( .A(n927), .ZN(n643) );
  AOI22_X1 U574 ( .A1(data_in[2]), .A2(n823), .B1(n929), .B2(\mem[30][2] ), 
        .ZN(n927) );
  INV_X1 U575 ( .A(n926), .ZN(n642) );
  AOI22_X1 U576 ( .A1(data_in[3]), .A2(n823), .B1(n929), .B2(\mem[30][3] ), 
        .ZN(n926) );
  INV_X1 U577 ( .A(n925), .ZN(n641) );
  AOI22_X1 U578 ( .A1(data_in[4]), .A2(n823), .B1(n929), .B2(\mem[30][4] ), 
        .ZN(n925) );
  INV_X1 U579 ( .A(n924), .ZN(n640) );
  AOI22_X1 U580 ( .A1(data_in[5]), .A2(n823), .B1(n929), .B2(\mem[30][5] ), 
        .ZN(n924) );
  INV_X1 U581 ( .A(n923), .ZN(n639) );
  AOI22_X1 U582 ( .A1(data_in[6]), .A2(n823), .B1(n929), .B2(\mem[30][6] ), 
        .ZN(n923) );
  INV_X1 U583 ( .A(n922), .ZN(n638) );
  AOI22_X1 U584 ( .A1(data_in[7]), .A2(n823), .B1(n929), .B2(\mem[30][7] ), 
        .ZN(n922) );
  INV_X1 U585 ( .A(n921), .ZN(n637) );
  AOI22_X1 U586 ( .A1(data_in[0]), .A2(n822), .B1(n920), .B2(\mem[31][0] ), 
        .ZN(n921) );
  INV_X1 U587 ( .A(n919), .ZN(n636) );
  AOI22_X1 U588 ( .A1(data_in[1]), .A2(n822), .B1(n920), .B2(\mem[31][1] ), 
        .ZN(n919) );
  INV_X1 U589 ( .A(n918), .ZN(n635) );
  AOI22_X1 U590 ( .A1(data_in[2]), .A2(n822), .B1(n920), .B2(\mem[31][2] ), 
        .ZN(n918) );
  INV_X1 U591 ( .A(n917), .ZN(n634) );
  AOI22_X1 U592 ( .A1(data_in[3]), .A2(n822), .B1(n920), .B2(\mem[31][3] ), 
        .ZN(n917) );
  INV_X1 U593 ( .A(n916), .ZN(n633) );
  AOI22_X1 U594 ( .A1(data_in[4]), .A2(n822), .B1(n920), .B2(\mem[31][4] ), 
        .ZN(n916) );
  INV_X1 U595 ( .A(n915), .ZN(n632) );
  AOI22_X1 U596 ( .A1(data_in[5]), .A2(n822), .B1(n920), .B2(\mem[31][5] ), 
        .ZN(n915) );
  INV_X1 U597 ( .A(n914), .ZN(n631) );
  AOI22_X1 U598 ( .A1(data_in[6]), .A2(n822), .B1(n920), .B2(\mem[31][6] ), 
        .ZN(n914) );
  INV_X1 U599 ( .A(n913), .ZN(n630) );
  AOI22_X1 U600 ( .A1(data_in[7]), .A2(n822), .B1(n920), .B2(\mem[31][7] ), 
        .ZN(n913) );
  MUX2_X1 U601 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n611), .Z(n1) );
  MUX2_X1 U602 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n611), .Z(n2) );
  MUX2_X1 U603 ( .A(n2), .B(n1), .S(n608), .Z(n3) );
  MUX2_X1 U604 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n611), .Z(n4) );
  MUX2_X1 U605 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n611), .Z(n5) );
  MUX2_X1 U606 ( .A(n5), .B(n4), .S(n608), .Z(n6) );
  MUX2_X1 U607 ( .A(n6), .B(n3), .S(n606), .Z(n7) );
  MUX2_X1 U608 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n611), .Z(n8) );
  MUX2_X1 U609 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n611), .Z(n9) );
  MUX2_X1 U610 ( .A(n9), .B(n8), .S(n608), .Z(n10) );
  MUX2_X1 U611 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n611), .Z(n11) );
  MUX2_X1 U612 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n611), .Z(n12) );
  MUX2_X1 U613 ( .A(n12), .B(n11), .S(n608), .Z(n13) );
  MUX2_X1 U614 ( .A(n13), .B(n10), .S(n606), .Z(n14) );
  MUX2_X1 U615 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U616 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n612), .Z(n16) );
  MUX2_X1 U617 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n612), .Z(n17) );
  MUX2_X1 U618 ( .A(n17), .B(n16), .S(n608), .Z(n18) );
  MUX2_X1 U619 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n612), .Z(n19) );
  MUX2_X1 U620 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n612), .Z(n20) );
  MUX2_X1 U621 ( .A(n20), .B(n19), .S(n609), .Z(n21) );
  MUX2_X1 U622 ( .A(n21), .B(n18), .S(n606), .Z(n22) );
  MUX2_X1 U623 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n612), .Z(n23) );
  MUX2_X1 U624 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n612), .Z(n24) );
  MUX2_X1 U625 ( .A(n24), .B(n23), .S(n610), .Z(n25) );
  MUX2_X1 U626 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n612), .Z(n26) );
  MUX2_X1 U627 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n612), .Z(n27) );
  MUX2_X1 U628 ( .A(n27), .B(n26), .S(N11), .Z(n28) );
  MUX2_X1 U629 ( .A(n28), .B(n25), .S(n606), .Z(n29) );
  MUX2_X1 U630 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U631 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U632 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n612), .Z(n31) );
  MUX2_X1 U633 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n612), .Z(n32) );
  MUX2_X1 U634 ( .A(n32), .B(n31), .S(n608), .Z(n33) );
  MUX2_X1 U635 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n612), .Z(n34) );
  MUX2_X1 U636 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n612), .Z(n35) );
  MUX2_X1 U637 ( .A(n35), .B(n34), .S(n608), .Z(n36) );
  MUX2_X1 U638 ( .A(n36), .B(n33), .S(n606), .Z(n37) );
  MUX2_X1 U639 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n613), .Z(n38) );
  MUX2_X1 U640 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n613), .Z(n39) );
  MUX2_X1 U641 ( .A(n39), .B(n38), .S(n608), .Z(n40) );
  MUX2_X1 U642 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n613), .Z(n41) );
  MUX2_X1 U643 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n613), .Z(n42) );
  MUX2_X1 U644 ( .A(n42), .B(n41), .S(n608), .Z(n43) );
  MUX2_X1 U645 ( .A(n43), .B(n40), .S(n606), .Z(n44) );
  MUX2_X1 U646 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U647 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n613), .Z(n46) );
  MUX2_X1 U648 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n613), .Z(n47) );
  MUX2_X1 U649 ( .A(n47), .B(n46), .S(n608), .Z(n48) );
  MUX2_X1 U650 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n613), .Z(n49) );
  MUX2_X1 U651 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n613), .Z(n50) );
  MUX2_X1 U652 ( .A(n50), .B(n49), .S(n608), .Z(n51) );
  MUX2_X1 U653 ( .A(n51), .B(n48), .S(n606), .Z(n52) );
  MUX2_X1 U654 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n613), .Z(n53) );
  MUX2_X1 U655 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n613), .Z(n54) );
  MUX2_X1 U656 ( .A(n54), .B(n53), .S(n608), .Z(n55) );
  MUX2_X1 U657 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n613), .Z(n56) );
  MUX2_X1 U658 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n613), .Z(n57) );
  MUX2_X1 U659 ( .A(n57), .B(n56), .S(n610), .Z(n58) );
  MUX2_X1 U660 ( .A(n58), .B(n55), .S(n606), .Z(n59) );
  MUX2_X1 U661 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U662 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U663 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n614), .Z(n61) );
  MUX2_X1 U664 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n614), .Z(n62) );
  MUX2_X1 U665 ( .A(n62), .B(n61), .S(n609), .Z(n63) );
  MUX2_X1 U666 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n614), .Z(n64) );
  MUX2_X1 U667 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n614), .Z(n65) );
  MUX2_X1 U668 ( .A(n65), .B(n64), .S(n609), .Z(n66) );
  MUX2_X1 U669 ( .A(n66), .B(n63), .S(n607), .Z(n67) );
  MUX2_X1 U670 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n614), .Z(n68) );
  MUX2_X1 U671 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n614), .Z(n69) );
  MUX2_X1 U672 ( .A(n69), .B(n68), .S(n609), .Z(n70) );
  MUX2_X1 U673 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n614), .Z(n71) );
  MUX2_X1 U674 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n614), .Z(n72) );
  MUX2_X1 U675 ( .A(n72), .B(n71), .S(n609), .Z(n73) );
  MUX2_X1 U676 ( .A(n73), .B(n70), .S(n607), .Z(n74) );
  MUX2_X1 U677 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U678 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n614), .Z(n76) );
  MUX2_X1 U679 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n614), .Z(n77) );
  MUX2_X1 U680 ( .A(n77), .B(n76), .S(n609), .Z(n78) );
  MUX2_X1 U681 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n614), .Z(n79) );
  MUX2_X1 U682 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n614), .Z(n80) );
  MUX2_X1 U683 ( .A(n80), .B(n79), .S(n609), .Z(n81) );
  MUX2_X1 U684 ( .A(n81), .B(n78), .S(n607), .Z(n82) );
  MUX2_X1 U685 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n615), .Z(n83) );
  MUX2_X1 U686 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n615), .Z(n84) );
  MUX2_X1 U687 ( .A(n84), .B(n83), .S(n609), .Z(n85) );
  MUX2_X1 U688 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n615), .Z(n86) );
  MUX2_X1 U689 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n615), .Z(n87) );
  MUX2_X1 U690 ( .A(n87), .B(n86), .S(n609), .Z(n88) );
  MUX2_X1 U691 ( .A(n88), .B(n85), .S(n607), .Z(n89) );
  MUX2_X1 U692 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U693 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U694 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n615), .Z(n91) );
  MUX2_X1 U695 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n615), .Z(n92) );
  MUX2_X1 U696 ( .A(n92), .B(n91), .S(n609), .Z(n93) );
  MUX2_X1 U697 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n615), .Z(n94) );
  MUX2_X1 U698 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n615), .Z(n95) );
  MUX2_X1 U699 ( .A(n95), .B(n94), .S(n609), .Z(n96) );
  MUX2_X1 U700 ( .A(n96), .B(n93), .S(n607), .Z(n97) );
  MUX2_X1 U701 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n615), .Z(n98) );
  MUX2_X1 U702 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n615), .Z(n99) );
  MUX2_X1 U703 ( .A(n99), .B(n98), .S(n609), .Z(n100) );
  MUX2_X1 U704 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n615), .Z(n101) );
  MUX2_X1 U705 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n615), .Z(n102) );
  MUX2_X1 U706 ( .A(n102), .B(n101), .S(n609), .Z(n103) );
  MUX2_X1 U707 ( .A(n103), .B(n100), .S(n607), .Z(n104) );
  MUX2_X1 U708 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U709 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n619), .Z(n106) );
  MUX2_X1 U710 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(N10), .Z(n107) );
  MUX2_X1 U711 ( .A(n107), .B(n106), .S(n610), .Z(n108) );
  MUX2_X1 U712 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(N10), .Z(n109) );
  MUX2_X1 U713 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n110) );
  MUX2_X1 U714 ( .A(n110), .B(n109), .S(n608), .Z(n111) );
  MUX2_X1 U715 ( .A(n111), .B(n108), .S(n607), .Z(n112) );
  MUX2_X1 U716 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n619), .Z(n113) );
  MUX2_X1 U717 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n618), .Z(n114) );
  MUX2_X1 U718 ( .A(n114), .B(n113), .S(n609), .Z(n115) );
  MUX2_X1 U719 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n618), .Z(n116) );
  MUX2_X1 U720 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n618), .Z(n117) );
  MUX2_X1 U721 ( .A(n117), .B(n116), .S(n610), .Z(n118) );
  MUX2_X1 U722 ( .A(n118), .B(n115), .S(n607), .Z(n119) );
  MUX2_X1 U723 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U724 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U725 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(N10), .Z(n121) );
  MUX2_X1 U726 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n619), .Z(n122) );
  MUX2_X1 U727 ( .A(n122), .B(n121), .S(n609), .Z(n123) );
  MUX2_X1 U728 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n618), .Z(n124) );
  MUX2_X1 U729 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n619), .Z(n125) );
  MUX2_X1 U730 ( .A(n125), .B(n124), .S(n608), .Z(n126) );
  MUX2_X1 U731 ( .A(n126), .B(n123), .S(n607), .Z(n127) );
  MUX2_X1 U732 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n611), .Z(n128) );
  MUX2_X1 U733 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n611), .Z(n129) );
  MUX2_X1 U734 ( .A(n129), .B(n128), .S(n609), .Z(n130) );
  MUX2_X1 U735 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n611), .Z(n131) );
  MUX2_X1 U736 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n618), .Z(n132) );
  MUX2_X1 U737 ( .A(n132), .B(n131), .S(n609), .Z(n133) );
  MUX2_X1 U738 ( .A(n133), .B(n130), .S(n607), .Z(n134) );
  MUX2_X1 U739 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U740 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n616), .Z(n136) );
  MUX2_X1 U741 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n619), .Z(n137) );
  MUX2_X1 U742 ( .A(n137), .B(n136), .S(N11), .Z(n138) );
  MUX2_X1 U743 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n614), .Z(n139) );
  MUX2_X1 U744 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n619), .Z(n140) );
  MUX2_X1 U745 ( .A(n140), .B(n139), .S(n610), .Z(n141) );
  MUX2_X1 U746 ( .A(n141), .B(n138), .S(n607), .Z(n142) );
  MUX2_X1 U747 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n611), .Z(n143) );
  MUX2_X1 U748 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n617), .Z(n144) );
  MUX2_X1 U749 ( .A(n144), .B(n143), .S(n609), .Z(n145) );
  MUX2_X1 U750 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n618), .Z(n146) );
  MUX2_X1 U751 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n147) );
  MUX2_X1 U752 ( .A(n147), .B(n146), .S(n608), .Z(n148) );
  MUX2_X1 U753 ( .A(n148), .B(n145), .S(n607), .Z(n149) );
  MUX2_X1 U754 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U755 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U756 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n616), .Z(n151) );
  MUX2_X1 U757 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n616), .Z(n152) );
  MUX2_X1 U758 ( .A(n152), .B(n151), .S(n610), .Z(n153) );
  MUX2_X1 U759 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n616), .Z(n154) );
  MUX2_X1 U760 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n616), .Z(n155) );
  MUX2_X1 U761 ( .A(n155), .B(n154), .S(n610), .Z(n156) );
  MUX2_X1 U762 ( .A(n156), .B(n153), .S(n606), .Z(n157) );
  MUX2_X1 U763 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n616), .Z(n158) );
  MUX2_X1 U764 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n616), .Z(n159) );
  MUX2_X1 U765 ( .A(n159), .B(n158), .S(n610), .Z(n160) );
  MUX2_X1 U766 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n616), .Z(n161) );
  MUX2_X1 U767 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n616), .Z(n162) );
  MUX2_X1 U768 ( .A(n162), .B(n161), .S(n610), .Z(n163) );
  MUX2_X1 U769 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U770 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U771 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n616), .Z(n166) );
  MUX2_X1 U772 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n616), .Z(n167) );
  MUX2_X1 U773 ( .A(n167), .B(n166), .S(n610), .Z(n168) );
  MUX2_X1 U774 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n616), .Z(n169) );
  MUX2_X1 U775 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n616), .Z(n170) );
  MUX2_X1 U776 ( .A(n170), .B(n169), .S(n610), .Z(n171) );
  MUX2_X1 U777 ( .A(n171), .B(n168), .S(n606), .Z(n172) );
  MUX2_X1 U778 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n617), .Z(n173) );
  MUX2_X1 U779 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n617), .Z(n174) );
  MUX2_X1 U780 ( .A(n174), .B(n173), .S(n610), .Z(n175) );
  MUX2_X1 U781 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n617), .Z(n176) );
  MUX2_X1 U782 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n617), .Z(n177) );
  MUX2_X1 U783 ( .A(n177), .B(n176), .S(n610), .Z(n178) );
  MUX2_X1 U784 ( .A(n178), .B(n175), .S(n606), .Z(n179) );
  MUX2_X1 U785 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U786 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U787 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n617), .Z(n181) );
  MUX2_X1 U788 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n617), .Z(n182) );
  MUX2_X1 U789 ( .A(n182), .B(n181), .S(n610), .Z(n183) );
  MUX2_X1 U790 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n617), .Z(n184) );
  MUX2_X1 U791 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n617), .Z(n185) );
  MUX2_X1 U792 ( .A(n185), .B(n184), .S(n610), .Z(n186) );
  MUX2_X1 U793 ( .A(n186), .B(n183), .S(n606), .Z(n187) );
  MUX2_X1 U794 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n617), .Z(n188) );
  MUX2_X1 U795 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n617), .Z(n189) );
  MUX2_X1 U796 ( .A(n189), .B(n188), .S(n610), .Z(n190) );
  MUX2_X1 U797 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n617), .Z(n191) );
  MUX2_X1 U798 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n617), .Z(n192) );
  MUX2_X1 U799 ( .A(n192), .B(n191), .S(n610), .Z(n193) );
  MUX2_X1 U800 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U801 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U802 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n618), .Z(n196) );
  MUX2_X1 U803 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n618), .Z(n197) );
  MUX2_X1 U804 ( .A(n197), .B(n196), .S(n608), .Z(n198) );
  MUX2_X1 U805 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n619), .Z(n199) );
  MUX2_X1 U806 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n619), .Z(n200) );
  MUX2_X1 U807 ( .A(n200), .B(n199), .S(N11), .Z(n201) );
  MUX2_X1 U808 ( .A(n201), .B(n198), .S(n606), .Z(n202) );
  MUX2_X1 U809 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n615), .Z(n203) );
  MUX2_X1 U810 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n619), .Z(n204) );
  MUX2_X1 U811 ( .A(n204), .B(n203), .S(n609), .Z(n205) );
  MUX2_X1 U812 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n618), .Z(n206) );
  MUX2_X1 U813 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n618), .Z(n207) );
  MUX2_X1 U814 ( .A(n207), .B(n206), .S(n610), .Z(n208) );
  MUX2_X1 U815 ( .A(n208), .B(n205), .S(n607), .Z(n209) );
  MUX2_X1 U816 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U817 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U818 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n614), .Z(n211) );
  MUX2_X1 U819 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n618), .Z(n212) );
  MUX2_X1 U820 ( .A(n212), .B(n211), .S(n608), .Z(n213) );
  MUX2_X1 U821 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n619), .Z(n214) );
  MUX2_X1 U822 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n619), .Z(n215) );
  MUX2_X1 U823 ( .A(n215), .B(n214), .S(n610), .Z(n216) );
  MUX2_X1 U824 ( .A(n216), .B(n213), .S(n606), .Z(n217) );
  MUX2_X1 U825 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n619), .Z(n218) );
  MUX2_X1 U826 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n619), .Z(n219) );
  MUX2_X1 U827 ( .A(n219), .B(n218), .S(n608), .Z(n220) );
  MUX2_X1 U828 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n612), .Z(n221) );
  MUX2_X1 U829 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n619), .Z(n222) );
  MUX2_X1 U830 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U831 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U832 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U833 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n616), .Z(n226) );
  MUX2_X1 U834 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n618), .Z(n227) );
  MUX2_X1 U835 ( .A(n227), .B(n226), .S(n610), .Z(n228) );
  MUX2_X1 U836 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n613), .Z(n229) );
  MUX2_X1 U837 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n617), .Z(n595) );
  MUX2_X1 U838 ( .A(n595), .B(n229), .S(N11), .Z(n596) );
  MUX2_X1 U839 ( .A(n596), .B(n228), .S(n607), .Z(n597) );
  MUX2_X1 U840 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n611), .Z(n598) );
  MUX2_X1 U841 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n618), .Z(n599) );
  MUX2_X1 U842 ( .A(n599), .B(n598), .S(n608), .Z(n600) );
  MUX2_X1 U843 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n619), .Z(n601) );
  MUX2_X1 U844 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n618), .Z(n602) );
  MUX2_X1 U845 ( .A(n602), .B(n601), .S(n608), .Z(n603) );
  MUX2_X1 U846 ( .A(n603), .B(n600), .S(n606), .Z(n604) );
  MUX2_X1 U847 ( .A(n604), .B(n597), .S(N13), .Z(n605) );
  MUX2_X1 U848 ( .A(n605), .B(n225), .S(N14), .Z(N15) );
  INV_X1 U849 ( .A(N10), .ZN(n620) );
  INV_X1 U850 ( .A(N11), .ZN(n621) );
  INV_X1 U851 ( .A(data_in[0]), .ZN(n622) );
  INV_X1 U852 ( .A(data_in[1]), .ZN(n623) );
  INV_X1 U853 ( .A(data_in[2]), .ZN(n624) );
  INV_X1 U854 ( .A(data_in[3]), .ZN(n625) );
  INV_X1 U855 ( .A(data_in[4]), .ZN(n626) );
  INV_X1 U856 ( .A(data_in[5]), .ZN(n627) );
  INV_X1 U857 ( .A(data_in[6]), .ZN(n628) );
  INV_X1 U858 ( .A(data_in[7]), .ZN(n629) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_1 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n630), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n631), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n632), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n633), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n634), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n635), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n636), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n637), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n638), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n639), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n640), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n641), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n642), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n643), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n644), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n645), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n646), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n647), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n648), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n649), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n650), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n651), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n652), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n653), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n654), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n655), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n656), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n657), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n658), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n659), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n660), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n661), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n662), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n663), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n664), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n665), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n666), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n667), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n668), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n669), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n670), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n671), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n672), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n673), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n674), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n675), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n676), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n677), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n678), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n679), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n680), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n681), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n682), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n683), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n684), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n685), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n686), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n687), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n688), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n689), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n690), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n691), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n692), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n693), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n694), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n695), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n696), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n697), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n698), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n699), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n700), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n701), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n702), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n703), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n704), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n705), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n706), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n707), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n708), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n709), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n710), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n711), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n712), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n713), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n714), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n715), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n716), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n717), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n718), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n719), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n720), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n721), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n722), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n723), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n724), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n725), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n726), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n727), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n728), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n729), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n730), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n731), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n732), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n733), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n734), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n735), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n736), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n737), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n738), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n739), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n740), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n741), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n742), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n743), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n744), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n745), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n746), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n747), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n748), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n749), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n750), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n751), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n752), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n753), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n754), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n755), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n756), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n757), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n758), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n759), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n760), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n761), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n762), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n763), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n764), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n765), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n766), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n767), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n768), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n769), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n770), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n771), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n772), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n773), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n774), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n775), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n776), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n777), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n778), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n779), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n780), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n781), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n782), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n783), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n784), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n785), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n786), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n787), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n788), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n789), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n790), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n791), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n792), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n793), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n794), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n795), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n796), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n797), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n798), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n799), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n800), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n801), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n802), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n803), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n804), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n805), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n806), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n807), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n808), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n809), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n810), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n811), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n812), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n813), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n814), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n815), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n816), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n817), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n818), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n819), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n820), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n821), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n849), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n850), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n851), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n852), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n853), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n854), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n855), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n856), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n857), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n858), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n859), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n860), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n861), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n862), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n863), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n864), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n865), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n866), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n867), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n868), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n869), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n870), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n871), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n872), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n873), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n874), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n875), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n876), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n877), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n878), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n879), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n880), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n881), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n882), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n883), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n884), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n885), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n886), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n887), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n888), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n889), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n890), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n891), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n892), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n893), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n894), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n895), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n896), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n897), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n898), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n899), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n900), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n901), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n902), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n903), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n904), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n905), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n906), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n907), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n908), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n909), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n910), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n911), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n912), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .QN(n2) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  NOR2_X1 U3 ( .A1(n846), .A2(addr[5]), .ZN(n1132) );
  AND3_X1 U4 ( .A1(n847), .A2(n848), .A3(n1132), .ZN(n1203) );
  AND3_X1 U5 ( .A1(n1132), .A2(n848), .A3(N13), .ZN(n1122) );
  AND3_X1 U6 ( .A1(n1132), .A2(n847), .A3(N14), .ZN(n1049) );
  AND3_X1 U7 ( .A1(N13), .A2(n1132), .A3(N14), .ZN(n976) );
  INV_X2 U8 ( .A(n2), .ZN(data_out[1]) );
  BUF_X1 U9 ( .A(n619), .Z(n617) );
  BUF_X1 U10 ( .A(n619), .Z(n618) );
  BUF_X1 U11 ( .A(N10), .Z(n615) );
  BUF_X1 U12 ( .A(n619), .Z(n616) );
  BUF_X1 U13 ( .A(N11), .Z(n612) );
  BUF_X1 U14 ( .A(N11), .Z(n613) );
  BUF_X1 U15 ( .A(N10), .Z(n619) );
  NOR3_X1 U16 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1204) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(n620), .ZN(n1193) );
  NOR3_X1 U18 ( .A1(N10), .A2(N12), .A3(n621), .ZN(n1183) );
  NOR3_X1 U19 ( .A1(n620), .A2(N12), .A3(n621), .ZN(n1173) );
  INV_X1 U20 ( .A(n1130), .ZN(n845) );
  INV_X1 U21 ( .A(n1120), .ZN(n844) );
  INV_X1 U22 ( .A(n1111), .ZN(n843) );
  INV_X1 U23 ( .A(n1102), .ZN(n842) );
  INV_X1 U24 ( .A(n1057), .ZN(n837) );
  INV_X1 U25 ( .A(n1047), .ZN(n836) );
  INV_X1 U26 ( .A(n1038), .ZN(n835) );
  INV_X1 U27 ( .A(n1029), .ZN(n834) );
  INV_X1 U28 ( .A(n984), .ZN(n829) );
  INV_X1 U29 ( .A(n974), .ZN(n828) );
  INV_X1 U30 ( .A(n965), .ZN(n827) );
  INV_X1 U31 ( .A(n956), .ZN(n826) );
  INV_X1 U32 ( .A(n1093), .ZN(n841) );
  INV_X1 U33 ( .A(n1084), .ZN(n840) );
  INV_X1 U34 ( .A(n1075), .ZN(n839) );
  INV_X1 U35 ( .A(n1066), .ZN(n838) );
  INV_X1 U36 ( .A(n947), .ZN(n825) );
  INV_X1 U37 ( .A(n938), .ZN(n824) );
  INV_X1 U38 ( .A(n929), .ZN(n823) );
  INV_X1 U39 ( .A(n920), .ZN(n822) );
  INV_X1 U40 ( .A(n1020), .ZN(n833) );
  INV_X1 U41 ( .A(n1011), .ZN(n832) );
  INV_X1 U42 ( .A(n1002), .ZN(n831) );
  INV_X1 U43 ( .A(n993), .ZN(n830) );
  BUF_X1 U44 ( .A(N12), .Z(n610) );
  INV_X1 U45 ( .A(N13), .ZN(n847) );
  AND3_X1 U46 ( .A1(n620), .A2(n621), .A3(N12), .ZN(n1163) );
  AND3_X1 U47 ( .A1(N10), .A2(n621), .A3(N12), .ZN(n1153) );
  AND3_X1 U48 ( .A1(N11), .A2(n620), .A3(N12), .ZN(n1143) );
  AND3_X1 U49 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1133) );
  BUF_X1 U50 ( .A(N12), .Z(n609) );
  INV_X1 U51 ( .A(N14), .ZN(n848) );
  NAND2_X1 U52 ( .A1(n1193), .A2(n1203), .ZN(n1202) );
  NAND2_X1 U53 ( .A1(n1183), .A2(n1203), .ZN(n1192) );
  NAND2_X1 U54 ( .A1(n1173), .A2(n1203), .ZN(n1182) );
  NAND2_X1 U55 ( .A1(n1163), .A2(n1203), .ZN(n1172) );
  NAND2_X1 U56 ( .A1(n1153), .A2(n1203), .ZN(n1162) );
  NAND2_X1 U57 ( .A1(n1143), .A2(n1203), .ZN(n1152) );
  NAND2_X1 U58 ( .A1(n1133), .A2(n1203), .ZN(n1142) );
  NAND2_X1 U59 ( .A1(n1204), .A2(n1203), .ZN(n1213) );
  NAND2_X1 U60 ( .A1(n1122), .A2(n1204), .ZN(n1130) );
  NAND2_X1 U61 ( .A1(n1122), .A2(n1193), .ZN(n1120) );
  NAND2_X1 U62 ( .A1(n1122), .A2(n1183), .ZN(n1111) );
  NAND2_X1 U63 ( .A1(n1122), .A2(n1173), .ZN(n1102) );
  NAND2_X1 U64 ( .A1(n1049), .A2(n1204), .ZN(n1057) );
  NAND2_X1 U65 ( .A1(n1049), .A2(n1193), .ZN(n1047) );
  NAND2_X1 U66 ( .A1(n1049), .A2(n1183), .ZN(n1038) );
  NAND2_X1 U67 ( .A1(n1049), .A2(n1173), .ZN(n1029) );
  NAND2_X1 U68 ( .A1(n976), .A2(n1204), .ZN(n984) );
  NAND2_X1 U69 ( .A1(n976), .A2(n1193), .ZN(n974) );
  NAND2_X1 U70 ( .A1(n976), .A2(n1183), .ZN(n965) );
  NAND2_X1 U71 ( .A1(n976), .A2(n1173), .ZN(n956) );
  NAND2_X1 U72 ( .A1(n1122), .A2(n1163), .ZN(n1093) );
  NAND2_X1 U73 ( .A1(n1122), .A2(n1153), .ZN(n1084) );
  NAND2_X1 U74 ( .A1(n1122), .A2(n1143), .ZN(n1075) );
  NAND2_X1 U75 ( .A1(n1122), .A2(n1133), .ZN(n1066) );
  NAND2_X1 U76 ( .A1(n1049), .A2(n1163), .ZN(n1020) );
  NAND2_X1 U77 ( .A1(n1049), .A2(n1153), .ZN(n1011) );
  NAND2_X1 U78 ( .A1(n1049), .A2(n1143), .ZN(n1002) );
  NAND2_X1 U79 ( .A1(n1049), .A2(n1133), .ZN(n993) );
  NAND2_X1 U80 ( .A1(n976), .A2(n1163), .ZN(n947) );
  NAND2_X1 U81 ( .A1(n976), .A2(n1153), .ZN(n938) );
  NAND2_X1 U82 ( .A1(n976), .A2(n1143), .ZN(n929) );
  NAND2_X1 U83 ( .A1(n976), .A2(n1133), .ZN(n920) );
  INV_X1 U84 ( .A(wr_en), .ZN(n846) );
  OAI21_X1 U85 ( .B1(n1213), .B2(n622), .A(n1212), .ZN(n912) );
  NAND2_X1 U86 ( .A1(\mem[0][0] ), .A2(n1213), .ZN(n1212) );
  OAI21_X1 U87 ( .B1(n1213), .B2(n623), .A(n1211), .ZN(n911) );
  NAND2_X1 U88 ( .A1(\mem[0][1] ), .A2(n1213), .ZN(n1211) );
  OAI21_X1 U89 ( .B1(n1213), .B2(n624), .A(n1210), .ZN(n910) );
  NAND2_X1 U90 ( .A1(\mem[0][2] ), .A2(n1213), .ZN(n1210) );
  OAI21_X1 U91 ( .B1(n1213), .B2(n625), .A(n1209), .ZN(n909) );
  NAND2_X1 U92 ( .A1(\mem[0][3] ), .A2(n1213), .ZN(n1209) );
  OAI21_X1 U93 ( .B1(n1213), .B2(n626), .A(n1208), .ZN(n908) );
  NAND2_X1 U94 ( .A1(\mem[0][4] ), .A2(n1213), .ZN(n1208) );
  OAI21_X1 U95 ( .B1(n1213), .B2(n627), .A(n1207), .ZN(n907) );
  NAND2_X1 U96 ( .A1(\mem[0][5] ), .A2(n1213), .ZN(n1207) );
  OAI21_X1 U97 ( .B1(n1213), .B2(n628), .A(n1206), .ZN(n906) );
  NAND2_X1 U98 ( .A1(\mem[0][6] ), .A2(n1213), .ZN(n1206) );
  OAI21_X1 U99 ( .B1(n1213), .B2(n629), .A(n1205), .ZN(n905) );
  NAND2_X1 U100 ( .A1(\mem[0][7] ), .A2(n1213), .ZN(n1205) );
  OAI21_X1 U101 ( .B1(n622), .B2(n1172), .A(n1171), .ZN(n880) );
  NAND2_X1 U102 ( .A1(\mem[4][0] ), .A2(n1172), .ZN(n1171) );
  OAI21_X1 U103 ( .B1(n623), .B2(n1172), .A(n1170), .ZN(n879) );
  NAND2_X1 U104 ( .A1(\mem[4][1] ), .A2(n1172), .ZN(n1170) );
  OAI21_X1 U105 ( .B1(n624), .B2(n1172), .A(n1169), .ZN(n878) );
  NAND2_X1 U106 ( .A1(\mem[4][2] ), .A2(n1172), .ZN(n1169) );
  OAI21_X1 U107 ( .B1(n625), .B2(n1172), .A(n1168), .ZN(n877) );
  NAND2_X1 U108 ( .A1(\mem[4][3] ), .A2(n1172), .ZN(n1168) );
  OAI21_X1 U109 ( .B1(n626), .B2(n1172), .A(n1167), .ZN(n876) );
  NAND2_X1 U110 ( .A1(\mem[4][4] ), .A2(n1172), .ZN(n1167) );
  OAI21_X1 U111 ( .B1(n627), .B2(n1172), .A(n1166), .ZN(n875) );
  NAND2_X1 U112 ( .A1(\mem[4][5] ), .A2(n1172), .ZN(n1166) );
  OAI21_X1 U113 ( .B1(n628), .B2(n1172), .A(n1165), .ZN(n874) );
  NAND2_X1 U114 ( .A1(\mem[4][6] ), .A2(n1172), .ZN(n1165) );
  OAI21_X1 U115 ( .B1(n629), .B2(n1172), .A(n1164), .ZN(n873) );
  NAND2_X1 U116 ( .A1(\mem[4][7] ), .A2(n1172), .ZN(n1164) );
  OAI21_X1 U117 ( .B1(n622), .B2(n1152), .A(n1151), .ZN(n864) );
  NAND2_X1 U118 ( .A1(\mem[6][0] ), .A2(n1152), .ZN(n1151) );
  OAI21_X1 U119 ( .B1(n623), .B2(n1152), .A(n1150), .ZN(n863) );
  NAND2_X1 U120 ( .A1(\mem[6][1] ), .A2(n1152), .ZN(n1150) );
  OAI21_X1 U121 ( .B1(n624), .B2(n1152), .A(n1149), .ZN(n862) );
  NAND2_X1 U122 ( .A1(\mem[6][2] ), .A2(n1152), .ZN(n1149) );
  OAI21_X1 U123 ( .B1(n625), .B2(n1152), .A(n1148), .ZN(n861) );
  NAND2_X1 U124 ( .A1(\mem[6][3] ), .A2(n1152), .ZN(n1148) );
  OAI21_X1 U125 ( .B1(n626), .B2(n1152), .A(n1147), .ZN(n860) );
  NAND2_X1 U126 ( .A1(\mem[6][4] ), .A2(n1152), .ZN(n1147) );
  OAI21_X1 U127 ( .B1(n627), .B2(n1152), .A(n1146), .ZN(n859) );
  NAND2_X1 U128 ( .A1(\mem[6][5] ), .A2(n1152), .ZN(n1146) );
  OAI21_X1 U129 ( .B1(n628), .B2(n1152), .A(n1145), .ZN(n858) );
  NAND2_X1 U130 ( .A1(\mem[6][6] ), .A2(n1152), .ZN(n1145) );
  OAI21_X1 U131 ( .B1(n629), .B2(n1152), .A(n1144), .ZN(n857) );
  NAND2_X1 U132 ( .A1(\mem[6][7] ), .A2(n1152), .ZN(n1144) );
  OAI21_X1 U133 ( .B1(n622), .B2(n1142), .A(n1141), .ZN(n856) );
  NAND2_X1 U134 ( .A1(\mem[7][0] ), .A2(n1142), .ZN(n1141) );
  OAI21_X1 U135 ( .B1(n623), .B2(n1142), .A(n1140), .ZN(n855) );
  NAND2_X1 U136 ( .A1(\mem[7][1] ), .A2(n1142), .ZN(n1140) );
  OAI21_X1 U137 ( .B1(n624), .B2(n1142), .A(n1139), .ZN(n854) );
  NAND2_X1 U138 ( .A1(\mem[7][2] ), .A2(n1142), .ZN(n1139) );
  OAI21_X1 U139 ( .B1(n625), .B2(n1142), .A(n1138), .ZN(n853) );
  NAND2_X1 U140 ( .A1(\mem[7][3] ), .A2(n1142), .ZN(n1138) );
  OAI21_X1 U141 ( .B1(n626), .B2(n1142), .A(n1137), .ZN(n852) );
  NAND2_X1 U142 ( .A1(\mem[7][4] ), .A2(n1142), .ZN(n1137) );
  OAI21_X1 U143 ( .B1(n627), .B2(n1142), .A(n1136), .ZN(n851) );
  NAND2_X1 U144 ( .A1(\mem[7][5] ), .A2(n1142), .ZN(n1136) );
  OAI21_X1 U145 ( .B1(n628), .B2(n1142), .A(n1135), .ZN(n850) );
  NAND2_X1 U146 ( .A1(\mem[7][6] ), .A2(n1142), .ZN(n1135) );
  OAI21_X1 U147 ( .B1(n629), .B2(n1142), .A(n1134), .ZN(n849) );
  NAND2_X1 U148 ( .A1(\mem[7][7] ), .A2(n1142), .ZN(n1134) );
  OAI21_X1 U149 ( .B1(n622), .B2(n1202), .A(n1201), .ZN(n904) );
  NAND2_X1 U150 ( .A1(\mem[1][0] ), .A2(n1202), .ZN(n1201) );
  OAI21_X1 U151 ( .B1(n623), .B2(n1202), .A(n1200), .ZN(n903) );
  NAND2_X1 U152 ( .A1(\mem[1][1] ), .A2(n1202), .ZN(n1200) );
  OAI21_X1 U153 ( .B1(n624), .B2(n1202), .A(n1199), .ZN(n902) );
  NAND2_X1 U154 ( .A1(\mem[1][2] ), .A2(n1202), .ZN(n1199) );
  OAI21_X1 U155 ( .B1(n625), .B2(n1202), .A(n1198), .ZN(n901) );
  NAND2_X1 U156 ( .A1(\mem[1][3] ), .A2(n1202), .ZN(n1198) );
  OAI21_X1 U157 ( .B1(n626), .B2(n1202), .A(n1197), .ZN(n900) );
  NAND2_X1 U158 ( .A1(\mem[1][4] ), .A2(n1202), .ZN(n1197) );
  OAI21_X1 U159 ( .B1(n627), .B2(n1202), .A(n1196), .ZN(n899) );
  NAND2_X1 U160 ( .A1(\mem[1][5] ), .A2(n1202), .ZN(n1196) );
  OAI21_X1 U161 ( .B1(n628), .B2(n1202), .A(n1195), .ZN(n898) );
  NAND2_X1 U162 ( .A1(\mem[1][6] ), .A2(n1202), .ZN(n1195) );
  OAI21_X1 U163 ( .B1(n629), .B2(n1202), .A(n1194), .ZN(n897) );
  NAND2_X1 U164 ( .A1(\mem[1][7] ), .A2(n1202), .ZN(n1194) );
  OAI21_X1 U165 ( .B1(n622), .B2(n1192), .A(n1191), .ZN(n896) );
  NAND2_X1 U166 ( .A1(\mem[2][0] ), .A2(n1192), .ZN(n1191) );
  OAI21_X1 U167 ( .B1(n623), .B2(n1192), .A(n1190), .ZN(n895) );
  NAND2_X1 U168 ( .A1(\mem[2][1] ), .A2(n1192), .ZN(n1190) );
  OAI21_X1 U169 ( .B1(n624), .B2(n1192), .A(n1189), .ZN(n894) );
  NAND2_X1 U170 ( .A1(\mem[2][2] ), .A2(n1192), .ZN(n1189) );
  OAI21_X1 U171 ( .B1(n625), .B2(n1192), .A(n1188), .ZN(n893) );
  NAND2_X1 U172 ( .A1(\mem[2][3] ), .A2(n1192), .ZN(n1188) );
  OAI21_X1 U173 ( .B1(n626), .B2(n1192), .A(n1187), .ZN(n892) );
  NAND2_X1 U174 ( .A1(\mem[2][4] ), .A2(n1192), .ZN(n1187) );
  OAI21_X1 U175 ( .B1(n627), .B2(n1192), .A(n1186), .ZN(n891) );
  NAND2_X1 U176 ( .A1(\mem[2][5] ), .A2(n1192), .ZN(n1186) );
  OAI21_X1 U177 ( .B1(n628), .B2(n1192), .A(n1185), .ZN(n890) );
  NAND2_X1 U178 ( .A1(\mem[2][6] ), .A2(n1192), .ZN(n1185) );
  OAI21_X1 U179 ( .B1(n629), .B2(n1192), .A(n1184), .ZN(n889) );
  NAND2_X1 U180 ( .A1(\mem[2][7] ), .A2(n1192), .ZN(n1184) );
  OAI21_X1 U181 ( .B1(n622), .B2(n1182), .A(n1181), .ZN(n888) );
  NAND2_X1 U182 ( .A1(\mem[3][0] ), .A2(n1182), .ZN(n1181) );
  OAI21_X1 U183 ( .B1(n623), .B2(n1182), .A(n1180), .ZN(n887) );
  NAND2_X1 U184 ( .A1(\mem[3][1] ), .A2(n1182), .ZN(n1180) );
  OAI21_X1 U185 ( .B1(n624), .B2(n1182), .A(n1179), .ZN(n886) );
  NAND2_X1 U186 ( .A1(\mem[3][2] ), .A2(n1182), .ZN(n1179) );
  OAI21_X1 U187 ( .B1(n625), .B2(n1182), .A(n1178), .ZN(n885) );
  NAND2_X1 U188 ( .A1(\mem[3][3] ), .A2(n1182), .ZN(n1178) );
  OAI21_X1 U189 ( .B1(n626), .B2(n1182), .A(n1177), .ZN(n884) );
  NAND2_X1 U190 ( .A1(\mem[3][4] ), .A2(n1182), .ZN(n1177) );
  OAI21_X1 U191 ( .B1(n627), .B2(n1182), .A(n1176), .ZN(n883) );
  NAND2_X1 U192 ( .A1(\mem[3][5] ), .A2(n1182), .ZN(n1176) );
  OAI21_X1 U193 ( .B1(n628), .B2(n1182), .A(n1175), .ZN(n882) );
  NAND2_X1 U194 ( .A1(\mem[3][6] ), .A2(n1182), .ZN(n1175) );
  OAI21_X1 U195 ( .B1(n629), .B2(n1182), .A(n1174), .ZN(n881) );
  NAND2_X1 U196 ( .A1(\mem[3][7] ), .A2(n1182), .ZN(n1174) );
  OAI21_X1 U197 ( .B1(n622), .B2(n1162), .A(n1161), .ZN(n872) );
  NAND2_X1 U198 ( .A1(\mem[5][0] ), .A2(n1162), .ZN(n1161) );
  OAI21_X1 U199 ( .B1(n623), .B2(n1162), .A(n1160), .ZN(n871) );
  NAND2_X1 U200 ( .A1(\mem[5][1] ), .A2(n1162), .ZN(n1160) );
  OAI21_X1 U201 ( .B1(n624), .B2(n1162), .A(n1159), .ZN(n870) );
  NAND2_X1 U202 ( .A1(\mem[5][2] ), .A2(n1162), .ZN(n1159) );
  OAI21_X1 U203 ( .B1(n625), .B2(n1162), .A(n1158), .ZN(n869) );
  NAND2_X1 U204 ( .A1(\mem[5][3] ), .A2(n1162), .ZN(n1158) );
  OAI21_X1 U205 ( .B1(n626), .B2(n1162), .A(n1157), .ZN(n868) );
  NAND2_X1 U206 ( .A1(\mem[5][4] ), .A2(n1162), .ZN(n1157) );
  OAI21_X1 U207 ( .B1(n627), .B2(n1162), .A(n1156), .ZN(n867) );
  NAND2_X1 U208 ( .A1(\mem[5][5] ), .A2(n1162), .ZN(n1156) );
  OAI21_X1 U209 ( .B1(n628), .B2(n1162), .A(n1155), .ZN(n866) );
  NAND2_X1 U210 ( .A1(\mem[5][6] ), .A2(n1162), .ZN(n1155) );
  OAI21_X1 U211 ( .B1(n629), .B2(n1162), .A(n1154), .ZN(n865) );
  NAND2_X1 U212 ( .A1(\mem[5][7] ), .A2(n1162), .ZN(n1154) );
  INV_X1 U213 ( .A(n1131), .ZN(n821) );
  AOI22_X1 U214 ( .A1(data_in[0]), .A2(n845), .B1(n1130), .B2(\mem[8][0] ), 
        .ZN(n1131) );
  INV_X1 U215 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U216 ( .A1(data_in[1]), .A2(n845), .B1(n1130), .B2(\mem[8][1] ), 
        .ZN(n1129) );
  INV_X1 U217 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U218 ( .A1(data_in[2]), .A2(n845), .B1(n1130), .B2(\mem[8][2] ), 
        .ZN(n1128) );
  INV_X1 U219 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U220 ( .A1(data_in[3]), .A2(n845), .B1(n1130), .B2(\mem[8][3] ), 
        .ZN(n1127) );
  INV_X1 U221 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U222 ( .A1(data_in[4]), .A2(n845), .B1(n1130), .B2(\mem[8][4] ), 
        .ZN(n1126) );
  INV_X1 U223 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U224 ( .A1(data_in[5]), .A2(n845), .B1(n1130), .B2(\mem[8][5] ), 
        .ZN(n1125) );
  INV_X1 U225 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U226 ( .A1(data_in[6]), .A2(n845), .B1(n1130), .B2(\mem[8][6] ), 
        .ZN(n1124) );
  INV_X1 U227 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U228 ( .A1(data_in[7]), .A2(n845), .B1(n1130), .B2(\mem[8][7] ), 
        .ZN(n1123) );
  INV_X1 U229 ( .A(n1121), .ZN(n813) );
  AOI22_X1 U230 ( .A1(data_in[0]), .A2(n844), .B1(n1120), .B2(\mem[9][0] ), 
        .ZN(n1121) );
  INV_X1 U231 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U232 ( .A1(data_in[1]), .A2(n844), .B1(n1120), .B2(\mem[9][1] ), 
        .ZN(n1119) );
  INV_X1 U233 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U234 ( .A1(data_in[2]), .A2(n844), .B1(n1120), .B2(\mem[9][2] ), 
        .ZN(n1118) );
  INV_X1 U235 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U236 ( .A1(data_in[3]), .A2(n844), .B1(n1120), .B2(\mem[9][3] ), 
        .ZN(n1117) );
  INV_X1 U237 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U238 ( .A1(data_in[4]), .A2(n844), .B1(n1120), .B2(\mem[9][4] ), 
        .ZN(n1116) );
  INV_X1 U239 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U240 ( .A1(data_in[5]), .A2(n844), .B1(n1120), .B2(\mem[9][5] ), 
        .ZN(n1115) );
  INV_X1 U241 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U242 ( .A1(data_in[6]), .A2(n844), .B1(n1120), .B2(\mem[9][6] ), 
        .ZN(n1114) );
  INV_X1 U243 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U244 ( .A1(data_in[7]), .A2(n844), .B1(n1120), .B2(\mem[9][7] ), 
        .ZN(n1113) );
  INV_X1 U245 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U246 ( .A1(data_in[0]), .A2(n843), .B1(n1111), .B2(\mem[10][0] ), 
        .ZN(n1112) );
  INV_X1 U247 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U248 ( .A1(data_in[1]), .A2(n843), .B1(n1111), .B2(\mem[10][1] ), 
        .ZN(n1110) );
  INV_X1 U249 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U250 ( .A1(data_in[2]), .A2(n843), .B1(n1111), .B2(\mem[10][2] ), 
        .ZN(n1109) );
  INV_X1 U251 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U252 ( .A1(data_in[3]), .A2(n843), .B1(n1111), .B2(\mem[10][3] ), 
        .ZN(n1108) );
  INV_X1 U253 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U254 ( .A1(data_in[4]), .A2(n843), .B1(n1111), .B2(\mem[10][4] ), 
        .ZN(n1107) );
  INV_X1 U255 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U256 ( .A1(data_in[5]), .A2(n843), .B1(n1111), .B2(\mem[10][5] ), 
        .ZN(n1106) );
  INV_X1 U257 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U258 ( .A1(data_in[6]), .A2(n843), .B1(n1111), .B2(\mem[10][6] ), 
        .ZN(n1105) );
  INV_X1 U259 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U260 ( .A1(data_in[7]), .A2(n843), .B1(n1111), .B2(\mem[10][7] ), 
        .ZN(n1104) );
  INV_X1 U261 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U262 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[11][0] ), 
        .ZN(n1103) );
  INV_X1 U263 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U264 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[11][1] ), 
        .ZN(n1101) );
  INV_X1 U265 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U266 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[11][2] ), 
        .ZN(n1100) );
  INV_X1 U267 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U268 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[11][3] ), 
        .ZN(n1099) );
  INV_X1 U269 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U270 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[11][4] ), 
        .ZN(n1098) );
  INV_X1 U271 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U272 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[11][5] ), 
        .ZN(n1097) );
  INV_X1 U273 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U274 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[11][6] ), 
        .ZN(n1096) );
  INV_X1 U275 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U276 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[11][7] ), 
        .ZN(n1095) );
  INV_X1 U277 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U278 ( .A1(data_in[0]), .A2(n841), .B1(n1093), .B2(\mem[12][0] ), 
        .ZN(n1094) );
  INV_X1 U279 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U280 ( .A1(data_in[1]), .A2(n841), .B1(n1093), .B2(\mem[12][1] ), 
        .ZN(n1092) );
  INV_X1 U281 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U282 ( .A1(data_in[2]), .A2(n841), .B1(n1093), .B2(\mem[12][2] ), 
        .ZN(n1091) );
  INV_X1 U283 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U284 ( .A1(data_in[3]), .A2(n841), .B1(n1093), .B2(\mem[12][3] ), 
        .ZN(n1090) );
  INV_X1 U285 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U286 ( .A1(data_in[4]), .A2(n841), .B1(n1093), .B2(\mem[12][4] ), 
        .ZN(n1089) );
  INV_X1 U287 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U288 ( .A1(data_in[5]), .A2(n841), .B1(n1093), .B2(\mem[12][5] ), 
        .ZN(n1088) );
  INV_X1 U289 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U290 ( .A1(data_in[6]), .A2(n841), .B1(n1093), .B2(\mem[12][6] ), 
        .ZN(n1087) );
  INV_X1 U291 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U292 ( .A1(data_in[7]), .A2(n841), .B1(n1093), .B2(\mem[12][7] ), 
        .ZN(n1086) );
  INV_X1 U293 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U294 ( .A1(data_in[0]), .A2(n840), .B1(n1084), .B2(\mem[13][0] ), 
        .ZN(n1085) );
  INV_X1 U295 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U296 ( .A1(data_in[1]), .A2(n840), .B1(n1084), .B2(\mem[13][1] ), 
        .ZN(n1083) );
  INV_X1 U297 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U298 ( .A1(data_in[2]), .A2(n840), .B1(n1084), .B2(\mem[13][2] ), 
        .ZN(n1082) );
  INV_X1 U299 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U300 ( .A1(data_in[3]), .A2(n840), .B1(n1084), .B2(\mem[13][3] ), 
        .ZN(n1081) );
  INV_X1 U301 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U302 ( .A1(data_in[4]), .A2(n840), .B1(n1084), .B2(\mem[13][4] ), 
        .ZN(n1080) );
  INV_X1 U303 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U304 ( .A1(data_in[5]), .A2(n840), .B1(n1084), .B2(\mem[13][5] ), 
        .ZN(n1079) );
  INV_X1 U305 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U306 ( .A1(data_in[6]), .A2(n840), .B1(n1084), .B2(\mem[13][6] ), 
        .ZN(n1078) );
  INV_X1 U307 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U308 ( .A1(data_in[7]), .A2(n840), .B1(n1084), .B2(\mem[13][7] ), 
        .ZN(n1077) );
  INV_X1 U309 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U310 ( .A1(data_in[0]), .A2(n839), .B1(n1075), .B2(\mem[14][0] ), 
        .ZN(n1076) );
  INV_X1 U311 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U312 ( .A1(data_in[1]), .A2(n839), .B1(n1075), .B2(\mem[14][1] ), 
        .ZN(n1074) );
  INV_X1 U313 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U314 ( .A1(data_in[2]), .A2(n839), .B1(n1075), .B2(\mem[14][2] ), 
        .ZN(n1073) );
  INV_X1 U315 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U316 ( .A1(data_in[3]), .A2(n839), .B1(n1075), .B2(\mem[14][3] ), 
        .ZN(n1072) );
  INV_X1 U317 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U318 ( .A1(data_in[4]), .A2(n839), .B1(n1075), .B2(\mem[14][4] ), 
        .ZN(n1071) );
  INV_X1 U319 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U320 ( .A1(data_in[5]), .A2(n839), .B1(n1075), .B2(\mem[14][5] ), 
        .ZN(n1070) );
  INV_X1 U321 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U322 ( .A1(data_in[6]), .A2(n839), .B1(n1075), .B2(\mem[14][6] ), 
        .ZN(n1069) );
  INV_X1 U323 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U324 ( .A1(data_in[7]), .A2(n839), .B1(n1075), .B2(\mem[14][7] ), 
        .ZN(n1068) );
  INV_X1 U325 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U326 ( .A1(data_in[0]), .A2(n838), .B1(n1066), .B2(\mem[15][0] ), 
        .ZN(n1067) );
  INV_X1 U327 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U328 ( .A1(data_in[1]), .A2(n838), .B1(n1066), .B2(\mem[15][1] ), 
        .ZN(n1065) );
  INV_X1 U329 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U330 ( .A1(data_in[2]), .A2(n838), .B1(n1066), .B2(\mem[15][2] ), 
        .ZN(n1064) );
  INV_X1 U331 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U332 ( .A1(data_in[3]), .A2(n838), .B1(n1066), .B2(\mem[15][3] ), 
        .ZN(n1063) );
  INV_X1 U333 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U334 ( .A1(data_in[4]), .A2(n838), .B1(n1066), .B2(\mem[15][4] ), 
        .ZN(n1062) );
  INV_X1 U335 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U336 ( .A1(data_in[5]), .A2(n838), .B1(n1066), .B2(\mem[15][5] ), 
        .ZN(n1061) );
  INV_X1 U337 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U338 ( .A1(data_in[6]), .A2(n838), .B1(n1066), .B2(\mem[15][6] ), 
        .ZN(n1060) );
  INV_X1 U339 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U340 ( .A1(data_in[7]), .A2(n838), .B1(n1066), .B2(\mem[15][7] ), 
        .ZN(n1059) );
  INV_X1 U341 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U342 ( .A1(data_in[0]), .A2(n837), .B1(n1057), .B2(\mem[16][0] ), 
        .ZN(n1058) );
  INV_X1 U343 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U344 ( .A1(data_in[1]), .A2(n837), .B1(n1057), .B2(\mem[16][1] ), 
        .ZN(n1056) );
  INV_X1 U345 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U346 ( .A1(data_in[2]), .A2(n837), .B1(n1057), .B2(\mem[16][2] ), 
        .ZN(n1055) );
  INV_X1 U347 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U348 ( .A1(data_in[3]), .A2(n837), .B1(n1057), .B2(\mem[16][3] ), 
        .ZN(n1054) );
  INV_X1 U349 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U350 ( .A1(data_in[4]), .A2(n837), .B1(n1057), .B2(\mem[16][4] ), 
        .ZN(n1053) );
  INV_X1 U351 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U352 ( .A1(data_in[5]), .A2(n837), .B1(n1057), .B2(\mem[16][5] ), 
        .ZN(n1052) );
  INV_X1 U353 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U354 ( .A1(data_in[6]), .A2(n837), .B1(n1057), .B2(\mem[16][6] ), 
        .ZN(n1051) );
  INV_X1 U355 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U356 ( .A1(data_in[7]), .A2(n837), .B1(n1057), .B2(\mem[16][7] ), 
        .ZN(n1050) );
  INV_X1 U357 ( .A(n1048), .ZN(n749) );
  AOI22_X1 U358 ( .A1(data_in[0]), .A2(n836), .B1(n1047), .B2(\mem[17][0] ), 
        .ZN(n1048) );
  INV_X1 U359 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U360 ( .A1(data_in[1]), .A2(n836), .B1(n1047), .B2(\mem[17][1] ), 
        .ZN(n1046) );
  INV_X1 U361 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U362 ( .A1(data_in[2]), .A2(n836), .B1(n1047), .B2(\mem[17][2] ), 
        .ZN(n1045) );
  INV_X1 U363 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U364 ( .A1(data_in[3]), .A2(n836), .B1(n1047), .B2(\mem[17][3] ), 
        .ZN(n1044) );
  INV_X1 U365 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U366 ( .A1(data_in[4]), .A2(n836), .B1(n1047), .B2(\mem[17][4] ), 
        .ZN(n1043) );
  INV_X1 U367 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U368 ( .A1(data_in[5]), .A2(n836), .B1(n1047), .B2(\mem[17][5] ), 
        .ZN(n1042) );
  INV_X1 U369 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U370 ( .A1(data_in[6]), .A2(n836), .B1(n1047), .B2(\mem[17][6] ), 
        .ZN(n1041) );
  INV_X1 U371 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U372 ( .A1(data_in[7]), .A2(n836), .B1(n1047), .B2(\mem[17][7] ), 
        .ZN(n1040) );
  INV_X1 U373 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U374 ( .A1(data_in[0]), .A2(n835), .B1(n1038), .B2(\mem[18][0] ), 
        .ZN(n1039) );
  INV_X1 U375 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U376 ( .A1(data_in[1]), .A2(n835), .B1(n1038), .B2(\mem[18][1] ), 
        .ZN(n1037) );
  INV_X1 U377 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U378 ( .A1(data_in[2]), .A2(n835), .B1(n1038), .B2(\mem[18][2] ), 
        .ZN(n1036) );
  INV_X1 U379 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U380 ( .A1(data_in[3]), .A2(n835), .B1(n1038), .B2(\mem[18][3] ), 
        .ZN(n1035) );
  INV_X1 U381 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U382 ( .A1(data_in[4]), .A2(n835), .B1(n1038), .B2(\mem[18][4] ), 
        .ZN(n1034) );
  INV_X1 U383 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U384 ( .A1(data_in[5]), .A2(n835), .B1(n1038), .B2(\mem[18][5] ), 
        .ZN(n1033) );
  INV_X1 U385 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U386 ( .A1(data_in[6]), .A2(n835), .B1(n1038), .B2(\mem[18][6] ), 
        .ZN(n1032) );
  INV_X1 U387 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U388 ( .A1(data_in[7]), .A2(n835), .B1(n1038), .B2(\mem[18][7] ), 
        .ZN(n1031) );
  INV_X1 U389 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U390 ( .A1(data_in[0]), .A2(n834), .B1(n1029), .B2(\mem[19][0] ), 
        .ZN(n1030) );
  INV_X1 U391 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U392 ( .A1(data_in[1]), .A2(n834), .B1(n1029), .B2(\mem[19][1] ), 
        .ZN(n1028) );
  INV_X1 U393 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U394 ( .A1(data_in[2]), .A2(n834), .B1(n1029), .B2(\mem[19][2] ), 
        .ZN(n1027) );
  INV_X1 U395 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U396 ( .A1(data_in[3]), .A2(n834), .B1(n1029), .B2(\mem[19][3] ), 
        .ZN(n1026) );
  INV_X1 U397 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U398 ( .A1(data_in[4]), .A2(n834), .B1(n1029), .B2(\mem[19][4] ), 
        .ZN(n1025) );
  INV_X1 U399 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U400 ( .A1(data_in[5]), .A2(n834), .B1(n1029), .B2(\mem[19][5] ), 
        .ZN(n1024) );
  INV_X1 U401 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U402 ( .A1(data_in[6]), .A2(n834), .B1(n1029), .B2(\mem[19][6] ), 
        .ZN(n1023) );
  INV_X1 U403 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U404 ( .A1(data_in[7]), .A2(n834), .B1(n1029), .B2(\mem[19][7] ), 
        .ZN(n1022) );
  INV_X1 U405 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U406 ( .A1(data_in[0]), .A2(n833), .B1(n1020), .B2(\mem[20][0] ), 
        .ZN(n1021) );
  INV_X1 U407 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U408 ( .A1(data_in[1]), .A2(n833), .B1(n1020), .B2(\mem[20][1] ), 
        .ZN(n1019) );
  INV_X1 U409 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U410 ( .A1(data_in[2]), .A2(n833), .B1(n1020), .B2(\mem[20][2] ), 
        .ZN(n1018) );
  INV_X1 U411 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U412 ( .A1(data_in[3]), .A2(n833), .B1(n1020), .B2(\mem[20][3] ), 
        .ZN(n1017) );
  INV_X1 U413 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U414 ( .A1(data_in[4]), .A2(n833), .B1(n1020), .B2(\mem[20][4] ), 
        .ZN(n1016) );
  INV_X1 U415 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U416 ( .A1(data_in[5]), .A2(n833), .B1(n1020), .B2(\mem[20][5] ), 
        .ZN(n1015) );
  INV_X1 U417 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U418 ( .A1(data_in[6]), .A2(n833), .B1(n1020), .B2(\mem[20][6] ), 
        .ZN(n1014) );
  INV_X1 U419 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U420 ( .A1(data_in[7]), .A2(n833), .B1(n1020), .B2(\mem[20][7] ), 
        .ZN(n1013) );
  INV_X1 U421 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U422 ( .A1(data_in[0]), .A2(n832), .B1(n1011), .B2(\mem[21][0] ), 
        .ZN(n1012) );
  INV_X1 U423 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U424 ( .A1(data_in[1]), .A2(n832), .B1(n1011), .B2(\mem[21][1] ), 
        .ZN(n1010) );
  INV_X1 U425 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U426 ( .A1(data_in[2]), .A2(n832), .B1(n1011), .B2(\mem[21][2] ), 
        .ZN(n1009) );
  INV_X1 U427 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U428 ( .A1(data_in[3]), .A2(n832), .B1(n1011), .B2(\mem[21][3] ), 
        .ZN(n1008) );
  INV_X1 U429 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U430 ( .A1(data_in[4]), .A2(n832), .B1(n1011), .B2(\mem[21][4] ), 
        .ZN(n1007) );
  INV_X1 U431 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U432 ( .A1(data_in[5]), .A2(n832), .B1(n1011), .B2(\mem[21][5] ), 
        .ZN(n1006) );
  INV_X1 U433 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U434 ( .A1(data_in[6]), .A2(n832), .B1(n1011), .B2(\mem[21][6] ), 
        .ZN(n1005) );
  INV_X1 U435 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U436 ( .A1(data_in[7]), .A2(n832), .B1(n1011), .B2(\mem[21][7] ), 
        .ZN(n1004) );
  INV_X1 U437 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U438 ( .A1(data_in[0]), .A2(n831), .B1(n1002), .B2(\mem[22][0] ), 
        .ZN(n1003) );
  INV_X1 U439 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U440 ( .A1(data_in[1]), .A2(n831), .B1(n1002), .B2(\mem[22][1] ), 
        .ZN(n1001) );
  INV_X1 U441 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U442 ( .A1(data_in[2]), .A2(n831), .B1(n1002), .B2(\mem[22][2] ), 
        .ZN(n1000) );
  INV_X1 U443 ( .A(n999), .ZN(n706) );
  AOI22_X1 U444 ( .A1(data_in[3]), .A2(n831), .B1(n1002), .B2(\mem[22][3] ), 
        .ZN(n999) );
  INV_X1 U445 ( .A(n998), .ZN(n705) );
  AOI22_X1 U446 ( .A1(data_in[4]), .A2(n831), .B1(n1002), .B2(\mem[22][4] ), 
        .ZN(n998) );
  INV_X1 U447 ( .A(n997), .ZN(n704) );
  AOI22_X1 U448 ( .A1(data_in[5]), .A2(n831), .B1(n1002), .B2(\mem[22][5] ), 
        .ZN(n997) );
  INV_X1 U449 ( .A(n996), .ZN(n703) );
  AOI22_X1 U450 ( .A1(data_in[6]), .A2(n831), .B1(n1002), .B2(\mem[22][6] ), 
        .ZN(n996) );
  INV_X1 U451 ( .A(n995), .ZN(n702) );
  AOI22_X1 U452 ( .A1(data_in[7]), .A2(n831), .B1(n1002), .B2(\mem[22][7] ), 
        .ZN(n995) );
  INV_X1 U453 ( .A(n994), .ZN(n701) );
  AOI22_X1 U454 ( .A1(data_in[0]), .A2(n830), .B1(n993), .B2(\mem[23][0] ), 
        .ZN(n994) );
  INV_X1 U455 ( .A(n992), .ZN(n700) );
  AOI22_X1 U456 ( .A1(data_in[1]), .A2(n830), .B1(n993), .B2(\mem[23][1] ), 
        .ZN(n992) );
  INV_X1 U457 ( .A(n991), .ZN(n699) );
  AOI22_X1 U458 ( .A1(data_in[2]), .A2(n830), .B1(n993), .B2(\mem[23][2] ), 
        .ZN(n991) );
  INV_X1 U459 ( .A(n990), .ZN(n698) );
  AOI22_X1 U460 ( .A1(data_in[3]), .A2(n830), .B1(n993), .B2(\mem[23][3] ), 
        .ZN(n990) );
  INV_X1 U461 ( .A(n989), .ZN(n697) );
  AOI22_X1 U462 ( .A1(data_in[4]), .A2(n830), .B1(n993), .B2(\mem[23][4] ), 
        .ZN(n989) );
  INV_X1 U463 ( .A(n988), .ZN(n696) );
  AOI22_X1 U464 ( .A1(data_in[5]), .A2(n830), .B1(n993), .B2(\mem[23][5] ), 
        .ZN(n988) );
  INV_X1 U465 ( .A(n987), .ZN(n695) );
  AOI22_X1 U466 ( .A1(data_in[6]), .A2(n830), .B1(n993), .B2(\mem[23][6] ), 
        .ZN(n987) );
  INV_X1 U467 ( .A(n986), .ZN(n694) );
  AOI22_X1 U468 ( .A1(data_in[7]), .A2(n830), .B1(n993), .B2(\mem[23][7] ), 
        .ZN(n986) );
  INV_X1 U469 ( .A(n985), .ZN(n693) );
  AOI22_X1 U470 ( .A1(data_in[0]), .A2(n829), .B1(n984), .B2(\mem[24][0] ), 
        .ZN(n985) );
  INV_X1 U471 ( .A(n983), .ZN(n692) );
  AOI22_X1 U472 ( .A1(data_in[1]), .A2(n829), .B1(n984), .B2(\mem[24][1] ), 
        .ZN(n983) );
  INV_X1 U473 ( .A(n982), .ZN(n691) );
  AOI22_X1 U474 ( .A1(data_in[2]), .A2(n829), .B1(n984), .B2(\mem[24][2] ), 
        .ZN(n982) );
  INV_X1 U475 ( .A(n981), .ZN(n690) );
  AOI22_X1 U476 ( .A1(data_in[3]), .A2(n829), .B1(n984), .B2(\mem[24][3] ), 
        .ZN(n981) );
  INV_X1 U477 ( .A(n980), .ZN(n689) );
  AOI22_X1 U478 ( .A1(data_in[4]), .A2(n829), .B1(n984), .B2(\mem[24][4] ), 
        .ZN(n980) );
  INV_X1 U479 ( .A(n979), .ZN(n688) );
  AOI22_X1 U480 ( .A1(data_in[5]), .A2(n829), .B1(n984), .B2(\mem[24][5] ), 
        .ZN(n979) );
  INV_X1 U481 ( .A(n978), .ZN(n687) );
  AOI22_X1 U482 ( .A1(data_in[6]), .A2(n829), .B1(n984), .B2(\mem[24][6] ), 
        .ZN(n978) );
  INV_X1 U483 ( .A(n977), .ZN(n686) );
  AOI22_X1 U484 ( .A1(data_in[7]), .A2(n829), .B1(n984), .B2(\mem[24][7] ), 
        .ZN(n977) );
  INV_X1 U485 ( .A(n975), .ZN(n685) );
  AOI22_X1 U486 ( .A1(data_in[0]), .A2(n828), .B1(n974), .B2(\mem[25][0] ), 
        .ZN(n975) );
  INV_X1 U487 ( .A(n973), .ZN(n684) );
  AOI22_X1 U488 ( .A1(data_in[1]), .A2(n828), .B1(n974), .B2(\mem[25][1] ), 
        .ZN(n973) );
  INV_X1 U489 ( .A(n972), .ZN(n683) );
  AOI22_X1 U490 ( .A1(data_in[2]), .A2(n828), .B1(n974), .B2(\mem[25][2] ), 
        .ZN(n972) );
  INV_X1 U491 ( .A(n971), .ZN(n682) );
  AOI22_X1 U492 ( .A1(data_in[3]), .A2(n828), .B1(n974), .B2(\mem[25][3] ), 
        .ZN(n971) );
  INV_X1 U493 ( .A(n970), .ZN(n681) );
  AOI22_X1 U494 ( .A1(data_in[4]), .A2(n828), .B1(n974), .B2(\mem[25][4] ), 
        .ZN(n970) );
  INV_X1 U495 ( .A(n969), .ZN(n680) );
  AOI22_X1 U496 ( .A1(data_in[5]), .A2(n828), .B1(n974), .B2(\mem[25][5] ), 
        .ZN(n969) );
  INV_X1 U497 ( .A(n968), .ZN(n679) );
  AOI22_X1 U498 ( .A1(data_in[6]), .A2(n828), .B1(n974), .B2(\mem[25][6] ), 
        .ZN(n968) );
  INV_X1 U499 ( .A(n967), .ZN(n678) );
  AOI22_X1 U500 ( .A1(data_in[7]), .A2(n828), .B1(n974), .B2(\mem[25][7] ), 
        .ZN(n967) );
  INV_X1 U501 ( .A(n966), .ZN(n677) );
  AOI22_X1 U502 ( .A1(data_in[0]), .A2(n827), .B1(n965), .B2(\mem[26][0] ), 
        .ZN(n966) );
  INV_X1 U503 ( .A(n964), .ZN(n676) );
  AOI22_X1 U504 ( .A1(data_in[1]), .A2(n827), .B1(n965), .B2(\mem[26][1] ), 
        .ZN(n964) );
  INV_X1 U505 ( .A(n963), .ZN(n675) );
  AOI22_X1 U506 ( .A1(data_in[2]), .A2(n827), .B1(n965), .B2(\mem[26][2] ), 
        .ZN(n963) );
  INV_X1 U507 ( .A(n962), .ZN(n674) );
  AOI22_X1 U508 ( .A1(data_in[3]), .A2(n827), .B1(n965), .B2(\mem[26][3] ), 
        .ZN(n962) );
  INV_X1 U509 ( .A(n961), .ZN(n673) );
  AOI22_X1 U510 ( .A1(data_in[4]), .A2(n827), .B1(n965), .B2(\mem[26][4] ), 
        .ZN(n961) );
  INV_X1 U511 ( .A(n960), .ZN(n672) );
  AOI22_X1 U512 ( .A1(data_in[5]), .A2(n827), .B1(n965), .B2(\mem[26][5] ), 
        .ZN(n960) );
  INV_X1 U513 ( .A(n959), .ZN(n671) );
  AOI22_X1 U514 ( .A1(data_in[6]), .A2(n827), .B1(n965), .B2(\mem[26][6] ), 
        .ZN(n959) );
  INV_X1 U515 ( .A(n958), .ZN(n670) );
  AOI22_X1 U516 ( .A1(data_in[7]), .A2(n827), .B1(n965), .B2(\mem[26][7] ), 
        .ZN(n958) );
  INV_X1 U517 ( .A(n957), .ZN(n669) );
  AOI22_X1 U518 ( .A1(data_in[0]), .A2(n826), .B1(n956), .B2(\mem[27][0] ), 
        .ZN(n957) );
  INV_X1 U519 ( .A(n955), .ZN(n668) );
  AOI22_X1 U520 ( .A1(data_in[1]), .A2(n826), .B1(n956), .B2(\mem[27][1] ), 
        .ZN(n955) );
  INV_X1 U521 ( .A(n954), .ZN(n667) );
  AOI22_X1 U522 ( .A1(data_in[2]), .A2(n826), .B1(n956), .B2(\mem[27][2] ), 
        .ZN(n954) );
  INV_X1 U523 ( .A(n953), .ZN(n666) );
  AOI22_X1 U524 ( .A1(data_in[3]), .A2(n826), .B1(n956), .B2(\mem[27][3] ), 
        .ZN(n953) );
  INV_X1 U525 ( .A(n952), .ZN(n665) );
  AOI22_X1 U526 ( .A1(data_in[4]), .A2(n826), .B1(n956), .B2(\mem[27][4] ), 
        .ZN(n952) );
  INV_X1 U527 ( .A(n951), .ZN(n664) );
  AOI22_X1 U528 ( .A1(data_in[5]), .A2(n826), .B1(n956), .B2(\mem[27][5] ), 
        .ZN(n951) );
  INV_X1 U529 ( .A(n950), .ZN(n663) );
  AOI22_X1 U530 ( .A1(data_in[6]), .A2(n826), .B1(n956), .B2(\mem[27][6] ), 
        .ZN(n950) );
  INV_X1 U531 ( .A(n949), .ZN(n662) );
  AOI22_X1 U532 ( .A1(data_in[7]), .A2(n826), .B1(n956), .B2(\mem[27][7] ), 
        .ZN(n949) );
  INV_X1 U533 ( .A(n948), .ZN(n661) );
  AOI22_X1 U534 ( .A1(data_in[0]), .A2(n825), .B1(n947), .B2(\mem[28][0] ), 
        .ZN(n948) );
  INV_X1 U535 ( .A(n946), .ZN(n660) );
  AOI22_X1 U536 ( .A1(data_in[1]), .A2(n825), .B1(n947), .B2(\mem[28][1] ), 
        .ZN(n946) );
  INV_X1 U537 ( .A(n945), .ZN(n659) );
  AOI22_X1 U538 ( .A1(data_in[2]), .A2(n825), .B1(n947), .B2(\mem[28][2] ), 
        .ZN(n945) );
  INV_X1 U539 ( .A(n944), .ZN(n658) );
  AOI22_X1 U540 ( .A1(data_in[3]), .A2(n825), .B1(n947), .B2(\mem[28][3] ), 
        .ZN(n944) );
  INV_X1 U541 ( .A(n943), .ZN(n657) );
  AOI22_X1 U542 ( .A1(data_in[4]), .A2(n825), .B1(n947), .B2(\mem[28][4] ), 
        .ZN(n943) );
  INV_X1 U543 ( .A(n942), .ZN(n656) );
  AOI22_X1 U544 ( .A1(data_in[5]), .A2(n825), .B1(n947), .B2(\mem[28][5] ), 
        .ZN(n942) );
  INV_X1 U545 ( .A(n941), .ZN(n655) );
  AOI22_X1 U546 ( .A1(data_in[6]), .A2(n825), .B1(n947), .B2(\mem[28][6] ), 
        .ZN(n941) );
  INV_X1 U547 ( .A(n940), .ZN(n654) );
  AOI22_X1 U548 ( .A1(data_in[7]), .A2(n825), .B1(n947), .B2(\mem[28][7] ), 
        .ZN(n940) );
  INV_X1 U549 ( .A(n939), .ZN(n653) );
  AOI22_X1 U550 ( .A1(data_in[0]), .A2(n824), .B1(n938), .B2(\mem[29][0] ), 
        .ZN(n939) );
  INV_X1 U551 ( .A(n937), .ZN(n652) );
  AOI22_X1 U552 ( .A1(data_in[1]), .A2(n824), .B1(n938), .B2(\mem[29][1] ), 
        .ZN(n937) );
  INV_X1 U553 ( .A(n936), .ZN(n651) );
  AOI22_X1 U554 ( .A1(data_in[2]), .A2(n824), .B1(n938), .B2(\mem[29][2] ), 
        .ZN(n936) );
  INV_X1 U555 ( .A(n935), .ZN(n650) );
  AOI22_X1 U556 ( .A1(data_in[3]), .A2(n824), .B1(n938), .B2(\mem[29][3] ), 
        .ZN(n935) );
  INV_X1 U557 ( .A(n934), .ZN(n649) );
  AOI22_X1 U558 ( .A1(data_in[4]), .A2(n824), .B1(n938), .B2(\mem[29][4] ), 
        .ZN(n934) );
  INV_X1 U559 ( .A(n933), .ZN(n648) );
  AOI22_X1 U560 ( .A1(data_in[5]), .A2(n824), .B1(n938), .B2(\mem[29][5] ), 
        .ZN(n933) );
  INV_X1 U561 ( .A(n932), .ZN(n647) );
  AOI22_X1 U562 ( .A1(data_in[6]), .A2(n824), .B1(n938), .B2(\mem[29][6] ), 
        .ZN(n932) );
  INV_X1 U563 ( .A(n931), .ZN(n646) );
  AOI22_X1 U564 ( .A1(data_in[7]), .A2(n824), .B1(n938), .B2(\mem[29][7] ), 
        .ZN(n931) );
  INV_X1 U565 ( .A(n930), .ZN(n645) );
  AOI22_X1 U566 ( .A1(data_in[0]), .A2(n823), .B1(n929), .B2(\mem[30][0] ), 
        .ZN(n930) );
  INV_X1 U567 ( .A(n928), .ZN(n644) );
  AOI22_X1 U568 ( .A1(data_in[1]), .A2(n823), .B1(n929), .B2(\mem[30][1] ), 
        .ZN(n928) );
  INV_X1 U569 ( .A(n927), .ZN(n643) );
  AOI22_X1 U570 ( .A1(data_in[2]), .A2(n823), .B1(n929), .B2(\mem[30][2] ), 
        .ZN(n927) );
  INV_X1 U571 ( .A(n926), .ZN(n642) );
  AOI22_X1 U572 ( .A1(data_in[3]), .A2(n823), .B1(n929), .B2(\mem[30][3] ), 
        .ZN(n926) );
  INV_X1 U573 ( .A(n925), .ZN(n641) );
  AOI22_X1 U574 ( .A1(data_in[4]), .A2(n823), .B1(n929), .B2(\mem[30][4] ), 
        .ZN(n925) );
  INV_X1 U575 ( .A(n924), .ZN(n640) );
  AOI22_X1 U576 ( .A1(data_in[5]), .A2(n823), .B1(n929), .B2(\mem[30][5] ), 
        .ZN(n924) );
  INV_X1 U577 ( .A(n923), .ZN(n639) );
  AOI22_X1 U578 ( .A1(data_in[6]), .A2(n823), .B1(n929), .B2(\mem[30][6] ), 
        .ZN(n923) );
  INV_X1 U579 ( .A(n922), .ZN(n638) );
  AOI22_X1 U580 ( .A1(data_in[7]), .A2(n823), .B1(n929), .B2(\mem[30][7] ), 
        .ZN(n922) );
  INV_X1 U581 ( .A(n921), .ZN(n637) );
  AOI22_X1 U582 ( .A1(data_in[0]), .A2(n822), .B1(n920), .B2(\mem[31][0] ), 
        .ZN(n921) );
  INV_X1 U583 ( .A(n919), .ZN(n636) );
  AOI22_X1 U584 ( .A1(data_in[1]), .A2(n822), .B1(n920), .B2(\mem[31][1] ), 
        .ZN(n919) );
  INV_X1 U585 ( .A(n918), .ZN(n635) );
  AOI22_X1 U586 ( .A1(data_in[2]), .A2(n822), .B1(n920), .B2(\mem[31][2] ), 
        .ZN(n918) );
  INV_X1 U587 ( .A(n917), .ZN(n634) );
  AOI22_X1 U588 ( .A1(data_in[3]), .A2(n822), .B1(n920), .B2(\mem[31][3] ), 
        .ZN(n917) );
  INV_X1 U589 ( .A(n916), .ZN(n633) );
  AOI22_X1 U590 ( .A1(data_in[4]), .A2(n822), .B1(n920), .B2(\mem[31][4] ), 
        .ZN(n916) );
  INV_X1 U591 ( .A(n915), .ZN(n632) );
  AOI22_X1 U592 ( .A1(data_in[5]), .A2(n822), .B1(n920), .B2(\mem[31][5] ), 
        .ZN(n915) );
  INV_X1 U593 ( .A(n914), .ZN(n631) );
  AOI22_X1 U594 ( .A1(data_in[6]), .A2(n822), .B1(n920), .B2(\mem[31][6] ), 
        .ZN(n914) );
  INV_X1 U595 ( .A(n913), .ZN(n630) );
  AOI22_X1 U596 ( .A1(data_in[7]), .A2(n822), .B1(n920), .B2(\mem[31][7] ), 
        .ZN(n913) );
  MUX2_X1 U597 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n614), .Z(n4) );
  MUX2_X1 U598 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n614), .Z(n5) );
  MUX2_X1 U599 ( .A(n5), .B(n4), .S(n611), .Z(n6) );
  MUX2_X1 U600 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n614), .Z(n7) );
  MUX2_X1 U601 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n614), .Z(n8) );
  MUX2_X1 U602 ( .A(n8), .B(n7), .S(n611), .Z(n9) );
  MUX2_X1 U603 ( .A(n9), .B(n6), .S(n609), .Z(n10) );
  MUX2_X1 U604 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n614), .Z(n11) );
  MUX2_X1 U605 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n614), .Z(n12) );
  MUX2_X1 U606 ( .A(n12), .B(n11), .S(n611), .Z(n13) );
  MUX2_X1 U607 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n614), .Z(n14) );
  MUX2_X1 U608 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n614), .Z(n15) );
  MUX2_X1 U609 ( .A(n15), .B(n14), .S(n611), .Z(n16) );
  MUX2_X1 U610 ( .A(n16), .B(n13), .S(n609), .Z(n17) );
  MUX2_X1 U611 ( .A(n17), .B(n10), .S(N13), .Z(n18) );
  MUX2_X1 U612 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n615), .Z(n19) );
  MUX2_X1 U613 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(N10), .Z(n20) );
  MUX2_X1 U614 ( .A(n20), .B(n19), .S(n613), .Z(n21) );
  MUX2_X1 U615 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n614), .Z(n22) );
  MUX2_X1 U616 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n614), .Z(n23) );
  MUX2_X1 U617 ( .A(n23), .B(n22), .S(n611), .Z(n24) );
  MUX2_X1 U618 ( .A(n24), .B(n21), .S(n609), .Z(n25) );
  MUX2_X1 U619 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n619), .Z(n26) );
  MUX2_X1 U620 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n27) );
  MUX2_X1 U621 ( .A(n27), .B(n26), .S(N11), .Z(n28) );
  MUX2_X1 U622 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n29) );
  MUX2_X1 U623 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n30) );
  MUX2_X1 U624 ( .A(n30), .B(n29), .S(n613), .Z(n31) );
  MUX2_X1 U625 ( .A(n31), .B(n28), .S(n609), .Z(n32) );
  MUX2_X1 U626 ( .A(n32), .B(n25), .S(N13), .Z(n33) );
  MUX2_X1 U627 ( .A(n33), .B(n18), .S(N14), .Z(N22) );
  MUX2_X1 U628 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n614), .Z(n34) );
  MUX2_X1 U629 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n619), .Z(n35) );
  MUX2_X1 U630 ( .A(n35), .B(n34), .S(n612), .Z(n36) );
  MUX2_X1 U631 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n614), .Z(n37) );
  MUX2_X1 U632 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n615), .Z(n38) );
  MUX2_X1 U633 ( .A(n38), .B(n37), .S(N11), .Z(n39) );
  MUX2_X1 U634 ( .A(n39), .B(n36), .S(n609), .Z(n40) );
  MUX2_X1 U635 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n615), .Z(n41) );
  MUX2_X1 U636 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n619), .Z(n42) );
  MUX2_X1 U637 ( .A(n42), .B(n41), .S(n611), .Z(n43) );
  MUX2_X1 U638 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n617), .Z(n44) );
  MUX2_X1 U639 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n618), .Z(n45) );
  MUX2_X1 U640 ( .A(n45), .B(n44), .S(N11), .Z(n46) );
  MUX2_X1 U641 ( .A(n46), .B(n43), .S(n609), .Z(n47) );
  MUX2_X1 U642 ( .A(n47), .B(n40), .S(N13), .Z(n48) );
  MUX2_X1 U643 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n619), .Z(n49) );
  MUX2_X1 U644 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n616), .Z(n50) );
  MUX2_X1 U645 ( .A(n50), .B(n49), .S(n611), .Z(n51) );
  MUX2_X1 U646 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n619), .Z(n52) );
  MUX2_X1 U647 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n619), .Z(n53) );
  MUX2_X1 U648 ( .A(n53), .B(n52), .S(n612), .Z(n54) );
  MUX2_X1 U649 ( .A(n54), .B(n51), .S(n609), .Z(n55) );
  MUX2_X1 U650 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n619), .Z(n56) );
  MUX2_X1 U651 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n57) );
  MUX2_X1 U652 ( .A(n57), .B(n56), .S(n613), .Z(n58) );
  MUX2_X1 U653 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n618), .Z(n59) );
  MUX2_X1 U654 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n619), .Z(n60) );
  MUX2_X1 U655 ( .A(n60), .B(n59), .S(n612), .Z(n61) );
  MUX2_X1 U656 ( .A(n61), .B(n58), .S(n609), .Z(n62) );
  MUX2_X1 U657 ( .A(n62), .B(n55), .S(N13), .Z(n63) );
  MUX2_X1 U658 ( .A(n63), .B(n48), .S(N14), .Z(N21) );
  MUX2_X1 U659 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n615), .Z(n64) );
  MUX2_X1 U660 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n615), .Z(n65) );
  MUX2_X1 U661 ( .A(n65), .B(n64), .S(n611), .Z(n66) );
  MUX2_X1 U662 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n615), .Z(n67) );
  MUX2_X1 U663 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n615), .Z(n68) );
  MUX2_X1 U664 ( .A(n68), .B(n67), .S(n611), .Z(n69) );
  MUX2_X1 U665 ( .A(n69), .B(n66), .S(n609), .Z(n70) );
  MUX2_X1 U666 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n615), .Z(n71) );
  MUX2_X1 U667 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n615), .Z(n72) );
  MUX2_X1 U668 ( .A(n72), .B(n71), .S(n611), .Z(n73) );
  MUX2_X1 U669 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n615), .Z(n74) );
  MUX2_X1 U670 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n615), .Z(n75) );
  MUX2_X1 U671 ( .A(n75), .B(n74), .S(n611), .Z(n76) );
  MUX2_X1 U672 ( .A(n76), .B(n73), .S(n610), .Z(n77) );
  MUX2_X1 U673 ( .A(n77), .B(n70), .S(N13), .Z(n78) );
  MUX2_X1 U674 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n615), .Z(n79) );
  MUX2_X1 U675 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n615), .Z(n80) );
  MUX2_X1 U676 ( .A(n80), .B(n79), .S(n611), .Z(n81) );
  MUX2_X1 U677 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n615), .Z(n82) );
  MUX2_X1 U678 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n615), .Z(n83) );
  MUX2_X1 U679 ( .A(n83), .B(n82), .S(n613), .Z(n84) );
  MUX2_X1 U680 ( .A(n84), .B(n81), .S(n609), .Z(n85) );
  MUX2_X1 U681 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n616), .Z(n86) );
  MUX2_X1 U682 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n616), .Z(n87) );
  MUX2_X1 U683 ( .A(n87), .B(n86), .S(n612), .Z(n88) );
  MUX2_X1 U684 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n616), .Z(n89) );
  MUX2_X1 U685 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n616), .Z(n90) );
  MUX2_X1 U686 ( .A(n90), .B(n89), .S(n611), .Z(n91) );
  MUX2_X1 U687 ( .A(n91), .B(n88), .S(n609), .Z(n92) );
  MUX2_X1 U688 ( .A(n92), .B(n85), .S(N13), .Z(n93) );
  MUX2_X1 U689 ( .A(n93), .B(n78), .S(N14), .Z(N20) );
  MUX2_X1 U690 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n616), .Z(n94) );
  MUX2_X1 U691 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n616), .Z(n95) );
  MUX2_X1 U692 ( .A(n95), .B(n94), .S(n611), .Z(n96) );
  MUX2_X1 U693 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n616), .Z(n97) );
  MUX2_X1 U694 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n616), .Z(n98) );
  MUX2_X1 U695 ( .A(n98), .B(n97), .S(n611), .Z(n99) );
  MUX2_X1 U696 ( .A(n99), .B(n96), .S(n609), .Z(n100) );
  MUX2_X1 U697 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n616), .Z(n101) );
  MUX2_X1 U698 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n616), .Z(n102) );
  MUX2_X1 U699 ( .A(n102), .B(n101), .S(n611), .Z(n103) );
  MUX2_X1 U700 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n616), .Z(n104) );
  MUX2_X1 U701 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n616), .Z(n105) );
  MUX2_X1 U702 ( .A(n105), .B(n104), .S(N11), .Z(n106) );
  MUX2_X1 U703 ( .A(n106), .B(n103), .S(n609), .Z(n107) );
  MUX2_X1 U704 ( .A(n107), .B(n100), .S(N13), .Z(n108) );
  MUX2_X1 U705 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n619), .Z(n109) );
  MUX2_X1 U706 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n619), .Z(n110) );
  MUX2_X1 U707 ( .A(n110), .B(n109), .S(n612), .Z(n111) );
  MUX2_X1 U708 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n619), .Z(n112) );
  MUX2_X1 U709 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n619), .Z(n113) );
  MUX2_X1 U710 ( .A(n113), .B(n112), .S(n612), .Z(n114) );
  MUX2_X1 U711 ( .A(n114), .B(n111), .S(n610), .Z(n115) );
  MUX2_X1 U712 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n619), .Z(n116) );
  MUX2_X1 U713 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n619), .Z(n117) );
  MUX2_X1 U714 ( .A(n117), .B(n116), .S(n612), .Z(n118) );
  MUX2_X1 U715 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n619), .Z(n119) );
  MUX2_X1 U716 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n617), .Z(n120) );
  MUX2_X1 U717 ( .A(n120), .B(n119), .S(n612), .Z(n121) );
  MUX2_X1 U718 ( .A(n121), .B(n118), .S(n610), .Z(n122) );
  MUX2_X1 U719 ( .A(n122), .B(n115), .S(N13), .Z(n123) );
  MUX2_X1 U720 ( .A(n123), .B(n108), .S(N14), .Z(N19) );
  MUX2_X1 U721 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n616), .Z(n124) );
  MUX2_X1 U722 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n619), .Z(n125) );
  MUX2_X1 U723 ( .A(n125), .B(n124), .S(n612), .Z(n126) );
  MUX2_X1 U724 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n619), .Z(n127) );
  MUX2_X1 U725 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n619), .Z(n128) );
  MUX2_X1 U726 ( .A(n128), .B(n127), .S(n612), .Z(n129) );
  MUX2_X1 U727 ( .A(n129), .B(n126), .S(n609), .Z(n130) );
  MUX2_X1 U728 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n615), .Z(n131) );
  MUX2_X1 U729 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n614), .Z(n132) );
  MUX2_X1 U730 ( .A(n132), .B(n131), .S(n612), .Z(n133) );
  MUX2_X1 U731 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n615), .Z(n134) );
  MUX2_X1 U732 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n618), .Z(n135) );
  MUX2_X1 U733 ( .A(n135), .B(n134), .S(n612), .Z(n136) );
  MUX2_X1 U734 ( .A(n136), .B(n133), .S(n610), .Z(n137) );
  MUX2_X1 U735 ( .A(n137), .B(n130), .S(N13), .Z(n138) );
  MUX2_X1 U736 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n614), .Z(n139) );
  MUX2_X1 U737 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n614), .Z(n140) );
  MUX2_X1 U738 ( .A(n140), .B(n139), .S(n612), .Z(n141) );
  MUX2_X1 U739 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n614), .Z(n142) );
  MUX2_X1 U740 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n617), .Z(n143) );
  MUX2_X1 U741 ( .A(n143), .B(n142), .S(n612), .Z(n144) );
  MUX2_X1 U742 ( .A(n144), .B(n141), .S(n609), .Z(n145) );
  MUX2_X1 U743 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n614), .Z(n146) );
  MUX2_X1 U744 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n619), .Z(n147) );
  MUX2_X1 U745 ( .A(n147), .B(n146), .S(n612), .Z(n148) );
  MUX2_X1 U746 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n619), .Z(n149) );
  MUX2_X1 U747 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n619), .Z(n150) );
  MUX2_X1 U748 ( .A(n150), .B(n149), .S(n612), .Z(n151) );
  MUX2_X1 U749 ( .A(n151), .B(n148), .S(n609), .Z(n152) );
  MUX2_X1 U750 ( .A(n152), .B(n145), .S(N13), .Z(n153) );
  MUX2_X1 U751 ( .A(n153), .B(n138), .S(N14), .Z(N18) );
  MUX2_X1 U752 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n615), .Z(n154) );
  MUX2_X1 U753 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n614), .Z(n155) );
  MUX2_X1 U754 ( .A(n155), .B(n154), .S(n613), .Z(n156) );
  MUX2_X1 U755 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n615), .Z(n157) );
  MUX2_X1 U756 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n614), .Z(n158) );
  MUX2_X1 U757 ( .A(n158), .B(n157), .S(n613), .Z(n159) );
  MUX2_X1 U758 ( .A(n159), .B(n156), .S(n610), .Z(n160) );
  MUX2_X1 U759 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n615), .Z(n161) );
  MUX2_X1 U760 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n614), .Z(n162) );
  MUX2_X1 U761 ( .A(n162), .B(n161), .S(n613), .Z(n163) );
  MUX2_X1 U762 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n615), .Z(n164) );
  MUX2_X1 U763 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n614), .Z(n165) );
  MUX2_X1 U764 ( .A(n165), .B(n164), .S(n613), .Z(n166) );
  MUX2_X1 U765 ( .A(n166), .B(n163), .S(n610), .Z(n167) );
  MUX2_X1 U766 ( .A(n167), .B(n160), .S(N13), .Z(n168) );
  MUX2_X1 U767 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n614), .Z(n169) );
  MUX2_X1 U768 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n615), .Z(n170) );
  MUX2_X1 U769 ( .A(n170), .B(n169), .S(n613), .Z(n171) );
  MUX2_X1 U770 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n614), .Z(n172) );
  MUX2_X1 U771 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n615), .Z(n173) );
  MUX2_X1 U772 ( .A(n173), .B(n172), .S(n613), .Z(n174) );
  MUX2_X1 U773 ( .A(n174), .B(n171), .S(n610), .Z(n175) );
  MUX2_X1 U774 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n617), .Z(n176) );
  MUX2_X1 U775 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n617), .Z(n177) );
  MUX2_X1 U776 ( .A(n177), .B(n176), .S(n613), .Z(n178) );
  MUX2_X1 U777 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n617), .Z(n179) );
  MUX2_X1 U778 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n617), .Z(n180) );
  MUX2_X1 U779 ( .A(n180), .B(n179), .S(n613), .Z(n181) );
  MUX2_X1 U780 ( .A(n181), .B(n178), .S(n610), .Z(n182) );
  MUX2_X1 U781 ( .A(n182), .B(n175), .S(N13), .Z(n183) );
  MUX2_X1 U782 ( .A(n183), .B(n168), .S(N14), .Z(N17) );
  MUX2_X1 U783 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n617), .Z(n184) );
  MUX2_X1 U784 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n617), .Z(n185) );
  MUX2_X1 U785 ( .A(n185), .B(n184), .S(n613), .Z(n186) );
  MUX2_X1 U786 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n617), .Z(n187) );
  MUX2_X1 U787 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n617), .Z(n188) );
  MUX2_X1 U788 ( .A(n188), .B(n187), .S(n613), .Z(n189) );
  MUX2_X1 U789 ( .A(n189), .B(n186), .S(n610), .Z(n190) );
  MUX2_X1 U790 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n617), .Z(n191) );
  MUX2_X1 U791 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n617), .Z(n192) );
  MUX2_X1 U792 ( .A(n192), .B(n191), .S(n613), .Z(n193) );
  MUX2_X1 U793 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n617), .Z(n194) );
  MUX2_X1 U794 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n617), .Z(n195) );
  MUX2_X1 U795 ( .A(n195), .B(n194), .S(n613), .Z(n196) );
  MUX2_X1 U796 ( .A(n196), .B(n193), .S(n610), .Z(n197) );
  MUX2_X1 U797 ( .A(n197), .B(n190), .S(N13), .Z(n198) );
  MUX2_X1 U798 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n618), .Z(n199) );
  MUX2_X1 U799 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n618), .Z(n200) );
  MUX2_X1 U800 ( .A(n200), .B(n199), .S(n613), .Z(n201) );
  MUX2_X1 U801 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n618), .Z(n202) );
  MUX2_X1 U802 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n618), .Z(n203) );
  MUX2_X1 U803 ( .A(n203), .B(n202), .S(n613), .Z(n204) );
  MUX2_X1 U804 ( .A(n204), .B(n201), .S(n610), .Z(n205) );
  MUX2_X1 U805 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n618), .Z(n206) );
  MUX2_X1 U806 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n618), .Z(n207) );
  MUX2_X1 U807 ( .A(n207), .B(n206), .S(n613), .Z(n208) );
  MUX2_X1 U808 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n618), .Z(n209) );
  MUX2_X1 U809 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n618), .Z(n210) );
  MUX2_X1 U810 ( .A(n210), .B(n209), .S(n611), .Z(n211) );
  MUX2_X1 U811 ( .A(n211), .B(n208), .S(n610), .Z(n212) );
  MUX2_X1 U812 ( .A(n212), .B(n205), .S(N13), .Z(n213) );
  MUX2_X1 U813 ( .A(n213), .B(n198), .S(N14), .Z(N16) );
  MUX2_X1 U814 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n618), .Z(n214) );
  MUX2_X1 U815 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n618), .Z(n215) );
  MUX2_X1 U816 ( .A(n215), .B(n214), .S(n612), .Z(n216) );
  MUX2_X1 U817 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n618), .Z(n217) );
  MUX2_X1 U818 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n618), .Z(n218) );
  MUX2_X1 U819 ( .A(n218), .B(n217), .S(N11), .Z(n219) );
  MUX2_X1 U820 ( .A(n219), .B(n216), .S(n610), .Z(n220) );
  MUX2_X1 U821 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n616), .Z(n221) );
  MUX2_X1 U822 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n618), .Z(n222) );
  MUX2_X1 U823 ( .A(n222), .B(n221), .S(n611), .Z(n223) );
  MUX2_X1 U824 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n618), .Z(n224) );
  MUX2_X1 U825 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n617), .Z(n225) );
  MUX2_X1 U826 ( .A(n225), .B(n224), .S(n613), .Z(n226) );
  MUX2_X1 U827 ( .A(n226), .B(n223), .S(n610), .Z(n227) );
  MUX2_X1 U828 ( .A(n227), .B(n220), .S(N13), .Z(n228) );
  MUX2_X1 U829 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n617), .Z(n229) );
  MUX2_X1 U830 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n618), .Z(n595) );
  MUX2_X1 U831 ( .A(n595), .B(n229), .S(n612), .Z(n596) );
  MUX2_X1 U832 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n616), .Z(n597) );
  MUX2_X1 U833 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n616), .Z(n598) );
  MUX2_X1 U834 ( .A(n598), .B(n597), .S(n612), .Z(n599) );
  MUX2_X1 U835 ( .A(n599), .B(n596), .S(n610), .Z(n600) );
  MUX2_X1 U836 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n617), .Z(n601) );
  MUX2_X1 U837 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n617), .Z(n602) );
  MUX2_X1 U838 ( .A(n602), .B(n601), .S(n612), .Z(n603) );
  MUX2_X1 U839 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n616), .Z(n604) );
  MUX2_X1 U840 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n618), .Z(n605) );
  MUX2_X1 U841 ( .A(n605), .B(n604), .S(n613), .Z(n606) );
  MUX2_X1 U842 ( .A(n606), .B(n603), .S(n610), .Z(n607) );
  MUX2_X1 U843 ( .A(n607), .B(n600), .S(N13), .Z(n608) );
  MUX2_X1 U844 ( .A(n608), .B(n228), .S(N14), .Z(N15) );
  CLKBUF_X1 U845 ( .A(N11), .Z(n611) );
  CLKBUF_X1 U846 ( .A(N10), .Z(n614) );
  INV_X1 U847 ( .A(N10), .ZN(n620) );
  INV_X1 U848 ( .A(N11), .ZN(n621) );
  INV_X1 U849 ( .A(data_in[0]), .ZN(n622) );
  INV_X1 U850 ( .A(data_in[1]), .ZN(n623) );
  INV_X1 U851 ( .A(data_in[2]), .ZN(n624) );
  INV_X1 U852 ( .A(data_in[3]), .ZN(n625) );
  INV_X1 U853 ( .A(data_in[4]), .ZN(n626) );
  INV_X1 U854 ( .A(data_in[5]), .ZN(n627) );
  INV_X1 U855 ( .A(data_in[6]), .ZN(n628) );
  INV_X1 U856 ( .A(data_in[7]), .ZN(n629) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6_0 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, n2,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .QN(n2) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n630), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n631), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n632), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n633), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n634), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n635), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n636), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n637), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n638), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n639), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n640), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n641), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n642), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n643), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n644), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n645), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n646), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n647), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n648), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n649), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n650), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n651), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n652), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n653), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n654), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n655), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n656), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n657), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n658), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n659), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n660), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n661), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n662), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n663), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n664), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n665), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n666), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n667), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n668), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n669), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n670), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n671), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n672), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n673), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n674), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n675), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n676), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n677), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n678), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n679), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n680), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n681), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n682), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n683), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n684), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n685), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n686), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n687), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n688), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n689), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n690), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n691), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n692), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n693), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n694), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n695), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n696), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n697), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n698), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n699), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n700), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n701), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n702), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n703), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n704), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n705), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n706), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n707), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n708), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n709), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n710), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n711), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n712), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n713), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n714), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n715), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n716), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n717), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n718), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n719), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n720), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n721), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n722), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n723), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n724), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n725), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n726), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n727), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n728), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n729), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n730), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n731), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n732), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n733), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n734), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n735), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n736), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n737), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n738), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n739), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n740), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n741), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n742), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n743), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n744), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n745), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n746), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n747), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n748), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n749), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n750), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n751), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n752), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n753), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n754), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n755), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n756), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n757), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n758), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n759), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n760), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n761), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n762), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n763), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n764), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n765), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n766), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n767), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n768), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n769), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n770), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n771), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n772), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n773), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n774), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n775), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n776), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n777), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n778), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n779), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n780), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n781), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n782), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n783), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n784), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n785), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n786), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n787), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n788), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n789), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n790), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n791), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n792), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n793), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n794), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n795), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n796), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n797), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n798), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n799), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n800), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n801), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n802), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n803), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n804), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n805), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n806), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n807), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n808), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n809), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n810), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n811), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n812), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n813), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n814), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n815), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n816), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n817), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n818), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n819), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n820), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n821), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n849), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n850), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n851), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n852), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n853), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n854), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n855), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n856), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n857), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n858), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n859), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n860), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n861), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n862), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n863), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n864), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n865), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n866), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n867), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n868), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n869), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n870), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n871), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n872), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n873), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n874), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n875), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n876), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n877), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n878), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n879), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n880), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n881), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n882), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n883), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n884), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n885), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n886), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n887), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n888), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n889), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n890), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n891), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n892), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n893), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n894), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n895), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n896), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n897), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n898), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n899), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n900), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n901), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n902), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n903), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n904), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n905), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n906), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n907), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n908), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n909), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n910), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n911), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n912), .CK(clk), .Q(\mem[0][0] ) );
  SDFF_X1 \data_out_reg[1]  ( .D(n48), .SI(n63), .SE(n847), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n18), .SI(n33), .SE(n847), .CK(clk), .Q(
        data_out[0]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n93), .SI(n78), .SE(N14), .CK(clk), .Q(
        data_out[2]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  BUF_X1 U3 ( .A(N10), .Z(n614) );
  INV_X2 U4 ( .A(n2), .ZN(data_out[4]) );
  BUF_X1 U5 ( .A(n619), .Z(n617) );
  BUF_X1 U6 ( .A(n619), .Z(n618) );
  BUF_X1 U7 ( .A(n619), .Z(n615) );
  BUF_X1 U8 ( .A(N10), .Z(n616) );
  BUF_X1 U9 ( .A(N11), .Z(n611) );
  BUF_X1 U10 ( .A(N11), .Z(n612) );
  BUF_X1 U11 ( .A(N11), .Z(n613) );
  BUF_X1 U12 ( .A(N10), .Z(n619) );
  INV_X1 U13 ( .A(n1130), .ZN(n845) );
  INV_X1 U14 ( .A(n1120), .ZN(n824) );
  INV_X1 U15 ( .A(n1111), .ZN(n842) );
  INV_X1 U16 ( .A(n1102), .ZN(n827) );
  INV_X1 U17 ( .A(n1057), .ZN(n844) );
  INV_X1 U18 ( .A(n1047), .ZN(n823) );
  INV_X1 U19 ( .A(n1038), .ZN(n841) );
  INV_X1 U20 ( .A(n1029), .ZN(n826) );
  INV_X1 U21 ( .A(n984), .ZN(n843) );
  INV_X1 U22 ( .A(n974), .ZN(n822) );
  INV_X1 U23 ( .A(n965), .ZN(n840) );
  INV_X1 U24 ( .A(n956), .ZN(n825) );
  INV_X1 U25 ( .A(n1093), .ZN(n830) );
  INV_X1 U26 ( .A(n1084), .ZN(n839) );
  INV_X1 U27 ( .A(n1075), .ZN(n833) );
  INV_X1 U28 ( .A(n1066), .ZN(n836) );
  INV_X1 U29 ( .A(n947), .ZN(n828) );
  INV_X1 U30 ( .A(n938), .ZN(n837) );
  INV_X1 U31 ( .A(n929), .ZN(n831) );
  INV_X1 U32 ( .A(n920), .ZN(n834) );
  INV_X1 U33 ( .A(n1020), .ZN(n829) );
  INV_X1 U34 ( .A(n1011), .ZN(n838) );
  INV_X1 U35 ( .A(n1002), .ZN(n832) );
  INV_X1 U36 ( .A(n993), .ZN(n835) );
  NAND2_X1 U37 ( .A1(n1193), .A2(n1203), .ZN(n1202) );
  NAND2_X1 U38 ( .A1(n1183), .A2(n1203), .ZN(n1192) );
  NAND2_X1 U39 ( .A1(n1173), .A2(n1203), .ZN(n1182) );
  NAND2_X1 U40 ( .A1(n1163), .A2(n1203), .ZN(n1172) );
  NAND2_X1 U41 ( .A1(n1153), .A2(n1203), .ZN(n1162) );
  NAND2_X1 U42 ( .A1(n1143), .A2(n1203), .ZN(n1152) );
  NAND2_X1 U43 ( .A1(n1133), .A2(n1203), .ZN(n1142) );
  NAND2_X1 U44 ( .A1(n1204), .A2(n1203), .ZN(n1213) );
  NOR3_X1 U45 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1204) );
  NOR3_X1 U46 ( .A1(N11), .A2(N12), .A3(n620), .ZN(n1193) );
  NOR3_X1 U47 ( .A1(N10), .A2(N12), .A3(n621), .ZN(n1183) );
  NOR3_X1 U48 ( .A1(n620), .A2(N12), .A3(n621), .ZN(n1173) );
  NAND2_X1 U49 ( .A1(n1122), .A2(n1204), .ZN(n1130) );
  NAND2_X1 U50 ( .A1(n1122), .A2(n1193), .ZN(n1120) );
  NAND2_X1 U51 ( .A1(n1122), .A2(n1183), .ZN(n1111) );
  NAND2_X1 U52 ( .A1(n1122), .A2(n1173), .ZN(n1102) );
  NAND2_X1 U53 ( .A1(n1049), .A2(n1204), .ZN(n1057) );
  NAND2_X1 U54 ( .A1(n1049), .A2(n1193), .ZN(n1047) );
  NAND2_X1 U55 ( .A1(n1049), .A2(n1183), .ZN(n1038) );
  NAND2_X1 U56 ( .A1(n1049), .A2(n1173), .ZN(n1029) );
  NAND2_X1 U57 ( .A1(n976), .A2(n1204), .ZN(n984) );
  NAND2_X1 U58 ( .A1(n976), .A2(n1193), .ZN(n974) );
  NAND2_X1 U59 ( .A1(n976), .A2(n1183), .ZN(n965) );
  NAND2_X1 U60 ( .A1(n976), .A2(n1173), .ZN(n956) );
  NAND2_X1 U61 ( .A1(n1122), .A2(n1163), .ZN(n1093) );
  NAND2_X1 U62 ( .A1(n1122), .A2(n1153), .ZN(n1084) );
  NAND2_X1 U63 ( .A1(n1122), .A2(n1143), .ZN(n1075) );
  NAND2_X1 U64 ( .A1(n1122), .A2(n1133), .ZN(n1066) );
  NAND2_X1 U65 ( .A1(n1049), .A2(n1163), .ZN(n1020) );
  NAND2_X1 U66 ( .A1(n1049), .A2(n1153), .ZN(n1011) );
  NAND2_X1 U67 ( .A1(n1049), .A2(n1143), .ZN(n1002) );
  NAND2_X1 U68 ( .A1(n1049), .A2(n1133), .ZN(n993) );
  NAND2_X1 U69 ( .A1(n976), .A2(n1163), .ZN(n947) );
  NAND2_X1 U70 ( .A1(n976), .A2(n1153), .ZN(n938) );
  NAND2_X1 U71 ( .A1(n976), .A2(n1143), .ZN(n929) );
  NAND2_X1 U72 ( .A1(n976), .A2(n1133), .ZN(n920) );
  BUF_X1 U73 ( .A(N12), .Z(n610) );
  INV_X1 U74 ( .A(N13), .ZN(n846) );
  AND3_X1 U75 ( .A1(n620), .A2(n621), .A3(N12), .ZN(n1163) );
  AND3_X1 U76 ( .A1(N10), .A2(n621), .A3(N12), .ZN(n1153) );
  AND3_X1 U77 ( .A1(N11), .A2(n620), .A3(N12), .ZN(n1143) );
  AND3_X1 U78 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n1133) );
  BUF_X1 U79 ( .A(N12), .Z(n609) );
  INV_X1 U80 ( .A(N14), .ZN(n847) );
  AND3_X1 U81 ( .A1(n846), .A2(n847), .A3(n1132), .ZN(n1203) );
  AND3_X1 U82 ( .A1(N13), .A2(n1132), .A3(N14), .ZN(n976) );
  AND3_X1 U83 ( .A1(n1132), .A2(n847), .A3(N13), .ZN(n1122) );
  AND3_X1 U84 ( .A1(n1132), .A2(n846), .A3(N14), .ZN(n1049) );
  NOR2_X1 U85 ( .A1(n848), .A2(addr[5]), .ZN(n1132) );
  INV_X1 U86 ( .A(wr_en), .ZN(n848) );
  OAI21_X1 U87 ( .B1(n622), .B2(n1172), .A(n1171), .ZN(n880) );
  NAND2_X1 U88 ( .A1(\mem[4][0] ), .A2(n1172), .ZN(n1171) );
  OAI21_X1 U89 ( .B1(n623), .B2(n1172), .A(n1170), .ZN(n879) );
  NAND2_X1 U90 ( .A1(\mem[4][1] ), .A2(n1172), .ZN(n1170) );
  OAI21_X1 U91 ( .B1(n624), .B2(n1172), .A(n1169), .ZN(n878) );
  NAND2_X1 U92 ( .A1(\mem[4][2] ), .A2(n1172), .ZN(n1169) );
  OAI21_X1 U93 ( .B1(n625), .B2(n1172), .A(n1168), .ZN(n877) );
  NAND2_X1 U94 ( .A1(\mem[4][3] ), .A2(n1172), .ZN(n1168) );
  OAI21_X1 U95 ( .B1(n626), .B2(n1172), .A(n1167), .ZN(n876) );
  NAND2_X1 U96 ( .A1(\mem[4][4] ), .A2(n1172), .ZN(n1167) );
  OAI21_X1 U97 ( .B1(n627), .B2(n1172), .A(n1166), .ZN(n875) );
  NAND2_X1 U98 ( .A1(\mem[4][5] ), .A2(n1172), .ZN(n1166) );
  OAI21_X1 U99 ( .B1(n628), .B2(n1172), .A(n1165), .ZN(n874) );
  NAND2_X1 U100 ( .A1(\mem[4][6] ), .A2(n1172), .ZN(n1165) );
  OAI21_X1 U101 ( .B1(n629), .B2(n1172), .A(n1164), .ZN(n873) );
  NAND2_X1 U102 ( .A1(\mem[4][7] ), .A2(n1172), .ZN(n1164) );
  OAI21_X1 U103 ( .B1(n622), .B2(n1152), .A(n1151), .ZN(n864) );
  NAND2_X1 U104 ( .A1(\mem[6][0] ), .A2(n1152), .ZN(n1151) );
  OAI21_X1 U105 ( .B1(n623), .B2(n1152), .A(n1150), .ZN(n863) );
  NAND2_X1 U106 ( .A1(\mem[6][1] ), .A2(n1152), .ZN(n1150) );
  OAI21_X1 U107 ( .B1(n624), .B2(n1152), .A(n1149), .ZN(n862) );
  NAND2_X1 U108 ( .A1(\mem[6][2] ), .A2(n1152), .ZN(n1149) );
  OAI21_X1 U109 ( .B1(n625), .B2(n1152), .A(n1148), .ZN(n861) );
  NAND2_X1 U110 ( .A1(\mem[6][3] ), .A2(n1152), .ZN(n1148) );
  OAI21_X1 U111 ( .B1(n626), .B2(n1152), .A(n1147), .ZN(n860) );
  NAND2_X1 U112 ( .A1(\mem[6][4] ), .A2(n1152), .ZN(n1147) );
  OAI21_X1 U113 ( .B1(n627), .B2(n1152), .A(n1146), .ZN(n859) );
  NAND2_X1 U114 ( .A1(\mem[6][5] ), .A2(n1152), .ZN(n1146) );
  OAI21_X1 U115 ( .B1(n628), .B2(n1152), .A(n1145), .ZN(n858) );
  NAND2_X1 U116 ( .A1(\mem[6][6] ), .A2(n1152), .ZN(n1145) );
  OAI21_X1 U117 ( .B1(n629), .B2(n1152), .A(n1144), .ZN(n857) );
  NAND2_X1 U118 ( .A1(\mem[6][7] ), .A2(n1152), .ZN(n1144) );
  OAI21_X1 U119 ( .B1(n622), .B2(n1142), .A(n1141), .ZN(n856) );
  NAND2_X1 U120 ( .A1(\mem[7][0] ), .A2(n1142), .ZN(n1141) );
  OAI21_X1 U121 ( .B1(n623), .B2(n1142), .A(n1140), .ZN(n855) );
  NAND2_X1 U122 ( .A1(\mem[7][1] ), .A2(n1142), .ZN(n1140) );
  OAI21_X1 U123 ( .B1(n624), .B2(n1142), .A(n1139), .ZN(n854) );
  NAND2_X1 U124 ( .A1(\mem[7][2] ), .A2(n1142), .ZN(n1139) );
  OAI21_X1 U125 ( .B1(n625), .B2(n1142), .A(n1138), .ZN(n853) );
  NAND2_X1 U126 ( .A1(\mem[7][3] ), .A2(n1142), .ZN(n1138) );
  OAI21_X1 U127 ( .B1(n626), .B2(n1142), .A(n1137), .ZN(n852) );
  NAND2_X1 U128 ( .A1(\mem[7][4] ), .A2(n1142), .ZN(n1137) );
  OAI21_X1 U129 ( .B1(n627), .B2(n1142), .A(n1136), .ZN(n851) );
  NAND2_X1 U130 ( .A1(\mem[7][5] ), .A2(n1142), .ZN(n1136) );
  OAI21_X1 U131 ( .B1(n628), .B2(n1142), .A(n1135), .ZN(n850) );
  NAND2_X1 U132 ( .A1(\mem[7][6] ), .A2(n1142), .ZN(n1135) );
  OAI21_X1 U133 ( .B1(n629), .B2(n1142), .A(n1134), .ZN(n849) );
  NAND2_X1 U134 ( .A1(\mem[7][7] ), .A2(n1142), .ZN(n1134) );
  OAI21_X1 U135 ( .B1(n622), .B2(n1202), .A(n1201), .ZN(n904) );
  NAND2_X1 U136 ( .A1(\mem[1][0] ), .A2(n1202), .ZN(n1201) );
  OAI21_X1 U137 ( .B1(n623), .B2(n1202), .A(n1200), .ZN(n903) );
  NAND2_X1 U138 ( .A1(\mem[1][1] ), .A2(n1202), .ZN(n1200) );
  OAI21_X1 U139 ( .B1(n624), .B2(n1202), .A(n1199), .ZN(n902) );
  NAND2_X1 U140 ( .A1(\mem[1][2] ), .A2(n1202), .ZN(n1199) );
  OAI21_X1 U141 ( .B1(n625), .B2(n1202), .A(n1198), .ZN(n901) );
  NAND2_X1 U142 ( .A1(\mem[1][3] ), .A2(n1202), .ZN(n1198) );
  OAI21_X1 U143 ( .B1(n626), .B2(n1202), .A(n1197), .ZN(n900) );
  NAND2_X1 U144 ( .A1(\mem[1][4] ), .A2(n1202), .ZN(n1197) );
  OAI21_X1 U145 ( .B1(n627), .B2(n1202), .A(n1196), .ZN(n899) );
  NAND2_X1 U146 ( .A1(\mem[1][5] ), .A2(n1202), .ZN(n1196) );
  OAI21_X1 U147 ( .B1(n628), .B2(n1202), .A(n1195), .ZN(n898) );
  NAND2_X1 U148 ( .A1(\mem[1][6] ), .A2(n1202), .ZN(n1195) );
  OAI21_X1 U149 ( .B1(n629), .B2(n1202), .A(n1194), .ZN(n897) );
  NAND2_X1 U150 ( .A1(\mem[1][7] ), .A2(n1202), .ZN(n1194) );
  OAI21_X1 U151 ( .B1(n622), .B2(n1192), .A(n1191), .ZN(n896) );
  NAND2_X1 U152 ( .A1(\mem[2][0] ), .A2(n1192), .ZN(n1191) );
  OAI21_X1 U153 ( .B1(n623), .B2(n1192), .A(n1190), .ZN(n895) );
  NAND2_X1 U154 ( .A1(\mem[2][1] ), .A2(n1192), .ZN(n1190) );
  OAI21_X1 U155 ( .B1(n624), .B2(n1192), .A(n1189), .ZN(n894) );
  NAND2_X1 U156 ( .A1(\mem[2][2] ), .A2(n1192), .ZN(n1189) );
  OAI21_X1 U157 ( .B1(n625), .B2(n1192), .A(n1188), .ZN(n893) );
  NAND2_X1 U158 ( .A1(\mem[2][3] ), .A2(n1192), .ZN(n1188) );
  OAI21_X1 U159 ( .B1(n626), .B2(n1192), .A(n1187), .ZN(n892) );
  NAND2_X1 U160 ( .A1(\mem[2][4] ), .A2(n1192), .ZN(n1187) );
  OAI21_X1 U161 ( .B1(n627), .B2(n1192), .A(n1186), .ZN(n891) );
  NAND2_X1 U162 ( .A1(\mem[2][5] ), .A2(n1192), .ZN(n1186) );
  OAI21_X1 U163 ( .B1(n628), .B2(n1192), .A(n1185), .ZN(n890) );
  NAND2_X1 U164 ( .A1(\mem[2][6] ), .A2(n1192), .ZN(n1185) );
  OAI21_X1 U165 ( .B1(n629), .B2(n1192), .A(n1184), .ZN(n889) );
  NAND2_X1 U166 ( .A1(\mem[2][7] ), .A2(n1192), .ZN(n1184) );
  OAI21_X1 U167 ( .B1(n622), .B2(n1182), .A(n1181), .ZN(n888) );
  NAND2_X1 U168 ( .A1(\mem[3][0] ), .A2(n1182), .ZN(n1181) );
  OAI21_X1 U169 ( .B1(n623), .B2(n1182), .A(n1180), .ZN(n887) );
  NAND2_X1 U170 ( .A1(\mem[3][1] ), .A2(n1182), .ZN(n1180) );
  OAI21_X1 U171 ( .B1(n624), .B2(n1182), .A(n1179), .ZN(n886) );
  NAND2_X1 U172 ( .A1(\mem[3][2] ), .A2(n1182), .ZN(n1179) );
  OAI21_X1 U173 ( .B1(n625), .B2(n1182), .A(n1178), .ZN(n885) );
  NAND2_X1 U174 ( .A1(\mem[3][3] ), .A2(n1182), .ZN(n1178) );
  OAI21_X1 U175 ( .B1(n626), .B2(n1182), .A(n1177), .ZN(n884) );
  NAND2_X1 U176 ( .A1(\mem[3][4] ), .A2(n1182), .ZN(n1177) );
  OAI21_X1 U177 ( .B1(n627), .B2(n1182), .A(n1176), .ZN(n883) );
  NAND2_X1 U178 ( .A1(\mem[3][5] ), .A2(n1182), .ZN(n1176) );
  OAI21_X1 U179 ( .B1(n628), .B2(n1182), .A(n1175), .ZN(n882) );
  NAND2_X1 U180 ( .A1(\mem[3][6] ), .A2(n1182), .ZN(n1175) );
  OAI21_X1 U181 ( .B1(n629), .B2(n1182), .A(n1174), .ZN(n881) );
  NAND2_X1 U182 ( .A1(\mem[3][7] ), .A2(n1182), .ZN(n1174) );
  OAI21_X1 U183 ( .B1(n622), .B2(n1162), .A(n1161), .ZN(n872) );
  NAND2_X1 U184 ( .A1(\mem[5][0] ), .A2(n1162), .ZN(n1161) );
  OAI21_X1 U185 ( .B1(n623), .B2(n1162), .A(n1160), .ZN(n871) );
  NAND2_X1 U186 ( .A1(\mem[5][1] ), .A2(n1162), .ZN(n1160) );
  OAI21_X1 U187 ( .B1(n624), .B2(n1162), .A(n1159), .ZN(n870) );
  NAND2_X1 U188 ( .A1(\mem[5][2] ), .A2(n1162), .ZN(n1159) );
  OAI21_X1 U189 ( .B1(n625), .B2(n1162), .A(n1158), .ZN(n869) );
  NAND2_X1 U190 ( .A1(\mem[5][3] ), .A2(n1162), .ZN(n1158) );
  OAI21_X1 U191 ( .B1(n626), .B2(n1162), .A(n1157), .ZN(n868) );
  NAND2_X1 U192 ( .A1(\mem[5][4] ), .A2(n1162), .ZN(n1157) );
  OAI21_X1 U193 ( .B1(n627), .B2(n1162), .A(n1156), .ZN(n867) );
  NAND2_X1 U194 ( .A1(\mem[5][5] ), .A2(n1162), .ZN(n1156) );
  OAI21_X1 U195 ( .B1(n628), .B2(n1162), .A(n1155), .ZN(n866) );
  NAND2_X1 U196 ( .A1(\mem[5][6] ), .A2(n1162), .ZN(n1155) );
  OAI21_X1 U197 ( .B1(n629), .B2(n1162), .A(n1154), .ZN(n865) );
  NAND2_X1 U198 ( .A1(\mem[5][7] ), .A2(n1162), .ZN(n1154) );
  OAI21_X1 U199 ( .B1(n1213), .B2(n622), .A(n1212), .ZN(n912) );
  NAND2_X1 U200 ( .A1(\mem[0][0] ), .A2(n1213), .ZN(n1212) );
  OAI21_X1 U201 ( .B1(n1213), .B2(n623), .A(n1211), .ZN(n911) );
  NAND2_X1 U202 ( .A1(\mem[0][1] ), .A2(n1213), .ZN(n1211) );
  OAI21_X1 U203 ( .B1(n1213), .B2(n624), .A(n1210), .ZN(n910) );
  NAND2_X1 U204 ( .A1(\mem[0][2] ), .A2(n1213), .ZN(n1210) );
  OAI21_X1 U205 ( .B1(n1213), .B2(n625), .A(n1209), .ZN(n909) );
  NAND2_X1 U206 ( .A1(\mem[0][3] ), .A2(n1213), .ZN(n1209) );
  OAI21_X1 U207 ( .B1(n1213), .B2(n626), .A(n1208), .ZN(n908) );
  NAND2_X1 U208 ( .A1(\mem[0][4] ), .A2(n1213), .ZN(n1208) );
  OAI21_X1 U209 ( .B1(n1213), .B2(n627), .A(n1207), .ZN(n907) );
  NAND2_X1 U210 ( .A1(\mem[0][5] ), .A2(n1213), .ZN(n1207) );
  OAI21_X1 U211 ( .B1(n1213), .B2(n628), .A(n1206), .ZN(n906) );
  NAND2_X1 U212 ( .A1(\mem[0][6] ), .A2(n1213), .ZN(n1206) );
  OAI21_X1 U213 ( .B1(n1213), .B2(n629), .A(n1205), .ZN(n905) );
  NAND2_X1 U214 ( .A1(\mem[0][7] ), .A2(n1213), .ZN(n1205) );
  INV_X1 U215 ( .A(n1131), .ZN(n821) );
  AOI22_X1 U216 ( .A1(data_in[0]), .A2(n845), .B1(n1130), .B2(\mem[8][0] ), 
        .ZN(n1131) );
  INV_X1 U217 ( .A(n1129), .ZN(n820) );
  AOI22_X1 U218 ( .A1(data_in[1]), .A2(n845), .B1(n1130), .B2(\mem[8][1] ), 
        .ZN(n1129) );
  INV_X1 U219 ( .A(n1128), .ZN(n819) );
  AOI22_X1 U220 ( .A1(data_in[2]), .A2(n845), .B1(n1130), .B2(\mem[8][2] ), 
        .ZN(n1128) );
  INV_X1 U221 ( .A(n1127), .ZN(n818) );
  AOI22_X1 U222 ( .A1(data_in[3]), .A2(n845), .B1(n1130), .B2(\mem[8][3] ), 
        .ZN(n1127) );
  INV_X1 U223 ( .A(n1126), .ZN(n817) );
  AOI22_X1 U224 ( .A1(data_in[4]), .A2(n845), .B1(n1130), .B2(\mem[8][4] ), 
        .ZN(n1126) );
  INV_X1 U225 ( .A(n1125), .ZN(n816) );
  AOI22_X1 U226 ( .A1(data_in[5]), .A2(n845), .B1(n1130), .B2(\mem[8][5] ), 
        .ZN(n1125) );
  INV_X1 U227 ( .A(n1124), .ZN(n815) );
  AOI22_X1 U228 ( .A1(data_in[6]), .A2(n845), .B1(n1130), .B2(\mem[8][6] ), 
        .ZN(n1124) );
  INV_X1 U229 ( .A(n1123), .ZN(n814) );
  AOI22_X1 U230 ( .A1(data_in[7]), .A2(n845), .B1(n1130), .B2(\mem[8][7] ), 
        .ZN(n1123) );
  INV_X1 U231 ( .A(n1121), .ZN(n813) );
  AOI22_X1 U232 ( .A1(data_in[0]), .A2(n824), .B1(n1120), .B2(\mem[9][0] ), 
        .ZN(n1121) );
  INV_X1 U233 ( .A(n1119), .ZN(n812) );
  AOI22_X1 U234 ( .A1(data_in[1]), .A2(n824), .B1(n1120), .B2(\mem[9][1] ), 
        .ZN(n1119) );
  INV_X1 U235 ( .A(n1118), .ZN(n811) );
  AOI22_X1 U236 ( .A1(data_in[2]), .A2(n824), .B1(n1120), .B2(\mem[9][2] ), 
        .ZN(n1118) );
  INV_X1 U237 ( .A(n1117), .ZN(n810) );
  AOI22_X1 U238 ( .A1(data_in[3]), .A2(n824), .B1(n1120), .B2(\mem[9][3] ), 
        .ZN(n1117) );
  INV_X1 U239 ( .A(n1116), .ZN(n809) );
  AOI22_X1 U240 ( .A1(data_in[4]), .A2(n824), .B1(n1120), .B2(\mem[9][4] ), 
        .ZN(n1116) );
  INV_X1 U241 ( .A(n1115), .ZN(n808) );
  AOI22_X1 U242 ( .A1(data_in[5]), .A2(n824), .B1(n1120), .B2(\mem[9][5] ), 
        .ZN(n1115) );
  INV_X1 U243 ( .A(n1114), .ZN(n807) );
  AOI22_X1 U244 ( .A1(data_in[6]), .A2(n824), .B1(n1120), .B2(\mem[9][6] ), 
        .ZN(n1114) );
  INV_X1 U245 ( .A(n1113), .ZN(n806) );
  AOI22_X1 U246 ( .A1(data_in[7]), .A2(n824), .B1(n1120), .B2(\mem[9][7] ), 
        .ZN(n1113) );
  INV_X1 U247 ( .A(n1112), .ZN(n805) );
  AOI22_X1 U248 ( .A1(data_in[0]), .A2(n842), .B1(n1111), .B2(\mem[10][0] ), 
        .ZN(n1112) );
  INV_X1 U249 ( .A(n1110), .ZN(n804) );
  AOI22_X1 U250 ( .A1(data_in[1]), .A2(n842), .B1(n1111), .B2(\mem[10][1] ), 
        .ZN(n1110) );
  INV_X1 U251 ( .A(n1109), .ZN(n803) );
  AOI22_X1 U252 ( .A1(data_in[2]), .A2(n842), .B1(n1111), .B2(\mem[10][2] ), 
        .ZN(n1109) );
  INV_X1 U253 ( .A(n1108), .ZN(n802) );
  AOI22_X1 U254 ( .A1(data_in[3]), .A2(n842), .B1(n1111), .B2(\mem[10][3] ), 
        .ZN(n1108) );
  INV_X1 U255 ( .A(n1107), .ZN(n801) );
  AOI22_X1 U256 ( .A1(data_in[4]), .A2(n842), .B1(n1111), .B2(\mem[10][4] ), 
        .ZN(n1107) );
  INV_X1 U257 ( .A(n1106), .ZN(n800) );
  AOI22_X1 U258 ( .A1(data_in[5]), .A2(n842), .B1(n1111), .B2(\mem[10][5] ), 
        .ZN(n1106) );
  INV_X1 U259 ( .A(n1105), .ZN(n799) );
  AOI22_X1 U260 ( .A1(data_in[6]), .A2(n842), .B1(n1111), .B2(\mem[10][6] ), 
        .ZN(n1105) );
  INV_X1 U261 ( .A(n1104), .ZN(n798) );
  AOI22_X1 U262 ( .A1(data_in[7]), .A2(n842), .B1(n1111), .B2(\mem[10][7] ), 
        .ZN(n1104) );
  INV_X1 U263 ( .A(n1103), .ZN(n797) );
  AOI22_X1 U264 ( .A1(data_in[0]), .A2(n827), .B1(n1102), .B2(\mem[11][0] ), 
        .ZN(n1103) );
  INV_X1 U265 ( .A(n1101), .ZN(n796) );
  AOI22_X1 U266 ( .A1(data_in[1]), .A2(n827), .B1(n1102), .B2(\mem[11][1] ), 
        .ZN(n1101) );
  INV_X1 U267 ( .A(n1100), .ZN(n795) );
  AOI22_X1 U268 ( .A1(data_in[2]), .A2(n827), .B1(n1102), .B2(\mem[11][2] ), 
        .ZN(n1100) );
  INV_X1 U269 ( .A(n1099), .ZN(n794) );
  AOI22_X1 U270 ( .A1(data_in[3]), .A2(n827), .B1(n1102), .B2(\mem[11][3] ), 
        .ZN(n1099) );
  INV_X1 U271 ( .A(n1098), .ZN(n793) );
  AOI22_X1 U272 ( .A1(data_in[4]), .A2(n827), .B1(n1102), .B2(\mem[11][4] ), 
        .ZN(n1098) );
  INV_X1 U273 ( .A(n1097), .ZN(n792) );
  AOI22_X1 U274 ( .A1(data_in[5]), .A2(n827), .B1(n1102), .B2(\mem[11][5] ), 
        .ZN(n1097) );
  INV_X1 U275 ( .A(n1096), .ZN(n791) );
  AOI22_X1 U276 ( .A1(data_in[6]), .A2(n827), .B1(n1102), .B2(\mem[11][6] ), 
        .ZN(n1096) );
  INV_X1 U277 ( .A(n1095), .ZN(n790) );
  AOI22_X1 U278 ( .A1(data_in[7]), .A2(n827), .B1(n1102), .B2(\mem[11][7] ), 
        .ZN(n1095) );
  INV_X1 U279 ( .A(n1094), .ZN(n789) );
  AOI22_X1 U280 ( .A1(data_in[0]), .A2(n830), .B1(n1093), .B2(\mem[12][0] ), 
        .ZN(n1094) );
  INV_X1 U281 ( .A(n1092), .ZN(n788) );
  AOI22_X1 U282 ( .A1(data_in[1]), .A2(n830), .B1(n1093), .B2(\mem[12][1] ), 
        .ZN(n1092) );
  INV_X1 U283 ( .A(n1091), .ZN(n787) );
  AOI22_X1 U284 ( .A1(data_in[2]), .A2(n830), .B1(n1093), .B2(\mem[12][2] ), 
        .ZN(n1091) );
  INV_X1 U285 ( .A(n1090), .ZN(n786) );
  AOI22_X1 U286 ( .A1(data_in[3]), .A2(n830), .B1(n1093), .B2(\mem[12][3] ), 
        .ZN(n1090) );
  INV_X1 U287 ( .A(n1089), .ZN(n785) );
  AOI22_X1 U288 ( .A1(data_in[4]), .A2(n830), .B1(n1093), .B2(\mem[12][4] ), 
        .ZN(n1089) );
  INV_X1 U289 ( .A(n1088), .ZN(n784) );
  AOI22_X1 U290 ( .A1(data_in[5]), .A2(n830), .B1(n1093), .B2(\mem[12][5] ), 
        .ZN(n1088) );
  INV_X1 U291 ( .A(n1087), .ZN(n783) );
  AOI22_X1 U292 ( .A1(data_in[6]), .A2(n830), .B1(n1093), .B2(\mem[12][6] ), 
        .ZN(n1087) );
  INV_X1 U293 ( .A(n1086), .ZN(n782) );
  AOI22_X1 U294 ( .A1(data_in[7]), .A2(n830), .B1(n1093), .B2(\mem[12][7] ), 
        .ZN(n1086) );
  INV_X1 U295 ( .A(n1085), .ZN(n781) );
  AOI22_X1 U296 ( .A1(data_in[0]), .A2(n839), .B1(n1084), .B2(\mem[13][0] ), 
        .ZN(n1085) );
  INV_X1 U297 ( .A(n1083), .ZN(n780) );
  AOI22_X1 U298 ( .A1(data_in[1]), .A2(n839), .B1(n1084), .B2(\mem[13][1] ), 
        .ZN(n1083) );
  INV_X1 U299 ( .A(n1082), .ZN(n779) );
  AOI22_X1 U300 ( .A1(data_in[2]), .A2(n839), .B1(n1084), .B2(\mem[13][2] ), 
        .ZN(n1082) );
  INV_X1 U301 ( .A(n1081), .ZN(n778) );
  AOI22_X1 U302 ( .A1(data_in[3]), .A2(n839), .B1(n1084), .B2(\mem[13][3] ), 
        .ZN(n1081) );
  INV_X1 U303 ( .A(n1080), .ZN(n777) );
  AOI22_X1 U304 ( .A1(data_in[4]), .A2(n839), .B1(n1084), .B2(\mem[13][4] ), 
        .ZN(n1080) );
  INV_X1 U305 ( .A(n1079), .ZN(n776) );
  AOI22_X1 U306 ( .A1(data_in[5]), .A2(n839), .B1(n1084), .B2(\mem[13][5] ), 
        .ZN(n1079) );
  INV_X1 U307 ( .A(n1078), .ZN(n775) );
  AOI22_X1 U308 ( .A1(data_in[6]), .A2(n839), .B1(n1084), .B2(\mem[13][6] ), 
        .ZN(n1078) );
  INV_X1 U309 ( .A(n1077), .ZN(n774) );
  AOI22_X1 U310 ( .A1(data_in[7]), .A2(n839), .B1(n1084), .B2(\mem[13][7] ), 
        .ZN(n1077) );
  INV_X1 U311 ( .A(n1076), .ZN(n773) );
  AOI22_X1 U312 ( .A1(data_in[0]), .A2(n833), .B1(n1075), .B2(\mem[14][0] ), 
        .ZN(n1076) );
  INV_X1 U313 ( .A(n1074), .ZN(n772) );
  AOI22_X1 U314 ( .A1(data_in[1]), .A2(n833), .B1(n1075), .B2(\mem[14][1] ), 
        .ZN(n1074) );
  INV_X1 U315 ( .A(n1073), .ZN(n771) );
  AOI22_X1 U316 ( .A1(data_in[2]), .A2(n833), .B1(n1075), .B2(\mem[14][2] ), 
        .ZN(n1073) );
  INV_X1 U317 ( .A(n1072), .ZN(n770) );
  AOI22_X1 U318 ( .A1(data_in[3]), .A2(n833), .B1(n1075), .B2(\mem[14][3] ), 
        .ZN(n1072) );
  INV_X1 U319 ( .A(n1071), .ZN(n769) );
  AOI22_X1 U320 ( .A1(data_in[4]), .A2(n833), .B1(n1075), .B2(\mem[14][4] ), 
        .ZN(n1071) );
  INV_X1 U321 ( .A(n1070), .ZN(n768) );
  AOI22_X1 U322 ( .A1(data_in[5]), .A2(n833), .B1(n1075), .B2(\mem[14][5] ), 
        .ZN(n1070) );
  INV_X1 U323 ( .A(n1069), .ZN(n767) );
  AOI22_X1 U324 ( .A1(data_in[6]), .A2(n833), .B1(n1075), .B2(\mem[14][6] ), 
        .ZN(n1069) );
  INV_X1 U325 ( .A(n1068), .ZN(n766) );
  AOI22_X1 U326 ( .A1(data_in[7]), .A2(n833), .B1(n1075), .B2(\mem[14][7] ), 
        .ZN(n1068) );
  INV_X1 U327 ( .A(n1067), .ZN(n765) );
  AOI22_X1 U328 ( .A1(data_in[0]), .A2(n836), .B1(n1066), .B2(\mem[15][0] ), 
        .ZN(n1067) );
  INV_X1 U329 ( .A(n1065), .ZN(n764) );
  AOI22_X1 U330 ( .A1(data_in[1]), .A2(n836), .B1(n1066), .B2(\mem[15][1] ), 
        .ZN(n1065) );
  INV_X1 U331 ( .A(n1064), .ZN(n763) );
  AOI22_X1 U332 ( .A1(data_in[2]), .A2(n836), .B1(n1066), .B2(\mem[15][2] ), 
        .ZN(n1064) );
  INV_X1 U333 ( .A(n1063), .ZN(n762) );
  AOI22_X1 U334 ( .A1(data_in[3]), .A2(n836), .B1(n1066), .B2(\mem[15][3] ), 
        .ZN(n1063) );
  INV_X1 U335 ( .A(n1062), .ZN(n761) );
  AOI22_X1 U336 ( .A1(data_in[4]), .A2(n836), .B1(n1066), .B2(\mem[15][4] ), 
        .ZN(n1062) );
  INV_X1 U337 ( .A(n1061), .ZN(n760) );
  AOI22_X1 U338 ( .A1(data_in[5]), .A2(n836), .B1(n1066), .B2(\mem[15][5] ), 
        .ZN(n1061) );
  INV_X1 U339 ( .A(n1060), .ZN(n759) );
  AOI22_X1 U340 ( .A1(data_in[6]), .A2(n836), .B1(n1066), .B2(\mem[15][6] ), 
        .ZN(n1060) );
  INV_X1 U341 ( .A(n1059), .ZN(n758) );
  AOI22_X1 U342 ( .A1(data_in[7]), .A2(n836), .B1(n1066), .B2(\mem[15][7] ), 
        .ZN(n1059) );
  INV_X1 U343 ( .A(n1058), .ZN(n757) );
  AOI22_X1 U344 ( .A1(data_in[0]), .A2(n844), .B1(n1057), .B2(\mem[16][0] ), 
        .ZN(n1058) );
  INV_X1 U345 ( .A(n1056), .ZN(n756) );
  AOI22_X1 U346 ( .A1(data_in[1]), .A2(n844), .B1(n1057), .B2(\mem[16][1] ), 
        .ZN(n1056) );
  INV_X1 U347 ( .A(n1055), .ZN(n755) );
  AOI22_X1 U348 ( .A1(data_in[2]), .A2(n844), .B1(n1057), .B2(\mem[16][2] ), 
        .ZN(n1055) );
  INV_X1 U349 ( .A(n1054), .ZN(n754) );
  AOI22_X1 U350 ( .A1(data_in[3]), .A2(n844), .B1(n1057), .B2(\mem[16][3] ), 
        .ZN(n1054) );
  INV_X1 U351 ( .A(n1053), .ZN(n753) );
  AOI22_X1 U352 ( .A1(data_in[4]), .A2(n844), .B1(n1057), .B2(\mem[16][4] ), 
        .ZN(n1053) );
  INV_X1 U353 ( .A(n1052), .ZN(n752) );
  AOI22_X1 U354 ( .A1(data_in[5]), .A2(n844), .B1(n1057), .B2(\mem[16][5] ), 
        .ZN(n1052) );
  INV_X1 U355 ( .A(n1051), .ZN(n751) );
  AOI22_X1 U356 ( .A1(data_in[6]), .A2(n844), .B1(n1057), .B2(\mem[16][6] ), 
        .ZN(n1051) );
  INV_X1 U357 ( .A(n1050), .ZN(n750) );
  AOI22_X1 U358 ( .A1(data_in[7]), .A2(n844), .B1(n1057), .B2(\mem[16][7] ), 
        .ZN(n1050) );
  INV_X1 U359 ( .A(n1048), .ZN(n749) );
  AOI22_X1 U360 ( .A1(data_in[0]), .A2(n823), .B1(n1047), .B2(\mem[17][0] ), 
        .ZN(n1048) );
  INV_X1 U361 ( .A(n1046), .ZN(n748) );
  AOI22_X1 U362 ( .A1(data_in[1]), .A2(n823), .B1(n1047), .B2(\mem[17][1] ), 
        .ZN(n1046) );
  INV_X1 U363 ( .A(n1045), .ZN(n747) );
  AOI22_X1 U364 ( .A1(data_in[2]), .A2(n823), .B1(n1047), .B2(\mem[17][2] ), 
        .ZN(n1045) );
  INV_X1 U365 ( .A(n1044), .ZN(n746) );
  AOI22_X1 U366 ( .A1(data_in[3]), .A2(n823), .B1(n1047), .B2(\mem[17][3] ), 
        .ZN(n1044) );
  INV_X1 U367 ( .A(n1043), .ZN(n745) );
  AOI22_X1 U368 ( .A1(data_in[4]), .A2(n823), .B1(n1047), .B2(\mem[17][4] ), 
        .ZN(n1043) );
  INV_X1 U369 ( .A(n1042), .ZN(n744) );
  AOI22_X1 U370 ( .A1(data_in[5]), .A2(n823), .B1(n1047), .B2(\mem[17][5] ), 
        .ZN(n1042) );
  INV_X1 U371 ( .A(n1041), .ZN(n743) );
  AOI22_X1 U372 ( .A1(data_in[6]), .A2(n823), .B1(n1047), .B2(\mem[17][6] ), 
        .ZN(n1041) );
  INV_X1 U373 ( .A(n1040), .ZN(n742) );
  AOI22_X1 U374 ( .A1(data_in[7]), .A2(n823), .B1(n1047), .B2(\mem[17][7] ), 
        .ZN(n1040) );
  INV_X1 U375 ( .A(n1039), .ZN(n741) );
  AOI22_X1 U376 ( .A1(data_in[0]), .A2(n841), .B1(n1038), .B2(\mem[18][0] ), 
        .ZN(n1039) );
  INV_X1 U377 ( .A(n1037), .ZN(n740) );
  AOI22_X1 U378 ( .A1(data_in[1]), .A2(n841), .B1(n1038), .B2(\mem[18][1] ), 
        .ZN(n1037) );
  INV_X1 U379 ( .A(n1036), .ZN(n739) );
  AOI22_X1 U380 ( .A1(data_in[2]), .A2(n841), .B1(n1038), .B2(\mem[18][2] ), 
        .ZN(n1036) );
  INV_X1 U381 ( .A(n1035), .ZN(n738) );
  AOI22_X1 U382 ( .A1(data_in[3]), .A2(n841), .B1(n1038), .B2(\mem[18][3] ), 
        .ZN(n1035) );
  INV_X1 U383 ( .A(n1034), .ZN(n737) );
  AOI22_X1 U384 ( .A1(data_in[4]), .A2(n841), .B1(n1038), .B2(\mem[18][4] ), 
        .ZN(n1034) );
  INV_X1 U385 ( .A(n1033), .ZN(n736) );
  AOI22_X1 U386 ( .A1(data_in[5]), .A2(n841), .B1(n1038), .B2(\mem[18][5] ), 
        .ZN(n1033) );
  INV_X1 U387 ( .A(n1032), .ZN(n735) );
  AOI22_X1 U388 ( .A1(data_in[6]), .A2(n841), .B1(n1038), .B2(\mem[18][6] ), 
        .ZN(n1032) );
  INV_X1 U389 ( .A(n1031), .ZN(n734) );
  AOI22_X1 U390 ( .A1(data_in[7]), .A2(n841), .B1(n1038), .B2(\mem[18][7] ), 
        .ZN(n1031) );
  INV_X1 U391 ( .A(n1030), .ZN(n733) );
  AOI22_X1 U392 ( .A1(data_in[0]), .A2(n826), .B1(n1029), .B2(\mem[19][0] ), 
        .ZN(n1030) );
  INV_X1 U393 ( .A(n1028), .ZN(n732) );
  AOI22_X1 U394 ( .A1(data_in[1]), .A2(n826), .B1(n1029), .B2(\mem[19][1] ), 
        .ZN(n1028) );
  INV_X1 U395 ( .A(n1027), .ZN(n731) );
  AOI22_X1 U396 ( .A1(data_in[2]), .A2(n826), .B1(n1029), .B2(\mem[19][2] ), 
        .ZN(n1027) );
  INV_X1 U397 ( .A(n1026), .ZN(n730) );
  AOI22_X1 U398 ( .A1(data_in[3]), .A2(n826), .B1(n1029), .B2(\mem[19][3] ), 
        .ZN(n1026) );
  INV_X1 U399 ( .A(n1025), .ZN(n729) );
  AOI22_X1 U400 ( .A1(data_in[4]), .A2(n826), .B1(n1029), .B2(\mem[19][4] ), 
        .ZN(n1025) );
  INV_X1 U401 ( .A(n1024), .ZN(n728) );
  AOI22_X1 U402 ( .A1(data_in[5]), .A2(n826), .B1(n1029), .B2(\mem[19][5] ), 
        .ZN(n1024) );
  INV_X1 U403 ( .A(n1023), .ZN(n727) );
  AOI22_X1 U404 ( .A1(data_in[6]), .A2(n826), .B1(n1029), .B2(\mem[19][6] ), 
        .ZN(n1023) );
  INV_X1 U405 ( .A(n1022), .ZN(n726) );
  AOI22_X1 U406 ( .A1(data_in[7]), .A2(n826), .B1(n1029), .B2(\mem[19][7] ), 
        .ZN(n1022) );
  INV_X1 U407 ( .A(n1021), .ZN(n725) );
  AOI22_X1 U408 ( .A1(data_in[0]), .A2(n829), .B1(n1020), .B2(\mem[20][0] ), 
        .ZN(n1021) );
  INV_X1 U409 ( .A(n1019), .ZN(n724) );
  AOI22_X1 U410 ( .A1(data_in[1]), .A2(n829), .B1(n1020), .B2(\mem[20][1] ), 
        .ZN(n1019) );
  INV_X1 U411 ( .A(n1018), .ZN(n723) );
  AOI22_X1 U412 ( .A1(data_in[2]), .A2(n829), .B1(n1020), .B2(\mem[20][2] ), 
        .ZN(n1018) );
  INV_X1 U413 ( .A(n1017), .ZN(n722) );
  AOI22_X1 U414 ( .A1(data_in[3]), .A2(n829), .B1(n1020), .B2(\mem[20][3] ), 
        .ZN(n1017) );
  INV_X1 U415 ( .A(n1016), .ZN(n721) );
  AOI22_X1 U416 ( .A1(data_in[4]), .A2(n829), .B1(n1020), .B2(\mem[20][4] ), 
        .ZN(n1016) );
  INV_X1 U417 ( .A(n1015), .ZN(n720) );
  AOI22_X1 U418 ( .A1(data_in[5]), .A2(n829), .B1(n1020), .B2(\mem[20][5] ), 
        .ZN(n1015) );
  INV_X1 U419 ( .A(n1014), .ZN(n719) );
  AOI22_X1 U420 ( .A1(data_in[6]), .A2(n829), .B1(n1020), .B2(\mem[20][6] ), 
        .ZN(n1014) );
  INV_X1 U421 ( .A(n1013), .ZN(n718) );
  AOI22_X1 U422 ( .A1(data_in[7]), .A2(n829), .B1(n1020), .B2(\mem[20][7] ), 
        .ZN(n1013) );
  INV_X1 U423 ( .A(n1012), .ZN(n717) );
  AOI22_X1 U424 ( .A1(data_in[0]), .A2(n838), .B1(n1011), .B2(\mem[21][0] ), 
        .ZN(n1012) );
  INV_X1 U425 ( .A(n1010), .ZN(n716) );
  AOI22_X1 U426 ( .A1(data_in[1]), .A2(n838), .B1(n1011), .B2(\mem[21][1] ), 
        .ZN(n1010) );
  INV_X1 U427 ( .A(n1009), .ZN(n715) );
  AOI22_X1 U428 ( .A1(data_in[2]), .A2(n838), .B1(n1011), .B2(\mem[21][2] ), 
        .ZN(n1009) );
  INV_X1 U429 ( .A(n1008), .ZN(n714) );
  AOI22_X1 U430 ( .A1(data_in[3]), .A2(n838), .B1(n1011), .B2(\mem[21][3] ), 
        .ZN(n1008) );
  INV_X1 U431 ( .A(n1007), .ZN(n713) );
  AOI22_X1 U432 ( .A1(data_in[4]), .A2(n838), .B1(n1011), .B2(\mem[21][4] ), 
        .ZN(n1007) );
  INV_X1 U433 ( .A(n1006), .ZN(n712) );
  AOI22_X1 U434 ( .A1(data_in[5]), .A2(n838), .B1(n1011), .B2(\mem[21][5] ), 
        .ZN(n1006) );
  INV_X1 U435 ( .A(n1005), .ZN(n711) );
  AOI22_X1 U436 ( .A1(data_in[6]), .A2(n838), .B1(n1011), .B2(\mem[21][6] ), 
        .ZN(n1005) );
  INV_X1 U437 ( .A(n1004), .ZN(n710) );
  AOI22_X1 U438 ( .A1(data_in[7]), .A2(n838), .B1(n1011), .B2(\mem[21][7] ), 
        .ZN(n1004) );
  INV_X1 U439 ( .A(n1003), .ZN(n709) );
  AOI22_X1 U440 ( .A1(data_in[0]), .A2(n832), .B1(n1002), .B2(\mem[22][0] ), 
        .ZN(n1003) );
  INV_X1 U441 ( .A(n1001), .ZN(n708) );
  AOI22_X1 U442 ( .A1(data_in[1]), .A2(n832), .B1(n1002), .B2(\mem[22][1] ), 
        .ZN(n1001) );
  INV_X1 U443 ( .A(n1000), .ZN(n707) );
  AOI22_X1 U444 ( .A1(data_in[2]), .A2(n832), .B1(n1002), .B2(\mem[22][2] ), 
        .ZN(n1000) );
  INV_X1 U445 ( .A(n999), .ZN(n706) );
  AOI22_X1 U446 ( .A1(data_in[3]), .A2(n832), .B1(n1002), .B2(\mem[22][3] ), 
        .ZN(n999) );
  INV_X1 U447 ( .A(n998), .ZN(n705) );
  AOI22_X1 U448 ( .A1(data_in[4]), .A2(n832), .B1(n1002), .B2(\mem[22][4] ), 
        .ZN(n998) );
  INV_X1 U449 ( .A(n997), .ZN(n704) );
  AOI22_X1 U450 ( .A1(data_in[5]), .A2(n832), .B1(n1002), .B2(\mem[22][5] ), 
        .ZN(n997) );
  INV_X1 U451 ( .A(n996), .ZN(n703) );
  AOI22_X1 U452 ( .A1(data_in[6]), .A2(n832), .B1(n1002), .B2(\mem[22][6] ), 
        .ZN(n996) );
  INV_X1 U453 ( .A(n995), .ZN(n702) );
  AOI22_X1 U454 ( .A1(data_in[7]), .A2(n832), .B1(n1002), .B2(\mem[22][7] ), 
        .ZN(n995) );
  INV_X1 U455 ( .A(n994), .ZN(n701) );
  AOI22_X1 U456 ( .A1(data_in[0]), .A2(n835), .B1(n993), .B2(\mem[23][0] ), 
        .ZN(n994) );
  INV_X1 U457 ( .A(n992), .ZN(n700) );
  AOI22_X1 U458 ( .A1(data_in[1]), .A2(n835), .B1(n993), .B2(\mem[23][1] ), 
        .ZN(n992) );
  INV_X1 U459 ( .A(n991), .ZN(n699) );
  AOI22_X1 U460 ( .A1(data_in[2]), .A2(n835), .B1(n993), .B2(\mem[23][2] ), 
        .ZN(n991) );
  INV_X1 U461 ( .A(n990), .ZN(n698) );
  AOI22_X1 U462 ( .A1(data_in[3]), .A2(n835), .B1(n993), .B2(\mem[23][3] ), 
        .ZN(n990) );
  INV_X1 U463 ( .A(n989), .ZN(n697) );
  AOI22_X1 U464 ( .A1(data_in[4]), .A2(n835), .B1(n993), .B2(\mem[23][4] ), 
        .ZN(n989) );
  INV_X1 U465 ( .A(n988), .ZN(n696) );
  AOI22_X1 U466 ( .A1(data_in[5]), .A2(n835), .B1(n993), .B2(\mem[23][5] ), 
        .ZN(n988) );
  INV_X1 U467 ( .A(n987), .ZN(n695) );
  AOI22_X1 U468 ( .A1(data_in[6]), .A2(n835), .B1(n993), .B2(\mem[23][6] ), 
        .ZN(n987) );
  INV_X1 U469 ( .A(n986), .ZN(n694) );
  AOI22_X1 U470 ( .A1(data_in[7]), .A2(n835), .B1(n993), .B2(\mem[23][7] ), 
        .ZN(n986) );
  INV_X1 U471 ( .A(n985), .ZN(n693) );
  AOI22_X1 U472 ( .A1(data_in[0]), .A2(n843), .B1(n984), .B2(\mem[24][0] ), 
        .ZN(n985) );
  INV_X1 U473 ( .A(n983), .ZN(n692) );
  AOI22_X1 U474 ( .A1(data_in[1]), .A2(n843), .B1(n984), .B2(\mem[24][1] ), 
        .ZN(n983) );
  INV_X1 U475 ( .A(n982), .ZN(n691) );
  AOI22_X1 U476 ( .A1(data_in[2]), .A2(n843), .B1(n984), .B2(\mem[24][2] ), 
        .ZN(n982) );
  INV_X1 U477 ( .A(n981), .ZN(n690) );
  AOI22_X1 U478 ( .A1(data_in[3]), .A2(n843), .B1(n984), .B2(\mem[24][3] ), 
        .ZN(n981) );
  INV_X1 U479 ( .A(n980), .ZN(n689) );
  AOI22_X1 U480 ( .A1(data_in[4]), .A2(n843), .B1(n984), .B2(\mem[24][4] ), 
        .ZN(n980) );
  INV_X1 U481 ( .A(n979), .ZN(n688) );
  AOI22_X1 U482 ( .A1(data_in[5]), .A2(n843), .B1(n984), .B2(\mem[24][5] ), 
        .ZN(n979) );
  INV_X1 U483 ( .A(n978), .ZN(n687) );
  AOI22_X1 U484 ( .A1(data_in[6]), .A2(n843), .B1(n984), .B2(\mem[24][6] ), 
        .ZN(n978) );
  INV_X1 U485 ( .A(n977), .ZN(n686) );
  AOI22_X1 U486 ( .A1(data_in[7]), .A2(n843), .B1(n984), .B2(\mem[24][7] ), 
        .ZN(n977) );
  INV_X1 U487 ( .A(n975), .ZN(n685) );
  AOI22_X1 U488 ( .A1(data_in[0]), .A2(n822), .B1(n974), .B2(\mem[25][0] ), 
        .ZN(n975) );
  INV_X1 U489 ( .A(n973), .ZN(n684) );
  AOI22_X1 U490 ( .A1(data_in[1]), .A2(n822), .B1(n974), .B2(\mem[25][1] ), 
        .ZN(n973) );
  INV_X1 U491 ( .A(n972), .ZN(n683) );
  AOI22_X1 U492 ( .A1(data_in[2]), .A2(n822), .B1(n974), .B2(\mem[25][2] ), 
        .ZN(n972) );
  INV_X1 U493 ( .A(n971), .ZN(n682) );
  AOI22_X1 U494 ( .A1(data_in[3]), .A2(n822), .B1(n974), .B2(\mem[25][3] ), 
        .ZN(n971) );
  INV_X1 U495 ( .A(n970), .ZN(n681) );
  AOI22_X1 U496 ( .A1(data_in[4]), .A2(n822), .B1(n974), .B2(\mem[25][4] ), 
        .ZN(n970) );
  INV_X1 U497 ( .A(n969), .ZN(n680) );
  AOI22_X1 U498 ( .A1(data_in[5]), .A2(n822), .B1(n974), .B2(\mem[25][5] ), 
        .ZN(n969) );
  INV_X1 U499 ( .A(n968), .ZN(n679) );
  AOI22_X1 U500 ( .A1(data_in[6]), .A2(n822), .B1(n974), .B2(\mem[25][6] ), 
        .ZN(n968) );
  INV_X1 U501 ( .A(n967), .ZN(n678) );
  AOI22_X1 U502 ( .A1(data_in[7]), .A2(n822), .B1(n974), .B2(\mem[25][7] ), 
        .ZN(n967) );
  INV_X1 U503 ( .A(n966), .ZN(n677) );
  AOI22_X1 U504 ( .A1(data_in[0]), .A2(n840), .B1(n965), .B2(\mem[26][0] ), 
        .ZN(n966) );
  INV_X1 U505 ( .A(n964), .ZN(n676) );
  AOI22_X1 U506 ( .A1(data_in[1]), .A2(n840), .B1(n965), .B2(\mem[26][1] ), 
        .ZN(n964) );
  INV_X1 U507 ( .A(n963), .ZN(n675) );
  AOI22_X1 U508 ( .A1(data_in[2]), .A2(n840), .B1(n965), .B2(\mem[26][2] ), 
        .ZN(n963) );
  INV_X1 U509 ( .A(n962), .ZN(n674) );
  AOI22_X1 U510 ( .A1(data_in[3]), .A2(n840), .B1(n965), .B2(\mem[26][3] ), 
        .ZN(n962) );
  INV_X1 U511 ( .A(n961), .ZN(n673) );
  AOI22_X1 U512 ( .A1(data_in[4]), .A2(n840), .B1(n965), .B2(\mem[26][4] ), 
        .ZN(n961) );
  INV_X1 U513 ( .A(n960), .ZN(n672) );
  AOI22_X1 U514 ( .A1(data_in[5]), .A2(n840), .B1(n965), .B2(\mem[26][5] ), 
        .ZN(n960) );
  INV_X1 U515 ( .A(n959), .ZN(n671) );
  AOI22_X1 U516 ( .A1(data_in[6]), .A2(n840), .B1(n965), .B2(\mem[26][6] ), 
        .ZN(n959) );
  INV_X1 U517 ( .A(n958), .ZN(n670) );
  AOI22_X1 U518 ( .A1(data_in[7]), .A2(n840), .B1(n965), .B2(\mem[26][7] ), 
        .ZN(n958) );
  INV_X1 U519 ( .A(n957), .ZN(n669) );
  AOI22_X1 U520 ( .A1(data_in[0]), .A2(n825), .B1(n956), .B2(\mem[27][0] ), 
        .ZN(n957) );
  INV_X1 U521 ( .A(n955), .ZN(n668) );
  AOI22_X1 U522 ( .A1(data_in[1]), .A2(n825), .B1(n956), .B2(\mem[27][1] ), 
        .ZN(n955) );
  INV_X1 U523 ( .A(n954), .ZN(n667) );
  AOI22_X1 U524 ( .A1(data_in[2]), .A2(n825), .B1(n956), .B2(\mem[27][2] ), 
        .ZN(n954) );
  INV_X1 U525 ( .A(n953), .ZN(n666) );
  AOI22_X1 U526 ( .A1(data_in[3]), .A2(n825), .B1(n956), .B2(\mem[27][3] ), 
        .ZN(n953) );
  INV_X1 U527 ( .A(n952), .ZN(n665) );
  AOI22_X1 U528 ( .A1(data_in[4]), .A2(n825), .B1(n956), .B2(\mem[27][4] ), 
        .ZN(n952) );
  INV_X1 U529 ( .A(n951), .ZN(n664) );
  AOI22_X1 U530 ( .A1(data_in[5]), .A2(n825), .B1(n956), .B2(\mem[27][5] ), 
        .ZN(n951) );
  INV_X1 U531 ( .A(n950), .ZN(n663) );
  AOI22_X1 U532 ( .A1(data_in[6]), .A2(n825), .B1(n956), .B2(\mem[27][6] ), 
        .ZN(n950) );
  INV_X1 U533 ( .A(n949), .ZN(n662) );
  AOI22_X1 U534 ( .A1(data_in[7]), .A2(n825), .B1(n956), .B2(\mem[27][7] ), 
        .ZN(n949) );
  INV_X1 U535 ( .A(n948), .ZN(n661) );
  AOI22_X1 U536 ( .A1(data_in[0]), .A2(n828), .B1(n947), .B2(\mem[28][0] ), 
        .ZN(n948) );
  INV_X1 U537 ( .A(n946), .ZN(n660) );
  AOI22_X1 U538 ( .A1(data_in[1]), .A2(n828), .B1(n947), .B2(\mem[28][1] ), 
        .ZN(n946) );
  INV_X1 U539 ( .A(n945), .ZN(n659) );
  AOI22_X1 U540 ( .A1(data_in[2]), .A2(n828), .B1(n947), .B2(\mem[28][2] ), 
        .ZN(n945) );
  INV_X1 U541 ( .A(n944), .ZN(n658) );
  AOI22_X1 U542 ( .A1(data_in[3]), .A2(n828), .B1(n947), .B2(\mem[28][3] ), 
        .ZN(n944) );
  INV_X1 U543 ( .A(n943), .ZN(n657) );
  AOI22_X1 U544 ( .A1(data_in[4]), .A2(n828), .B1(n947), .B2(\mem[28][4] ), 
        .ZN(n943) );
  INV_X1 U545 ( .A(n942), .ZN(n656) );
  AOI22_X1 U546 ( .A1(data_in[5]), .A2(n828), .B1(n947), .B2(\mem[28][5] ), 
        .ZN(n942) );
  INV_X1 U547 ( .A(n941), .ZN(n655) );
  AOI22_X1 U548 ( .A1(data_in[6]), .A2(n828), .B1(n947), .B2(\mem[28][6] ), 
        .ZN(n941) );
  INV_X1 U549 ( .A(n940), .ZN(n654) );
  AOI22_X1 U550 ( .A1(data_in[7]), .A2(n828), .B1(n947), .B2(\mem[28][7] ), 
        .ZN(n940) );
  INV_X1 U551 ( .A(n939), .ZN(n653) );
  AOI22_X1 U552 ( .A1(data_in[0]), .A2(n837), .B1(n938), .B2(\mem[29][0] ), 
        .ZN(n939) );
  INV_X1 U553 ( .A(n937), .ZN(n652) );
  AOI22_X1 U554 ( .A1(data_in[1]), .A2(n837), .B1(n938), .B2(\mem[29][1] ), 
        .ZN(n937) );
  INV_X1 U555 ( .A(n936), .ZN(n651) );
  AOI22_X1 U556 ( .A1(data_in[2]), .A2(n837), .B1(n938), .B2(\mem[29][2] ), 
        .ZN(n936) );
  INV_X1 U557 ( .A(n935), .ZN(n650) );
  AOI22_X1 U558 ( .A1(data_in[3]), .A2(n837), .B1(n938), .B2(\mem[29][3] ), 
        .ZN(n935) );
  INV_X1 U559 ( .A(n934), .ZN(n649) );
  AOI22_X1 U560 ( .A1(data_in[4]), .A2(n837), .B1(n938), .B2(\mem[29][4] ), 
        .ZN(n934) );
  INV_X1 U561 ( .A(n933), .ZN(n648) );
  AOI22_X1 U562 ( .A1(data_in[5]), .A2(n837), .B1(n938), .B2(\mem[29][5] ), 
        .ZN(n933) );
  INV_X1 U563 ( .A(n932), .ZN(n647) );
  AOI22_X1 U564 ( .A1(data_in[6]), .A2(n837), .B1(n938), .B2(\mem[29][6] ), 
        .ZN(n932) );
  INV_X1 U565 ( .A(n931), .ZN(n646) );
  AOI22_X1 U566 ( .A1(data_in[7]), .A2(n837), .B1(n938), .B2(\mem[29][7] ), 
        .ZN(n931) );
  INV_X1 U567 ( .A(n930), .ZN(n645) );
  AOI22_X1 U568 ( .A1(data_in[0]), .A2(n831), .B1(n929), .B2(\mem[30][0] ), 
        .ZN(n930) );
  INV_X1 U569 ( .A(n928), .ZN(n644) );
  AOI22_X1 U570 ( .A1(data_in[1]), .A2(n831), .B1(n929), .B2(\mem[30][1] ), 
        .ZN(n928) );
  INV_X1 U571 ( .A(n927), .ZN(n643) );
  AOI22_X1 U572 ( .A1(data_in[2]), .A2(n831), .B1(n929), .B2(\mem[30][2] ), 
        .ZN(n927) );
  INV_X1 U573 ( .A(n926), .ZN(n642) );
  AOI22_X1 U574 ( .A1(data_in[3]), .A2(n831), .B1(n929), .B2(\mem[30][3] ), 
        .ZN(n926) );
  INV_X1 U575 ( .A(n925), .ZN(n641) );
  AOI22_X1 U576 ( .A1(data_in[4]), .A2(n831), .B1(n929), .B2(\mem[30][4] ), 
        .ZN(n925) );
  INV_X1 U577 ( .A(n924), .ZN(n640) );
  AOI22_X1 U578 ( .A1(data_in[5]), .A2(n831), .B1(n929), .B2(\mem[30][5] ), 
        .ZN(n924) );
  INV_X1 U579 ( .A(n923), .ZN(n639) );
  AOI22_X1 U580 ( .A1(data_in[6]), .A2(n831), .B1(n929), .B2(\mem[30][6] ), 
        .ZN(n923) );
  INV_X1 U581 ( .A(n922), .ZN(n638) );
  AOI22_X1 U582 ( .A1(data_in[7]), .A2(n831), .B1(n929), .B2(\mem[30][7] ), 
        .ZN(n922) );
  INV_X1 U583 ( .A(n921), .ZN(n637) );
  AOI22_X1 U584 ( .A1(data_in[0]), .A2(n834), .B1(n920), .B2(\mem[31][0] ), 
        .ZN(n921) );
  INV_X1 U585 ( .A(n919), .ZN(n636) );
  AOI22_X1 U586 ( .A1(data_in[1]), .A2(n834), .B1(n920), .B2(\mem[31][1] ), 
        .ZN(n919) );
  INV_X1 U587 ( .A(n918), .ZN(n635) );
  AOI22_X1 U588 ( .A1(data_in[2]), .A2(n834), .B1(n920), .B2(\mem[31][2] ), 
        .ZN(n918) );
  INV_X1 U589 ( .A(n917), .ZN(n634) );
  AOI22_X1 U590 ( .A1(data_in[3]), .A2(n834), .B1(n920), .B2(\mem[31][3] ), 
        .ZN(n917) );
  INV_X1 U591 ( .A(n916), .ZN(n633) );
  AOI22_X1 U592 ( .A1(data_in[4]), .A2(n834), .B1(n920), .B2(\mem[31][4] ), 
        .ZN(n916) );
  INV_X1 U593 ( .A(n915), .ZN(n632) );
  AOI22_X1 U594 ( .A1(data_in[5]), .A2(n834), .B1(n920), .B2(\mem[31][5] ), 
        .ZN(n915) );
  INV_X1 U595 ( .A(n914), .ZN(n631) );
  AOI22_X1 U596 ( .A1(data_in[6]), .A2(n834), .B1(n920), .B2(\mem[31][6] ), 
        .ZN(n914) );
  INV_X1 U597 ( .A(n913), .ZN(n630) );
  AOI22_X1 U598 ( .A1(data_in[7]), .A2(n834), .B1(n920), .B2(\mem[31][7] ), 
        .ZN(n913) );
  MUX2_X1 U599 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n614), .Z(n4) );
  MUX2_X1 U600 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n614), .Z(n5) );
  MUX2_X1 U601 ( .A(n5), .B(n4), .S(n611), .Z(n6) );
  MUX2_X1 U602 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n614), .Z(n7) );
  MUX2_X1 U603 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n614), .Z(n8) );
  MUX2_X1 U604 ( .A(n8), .B(n7), .S(n611), .Z(n9) );
  MUX2_X1 U605 ( .A(n9), .B(n6), .S(n609), .Z(n10) );
  MUX2_X1 U606 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n614), .Z(n11) );
  MUX2_X1 U607 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n614), .Z(n12) );
  MUX2_X1 U608 ( .A(n12), .B(n11), .S(n611), .Z(n13) );
  MUX2_X1 U609 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n614), .Z(n14) );
  MUX2_X1 U610 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n614), .Z(n15) );
  MUX2_X1 U611 ( .A(n15), .B(n14), .S(n612), .Z(n16) );
  MUX2_X1 U612 ( .A(n16), .B(n13), .S(n609), .Z(n17) );
  MUX2_X1 U613 ( .A(n17), .B(n10), .S(N13), .Z(n18) );
  MUX2_X1 U614 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n616), .Z(n19) );
  MUX2_X1 U615 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n618), .Z(n20) );
  MUX2_X1 U616 ( .A(n20), .B(n19), .S(n611), .Z(n21) );
  MUX2_X1 U617 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n615), .Z(n22) );
  MUX2_X1 U618 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n23) );
  MUX2_X1 U619 ( .A(n23), .B(n22), .S(n611), .Z(n24) );
  MUX2_X1 U620 ( .A(n24), .B(n21), .S(n609), .Z(n25) );
  MUX2_X1 U621 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n616), .Z(n26) );
  MUX2_X1 U622 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n27) );
  MUX2_X1 U623 ( .A(n27), .B(n26), .S(n611), .Z(n28) );
  MUX2_X1 U624 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n619), .Z(n29) );
  MUX2_X1 U625 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n30) );
  MUX2_X1 U626 ( .A(n30), .B(n29), .S(n611), .Z(n31) );
  MUX2_X1 U627 ( .A(n31), .B(n28), .S(n609), .Z(n32) );
  MUX2_X1 U628 ( .A(n32), .B(n25), .S(N13), .Z(n33) );
  MUX2_X1 U629 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(N10), .Z(n34) );
  MUX2_X1 U630 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n618), .Z(n35) );
  MUX2_X1 U631 ( .A(n35), .B(n34), .S(n611), .Z(n36) );
  MUX2_X1 U632 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n619), .Z(n37) );
  MUX2_X1 U633 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n619), .Z(n38) );
  MUX2_X1 U634 ( .A(n38), .B(n37), .S(n611), .Z(n39) );
  MUX2_X1 U635 ( .A(n39), .B(n36), .S(n609), .Z(n40) );
  MUX2_X1 U636 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n619), .Z(n41) );
  MUX2_X1 U637 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n615), .Z(n42) );
  MUX2_X1 U638 ( .A(n42), .B(n41), .S(n611), .Z(n43) );
  MUX2_X1 U639 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n614), .Z(n44) );
  MUX2_X1 U640 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n619), .Z(n45) );
  MUX2_X1 U641 ( .A(n45), .B(n44), .S(n611), .Z(n46) );
  MUX2_X1 U642 ( .A(n46), .B(n43), .S(n609), .Z(n47) );
  MUX2_X1 U643 ( .A(n47), .B(n40), .S(N13), .Z(n48) );
  MUX2_X1 U644 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n614), .Z(n49) );
  MUX2_X1 U645 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n614), .Z(n50) );
  MUX2_X1 U646 ( .A(n50), .B(n49), .S(n611), .Z(n51) );
  MUX2_X1 U647 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n614), .Z(n52) );
  MUX2_X1 U648 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(N10), .Z(n53) );
  MUX2_X1 U649 ( .A(n53), .B(n52), .S(n611), .Z(n54) );
  MUX2_X1 U650 ( .A(n54), .B(n51), .S(n609), .Z(n55) );
  MUX2_X1 U651 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n614), .Z(n56) );
  MUX2_X1 U652 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n614), .Z(n57) );
  MUX2_X1 U653 ( .A(n57), .B(n56), .S(n611), .Z(n58) );
  MUX2_X1 U654 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n615), .Z(n59) );
  MUX2_X1 U655 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n615), .Z(n60) );
  MUX2_X1 U656 ( .A(n60), .B(n59), .S(n611), .Z(n61) );
  MUX2_X1 U657 ( .A(n61), .B(n58), .S(n609), .Z(n62) );
  MUX2_X1 U658 ( .A(n62), .B(n55), .S(N13), .Z(n63) );
  MUX2_X1 U659 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n615), .Z(n64) );
  MUX2_X1 U660 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n615), .Z(n65) );
  MUX2_X1 U661 ( .A(n65), .B(n64), .S(n612), .Z(n66) );
  MUX2_X1 U662 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n615), .Z(n67) );
  MUX2_X1 U663 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n615), .Z(n68) );
  MUX2_X1 U664 ( .A(n68), .B(n67), .S(n612), .Z(n69) );
  MUX2_X1 U665 ( .A(n69), .B(n66), .S(n610), .Z(n70) );
  MUX2_X1 U666 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n615), .Z(n71) );
  MUX2_X1 U667 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n615), .Z(n72) );
  MUX2_X1 U668 ( .A(n72), .B(n71), .S(n612), .Z(n73) );
  MUX2_X1 U669 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n615), .Z(n74) );
  MUX2_X1 U670 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n615), .Z(n75) );
  MUX2_X1 U671 ( .A(n75), .B(n74), .S(n612), .Z(n76) );
  MUX2_X1 U672 ( .A(n76), .B(n73), .S(n610), .Z(n77) );
  MUX2_X1 U673 ( .A(n77), .B(n70), .S(N13), .Z(n78) );
  MUX2_X1 U674 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n615), .Z(n79) );
  MUX2_X1 U675 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n615), .Z(n80) );
  MUX2_X1 U676 ( .A(n80), .B(n79), .S(n612), .Z(n81) );
  MUX2_X1 U677 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n615), .Z(n82) );
  MUX2_X1 U678 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n615), .Z(n83) );
  MUX2_X1 U679 ( .A(n83), .B(n82), .S(n612), .Z(n84) );
  MUX2_X1 U680 ( .A(n84), .B(n81), .S(n610), .Z(n85) );
  MUX2_X1 U681 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n616), .Z(n86) );
  MUX2_X1 U682 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n616), .Z(n87) );
  MUX2_X1 U683 ( .A(n87), .B(n86), .S(n612), .Z(n88) );
  MUX2_X1 U684 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n616), .Z(n89) );
  MUX2_X1 U685 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n616), .Z(n90) );
  MUX2_X1 U686 ( .A(n90), .B(n89), .S(n612), .Z(n91) );
  MUX2_X1 U687 ( .A(n91), .B(n88), .S(n610), .Z(n92) );
  MUX2_X1 U688 ( .A(n92), .B(n85), .S(N13), .Z(n93) );
  MUX2_X1 U689 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n616), .Z(n94) );
  MUX2_X1 U690 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n616), .Z(n95) );
  MUX2_X1 U691 ( .A(n95), .B(n94), .S(n612), .Z(n96) );
  MUX2_X1 U692 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n616), .Z(n97) );
  MUX2_X1 U693 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n616), .Z(n98) );
  MUX2_X1 U694 ( .A(n98), .B(n97), .S(n612), .Z(n99) );
  MUX2_X1 U695 ( .A(n99), .B(n96), .S(n610), .Z(n100) );
  MUX2_X1 U696 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n616), .Z(n101) );
  MUX2_X1 U697 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n616), .Z(n102) );
  MUX2_X1 U698 ( .A(n102), .B(n101), .S(n612), .Z(n103) );
  MUX2_X1 U699 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n616), .Z(n104) );
  MUX2_X1 U700 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n616), .Z(n105) );
  MUX2_X1 U701 ( .A(n105), .B(n104), .S(n612), .Z(n106) );
  MUX2_X1 U702 ( .A(n106), .B(n103), .S(n610), .Z(n107) );
  MUX2_X1 U703 ( .A(n107), .B(n100), .S(N13), .Z(n108) );
  MUX2_X1 U704 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n619), .Z(n109) );
  MUX2_X1 U705 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n619), .Z(n110) );
  MUX2_X1 U706 ( .A(n110), .B(n109), .S(n613), .Z(n111) );
  MUX2_X1 U707 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n619), .Z(n112) );
  MUX2_X1 U708 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n619), .Z(n113) );
  MUX2_X1 U709 ( .A(n113), .B(n112), .S(n613), .Z(n114) );
  MUX2_X1 U710 ( .A(n114), .B(n111), .S(n610), .Z(n115) );
  MUX2_X1 U711 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n619), .Z(n116) );
  MUX2_X1 U712 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n619), .Z(n117) );
  MUX2_X1 U713 ( .A(n117), .B(n116), .S(n613), .Z(n118) );
  MUX2_X1 U714 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n619), .Z(n119) );
  MUX2_X1 U715 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n619), .Z(n120) );
  MUX2_X1 U716 ( .A(n120), .B(n119), .S(n613), .Z(n121) );
  MUX2_X1 U717 ( .A(n121), .B(n118), .S(n610), .Z(n122) );
  MUX2_X1 U718 ( .A(n122), .B(n115), .S(N13), .Z(n123) );
  MUX2_X1 U719 ( .A(n123), .B(n108), .S(N14), .Z(N19) );
  MUX2_X1 U720 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n619), .Z(n124) );
  MUX2_X1 U721 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n619), .Z(n125) );
  MUX2_X1 U722 ( .A(n125), .B(n124), .S(n613), .Z(n126) );
  MUX2_X1 U723 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n619), .Z(n127) );
  MUX2_X1 U724 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n619), .Z(n128) );
  MUX2_X1 U725 ( .A(n128), .B(n127), .S(n613), .Z(n129) );
  MUX2_X1 U726 ( .A(n129), .B(n126), .S(n610), .Z(n130) );
  MUX2_X1 U727 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n616), .Z(n131) );
  MUX2_X1 U728 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n617), .Z(n132) );
  MUX2_X1 U729 ( .A(n132), .B(n131), .S(n613), .Z(n133) );
  MUX2_X1 U730 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n614), .Z(n134) );
  MUX2_X1 U731 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n619), .Z(n135) );
  MUX2_X1 U732 ( .A(n135), .B(n134), .S(n613), .Z(n136) );
  MUX2_X1 U733 ( .A(n136), .B(n133), .S(n610), .Z(n137) );
  MUX2_X1 U734 ( .A(n137), .B(n130), .S(N13), .Z(n138) );
  MUX2_X1 U735 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n614), .Z(n139) );
  MUX2_X1 U736 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n616), .Z(n140) );
  MUX2_X1 U737 ( .A(n140), .B(n139), .S(n613), .Z(n141) );
  MUX2_X1 U738 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n614), .Z(n142) );
  MUX2_X1 U739 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n618), .Z(n143) );
  MUX2_X1 U740 ( .A(n143), .B(n142), .S(n613), .Z(n144) );
  MUX2_X1 U741 ( .A(n144), .B(n141), .S(n610), .Z(n145) );
  MUX2_X1 U742 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n616), .Z(n146) );
  MUX2_X1 U743 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n618), .Z(n147) );
  MUX2_X1 U744 ( .A(n147), .B(n146), .S(n613), .Z(n148) );
  MUX2_X1 U745 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n617), .Z(n149) );
  MUX2_X1 U746 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n619), .Z(n150) );
  MUX2_X1 U747 ( .A(n150), .B(n149), .S(n613), .Z(n151) );
  MUX2_X1 U748 ( .A(n151), .B(n148), .S(n610), .Z(n152) );
  MUX2_X1 U749 ( .A(n152), .B(n145), .S(N13), .Z(n153) );
  MUX2_X1 U750 ( .A(n153), .B(n138), .S(N14), .Z(N18) );
  MUX2_X1 U751 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n616), .Z(n154) );
  MUX2_X1 U752 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n614), .Z(n155) );
  MUX2_X1 U753 ( .A(n155), .B(n154), .S(n612), .Z(n156) );
  MUX2_X1 U754 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n614), .Z(n157) );
  MUX2_X1 U755 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n614), .Z(n158) );
  MUX2_X1 U756 ( .A(n158), .B(n157), .S(n611), .Z(n159) );
  MUX2_X1 U757 ( .A(n159), .B(n156), .S(n609), .Z(n160) );
  MUX2_X1 U758 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n616), .Z(n161) );
  MUX2_X1 U759 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n616), .Z(n162) );
  MUX2_X1 U760 ( .A(n162), .B(n161), .S(n612), .Z(n163) );
  MUX2_X1 U761 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n614), .Z(n164) );
  MUX2_X1 U762 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n616), .Z(n165) );
  MUX2_X1 U763 ( .A(n165), .B(n164), .S(n613), .Z(n166) );
  MUX2_X1 U764 ( .A(n166), .B(n163), .S(n610), .Z(n167) );
  MUX2_X1 U765 ( .A(n167), .B(n160), .S(N13), .Z(n168) );
  MUX2_X1 U766 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n614), .Z(n169) );
  MUX2_X1 U767 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n616), .Z(n170) );
  MUX2_X1 U768 ( .A(n170), .B(n169), .S(n611), .Z(n171) );
  MUX2_X1 U769 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n616), .Z(n172) );
  MUX2_X1 U770 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n614), .Z(n173) );
  MUX2_X1 U771 ( .A(n173), .B(n172), .S(n612), .Z(n174) );
  MUX2_X1 U772 ( .A(n174), .B(n171), .S(n609), .Z(n175) );
  MUX2_X1 U773 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n617), .Z(n176) );
  MUX2_X1 U774 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n617), .Z(n177) );
  MUX2_X1 U775 ( .A(n177), .B(n176), .S(n613), .Z(n178) );
  MUX2_X1 U776 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n617), .Z(n179) );
  MUX2_X1 U777 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n617), .Z(n180) );
  MUX2_X1 U778 ( .A(n180), .B(n179), .S(n612), .Z(n181) );
  MUX2_X1 U779 ( .A(n181), .B(n178), .S(n609), .Z(n182) );
  MUX2_X1 U780 ( .A(n182), .B(n175), .S(N13), .Z(n183) );
  MUX2_X1 U781 ( .A(n183), .B(n168), .S(N14), .Z(N17) );
  MUX2_X1 U782 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n617), .Z(n184) );
  MUX2_X1 U783 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n617), .Z(n185) );
  MUX2_X1 U784 ( .A(n185), .B(n184), .S(n613), .Z(n186) );
  MUX2_X1 U785 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n617), .Z(n187) );
  MUX2_X1 U786 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n617), .Z(n188) );
  MUX2_X1 U787 ( .A(n188), .B(n187), .S(n612), .Z(n189) );
  MUX2_X1 U788 ( .A(n189), .B(n186), .S(n609), .Z(n190) );
  MUX2_X1 U789 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n617), .Z(n191) );
  MUX2_X1 U790 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n617), .Z(n192) );
  MUX2_X1 U791 ( .A(n192), .B(n191), .S(n613), .Z(n193) );
  MUX2_X1 U792 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n617), .Z(n194) );
  MUX2_X1 U793 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n617), .Z(n195) );
  MUX2_X1 U794 ( .A(n195), .B(n194), .S(n611), .Z(n196) );
  MUX2_X1 U795 ( .A(n196), .B(n193), .S(n610), .Z(n197) );
  MUX2_X1 U796 ( .A(n197), .B(n190), .S(N13), .Z(n198) );
  MUX2_X1 U797 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n618), .Z(n199) );
  MUX2_X1 U798 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n618), .Z(n200) );
  MUX2_X1 U799 ( .A(n200), .B(n199), .S(N11), .Z(n201) );
  MUX2_X1 U800 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n618), .Z(n202) );
  MUX2_X1 U801 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n618), .Z(n203) );
  MUX2_X1 U802 ( .A(n203), .B(n202), .S(N11), .Z(n204) );
  MUX2_X1 U803 ( .A(n204), .B(n201), .S(n609), .Z(n205) );
  MUX2_X1 U804 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n618), .Z(n206) );
  MUX2_X1 U805 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n618), .Z(n207) );
  MUX2_X1 U806 ( .A(n207), .B(n206), .S(n612), .Z(n208) );
  MUX2_X1 U807 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n618), .Z(n209) );
  MUX2_X1 U808 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n618), .Z(n210) );
  MUX2_X1 U809 ( .A(n210), .B(n209), .S(n612), .Z(n211) );
  MUX2_X1 U810 ( .A(n211), .B(n208), .S(n609), .Z(n212) );
  MUX2_X1 U811 ( .A(n212), .B(n205), .S(N13), .Z(n213) );
  MUX2_X1 U812 ( .A(n213), .B(n198), .S(N14), .Z(N16) );
  MUX2_X1 U813 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n618), .Z(n214) );
  MUX2_X1 U814 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n618), .Z(n215) );
  MUX2_X1 U815 ( .A(n215), .B(n214), .S(n613), .Z(n216) );
  MUX2_X1 U816 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n618), .Z(n217) );
  MUX2_X1 U817 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n618), .Z(n218) );
  MUX2_X1 U818 ( .A(n218), .B(n217), .S(n613), .Z(n219) );
  MUX2_X1 U819 ( .A(n219), .B(n216), .S(n609), .Z(n220) );
  MUX2_X1 U820 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n619), .Z(n221) );
  MUX2_X1 U821 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n615), .Z(n222) );
  MUX2_X1 U822 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U823 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n618), .Z(n224) );
  MUX2_X1 U824 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n617), .Z(n225) );
  MUX2_X1 U825 ( .A(n225), .B(n224), .S(n613), .Z(n226) );
  MUX2_X1 U826 ( .A(n226), .B(n223), .S(n609), .Z(n227) );
  MUX2_X1 U827 ( .A(n227), .B(n220), .S(N13), .Z(n228) );
  MUX2_X1 U828 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n619), .Z(n229) );
  MUX2_X1 U829 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n617), .Z(n595) );
  MUX2_X1 U830 ( .A(n595), .B(n229), .S(n611), .Z(n596) );
  MUX2_X1 U831 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n618), .Z(n597) );
  MUX2_X1 U832 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n617), .Z(n598) );
  MUX2_X1 U833 ( .A(n598), .B(n597), .S(N11), .Z(n599) );
  MUX2_X1 U834 ( .A(n599), .B(n596), .S(n610), .Z(n600) );
  MUX2_X1 U835 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n617), .Z(n601) );
  MUX2_X1 U836 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n615), .Z(n602) );
  MUX2_X1 U837 ( .A(n602), .B(n601), .S(n611), .Z(n603) );
  MUX2_X1 U838 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n618), .Z(n604) );
  MUX2_X1 U839 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n615), .Z(n605) );
  MUX2_X1 U840 ( .A(n605), .B(n604), .S(n613), .Z(n606) );
  MUX2_X1 U841 ( .A(n606), .B(n603), .S(n610), .Z(n607) );
  MUX2_X1 U842 ( .A(n607), .B(n600), .S(N13), .Z(n608) );
  MUX2_X1 U843 ( .A(n608), .B(n228), .S(N14), .Z(N15) );
  INV_X1 U844 ( .A(N10), .ZN(n620) );
  INV_X1 U845 ( .A(N11), .ZN(n621) );
  INV_X1 U846 ( .A(data_in[0]), .ZN(n622) );
  INV_X1 U847 ( .A(data_in[1]), .ZN(n623) );
  INV_X1 U848 ( .A(data_in[2]), .ZN(n624) );
  INV_X1 U849 ( .A(data_in[3]), .ZN(n625) );
  INV_X1 U850 ( .A(data_in[4]), .ZN(n626) );
  INV_X1 U851 ( .A(data_in[5]), .ZN(n627) );
  INV_X1 U852 ( .A(data_in[6]), .ZN(n628) );
  INV_X1 U853 ( .A(data_in[7]), .ZN(n629) );
endmodule


module mac_31_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70;
  wire   [15:1] carry;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKBUF_X1 U1 ( .A(carry[12]), .Z(n1) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n70) );
  XOR2_X1 U3 ( .A(B[15]), .B(A[15]), .Z(n2) );
  XOR2_X1 U4 ( .A(carry[15]), .B(n2), .Z(SUM[15]) );
  XOR2_X1 U5 ( .A(B[3]), .B(A[3]), .Z(n3) );
  XOR2_X1 U6 ( .A(carry[3]), .B(n3), .Z(SUM[3]) );
  NAND2_X1 U7 ( .A1(carry[3]), .A2(B[3]), .ZN(n4) );
  NAND2_X1 U8 ( .A1(carry[3]), .A2(A[3]), .ZN(n5) );
  NAND2_X1 U9 ( .A1(B[3]), .A2(A[3]), .ZN(n6) );
  NAND3_X1 U10 ( .A1(n4), .A2(n5), .A3(n6), .ZN(carry[4]) );
  NAND2_X1 U11 ( .A1(n20), .A2(B[9]), .ZN(n7) );
  CLKBUF_X1 U12 ( .A(n7), .Z(n8) );
  CLKBUF_X1 U13 ( .A(n45), .Z(n9) );
  XOR2_X1 U14 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR2_X1 U15 ( .A(carry[5]), .B(n10), .Z(SUM[5]) );
  NAND2_X1 U16 ( .A1(carry[5]), .A2(B[5]), .ZN(n11) );
  NAND2_X1 U17 ( .A1(carry[5]), .A2(A[5]), .ZN(n12) );
  NAND2_X1 U18 ( .A1(B[5]), .A2(A[5]), .ZN(n13) );
  NAND3_X1 U19 ( .A1(n11), .A2(n12), .A3(n13), .ZN(carry[6]) );
  XOR2_X1 U20 ( .A(B[11]), .B(A[11]), .Z(n14) );
  XOR2_X1 U21 ( .A(carry[11]), .B(n14), .Z(SUM[11]) );
  NAND2_X1 U22 ( .A1(carry[11]), .A2(B[11]), .ZN(n15) );
  NAND2_X1 U23 ( .A1(carry[11]), .A2(A[11]), .ZN(n16) );
  NAND2_X1 U24 ( .A1(B[11]), .A2(A[11]), .ZN(n17) );
  NAND3_X1 U25 ( .A1(n15), .A2(n16), .A3(n17), .ZN(carry[12]) );
  NAND3_X1 U26 ( .A1(n23), .A2(n22), .A3(n24), .ZN(n18) );
  NAND3_X1 U27 ( .A1(n40), .A2(n41), .A3(n42), .ZN(n19) );
  NAND3_X1 U28 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n20) );
  XOR2_X1 U29 ( .A(B[6]), .B(A[6]), .Z(n21) );
  XOR2_X1 U30 ( .A(carry[6]), .B(n21), .Z(SUM[6]) );
  NAND2_X1 U31 ( .A1(carry[6]), .A2(B[6]), .ZN(n22) );
  NAND2_X1 U32 ( .A1(carry[6]), .A2(A[6]), .ZN(n23) );
  NAND2_X1 U33 ( .A1(B[6]), .A2(A[6]), .ZN(n24) );
  NAND3_X1 U34 ( .A1(n22), .A2(n23), .A3(n24), .ZN(carry[7]) );
  NAND3_X1 U35 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n25) );
  XOR2_X1 U36 ( .A(B[12]), .B(A[12]), .Z(n26) );
  XOR2_X1 U37 ( .A(n1), .B(n26), .Z(SUM[12]) );
  NAND2_X1 U38 ( .A1(carry[12]), .A2(B[12]), .ZN(n27) );
  NAND2_X1 U39 ( .A1(carry[12]), .A2(A[12]), .ZN(n28) );
  NAND2_X1 U40 ( .A1(B[12]), .A2(A[12]), .ZN(n29) );
  NAND3_X1 U41 ( .A1(n27), .A2(n28), .A3(n29), .ZN(carry[13]) );
  CLKBUF_X1 U42 ( .A(n19), .Z(n30) );
  NAND3_X1 U43 ( .A1(n44), .A2(n45), .A3(n46), .ZN(n31) );
  NAND3_X1 U44 ( .A1(n44), .A2(n9), .A3(n46), .ZN(n32) );
  NAND3_X1 U45 ( .A1(n7), .A2(n60), .A3(n61), .ZN(n33) );
  NAND3_X1 U46 ( .A1(n8), .A2(n60), .A3(n61), .ZN(n34) );
  XOR2_X1 U47 ( .A(B[10]), .B(A[10]), .Z(n35) );
  XOR2_X1 U48 ( .A(n34), .B(n35), .Z(SUM[10]) );
  NAND2_X1 U49 ( .A1(n33), .A2(B[10]), .ZN(n36) );
  NAND2_X1 U50 ( .A1(carry[10]), .A2(A[10]), .ZN(n37) );
  NAND2_X1 U51 ( .A1(B[10]), .A2(A[10]), .ZN(n38) );
  NAND3_X1 U52 ( .A1(n36), .A2(n37), .A3(n38), .ZN(carry[11]) );
  XOR2_X1 U53 ( .A(B[13]), .B(A[13]), .Z(n39) );
  XOR2_X1 U54 ( .A(carry[13]), .B(n39), .Z(SUM[13]) );
  NAND2_X1 U55 ( .A1(n25), .A2(B[13]), .ZN(n40) );
  NAND2_X1 U56 ( .A1(n25), .A2(A[13]), .ZN(n41) );
  NAND2_X1 U57 ( .A1(B[13]), .A2(A[13]), .ZN(n42) );
  NAND3_X1 U58 ( .A1(n40), .A2(n41), .A3(n42), .ZN(carry[14]) );
  XOR2_X1 U59 ( .A(B[7]), .B(A[7]), .Z(n43) );
  XOR2_X1 U60 ( .A(carry[7]), .B(n43), .Z(SUM[7]) );
  NAND2_X1 U61 ( .A1(n18), .A2(B[7]), .ZN(n44) );
  NAND2_X1 U62 ( .A1(carry[7]), .A2(A[7]), .ZN(n45) );
  NAND2_X1 U63 ( .A1(B[7]), .A2(A[7]), .ZN(n46) );
  NAND3_X1 U64 ( .A1(n45), .A2(n44), .A3(n46), .ZN(carry[8]) );
  NAND3_X1 U65 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n47) );
  NAND3_X1 U66 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n48) );
  XOR2_X1 U67 ( .A(B[14]), .B(A[14]), .Z(n49) );
  XOR2_X1 U68 ( .A(n30), .B(n49), .Z(SUM[14]) );
  NAND2_X1 U69 ( .A1(n19), .A2(B[14]), .ZN(n50) );
  NAND2_X1 U70 ( .A1(carry[14]), .A2(A[14]), .ZN(n51) );
  NAND2_X1 U71 ( .A1(B[14]), .A2(A[14]), .ZN(n52) );
  NAND3_X1 U72 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[15]) );
  CLKBUF_X1 U73 ( .A(n20), .Z(n53) );
  XOR2_X1 U74 ( .A(B[8]), .B(A[8]), .Z(n54) );
  XOR2_X1 U75 ( .A(n32), .B(n54), .Z(SUM[8]) );
  NAND2_X1 U76 ( .A1(n31), .A2(B[8]), .ZN(n55) );
  NAND2_X1 U77 ( .A1(carry[8]), .A2(A[8]), .ZN(n56) );
  NAND2_X1 U78 ( .A1(B[8]), .A2(A[8]), .ZN(n57) );
  NAND3_X1 U79 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[9]) );
  XOR2_X1 U80 ( .A(B[9]), .B(A[9]), .Z(n58) );
  XOR2_X1 U81 ( .A(n53), .B(n58), .Z(SUM[9]) );
  NAND2_X1 U82 ( .A1(n20), .A2(B[9]), .ZN(n59) );
  NAND2_X1 U83 ( .A1(carry[9]), .A2(A[9]), .ZN(n60) );
  NAND2_X1 U84 ( .A1(B[9]), .A2(A[9]), .ZN(n61) );
  NAND3_X1 U85 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[10]) );
  XOR2_X1 U86 ( .A(B[1]), .B(A[1]), .Z(n62) );
  XOR2_X1 U87 ( .A(n70), .B(n62), .Z(SUM[1]) );
  NAND2_X1 U88 ( .A1(n70), .A2(B[1]), .ZN(n63) );
  NAND2_X1 U89 ( .A1(n70), .A2(A[1]), .ZN(n64) );
  NAND2_X1 U90 ( .A1(B[1]), .A2(A[1]), .ZN(n65) );
  NAND3_X1 U91 ( .A1(n63), .A2(n64), .A3(n65), .ZN(carry[2]) );
  XOR2_X1 U92 ( .A(B[2]), .B(A[2]), .Z(n66) );
  XOR2_X1 U93 ( .A(n48), .B(n66), .Z(SUM[2]) );
  NAND2_X1 U94 ( .A1(n47), .A2(B[2]), .ZN(n67) );
  NAND2_X1 U95 ( .A1(carry[2]), .A2(A[2]), .ZN(n68) );
  NAND2_X1 U96 ( .A1(B[2]), .A2(A[2]), .ZN(n69) );
  NAND3_X1 U97 ( .A1(n67), .A2(n68), .A3(n69), .ZN(carry[3]) );
  XOR2_X1 U98 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_31_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n308), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n307), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n306), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n305), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n304), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  INV_X1 U157 ( .A(a[4]), .ZN(n232) );
  BUF_X1 U158 ( .A(n303), .Z(n293) );
  CLKBUF_X1 U159 ( .A(n56), .Z(n206) );
  AND2_X1 U160 ( .A1(n212), .A2(n102), .ZN(n207) );
  CLKBUF_X1 U161 ( .A(n300), .Z(n208) );
  NAND2_X1 U162 ( .A1(n245), .A2(n18), .ZN(n209) );
  CLKBUF_X1 U163 ( .A(n244), .Z(n210) );
  NAND3_X1 U164 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n211) );
  XOR2_X1 U165 ( .A(n95), .B(n102), .Z(n56) );
  OAI22_X1 U166 ( .A1(n322), .A2(n323), .B1(n252), .B2(n324), .ZN(n212) );
  XOR2_X1 U167 ( .A(n100), .B(n93), .Z(n213) );
  XOR2_X1 U168 ( .A(n52), .B(n213), .Z(n50) );
  NAND2_X1 U169 ( .A1(n52), .A2(n100), .ZN(n214) );
  NAND2_X1 U170 ( .A1(n52), .A2(n93), .ZN(n215) );
  NAND2_X1 U171 ( .A1(n100), .A2(n93), .ZN(n216) );
  NAND3_X1 U172 ( .A1(n214), .A2(n215), .A3(n216), .ZN(n49) );
  NAND3_X1 U173 ( .A1(n299), .A2(n300), .A3(n301), .ZN(n217) );
  NAND3_X1 U174 ( .A1(n299), .A2(n208), .A3(n301), .ZN(n218) );
  CLKBUF_X1 U175 ( .A(n211), .Z(n219) );
  INV_X1 U176 ( .A(n303), .ZN(n220) );
  INV_X1 U177 ( .A(n303), .ZN(n302) );
  CLKBUF_X1 U178 ( .A(n261), .Z(n221) );
  CLKBUF_X1 U179 ( .A(n238), .Z(n222) );
  NAND2_X1 U180 ( .A1(n17), .A2(n251), .ZN(n223) );
  CLKBUF_X1 U181 ( .A(n209), .Z(n224) );
  XOR2_X1 U182 ( .A(n46), .B(n49), .Z(n225) );
  XOR2_X1 U183 ( .A(n218), .B(n225), .Z(product[6]) );
  NAND2_X1 U184 ( .A1(n217), .A2(n46), .ZN(n226) );
  NAND2_X1 U185 ( .A1(n10), .A2(n49), .ZN(n227) );
  NAND2_X1 U186 ( .A1(n46), .A2(n49), .ZN(n228) );
  NAND3_X1 U187 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n9) );
  CLKBUF_X1 U188 ( .A(n289), .Z(n229) );
  NAND3_X1 U189 ( .A1(n209), .A2(n268), .A3(n269), .ZN(n230) );
  NAND3_X1 U190 ( .A1(n224), .A2(n268), .A3(n269), .ZN(n231) );
  NAND2_X1 U191 ( .A1(a[4]), .A2(a[3]), .ZN(n233) );
  NAND2_X1 U192 ( .A1(n232), .A2(n313), .ZN(n234) );
  NAND2_X2 U193 ( .A1(n233), .A2(n234), .ZN(n331) );
  CLKBUF_X1 U194 ( .A(n245), .Z(n235) );
  AND2_X1 U195 ( .A1(n104), .A2(n72), .ZN(n236) );
  NAND3_X1 U196 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n237) );
  NAND3_X1 U197 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n238) );
  NAND3_X1 U198 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n239) );
  XOR2_X1 U199 ( .A(n40), .B(n45), .Z(n240) );
  XOR2_X1 U200 ( .A(n219), .B(n240), .Z(product[7]) );
  NAND2_X1 U201 ( .A1(n211), .A2(n40), .ZN(n241) );
  NAND2_X1 U202 ( .A1(n9), .A2(n45), .ZN(n242) );
  NAND2_X1 U203 ( .A1(n40), .A2(n45), .ZN(n243) );
  NAND3_X1 U204 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n8) );
  NAND3_X1 U205 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n244) );
  NAND3_X1 U206 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n245) );
  CLKBUF_X1 U207 ( .A(n7), .Z(n246) );
  XOR2_X1 U208 ( .A(n23), .B(n20), .Z(n247) );
  XOR2_X1 U209 ( .A(n210), .B(n247), .Z(product[11]) );
  NAND2_X1 U210 ( .A1(n244), .A2(n23), .ZN(n248) );
  NAND2_X1 U211 ( .A1(n5), .A2(n20), .ZN(n249) );
  NAND2_X1 U212 ( .A1(n23), .A2(n20), .ZN(n250) );
  NAND3_X1 U213 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n4) );
  NAND3_X1 U214 ( .A1(n267), .A2(n268), .A3(n269), .ZN(n251) );
  XNOR2_X1 U215 ( .A(a[2]), .B(a[1]), .ZN(n252) );
  XNOR2_X1 U216 ( .A(a[2]), .B(a[1]), .ZN(n321) );
  XOR2_X1 U217 ( .A(n34), .B(n39), .Z(n253) );
  XOR2_X1 U218 ( .A(n239), .B(n253), .Z(product[8]) );
  NAND2_X1 U219 ( .A1(n8), .A2(n34), .ZN(n254) );
  NAND2_X1 U220 ( .A1(n8), .A2(n39), .ZN(n255) );
  NAND2_X1 U221 ( .A1(n34), .A2(n39), .ZN(n256) );
  NAND3_X1 U222 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n7) );
  XOR2_X1 U223 ( .A(n103), .B(n96), .Z(n257) );
  XOR2_X1 U224 ( .A(n236), .B(n257), .Z(product[2]) );
  NAND2_X1 U225 ( .A1(n236), .A2(n103), .ZN(n258) );
  NAND2_X1 U226 ( .A1(n14), .A2(n96), .ZN(n259) );
  NAND2_X1 U227 ( .A1(n103), .A2(n96), .ZN(n260) );
  NAND3_X1 U228 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n13) );
  NAND3_X1 U229 ( .A1(n264), .A2(n263), .A3(n265), .ZN(n261) );
  NAND2_X2 U230 ( .A1(n331), .A2(n360), .ZN(n333) );
  XOR2_X1 U231 ( .A(n33), .B(n28), .Z(n262) );
  XOR2_X1 U232 ( .A(n246), .B(n262), .Z(product[9]) );
  NAND2_X1 U233 ( .A1(n237), .A2(n33), .ZN(n263) );
  NAND2_X1 U234 ( .A1(n7), .A2(n28), .ZN(n264) );
  NAND2_X1 U235 ( .A1(n33), .A2(n28), .ZN(n265) );
  NAND3_X1 U236 ( .A1(n264), .A2(n263), .A3(n265), .ZN(n6) );
  XOR2_X1 U237 ( .A(n18), .B(n19), .Z(n266) );
  XOR2_X1 U238 ( .A(n235), .B(n266), .Z(product[12]) );
  NAND2_X1 U239 ( .A1(n245), .A2(n18), .ZN(n267) );
  NAND2_X1 U240 ( .A1(n4), .A2(n19), .ZN(n268) );
  NAND2_X1 U241 ( .A1(n18), .A2(n19), .ZN(n269) );
  XOR2_X1 U242 ( .A(n27), .B(n24), .Z(n270) );
  XOR2_X1 U243 ( .A(n221), .B(n270), .Z(product[10]) );
  NAND2_X1 U244 ( .A1(n261), .A2(n27), .ZN(n271) );
  NAND2_X1 U245 ( .A1(n6), .A2(n24), .ZN(n272) );
  NAND2_X1 U246 ( .A1(n27), .A2(n24), .ZN(n273) );
  NAND3_X1 U247 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n5) );
  XNOR2_X1 U248 ( .A(n274), .B(n280), .ZN(product[14]) );
  XNOR2_X1 U249 ( .A(n310), .B(n15), .ZN(n274) );
  AND3_X1 U250 ( .A1(n287), .A2(n286), .A3(n285), .ZN(product[15]) );
  NAND3_X1 U251 ( .A1(n295), .A2(n296), .A3(n297), .ZN(n276) );
  NAND3_X1 U252 ( .A1(n289), .A2(n290), .A3(n291), .ZN(n277) );
  NAND3_X1 U253 ( .A1(n229), .A2(n290), .A3(n291), .ZN(n278) );
  NAND3_X1 U254 ( .A1(n284), .A2(n283), .A3(n282), .ZN(n279) );
  NAND3_X1 U255 ( .A1(n284), .A2(n223), .A3(n282), .ZN(n280) );
  XOR2_X1 U256 ( .A(n17), .B(n309), .Z(n281) );
  XOR2_X1 U257 ( .A(n281), .B(n231), .Z(product[13]) );
  NAND2_X1 U258 ( .A1(n17), .A2(n309), .ZN(n282) );
  NAND2_X1 U259 ( .A1(n17), .A2(n251), .ZN(n283) );
  NAND2_X1 U260 ( .A1(n230), .A2(n309), .ZN(n284) );
  NAND3_X1 U261 ( .A1(n223), .A2(n282), .A3(n284), .ZN(n2) );
  NAND2_X1 U262 ( .A1(n310), .A2(n15), .ZN(n285) );
  NAND2_X1 U263 ( .A1(n2), .A2(n310), .ZN(n286) );
  NAND2_X1 U264 ( .A1(n15), .A2(n279), .ZN(n287) );
  XOR2_X1 U265 ( .A(n206), .B(n71), .Z(n288) );
  XOR2_X1 U266 ( .A(n222), .B(n288), .Z(product[3]) );
  NAND2_X1 U267 ( .A1(n238), .A2(n56), .ZN(n289) );
  NAND2_X1 U268 ( .A1(n13), .A2(n71), .ZN(n290) );
  NAND2_X1 U269 ( .A1(n56), .A2(n71), .ZN(n291) );
  NAND3_X1 U270 ( .A1(n289), .A2(n290), .A3(n291), .ZN(n12) );
  CLKBUF_X1 U271 ( .A(n11), .Z(n292) );
  INV_X1 U272 ( .A(n15), .ZN(n309) );
  INV_X1 U273 ( .A(n21), .ZN(n307) );
  INV_X1 U274 ( .A(n340), .ZN(n308) );
  INV_X1 U275 ( .A(n320), .ZN(n304) );
  INV_X1 U276 ( .A(n329), .ZN(n306) );
  INV_X1 U277 ( .A(n351), .ZN(n310) );
  INV_X1 U278 ( .A(n31), .ZN(n305) );
  INV_X1 U279 ( .A(a[0]), .ZN(n315) );
  INV_X1 U280 ( .A(a[5]), .ZN(n312) );
  INV_X1 U281 ( .A(a[7]), .ZN(n311) );
  INV_X1 U282 ( .A(b[0]), .ZN(n303) );
  XOR2_X1 U283 ( .A(n54), .B(n207), .Z(n294) );
  XOR2_X1 U284 ( .A(n278), .B(n294), .Z(product[4]) );
  NAND2_X1 U285 ( .A1(n277), .A2(n54), .ZN(n295) );
  NAND2_X1 U286 ( .A1(n12), .A2(n207), .ZN(n296) );
  NAND2_X1 U287 ( .A1(n54), .A2(n207), .ZN(n297) );
  NAND3_X1 U288 ( .A1(n295), .A2(n296), .A3(n297), .ZN(n11) );
  XOR2_X1 U289 ( .A(n50), .B(n53), .Z(n298) );
  XOR2_X1 U290 ( .A(n292), .B(n298), .Z(product[5]) );
  NAND2_X1 U291 ( .A1(n276), .A2(n50), .ZN(n299) );
  NAND2_X1 U292 ( .A1(n11), .A2(n53), .ZN(n300) );
  NAND2_X1 U293 ( .A1(n50), .A2(n53), .ZN(n301) );
  NAND3_X1 U294 ( .A1(n299), .A2(n300), .A3(n301), .ZN(n10) );
  INV_X1 U295 ( .A(a[3]), .ZN(n313) );
  INV_X1 U296 ( .A(a[1]), .ZN(n314) );
  NAND2_X2 U297 ( .A1(n321), .A2(n359), .ZN(n323) );
  XOR2_X2 U298 ( .A(a[6]), .B(n312), .Z(n342) );
  NOR2_X1 U299 ( .A1(n315), .A2(n293), .ZN(product[0]) );
  OAI22_X1 U300 ( .A1(n316), .A2(n317), .B1(n318), .B2(n315), .ZN(n99) );
  OAI22_X1 U301 ( .A1(n318), .A2(n317), .B1(n319), .B2(n315), .ZN(n98) );
  XNOR2_X1 U302 ( .A(b[6]), .B(a[1]), .ZN(n318) );
  OAI22_X1 U303 ( .A1(n315), .A2(n319), .B1(n317), .B2(n319), .ZN(n320) );
  XNOR2_X1 U304 ( .A(b[7]), .B(a[1]), .ZN(n319) );
  NOR2_X1 U305 ( .A1(n252), .A2(n293), .ZN(n96) );
  OAI22_X1 U306 ( .A1(n322), .A2(n323), .B1(n252), .B2(n324), .ZN(n95) );
  XNOR2_X1 U307 ( .A(a[3]), .B(n302), .ZN(n322) );
  OAI22_X1 U308 ( .A1(n324), .A2(n323), .B1(n252), .B2(n325), .ZN(n94) );
  XNOR2_X1 U309 ( .A(b[1]), .B(a[3]), .ZN(n324) );
  OAI22_X1 U310 ( .A1(n325), .A2(n323), .B1(n252), .B2(n326), .ZN(n93) );
  XNOR2_X1 U311 ( .A(b[2]), .B(a[3]), .ZN(n325) );
  OAI22_X1 U312 ( .A1(n326), .A2(n323), .B1(n252), .B2(n327), .ZN(n92) );
  XNOR2_X1 U313 ( .A(b[3]), .B(a[3]), .ZN(n326) );
  OAI22_X1 U314 ( .A1(n327), .A2(n323), .B1(n252), .B2(n328), .ZN(n91) );
  XNOR2_X1 U315 ( .A(b[4]), .B(a[3]), .ZN(n327) );
  OAI22_X1 U316 ( .A1(n330), .A2(n252), .B1(n323), .B2(n330), .ZN(n329) );
  NOR2_X1 U317 ( .A1(n331), .A2(n293), .ZN(n88) );
  OAI22_X1 U318 ( .A1(n332), .A2(n333), .B1(n331), .B2(n334), .ZN(n87) );
  XNOR2_X1 U319 ( .A(a[5]), .B(n220), .ZN(n332) );
  OAI22_X1 U320 ( .A1(n334), .A2(n333), .B1(n331), .B2(n335), .ZN(n86) );
  XNOR2_X1 U321 ( .A(b[1]), .B(a[5]), .ZN(n334) );
  OAI22_X1 U322 ( .A1(n335), .A2(n333), .B1(n331), .B2(n336), .ZN(n85) );
  XNOR2_X1 U323 ( .A(b[2]), .B(a[5]), .ZN(n335) );
  OAI22_X1 U324 ( .A1(n336), .A2(n333), .B1(n331), .B2(n337), .ZN(n84) );
  XNOR2_X1 U325 ( .A(b[3]), .B(a[5]), .ZN(n336) );
  OAI22_X1 U326 ( .A1(n337), .A2(n333), .B1(n331), .B2(n338), .ZN(n83) );
  XNOR2_X1 U327 ( .A(b[4]), .B(a[5]), .ZN(n337) );
  OAI22_X1 U328 ( .A1(n338), .A2(n333), .B1(n331), .B2(n339), .ZN(n82) );
  XNOR2_X1 U329 ( .A(b[5]), .B(a[5]), .ZN(n338) );
  OAI22_X1 U330 ( .A1(n341), .A2(n331), .B1(n333), .B2(n341), .ZN(n340) );
  NOR2_X1 U331 ( .A1(n342), .A2(n293), .ZN(n80) );
  OAI22_X1 U332 ( .A1(n343), .A2(n344), .B1(n342), .B2(n345), .ZN(n79) );
  XNOR2_X1 U333 ( .A(a[7]), .B(n220), .ZN(n343) );
  OAI22_X1 U334 ( .A1(n346), .A2(n344), .B1(n342), .B2(n347), .ZN(n77) );
  OAI22_X1 U335 ( .A1(n347), .A2(n344), .B1(n342), .B2(n348), .ZN(n76) );
  XNOR2_X1 U336 ( .A(b[3]), .B(a[7]), .ZN(n347) );
  OAI22_X1 U337 ( .A1(n348), .A2(n344), .B1(n342), .B2(n349), .ZN(n75) );
  XNOR2_X1 U338 ( .A(b[4]), .B(a[7]), .ZN(n348) );
  OAI22_X1 U339 ( .A1(n349), .A2(n344), .B1(n342), .B2(n350), .ZN(n74) );
  XNOR2_X1 U340 ( .A(b[5]), .B(a[7]), .ZN(n349) );
  OAI22_X1 U341 ( .A1(n352), .A2(n342), .B1(n344), .B2(n352), .ZN(n351) );
  OAI21_X1 U342 ( .B1(n220), .B2(n314), .A(n317), .ZN(n72) );
  OAI21_X1 U343 ( .B1(n313), .B2(n323), .A(n353), .ZN(n71) );
  OR3_X1 U344 ( .A1(n252), .A2(n220), .A3(n313), .ZN(n353) );
  OAI21_X1 U345 ( .B1(n312), .B2(n333), .A(n354), .ZN(n70) );
  OR3_X1 U346 ( .A1(n331), .A2(n302), .A3(n312), .ZN(n354) );
  OAI21_X1 U347 ( .B1(n311), .B2(n344), .A(n355), .ZN(n69) );
  OR3_X1 U348 ( .A1(n342), .A2(n220), .A3(n311), .ZN(n355) );
  XNOR2_X1 U349 ( .A(n356), .B(n357), .ZN(n38) );
  OR2_X1 U350 ( .A1(n356), .A2(n357), .ZN(n37) );
  OAI22_X1 U351 ( .A1(n328), .A2(n323), .B1(n252), .B2(n358), .ZN(n357) );
  XNOR2_X1 U352 ( .A(b[5]), .B(a[3]), .ZN(n328) );
  OAI22_X1 U353 ( .A1(n345), .A2(n344), .B1(n342), .B2(n346), .ZN(n356) );
  XNOR2_X1 U354 ( .A(b[2]), .B(a[7]), .ZN(n346) );
  XNOR2_X1 U355 ( .A(b[1]), .B(a[7]), .ZN(n345) );
  OAI22_X1 U356 ( .A1(n358), .A2(n323), .B1(n252), .B2(n330), .ZN(n31) );
  XNOR2_X1 U357 ( .A(b[7]), .B(a[3]), .ZN(n330) );
  XNOR2_X1 U358 ( .A(n313), .B(a[2]), .ZN(n359) );
  XNOR2_X1 U359 ( .A(b[6]), .B(a[3]), .ZN(n358) );
  OAI22_X1 U360 ( .A1(n339), .A2(n333), .B1(n331), .B2(n341), .ZN(n21) );
  XNOR2_X1 U361 ( .A(b[7]), .B(a[5]), .ZN(n341) );
  XNOR2_X1 U362 ( .A(n312), .B(a[4]), .ZN(n360) );
  XNOR2_X1 U363 ( .A(b[6]), .B(a[5]), .ZN(n339) );
  OAI22_X1 U364 ( .A1(n350), .A2(n344), .B1(n342), .B2(n352), .ZN(n15) );
  XNOR2_X1 U365 ( .A(b[7]), .B(a[7]), .ZN(n352) );
  NAND2_X1 U366 ( .A1(n342), .A2(n361), .ZN(n344) );
  XNOR2_X1 U367 ( .A(n311), .B(a[6]), .ZN(n361) );
  XNOR2_X1 U368 ( .A(b[6]), .B(a[7]), .ZN(n350) );
  OAI22_X1 U369 ( .A1(n220), .A2(n317), .B1(n362), .B2(n315), .ZN(n104) );
  OAI22_X1 U370 ( .A1(n362), .A2(n317), .B1(n363), .B2(n315), .ZN(n103) );
  XNOR2_X1 U371 ( .A(b[1]), .B(a[1]), .ZN(n362) );
  OAI22_X1 U372 ( .A1(n363), .A2(n317), .B1(n364), .B2(n315), .ZN(n102) );
  XNOR2_X1 U373 ( .A(b[2]), .B(a[1]), .ZN(n363) );
  OAI22_X1 U374 ( .A1(n364), .A2(n317), .B1(n365), .B2(n315), .ZN(n101) );
  XNOR2_X1 U375 ( .A(b[3]), .B(a[1]), .ZN(n364) );
  OAI22_X1 U376 ( .A1(n365), .A2(n317), .B1(n316), .B2(n315), .ZN(n100) );
  XNOR2_X1 U377 ( .A(b[5]), .B(a[1]), .ZN(n316) );
  NAND2_X1 U378 ( .A1(a[1]), .A2(n315), .ZN(n317) );
  XNOR2_X1 U379 ( .A(b[4]), .B(a[1]), .ZN(n365) );
endmodule


module mac_31 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_31_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_31_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_30_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61;
  wire   [15:1] carry;

  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CLKBUF_X1 U1 ( .A(carry[13]), .Z(n1) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n61) );
  XNOR2_X1 U3 ( .A(B[15]), .B(A[15]), .ZN(n2) );
  XOR2_X1 U4 ( .A(B[11]), .B(A[11]), .Z(n3) );
  XOR2_X1 U5 ( .A(carry[11]), .B(n3), .Z(SUM[11]) );
  NAND2_X1 U6 ( .A1(carry[11]), .A2(B[11]), .ZN(n4) );
  NAND2_X1 U7 ( .A1(carry[11]), .A2(A[11]), .ZN(n5) );
  NAND2_X1 U8 ( .A1(B[11]), .A2(A[11]), .ZN(n6) );
  NAND3_X1 U9 ( .A1(n4), .A2(n5), .A3(n6), .ZN(carry[12]) );
  NAND3_X1 U10 ( .A1(n35), .A2(n36), .A3(n37), .ZN(n7) );
  CLKBUF_X1 U11 ( .A(n26), .Z(n8) );
  CLKBUF_X1 U12 ( .A(A[0]), .Z(n9) );
  XOR2_X1 U13 ( .A(B[10]), .B(A[10]), .Z(n10) );
  XOR2_X1 U14 ( .A(carry[10]), .B(n10), .Z(SUM[10]) );
  NAND2_X1 U15 ( .A1(carry[10]), .A2(B[10]), .ZN(n11) );
  NAND2_X1 U16 ( .A1(carry[10]), .A2(A[10]), .ZN(n12) );
  NAND2_X1 U17 ( .A1(B[10]), .A2(A[10]), .ZN(n13) );
  NAND3_X1 U18 ( .A1(n11), .A2(n12), .A3(n13), .ZN(carry[11]) );
  CLKBUF_X1 U19 ( .A(n32), .Z(n14) );
  CLKBUF_X1 U20 ( .A(carry[6]), .Z(n15) );
  CLKBUF_X1 U21 ( .A(carry[12]), .Z(n16) );
  XNOR2_X1 U22 ( .A(carry[15]), .B(n2), .ZN(SUM[15]) );
  NAND3_X1 U23 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n17) );
  NAND3_X1 U24 ( .A1(n25), .A2(n8), .A3(n27), .ZN(n18) );
  NAND3_X1 U25 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n19) );
  XOR2_X1 U26 ( .A(B[12]), .B(A[12]), .Z(n20) );
  XOR2_X1 U27 ( .A(n16), .B(n20), .Z(SUM[12]) );
  NAND2_X1 U28 ( .A1(carry[12]), .A2(B[12]), .ZN(n21) );
  NAND2_X1 U29 ( .A1(carry[12]), .A2(A[12]), .ZN(n22) );
  NAND2_X1 U30 ( .A1(B[12]), .A2(A[12]), .ZN(n23) );
  NAND3_X1 U31 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[13]) );
  XOR2_X1 U32 ( .A(B[6]), .B(A[6]), .Z(n24) );
  XOR2_X1 U33 ( .A(n15), .B(n24), .Z(SUM[6]) );
  NAND2_X1 U34 ( .A1(carry[6]), .A2(B[6]), .ZN(n25) );
  NAND2_X1 U35 ( .A1(carry[6]), .A2(A[6]), .ZN(n26) );
  NAND2_X1 U36 ( .A1(B[6]), .A2(A[6]), .ZN(n27) );
  NAND3_X1 U37 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[7]) );
  NAND3_X1 U38 ( .A1(n31), .A2(n14), .A3(n33), .ZN(n28) );
  NAND3_X1 U39 ( .A1(n35), .A2(n36), .A3(n37), .ZN(n29) );
  XOR2_X1 U40 ( .A(B[13]), .B(A[13]), .Z(n30) );
  XOR2_X1 U41 ( .A(n1), .B(n30), .Z(SUM[13]) );
  NAND2_X1 U42 ( .A1(carry[13]), .A2(B[13]), .ZN(n31) );
  NAND2_X1 U43 ( .A1(carry[13]), .A2(A[13]), .ZN(n32) );
  NAND2_X1 U44 ( .A1(B[13]), .A2(A[13]), .ZN(n33) );
  NAND3_X1 U45 ( .A1(n31), .A2(n32), .A3(n33), .ZN(carry[14]) );
  XOR2_X1 U46 ( .A(B[7]), .B(A[7]), .Z(n34) );
  XOR2_X1 U47 ( .A(n18), .B(n34), .Z(SUM[7]) );
  NAND2_X1 U48 ( .A1(n17), .A2(B[7]), .ZN(n35) );
  NAND2_X1 U49 ( .A1(carry[7]), .A2(A[7]), .ZN(n36) );
  NAND2_X1 U50 ( .A1(B[7]), .A2(A[7]), .ZN(n37) );
  NAND3_X1 U51 ( .A1(n35), .A2(n36), .A3(n37), .ZN(carry[8]) );
  NAND3_X1 U52 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n38) );
  NAND3_X1 U53 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n39) );
  XOR2_X1 U54 ( .A(B[14]), .B(A[14]), .Z(n40) );
  XOR2_X1 U55 ( .A(n28), .B(n40), .Z(SUM[14]) );
  NAND2_X1 U56 ( .A1(carry[14]), .A2(B[14]), .ZN(n41) );
  NAND2_X1 U57 ( .A1(carry[14]), .A2(A[14]), .ZN(n42) );
  NAND2_X1 U58 ( .A1(B[14]), .A2(A[14]), .ZN(n43) );
  NAND3_X1 U59 ( .A1(n41), .A2(n42), .A3(n43), .ZN(carry[15]) );
  CLKBUF_X1 U60 ( .A(n19), .Z(n44) );
  XOR2_X1 U61 ( .A(B[8]), .B(A[8]), .Z(n45) );
  XOR2_X1 U62 ( .A(n7), .B(n45), .Z(SUM[8]) );
  NAND2_X1 U63 ( .A1(carry[8]), .A2(B[8]), .ZN(n46) );
  NAND2_X1 U64 ( .A1(n29), .A2(A[8]), .ZN(n47) );
  NAND2_X1 U65 ( .A1(B[8]), .A2(A[8]), .ZN(n48) );
  NAND3_X1 U66 ( .A1(n47), .A2(n46), .A3(n48), .ZN(carry[9]) );
  XOR2_X1 U67 ( .A(B[9]), .B(A[9]), .Z(n49) );
  XOR2_X1 U68 ( .A(n44), .B(n49), .Z(SUM[9]) );
  NAND2_X1 U69 ( .A1(n19), .A2(B[9]), .ZN(n50) );
  NAND2_X1 U70 ( .A1(carry[9]), .A2(A[9]), .ZN(n51) );
  NAND2_X1 U71 ( .A1(B[9]), .A2(A[9]), .ZN(n52) );
  NAND3_X1 U72 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[10]) );
  XOR2_X1 U73 ( .A(B[1]), .B(A[1]), .Z(n53) );
  XOR2_X1 U74 ( .A(n61), .B(n53), .Z(SUM[1]) );
  NAND2_X1 U75 ( .A1(n61), .A2(B[1]), .ZN(n54) );
  NAND2_X1 U76 ( .A1(n61), .A2(A[1]), .ZN(n55) );
  NAND2_X1 U77 ( .A1(B[1]), .A2(A[1]), .ZN(n56) );
  NAND3_X1 U78 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[2]) );
  XOR2_X1 U79 ( .A(B[2]), .B(A[2]), .Z(n57) );
  XOR2_X1 U80 ( .A(n39), .B(n57), .Z(SUM[2]) );
  NAND2_X1 U81 ( .A1(n38), .A2(B[2]), .ZN(n58) );
  NAND2_X1 U82 ( .A1(carry[2]), .A2(A[2]), .ZN(n59) );
  NAND2_X1 U83 ( .A1(B[2]), .A2(A[2]), .ZN(n60) );
  NAND3_X1 U84 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[3]) );
  XOR2_X1 U85 ( .A(B[0]), .B(n9), .Z(SUM[0]) );
endmodule


module mac_30_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n304), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n303), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n307), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n306), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n309), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n94), .B(n88), .CI(n101), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n102), .B(n95), .CO(n55), .S(n56) );
  NAND2_X1 U157 ( .A1(n317), .A2(n355), .ZN(n319) );
  NAND2_X1 U158 ( .A1(n327), .A2(n356), .ZN(n329) );
  CLKBUF_X1 U159 ( .A(n228), .Z(n206) );
  NAND2_X1 U160 ( .A1(n221), .A2(n46), .ZN(n207) );
  CLKBUF_X1 U161 ( .A(n207), .Z(n208) );
  INV_X1 U162 ( .A(a[5]), .ZN(n209) );
  CLKBUF_X1 U163 ( .A(n358), .Z(n210) );
  NAND2_X1 U164 ( .A1(n225), .A2(n34), .ZN(n211) );
  CLKBUF_X1 U165 ( .A(n3), .Z(n212) );
  CLKBUF_X1 U166 ( .A(n246), .Z(n213) );
  NAND3_X1 U167 ( .A1(n207), .A2(n249), .A3(n250), .ZN(n214) );
  NAND3_X1 U168 ( .A1(n208), .A2(n249), .A3(n250), .ZN(n215) );
  NAND3_X1 U169 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n216) );
  NAND3_X1 U170 ( .A1(n227), .A2(n206), .A3(n229), .ZN(n217) );
  XOR2_X1 U171 ( .A(a[3]), .B(a[2]), .Z(n355) );
  CLKBUF_X1 U172 ( .A(n286), .Z(n218) );
  CLKBUF_X1 U173 ( .A(n285), .Z(n219) );
  CLKBUF_X1 U174 ( .A(n56), .Z(n220) );
  XOR2_X2 U175 ( .A(a[6]), .B(n305), .Z(n338) );
  NAND3_X1 U176 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n221) );
  NAND3_X1 U177 ( .A1(n287), .A2(n286), .A3(n285), .ZN(n222) );
  NAND3_X1 U178 ( .A1(n287), .A2(n218), .A3(n219), .ZN(n223) );
  CLKBUF_X1 U179 ( .A(n221), .Z(n224) );
  NAND3_X1 U180 ( .A1(n239), .A2(n238), .A3(n240), .ZN(n225) );
  XOR2_X1 U181 ( .A(n54), .B(n55), .Z(n226) );
  XOR2_X1 U182 ( .A(n223), .B(n226), .Z(product[4]) );
  NAND2_X1 U183 ( .A1(n222), .A2(n54), .ZN(n227) );
  NAND2_X1 U184 ( .A1(n12), .A2(n55), .ZN(n228) );
  NAND2_X1 U185 ( .A1(n54), .A2(n55), .ZN(n229) );
  NAND3_X1 U186 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n11) );
  CLKBUF_X1 U187 ( .A(n225), .Z(n230) );
  NAND2_X1 U188 ( .A1(n14), .A2(n96), .ZN(n231) );
  AND2_X1 U189 ( .A1(n104), .A2(n72), .ZN(n232) );
  XOR2_X1 U190 ( .A(n50), .B(n53), .Z(n233) );
  XOR2_X1 U191 ( .A(n217), .B(n233), .Z(product[5]) );
  NAND2_X1 U192 ( .A1(n11), .A2(n50), .ZN(n234) );
  NAND2_X1 U193 ( .A1(n216), .A2(n53), .ZN(n235) );
  NAND2_X1 U194 ( .A1(n50), .A2(n53), .ZN(n236) );
  NAND3_X1 U195 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n10) );
  XNOR2_X1 U196 ( .A(a[2]), .B(a[1]), .ZN(n317) );
  XOR2_X1 U197 ( .A(n40), .B(n45), .Z(n237) );
  XOR2_X1 U198 ( .A(n215), .B(n237), .Z(product[7]) );
  NAND2_X1 U199 ( .A1(n9), .A2(n40), .ZN(n238) );
  NAND2_X1 U200 ( .A1(n214), .A2(n45), .ZN(n239) );
  NAND2_X1 U201 ( .A1(n40), .A2(n45), .ZN(n240) );
  NAND3_X1 U202 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n8) );
  XNOR2_X1 U203 ( .A(a[4]), .B(a[3]), .ZN(n241) );
  XNOR2_X1 U204 ( .A(a[4]), .B(a[3]), .ZN(n242) );
  XNOR2_X1 U205 ( .A(a[4]), .B(a[3]), .ZN(n327) );
  NAND3_X1 U206 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n243) );
  NAND3_X1 U207 ( .A1(n211), .A2(n261), .A3(n262), .ZN(n244) );
  NAND3_X1 U208 ( .A1(n211), .A2(n261), .A3(n262), .ZN(n245) );
  NAND3_X1 U209 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n246) );
  XOR2_X1 U210 ( .A(n46), .B(n49), .Z(n247) );
  XOR2_X1 U211 ( .A(n224), .B(n247), .Z(product[6]) );
  NAND2_X1 U212 ( .A1(n221), .A2(n46), .ZN(n248) );
  NAND2_X1 U213 ( .A1(n10), .A2(n49), .ZN(n249) );
  NAND2_X1 U214 ( .A1(n46), .A2(n49), .ZN(n250) );
  NAND3_X1 U215 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n9) );
  CLKBUF_X1 U216 ( .A(n274), .Z(n251) );
  CLKBUF_X1 U217 ( .A(n243), .Z(n252) );
  INV_X1 U218 ( .A(b[0]), .ZN(n253) );
  XOR2_X1 U219 ( .A(n33), .B(n28), .Z(n254) );
  XOR2_X1 U220 ( .A(n245), .B(n254), .Z(product[9]) );
  NAND2_X1 U221 ( .A1(n244), .A2(n33), .ZN(n255) );
  NAND2_X1 U222 ( .A1(n7), .A2(n28), .ZN(n256) );
  NAND2_X1 U223 ( .A1(n33), .A2(n28), .ZN(n257) );
  NAND3_X1 U224 ( .A1(n256), .A2(n255), .A3(n257), .ZN(n6) );
  XNOR2_X1 U225 ( .A(n258), .B(n2), .ZN(product[14]) );
  XNOR2_X1 U226 ( .A(n301), .B(n15), .ZN(n258) );
  XOR2_X1 U227 ( .A(n34), .B(n39), .Z(n259) );
  XOR2_X1 U228 ( .A(n230), .B(n259), .Z(product[8]) );
  NAND2_X1 U229 ( .A1(n225), .A2(n34), .ZN(n260) );
  NAND2_X1 U230 ( .A1(n8), .A2(n39), .ZN(n261) );
  NAND2_X1 U231 ( .A1(n34), .A2(n39), .ZN(n262) );
  NAND3_X1 U232 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n7) );
  XOR2_X1 U233 ( .A(n27), .B(n24), .Z(n263) );
  XOR2_X1 U234 ( .A(n252), .B(n263), .Z(product[10]) );
  NAND2_X1 U235 ( .A1(n243), .A2(n27), .ZN(n264) );
  NAND2_X1 U236 ( .A1(n6), .A2(n24), .ZN(n265) );
  NAND2_X1 U237 ( .A1(n27), .A2(n24), .ZN(n266) );
  NAND3_X1 U238 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n5) );
  NAND3_X1 U239 ( .A1(n282), .A2(n231), .A3(n281), .ZN(n267) );
  NAND3_X1 U240 ( .A1(n282), .A2(n231), .A3(n281), .ZN(n268) );
  NAND3_X1 U241 ( .A1(n274), .A2(n273), .A3(n275), .ZN(n269) );
  NAND3_X1 U242 ( .A1(n273), .A2(n251), .A3(n275), .ZN(n270) );
  NAND3_X1 U243 ( .A1(n278), .A2(n277), .A3(n279), .ZN(n271) );
  XOR2_X1 U244 ( .A(n20), .B(n23), .Z(n272) );
  XOR2_X1 U245 ( .A(n272), .B(n213), .Z(product[11]) );
  NAND2_X1 U246 ( .A1(n20), .A2(n23), .ZN(n273) );
  NAND2_X1 U247 ( .A1(n20), .A2(n246), .ZN(n274) );
  NAND2_X1 U248 ( .A1(n23), .A2(n5), .ZN(n275) );
  XOR2_X1 U249 ( .A(n19), .B(n18), .Z(n276) );
  XOR2_X1 U250 ( .A(n276), .B(n270), .Z(product[12]) );
  NAND2_X1 U251 ( .A1(n19), .A2(n18), .ZN(n277) );
  NAND2_X1 U252 ( .A1(n269), .A2(n19), .ZN(n278) );
  NAND2_X1 U253 ( .A1(n269), .A2(n18), .ZN(n279) );
  NAND3_X1 U254 ( .A1(n279), .A2(n278), .A3(n277), .ZN(n3) );
  XOR2_X1 U255 ( .A(n103), .B(n96), .Z(n280) );
  XOR2_X1 U256 ( .A(n280), .B(n232), .Z(product[2]) );
  NAND2_X1 U257 ( .A1(n103), .A2(n96), .ZN(n281) );
  NAND2_X1 U258 ( .A1(n103), .A2(n232), .ZN(n282) );
  NAND2_X1 U259 ( .A1(n14), .A2(n96), .ZN(n283) );
  NAND3_X1 U260 ( .A1(n283), .A2(n282), .A3(n281), .ZN(n13) );
  XOR2_X1 U261 ( .A(n220), .B(n71), .Z(n284) );
  XOR2_X1 U262 ( .A(n284), .B(n268), .Z(product[3]) );
  NAND2_X1 U263 ( .A1(n56), .A2(n71), .ZN(n285) );
  NAND2_X1 U264 ( .A1(n56), .A2(n13), .ZN(n286) );
  NAND2_X1 U265 ( .A1(n267), .A2(n71), .ZN(n287) );
  NAND3_X1 U266 ( .A1(n287), .A2(n286), .A3(n285), .ZN(n12) );
  INV_X2 U267 ( .A(n253), .ZN(n299) );
  NAND3_X1 U268 ( .A1(n295), .A2(n294), .A3(n293), .ZN(n288) );
  XOR2_X1 U269 ( .A(a[2]), .B(n310), .Z(n289) );
  XOR2_X1 U270 ( .A(a[2]), .B(n310), .Z(n290) );
  INV_X1 U271 ( .A(n15), .ZN(n300) );
  AND3_X1 U272 ( .A1(n298), .A2(n297), .A3(n296), .ZN(product[15]) );
  INV_X1 U273 ( .A(n347), .ZN(n301) );
  INV_X1 U274 ( .A(n21), .ZN(n303) );
  INV_X1 U275 ( .A(n336), .ZN(n304) );
  INV_X1 U276 ( .A(n316), .ZN(n309) );
  INV_X1 U277 ( .A(n325), .ZN(n307) );
  INV_X1 U278 ( .A(n31), .ZN(n306) );
  INV_X1 U279 ( .A(a[0]), .ZN(n311) );
  INV_X1 U280 ( .A(a[5]), .ZN(n305) );
  INV_X1 U281 ( .A(a[7]), .ZN(n302) );
  INV_X1 U282 ( .A(a[3]), .ZN(n308) );
  XOR2_X1 U283 ( .A(n17), .B(n300), .Z(n292) );
  XOR2_X1 U284 ( .A(n212), .B(n292), .Z(product[13]) );
  NAND2_X1 U285 ( .A1(n17), .A2(n300), .ZN(n293) );
  NAND2_X1 U286 ( .A1(n17), .A2(n271), .ZN(n294) );
  NAND2_X1 U287 ( .A1(n3), .A2(n300), .ZN(n295) );
  NAND3_X1 U288 ( .A1(n295), .A2(n294), .A3(n293), .ZN(n2) );
  NAND2_X1 U289 ( .A1(n301), .A2(n15), .ZN(n296) );
  NAND2_X1 U290 ( .A1(n288), .A2(n301), .ZN(n297) );
  NAND2_X1 U291 ( .A1(n288), .A2(n15), .ZN(n298) );
  INV_X1 U292 ( .A(a[1]), .ZN(n310) );
  NOR2_X1 U293 ( .A1(n311), .A2(n253), .ZN(product[0]) );
  OAI22_X1 U294 ( .A1(n312), .A2(n313), .B1(n314), .B2(n311), .ZN(n99) );
  OAI22_X1 U295 ( .A1(n314), .A2(n313), .B1(n315), .B2(n311), .ZN(n98) );
  XNOR2_X1 U296 ( .A(b[6]), .B(a[1]), .ZN(n314) );
  OAI22_X1 U297 ( .A1(n311), .A2(n315), .B1(n313), .B2(n315), .ZN(n316) );
  XNOR2_X1 U298 ( .A(b[7]), .B(a[1]), .ZN(n315) );
  NOR2_X1 U299 ( .A1(n290), .A2(n253), .ZN(n96) );
  OAI22_X1 U300 ( .A1(n318), .A2(n319), .B1(n290), .B2(n320), .ZN(n95) );
  XNOR2_X1 U301 ( .A(a[3]), .B(n299), .ZN(n318) );
  OAI22_X1 U302 ( .A1(n320), .A2(n319), .B1(n290), .B2(n321), .ZN(n94) );
  XNOR2_X1 U303 ( .A(b[1]), .B(a[3]), .ZN(n320) );
  OAI22_X1 U304 ( .A1(n321), .A2(n319), .B1(n289), .B2(n322), .ZN(n93) );
  XNOR2_X1 U305 ( .A(b[2]), .B(a[3]), .ZN(n321) );
  OAI22_X1 U306 ( .A1(n322), .A2(n319), .B1(n289), .B2(n323), .ZN(n92) );
  XNOR2_X1 U307 ( .A(b[3]), .B(a[3]), .ZN(n322) );
  OAI22_X1 U308 ( .A1(n323), .A2(n319), .B1(n289), .B2(n324), .ZN(n91) );
  XNOR2_X1 U309 ( .A(b[4]), .B(a[3]), .ZN(n323) );
  OAI22_X1 U310 ( .A1(n326), .A2(n289), .B1(n319), .B2(n326), .ZN(n325) );
  NOR2_X1 U311 ( .A1(n242), .A2(n253), .ZN(n88) );
  OAI22_X1 U312 ( .A1(n328), .A2(n329), .B1(n241), .B2(n330), .ZN(n87) );
  XNOR2_X1 U313 ( .A(a[5]), .B(n299), .ZN(n328) );
  OAI22_X1 U314 ( .A1(n330), .A2(n329), .B1(n242), .B2(n331), .ZN(n86) );
  XNOR2_X1 U315 ( .A(b[1]), .B(a[5]), .ZN(n330) );
  OAI22_X1 U316 ( .A1(n331), .A2(n329), .B1(n241), .B2(n332), .ZN(n85) );
  XNOR2_X1 U317 ( .A(b[2]), .B(a[5]), .ZN(n331) );
  OAI22_X1 U318 ( .A1(n332), .A2(n329), .B1(n241), .B2(n333), .ZN(n84) );
  XNOR2_X1 U319 ( .A(b[3]), .B(a[5]), .ZN(n332) );
  OAI22_X1 U320 ( .A1(n333), .A2(n329), .B1(n242), .B2(n334), .ZN(n83) );
  XNOR2_X1 U321 ( .A(b[4]), .B(a[5]), .ZN(n333) );
  OAI22_X1 U322 ( .A1(n334), .A2(n329), .B1(n241), .B2(n335), .ZN(n82) );
  XNOR2_X1 U323 ( .A(b[5]), .B(a[5]), .ZN(n334) );
  OAI22_X1 U324 ( .A1(n337), .A2(n241), .B1(n329), .B2(n337), .ZN(n336) );
  NOR2_X1 U325 ( .A1(n338), .A2(n253), .ZN(n80) );
  OAI22_X1 U326 ( .A1(n339), .A2(n340), .B1(n338), .B2(n341), .ZN(n79) );
  XNOR2_X1 U327 ( .A(a[7]), .B(n299), .ZN(n339) );
  OAI22_X1 U328 ( .A1(n342), .A2(n340), .B1(n338), .B2(n343), .ZN(n77) );
  OAI22_X1 U329 ( .A1(n343), .A2(n340), .B1(n338), .B2(n344), .ZN(n76) );
  XNOR2_X1 U330 ( .A(b[3]), .B(a[7]), .ZN(n343) );
  OAI22_X1 U331 ( .A1(n344), .A2(n340), .B1(n338), .B2(n345), .ZN(n75) );
  XNOR2_X1 U332 ( .A(b[4]), .B(a[7]), .ZN(n344) );
  OAI22_X1 U333 ( .A1(n345), .A2(n340), .B1(n338), .B2(n346), .ZN(n74) );
  XNOR2_X1 U334 ( .A(b[5]), .B(a[7]), .ZN(n345) );
  OAI22_X1 U335 ( .A1(n348), .A2(n338), .B1(n340), .B2(n348), .ZN(n347) );
  OAI21_X1 U336 ( .B1(n299), .B2(n310), .A(n313), .ZN(n72) );
  OAI21_X1 U337 ( .B1(n308), .B2(n319), .A(n349), .ZN(n71) );
  OR3_X1 U338 ( .A1(n289), .A2(n299), .A3(n308), .ZN(n349) );
  OAI21_X1 U339 ( .B1(n305), .B2(n329), .A(n350), .ZN(n70) );
  OR3_X1 U340 ( .A1(n242), .A2(n299), .A3(n305), .ZN(n350) );
  OAI21_X1 U341 ( .B1(n302), .B2(n340), .A(n351), .ZN(n69) );
  OR3_X1 U342 ( .A1(n338), .A2(n299), .A3(n302), .ZN(n351) );
  XNOR2_X1 U343 ( .A(n352), .B(n353), .ZN(n38) );
  OR2_X1 U344 ( .A1(n352), .A2(n353), .ZN(n37) );
  OAI22_X1 U345 ( .A1(n324), .A2(n319), .B1(n289), .B2(n354), .ZN(n353) );
  XNOR2_X1 U346 ( .A(b[5]), .B(a[3]), .ZN(n324) );
  OAI22_X1 U347 ( .A1(n341), .A2(n340), .B1(n338), .B2(n342), .ZN(n352) );
  XNOR2_X1 U348 ( .A(b[2]), .B(a[7]), .ZN(n342) );
  XNOR2_X1 U349 ( .A(b[1]), .B(a[7]), .ZN(n341) );
  OAI22_X1 U350 ( .A1(n354), .A2(n319), .B1(n289), .B2(n326), .ZN(n31) );
  XNOR2_X1 U351 ( .A(b[7]), .B(a[3]), .ZN(n326) );
  XNOR2_X1 U352 ( .A(b[6]), .B(a[3]), .ZN(n354) );
  OAI22_X1 U353 ( .A1(n335), .A2(n329), .B1(n242), .B2(n337), .ZN(n21) );
  XNOR2_X1 U354 ( .A(b[7]), .B(a[5]), .ZN(n337) );
  XNOR2_X1 U355 ( .A(n209), .B(a[4]), .ZN(n356) );
  XNOR2_X1 U356 ( .A(b[6]), .B(a[5]), .ZN(n335) );
  OAI22_X1 U357 ( .A1(n346), .A2(n340), .B1(n338), .B2(n348), .ZN(n15) );
  XNOR2_X1 U358 ( .A(b[7]), .B(a[7]), .ZN(n348) );
  NAND2_X1 U359 ( .A1(n338), .A2(n357), .ZN(n340) );
  XNOR2_X1 U360 ( .A(n302), .B(a[6]), .ZN(n357) );
  XNOR2_X1 U361 ( .A(b[6]), .B(a[7]), .ZN(n346) );
  OAI22_X1 U362 ( .A1(n299), .A2(n313), .B1(n358), .B2(n311), .ZN(n104) );
  OAI22_X1 U363 ( .A1(n210), .A2(n313), .B1(n359), .B2(n311), .ZN(n103) );
  XNOR2_X1 U364 ( .A(b[1]), .B(a[1]), .ZN(n358) );
  OAI22_X1 U365 ( .A1(n359), .A2(n313), .B1(n360), .B2(n311), .ZN(n102) );
  XNOR2_X1 U366 ( .A(b[2]), .B(a[1]), .ZN(n359) );
  OAI22_X1 U367 ( .A1(n313), .A2(n360), .B1(n361), .B2(n311), .ZN(n101) );
  XNOR2_X1 U368 ( .A(b[3]), .B(a[1]), .ZN(n360) );
  OAI22_X1 U369 ( .A1(n361), .A2(n313), .B1(n312), .B2(n311), .ZN(n100) );
  XNOR2_X1 U370 ( .A(b[5]), .B(a[1]), .ZN(n312) );
  NAND2_X1 U371 ( .A1(a[1]), .A2(n311), .ZN(n313) );
  XNOR2_X1 U372 ( .A(b[4]), .B(a[1]), .ZN(n361) );
endmodule


module mac_30 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   n6, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, n2, n4;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(n6), .QN(n2) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_30_DW01_add_0 add_356 ( .A(pipeline), .B({mac_out[15:1], n6}), .CI(1'b0), 
        .SUM(sum) );
  mac_30_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n4), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n4), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n4), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n4), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n4), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n4), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n4), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n4), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n4), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n4), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n4), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n4), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n4), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n4), .ZN(N6) );
  INV_X1 U18 ( .A(n2), .ZN(mac_out[0]) );
  AND2_X1 U19 ( .A1(sum[0]), .A2(n4), .ZN(N3) );
  AND2_X1 U20 ( .A1(sum[15]), .A2(n4), .ZN(N18) );
  INV_X1 U21 ( .A(clear_acc), .ZN(n4) );
endmodule


module mac_29_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72;
  wire   [15:1] carry;

  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n72) );
  NAND3_X1 U2 ( .A1(n15), .A2(n16), .A3(n17), .ZN(n1) );
  NAND3_X1 U3 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n2) );
  NAND3_X1 U4 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n3) );
  NAND3_X1 U5 ( .A1(n11), .A2(n12), .A3(n13), .ZN(n4) );
  NAND3_X1 U6 ( .A1(n11), .A2(n12), .A3(n13), .ZN(n5) );
  NAND3_X1 U7 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n6) );
  NAND3_X1 U8 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n7) );
  NAND3_X1 U9 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n8) );
  XOR2_X1 U10 ( .A(B[15]), .B(A[15]), .Z(n9) );
  XOR2_X1 U11 ( .A(carry[15]), .B(n9), .Z(SUM[15]) );
  XOR2_X1 U12 ( .A(B[10]), .B(A[10]), .Z(n10) );
  XOR2_X1 U13 ( .A(carry[10]), .B(n10), .Z(SUM[10]) );
  NAND2_X1 U14 ( .A1(n3), .A2(B[10]), .ZN(n11) );
  NAND2_X1 U15 ( .A1(n2), .A2(A[10]), .ZN(n12) );
  NAND2_X1 U16 ( .A1(B[10]), .A2(A[10]), .ZN(n13) );
  NAND3_X1 U17 ( .A1(n11), .A2(n12), .A3(n13), .ZN(carry[11]) );
  XOR2_X1 U18 ( .A(B[11]), .B(A[11]), .Z(n14) );
  XOR2_X1 U19 ( .A(carry[11]), .B(n14), .Z(SUM[11]) );
  NAND2_X1 U20 ( .A1(n5), .A2(B[11]), .ZN(n15) );
  NAND2_X1 U21 ( .A1(n4), .A2(A[11]), .ZN(n16) );
  NAND2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n17) );
  NAND3_X1 U23 ( .A1(n15), .A2(n16), .A3(n17), .ZN(carry[12]) );
  XOR2_X1 U24 ( .A(B[4]), .B(A[4]), .Z(n18) );
  XOR2_X1 U25 ( .A(carry[4]), .B(n18), .Z(SUM[4]) );
  NAND2_X1 U26 ( .A1(carry[4]), .A2(B[4]), .ZN(n19) );
  NAND2_X1 U27 ( .A1(carry[4]), .A2(A[4]), .ZN(n20) );
  NAND2_X1 U28 ( .A1(B[4]), .A2(A[4]), .ZN(n21) );
  NAND3_X1 U29 ( .A1(n19), .A2(n20), .A3(n21), .ZN(carry[5]) );
  NAND3_X1 U30 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n22) );
  NAND3_X1 U31 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n23) );
  XOR2_X1 U32 ( .A(B[9]), .B(A[9]), .Z(n24) );
  XOR2_X1 U33 ( .A(n23), .B(n24), .Z(SUM[9]) );
  NAND2_X1 U34 ( .A1(n22), .A2(B[9]), .ZN(n25) );
  NAND2_X1 U35 ( .A1(carry[9]), .A2(A[9]), .ZN(n26) );
  NAND2_X1 U36 ( .A1(B[9]), .A2(A[9]), .ZN(n27) );
  NAND3_X1 U37 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[10]) );
  XOR2_X1 U38 ( .A(B[2]), .B(A[2]), .Z(n28) );
  XOR2_X1 U39 ( .A(carry[2]), .B(n28), .Z(SUM[2]) );
  NAND2_X1 U40 ( .A1(n7), .A2(B[2]), .ZN(n29) );
  NAND2_X1 U41 ( .A1(n6), .A2(A[2]), .ZN(n30) );
  NAND2_X1 U42 ( .A1(B[2]), .A2(A[2]), .ZN(n31) );
  NAND3_X1 U43 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[3]) );
  XOR2_X1 U44 ( .A(B[3]), .B(A[3]), .Z(n32) );
  XOR2_X1 U45 ( .A(n8), .B(n32), .Z(SUM[3]) );
  NAND2_X1 U46 ( .A1(n8), .A2(B[3]), .ZN(n33) );
  NAND2_X1 U47 ( .A1(carry[3]), .A2(A[3]), .ZN(n34) );
  NAND2_X1 U48 ( .A1(B[3]), .A2(A[3]), .ZN(n35) );
  NAND3_X1 U49 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[4]) );
  XOR2_X1 U50 ( .A(B[5]), .B(A[5]), .Z(n36) );
  XOR2_X1 U51 ( .A(carry[5]), .B(n36), .Z(SUM[5]) );
  NAND2_X1 U52 ( .A1(carry[5]), .A2(B[5]), .ZN(n37) );
  NAND2_X1 U53 ( .A1(carry[5]), .A2(A[5]), .ZN(n38) );
  NAND2_X1 U54 ( .A1(B[5]), .A2(A[5]), .ZN(n39) );
  NAND3_X1 U55 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[6]) );
  NAND3_X1 U56 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n40) );
  XOR2_X1 U57 ( .A(B[12]), .B(A[12]), .Z(n41) );
  XOR2_X1 U58 ( .A(n1), .B(n41), .Z(SUM[12]) );
  NAND2_X1 U59 ( .A1(n1), .A2(B[12]), .ZN(n42) );
  NAND2_X1 U60 ( .A1(carry[12]), .A2(A[12]), .ZN(n43) );
  NAND2_X1 U61 ( .A1(B[12]), .A2(A[12]), .ZN(n44) );
  NAND3_X1 U62 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[13]) );
  NAND3_X1 U63 ( .A1(n57), .A2(n58), .A3(n59), .ZN(n45) );
  NAND3_X1 U64 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n46) );
  NAND3_X1 U65 ( .A1(n69), .A2(n70), .A3(n71), .ZN(n47) );
  XOR2_X1 U66 ( .A(B[8]), .B(A[8]), .Z(n48) );
  XOR2_X1 U67 ( .A(carry[8]), .B(n48), .Z(SUM[8]) );
  NAND2_X1 U68 ( .A1(n47), .A2(B[8]), .ZN(n49) );
  NAND2_X1 U69 ( .A1(n47), .A2(A[8]), .ZN(n50) );
  NAND2_X1 U70 ( .A1(B[8]), .A2(A[8]), .ZN(n51) );
  NAND3_X1 U71 ( .A1(n49), .A2(n50), .A3(n51), .ZN(carry[9]) );
  XOR2_X1 U72 ( .A(B[1]), .B(A[1]), .Z(n52) );
  XOR2_X1 U73 ( .A(n72), .B(n52), .Z(SUM[1]) );
  NAND2_X1 U74 ( .A1(n72), .A2(B[1]), .ZN(n53) );
  NAND2_X1 U75 ( .A1(n72), .A2(A[1]), .ZN(n54) );
  NAND2_X1 U76 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  NAND3_X1 U77 ( .A1(n53), .A2(n54), .A3(n55), .ZN(carry[2]) );
  XOR2_X1 U78 ( .A(B[13]), .B(A[13]), .Z(n56) );
  XOR2_X1 U79 ( .A(carry[13]), .B(n56), .Z(SUM[13]) );
  NAND2_X1 U80 ( .A1(n40), .A2(B[13]), .ZN(n57) );
  NAND2_X1 U81 ( .A1(n40), .A2(A[13]), .ZN(n58) );
  NAND2_X1 U82 ( .A1(B[13]), .A2(A[13]), .ZN(n59) );
  NAND3_X1 U83 ( .A1(n58), .A2(n57), .A3(n59), .ZN(carry[14]) );
  XOR2_X1 U84 ( .A(B[6]), .B(A[6]), .Z(n60) );
  XOR2_X1 U85 ( .A(carry[6]), .B(n60), .Z(SUM[6]) );
  NAND2_X1 U86 ( .A1(carry[6]), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U87 ( .A1(carry[6]), .A2(A[6]), .ZN(n62) );
  NAND2_X1 U88 ( .A1(B[6]), .A2(A[6]), .ZN(n63) );
  NAND3_X1 U89 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[7]) );
  XOR2_X1 U90 ( .A(B[14]), .B(A[14]), .Z(n64) );
  XOR2_X1 U91 ( .A(n45), .B(n64), .Z(SUM[14]) );
  NAND2_X1 U92 ( .A1(n45), .A2(B[14]), .ZN(n65) );
  NAND2_X1 U93 ( .A1(carry[14]), .A2(A[14]), .ZN(n66) );
  NAND2_X1 U94 ( .A1(B[14]), .A2(A[14]), .ZN(n67) );
  NAND3_X1 U95 ( .A1(n65), .A2(n66), .A3(n67), .ZN(carry[15]) );
  XOR2_X1 U96 ( .A(B[7]), .B(A[7]), .Z(n68) );
  XOR2_X1 U97 ( .A(n46), .B(n68), .Z(SUM[7]) );
  NAND2_X1 U98 ( .A1(carry[7]), .A2(B[7]), .ZN(n69) );
  NAND2_X1 U99 ( .A1(carry[7]), .A2(A[7]), .ZN(n70) );
  NAND2_X1 U100 ( .A1(B[7]), .A2(A[7]), .ZN(n71) );
  NAND3_X1 U101 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[8]) );
  XOR2_X1 U102 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_29_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n316), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n315), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n319), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n318), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n321), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  NAND2_X2 U157 ( .A1(n339), .A2(n368), .ZN(n341) );
  BUF_X1 U158 ( .A(n311), .Z(n274) );
  AND2_X1 U159 ( .A1(n209), .A2(n102), .ZN(n206) );
  CLKBUF_X1 U160 ( .A(n46), .Z(n207) );
  XNOR2_X1 U161 ( .A(b[3]), .B(a[1]), .ZN(n208) );
  OAI22_X1 U162 ( .A1(n330), .A2(n331), .B1(n293), .B2(n332), .ZN(n209) );
  XOR2_X1 U163 ( .A(a[5]), .B(a[4]), .Z(n368) );
  CLKBUF_X1 U164 ( .A(b[3]), .Z(n210) );
  XOR2_X1 U165 ( .A(n207), .B(n49), .Z(n211) );
  XOR2_X1 U166 ( .A(n10), .B(n211), .Z(product[6]) );
  NAND2_X1 U167 ( .A1(n10), .A2(n46), .ZN(n212) );
  NAND2_X1 U168 ( .A1(n10), .A2(n49), .ZN(n213) );
  NAND2_X1 U169 ( .A1(n46), .A2(n49), .ZN(n214) );
  NAND3_X1 U170 ( .A1(n212), .A2(n213), .A3(n214), .ZN(n9) );
  NAND2_X2 U171 ( .A1(n236), .A2(n237), .ZN(n215) );
  NAND2_X1 U172 ( .A1(n236), .A2(n237), .ZN(n339) );
  CLKBUF_X1 U173 ( .A(n56), .Z(n216) );
  NAND2_X1 U174 ( .A1(n14), .A2(n96), .ZN(n217) );
  NAND2_X1 U175 ( .A1(n4), .A2(n18), .ZN(n218) );
  AND2_X1 U176 ( .A1(n104), .A2(n72), .ZN(n219) );
  NAND2_X1 U177 ( .A1(n256), .A2(n33), .ZN(n220) );
  NAND3_X1 U178 ( .A1(n290), .A2(n289), .A3(n291), .ZN(n221) );
  NAND2_X1 U179 ( .A1(n3), .A2(n17), .ZN(n222) );
  NAND2_X1 U180 ( .A1(n223), .A2(n20), .ZN(n305) );
  NAND3_X1 U181 ( .A1(n300), .A2(n299), .A3(n301), .ZN(n223) );
  XOR2_X2 U182 ( .A(a[6]), .B(n317), .Z(n350) );
  CLKBUF_X1 U183 ( .A(n240), .Z(n224) );
  CLKBUF_X1 U184 ( .A(n9), .Z(n225) );
  CLKBUF_X1 U185 ( .A(n268), .Z(n226) );
  CLKBUF_X1 U186 ( .A(n218), .Z(n227) );
  NAND3_X1 U187 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n228) );
  NAND3_X1 U188 ( .A1(n239), .A2(n224), .A3(n241), .ZN(n229) );
  XNOR2_X1 U189 ( .A(a[2]), .B(a[1]), .ZN(n329) );
  CLKBUF_X1 U190 ( .A(n306), .Z(n230) );
  NAND3_X1 U191 ( .A1(n263), .A2(n264), .A3(n265), .ZN(n231) );
  CLKBUF_X1 U192 ( .A(n221), .Z(n232) );
  CLKBUF_X1 U193 ( .A(n308), .Z(n233) );
  NAND2_X1 U194 ( .A1(a[4]), .A2(a[3]), .ZN(n236) );
  NAND2_X1 U195 ( .A1(n234), .A2(n235), .ZN(n237) );
  INV_X1 U196 ( .A(a[4]), .ZN(n234) );
  INV_X1 U197 ( .A(a[3]), .ZN(n235) );
  XOR2_X1 U198 ( .A(n40), .B(n45), .Z(n238) );
  XOR2_X1 U199 ( .A(n225), .B(n238), .Z(product[7]) );
  NAND2_X1 U200 ( .A1(n9), .A2(n40), .ZN(n239) );
  NAND2_X1 U201 ( .A1(n9), .A2(n45), .ZN(n240) );
  NAND2_X1 U202 ( .A1(n40), .A2(n45), .ZN(n241) );
  NAND3_X1 U203 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n8) );
  NAND3_X1 U204 ( .A1(n217), .A2(n251), .A3(n253), .ZN(n242) );
  NAND3_X1 U205 ( .A1(n251), .A2(n217), .A3(n253), .ZN(n243) );
  CLKBUF_X1 U206 ( .A(n231), .Z(n244) );
  NAND3_X1 U207 ( .A1(n307), .A2(n233), .A3(n227), .ZN(n245) );
  CLKBUF_X1 U208 ( .A(n12), .Z(n246) );
  XNOR2_X1 U209 ( .A(n247), .B(n273), .ZN(product[14]) );
  XNOR2_X1 U210 ( .A(n313), .B(n15), .ZN(n247) );
  AND3_X1 U211 ( .A1(n281), .A2(n280), .A3(n279), .ZN(product[15]) );
  NAND2_X1 U212 ( .A1(n287), .A2(n24), .ZN(n249) );
  XOR2_X1 U213 ( .A(n103), .B(n96), .Z(n250) );
  XOR2_X1 U214 ( .A(n219), .B(n250), .Z(product[2]) );
  NAND2_X1 U215 ( .A1(n219), .A2(n103), .ZN(n251) );
  NAND2_X1 U216 ( .A1(n14), .A2(n96), .ZN(n252) );
  NAND2_X1 U217 ( .A1(n103), .A2(n96), .ZN(n253) );
  NAND3_X1 U218 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n13) );
  NAND3_X1 U219 ( .A1(n259), .A2(n261), .A3(n260), .ZN(n254) );
  NAND2_X1 U220 ( .A1(n221), .A2(n27), .ZN(n255) );
  NAND3_X1 U221 ( .A1(n267), .A2(n268), .A3(n269), .ZN(n256) );
  NAND3_X1 U222 ( .A1(n267), .A2(n226), .A3(n269), .ZN(n257) );
  XOR2_X1 U223 ( .A(n216), .B(n71), .Z(n258) );
  XOR2_X1 U224 ( .A(n243), .B(n258), .Z(product[3]) );
  NAND2_X1 U225 ( .A1(n242), .A2(n56), .ZN(n259) );
  NAND2_X1 U226 ( .A1(n13), .A2(n71), .ZN(n260) );
  NAND2_X1 U227 ( .A1(n56), .A2(n71), .ZN(n261) );
  NAND3_X1 U228 ( .A1(n259), .A2(n261), .A3(n260), .ZN(n12) );
  XOR2_X1 U229 ( .A(n54), .B(n206), .Z(n262) );
  XOR2_X1 U230 ( .A(n246), .B(n262), .Z(product[4]) );
  NAND2_X1 U231 ( .A1(n12), .A2(n54), .ZN(n263) );
  NAND2_X1 U232 ( .A1(n254), .A2(n206), .ZN(n264) );
  NAND2_X1 U233 ( .A1(n54), .A2(n206), .ZN(n265) );
  NAND3_X1 U234 ( .A1(n263), .A2(n264), .A3(n265), .ZN(n11) );
  XOR2_X1 U235 ( .A(n34), .B(n39), .Z(n266) );
  XOR2_X1 U236 ( .A(n229), .B(n266), .Z(product[8]) );
  NAND2_X1 U237 ( .A1(n228), .A2(n34), .ZN(n267) );
  NAND2_X1 U238 ( .A1(n8), .A2(n39), .ZN(n268) );
  NAND2_X1 U239 ( .A1(n34), .A2(n39), .ZN(n269) );
  NAND3_X1 U240 ( .A1(n267), .A2(n268), .A3(n269), .ZN(n7) );
  NAND3_X1 U241 ( .A1(n308), .A2(n307), .A3(n309), .ZN(n270) );
  INV_X1 U242 ( .A(n311), .ZN(n271) );
  NAND3_X1 U243 ( .A1(n222), .A2(n278), .A3(n276), .ZN(n272) );
  NAND3_X1 U244 ( .A1(n222), .A2(n276), .A3(n278), .ZN(n273) );
  INV_X1 U245 ( .A(n311), .ZN(n310) );
  XOR2_X1 U246 ( .A(n17), .B(n312), .Z(n275) );
  XOR2_X1 U247 ( .A(n275), .B(n245), .Z(product[13]) );
  NAND2_X1 U248 ( .A1(n17), .A2(n312), .ZN(n276) );
  NAND2_X1 U249 ( .A1(n3), .A2(n17), .ZN(n277) );
  NAND2_X1 U250 ( .A1(n312), .A2(n270), .ZN(n278) );
  NAND3_X1 U251 ( .A1(n278), .A2(n276), .A3(n277), .ZN(n2) );
  NAND2_X1 U252 ( .A1(n313), .A2(n15), .ZN(n279) );
  NAND2_X1 U253 ( .A1(n2), .A2(n313), .ZN(n280) );
  NAND2_X1 U254 ( .A1(n272), .A2(n15), .ZN(n281) );
  XOR2_X1 U255 ( .A(n50), .B(n53), .Z(n282) );
  XOR2_X1 U256 ( .A(n244), .B(n282), .Z(product[5]) );
  NAND2_X1 U257 ( .A1(n231), .A2(n50), .ZN(n283) );
  NAND2_X1 U258 ( .A1(n11), .A2(n53), .ZN(n284) );
  NAND2_X1 U259 ( .A1(n50), .A2(n53), .ZN(n285) );
  NAND3_X1 U260 ( .A1(n283), .A2(n284), .A3(n285), .ZN(n10) );
  CLKBUF_X1 U261 ( .A(n255), .Z(n286) );
  NAND3_X1 U262 ( .A1(n290), .A2(n220), .A3(n291), .ZN(n287) );
  XOR2_X1 U263 ( .A(n95), .B(n102), .Z(n56) );
  NAND2_X2 U264 ( .A1(n329), .A2(n367), .ZN(n331) );
  XOR2_X1 U265 ( .A(n33), .B(n28), .Z(n288) );
  XOR2_X1 U266 ( .A(n257), .B(n288), .Z(product[9]) );
  NAND2_X1 U267 ( .A1(n256), .A2(n33), .ZN(n289) );
  NAND2_X1 U268 ( .A1(n7), .A2(n28), .ZN(n290) );
  NAND2_X1 U269 ( .A1(n33), .A2(n28), .ZN(n291) );
  NAND3_X1 U270 ( .A1(n220), .A2(n290), .A3(n291), .ZN(n6) );
  XOR2_X1 U271 ( .A(a[2]), .B(n322), .Z(n292) );
  XOR2_X1 U272 ( .A(a[2]), .B(n322), .Z(n293) );
  XNOR2_X1 U273 ( .A(n294), .B(n303), .ZN(product[12]) );
  XNOR2_X1 U274 ( .A(n19), .B(n18), .ZN(n294) );
  XNOR2_X1 U275 ( .A(n295), .B(n297), .ZN(product[11]) );
  XNOR2_X1 U276 ( .A(n20), .B(n23), .ZN(n295) );
  INV_X1 U277 ( .A(n15), .ZN(n312) );
  INV_X1 U278 ( .A(n337), .ZN(n319) );
  INV_X1 U279 ( .A(n348), .ZN(n316) );
  INV_X1 U280 ( .A(n21), .ZN(n315) );
  INV_X1 U281 ( .A(n328), .ZN(n321) );
  INV_X1 U282 ( .A(b[0]), .ZN(n311) );
  INV_X1 U283 ( .A(n359), .ZN(n313) );
  INV_X1 U284 ( .A(n31), .ZN(n318) );
  INV_X1 U285 ( .A(a[0]), .ZN(n323) );
  INV_X1 U286 ( .A(a[5]), .ZN(n317) );
  INV_X1 U287 ( .A(a[7]), .ZN(n314) );
  NAND3_X1 U288 ( .A1(n249), .A2(n255), .A3(n301), .ZN(n296) );
  NAND3_X1 U289 ( .A1(n249), .A2(n286), .A3(n301), .ZN(n297) );
  XOR2_X1 U290 ( .A(n24), .B(n27), .Z(n298) );
  XOR2_X1 U291 ( .A(n232), .B(n298), .Z(product[10]) );
  NAND2_X1 U292 ( .A1(n6), .A2(n24), .ZN(n299) );
  NAND2_X1 U293 ( .A1(n6), .A2(n27), .ZN(n300) );
  NAND2_X1 U294 ( .A1(n24), .A2(n27), .ZN(n301) );
  NAND3_X1 U295 ( .A1(n305), .A2(n306), .A3(n304), .ZN(n302) );
  NAND3_X1 U296 ( .A1(n304), .A2(n305), .A3(n230), .ZN(n303) );
  INV_X1 U297 ( .A(a[3]), .ZN(n320) );
  NAND2_X1 U298 ( .A1(n20), .A2(n23), .ZN(n304) );
  NAND2_X1 U299 ( .A1(n296), .A2(n23), .ZN(n306) );
  NAND3_X1 U300 ( .A1(n304), .A2(n305), .A3(n306), .ZN(n4) );
  NAND2_X1 U301 ( .A1(n19), .A2(n18), .ZN(n307) );
  NAND2_X1 U302 ( .A1(n302), .A2(n19), .ZN(n308) );
  NAND2_X1 U303 ( .A1(n4), .A2(n18), .ZN(n309) );
  NAND3_X1 U304 ( .A1(n218), .A2(n308), .A3(n307), .ZN(n3) );
  INV_X1 U305 ( .A(a[1]), .ZN(n322) );
  NOR2_X1 U306 ( .A1(n323), .A2(n274), .ZN(product[0]) );
  OAI22_X1 U307 ( .A1(n324), .A2(n325), .B1(n326), .B2(n323), .ZN(n99) );
  OAI22_X1 U308 ( .A1(n326), .A2(n325), .B1(n327), .B2(n323), .ZN(n98) );
  XNOR2_X1 U309 ( .A(b[6]), .B(a[1]), .ZN(n326) );
  OAI22_X1 U310 ( .A1(n323), .A2(n327), .B1(n325), .B2(n327), .ZN(n328) );
  XNOR2_X1 U311 ( .A(b[7]), .B(a[1]), .ZN(n327) );
  NOR2_X1 U312 ( .A1(n292), .A2(n274), .ZN(n96) );
  OAI22_X1 U313 ( .A1(n330), .A2(n331), .B1(n293), .B2(n332), .ZN(n95) );
  XNOR2_X1 U314 ( .A(a[3]), .B(n310), .ZN(n330) );
  OAI22_X1 U315 ( .A1(n332), .A2(n331), .B1(n293), .B2(n333), .ZN(n94) );
  XNOR2_X1 U316 ( .A(b[1]), .B(a[3]), .ZN(n332) );
  OAI22_X1 U317 ( .A1(n333), .A2(n331), .B1(n292), .B2(n334), .ZN(n93) );
  XNOR2_X1 U318 ( .A(b[2]), .B(a[3]), .ZN(n333) );
  OAI22_X1 U319 ( .A1(n334), .A2(n331), .B1(n293), .B2(n335), .ZN(n92) );
  XNOR2_X1 U320 ( .A(n210), .B(a[3]), .ZN(n334) );
  OAI22_X1 U321 ( .A1(n335), .A2(n331), .B1(n293), .B2(n336), .ZN(n91) );
  XNOR2_X1 U322 ( .A(b[4]), .B(a[3]), .ZN(n335) );
  OAI22_X1 U323 ( .A1(n338), .A2(n292), .B1(n331), .B2(n338), .ZN(n337) );
  NOR2_X1 U324 ( .A1(n215), .A2(n274), .ZN(n88) );
  OAI22_X1 U325 ( .A1(n340), .A2(n341), .B1(n215), .B2(n342), .ZN(n87) );
  XNOR2_X1 U326 ( .A(a[5]), .B(n271), .ZN(n340) );
  OAI22_X1 U327 ( .A1(n342), .A2(n341), .B1(n215), .B2(n343), .ZN(n86) );
  XNOR2_X1 U328 ( .A(b[1]), .B(a[5]), .ZN(n342) );
  OAI22_X1 U329 ( .A1(n343), .A2(n341), .B1(n215), .B2(n344), .ZN(n85) );
  XNOR2_X1 U330 ( .A(b[2]), .B(a[5]), .ZN(n343) );
  OAI22_X1 U331 ( .A1(n344), .A2(n341), .B1(n215), .B2(n345), .ZN(n84) );
  XNOR2_X1 U332 ( .A(n210), .B(a[5]), .ZN(n344) );
  OAI22_X1 U333 ( .A1(n345), .A2(n341), .B1(n215), .B2(n346), .ZN(n83) );
  XNOR2_X1 U334 ( .A(b[4]), .B(a[5]), .ZN(n345) );
  OAI22_X1 U335 ( .A1(n346), .A2(n341), .B1(n215), .B2(n347), .ZN(n82) );
  XNOR2_X1 U336 ( .A(b[5]), .B(a[5]), .ZN(n346) );
  OAI22_X1 U337 ( .A1(n349), .A2(n215), .B1(n341), .B2(n349), .ZN(n348) );
  NOR2_X1 U338 ( .A1(n350), .A2(n274), .ZN(n80) );
  OAI22_X1 U339 ( .A1(n351), .A2(n352), .B1(n350), .B2(n353), .ZN(n79) );
  XNOR2_X1 U340 ( .A(a[7]), .B(n271), .ZN(n351) );
  OAI22_X1 U341 ( .A1(n354), .A2(n352), .B1(n350), .B2(n355), .ZN(n77) );
  OAI22_X1 U342 ( .A1(n355), .A2(n352), .B1(n350), .B2(n356), .ZN(n76) );
  XNOR2_X1 U343 ( .A(n210), .B(a[7]), .ZN(n355) );
  OAI22_X1 U344 ( .A1(n356), .A2(n352), .B1(n350), .B2(n357), .ZN(n75) );
  XNOR2_X1 U345 ( .A(b[4]), .B(a[7]), .ZN(n356) );
  OAI22_X1 U346 ( .A1(n357), .A2(n352), .B1(n350), .B2(n358), .ZN(n74) );
  XNOR2_X1 U347 ( .A(b[5]), .B(a[7]), .ZN(n357) );
  OAI22_X1 U348 ( .A1(n360), .A2(n350), .B1(n352), .B2(n360), .ZN(n359) );
  OAI21_X1 U349 ( .B1(n310), .B2(n322), .A(n325), .ZN(n72) );
  OAI21_X1 U350 ( .B1(n320), .B2(n331), .A(n361), .ZN(n71) );
  OR3_X1 U351 ( .A1(n292), .A2(n271), .A3(n320), .ZN(n361) );
  OAI21_X1 U352 ( .B1(n317), .B2(n341), .A(n362), .ZN(n70) );
  OR3_X1 U353 ( .A1(n339), .A2(n271), .A3(n317), .ZN(n362) );
  OAI21_X1 U354 ( .B1(n314), .B2(n352), .A(n363), .ZN(n69) );
  OR3_X1 U355 ( .A1(n350), .A2(n271), .A3(n314), .ZN(n363) );
  XNOR2_X1 U356 ( .A(n364), .B(n365), .ZN(n38) );
  OR2_X1 U357 ( .A1(n364), .A2(n365), .ZN(n37) );
  OAI22_X1 U358 ( .A1(n336), .A2(n331), .B1(n292), .B2(n366), .ZN(n365) );
  XNOR2_X1 U359 ( .A(b[5]), .B(a[3]), .ZN(n336) );
  OAI22_X1 U360 ( .A1(n353), .A2(n352), .B1(n350), .B2(n354), .ZN(n364) );
  XNOR2_X1 U361 ( .A(b[2]), .B(a[7]), .ZN(n354) );
  XNOR2_X1 U362 ( .A(b[1]), .B(a[7]), .ZN(n353) );
  OAI22_X1 U363 ( .A1(n366), .A2(n331), .B1(n293), .B2(n338), .ZN(n31) );
  XNOR2_X1 U364 ( .A(b[7]), .B(a[3]), .ZN(n338) );
  XNOR2_X1 U365 ( .A(n320), .B(a[2]), .ZN(n367) );
  XNOR2_X1 U366 ( .A(b[6]), .B(a[3]), .ZN(n366) );
  OAI22_X1 U367 ( .A1(n347), .A2(n341), .B1(n215), .B2(n349), .ZN(n21) );
  XNOR2_X1 U368 ( .A(b[7]), .B(a[5]), .ZN(n349) );
  XNOR2_X1 U369 ( .A(b[6]), .B(a[5]), .ZN(n347) );
  OAI22_X1 U370 ( .A1(n358), .A2(n352), .B1(n350), .B2(n360), .ZN(n15) );
  XNOR2_X1 U371 ( .A(b[7]), .B(a[7]), .ZN(n360) );
  NAND2_X1 U372 ( .A1(n350), .A2(n369), .ZN(n352) );
  XNOR2_X1 U373 ( .A(n314), .B(a[6]), .ZN(n369) );
  XNOR2_X1 U374 ( .A(b[6]), .B(a[7]), .ZN(n358) );
  OAI22_X1 U375 ( .A1(n310), .A2(n325), .B1(n370), .B2(n323), .ZN(n104) );
  OAI22_X1 U376 ( .A1(n370), .A2(n325), .B1(n371), .B2(n323), .ZN(n103) );
  XNOR2_X1 U377 ( .A(b[1]), .B(a[1]), .ZN(n370) );
  OAI22_X1 U378 ( .A1(n371), .A2(n325), .B1(n372), .B2(n323), .ZN(n102) );
  XNOR2_X1 U379 ( .A(b[2]), .B(a[1]), .ZN(n371) );
  OAI22_X1 U380 ( .A1(n325), .A2(n208), .B1(n373), .B2(n323), .ZN(n101) );
  XNOR2_X1 U381 ( .A(b[3]), .B(a[1]), .ZN(n372) );
  OAI22_X1 U382 ( .A1(n373), .A2(n325), .B1(n324), .B2(n323), .ZN(n100) );
  XNOR2_X1 U383 ( .A(b[5]), .B(a[1]), .ZN(n324) );
  NAND2_X1 U384 ( .A1(a[1]), .A2(n323), .ZN(n325) );
  XNOR2_X1 U385 ( .A(b[4]), .B(a[1]), .ZN(n373) );
endmodule


module mac_29 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_29_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_29_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X2 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_28_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;
  wire   [15:1] carry;

  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n76), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[15]), .B(A[15]), .Z(n1) );
  XOR2_X1 U2 ( .A(carry[15]), .B(n1), .Z(SUM[15]) );
  FA_X1 U3 ( .A(A[1]), .B(B[1]), .CI(n76), .CO(n2) );
  FA_X1 U4 ( .A(A[1]), .B(B[1]), .CI(n76), .CO(n3) );
  AND2_X2 U5 ( .A1(B[0]), .A2(A[0]), .ZN(n76) );
  NAND3_X1 U6 ( .A1(n15), .A2(n16), .A3(n17), .ZN(n4) );
  NAND3_X1 U7 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n5) );
  NAND3_X1 U8 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n6) );
  NAND3_X1 U9 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n7) );
  NAND3_X1 U10 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n8) );
  NAND3_X1 U11 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n9) );
  NAND3_X1 U12 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n10) );
  NAND3_X1 U13 ( .A1(n20), .A2(n19), .A3(n21), .ZN(n11) );
  NAND3_X1 U14 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n12) );
  NAND3_X1 U15 ( .A1(n35), .A2(n36), .A3(n37), .ZN(n13) );
  XOR2_X1 U16 ( .A(B[10]), .B(A[10]), .Z(n14) );
  XOR2_X1 U17 ( .A(n6), .B(n14), .Z(SUM[10]) );
  NAND2_X1 U18 ( .A1(n5), .A2(B[10]), .ZN(n15) );
  NAND2_X1 U19 ( .A1(carry[10]), .A2(A[10]), .ZN(n16) );
  NAND2_X1 U20 ( .A1(B[10]), .A2(A[10]), .ZN(n17) );
  NAND3_X1 U21 ( .A1(n15), .A2(n16), .A3(n17), .ZN(carry[11]) );
  XOR2_X1 U22 ( .A(B[4]), .B(A[4]), .Z(n18) );
  XOR2_X1 U23 ( .A(n8), .B(n18), .Z(SUM[4]) );
  NAND2_X1 U24 ( .A1(n7), .A2(B[4]), .ZN(n19) );
  NAND2_X1 U25 ( .A1(carry[4]), .A2(A[4]), .ZN(n20) );
  NAND2_X1 U26 ( .A1(B[4]), .A2(A[4]), .ZN(n21) );
  NAND3_X1 U27 ( .A1(n19), .A2(n20), .A3(n21), .ZN(carry[5]) );
  NAND3_X1 U28 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n22) );
  NAND3_X1 U29 ( .A1(n35), .A2(n36), .A3(n37), .ZN(n23) );
  NAND3_X1 U30 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n24) );
  NAND3_X1 U31 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n25) );
  XOR2_X1 U32 ( .A(B[11]), .B(A[11]), .Z(n26) );
  XOR2_X1 U33 ( .A(n4), .B(n26), .Z(SUM[11]) );
  NAND2_X1 U34 ( .A1(n4), .A2(B[11]), .ZN(n27) );
  NAND2_X1 U35 ( .A1(carry[11]), .A2(A[11]), .ZN(n28) );
  NAND2_X1 U36 ( .A1(B[11]), .A2(A[11]), .ZN(n29) );
  NAND3_X1 U37 ( .A1(n27), .A2(n28), .A3(n29), .ZN(carry[12]) );
  NAND3_X1 U38 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n30) );
  NAND3_X1 U39 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n31) );
  NAND3_X1 U40 ( .A1(n73), .A2(n74), .A3(n75), .ZN(n32) );
  NAND3_X1 U41 ( .A1(n73), .A2(n74), .A3(n75), .ZN(n33) );
  XOR2_X1 U42 ( .A(B[8]), .B(A[8]), .Z(n34) );
  XOR2_X1 U43 ( .A(n33), .B(n34), .Z(SUM[8]) );
  NAND2_X1 U44 ( .A1(n32), .A2(B[8]), .ZN(n35) );
  NAND2_X1 U45 ( .A1(carry[8]), .A2(A[8]), .ZN(n36) );
  NAND2_X1 U46 ( .A1(B[8]), .A2(A[8]), .ZN(n37) );
  NAND3_X1 U47 ( .A1(n35), .A2(n36), .A3(n37), .ZN(carry[9]) );
  XOR2_X1 U48 ( .A(B[9]), .B(A[9]), .Z(n38) );
  XOR2_X1 U49 ( .A(n23), .B(n38), .Z(SUM[9]) );
  NAND2_X1 U50 ( .A1(n13), .A2(B[9]), .ZN(n39) );
  NAND2_X1 U51 ( .A1(carry[9]), .A2(A[9]), .ZN(n40) );
  NAND2_X1 U52 ( .A1(B[9]), .A2(A[9]), .ZN(n41) );
  NAND3_X1 U53 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[10]) );
  XOR2_X1 U54 ( .A(B[2]), .B(A[2]), .Z(n42) );
  XOR2_X1 U55 ( .A(n3), .B(n42), .Z(SUM[2]) );
  NAND2_X1 U56 ( .A1(n2), .A2(B[2]), .ZN(n43) );
  NAND2_X1 U57 ( .A1(carry[2]), .A2(A[2]), .ZN(n44) );
  NAND2_X1 U58 ( .A1(B[2]), .A2(A[2]), .ZN(n45) );
  NAND3_X1 U59 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[3]) );
  XOR2_X1 U60 ( .A(B[3]), .B(A[3]), .Z(n46) );
  XOR2_X1 U61 ( .A(n25), .B(n46), .Z(SUM[3]) );
  NAND2_X1 U62 ( .A1(n24), .A2(B[3]), .ZN(n47) );
  NAND2_X1 U63 ( .A1(carry[3]), .A2(A[3]), .ZN(n48) );
  NAND2_X1 U64 ( .A1(B[3]), .A2(A[3]), .ZN(n49) );
  NAND3_X1 U65 ( .A1(n47), .A2(n48), .A3(n49), .ZN(carry[4]) );
  XOR2_X1 U66 ( .A(B[12]), .B(A[12]), .Z(n50) );
  XOR2_X1 U67 ( .A(n10), .B(n50), .Z(SUM[12]) );
  NAND2_X1 U68 ( .A1(n10), .A2(B[12]), .ZN(n51) );
  NAND2_X1 U69 ( .A1(carry[12]), .A2(A[12]), .ZN(n52) );
  NAND2_X1 U70 ( .A1(B[12]), .A2(A[12]), .ZN(n53) );
  NAND3_X1 U71 ( .A1(n51), .A2(n52), .A3(n53), .ZN(carry[13]) );
  XOR2_X1 U72 ( .A(B[5]), .B(A[5]), .Z(n54) );
  XOR2_X1 U73 ( .A(n11), .B(n54), .Z(SUM[5]) );
  NAND2_X1 U74 ( .A1(n11), .A2(B[5]), .ZN(n55) );
  NAND2_X1 U75 ( .A1(carry[5]), .A2(A[5]), .ZN(n56) );
  NAND2_X1 U76 ( .A1(B[5]), .A2(A[5]), .ZN(n57) );
  NAND3_X1 U77 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[6]) );
  NAND3_X1 U78 ( .A1(n62), .A2(n61), .A3(n63), .ZN(n58) );
  NAND3_X1 U79 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n59) );
  XOR2_X1 U80 ( .A(B[13]), .B(A[13]), .Z(n60) );
  XOR2_X1 U81 ( .A(carry[13]), .B(n60), .Z(SUM[13]) );
  NAND2_X1 U82 ( .A1(n9), .A2(B[13]), .ZN(n61) );
  NAND2_X1 U83 ( .A1(n22), .A2(A[13]), .ZN(n62) );
  NAND2_X1 U84 ( .A1(B[13]), .A2(A[13]), .ZN(n63) );
  NAND3_X1 U85 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[14]) );
  XOR2_X1 U86 ( .A(B[6]), .B(A[6]), .Z(n64) );
  XOR2_X1 U87 ( .A(n31), .B(n64), .Z(SUM[6]) );
  NAND2_X1 U88 ( .A1(n30), .A2(B[6]), .ZN(n65) );
  NAND2_X1 U89 ( .A1(carry[6]), .A2(A[6]), .ZN(n66) );
  NAND2_X1 U90 ( .A1(B[6]), .A2(A[6]), .ZN(n67) );
  NAND3_X1 U91 ( .A1(n65), .A2(n66), .A3(n67), .ZN(carry[7]) );
  XOR2_X1 U92 ( .A(B[14]), .B(A[14]), .Z(n68) );
  XOR2_X1 U93 ( .A(carry[14]), .B(n68), .Z(SUM[14]) );
  NAND2_X1 U94 ( .A1(carry[14]), .A2(B[14]), .ZN(n69) );
  NAND2_X1 U95 ( .A1(n58), .A2(A[14]), .ZN(n70) );
  NAND2_X1 U96 ( .A1(B[14]), .A2(A[14]), .ZN(n71) );
  NAND3_X1 U97 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[15]) );
  XOR2_X1 U98 ( .A(B[7]), .B(A[7]), .Z(n72) );
  XOR2_X1 U99 ( .A(n12), .B(n72), .Z(SUM[7]) );
  NAND2_X1 U100 ( .A1(carry[7]), .A2(B[7]), .ZN(n73) );
  NAND2_X1 U101 ( .A1(n59), .A2(A[7]), .ZN(n74) );
  NAND2_X1 U102 ( .A1(B[7]), .A2(A[7]), .ZN(n75) );
  NAND3_X1 U103 ( .A1(n73), .A2(n74), .A3(n75), .ZN(carry[8]) );
  XOR2_X1 U104 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_28_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n311), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n310), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n314), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n313), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n316), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U33 ( .A(n92), .B(n80), .CI(n99), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n94), .B(n88), .CI(n101), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n102), .B(n95), .CO(n55), .S(n56) );
  NAND3_X1 U157 ( .A1(n299), .A2(n300), .A3(n301), .ZN(n49) );
  NAND3_X1 U158 ( .A1(n295), .A2(n296), .A3(n294), .ZN(n206) );
  NAND3_X1 U159 ( .A1(n295), .A2(n296), .A3(n294), .ZN(n207) );
  AND3_X1 U160 ( .A1(n210), .A2(n211), .A3(n212), .ZN(product[15]) );
  XOR2_X1 U161 ( .A(n308), .B(n15), .Z(n209) );
  XOR2_X1 U162 ( .A(n2), .B(n209), .Z(product[14]) );
  NAND2_X1 U163 ( .A1(n207), .A2(n308), .ZN(n210) );
  NAND2_X1 U164 ( .A1(n206), .A2(n15), .ZN(n211) );
  NAND2_X1 U165 ( .A1(n308), .A2(n15), .ZN(n212) );
  NAND2_X1 U166 ( .A1(n234), .A2(n18), .ZN(n213) );
  XOR2_X1 U167 ( .A(a[3]), .B(a[2]), .Z(n362) );
  NAND2_X1 U168 ( .A1(n14), .A2(n96), .ZN(n214) );
  CLKBUF_X1 U169 ( .A(b[1]), .Z(n215) );
  INV_X1 U170 ( .A(n288), .ZN(n216) );
  CLKBUF_X1 U171 ( .A(b[1]), .Z(n217) );
  NAND2_X1 U172 ( .A1(n10), .A2(n49), .ZN(n218) );
  XOR2_X1 U173 ( .A(n51), .B(n86), .Z(n219) );
  XOR2_X1 U174 ( .A(n48), .B(n219), .Z(n46) );
  NAND2_X1 U175 ( .A1(n48), .A2(n51), .ZN(n220) );
  NAND2_X1 U176 ( .A1(n48), .A2(n86), .ZN(n221) );
  NAND2_X1 U177 ( .A1(n51), .A2(n86), .ZN(n222) );
  NAND3_X1 U178 ( .A1(n220), .A2(n221), .A3(n222), .ZN(n45) );
  NAND2_X1 U179 ( .A1(b[3]), .A2(a[1]), .ZN(n224) );
  NAND2_X1 U180 ( .A1(n223), .A2(n317), .ZN(n225) );
  NAND2_X1 U181 ( .A1(n224), .A2(n225), .ZN(n367) );
  INV_X1 U182 ( .A(b[3]), .ZN(n223) );
  CLKBUF_X1 U183 ( .A(b[3]), .Z(n226) );
  CLKBUF_X1 U184 ( .A(n12), .Z(n227) );
  AND2_X1 U185 ( .A1(n104), .A2(n72), .ZN(n228) );
  CLKBUF_X1 U186 ( .A(n236), .Z(n229) );
  NAND3_X1 U187 ( .A1(n218), .A2(n269), .A3(n271), .ZN(n230) );
  NAND3_X1 U188 ( .A1(n213), .A2(n291), .A3(n290), .ZN(n231) );
  NAND3_X1 U189 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n232) );
  NAND3_X1 U190 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n233) );
  NAND3_X1 U191 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n234) );
  NAND3_X1 U192 ( .A1(n239), .A2(n238), .A3(n240), .ZN(n235) );
  NAND3_X1 U193 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n236) );
  XOR2_X1 U194 ( .A(n103), .B(n96), .Z(n237) );
  XOR2_X1 U195 ( .A(n228), .B(n237), .Z(product[2]) );
  NAND2_X1 U196 ( .A1(n228), .A2(n103), .ZN(n238) );
  NAND2_X1 U197 ( .A1(n14), .A2(n96), .ZN(n239) );
  NAND2_X1 U198 ( .A1(n103), .A2(n96), .ZN(n240) );
  NAND3_X1 U199 ( .A1(n238), .A2(n214), .A3(n240), .ZN(n13) );
  XNOR2_X2 U200 ( .A(a[4]), .B(a[3]), .ZN(n334) );
  XOR2_X1 U201 ( .A(n23), .B(n20), .Z(n241) );
  XOR2_X1 U202 ( .A(n229), .B(n241), .Z(product[11]) );
  NAND2_X1 U203 ( .A1(n236), .A2(n23), .ZN(n242) );
  NAND2_X1 U204 ( .A1(n5), .A2(n20), .ZN(n243) );
  NAND2_X1 U205 ( .A1(n23), .A2(n20), .ZN(n244) );
  NAND3_X1 U206 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n4) );
  NAND3_X1 U207 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n245) );
  NAND3_X1 U208 ( .A1(n262), .A2(n264), .A3(n263), .ZN(n246) );
  NAND3_X1 U209 ( .A1(n269), .A2(n218), .A3(n271), .ZN(n247) );
  CLKBUF_X1 U210 ( .A(n232), .Z(n248) );
  NAND3_X1 U211 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n249) );
  XOR2_X1 U212 ( .A(n40), .B(n45), .Z(n250) );
  XOR2_X1 U213 ( .A(n247), .B(n250), .Z(product[7]) );
  NAND2_X1 U214 ( .A1(n230), .A2(n40), .ZN(n251) );
  NAND2_X1 U215 ( .A1(n9), .A2(n45), .ZN(n252) );
  NAND2_X1 U216 ( .A1(n40), .A2(n45), .ZN(n253) );
  NAND3_X1 U217 ( .A1(n252), .A2(n251), .A3(n253), .ZN(n8) );
  CLKBUF_X1 U218 ( .A(n234), .Z(n254) );
  CLKBUF_X1 U219 ( .A(n233), .Z(n255) );
  XNOR2_X1 U220 ( .A(n215), .B(a[1]), .ZN(n256) );
  XOR2_X1 U221 ( .A(n34), .B(n39), .Z(n257) );
  XOR2_X1 U222 ( .A(n248), .B(n257), .Z(product[8]) );
  NAND2_X1 U223 ( .A1(n232), .A2(n34), .ZN(n258) );
  NAND2_X1 U224 ( .A1(n8), .A2(n39), .ZN(n259) );
  NAND2_X1 U225 ( .A1(n34), .A2(n39), .ZN(n260) );
  XOR2_X1 U226 ( .A(n56), .B(n71), .Z(n261) );
  XOR2_X1 U227 ( .A(n235), .B(n261), .Z(product[3]) );
  NAND2_X1 U228 ( .A1(n235), .A2(n56), .ZN(n262) );
  NAND2_X1 U229 ( .A1(n13), .A2(n71), .ZN(n263) );
  NAND2_X1 U230 ( .A1(n56), .A2(n71), .ZN(n264) );
  NAND3_X1 U231 ( .A1(n262), .A2(n264), .A3(n263), .ZN(n12) );
  CLKBUF_X1 U232 ( .A(n249), .Z(n265) );
  NAND3_X1 U233 ( .A1(n302), .A2(n304), .A3(n303), .ZN(n266) );
  NAND3_X1 U234 ( .A1(n302), .A2(n303), .A3(n304), .ZN(n267) );
  XOR2_X1 U235 ( .A(n46), .B(n49), .Z(n268) );
  XOR2_X1 U236 ( .A(n267), .B(n268), .Z(product[6]) );
  NAND2_X1 U237 ( .A1(n266), .A2(n46), .ZN(n269) );
  NAND2_X1 U238 ( .A1(n10), .A2(n49), .ZN(n270) );
  NAND2_X1 U239 ( .A1(n46), .A2(n49), .ZN(n271) );
  NAND3_X1 U240 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n9) );
  XOR2_X1 U241 ( .A(n33), .B(n28), .Z(n272) );
  XOR2_X1 U242 ( .A(n255), .B(n272), .Z(product[9]) );
  NAND2_X1 U243 ( .A1(n233), .A2(n33), .ZN(n273) );
  NAND2_X1 U244 ( .A1(n245), .A2(n28), .ZN(n274) );
  NAND2_X1 U245 ( .A1(n33), .A2(n28), .ZN(n275) );
  NAND3_X1 U246 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n6) );
  XNOR2_X2 U247 ( .A(a[2]), .B(a[1]), .ZN(n276) );
  XNOR2_X1 U248 ( .A(a[2]), .B(a[1]), .ZN(n324) );
  NAND2_X2 U249 ( .A1(n334), .A2(n363), .ZN(n336) );
  XOR2_X1 U250 ( .A(n24), .B(n27), .Z(n277) );
  XOR2_X1 U251 ( .A(n265), .B(n277), .Z(product[10]) );
  NAND2_X1 U252 ( .A1(n249), .A2(n24), .ZN(n278) );
  NAND2_X1 U253 ( .A1(n6), .A2(n27), .ZN(n279) );
  NAND2_X1 U254 ( .A1(n24), .A2(n27), .ZN(n280) );
  NAND3_X1 U255 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n5) );
  NAND3_X1 U256 ( .A1(n285), .A2(n284), .A3(n286), .ZN(n281) );
  NAND3_X1 U257 ( .A1(n284), .A2(n285), .A3(n286), .ZN(n282) );
  XOR2_X1 U258 ( .A(n54), .B(n55), .Z(n283) );
  XOR2_X1 U259 ( .A(n227), .B(n283), .Z(product[4]) );
  NAND2_X1 U260 ( .A1(n246), .A2(n54), .ZN(n284) );
  NAND2_X1 U261 ( .A1(n12), .A2(n55), .ZN(n285) );
  NAND2_X1 U262 ( .A1(n54), .A2(n55), .ZN(n286) );
  NAND3_X1 U263 ( .A1(n285), .A2(n284), .A3(n286), .ZN(n11) );
  NAND3_X1 U264 ( .A1(n213), .A2(n291), .A3(n290), .ZN(n287) );
  INV_X1 U265 ( .A(n306), .ZN(n288) );
  XOR2_X1 U266 ( .A(n297), .B(n52), .Z(n50) );
  INV_X1 U267 ( .A(n15), .ZN(n307) );
  INV_X1 U268 ( .A(n343), .ZN(n311) );
  INV_X1 U269 ( .A(n21), .ZN(n310) );
  INV_X1 U270 ( .A(n323), .ZN(n316) );
  INV_X1 U271 ( .A(n332), .ZN(n314) );
  INV_X1 U272 ( .A(b[0]), .ZN(n306) );
  INV_X1 U273 ( .A(n354), .ZN(n308) );
  INV_X1 U274 ( .A(n31), .ZN(n313) );
  INV_X1 U275 ( .A(a[0]), .ZN(n318) );
  INV_X1 U276 ( .A(a[5]), .ZN(n312) );
  INV_X1 U277 ( .A(a[7]), .ZN(n309) );
  XOR2_X1 U278 ( .A(n19), .B(n18), .Z(n289) );
  XOR2_X1 U279 ( .A(n289), .B(n254), .Z(product[12]) );
  NAND2_X1 U280 ( .A1(n19), .A2(n18), .ZN(n290) );
  NAND2_X1 U281 ( .A1(n19), .A2(n4), .ZN(n291) );
  NAND2_X1 U282 ( .A1(n234), .A2(n18), .ZN(n292) );
  NAND3_X1 U283 ( .A1(n292), .A2(n291), .A3(n290), .ZN(n3) );
  XOR2_X1 U284 ( .A(n17), .B(n307), .Z(n293) );
  XOR2_X1 U285 ( .A(n293), .B(n287), .Z(product[13]) );
  NAND2_X1 U286 ( .A1(n17), .A2(n307), .ZN(n294) );
  NAND2_X1 U287 ( .A1(n231), .A2(n17), .ZN(n295) );
  NAND2_X1 U288 ( .A1(n3), .A2(n307), .ZN(n296) );
  NAND3_X1 U289 ( .A1(n295), .A2(n296), .A3(n294), .ZN(n2) );
  XOR2_X1 U290 ( .A(n93), .B(n100), .Z(n297) );
  XOR2_X1 U291 ( .A(n53), .B(n282), .Z(n298) );
  XOR2_X1 U292 ( .A(n298), .B(n50), .Z(product[5]) );
  NAND2_X1 U293 ( .A1(n93), .A2(n100), .ZN(n299) );
  NAND2_X1 U294 ( .A1(n93), .A2(n52), .ZN(n300) );
  NAND2_X1 U295 ( .A1(n100), .A2(n52), .ZN(n301) );
  NAND2_X1 U296 ( .A1(n53), .A2(n281), .ZN(n302) );
  NAND2_X1 U297 ( .A1(n53), .A2(n50), .ZN(n303) );
  NAND2_X1 U298 ( .A1(n11), .A2(n50), .ZN(n304) );
  NAND3_X1 U299 ( .A1(n302), .A2(n304), .A3(n303), .ZN(n10) );
  INV_X1 U300 ( .A(a[3]), .ZN(n315) );
  INV_X1 U301 ( .A(a[1]), .ZN(n317) );
  NAND2_X2 U302 ( .A1(n324), .A2(n362), .ZN(n326) );
  XOR2_X2 U303 ( .A(a[6]), .B(n312), .Z(n345) );
  INV_X1 U304 ( .A(n306), .ZN(n305) );
  NOR2_X1 U305 ( .A1(n318), .A2(n216), .ZN(product[0]) );
  OAI22_X1 U306 ( .A1(n319), .A2(n320), .B1(n321), .B2(n318), .ZN(n99) );
  OAI22_X1 U307 ( .A1(n321), .A2(n320), .B1(n322), .B2(n318), .ZN(n98) );
  XNOR2_X1 U308 ( .A(b[6]), .B(a[1]), .ZN(n321) );
  OAI22_X1 U309 ( .A1(n318), .A2(n322), .B1(n320), .B2(n322), .ZN(n323) );
  XNOR2_X1 U310 ( .A(b[7]), .B(a[1]), .ZN(n322) );
  NOR2_X1 U311 ( .A1(n276), .A2(n216), .ZN(n96) );
  OAI22_X1 U312 ( .A1(n325), .A2(n326), .B1(n276), .B2(n327), .ZN(n95) );
  XNOR2_X1 U313 ( .A(a[3]), .B(n305), .ZN(n325) );
  OAI22_X1 U314 ( .A1(n327), .A2(n326), .B1(n276), .B2(n328), .ZN(n94) );
  XNOR2_X1 U315 ( .A(b[1]), .B(a[3]), .ZN(n327) );
  OAI22_X1 U316 ( .A1(n328), .A2(n326), .B1(n276), .B2(n329), .ZN(n93) );
  XNOR2_X1 U317 ( .A(b[2]), .B(a[3]), .ZN(n328) );
  OAI22_X1 U318 ( .A1(n329), .A2(n326), .B1(n276), .B2(n330), .ZN(n92) );
  XNOR2_X1 U319 ( .A(n226), .B(a[3]), .ZN(n329) );
  OAI22_X1 U320 ( .A1(n330), .A2(n326), .B1(n276), .B2(n331), .ZN(n91) );
  XNOR2_X1 U321 ( .A(b[4]), .B(a[3]), .ZN(n330) );
  OAI22_X1 U322 ( .A1(n333), .A2(n276), .B1(n326), .B2(n333), .ZN(n332) );
  NOR2_X1 U323 ( .A1(n334), .A2(n216), .ZN(n88) );
  OAI22_X1 U324 ( .A1(n335), .A2(n336), .B1(n334), .B2(n337), .ZN(n87) );
  XNOR2_X1 U325 ( .A(a[5]), .B(n288), .ZN(n335) );
  OAI22_X1 U326 ( .A1(n337), .A2(n336), .B1(n334), .B2(n338), .ZN(n86) );
  XNOR2_X1 U327 ( .A(a[5]), .B(n217), .ZN(n337) );
  OAI22_X1 U328 ( .A1(n338), .A2(n336), .B1(n334), .B2(n339), .ZN(n85) );
  XNOR2_X1 U329 ( .A(b[2]), .B(a[5]), .ZN(n338) );
  OAI22_X1 U330 ( .A1(n339), .A2(n336), .B1(n334), .B2(n340), .ZN(n84) );
  XNOR2_X1 U331 ( .A(n226), .B(a[5]), .ZN(n339) );
  OAI22_X1 U332 ( .A1(n340), .A2(n336), .B1(n334), .B2(n341), .ZN(n83) );
  XNOR2_X1 U333 ( .A(b[4]), .B(a[5]), .ZN(n340) );
  OAI22_X1 U334 ( .A1(n341), .A2(n336), .B1(n334), .B2(n342), .ZN(n82) );
  XNOR2_X1 U335 ( .A(b[5]), .B(a[5]), .ZN(n341) );
  OAI22_X1 U336 ( .A1(n344), .A2(n334), .B1(n336), .B2(n344), .ZN(n343) );
  NOR2_X1 U337 ( .A1(n345), .A2(n216), .ZN(n80) );
  OAI22_X1 U338 ( .A1(n346), .A2(n347), .B1(n345), .B2(n348), .ZN(n79) );
  XNOR2_X1 U339 ( .A(a[7]), .B(n288), .ZN(n346) );
  OAI22_X1 U340 ( .A1(n349), .A2(n347), .B1(n345), .B2(n350), .ZN(n77) );
  OAI22_X1 U341 ( .A1(n350), .A2(n347), .B1(n345), .B2(n351), .ZN(n76) );
  XNOR2_X1 U342 ( .A(n226), .B(a[7]), .ZN(n350) );
  OAI22_X1 U343 ( .A1(n351), .A2(n347), .B1(n345), .B2(n352), .ZN(n75) );
  XNOR2_X1 U344 ( .A(b[4]), .B(a[7]), .ZN(n351) );
  OAI22_X1 U345 ( .A1(n352), .A2(n347), .B1(n345), .B2(n353), .ZN(n74) );
  XNOR2_X1 U346 ( .A(b[5]), .B(a[7]), .ZN(n352) );
  OAI22_X1 U347 ( .A1(n355), .A2(n345), .B1(n347), .B2(n355), .ZN(n354) );
  OAI21_X1 U348 ( .B1(n305), .B2(n317), .A(n320), .ZN(n72) );
  OAI21_X1 U349 ( .B1(n315), .B2(n326), .A(n356), .ZN(n71) );
  OR3_X1 U350 ( .A1(n276), .A2(n288), .A3(n315), .ZN(n356) );
  OAI21_X1 U351 ( .B1(n312), .B2(n336), .A(n357), .ZN(n70) );
  OR3_X1 U352 ( .A1(n334), .A2(n288), .A3(n312), .ZN(n357) );
  OAI21_X1 U353 ( .B1(n309), .B2(n347), .A(n358), .ZN(n69) );
  OR3_X1 U354 ( .A1(n345), .A2(n288), .A3(n309), .ZN(n358) );
  XNOR2_X1 U355 ( .A(n359), .B(n360), .ZN(n38) );
  OR2_X1 U356 ( .A1(n359), .A2(n360), .ZN(n37) );
  OAI22_X1 U357 ( .A1(n331), .A2(n326), .B1(n276), .B2(n361), .ZN(n360) );
  XNOR2_X1 U358 ( .A(b[5]), .B(a[3]), .ZN(n331) );
  OAI22_X1 U359 ( .A1(n348), .A2(n347), .B1(n345), .B2(n349), .ZN(n359) );
  XNOR2_X1 U360 ( .A(b[2]), .B(a[7]), .ZN(n349) );
  XNOR2_X1 U361 ( .A(n217), .B(a[7]), .ZN(n348) );
  OAI22_X1 U362 ( .A1(n361), .A2(n326), .B1(n276), .B2(n333), .ZN(n31) );
  XNOR2_X1 U363 ( .A(b[7]), .B(a[3]), .ZN(n333) );
  XNOR2_X1 U364 ( .A(b[6]), .B(a[3]), .ZN(n361) );
  OAI22_X1 U365 ( .A1(n342), .A2(n336), .B1(n334), .B2(n344), .ZN(n21) );
  XNOR2_X1 U366 ( .A(b[7]), .B(a[5]), .ZN(n344) );
  XNOR2_X1 U367 ( .A(n312), .B(a[4]), .ZN(n363) );
  XNOR2_X1 U368 ( .A(b[6]), .B(a[5]), .ZN(n342) );
  OAI22_X1 U369 ( .A1(n353), .A2(n347), .B1(n345), .B2(n355), .ZN(n15) );
  XNOR2_X1 U370 ( .A(b[7]), .B(a[7]), .ZN(n355) );
  NAND2_X1 U371 ( .A1(n345), .A2(n364), .ZN(n347) );
  XNOR2_X1 U372 ( .A(n309), .B(a[6]), .ZN(n364) );
  XNOR2_X1 U373 ( .A(b[6]), .B(a[7]), .ZN(n353) );
  OAI22_X1 U374 ( .A1(n305), .A2(n320), .B1(n365), .B2(n318), .ZN(n104) );
  OAI22_X1 U375 ( .A1(n256), .A2(n320), .B1(n366), .B2(n318), .ZN(n103) );
  XNOR2_X1 U376 ( .A(b[1]), .B(a[1]), .ZN(n365) );
  OAI22_X1 U377 ( .A1(n366), .A2(n320), .B1(n367), .B2(n318), .ZN(n102) );
  XNOR2_X1 U378 ( .A(b[2]), .B(a[1]), .ZN(n366) );
  OAI22_X1 U379 ( .A1(n367), .A2(n320), .B1(n368), .B2(n318), .ZN(n101) );
  OAI22_X1 U380 ( .A1(n368), .A2(n320), .B1(n319), .B2(n318), .ZN(n100) );
  XNOR2_X1 U381 ( .A(b[5]), .B(a[1]), .ZN(n319) );
  NAND2_X1 U382 ( .A1(a[1]), .A2(n318), .ZN(n320) );
  XNOR2_X1 U383 ( .A(b[4]), .B(a[1]), .ZN(n368) );
endmodule


module mac_28 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_28_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_28_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_27_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;
  wire   [15:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .S(SUM[15]) );
  AND2_X2 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n85) );
  CLKBUF_X1 U2 ( .A(B[0]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(n79), .Z(n2) );
  CLKBUF_X1 U4 ( .A(n83), .Z(n3) );
  NAND3_X1 U5 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n4) );
  CLKBUF_X1 U6 ( .A(n35), .Z(n5) );
  CLKBUF_X1 U7 ( .A(n64), .Z(n6) );
  CLKBUF_X1 U8 ( .A(n71), .Z(n7) );
  NAND3_X1 U9 ( .A1(n12), .A2(n13), .A3(n14), .ZN(n8) );
  CLKBUF_X1 U10 ( .A(n4), .Z(n9) );
  NAND2_X1 U11 ( .A1(carry[12]), .A2(A[12]), .ZN(n10) );
  XOR2_X1 U12 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR2_X1 U13 ( .A(n9), .B(n11), .Z(SUM[5]) );
  NAND2_X1 U14 ( .A1(n4), .A2(B[5]), .ZN(n12) );
  NAND2_X1 U15 ( .A1(carry[5]), .A2(A[5]), .ZN(n13) );
  NAND2_X1 U16 ( .A1(B[5]), .A2(A[5]), .ZN(n14) );
  NAND3_X1 U17 ( .A1(n12), .A2(n13), .A3(n14), .ZN(carry[6]) );
  CLKBUF_X1 U18 ( .A(n24), .Z(n15) );
  CLKBUF_X1 U19 ( .A(n20), .Z(n16) );
  CLKBUF_X1 U20 ( .A(n8), .Z(n17) );
  NAND3_X1 U21 ( .A1(n50), .A2(n10), .A3(n52), .ZN(n18) );
  NAND3_X1 U22 ( .A1(n50), .A2(n10), .A3(n52), .ZN(n19) );
  NAND3_X1 U23 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n20) );
  NAND3_X1 U24 ( .A1(n35), .A2(n36), .A3(n37), .ZN(n21) );
  NAND3_X1 U25 ( .A1(n5), .A2(n36), .A3(n37), .ZN(n22) );
  NAND3_X1 U26 ( .A1(n82), .A2(n3), .A3(n84), .ZN(n23) );
  NAND3_X1 U27 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n24) );
  XOR2_X1 U28 ( .A(B[3]), .B(A[3]), .Z(n25) );
  XOR2_X1 U29 ( .A(n23), .B(n25), .Z(SUM[3]) );
  NAND2_X1 U30 ( .A1(carry[3]), .A2(B[3]), .ZN(n26) );
  NAND2_X1 U31 ( .A1(carry[3]), .A2(A[3]), .ZN(n27) );
  NAND2_X1 U32 ( .A1(B[3]), .A2(A[3]), .ZN(n28) );
  NAND3_X1 U33 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[4]) );
  XOR2_X1 U34 ( .A(B[4]), .B(A[4]), .Z(n29) );
  XOR2_X1 U35 ( .A(n15), .B(n29), .Z(SUM[4]) );
  NAND2_X1 U36 ( .A1(n24), .A2(B[4]), .ZN(n30) );
  NAND2_X1 U37 ( .A1(carry[4]), .A2(A[4]), .ZN(n31) );
  NAND2_X1 U38 ( .A1(B[4]), .A2(A[4]), .ZN(n32) );
  NAND3_X1 U39 ( .A1(n30), .A2(n31), .A3(n32), .ZN(carry[5]) );
  NAND3_X1 U40 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n33) );
  XOR2_X1 U41 ( .A(B[6]), .B(A[6]), .Z(n34) );
  XOR2_X1 U42 ( .A(n17), .B(n34), .Z(SUM[6]) );
  NAND2_X1 U43 ( .A1(n8), .A2(B[6]), .ZN(n35) );
  NAND2_X1 U44 ( .A1(carry[6]), .A2(A[6]), .ZN(n36) );
  NAND2_X1 U45 ( .A1(B[6]), .A2(A[6]), .ZN(n37) );
  NAND3_X1 U46 ( .A1(n35), .A2(n36), .A3(n37), .ZN(carry[7]) );
  XOR2_X1 U47 ( .A(B[13]), .B(A[13]), .Z(n38) );
  XOR2_X1 U48 ( .A(n19), .B(n38), .Z(SUM[13]) );
  NAND2_X1 U49 ( .A1(n18), .A2(B[13]), .ZN(n39) );
  NAND2_X1 U50 ( .A1(carry[13]), .A2(A[13]), .ZN(n40) );
  NAND2_X1 U51 ( .A1(B[13]), .A2(A[13]), .ZN(n41) );
  NAND3_X1 U52 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[14]) );
  XOR2_X1 U53 ( .A(B[14]), .B(A[14]), .Z(n42) );
  XOR2_X1 U54 ( .A(n16), .B(n42), .Z(SUM[14]) );
  NAND2_X1 U55 ( .A1(n20), .A2(B[14]), .ZN(n43) );
  NAND2_X1 U56 ( .A1(carry[14]), .A2(A[14]), .ZN(n44) );
  NAND2_X1 U57 ( .A1(B[14]), .A2(A[14]), .ZN(n45) );
  NAND3_X1 U58 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[15]) );
  NAND3_X1 U59 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n46) );
  NAND3_X1 U60 ( .A1(n6), .A2(n65), .A3(n66), .ZN(n47) );
  NAND3_X1 U61 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n48) );
  XOR2_X1 U62 ( .A(B[12]), .B(A[12]), .Z(n49) );
  XOR2_X1 U63 ( .A(n47), .B(n49), .Z(SUM[12]) );
  NAND2_X1 U64 ( .A1(n46), .A2(B[12]), .ZN(n50) );
  NAND2_X1 U65 ( .A1(carry[12]), .A2(A[12]), .ZN(n51) );
  NAND2_X1 U66 ( .A1(B[12]), .A2(A[12]), .ZN(n52) );
  NAND3_X1 U67 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[13]) );
  XOR2_X1 U68 ( .A(B[7]), .B(A[7]), .Z(n53) );
  XOR2_X1 U69 ( .A(n22), .B(n53), .Z(SUM[7]) );
  NAND2_X1 U70 ( .A1(carry[7]), .A2(B[7]), .ZN(n54) );
  NAND2_X1 U71 ( .A1(n21), .A2(A[7]), .ZN(n55) );
  NAND2_X1 U72 ( .A1(B[7]), .A2(A[7]), .ZN(n56) );
  NAND3_X1 U73 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[8]) );
  CLKBUF_X1 U74 ( .A(n33), .Z(n57) );
  NAND3_X1 U75 ( .A1(n74), .A2(n75), .A3(n76), .ZN(n58) );
  XOR2_X1 U76 ( .A(B[10]), .B(A[10]), .Z(n59) );
  XOR2_X1 U77 ( .A(n58), .B(n59), .Z(SUM[10]) );
  NAND2_X1 U78 ( .A1(carry[10]), .A2(B[10]), .ZN(n60) );
  NAND2_X1 U79 ( .A1(carry[10]), .A2(A[10]), .ZN(n61) );
  NAND2_X1 U80 ( .A1(B[10]), .A2(A[10]), .ZN(n62) );
  NAND3_X1 U81 ( .A1(n61), .A2(n60), .A3(n62), .ZN(carry[11]) );
  XOR2_X1 U82 ( .A(B[11]), .B(A[11]), .Z(n63) );
  XOR2_X1 U83 ( .A(n57), .B(n63), .Z(SUM[11]) );
  NAND2_X1 U84 ( .A1(n33), .A2(B[11]), .ZN(n64) );
  NAND2_X1 U85 ( .A1(carry[11]), .A2(A[11]), .ZN(n65) );
  NAND2_X1 U86 ( .A1(B[11]), .A2(A[11]), .ZN(n66) );
  NAND3_X1 U87 ( .A1(n64), .A2(n65), .A3(n66), .ZN(carry[12]) );
  NAND3_X1 U88 ( .A1(n78), .A2(n2), .A3(n80), .ZN(n67) );
  NAND3_X1 U89 ( .A1(n70), .A2(n7), .A3(n72), .ZN(n68) );
  XOR2_X1 U90 ( .A(B[8]), .B(A[8]), .Z(n69) );
  XOR2_X1 U91 ( .A(carry[8]), .B(n69), .Z(SUM[8]) );
  NAND2_X1 U92 ( .A1(n48), .A2(B[8]), .ZN(n70) );
  NAND2_X1 U93 ( .A1(n48), .A2(A[8]), .ZN(n71) );
  NAND2_X1 U94 ( .A1(B[8]), .A2(A[8]), .ZN(n72) );
  NAND3_X1 U95 ( .A1(n70), .A2(n71), .A3(n72), .ZN(carry[9]) );
  XOR2_X1 U96 ( .A(B[9]), .B(A[9]), .Z(n73) );
  XOR2_X1 U97 ( .A(n68), .B(n73), .Z(SUM[9]) );
  NAND2_X1 U98 ( .A1(carry[9]), .A2(B[9]), .ZN(n74) );
  NAND2_X1 U99 ( .A1(carry[9]), .A2(A[9]), .ZN(n75) );
  NAND2_X1 U100 ( .A1(B[9]), .A2(A[9]), .ZN(n76) );
  NAND3_X1 U101 ( .A1(n74), .A2(n75), .A3(n76), .ZN(carry[10]) );
  XOR2_X1 U102 ( .A(B[1]), .B(A[1]), .Z(n77) );
  XOR2_X1 U103 ( .A(n85), .B(n77), .Z(SUM[1]) );
  NAND2_X1 U104 ( .A1(n85), .A2(B[1]), .ZN(n78) );
  NAND2_X1 U105 ( .A1(n85), .A2(A[1]), .ZN(n79) );
  NAND2_X1 U106 ( .A1(B[1]), .A2(A[1]), .ZN(n80) );
  NAND3_X1 U107 ( .A1(n78), .A2(n79), .A3(n80), .ZN(carry[2]) );
  XOR2_X1 U108 ( .A(B[2]), .B(A[2]), .Z(n81) );
  XOR2_X1 U109 ( .A(n67), .B(n81), .Z(SUM[2]) );
  NAND2_X1 U110 ( .A1(carry[2]), .A2(B[2]), .ZN(n82) );
  NAND2_X1 U111 ( .A1(carry[2]), .A2(A[2]), .ZN(n83) );
  NAND2_X1 U112 ( .A1(B[2]), .A2(A[2]), .ZN(n84) );
  NAND3_X1 U113 ( .A1(n82), .A2(n83), .A3(n84), .ZN(carry[3]) );
  XOR2_X1 U114 ( .A(n1), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_27_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18, n19,
         n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76, n77,
         n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94, n95,
         n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369;

  FA_X1 U10 ( .A(n46), .B(n49), .CI(n10), .CO(n9), .S(product[6]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n312), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n311), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n315), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n314), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n317), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n88), .B(n101), .CI(n94), .CO(n53), .S(n54) );
  NAND2_X1 U157 ( .A1(n325), .A2(n363), .ZN(n327) );
  AND2_X1 U158 ( .A1(n95), .A2(n102), .ZN(n206) );
  AND2_X1 U159 ( .A1(n104), .A2(n72), .ZN(n207) );
  NAND2_X1 U160 ( .A1(n263), .A2(n24), .ZN(n208) );
  BUF_X1 U161 ( .A(n245), .Z(n209) );
  CLKBUF_X1 U162 ( .A(b[1]), .Z(n245) );
  CLKBUF_X1 U163 ( .A(b[5]), .Z(n210) );
  CLKBUF_X1 U164 ( .A(b[4]), .Z(n211) );
  XOR2_X1 U165 ( .A(a[3]), .B(a[2]), .Z(n363) );
  XOR2_X1 U166 ( .A(n100), .B(n93), .Z(n212) );
  XOR2_X1 U167 ( .A(n52), .B(n212), .Z(n50) );
  NAND2_X1 U168 ( .A1(n52), .A2(n100), .ZN(n213) );
  NAND2_X1 U169 ( .A1(n52), .A2(n93), .ZN(n214) );
  NAND2_X1 U170 ( .A1(n100), .A2(n93), .ZN(n215) );
  NAND3_X1 U171 ( .A1(n213), .A2(n214), .A3(n215), .ZN(n49) );
  CLKBUF_X1 U172 ( .A(n265), .Z(n216) );
  CLKBUF_X1 U173 ( .A(n208), .Z(n217) );
  CLKBUF_X1 U174 ( .A(n9), .Z(n218) );
  NAND3_X1 U175 ( .A1(n208), .A2(n288), .A3(n290), .ZN(n219) );
  NAND3_X1 U176 ( .A1(n217), .A2(n288), .A3(n290), .ZN(n220) );
  CLKBUF_X1 U177 ( .A(n253), .Z(n221) );
  NAND2_X1 U178 ( .A1(n235), .A2(n19), .ZN(n222) );
  CLKBUF_X1 U179 ( .A(n252), .Z(n223) );
  CLKBUF_X1 U180 ( .A(b[1]), .Z(n224) );
  NAND2_X2 U181 ( .A1(n346), .A2(n365), .ZN(n348) );
  XOR2_X2 U182 ( .A(a[6]), .B(n313), .Z(n346) );
  CLKBUF_X1 U183 ( .A(n293), .Z(n225) );
  XNOR2_X1 U184 ( .A(a[2]), .B(a[1]), .ZN(n325) );
  CLKBUF_X1 U185 ( .A(n236), .Z(n226) );
  INV_X1 U186 ( .A(n307), .ZN(n227) );
  INV_X1 U187 ( .A(n307), .ZN(n228) );
  INV_X1 U188 ( .A(n306), .ZN(n229) );
  INV_X1 U189 ( .A(n307), .ZN(n306) );
  XOR2_X1 U190 ( .A(n95), .B(n102), .Z(n56) );
  CLKBUF_X1 U191 ( .A(n222), .Z(n230) );
  NAND2_X1 U192 ( .A1(a[4]), .A2(a[3]), .ZN(n232) );
  NAND2_X1 U193 ( .A1(n231), .A2(n316), .ZN(n233) );
  NAND2_X2 U194 ( .A1(n232), .A2(n233), .ZN(n335) );
  INV_X1 U195 ( .A(a[4]), .ZN(n231) );
  NAND3_X1 U196 ( .A1(n222), .A2(n304), .A3(n305), .ZN(n234) );
  NAND3_X1 U197 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n235) );
  NAND3_X1 U198 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n236) );
  NAND3_X1 U199 ( .A1(n274), .A2(n273), .A3(n275), .ZN(n237) );
  XOR2_X1 U200 ( .A(n40), .B(n45), .Z(n238) );
  XOR2_X1 U201 ( .A(n218), .B(n238), .Z(product[7]) );
  NAND2_X1 U202 ( .A1(n9), .A2(n40), .ZN(n239) );
  NAND2_X1 U203 ( .A1(n9), .A2(n45), .ZN(n240) );
  NAND2_X1 U204 ( .A1(n40), .A2(n45), .ZN(n241) );
  NAND3_X1 U205 ( .A1(n240), .A2(n239), .A3(n241), .ZN(n8) );
  CLKBUF_X1 U206 ( .A(n235), .Z(n242) );
  CLKBUF_X1 U207 ( .A(n56), .Z(n243) );
  XNOR2_X1 U208 ( .A(n245), .B(a[1]), .ZN(n244) );
  NAND3_X1 U209 ( .A1(n292), .A2(n293), .A3(n294), .ZN(n246) );
  NAND3_X1 U210 ( .A1(n292), .A2(n225), .A3(n294), .ZN(n247) );
  NAND3_X1 U211 ( .A1(n252), .A2(n253), .A3(n251), .ZN(n248) );
  NAND3_X1 U212 ( .A1(n251), .A2(n223), .A3(n221), .ZN(n249) );
  XOR2_X1 U213 ( .A(n54), .B(n206), .Z(n250) );
  XOR2_X1 U214 ( .A(n250), .B(n247), .Z(product[4]) );
  NAND2_X1 U215 ( .A1(n54), .A2(n206), .ZN(n251) );
  NAND2_X1 U216 ( .A1(n12), .A2(n54), .ZN(n252) );
  NAND2_X1 U217 ( .A1(n206), .A2(n246), .ZN(n253) );
  NAND3_X1 U218 ( .A1(n253), .A2(n252), .A3(n251), .ZN(n11) );
  XOR2_X1 U219 ( .A(n50), .B(n53), .Z(n254) );
  XOR2_X1 U220 ( .A(n254), .B(n249), .Z(product[5]) );
  NAND2_X1 U221 ( .A1(n50), .A2(n53), .ZN(n255) );
  NAND2_X1 U222 ( .A1(n248), .A2(n50), .ZN(n256) );
  NAND2_X1 U223 ( .A1(n11), .A2(n53), .ZN(n257) );
  NAND3_X1 U224 ( .A1(n256), .A2(n257), .A3(n255), .ZN(n10) );
  XOR2_X1 U225 ( .A(n20), .B(n23), .Z(n258) );
  XOR2_X1 U226 ( .A(n220), .B(n258), .Z(product[11]) );
  NAND2_X1 U227 ( .A1(n219), .A2(n20), .ZN(n259) );
  NAND2_X1 U228 ( .A1(n5), .A2(n23), .ZN(n260) );
  NAND2_X1 U229 ( .A1(n20), .A2(n23), .ZN(n261) );
  NAND3_X1 U230 ( .A1(n260), .A2(n259), .A3(n261), .ZN(n4) );
  NAND3_X1 U231 ( .A1(n230), .A2(n304), .A3(n305), .ZN(n262) );
  NAND3_X1 U232 ( .A1(n281), .A2(n280), .A3(n282), .ZN(n263) );
  NAND3_X1 U233 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n264) );
  NAND3_X1 U234 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n265) );
  NAND3_X1 U235 ( .A1(n274), .A2(n273), .A3(n275), .ZN(n266) );
  NAND3_X1 U236 ( .A1(n274), .A2(n273), .A3(n275), .ZN(n267) );
  XOR2_X1 U237 ( .A(n34), .B(n39), .Z(n268) );
  XOR2_X1 U238 ( .A(n226), .B(n268), .Z(product[8]) );
  NAND2_X1 U239 ( .A1(n236), .A2(n34), .ZN(n269) );
  NAND2_X1 U240 ( .A1(n8), .A2(n39), .ZN(n270) );
  NAND2_X1 U241 ( .A1(n34), .A2(n39), .ZN(n271) );
  XOR2_X1 U242 ( .A(n308), .B(n17), .Z(n272) );
  XOR2_X1 U243 ( .A(n262), .B(n272), .Z(product[13]) );
  NAND2_X1 U244 ( .A1(n3), .A2(n308), .ZN(n273) );
  NAND2_X1 U245 ( .A1(n234), .A2(n17), .ZN(n274) );
  NAND2_X1 U246 ( .A1(n308), .A2(n17), .ZN(n275) );
  NAND3_X1 U247 ( .A1(n284), .A2(n285), .A3(n286), .ZN(n276) );
  NAND3_X1 U248 ( .A1(n284), .A2(n285), .A3(n286), .ZN(n277) );
  CLKBUF_X1 U249 ( .A(n263), .Z(n278) );
  XOR2_X1 U250 ( .A(n33), .B(n28), .Z(n279) );
  XOR2_X1 U251 ( .A(n216), .B(n279), .Z(product[9]) );
  NAND2_X1 U252 ( .A1(n264), .A2(n33), .ZN(n280) );
  NAND2_X1 U253 ( .A1(n265), .A2(n28), .ZN(n281) );
  NAND2_X1 U254 ( .A1(n33), .A2(n28), .ZN(n282) );
  NAND3_X1 U255 ( .A1(n281), .A2(n280), .A3(n282), .ZN(n6) );
  XOR2_X1 U256 ( .A(n103), .B(n96), .Z(n283) );
  XOR2_X1 U257 ( .A(n207), .B(n283), .Z(product[2]) );
  NAND2_X1 U258 ( .A1(n207), .A2(n103), .ZN(n284) );
  NAND2_X1 U259 ( .A1(n14), .A2(n96), .ZN(n285) );
  NAND2_X1 U260 ( .A1(n103), .A2(n96), .ZN(n286) );
  NAND3_X1 U261 ( .A1(n284), .A2(n285), .A3(n286), .ZN(n13) );
  XOR2_X1 U262 ( .A(n27), .B(n24), .Z(n287) );
  XOR2_X1 U263 ( .A(n278), .B(n287), .Z(product[10]) );
  NAND2_X1 U264 ( .A1(n6), .A2(n27), .ZN(n288) );
  NAND2_X1 U265 ( .A1(n263), .A2(n24), .ZN(n289) );
  NAND2_X1 U266 ( .A1(n27), .A2(n24), .ZN(n290) );
  NAND3_X1 U267 ( .A1(n289), .A2(n288), .A3(n290), .ZN(n5) );
  XOR2_X1 U268 ( .A(n243), .B(n71), .Z(n291) );
  XOR2_X1 U269 ( .A(n277), .B(n291), .Z(product[3]) );
  NAND2_X1 U270 ( .A1(n276), .A2(n56), .ZN(n292) );
  NAND2_X1 U271 ( .A1(n13), .A2(n71), .ZN(n293) );
  NAND2_X1 U272 ( .A1(n56), .A2(n71), .ZN(n294) );
  NAND3_X1 U273 ( .A1(n292), .A2(n293), .A3(n294), .ZN(n12) );
  NAND2_X2 U274 ( .A1(n335), .A2(n364), .ZN(n337) );
  XOR2_X1 U275 ( .A(a[2]), .B(n318), .Z(n295) );
  XOR2_X1 U276 ( .A(a[2]), .B(n318), .Z(n296) );
  INV_X1 U277 ( .A(n15), .ZN(n308) );
  XNOR2_X1 U278 ( .A(n242), .B(n297), .ZN(product[12]) );
  XNOR2_X1 U279 ( .A(n19), .B(n18), .ZN(n297) );
  XNOR2_X1 U280 ( .A(n267), .B(n298), .ZN(product[14]) );
  XNOR2_X1 U281 ( .A(n309), .B(n15), .ZN(n298) );
  AND3_X1 U282 ( .A1(n301), .A2(n300), .A3(n302), .ZN(product[15]) );
  OAI22_X1 U283 ( .A1(n354), .A2(n348), .B1(n346), .B2(n356), .ZN(n15) );
  INV_X1 U284 ( .A(n333), .ZN(n315) );
  INV_X1 U285 ( .A(n344), .ZN(n312) );
  INV_X1 U286 ( .A(n21), .ZN(n311) );
  INV_X1 U287 ( .A(n324), .ZN(n317) );
  INV_X1 U288 ( .A(b[0]), .ZN(n307) );
  INV_X1 U289 ( .A(n31), .ZN(n314) );
  INV_X1 U290 ( .A(a[0]), .ZN(n319) );
  INV_X1 U291 ( .A(a[5]), .ZN(n313) );
  INV_X1 U292 ( .A(a[7]), .ZN(n310) );
  NAND2_X1 U293 ( .A1(n266), .A2(n309), .ZN(n300) );
  NAND2_X1 U294 ( .A1(n237), .A2(n15), .ZN(n301) );
  NAND2_X1 U295 ( .A1(n309), .A2(n15), .ZN(n302) );
  NAND2_X1 U296 ( .A1(n235), .A2(n19), .ZN(n303) );
  NAND2_X1 U297 ( .A1(n4), .A2(n18), .ZN(n304) );
  NAND2_X1 U298 ( .A1(n19), .A2(n18), .ZN(n305) );
  NAND3_X1 U299 ( .A1(n304), .A2(n303), .A3(n305), .ZN(n3) );
  INV_X1 U300 ( .A(n355), .ZN(n309) );
  INV_X1 U301 ( .A(a[3]), .ZN(n316) );
  INV_X1 U302 ( .A(a[1]), .ZN(n318) );
  NOR2_X1 U303 ( .A1(n319), .A2(n229), .ZN(product[0]) );
  OAI22_X1 U304 ( .A1(n320), .A2(n321), .B1(n322), .B2(n319), .ZN(n99) );
  OAI22_X1 U305 ( .A1(n322), .A2(n321), .B1(n323), .B2(n319), .ZN(n98) );
  XNOR2_X1 U306 ( .A(b[6]), .B(a[1]), .ZN(n322) );
  OAI22_X1 U307 ( .A1(n319), .A2(n323), .B1(n321), .B2(n323), .ZN(n324) );
  XNOR2_X1 U308 ( .A(b[7]), .B(a[1]), .ZN(n323) );
  NOR2_X1 U309 ( .A1(n295), .A2(n229), .ZN(n96) );
  OAI22_X1 U310 ( .A1(n326), .A2(n327), .B1(n296), .B2(n328), .ZN(n95) );
  XNOR2_X1 U311 ( .A(a[3]), .B(n228), .ZN(n326) );
  OAI22_X1 U312 ( .A1(n328), .A2(n327), .B1(n296), .B2(n329), .ZN(n94) );
  XNOR2_X1 U313 ( .A(n224), .B(a[3]), .ZN(n328) );
  OAI22_X1 U314 ( .A1(n329), .A2(n327), .B1(n295), .B2(n330), .ZN(n93) );
  XNOR2_X1 U315 ( .A(b[2]), .B(a[3]), .ZN(n329) );
  OAI22_X1 U316 ( .A1(n330), .A2(n327), .B1(n296), .B2(n331), .ZN(n92) );
  XNOR2_X1 U317 ( .A(b[3]), .B(a[3]), .ZN(n330) );
  OAI22_X1 U318 ( .A1(n331), .A2(n327), .B1(n296), .B2(n332), .ZN(n91) );
  XNOR2_X1 U319 ( .A(b[4]), .B(a[3]), .ZN(n331) );
  OAI22_X1 U320 ( .A1(n334), .A2(n295), .B1(n327), .B2(n334), .ZN(n333) );
  NOR2_X1 U321 ( .A1(n335), .A2(n229), .ZN(n88) );
  OAI22_X1 U322 ( .A1(n336), .A2(n337), .B1(n335), .B2(n338), .ZN(n87) );
  XNOR2_X1 U323 ( .A(a[5]), .B(n227), .ZN(n336) );
  OAI22_X1 U324 ( .A1(n338), .A2(n337), .B1(n335), .B2(n339), .ZN(n86) );
  XNOR2_X1 U325 ( .A(n209), .B(a[5]), .ZN(n338) );
  OAI22_X1 U326 ( .A1(n339), .A2(n337), .B1(n335), .B2(n340), .ZN(n85) );
  XNOR2_X1 U327 ( .A(b[2]), .B(a[5]), .ZN(n339) );
  OAI22_X1 U328 ( .A1(n340), .A2(n337), .B1(n335), .B2(n341), .ZN(n84) );
  XNOR2_X1 U329 ( .A(b[3]), .B(a[5]), .ZN(n340) );
  OAI22_X1 U330 ( .A1(n341), .A2(n337), .B1(n335), .B2(n342), .ZN(n83) );
  XNOR2_X1 U331 ( .A(n211), .B(a[5]), .ZN(n341) );
  OAI22_X1 U332 ( .A1(n342), .A2(n337), .B1(n335), .B2(n343), .ZN(n82) );
  XNOR2_X1 U333 ( .A(n210), .B(a[5]), .ZN(n342) );
  OAI22_X1 U334 ( .A1(n345), .A2(n335), .B1(n337), .B2(n345), .ZN(n344) );
  NOR2_X1 U335 ( .A1(n346), .A2(n229), .ZN(n80) );
  OAI22_X1 U336 ( .A1(n347), .A2(n348), .B1(n346), .B2(n349), .ZN(n79) );
  XNOR2_X1 U337 ( .A(a[7]), .B(n227), .ZN(n347) );
  OAI22_X1 U338 ( .A1(n350), .A2(n348), .B1(n346), .B2(n351), .ZN(n77) );
  OAI22_X1 U339 ( .A1(n351), .A2(n348), .B1(n346), .B2(n352), .ZN(n76) );
  XNOR2_X1 U340 ( .A(b[3]), .B(a[7]), .ZN(n351) );
  OAI22_X1 U341 ( .A1(n352), .A2(n348), .B1(n346), .B2(n353), .ZN(n75) );
  XNOR2_X1 U342 ( .A(n211), .B(a[7]), .ZN(n352) );
  OAI22_X1 U343 ( .A1(n353), .A2(n348), .B1(n346), .B2(n354), .ZN(n74) );
  XNOR2_X1 U344 ( .A(n210), .B(a[7]), .ZN(n353) );
  OAI22_X1 U345 ( .A1(n356), .A2(n346), .B1(n348), .B2(n356), .ZN(n355) );
  OAI21_X1 U346 ( .B1(n306), .B2(n318), .A(n321), .ZN(n72) );
  OAI21_X1 U347 ( .B1(n316), .B2(n327), .A(n357), .ZN(n71) );
  OR3_X1 U348 ( .A1(n295), .A2(n228), .A3(n316), .ZN(n357) );
  OAI21_X1 U349 ( .B1(n313), .B2(n337), .A(n358), .ZN(n70) );
  OR3_X1 U350 ( .A1(n335), .A2(n306), .A3(n313), .ZN(n358) );
  OAI21_X1 U351 ( .B1(n310), .B2(n348), .A(n359), .ZN(n69) );
  OR3_X1 U352 ( .A1(n346), .A2(n228), .A3(n310), .ZN(n359) );
  XNOR2_X1 U353 ( .A(n360), .B(n361), .ZN(n38) );
  OR2_X1 U354 ( .A1(n360), .A2(n361), .ZN(n37) );
  OAI22_X1 U355 ( .A1(n332), .A2(n327), .B1(n295), .B2(n362), .ZN(n361) );
  XNOR2_X1 U356 ( .A(n210), .B(a[3]), .ZN(n332) );
  OAI22_X1 U357 ( .A1(n349), .A2(n348), .B1(n346), .B2(n350), .ZN(n360) );
  XNOR2_X1 U358 ( .A(b[2]), .B(a[7]), .ZN(n350) );
  XNOR2_X1 U359 ( .A(n209), .B(a[7]), .ZN(n349) );
  OAI22_X1 U360 ( .A1(n362), .A2(n327), .B1(n296), .B2(n334), .ZN(n31) );
  XNOR2_X1 U361 ( .A(b[7]), .B(a[3]), .ZN(n334) );
  XNOR2_X1 U362 ( .A(b[6]), .B(a[3]), .ZN(n362) );
  OAI22_X1 U363 ( .A1(n343), .A2(n337), .B1(n335), .B2(n345), .ZN(n21) );
  XNOR2_X1 U364 ( .A(b[7]), .B(a[5]), .ZN(n345) );
  XNOR2_X1 U365 ( .A(n313), .B(a[4]), .ZN(n364) );
  XNOR2_X1 U366 ( .A(b[6]), .B(a[5]), .ZN(n343) );
  XNOR2_X1 U367 ( .A(b[7]), .B(a[7]), .ZN(n356) );
  XNOR2_X1 U368 ( .A(n310), .B(a[6]), .ZN(n365) );
  XNOR2_X1 U369 ( .A(b[6]), .B(a[7]), .ZN(n354) );
  OAI22_X1 U370 ( .A1(n227), .A2(n321), .B1(n366), .B2(n319), .ZN(n104) );
  OAI22_X1 U371 ( .A1(n244), .A2(n321), .B1(n367), .B2(n319), .ZN(n103) );
  XNOR2_X1 U372 ( .A(b[1]), .B(a[1]), .ZN(n366) );
  OAI22_X1 U373 ( .A1(n367), .A2(n321), .B1(n368), .B2(n319), .ZN(n102) );
  XNOR2_X1 U374 ( .A(b[2]), .B(a[1]), .ZN(n367) );
  OAI22_X1 U375 ( .A1(n368), .A2(n321), .B1(n369), .B2(n319), .ZN(n101) );
  XNOR2_X1 U376 ( .A(b[3]), .B(a[1]), .ZN(n368) );
  OAI22_X1 U377 ( .A1(n369), .A2(n321), .B1(n320), .B2(n319), .ZN(n100) );
  XNOR2_X1 U378 ( .A(b[5]), .B(a[1]), .ZN(n320) );
  NAND2_X1 U379 ( .A1(a[1]), .A2(n319), .ZN(n321) );
  XNOR2_X1 U380 ( .A(b[4]), .B(a[1]), .ZN(n369) );
endmodule


module mac_27 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_27_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_27_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X2 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_26_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;
  wire   [15:1] carry;

  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n71) );
  NAND3_X1 U2 ( .A1(n68), .A2(n69), .A3(n70), .ZN(n1) );
  NAND3_X1 U3 ( .A1(n68), .A2(n69), .A3(n70), .ZN(n2) );
  XOR2_X1 U4 ( .A(B[15]), .B(A[15]), .Z(n3) );
  XOR2_X1 U5 ( .A(carry[15]), .B(n3), .Z(SUM[15]) );
  NAND3_X1 U6 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n4) );
  NAND3_X1 U7 ( .A1(n8), .A2(n9), .A3(n10), .ZN(n5) );
  NAND3_X1 U8 ( .A1(n8), .A2(n9), .A3(n10), .ZN(n6) );
  XOR2_X1 U9 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR2_X1 U10 ( .A(carry[3]), .B(n7), .Z(SUM[3]) );
  NAND2_X1 U11 ( .A1(carry[3]), .A2(B[3]), .ZN(n8) );
  NAND2_X1 U12 ( .A1(carry[3]), .A2(A[3]), .ZN(n9) );
  NAND2_X1 U13 ( .A1(B[3]), .A2(A[3]), .ZN(n10) );
  NAND3_X1 U14 ( .A1(n8), .A2(n9), .A3(n10), .ZN(carry[4]) );
  NAND3_X1 U15 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n11) );
  NAND3_X1 U16 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n12) );
  NAND3_X1 U17 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n13) );
  NAND3_X1 U18 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n14) );
  NAND3_X1 U19 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n15) );
  NAND3_X1 U20 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n16) );
  XOR2_X1 U21 ( .A(B[4]), .B(A[4]), .Z(n17) );
  XOR2_X1 U22 ( .A(n6), .B(n17), .Z(SUM[4]) );
  NAND2_X1 U23 ( .A1(n5), .A2(B[4]), .ZN(n18) );
  NAND2_X1 U24 ( .A1(carry[4]), .A2(A[4]), .ZN(n19) );
  NAND2_X1 U25 ( .A1(B[4]), .A2(A[4]), .ZN(n20) );
  NAND3_X1 U26 ( .A1(n18), .A2(n19), .A3(n20), .ZN(carry[5]) );
  XOR2_X1 U27 ( .A(B[10]), .B(A[10]), .Z(n21) );
  XOR2_X1 U28 ( .A(n12), .B(n21), .Z(SUM[10]) );
  NAND2_X1 U29 ( .A1(n11), .A2(B[10]), .ZN(n22) );
  NAND2_X1 U30 ( .A1(carry[10]), .A2(A[10]), .ZN(n23) );
  NAND2_X1 U31 ( .A1(B[10]), .A2(A[10]), .ZN(n24) );
  NAND3_X1 U32 ( .A1(n22), .A2(n23), .A3(n24), .ZN(carry[11]) );
  NAND3_X1 U33 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n25) );
  NAND3_X1 U34 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n26) );
  NAND3_X1 U35 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n27) );
  NAND3_X1 U36 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n28) );
  XOR2_X1 U37 ( .A(B[11]), .B(A[11]), .Z(n29) );
  XOR2_X1 U38 ( .A(n14), .B(n29), .Z(SUM[11]) );
  NAND2_X1 U39 ( .A1(n13), .A2(B[11]), .ZN(n30) );
  NAND2_X1 U40 ( .A1(carry[11]), .A2(A[11]), .ZN(n31) );
  NAND2_X1 U41 ( .A1(B[11]), .A2(A[11]), .ZN(n32) );
  NAND3_X1 U42 ( .A1(n31), .A2(n30), .A3(n32), .ZN(carry[12]) );
  XOR2_X1 U43 ( .A(B[5]), .B(A[5]), .Z(n33) );
  XOR2_X1 U44 ( .A(n16), .B(n33), .Z(SUM[5]) );
  NAND2_X1 U45 ( .A1(n15), .A2(B[5]), .ZN(n34) );
  NAND2_X1 U46 ( .A1(carry[5]), .A2(A[5]), .ZN(n35) );
  NAND2_X1 U47 ( .A1(B[5]), .A2(A[5]), .ZN(n36) );
  NAND3_X1 U48 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[6]) );
  XOR2_X1 U49 ( .A(B[12]), .B(A[12]), .Z(n37) );
  XOR2_X1 U50 ( .A(n25), .B(n37), .Z(SUM[12]) );
  NAND2_X1 U51 ( .A1(n25), .A2(B[12]), .ZN(n38) );
  NAND2_X1 U52 ( .A1(carry[12]), .A2(A[12]), .ZN(n39) );
  NAND2_X1 U53 ( .A1(B[12]), .A2(A[12]), .ZN(n40) );
  NAND3_X1 U54 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[13]) );
  NAND3_X1 U55 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n41) );
  XOR2_X1 U56 ( .A(B[9]), .B(A[9]), .Z(n42) );
  XOR2_X1 U57 ( .A(carry[9]), .B(n42), .Z(SUM[9]) );
  NAND2_X1 U58 ( .A1(n41), .A2(B[9]), .ZN(n43) );
  NAND2_X1 U59 ( .A1(n41), .A2(A[9]), .ZN(n44) );
  NAND2_X1 U60 ( .A1(B[9]), .A2(A[9]), .ZN(n45) );
  NAND3_X1 U61 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[10]) );
  NAND3_X1 U62 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n46) );
  XOR2_X1 U63 ( .A(B[8]), .B(A[8]), .Z(n47) );
  XOR2_X1 U64 ( .A(carry[8]), .B(n47), .Z(SUM[8]) );
  NAND2_X1 U65 ( .A1(n2), .A2(B[8]), .ZN(n48) );
  NAND2_X1 U66 ( .A1(n1), .A2(A[8]), .ZN(n49) );
  NAND2_X1 U67 ( .A1(B[8]), .A2(A[8]), .ZN(n50) );
  NAND3_X1 U68 ( .A1(n48), .A2(n49), .A3(n50), .ZN(carry[9]) );
  XOR2_X1 U69 ( .A(B[1]), .B(A[1]), .Z(n51) );
  XOR2_X1 U70 ( .A(n71), .B(n51), .Z(SUM[1]) );
  NAND2_X1 U71 ( .A1(n71), .A2(B[1]), .ZN(n52) );
  NAND2_X1 U72 ( .A1(n71), .A2(A[1]), .ZN(n53) );
  NAND2_X1 U73 ( .A1(B[1]), .A2(A[1]), .ZN(n54) );
  NAND3_X1 U74 ( .A1(n52), .A2(n53), .A3(n54), .ZN(carry[2]) );
  XOR2_X1 U75 ( .A(B[13]), .B(A[13]), .Z(n55) );
  XOR2_X1 U76 ( .A(n26), .B(n55), .Z(SUM[13]) );
  NAND2_X1 U77 ( .A1(n26), .A2(B[13]), .ZN(n56) );
  NAND2_X1 U78 ( .A1(carry[13]), .A2(A[13]), .ZN(n57) );
  NAND2_X1 U79 ( .A1(B[13]), .A2(A[13]), .ZN(n58) );
  NAND3_X1 U80 ( .A1(n56), .A2(n57), .A3(n58), .ZN(carry[14]) );
  XOR2_X1 U81 ( .A(B[6]), .B(A[6]), .Z(n59) );
  XOR2_X1 U82 ( .A(n27), .B(n59), .Z(SUM[6]) );
  NAND2_X1 U83 ( .A1(n4), .A2(B[6]), .ZN(n60) );
  NAND2_X1 U84 ( .A1(carry[6]), .A2(A[6]), .ZN(n61) );
  NAND2_X1 U85 ( .A1(B[6]), .A2(A[6]), .ZN(n62) );
  NAND3_X1 U86 ( .A1(n61), .A2(n60), .A3(n62), .ZN(carry[7]) );
  XOR2_X1 U87 ( .A(B[14]), .B(A[14]), .Z(n63) );
  XOR2_X1 U88 ( .A(carry[14]), .B(n63), .Z(SUM[14]) );
  NAND2_X1 U89 ( .A1(carry[14]), .A2(B[14]), .ZN(n64) );
  NAND2_X1 U90 ( .A1(n46), .A2(A[14]), .ZN(n65) );
  NAND2_X1 U91 ( .A1(B[14]), .A2(A[14]), .ZN(n66) );
  NAND3_X1 U92 ( .A1(n64), .A2(n65), .A3(n66), .ZN(carry[15]) );
  XOR2_X1 U93 ( .A(B[7]), .B(A[7]), .Z(n67) );
  XOR2_X1 U94 ( .A(n28), .B(n67), .Z(SUM[7]) );
  NAND2_X1 U95 ( .A1(n28), .A2(B[7]), .ZN(n68) );
  NAND2_X1 U96 ( .A1(carry[7]), .A2(A[7]), .ZN(n69) );
  NAND2_X1 U97 ( .A1(B[7]), .A2(A[7]), .ZN(n70) );
  NAND3_X1 U98 ( .A1(n68), .A2(n69), .A3(n70), .ZN(carry[8]) );
  XOR2_X1 U99 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_26_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n317), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n316), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n320), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n319), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n322), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n88), .B(n101), .CI(n94), .CO(n53), .S(n54) );
  XOR2_X2 U157 ( .A(a[2]), .B(n323), .Z(n294) );
  OR3_X1 U158 ( .A1(n249), .A2(n311), .A3(n318), .ZN(n363) );
  NAND2_X1 U159 ( .A1(n330), .A2(n368), .ZN(n332) );
  NAND2_X1 U160 ( .A1(n340), .A2(n369), .ZN(n342) );
  AND2_X1 U161 ( .A1(n95), .A2(n102), .ZN(n206) );
  AND3_X1 U162 ( .A1(n223), .A2(n222), .A3(n224), .ZN(product[15]) );
  CLKBUF_X1 U163 ( .A(b[1]), .Z(n208) );
  XOR2_X1 U164 ( .A(n52), .B(n210), .Z(n50) );
  XOR2_X1 U165 ( .A(a[3]), .B(a[2]), .Z(n368) );
  CLKBUF_X1 U166 ( .A(b[3]), .Z(n209) );
  XOR2_X1 U167 ( .A(n100), .B(n93), .Z(n210) );
  NAND2_X1 U168 ( .A1(n52), .A2(n100), .ZN(n211) );
  NAND2_X1 U169 ( .A1(n52), .A2(n93), .ZN(n212) );
  NAND2_X1 U170 ( .A1(n100), .A2(n93), .ZN(n213) );
  NAND3_X1 U171 ( .A1(n211), .A2(n212), .A3(n213), .ZN(n49) );
  OR2_X1 U172 ( .A1(n341), .A2(n342), .ZN(n214) );
  OR2_X1 U173 ( .A1(n249), .A2(n343), .ZN(n215) );
  NAND2_X1 U174 ( .A1(n214), .A2(n215), .ZN(n87) );
  CLKBUF_X1 U175 ( .A(n56), .Z(n216) );
  CLKBUF_X1 U176 ( .A(b[1]), .Z(n217) );
  NAND2_X1 U177 ( .A1(n103), .A2(n14), .ZN(n218) );
  NAND3_X1 U178 ( .A1(n301), .A2(n300), .A3(n302), .ZN(n219) );
  NAND3_X1 U179 ( .A1(n301), .A2(n300), .A3(n302), .ZN(n220) );
  XOR2_X1 U180 ( .A(n314), .B(n15), .Z(n221) );
  XOR2_X1 U181 ( .A(n220), .B(n221), .Z(product[14]) );
  NAND2_X1 U182 ( .A1(n219), .A2(n314), .ZN(n222) );
  NAND2_X1 U183 ( .A1(n2), .A2(n15), .ZN(n223) );
  NAND2_X1 U184 ( .A1(n314), .A2(n15), .ZN(n224) );
  NAND2_X1 U185 ( .A1(n237), .A2(n20), .ZN(n225) );
  CLKBUF_X1 U186 ( .A(n218), .Z(n226) );
  AND2_X1 U187 ( .A1(n104), .A2(n72), .ZN(n227) );
  CLKBUF_X1 U188 ( .A(n251), .Z(n228) );
  NAND2_X1 U189 ( .A1(n257), .A2(n33), .ZN(n229) );
  CLKBUF_X1 U190 ( .A(n257), .Z(n230) );
  CLKBUF_X1 U191 ( .A(n225), .Z(n231) );
  NAND3_X1 U192 ( .A1(n256), .A2(n255), .A3(n254), .ZN(n232) );
  NAND3_X1 U193 ( .A1(n304), .A2(n305), .A3(n306), .ZN(n233) );
  CLKBUF_X1 U194 ( .A(n227), .Z(n234) );
  NAND2_X2 U195 ( .A1(n351), .A2(n370), .ZN(n353) );
  XOR2_X2 U196 ( .A(a[6]), .B(n318), .Z(n351) );
  NAND3_X1 U197 ( .A1(n298), .A2(n297), .A3(n296), .ZN(n235) );
  CLKBUF_X1 U198 ( .A(n229), .Z(n236) );
  NAND3_X1 U199 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n237) );
  NAND3_X1 U200 ( .A1(n266), .A2(n267), .A3(n265), .ZN(n238) );
  CLKBUF_X1 U201 ( .A(n309), .Z(n239) );
  CLKBUF_X1 U202 ( .A(n237), .Z(n240) );
  NAND3_X1 U203 ( .A1(n229), .A2(n277), .A3(n278), .ZN(n241) );
  NAND3_X1 U204 ( .A1(n236), .A2(n277), .A3(n278), .ZN(n242) );
  NAND3_X1 U205 ( .A1(n218), .A2(n263), .A3(n261), .ZN(n243) );
  NAND3_X1 U206 ( .A1(n261), .A2(n226), .A3(n263), .ZN(n244) );
  XOR2_X1 U207 ( .A(n27), .B(n24), .Z(n245) );
  XOR2_X1 U208 ( .A(n242), .B(n245), .Z(product[10]) );
  NAND2_X1 U209 ( .A1(n241), .A2(n27), .ZN(n246) );
  NAND2_X1 U210 ( .A1(n6), .A2(n24), .ZN(n247) );
  NAND2_X1 U211 ( .A1(n27), .A2(n24), .ZN(n248) );
  NAND3_X1 U212 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n5) );
  XNOR2_X1 U213 ( .A(a[4]), .B(a[3]), .ZN(n249) );
  XNOR2_X1 U214 ( .A(a[4]), .B(a[3]), .ZN(n340) );
  CLKBUF_X1 U215 ( .A(n232), .Z(n250) );
  NAND3_X1 U216 ( .A1(n280), .A2(n282), .A3(n281), .ZN(n251) );
  CLKBUF_X1 U217 ( .A(n12), .Z(n252) );
  XOR2_X1 U218 ( .A(n252), .B(n206), .Z(n253) );
  XOR2_X1 U219 ( .A(n54), .B(n253), .Z(product[4]) );
  NAND2_X1 U220 ( .A1(n54), .A2(n238), .ZN(n254) );
  NAND2_X1 U221 ( .A1(n54), .A2(n206), .ZN(n255) );
  NAND2_X1 U222 ( .A1(n12), .A2(n206), .ZN(n256) );
  NAND3_X1 U223 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n11) );
  NAND3_X1 U224 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n257) );
  NAND3_X1 U225 ( .A1(n309), .A2(n308), .A3(n310), .ZN(n258) );
  NAND3_X1 U226 ( .A1(n308), .A2(n239), .A3(n310), .ZN(n259) );
  XOR2_X1 U227 ( .A(n103), .B(n96), .Z(n260) );
  XOR2_X1 U228 ( .A(n260), .B(n234), .Z(product[2]) );
  NAND2_X1 U229 ( .A1(n103), .A2(n96), .ZN(n261) );
  NAND2_X1 U230 ( .A1(n103), .A2(n14), .ZN(n262) );
  NAND2_X1 U231 ( .A1(n96), .A2(n227), .ZN(n263) );
  NAND3_X1 U232 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n13) );
  XOR2_X1 U233 ( .A(n216), .B(n71), .Z(n264) );
  XOR2_X1 U234 ( .A(n264), .B(n244), .Z(product[3]) );
  NAND2_X1 U235 ( .A1(n56), .A2(n71), .ZN(n265) );
  NAND2_X1 U236 ( .A1(n56), .A2(n243), .ZN(n266) );
  NAND2_X1 U237 ( .A1(n71), .A2(n13), .ZN(n267) );
  NAND3_X1 U238 ( .A1(n266), .A2(n267), .A3(n265), .ZN(n12) );
  XOR2_X1 U239 ( .A(n34), .B(n39), .Z(n268) );
  XOR2_X1 U240 ( .A(n259), .B(n268), .Z(product[8]) );
  NAND2_X1 U241 ( .A1(n258), .A2(n34), .ZN(n269) );
  NAND2_X1 U242 ( .A1(n8), .A2(n39), .ZN(n270) );
  NAND2_X1 U243 ( .A1(n34), .A2(n39), .ZN(n271) );
  NAND3_X1 U244 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n7) );
  NAND3_X1 U245 ( .A1(n280), .A2(n281), .A3(n282), .ZN(n272) );
  NAND3_X1 U246 ( .A1(n286), .A2(n287), .A3(n288), .ZN(n273) );
  NAND3_X1 U247 ( .A1(n231), .A2(n287), .A3(n288), .ZN(n274) );
  XOR2_X1 U248 ( .A(n33), .B(n28), .Z(n275) );
  XOR2_X1 U249 ( .A(n230), .B(n275), .Z(product[9]) );
  NAND2_X1 U250 ( .A1(n257), .A2(n33), .ZN(n276) );
  NAND2_X1 U251 ( .A1(n7), .A2(n28), .ZN(n277) );
  NAND2_X1 U252 ( .A1(n33), .A2(n28), .ZN(n278) );
  NAND3_X1 U253 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n6) );
  XOR2_X1 U254 ( .A(n50), .B(n53), .Z(n279) );
  XOR2_X1 U255 ( .A(n250), .B(n279), .Z(product[5]) );
  NAND2_X1 U256 ( .A1(n232), .A2(n50), .ZN(n280) );
  NAND2_X1 U257 ( .A1(n11), .A2(n53), .ZN(n281) );
  NAND2_X1 U258 ( .A1(n50), .A2(n53), .ZN(n282) );
  CLKBUF_X1 U259 ( .A(n9), .Z(n283) );
  INV_X1 U260 ( .A(n312), .ZN(n284) );
  INV_X1 U261 ( .A(n312), .ZN(n311) );
  XNOR2_X1 U262 ( .A(a[2]), .B(a[1]), .ZN(n330) );
  XOR2_X1 U263 ( .A(n20), .B(n23), .Z(n285) );
  XOR2_X1 U264 ( .A(n240), .B(n285), .Z(product[11]) );
  NAND2_X1 U265 ( .A1(n237), .A2(n20), .ZN(n286) );
  NAND2_X1 U266 ( .A1(n5), .A2(n23), .ZN(n287) );
  NAND2_X1 U267 ( .A1(n20), .A2(n23), .ZN(n288) );
  NAND3_X1 U268 ( .A1(n225), .A2(n287), .A3(n288), .ZN(n4) );
  XOR2_X1 U269 ( .A(n102), .B(n95), .Z(n56) );
  NAND2_X1 U270 ( .A1(b[1]), .A2(a[1]), .ZN(n291) );
  NAND2_X1 U271 ( .A1(n289), .A2(n290), .ZN(n292) );
  NAND2_X1 U272 ( .A1(n291), .A2(n292), .ZN(n371) );
  INV_X1 U273 ( .A(b[1]), .ZN(n289) );
  INV_X1 U274 ( .A(a[1]), .ZN(n290) );
  XOR2_X1 U275 ( .A(a[2]), .B(n323), .Z(n293) );
  XOR2_X1 U276 ( .A(n283), .B(n307), .Z(product[7]) );
  INV_X1 U277 ( .A(n15), .ZN(n313) );
  INV_X1 U278 ( .A(n349), .ZN(n317) );
  INV_X1 U279 ( .A(n21), .ZN(n316) );
  INV_X1 U280 ( .A(n329), .ZN(n322) );
  INV_X1 U281 ( .A(n338), .ZN(n320) );
  INV_X1 U282 ( .A(b[0]), .ZN(n312) );
  INV_X1 U283 ( .A(n360), .ZN(n314) );
  INV_X1 U284 ( .A(n31), .ZN(n319) );
  INV_X1 U285 ( .A(a[0]), .ZN(n324) );
  INV_X1 U286 ( .A(a[5]), .ZN(n318) );
  INV_X1 U287 ( .A(a[7]), .ZN(n315) );
  XOR2_X1 U288 ( .A(n19), .B(n18), .Z(n295) );
  XOR2_X1 U289 ( .A(n295), .B(n274), .Z(product[12]) );
  NAND2_X1 U290 ( .A1(n19), .A2(n18), .ZN(n296) );
  NAND2_X1 U291 ( .A1(n19), .A2(n273), .ZN(n297) );
  NAND2_X1 U292 ( .A1(n18), .A2(n4), .ZN(n298) );
  NAND3_X1 U293 ( .A1(n298), .A2(n296), .A3(n297), .ZN(n3) );
  XOR2_X1 U294 ( .A(n17), .B(n313), .Z(n299) );
  XOR2_X1 U295 ( .A(n299), .B(n235), .Z(product[13]) );
  NAND2_X1 U296 ( .A1(n17), .A2(n313), .ZN(n300) );
  NAND2_X1 U297 ( .A1(n17), .A2(n235), .ZN(n301) );
  NAND2_X1 U298 ( .A1(n313), .A2(n3), .ZN(n302) );
  NAND3_X1 U299 ( .A1(n300), .A2(n301), .A3(n302), .ZN(n2) );
  INV_X1 U300 ( .A(a[3]), .ZN(n321) );
  XOR2_X1 U301 ( .A(n46), .B(n49), .Z(n303) );
  XOR2_X1 U302 ( .A(n228), .B(n303), .Z(product[6]) );
  NAND2_X1 U303 ( .A1(n251), .A2(n46), .ZN(n304) );
  NAND2_X1 U304 ( .A1(n272), .A2(n49), .ZN(n305) );
  NAND2_X1 U305 ( .A1(n46), .A2(n49), .ZN(n306) );
  NAND3_X1 U306 ( .A1(n304), .A2(n305), .A3(n306), .ZN(n9) );
  XOR2_X1 U307 ( .A(n40), .B(n45), .Z(n307) );
  NAND2_X1 U308 ( .A1(n233), .A2(n40), .ZN(n308) );
  NAND2_X1 U309 ( .A1(n9), .A2(n45), .ZN(n309) );
  NAND2_X1 U310 ( .A1(n40), .A2(n45), .ZN(n310) );
  NAND3_X1 U311 ( .A1(n309), .A2(n308), .A3(n310), .ZN(n8) );
  INV_X1 U312 ( .A(a[1]), .ZN(n323) );
  NOR2_X1 U313 ( .A1(n324), .A2(n312), .ZN(product[0]) );
  OAI22_X1 U314 ( .A1(n325), .A2(n326), .B1(n327), .B2(n324), .ZN(n99) );
  OAI22_X1 U315 ( .A1(n327), .A2(n326), .B1(n328), .B2(n324), .ZN(n98) );
  XNOR2_X1 U316 ( .A(b[6]), .B(a[1]), .ZN(n327) );
  OAI22_X1 U317 ( .A1(n324), .A2(n328), .B1(n326), .B2(n328), .ZN(n329) );
  XNOR2_X1 U318 ( .A(b[7]), .B(a[1]), .ZN(n328) );
  NOR2_X1 U319 ( .A1(n293), .A2(n312), .ZN(n96) );
  OAI22_X1 U320 ( .A1(n331), .A2(n332), .B1(n294), .B2(n333), .ZN(n95) );
  XNOR2_X1 U321 ( .A(a[3]), .B(n311), .ZN(n331) );
  OAI22_X1 U322 ( .A1(n333), .A2(n332), .B1(n294), .B2(n334), .ZN(n94) );
  XNOR2_X1 U323 ( .A(n208), .B(a[3]), .ZN(n333) );
  OAI22_X1 U324 ( .A1(n334), .A2(n332), .B1(n294), .B2(n335), .ZN(n93) );
  XNOR2_X1 U325 ( .A(b[2]), .B(a[3]), .ZN(n334) );
  OAI22_X1 U326 ( .A1(n335), .A2(n332), .B1(n293), .B2(n336), .ZN(n92) );
  XNOR2_X1 U327 ( .A(b[3]), .B(a[3]), .ZN(n335) );
  OAI22_X1 U328 ( .A1(n336), .A2(n332), .B1(n294), .B2(n337), .ZN(n91) );
  XNOR2_X1 U329 ( .A(b[4]), .B(a[3]), .ZN(n336) );
  OAI22_X1 U330 ( .A1(n339), .A2(n293), .B1(n332), .B2(n339), .ZN(n338) );
  NOR2_X1 U331 ( .A1(n249), .A2(n312), .ZN(n88) );
  XNOR2_X1 U332 ( .A(a[5]), .B(n284), .ZN(n341) );
  OAI22_X1 U333 ( .A1(n343), .A2(n342), .B1(n249), .B2(n344), .ZN(n86) );
  XNOR2_X1 U334 ( .A(n217), .B(a[5]), .ZN(n343) );
  OAI22_X1 U335 ( .A1(n344), .A2(n342), .B1(n249), .B2(n345), .ZN(n85) );
  XNOR2_X1 U336 ( .A(b[2]), .B(a[5]), .ZN(n344) );
  OAI22_X1 U337 ( .A1(n345), .A2(n342), .B1(n249), .B2(n346), .ZN(n84) );
  XNOR2_X1 U338 ( .A(n209), .B(a[5]), .ZN(n345) );
  OAI22_X1 U339 ( .A1(n346), .A2(n342), .B1(n249), .B2(n347), .ZN(n83) );
  XNOR2_X1 U340 ( .A(b[4]), .B(a[5]), .ZN(n346) );
  OAI22_X1 U341 ( .A1(n347), .A2(n342), .B1(n249), .B2(n348), .ZN(n82) );
  XNOR2_X1 U342 ( .A(b[5]), .B(a[5]), .ZN(n347) );
  OAI22_X1 U343 ( .A1(n350), .A2(n249), .B1(n342), .B2(n350), .ZN(n349) );
  NOR2_X1 U344 ( .A1(n351), .A2(n312), .ZN(n80) );
  OAI22_X1 U345 ( .A1(n352), .A2(n353), .B1(n351), .B2(n354), .ZN(n79) );
  XNOR2_X1 U346 ( .A(a[7]), .B(n284), .ZN(n352) );
  OAI22_X1 U347 ( .A1(n355), .A2(n353), .B1(n351), .B2(n356), .ZN(n77) );
  OAI22_X1 U348 ( .A1(n356), .A2(n353), .B1(n351), .B2(n357), .ZN(n76) );
  XNOR2_X1 U349 ( .A(n209), .B(a[7]), .ZN(n356) );
  OAI22_X1 U350 ( .A1(n357), .A2(n353), .B1(n351), .B2(n358), .ZN(n75) );
  XNOR2_X1 U351 ( .A(b[4]), .B(a[7]), .ZN(n357) );
  OAI22_X1 U352 ( .A1(n358), .A2(n353), .B1(n351), .B2(n359), .ZN(n74) );
  XNOR2_X1 U353 ( .A(b[5]), .B(a[7]), .ZN(n358) );
  OAI22_X1 U354 ( .A1(n361), .A2(n351), .B1(n353), .B2(n361), .ZN(n360) );
  OAI21_X1 U355 ( .B1(n311), .B2(n323), .A(n326), .ZN(n72) );
  OAI21_X1 U356 ( .B1(n321), .B2(n332), .A(n362), .ZN(n71) );
  OR3_X1 U357 ( .A1(n293), .A2(n284), .A3(n321), .ZN(n362) );
  OAI21_X1 U358 ( .B1(n318), .B2(n342), .A(n363), .ZN(n70) );
  OAI21_X1 U359 ( .B1(n315), .B2(n353), .A(n364), .ZN(n69) );
  OR3_X1 U360 ( .A1(n351), .A2(n284), .A3(n315), .ZN(n364) );
  XNOR2_X1 U361 ( .A(n365), .B(n366), .ZN(n38) );
  OR2_X1 U362 ( .A1(n365), .A2(n366), .ZN(n37) );
  OAI22_X1 U363 ( .A1(n337), .A2(n332), .B1(n293), .B2(n367), .ZN(n366) );
  XNOR2_X1 U364 ( .A(b[5]), .B(a[3]), .ZN(n337) );
  OAI22_X1 U365 ( .A1(n354), .A2(n353), .B1(n351), .B2(n355), .ZN(n365) );
  XNOR2_X1 U366 ( .A(b[2]), .B(a[7]), .ZN(n355) );
  XNOR2_X1 U367 ( .A(n217), .B(a[7]), .ZN(n354) );
  OAI22_X1 U368 ( .A1(n367), .A2(n332), .B1(n294), .B2(n339), .ZN(n31) );
  XNOR2_X1 U369 ( .A(b[7]), .B(a[3]), .ZN(n339) );
  XNOR2_X1 U370 ( .A(b[6]), .B(a[3]), .ZN(n367) );
  OAI22_X1 U371 ( .A1(n348), .A2(n342), .B1(n249), .B2(n350), .ZN(n21) );
  XNOR2_X1 U372 ( .A(b[7]), .B(a[5]), .ZN(n350) );
  XNOR2_X1 U373 ( .A(n318), .B(a[4]), .ZN(n369) );
  XNOR2_X1 U374 ( .A(b[6]), .B(a[5]), .ZN(n348) );
  OAI22_X1 U375 ( .A1(n359), .A2(n353), .B1(n351), .B2(n361), .ZN(n15) );
  XNOR2_X1 U376 ( .A(b[7]), .B(a[7]), .ZN(n361) );
  XNOR2_X1 U377 ( .A(n315), .B(a[6]), .ZN(n370) );
  XNOR2_X1 U378 ( .A(b[6]), .B(a[7]), .ZN(n359) );
  OAI22_X1 U379 ( .A1(n284), .A2(n326), .B1(n371), .B2(n324), .ZN(n104) );
  OAI22_X1 U380 ( .A1(n371), .A2(n326), .B1(n372), .B2(n324), .ZN(n103) );
  OAI22_X1 U381 ( .A1(n372), .A2(n326), .B1(n373), .B2(n324), .ZN(n102) );
  XNOR2_X1 U382 ( .A(b[2]), .B(a[1]), .ZN(n372) );
  OAI22_X1 U383 ( .A1(n326), .A2(n373), .B1(n374), .B2(n324), .ZN(n101) );
  XNOR2_X1 U384 ( .A(b[3]), .B(a[1]), .ZN(n373) );
  OAI22_X1 U385 ( .A1(n374), .A2(n326), .B1(n325), .B2(n324), .ZN(n100) );
  XNOR2_X1 U386 ( .A(b[5]), .B(a[1]), .ZN(n325) );
  NAND2_X1 U387 ( .A1(a[1]), .A2(n324), .ZN(n326) );
  XNOR2_X1 U388 ( .A(b[4]), .B(a[1]), .ZN(n374) );
endmodule


module mac_26 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_26_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_26_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_25_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  wire   [15:1] carry;

  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n64) );
  CLKBUF_X1 U2 ( .A(carry[3]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(carry[10]), .Z(n2) );
  NAND3_X1 U4 ( .A1(n7), .A2(n8), .A3(n9), .ZN(n3) );
  NAND3_X1 U5 ( .A1(n7), .A2(n8), .A3(n9), .ZN(n4) );
  XNOR2_X1 U6 ( .A(B[15]), .B(A[15]), .ZN(n5) );
  XOR2_X1 U7 ( .A(B[10]), .B(A[10]), .Z(n6) );
  XOR2_X1 U8 ( .A(n2), .B(n6), .Z(SUM[10]) );
  NAND2_X1 U9 ( .A1(carry[10]), .A2(B[10]), .ZN(n7) );
  NAND2_X1 U10 ( .A1(carry[10]), .A2(A[10]), .ZN(n8) );
  NAND2_X1 U11 ( .A1(B[10]), .A2(A[10]), .ZN(n9) );
  NAND3_X1 U12 ( .A1(n7), .A2(n8), .A3(n9), .ZN(carry[11]) );
  NAND3_X1 U13 ( .A1(n16), .A2(n17), .A3(n18), .ZN(n10) );
  XOR2_X1 U14 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR2_X1 U15 ( .A(carry[2]), .B(n11), .Z(SUM[2]) );
  NAND2_X1 U16 ( .A1(carry[2]), .A2(B[2]), .ZN(n12) );
  NAND2_X1 U17 ( .A1(carry[2]), .A2(A[2]), .ZN(n13) );
  NAND2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n14) );
  NAND3_X1 U19 ( .A1(n12), .A2(n13), .A3(n14), .ZN(carry[3]) );
  XOR2_X1 U20 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR2_X1 U21 ( .A(n1), .B(n15), .Z(SUM[3]) );
  NAND2_X1 U22 ( .A1(carry[3]), .A2(B[3]), .ZN(n16) );
  NAND2_X1 U23 ( .A1(carry[3]), .A2(A[3]), .ZN(n17) );
  NAND2_X1 U24 ( .A1(B[3]), .A2(A[3]), .ZN(n18) );
  NAND3_X1 U25 ( .A1(n16), .A2(n17), .A3(n18), .ZN(carry[4]) );
  NAND3_X1 U26 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n19) );
  NAND3_X1 U27 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n20) );
  NAND3_X1 U28 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n21) );
  NAND3_X1 U29 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n22) );
  NAND3_X1 U30 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n23) );
  NAND3_X1 U31 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n24) );
  XOR2_X1 U32 ( .A(B[1]), .B(A[1]), .Z(n25) );
  XOR2_X1 U33 ( .A(n64), .B(n25), .Z(SUM[1]) );
  NAND2_X1 U34 ( .A1(n64), .A2(B[1]), .ZN(n26) );
  NAND2_X1 U35 ( .A1(n64), .A2(A[1]), .ZN(n27) );
  NAND2_X1 U36 ( .A1(B[1]), .A2(A[1]), .ZN(n28) );
  NAND3_X1 U37 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[2]) );
  XOR2_X1 U38 ( .A(B[11]), .B(A[11]), .Z(n29) );
  XOR2_X1 U39 ( .A(carry[11]), .B(n29), .Z(SUM[11]) );
  NAND2_X1 U40 ( .A1(n4), .A2(B[11]), .ZN(n30) );
  NAND2_X1 U41 ( .A1(n3), .A2(A[11]), .ZN(n31) );
  NAND2_X1 U42 ( .A1(B[11]), .A2(A[11]), .ZN(n32) );
  NAND3_X1 U43 ( .A1(n30), .A2(n31), .A3(n32), .ZN(carry[12]) );
  XOR2_X1 U44 ( .A(B[4]), .B(A[4]), .Z(n33) );
  XOR2_X1 U45 ( .A(n10), .B(n33), .Z(SUM[4]) );
  NAND2_X1 U46 ( .A1(n10), .A2(B[4]), .ZN(n34) );
  NAND2_X1 U47 ( .A1(carry[4]), .A2(A[4]), .ZN(n35) );
  NAND2_X1 U48 ( .A1(B[4]), .A2(A[4]), .ZN(n36) );
  NAND3_X1 U49 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[5]) );
  XNOR2_X1 U50 ( .A(carry[15]), .B(n5), .ZN(SUM[15]) );
  XOR2_X1 U51 ( .A(B[12]), .B(A[12]), .Z(n37) );
  XOR2_X1 U52 ( .A(n20), .B(n37), .Z(SUM[12]) );
  NAND2_X1 U53 ( .A1(n19), .A2(B[12]), .ZN(n38) );
  NAND2_X1 U54 ( .A1(carry[12]), .A2(A[12]), .ZN(n39) );
  NAND2_X1 U55 ( .A1(B[12]), .A2(A[12]), .ZN(n40) );
  NAND3_X1 U56 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[13]) );
  XOR2_X1 U57 ( .A(B[5]), .B(A[5]), .Z(n41) );
  XOR2_X1 U58 ( .A(n22), .B(n41), .Z(SUM[5]) );
  NAND2_X1 U59 ( .A1(n22), .A2(B[5]), .ZN(n42) );
  NAND2_X1 U60 ( .A1(carry[5]), .A2(A[5]), .ZN(n43) );
  NAND2_X1 U61 ( .A1(B[5]), .A2(A[5]), .ZN(n44) );
  NAND3_X1 U62 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[6]) );
  NAND3_X1 U63 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n45) );
  NAND3_X1 U64 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n46) );
  NAND3_X1 U65 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n47) );
  XOR2_X1 U66 ( .A(B[13]), .B(A[13]), .Z(n48) );
  XOR2_X1 U67 ( .A(n21), .B(n48), .Z(SUM[13]) );
  NAND2_X1 U68 ( .A1(n21), .A2(B[13]), .ZN(n49) );
  NAND2_X1 U69 ( .A1(carry[13]), .A2(A[13]), .ZN(n50) );
  NAND2_X1 U70 ( .A1(B[13]), .A2(A[13]), .ZN(n51) );
  NAND3_X1 U71 ( .A1(n49), .A2(n50), .A3(n51), .ZN(carry[14]) );
  XOR2_X1 U72 ( .A(B[6]), .B(A[6]), .Z(n52) );
  XOR2_X1 U73 ( .A(n24), .B(n52), .Z(SUM[6]) );
  NAND2_X1 U74 ( .A1(n23), .A2(B[6]), .ZN(n53) );
  NAND2_X1 U75 ( .A1(carry[6]), .A2(A[6]), .ZN(n54) );
  NAND2_X1 U76 ( .A1(B[6]), .A2(A[6]), .ZN(n55) );
  NAND3_X1 U77 ( .A1(n53), .A2(n54), .A3(n55), .ZN(carry[7]) );
  XOR2_X1 U78 ( .A(B[14]), .B(A[14]), .Z(n56) );
  XOR2_X1 U79 ( .A(n46), .B(n56), .Z(SUM[14]) );
  NAND2_X1 U80 ( .A1(n45), .A2(B[14]), .ZN(n57) );
  NAND2_X1 U81 ( .A1(carry[14]), .A2(A[14]), .ZN(n58) );
  NAND2_X1 U82 ( .A1(B[14]), .A2(A[14]), .ZN(n59) );
  NAND3_X1 U83 ( .A1(n57), .A2(n58), .A3(n59), .ZN(carry[15]) );
  XOR2_X1 U84 ( .A(B[7]), .B(A[7]), .Z(n60) );
  XOR2_X1 U85 ( .A(carry[7]), .B(n60), .Z(SUM[7]) );
  NAND2_X1 U86 ( .A1(n47), .A2(B[7]), .ZN(n61) );
  NAND2_X1 U87 ( .A1(n47), .A2(A[7]), .ZN(n62) );
  NAND2_X1 U88 ( .A1(B[7]), .A2(A[7]), .ZN(n63) );
  NAND3_X1 U89 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[8]) );
  XOR2_X1 U90 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_25_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n316), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n315), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n319), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n318), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n321), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  AND2_X1 U157 ( .A1(n210), .A2(n102), .ZN(n206) );
  CLKBUF_X1 U158 ( .A(n339), .Z(n207) );
  NAND2_X1 U159 ( .A1(n251), .A2(n40), .ZN(n208) );
  NAND2_X1 U160 ( .A1(n225), .A2(n28), .ZN(n209) );
  OAI22_X1 U161 ( .A1(n330), .A2(n331), .B1(n292), .B2(n332), .ZN(n210) );
  CLKBUF_X1 U162 ( .A(n56), .Z(n211) );
  CLKBUF_X1 U163 ( .A(n301), .Z(n212) );
  CLKBUF_X1 U164 ( .A(n264), .Z(n213) );
  NAND3_X1 U165 ( .A1(n300), .A2(n301), .A3(n302), .ZN(n214) );
  XNOR2_X1 U166 ( .A(a[4]), .B(a[3]), .ZN(n339) );
  CLKBUF_X1 U167 ( .A(n305), .Z(n215) );
  CLKBUF_X1 U168 ( .A(n209), .Z(n216) );
  CLKBUF_X1 U169 ( .A(b[1]), .Z(n217) );
  CLKBUF_X1 U170 ( .A(n262), .Z(n218) );
  CLKBUF_X1 U171 ( .A(b[1]), .Z(n219) );
  CLKBUF_X1 U172 ( .A(n225), .Z(n220) );
  AND2_X1 U173 ( .A1(n104), .A2(n72), .ZN(n221) );
  CLKBUF_X1 U174 ( .A(n208), .Z(n222) );
  NAND3_X1 U175 ( .A1(n208), .A2(n282), .A3(n283), .ZN(n223) );
  NAND3_X1 U176 ( .A1(n222), .A2(n282), .A3(n283), .ZN(n224) );
  NAND3_X1 U177 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n225) );
  XOR2_X1 U178 ( .A(n34), .B(n39), .Z(n226) );
  XOR2_X1 U179 ( .A(n224), .B(n226), .Z(product[8]) );
  NAND2_X1 U180 ( .A1(n223), .A2(n34), .ZN(n227) );
  NAND2_X1 U181 ( .A1(n8), .A2(n39), .ZN(n228) );
  NAND2_X1 U182 ( .A1(n34), .A2(n39), .ZN(n229) );
  NAND3_X1 U183 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n7) );
  NAND3_X1 U184 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n230) );
  XOR2_X1 U185 ( .A(n100), .B(n93), .Z(n231) );
  XOR2_X1 U186 ( .A(n52), .B(n231), .Z(n50) );
  NAND2_X1 U187 ( .A1(n237), .A2(n100), .ZN(n232) );
  NAND2_X1 U188 ( .A1(n237), .A2(n93), .ZN(n233) );
  NAND2_X1 U189 ( .A1(n100), .A2(n93), .ZN(n234) );
  NAND3_X1 U190 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n49) );
  NAND3_X1 U191 ( .A1(n254), .A2(n253), .A3(n255), .ZN(n235) );
  NAND3_X1 U192 ( .A1(n216), .A2(n253), .A3(n255), .ZN(n236) );
  CLKBUF_X1 U193 ( .A(n52), .Z(n237) );
  CLKBUF_X1 U194 ( .A(n273), .Z(n238) );
  NAND3_X1 U195 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n239) );
  NAND3_X1 U196 ( .A1(n218), .A2(n263), .A3(n213), .ZN(n240) );
  NAND2_X2 U197 ( .A1(n350), .A2(n369), .ZN(n352) );
  XOR2_X2 U198 ( .A(a[6]), .B(n317), .Z(n350) );
  CLKBUF_X1 U199 ( .A(n251), .Z(n241) );
  XOR2_X1 U200 ( .A(n103), .B(n96), .Z(n242) );
  XOR2_X1 U201 ( .A(n221), .B(n242), .Z(product[2]) );
  NAND2_X1 U202 ( .A1(n221), .A2(n103), .ZN(n243) );
  NAND2_X1 U203 ( .A1(n14), .A2(n96), .ZN(n244) );
  NAND2_X1 U204 ( .A1(n103), .A2(n96), .ZN(n245) );
  NAND3_X1 U205 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n13) );
  CLKBUF_X1 U206 ( .A(n219), .Z(n246) );
  CLKBUF_X1 U207 ( .A(n309), .Z(n247) );
  CLKBUF_X1 U208 ( .A(n274), .Z(n248) );
  NAND3_X1 U209 ( .A1(n308), .A2(n309), .A3(n310), .ZN(n249) );
  NAND3_X1 U210 ( .A1(n308), .A2(n247), .A3(n310), .ZN(n250) );
  NAND3_X1 U211 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n251) );
  XOR2_X1 U212 ( .A(n33), .B(n28), .Z(n252) );
  XOR2_X1 U213 ( .A(n220), .B(n252), .Z(product[9]) );
  NAND2_X1 U214 ( .A1(n7), .A2(n33), .ZN(n253) );
  NAND2_X1 U215 ( .A1(n225), .A2(n28), .ZN(n254) );
  NAND2_X1 U216 ( .A1(n33), .A2(n28), .ZN(n255) );
  NAND3_X1 U217 ( .A1(n209), .A2(n253), .A3(n255), .ZN(n6) );
  NAND3_X1 U218 ( .A1(n289), .A2(n288), .A3(n290), .ZN(n256) );
  XOR2_X1 U219 ( .A(n46), .B(n49), .Z(n257) );
  XOR2_X1 U220 ( .A(n250), .B(n257), .Z(product[6]) );
  NAND2_X1 U221 ( .A1(n249), .A2(n46), .ZN(n258) );
  NAND2_X1 U222 ( .A1(n10), .A2(n49), .ZN(n259) );
  NAND2_X1 U223 ( .A1(n46), .A2(n49), .ZN(n260) );
  NAND3_X1 U224 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n9) );
  XOR2_X1 U225 ( .A(n211), .B(n71), .Z(n261) );
  XOR2_X1 U226 ( .A(n230), .B(n261), .Z(product[3]) );
  NAND2_X1 U227 ( .A1(n230), .A2(n56), .ZN(n262) );
  NAND2_X1 U228 ( .A1(n13), .A2(n71), .ZN(n263) );
  NAND2_X1 U229 ( .A1(n56), .A2(n71), .ZN(n264) );
  NAND3_X1 U230 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n12) );
  NAND3_X1 U231 ( .A1(n300), .A2(n301), .A3(n302), .ZN(n265) );
  NAND3_X1 U232 ( .A1(n212), .A2(n300), .A3(n302), .ZN(n266) );
  NAND3_X1 U233 ( .A1(n274), .A2(n273), .A3(n275), .ZN(n267) );
  NAND3_X1 U234 ( .A1(n238), .A2(n248), .A3(n275), .ZN(n268) );
  NAND3_X1 U235 ( .A1(n278), .A2(n277), .A3(n279), .ZN(n269) );
  INV_X1 U236 ( .A(n311), .ZN(n270) );
  INV_X1 U237 ( .A(n311), .ZN(n271) );
  XOR2_X1 U238 ( .A(n20), .B(n23), .Z(n272) );
  XOR2_X1 U239 ( .A(n5), .B(n272), .Z(product[11]) );
  NAND2_X1 U240 ( .A1(n256), .A2(n20), .ZN(n273) );
  NAND2_X1 U241 ( .A1(n256), .A2(n23), .ZN(n274) );
  NAND2_X1 U242 ( .A1(n20), .A2(n23), .ZN(n275) );
  NAND3_X1 U243 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n4) );
  XOR2_X1 U244 ( .A(n312), .B(n17), .Z(n276) );
  XOR2_X1 U245 ( .A(n266), .B(n276), .Z(product[13]) );
  NAND2_X1 U246 ( .A1(n214), .A2(n312), .ZN(n277) );
  NAND2_X1 U247 ( .A1(n265), .A2(n17), .ZN(n278) );
  NAND2_X1 U248 ( .A1(n312), .A2(n17), .ZN(n279) );
  NAND3_X1 U249 ( .A1(n277), .A2(n278), .A3(n279), .ZN(n2) );
  XOR2_X1 U250 ( .A(n40), .B(n45), .Z(n280) );
  XOR2_X1 U251 ( .A(n241), .B(n280), .Z(product[7]) );
  NAND2_X1 U252 ( .A1(n251), .A2(n40), .ZN(n281) );
  NAND2_X1 U253 ( .A1(n9), .A2(n45), .ZN(n282) );
  NAND2_X1 U254 ( .A1(n40), .A2(n45), .ZN(n283) );
  NAND3_X1 U255 ( .A1(n281), .A2(n282), .A3(n283), .ZN(n8) );
  NAND3_X1 U256 ( .A1(n306), .A2(n305), .A3(n304), .ZN(n284) );
  NAND3_X1 U257 ( .A1(n304), .A2(n215), .A3(n306), .ZN(n285) );
  XNOR2_X1 U258 ( .A(n219), .B(n291), .ZN(n286) );
  XOR2_X1 U259 ( .A(n27), .B(n24), .Z(n287) );
  XOR2_X1 U260 ( .A(n236), .B(n287), .Z(product[10]) );
  NAND2_X1 U261 ( .A1(n235), .A2(n27), .ZN(n288) );
  NAND2_X1 U262 ( .A1(n6), .A2(n24), .ZN(n289) );
  NAND2_X1 U263 ( .A1(n27), .A2(n24), .ZN(n290) );
  NAND3_X1 U264 ( .A1(n288), .A2(n289), .A3(n290), .ZN(n5) );
  XOR2_X1 U265 ( .A(n95), .B(n102), .Z(n56) );
  BUF_X2 U266 ( .A(a[1]), .Z(n291) );
  NAND2_X2 U267 ( .A1(n339), .A2(n368), .ZN(n341) );
  NAND2_X2 U268 ( .A1(n329), .A2(n367), .ZN(n331) );
  XOR2_X1 U269 ( .A(a[2]), .B(n322), .Z(n292) );
  XOR2_X1 U270 ( .A(a[2]), .B(n322), .Z(n293) );
  INV_X1 U271 ( .A(n15), .ZN(n312) );
  XNOR2_X1 U272 ( .A(n268), .B(n294), .ZN(product[12]) );
  XNOR2_X1 U273 ( .A(n19), .B(n18), .ZN(n294) );
  XNOR2_X1 U274 ( .A(n2), .B(n295), .ZN(product[14]) );
  XNOR2_X1 U275 ( .A(n313), .B(n15), .ZN(n295) );
  AND3_X1 U276 ( .A1(n298), .A2(n297), .A3(n299), .ZN(product[15]) );
  INV_X1 U277 ( .A(n348), .ZN(n316) );
  INV_X1 U278 ( .A(n21), .ZN(n315) );
  INV_X1 U279 ( .A(n328), .ZN(n321) );
  INV_X1 U280 ( .A(n337), .ZN(n319) );
  INV_X1 U281 ( .A(n31), .ZN(n318) );
  INV_X1 U282 ( .A(b[0]), .ZN(n311) );
  XOR2_X1 U283 ( .A(a[2]), .B(n322), .Z(n329) );
  INV_X1 U284 ( .A(a[0]), .ZN(n323) );
  INV_X1 U285 ( .A(a[5]), .ZN(n317) );
  INV_X1 U286 ( .A(a[7]), .ZN(n314) );
  NAND2_X1 U287 ( .A1(n269), .A2(n313), .ZN(n297) );
  NAND2_X1 U288 ( .A1(n2), .A2(n15), .ZN(n298) );
  NAND2_X1 U289 ( .A1(n313), .A2(n15), .ZN(n299) );
  NAND2_X1 U290 ( .A1(n4), .A2(n19), .ZN(n300) );
  NAND2_X1 U291 ( .A1(n267), .A2(n18), .ZN(n301) );
  NAND2_X1 U292 ( .A1(n19), .A2(n18), .ZN(n302) );
  INV_X1 U293 ( .A(n359), .ZN(n313) );
  INV_X1 U294 ( .A(a[3]), .ZN(n320) );
  XOR2_X1 U295 ( .A(n54), .B(n206), .Z(n303) );
  XOR2_X1 U296 ( .A(n303), .B(n240), .Z(product[4]) );
  NAND2_X1 U297 ( .A1(n54), .A2(n206), .ZN(n304) );
  NAND2_X1 U298 ( .A1(n54), .A2(n12), .ZN(n305) );
  NAND2_X1 U299 ( .A1(n206), .A2(n239), .ZN(n306) );
  NAND3_X1 U300 ( .A1(n306), .A2(n305), .A3(n304), .ZN(n11) );
  XOR2_X1 U301 ( .A(n50), .B(n53), .Z(n307) );
  XOR2_X1 U302 ( .A(n307), .B(n285), .Z(product[5]) );
  NAND2_X1 U303 ( .A1(n50), .A2(n53), .ZN(n308) );
  NAND2_X1 U304 ( .A1(n284), .A2(n50), .ZN(n309) );
  NAND2_X1 U305 ( .A1(n11), .A2(n53), .ZN(n310) );
  NAND3_X1 U306 ( .A1(n310), .A2(n309), .A3(n308), .ZN(n10) );
  INV_X1 U307 ( .A(a[1]), .ZN(n322) );
  NOR2_X1 U308 ( .A1(n323), .A2(n311), .ZN(product[0]) );
  OAI22_X1 U309 ( .A1(n324), .A2(n325), .B1(n326), .B2(n323), .ZN(n99) );
  OAI22_X1 U310 ( .A1(n326), .A2(n325), .B1(n327), .B2(n323), .ZN(n98) );
  XNOR2_X1 U311 ( .A(b[6]), .B(n291), .ZN(n326) );
  OAI22_X1 U312 ( .A1(n323), .A2(n327), .B1(n325), .B2(n327), .ZN(n328) );
  XNOR2_X1 U313 ( .A(b[7]), .B(n291), .ZN(n327) );
  NOR2_X1 U314 ( .A1(n293), .A2(n311), .ZN(n96) );
  OAI22_X1 U315 ( .A1(n330), .A2(n331), .B1(n292), .B2(n332), .ZN(n95) );
  XNOR2_X1 U316 ( .A(a[3]), .B(b[0]), .ZN(n330) );
  OAI22_X1 U317 ( .A1(n332), .A2(n331), .B1(n292), .B2(n333), .ZN(n94) );
  XNOR2_X1 U318 ( .A(n217), .B(a[3]), .ZN(n332) );
  OAI22_X1 U319 ( .A1(n333), .A2(n331), .B1(n292), .B2(n334), .ZN(n93) );
  XNOR2_X1 U320 ( .A(b[2]), .B(a[3]), .ZN(n333) );
  OAI22_X1 U321 ( .A1(n334), .A2(n331), .B1(n293), .B2(n335), .ZN(n92) );
  XNOR2_X1 U322 ( .A(b[3]), .B(a[3]), .ZN(n334) );
  OAI22_X1 U323 ( .A1(n335), .A2(n331), .B1(n293), .B2(n336), .ZN(n91) );
  XNOR2_X1 U324 ( .A(b[4]), .B(a[3]), .ZN(n335) );
  OAI22_X1 U325 ( .A1(n338), .A2(n292), .B1(n331), .B2(n338), .ZN(n337) );
  NOR2_X1 U326 ( .A1(n339), .A2(n311), .ZN(n88) );
  OAI22_X1 U327 ( .A1(n340), .A2(n341), .B1(n339), .B2(n342), .ZN(n87) );
  XNOR2_X1 U328 ( .A(a[5]), .B(n270), .ZN(n340) );
  OAI22_X1 U329 ( .A1(n342), .A2(n341), .B1(n339), .B2(n343), .ZN(n86) );
  XNOR2_X1 U330 ( .A(n246), .B(a[5]), .ZN(n342) );
  OAI22_X1 U331 ( .A1(n343), .A2(n341), .B1(n339), .B2(n344), .ZN(n85) );
  XNOR2_X1 U332 ( .A(b[2]), .B(a[5]), .ZN(n343) );
  OAI22_X1 U333 ( .A1(n344), .A2(n341), .B1(n339), .B2(n345), .ZN(n84) );
  XNOR2_X1 U334 ( .A(b[3]), .B(a[5]), .ZN(n344) );
  OAI22_X1 U335 ( .A1(n345), .A2(n341), .B1(n339), .B2(n346), .ZN(n83) );
  XNOR2_X1 U336 ( .A(b[4]), .B(a[5]), .ZN(n345) );
  OAI22_X1 U337 ( .A1(n346), .A2(n341), .B1(n339), .B2(n347), .ZN(n82) );
  XNOR2_X1 U338 ( .A(b[5]), .B(a[5]), .ZN(n346) );
  OAI22_X1 U339 ( .A1(n349), .A2(n207), .B1(n341), .B2(n349), .ZN(n348) );
  NOR2_X1 U340 ( .A1(n350), .A2(n311), .ZN(n80) );
  OAI22_X1 U341 ( .A1(n351), .A2(n352), .B1(n350), .B2(n353), .ZN(n79) );
  XNOR2_X1 U342 ( .A(a[7]), .B(n270), .ZN(n351) );
  OAI22_X1 U343 ( .A1(n354), .A2(n352), .B1(n350), .B2(n355), .ZN(n77) );
  OAI22_X1 U344 ( .A1(n355), .A2(n352), .B1(n350), .B2(n356), .ZN(n76) );
  XNOR2_X1 U345 ( .A(b[3]), .B(a[7]), .ZN(n355) );
  OAI22_X1 U346 ( .A1(n356), .A2(n352), .B1(n350), .B2(n357), .ZN(n75) );
  XNOR2_X1 U347 ( .A(b[4]), .B(a[7]), .ZN(n356) );
  OAI22_X1 U348 ( .A1(n357), .A2(n352), .B1(n350), .B2(n358), .ZN(n74) );
  XNOR2_X1 U349 ( .A(b[5]), .B(a[7]), .ZN(n357) );
  OAI22_X1 U350 ( .A1(n360), .A2(n350), .B1(n352), .B2(n360), .ZN(n359) );
  OAI21_X1 U351 ( .B1(n270), .B2(n322), .A(n325), .ZN(n72) );
  OAI21_X1 U352 ( .B1(n320), .B2(n331), .A(n361), .ZN(n71) );
  OR3_X1 U353 ( .A1(n293), .A2(n271), .A3(n320), .ZN(n361) );
  OAI21_X1 U354 ( .B1(n317), .B2(n341), .A(n362), .ZN(n70) );
  OR3_X1 U355 ( .A1(n339), .A2(n271), .A3(n317), .ZN(n362) );
  OAI21_X1 U356 ( .B1(n314), .B2(n352), .A(n363), .ZN(n69) );
  OR3_X1 U357 ( .A1(n350), .A2(n271), .A3(n314), .ZN(n363) );
  XNOR2_X1 U358 ( .A(n364), .B(n365), .ZN(n38) );
  OR2_X1 U359 ( .A1(n364), .A2(n365), .ZN(n37) );
  OAI22_X1 U360 ( .A1(n336), .A2(n331), .B1(n292), .B2(n366), .ZN(n365) );
  XNOR2_X1 U361 ( .A(b[5]), .B(a[3]), .ZN(n336) );
  OAI22_X1 U362 ( .A1(n353), .A2(n352), .B1(n350), .B2(n354), .ZN(n364) );
  XNOR2_X1 U363 ( .A(b[2]), .B(a[7]), .ZN(n354) );
  XNOR2_X1 U364 ( .A(n246), .B(a[7]), .ZN(n353) );
  OAI22_X1 U365 ( .A1(n366), .A2(n331), .B1(n293), .B2(n338), .ZN(n31) );
  XNOR2_X1 U366 ( .A(b[7]), .B(a[3]), .ZN(n338) );
  XNOR2_X1 U367 ( .A(n320), .B(a[2]), .ZN(n367) );
  XNOR2_X1 U368 ( .A(b[6]), .B(a[3]), .ZN(n366) );
  OAI22_X1 U369 ( .A1(n347), .A2(n341), .B1(n207), .B2(n349), .ZN(n21) );
  XNOR2_X1 U370 ( .A(b[7]), .B(a[5]), .ZN(n349) );
  XNOR2_X1 U371 ( .A(n317), .B(a[4]), .ZN(n368) );
  XNOR2_X1 U372 ( .A(b[6]), .B(a[5]), .ZN(n347) );
  OAI22_X1 U373 ( .A1(n358), .A2(n352), .B1(n350), .B2(n360), .ZN(n15) );
  XNOR2_X1 U374 ( .A(b[7]), .B(a[7]), .ZN(n360) );
  XNOR2_X1 U375 ( .A(n314), .B(a[6]), .ZN(n369) );
  XNOR2_X1 U376 ( .A(b[6]), .B(a[7]), .ZN(n358) );
  OAI22_X1 U377 ( .A1(n271), .A2(n325), .B1(n370), .B2(n323), .ZN(n104) );
  OAI22_X1 U378 ( .A1(n286), .A2(n325), .B1(n371), .B2(n323), .ZN(n103) );
  XNOR2_X1 U379 ( .A(b[1]), .B(n291), .ZN(n370) );
  OAI22_X1 U380 ( .A1(n371), .A2(n325), .B1(n372), .B2(n323), .ZN(n102) );
  XNOR2_X1 U381 ( .A(b[2]), .B(n291), .ZN(n371) );
  OAI22_X1 U382 ( .A1(n372), .A2(n325), .B1(n373), .B2(n323), .ZN(n101) );
  XNOR2_X1 U383 ( .A(b[3]), .B(n291), .ZN(n372) );
  OAI22_X1 U384 ( .A1(n373), .A2(n325), .B1(n324), .B2(n323), .ZN(n100) );
  XNOR2_X1 U385 ( .A(b[5]), .B(n291), .ZN(n324) );
  NAND2_X1 U386 ( .A1(n291), .A2(n323), .ZN(n325) );
  XNOR2_X1 U387 ( .A(b[4]), .B(n291), .ZN(n373) );
endmodule


module mac_25 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_25_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_25_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X2 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_24_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;
  wire   [15:1] carry;

  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n76) );
  XOR2_X1 U2 ( .A(B[15]), .B(A[15]), .Z(n1) );
  XOR2_X1 U3 ( .A(carry[15]), .B(n1), .Z(SUM[15]) );
  NAND3_X1 U4 ( .A1(n32), .A2(n33), .A3(n34), .ZN(n2) );
  NAND3_X1 U5 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n3) );
  NAND3_X1 U6 ( .A1(n7), .A2(n8), .A3(n9), .ZN(n4) );
  NAND2_X1 U7 ( .A1(n30), .A2(B[9]), .ZN(n5) );
  XOR2_X1 U8 ( .A(B[3]), .B(A[3]), .Z(n6) );
  XOR2_X1 U9 ( .A(carry[3]), .B(n6), .Z(SUM[3]) );
  NAND2_X1 U10 ( .A1(carry[3]), .A2(B[3]), .ZN(n7) );
  NAND2_X1 U11 ( .A1(carry[3]), .A2(A[3]), .ZN(n8) );
  NAND2_X1 U12 ( .A1(B[3]), .A2(A[3]), .ZN(n9) );
  NAND3_X1 U13 ( .A1(n7), .A2(n8), .A3(n9), .ZN(carry[4]) );
  NAND3_X1 U14 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n10) );
  NAND3_X1 U15 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n11) );
  NAND3_X1 U16 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n12) );
  NAND3_X1 U17 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n13) );
  NAND3_X1 U18 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n14) );
  NAND3_X1 U19 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n15) );
  XOR2_X1 U20 ( .A(B[4]), .B(A[4]), .Z(n16) );
  XOR2_X1 U21 ( .A(n4), .B(n16), .Z(SUM[4]) );
  NAND2_X1 U22 ( .A1(n4), .A2(B[4]), .ZN(n17) );
  NAND2_X1 U23 ( .A1(carry[4]), .A2(A[4]), .ZN(n18) );
  NAND2_X1 U24 ( .A1(B[4]), .A2(A[4]), .ZN(n19) );
  NAND3_X1 U25 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[5]) );
  XOR2_X1 U26 ( .A(B[11]), .B(A[11]), .Z(n20) );
  XOR2_X1 U27 ( .A(n13), .B(n20), .Z(SUM[11]) );
  NAND2_X1 U28 ( .A1(n12), .A2(B[11]), .ZN(n21) );
  NAND2_X1 U29 ( .A1(carry[11]), .A2(A[11]), .ZN(n22) );
  NAND2_X1 U30 ( .A1(B[11]), .A2(A[11]), .ZN(n23) );
  NAND3_X1 U31 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[12]) );
  NAND3_X1 U32 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n24) );
  XOR2_X1 U33 ( .A(B[5]), .B(A[5]), .Z(n25) );
  XOR2_X1 U34 ( .A(n11), .B(n25), .Z(SUM[5]) );
  NAND2_X1 U35 ( .A1(n10), .A2(B[5]), .ZN(n26) );
  NAND2_X1 U36 ( .A1(carry[5]), .A2(A[5]), .ZN(n27) );
  NAND2_X1 U37 ( .A1(B[5]), .A2(A[5]), .ZN(n28) );
  NAND3_X1 U38 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[6]) );
  NAND3_X1 U39 ( .A1(n32), .A2(n33), .A3(n34), .ZN(n29) );
  NAND3_X1 U40 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n30) );
  XOR2_X1 U41 ( .A(B[12]), .B(A[12]), .Z(n31) );
  XOR2_X1 U42 ( .A(n3), .B(n31), .Z(SUM[12]) );
  NAND2_X1 U43 ( .A1(n3), .A2(B[12]), .ZN(n32) );
  NAND2_X1 U44 ( .A1(carry[12]), .A2(A[12]), .ZN(n33) );
  NAND2_X1 U45 ( .A1(B[12]), .A2(A[12]), .ZN(n34) );
  NAND3_X1 U46 ( .A1(n32), .A2(n33), .A3(n34), .ZN(carry[13]) );
  XOR2_X1 U47 ( .A(B[6]), .B(A[6]), .Z(n35) );
  XOR2_X1 U48 ( .A(n14), .B(n35), .Z(SUM[6]) );
  NAND2_X1 U49 ( .A1(n14), .A2(B[6]), .ZN(n36) );
  NAND2_X1 U50 ( .A1(carry[6]), .A2(A[6]), .ZN(n37) );
  NAND2_X1 U51 ( .A1(B[6]), .A2(A[6]), .ZN(n38) );
  NAND3_X1 U52 ( .A1(n36), .A2(n37), .A3(n38), .ZN(carry[7]) );
  NAND3_X1 U53 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n39) );
  NAND3_X1 U54 ( .A1(n5), .A2(n66), .A3(n67), .ZN(n40) );
  NAND3_X1 U55 ( .A1(n5), .A2(n66), .A3(n67), .ZN(n41) );
  XOR2_X1 U56 ( .A(B[10]), .B(A[10]), .Z(n42) );
  XOR2_X1 U57 ( .A(n41), .B(n42), .Z(SUM[10]) );
  NAND2_X1 U58 ( .A1(n40), .A2(B[10]), .ZN(n43) );
  NAND2_X1 U59 ( .A1(carry[10]), .A2(A[10]), .ZN(n44) );
  NAND2_X1 U60 ( .A1(B[10]), .A2(A[10]), .ZN(n45) );
  NAND3_X1 U61 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[11]) );
  XOR2_X1 U62 ( .A(B[13]), .B(A[13]), .Z(n46) );
  XOR2_X1 U63 ( .A(n2), .B(n46), .Z(SUM[13]) );
  NAND2_X1 U64 ( .A1(carry[13]), .A2(B[13]), .ZN(n47) );
  NAND2_X1 U65 ( .A1(n29), .A2(A[13]), .ZN(n48) );
  NAND2_X1 U66 ( .A1(B[13]), .A2(A[13]), .ZN(n49) );
  NAND3_X1 U67 ( .A1(n48), .A2(n47), .A3(n49), .ZN(carry[14]) );
  XOR2_X1 U68 ( .A(B[7]), .B(A[7]), .Z(n50) );
  XOR2_X1 U69 ( .A(n15), .B(n50), .Z(SUM[7]) );
  NAND2_X1 U70 ( .A1(n15), .A2(B[7]), .ZN(n51) );
  NAND2_X1 U71 ( .A1(carry[7]), .A2(A[7]), .ZN(n52) );
  NAND2_X1 U72 ( .A1(B[7]), .A2(A[7]), .ZN(n53) );
  NAND3_X1 U73 ( .A1(n51), .A2(n52), .A3(n53), .ZN(carry[8]) );
  NAND3_X1 U74 ( .A1(n69), .A2(n70), .A3(n71), .ZN(n54) );
  NAND3_X1 U75 ( .A1(n69), .A2(n70), .A3(n71), .ZN(n55) );
  XOR2_X1 U76 ( .A(B[14]), .B(A[14]), .Z(n56) );
  XOR2_X1 U77 ( .A(n39), .B(n56), .Z(SUM[14]) );
  NAND2_X1 U78 ( .A1(n39), .A2(B[14]), .ZN(n57) );
  NAND2_X1 U79 ( .A1(carry[14]), .A2(A[14]), .ZN(n58) );
  NAND2_X1 U80 ( .A1(B[14]), .A2(A[14]), .ZN(n59) );
  NAND3_X1 U81 ( .A1(n57), .A2(n58), .A3(n59), .ZN(carry[15]) );
  XOR2_X1 U82 ( .A(B[8]), .B(A[8]), .Z(n60) );
  XOR2_X1 U83 ( .A(n24), .B(n60), .Z(SUM[8]) );
  NAND2_X1 U84 ( .A1(n24), .A2(B[8]), .ZN(n61) );
  NAND2_X1 U85 ( .A1(carry[8]), .A2(A[8]), .ZN(n62) );
  NAND2_X1 U86 ( .A1(B[8]), .A2(A[8]), .ZN(n63) );
  NAND3_X1 U87 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[9]) );
  XOR2_X1 U88 ( .A(B[9]), .B(A[9]), .Z(n64) );
  XOR2_X1 U89 ( .A(n30), .B(n64), .Z(SUM[9]) );
  NAND2_X1 U90 ( .A1(n30), .A2(B[9]), .ZN(n65) );
  NAND2_X1 U91 ( .A1(carry[9]), .A2(A[9]), .ZN(n66) );
  NAND2_X1 U92 ( .A1(B[9]), .A2(A[9]), .ZN(n67) );
  NAND3_X1 U93 ( .A1(n65), .A2(n66), .A3(n67), .ZN(carry[10]) );
  XOR2_X1 U94 ( .A(B[1]), .B(A[1]), .Z(n68) );
  XOR2_X1 U95 ( .A(n76), .B(n68), .Z(SUM[1]) );
  NAND2_X1 U96 ( .A1(n76), .A2(B[1]), .ZN(n69) );
  NAND2_X1 U97 ( .A1(n76), .A2(A[1]), .ZN(n70) );
  NAND2_X1 U98 ( .A1(B[1]), .A2(A[1]), .ZN(n71) );
  NAND3_X1 U99 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[2]) );
  XOR2_X1 U100 ( .A(B[2]), .B(A[2]), .Z(n72) );
  XOR2_X1 U101 ( .A(n55), .B(n72), .Z(SUM[2]) );
  NAND2_X1 U102 ( .A1(n54), .A2(B[2]), .ZN(n73) );
  NAND2_X1 U103 ( .A1(carry[2]), .A2(A[2]), .ZN(n74) );
  NAND2_X1 U104 ( .A1(B[2]), .A2(A[2]), .ZN(n75) );
  NAND3_X1 U105 ( .A1(n73), .A2(n74), .A3(n75), .ZN(carry[3]) );
  XOR2_X1 U106 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_24_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n311), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n310), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n314), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n313), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n316), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  AND2_X1 U157 ( .A1(n104), .A2(n72), .ZN(n206) );
  AND2_X1 U158 ( .A1(n104), .A2(n72), .ZN(n207) );
  AND2_X1 U159 ( .A1(n95), .A2(n102), .ZN(n208) );
  CLKBUF_X1 U160 ( .A(b[1]), .Z(n209) );
  INV_X1 U161 ( .A(n315), .ZN(n210) );
  CLKBUF_X1 U162 ( .A(n238), .Z(n211) );
  NAND3_X1 U163 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n212) );
  NAND2_X1 U164 ( .A1(n231), .A2(n18), .ZN(n213) );
  NAND2_X1 U165 ( .A1(n4), .A2(n19), .ZN(n214) );
  NAND3_X1 U166 ( .A1(n213), .A2(n214), .A3(n297), .ZN(n215) );
  XOR2_X1 U167 ( .A(n95), .B(n102), .Z(n56) );
  CLKBUF_X1 U168 ( .A(n56), .Z(n216) );
  CLKBUF_X1 U169 ( .A(n260), .Z(n217) );
  XNOR2_X1 U170 ( .A(a[6]), .B(a[5]), .ZN(n345) );
  XNOR2_X1 U171 ( .A(a[6]), .B(a[5]), .ZN(n218) );
  CLKBUF_X1 U172 ( .A(n209), .Z(n219) );
  NAND3_X1 U173 ( .A1(n217), .A2(n261), .A3(n262), .ZN(n220) );
  CLKBUF_X1 U174 ( .A(n5), .Z(n221) );
  NAND3_X1 U175 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n222) );
  CLKBUF_X1 U176 ( .A(n280), .Z(n223) );
  NAND2_X1 U177 ( .A1(a[4]), .A2(a[3]), .ZN(n226) );
  NAND2_X1 U178 ( .A1(n224), .A2(n225), .ZN(n227) );
  NAND2_X2 U179 ( .A1(n226), .A2(n227), .ZN(n334) );
  INV_X1 U180 ( .A(a[4]), .ZN(n224) );
  INV_X1 U181 ( .A(a[3]), .ZN(n225) );
  NAND2_X1 U182 ( .A1(b[1]), .A2(a[1]), .ZN(n229) );
  NAND2_X1 U183 ( .A1(n228), .A2(n317), .ZN(n230) );
  NAND2_X1 U184 ( .A1(n229), .A2(n230), .ZN(n365) );
  INV_X1 U185 ( .A(b[1]), .ZN(n228) );
  NAND3_X1 U186 ( .A1(n280), .A2(n281), .A3(n282), .ZN(n231) );
  NAND3_X1 U187 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n232) );
  NAND3_X1 U188 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n233) );
  NAND3_X1 U189 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n234) );
  XOR2_X1 U190 ( .A(n216), .B(n71), .Z(n235) );
  XOR2_X1 U191 ( .A(n232), .B(n235), .Z(product[3]) );
  NAND2_X1 U192 ( .A1(n56), .A2(n232), .ZN(n236) );
  NAND2_X1 U193 ( .A1(n13), .A2(n71), .ZN(n237) );
  NAND2_X1 U194 ( .A1(n56), .A2(n71), .ZN(n238) );
  NAND3_X1 U195 ( .A1(n236), .A2(n237), .A3(n211), .ZN(n12) );
  NAND3_X1 U196 ( .A1(n276), .A2(n275), .A3(n277), .ZN(n239) );
  CLKBUF_X1 U197 ( .A(n222), .Z(n240) );
  CLKBUF_X1 U198 ( .A(n234), .Z(n241) );
  CLKBUF_X1 U199 ( .A(n7), .Z(n242) );
  NAND3_X1 U200 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n243) );
  XOR2_X1 U201 ( .A(n54), .B(n208), .Z(n244) );
  XOR2_X1 U202 ( .A(n12), .B(n244), .Z(product[4]) );
  NAND2_X1 U203 ( .A1(n212), .A2(n54), .ZN(n245) );
  NAND2_X1 U204 ( .A1(n233), .A2(n208), .ZN(n246) );
  NAND2_X1 U205 ( .A1(n54), .A2(n208), .ZN(n247) );
  NAND3_X1 U206 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n11) );
  XOR2_X1 U207 ( .A(n50), .B(n53), .Z(n248) );
  XOR2_X1 U208 ( .A(n241), .B(n248), .Z(product[5]) );
  NAND2_X1 U209 ( .A1(n234), .A2(n50), .ZN(n249) );
  NAND2_X1 U210 ( .A1(n11), .A2(n53), .ZN(n250) );
  NAND2_X1 U211 ( .A1(n50), .A2(n53), .ZN(n251) );
  NAND3_X1 U212 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n10) );
  NAND3_X1 U213 ( .A1(n272), .A2(n271), .A3(n273), .ZN(n252) );
  NAND3_X1 U214 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n253) );
  XOR2_X1 U215 ( .A(n103), .B(n96), .Z(n254) );
  XOR2_X1 U216 ( .A(n14), .B(n254), .Z(product[2]) );
  NAND2_X1 U217 ( .A1(n207), .A2(n103), .ZN(n255) );
  NAND2_X1 U218 ( .A1(n206), .A2(n96), .ZN(n256) );
  NAND2_X1 U219 ( .A1(n103), .A2(n96), .ZN(n257) );
  NAND3_X1 U220 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n13) );
  CLKBUF_X1 U221 ( .A(n214), .Z(n258) );
  XOR2_X1 U222 ( .A(n46), .B(n49), .Z(n259) );
  XOR2_X1 U223 ( .A(n240), .B(n259), .Z(product[6]) );
  NAND2_X1 U224 ( .A1(n222), .A2(n46), .ZN(n260) );
  NAND2_X1 U225 ( .A1(n10), .A2(n49), .ZN(n261) );
  NAND2_X1 U226 ( .A1(n46), .A2(n49), .ZN(n262) );
  NAND3_X1 U227 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n9) );
  NAND3_X1 U228 ( .A1(n285), .A2(n286), .A3(n287), .ZN(n263) );
  CLKBUF_X1 U229 ( .A(n6), .Z(n264) );
  XOR2_X1 U230 ( .A(n33), .B(n28), .Z(n265) );
  XOR2_X1 U231 ( .A(n242), .B(n265), .Z(product[9]) );
  NAND2_X1 U232 ( .A1(n263), .A2(n33), .ZN(n266) );
  NAND2_X1 U233 ( .A1(n7), .A2(n28), .ZN(n267) );
  NAND2_X1 U234 ( .A1(n33), .A2(n28), .ZN(n268) );
  NAND3_X1 U235 ( .A1(n267), .A2(n266), .A3(n268), .ZN(n6) );
  CLKBUF_X1 U236 ( .A(n239), .Z(n269) );
  XOR2_X1 U237 ( .A(n27), .B(n24), .Z(n270) );
  XOR2_X1 U238 ( .A(n264), .B(n270), .Z(product[10]) );
  NAND2_X1 U239 ( .A1(n243), .A2(n27), .ZN(n271) );
  NAND2_X1 U240 ( .A1(n6), .A2(n24), .ZN(n272) );
  NAND2_X1 U241 ( .A1(n27), .A2(n24), .ZN(n273) );
  NAND3_X1 U242 ( .A1(n272), .A2(n271), .A3(n273), .ZN(n5) );
  XOR2_X1 U243 ( .A(n40), .B(n45), .Z(n274) );
  XOR2_X1 U244 ( .A(n220), .B(n274), .Z(product[7]) );
  NAND2_X1 U245 ( .A1(n9), .A2(n40), .ZN(n275) );
  NAND2_X1 U246 ( .A1(n253), .A2(n45), .ZN(n276) );
  NAND2_X1 U247 ( .A1(n40), .A2(n45), .ZN(n277) );
  NAND3_X1 U248 ( .A1(n275), .A2(n276), .A3(n277), .ZN(n8) );
  NAND3_X1 U249 ( .A1(n223), .A2(n281), .A3(n282), .ZN(n278) );
  XOR2_X1 U250 ( .A(n20), .B(n23), .Z(n279) );
  XOR2_X1 U251 ( .A(n221), .B(n279), .Z(product[11]) );
  NAND2_X1 U252 ( .A1(n5), .A2(n20), .ZN(n280) );
  NAND2_X1 U253 ( .A1(n252), .A2(n23), .ZN(n281) );
  NAND2_X1 U254 ( .A1(n20), .A2(n23), .ZN(n282) );
  NAND3_X1 U255 ( .A1(n280), .A2(n281), .A3(n282), .ZN(n4) );
  CLKBUF_X1 U256 ( .A(b[0]), .Z(n283) );
  XOR2_X1 U257 ( .A(a[3]), .B(n306), .Z(n325) );
  XNOR2_X1 U258 ( .A(a[2]), .B(a[1]), .ZN(n324) );
  NAND2_X2 U259 ( .A1(n324), .A2(n362), .ZN(n326) );
  NAND2_X2 U260 ( .A1(n334), .A2(n363), .ZN(n336) );
  XOR2_X1 U261 ( .A(n34), .B(n39), .Z(n284) );
  XOR2_X1 U262 ( .A(n269), .B(n284), .Z(product[8]) );
  NAND2_X1 U263 ( .A1(n239), .A2(n34), .ZN(n285) );
  NAND2_X1 U264 ( .A1(n8), .A2(n39), .ZN(n286) );
  NAND2_X1 U265 ( .A1(n34), .A2(n39), .ZN(n287) );
  NAND3_X1 U266 ( .A1(n285), .A2(n286), .A3(n287), .ZN(n7) );
  NAND3_X1 U267 ( .A1(n302), .A2(n301), .A3(n300), .ZN(n288) );
  NAND3_X1 U268 ( .A1(n213), .A2(n258), .A3(n297), .ZN(n289) );
  XOR2_X1 U269 ( .A(a[2]), .B(n317), .Z(n290) );
  XOR2_X1 U270 ( .A(a[2]), .B(n317), .Z(n291) );
  XNOR2_X1 U271 ( .A(n278), .B(n292), .ZN(product[12]) );
  XNOR2_X1 U272 ( .A(n19), .B(n18), .ZN(n292) );
  XNOR2_X1 U273 ( .A(n298), .B(n293), .ZN(product[14]) );
  XNOR2_X1 U274 ( .A(n308), .B(n15), .ZN(n293) );
  INV_X1 U275 ( .A(n15), .ZN(n307) );
  AND3_X1 U276 ( .A1(n305), .A2(n304), .A3(n303), .ZN(product[15]) );
  INV_X1 U277 ( .A(n354), .ZN(n308) );
  INV_X1 U278 ( .A(n343), .ZN(n311) );
  INV_X1 U279 ( .A(n21), .ZN(n310) );
  INV_X1 U280 ( .A(n323), .ZN(n316) );
  INV_X1 U281 ( .A(n332), .ZN(n314) );
  INV_X1 U282 ( .A(n31), .ZN(n313) );
  INV_X1 U283 ( .A(b[0]), .ZN(n306) );
  INV_X1 U284 ( .A(a[0]), .ZN(n318) );
  INV_X1 U285 ( .A(a[5]), .ZN(n312) );
  INV_X1 U286 ( .A(a[7]), .ZN(n309) );
  NAND2_X1 U287 ( .A1(n4), .A2(n19), .ZN(n295) );
  NAND2_X1 U288 ( .A1(n231), .A2(n18), .ZN(n296) );
  NAND2_X1 U289 ( .A1(n19), .A2(n18), .ZN(n297) );
  NAND3_X1 U290 ( .A1(n296), .A2(n295), .A3(n297), .ZN(n3) );
  NAND3_X1 U291 ( .A1(n301), .A2(n302), .A3(n300), .ZN(n298) );
  INV_X1 U292 ( .A(a[3]), .ZN(n315) );
  XOR2_X1 U293 ( .A(n17), .B(n307), .Z(n299) );
  XOR2_X1 U294 ( .A(n299), .B(n289), .Z(product[13]) );
  NAND2_X1 U295 ( .A1(n17), .A2(n307), .ZN(n300) );
  NAND2_X1 U296 ( .A1(n3), .A2(n17), .ZN(n301) );
  NAND2_X1 U297 ( .A1(n215), .A2(n307), .ZN(n302) );
  NAND2_X1 U298 ( .A1(n308), .A2(n15), .ZN(n303) );
  NAND2_X1 U299 ( .A1(n308), .A2(n288), .ZN(n304) );
  NAND2_X1 U300 ( .A1(n15), .A2(n288), .ZN(n305) );
  INV_X1 U301 ( .A(a[1]), .ZN(n317) );
  NOR2_X1 U302 ( .A1(n318), .A2(n306), .ZN(product[0]) );
  OAI22_X1 U303 ( .A1(n319), .A2(n320), .B1(n321), .B2(n318), .ZN(n99) );
  OAI22_X1 U304 ( .A1(n321), .A2(n320), .B1(n322), .B2(n318), .ZN(n98) );
  XNOR2_X1 U305 ( .A(b[6]), .B(a[1]), .ZN(n321) );
  OAI22_X1 U306 ( .A1(n318), .A2(n322), .B1(n320), .B2(n322), .ZN(n323) );
  XNOR2_X1 U307 ( .A(b[7]), .B(a[1]), .ZN(n322) );
  NOR2_X1 U308 ( .A1(n290), .A2(n306), .ZN(n96) );
  OAI22_X1 U309 ( .A1(n325), .A2(n326), .B1(n291), .B2(n327), .ZN(n95) );
  OAI22_X1 U310 ( .A1(n327), .A2(n326), .B1(n291), .B2(n328), .ZN(n94) );
  XNOR2_X1 U311 ( .A(n209), .B(a[3]), .ZN(n327) );
  OAI22_X1 U312 ( .A1(n328), .A2(n326), .B1(n290), .B2(n329), .ZN(n93) );
  XNOR2_X1 U313 ( .A(b[2]), .B(a[3]), .ZN(n328) );
  OAI22_X1 U314 ( .A1(n329), .A2(n326), .B1(n291), .B2(n330), .ZN(n92) );
  XNOR2_X1 U315 ( .A(b[3]), .B(n210), .ZN(n329) );
  OAI22_X1 U316 ( .A1(n330), .A2(n326), .B1(n291), .B2(n331), .ZN(n91) );
  XNOR2_X1 U317 ( .A(b[4]), .B(a[3]), .ZN(n330) );
  OAI22_X1 U318 ( .A1(n333), .A2(n290), .B1(n326), .B2(n333), .ZN(n332) );
  NOR2_X1 U319 ( .A1(n334), .A2(n306), .ZN(n88) );
  OAI22_X1 U320 ( .A1(n335), .A2(n336), .B1(n334), .B2(n337), .ZN(n87) );
  XNOR2_X1 U321 ( .A(a[5]), .B(n283), .ZN(n335) );
  OAI22_X1 U322 ( .A1(n337), .A2(n336), .B1(n334), .B2(n338), .ZN(n86) );
  XNOR2_X1 U323 ( .A(n209), .B(a[5]), .ZN(n337) );
  OAI22_X1 U324 ( .A1(n338), .A2(n336), .B1(n334), .B2(n339), .ZN(n85) );
  XNOR2_X1 U325 ( .A(b[2]), .B(a[5]), .ZN(n338) );
  OAI22_X1 U326 ( .A1(n339), .A2(n336), .B1(n334), .B2(n340), .ZN(n84) );
  XNOR2_X1 U327 ( .A(b[3]), .B(a[5]), .ZN(n339) );
  OAI22_X1 U328 ( .A1(n340), .A2(n336), .B1(n334), .B2(n341), .ZN(n83) );
  XNOR2_X1 U329 ( .A(b[4]), .B(a[5]), .ZN(n340) );
  OAI22_X1 U330 ( .A1(n341), .A2(n336), .B1(n334), .B2(n342), .ZN(n82) );
  XNOR2_X1 U331 ( .A(b[5]), .B(a[5]), .ZN(n341) );
  OAI22_X1 U332 ( .A1(n344), .A2(n334), .B1(n336), .B2(n344), .ZN(n343) );
  NOR2_X1 U333 ( .A1(n345), .A2(n306), .ZN(n80) );
  OAI22_X1 U334 ( .A1(n346), .A2(n347), .B1(n218), .B2(n348), .ZN(n79) );
  XNOR2_X1 U335 ( .A(a[7]), .B(n283), .ZN(n346) );
  OAI22_X1 U336 ( .A1(n349), .A2(n347), .B1(n218), .B2(n350), .ZN(n77) );
  OAI22_X1 U337 ( .A1(n350), .A2(n347), .B1(n218), .B2(n351), .ZN(n76) );
  XNOR2_X1 U338 ( .A(b[3]), .B(a[7]), .ZN(n350) );
  OAI22_X1 U339 ( .A1(n351), .A2(n347), .B1(n218), .B2(n352), .ZN(n75) );
  XNOR2_X1 U340 ( .A(b[4]), .B(a[7]), .ZN(n351) );
  OAI22_X1 U341 ( .A1(n352), .A2(n347), .B1(n218), .B2(n353), .ZN(n74) );
  XNOR2_X1 U342 ( .A(b[5]), .B(a[7]), .ZN(n352) );
  OAI22_X1 U343 ( .A1(n355), .A2(n218), .B1(n347), .B2(n355), .ZN(n354) );
  OAI21_X1 U344 ( .B1(n283), .B2(n317), .A(n320), .ZN(n72) );
  OAI21_X1 U345 ( .B1(n315), .B2(n326), .A(n356), .ZN(n71) );
  OR3_X1 U346 ( .A1(n290), .A2(n283), .A3(n315), .ZN(n356) );
  OAI21_X1 U347 ( .B1(n312), .B2(n336), .A(n357), .ZN(n70) );
  OR3_X1 U348 ( .A1(n334), .A2(n283), .A3(n312), .ZN(n357) );
  OAI21_X1 U349 ( .B1(n309), .B2(n347), .A(n358), .ZN(n69) );
  OR3_X1 U350 ( .A1(n218), .A2(n283), .A3(n309), .ZN(n358) );
  XNOR2_X1 U351 ( .A(n359), .B(n360), .ZN(n38) );
  OR2_X1 U352 ( .A1(n359), .A2(n360), .ZN(n37) );
  OAI22_X1 U353 ( .A1(n331), .A2(n326), .B1(n290), .B2(n361), .ZN(n360) );
  XNOR2_X1 U354 ( .A(b[5]), .B(n210), .ZN(n331) );
  OAI22_X1 U355 ( .A1(n348), .A2(n347), .B1(n218), .B2(n349), .ZN(n359) );
  XNOR2_X1 U356 ( .A(b[2]), .B(a[7]), .ZN(n349) );
  XNOR2_X1 U357 ( .A(n219), .B(a[7]), .ZN(n348) );
  OAI22_X1 U358 ( .A1(n361), .A2(n326), .B1(n291), .B2(n333), .ZN(n31) );
  XNOR2_X1 U359 ( .A(b[7]), .B(n210), .ZN(n333) );
  XNOR2_X1 U360 ( .A(n315), .B(a[2]), .ZN(n362) );
  XNOR2_X1 U361 ( .A(b[6]), .B(n210), .ZN(n361) );
  OAI22_X1 U362 ( .A1(n342), .A2(n336), .B1(n334), .B2(n344), .ZN(n21) );
  XNOR2_X1 U363 ( .A(b[7]), .B(a[5]), .ZN(n344) );
  XNOR2_X1 U364 ( .A(n312), .B(a[4]), .ZN(n363) );
  XNOR2_X1 U365 ( .A(b[6]), .B(a[5]), .ZN(n342) );
  OAI22_X1 U366 ( .A1(n353), .A2(n347), .B1(n218), .B2(n355), .ZN(n15) );
  XNOR2_X1 U367 ( .A(b[7]), .B(a[7]), .ZN(n355) );
  NAND2_X1 U368 ( .A1(n345), .A2(n364), .ZN(n347) );
  XNOR2_X1 U369 ( .A(n309), .B(a[6]), .ZN(n364) );
  XNOR2_X1 U370 ( .A(b[6]), .B(a[7]), .ZN(n353) );
  OAI22_X1 U371 ( .A1(n283), .A2(n320), .B1(n365), .B2(n318), .ZN(n104) );
  OAI22_X1 U372 ( .A1(n365), .A2(n320), .B1(n366), .B2(n318), .ZN(n103) );
  OAI22_X1 U373 ( .A1(n366), .A2(n320), .B1(n367), .B2(n318), .ZN(n102) );
  XNOR2_X1 U374 ( .A(b[2]), .B(a[1]), .ZN(n366) );
  OAI22_X1 U375 ( .A1(n320), .A2(n367), .B1(n368), .B2(n318), .ZN(n101) );
  XNOR2_X1 U376 ( .A(b[3]), .B(a[1]), .ZN(n367) );
  OAI22_X1 U377 ( .A1(n368), .A2(n320), .B1(n319), .B2(n318), .ZN(n100) );
  XNOR2_X1 U378 ( .A(b[5]), .B(a[1]), .ZN(n319) );
  NAND2_X1 U379 ( .A1(a[1]), .A2(n318), .ZN(n320) );
  XNOR2_X1 U380 ( .A(b[4]), .B(a[1]), .ZN(n368) );
endmodule


module mac_24 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  mac_24_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_24_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_23_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;
  wire   [15:1] carry;

  XOR2_X1 U1 ( .A(B[15]), .B(A[15]), .Z(n1) );
  XOR2_X1 U2 ( .A(carry[15]), .B(n1), .Z(SUM[15]) );
  NAND3_X1 U3 ( .A1(n15), .A2(n16), .A3(n17), .ZN(n2) );
  NAND3_X1 U4 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n3) );
  AND2_X1 U5 ( .A1(B[0]), .A2(A[0]), .ZN(n4) );
  AND2_X1 U6 ( .A1(B[0]), .A2(A[0]), .ZN(n5) );
  AND2_X1 U7 ( .A1(B[0]), .A2(A[0]), .ZN(n77) );
  NAND3_X1 U8 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n6) );
  NAND3_X1 U9 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n7) );
  NAND3_X1 U10 ( .A1(n11), .A2(n12), .A3(n13), .ZN(n8) );
  NAND3_X1 U11 ( .A1(n11), .A2(n12), .A3(n13), .ZN(n9) );
  XOR2_X1 U12 ( .A(B[9]), .B(A[9]), .Z(n10) );
  XOR2_X1 U13 ( .A(n7), .B(n10), .Z(SUM[9]) );
  NAND2_X1 U14 ( .A1(n6), .A2(B[9]), .ZN(n11) );
  NAND2_X1 U15 ( .A1(carry[9]), .A2(A[9]), .ZN(n12) );
  NAND2_X1 U16 ( .A1(B[9]), .A2(A[9]), .ZN(n13) );
  NAND3_X1 U17 ( .A1(n11), .A2(n12), .A3(n13), .ZN(carry[10]) );
  XOR2_X1 U18 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR2_X1 U19 ( .A(n3), .B(n14), .Z(SUM[2]) );
  NAND2_X1 U20 ( .A1(n3), .A2(B[2]), .ZN(n15) );
  NAND2_X1 U21 ( .A1(carry[2]), .A2(A[2]), .ZN(n16) );
  NAND2_X1 U22 ( .A1(B[2]), .A2(A[2]), .ZN(n17) );
  NAND3_X1 U23 ( .A1(n15), .A2(n16), .A3(n17), .ZN(carry[3]) );
  NAND3_X1 U24 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n18) );
  NAND3_X1 U25 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n19) );
  XOR2_X1 U26 ( .A(B[10]), .B(A[10]), .Z(n20) );
  XOR2_X1 U27 ( .A(n9), .B(n20), .Z(SUM[10]) );
  NAND2_X1 U28 ( .A1(n8), .A2(B[10]), .ZN(n21) );
  NAND2_X1 U29 ( .A1(carry[10]), .A2(A[10]), .ZN(n22) );
  NAND2_X1 U30 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
  NAND3_X1 U31 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n24) );
  XOR2_X1 U32 ( .A(B[3]), .B(A[3]), .Z(n25) );
  XOR2_X1 U33 ( .A(n2), .B(n25), .Z(SUM[3]) );
  NAND2_X1 U34 ( .A1(n2), .A2(B[3]), .ZN(n26) );
  NAND2_X1 U35 ( .A1(carry[3]), .A2(A[3]), .ZN(n27) );
  NAND2_X1 U36 ( .A1(B[3]), .A2(A[3]), .ZN(n28) );
  NAND3_X1 U37 ( .A1(n27), .A2(n26), .A3(n28), .ZN(carry[4]) );
  NAND3_X1 U38 ( .A1(n31), .A2(n32), .A3(n33), .ZN(n29) );
  XOR2_X1 U39 ( .A(B[4]), .B(A[4]), .Z(n30) );
  XOR2_X1 U40 ( .A(n24), .B(n30), .Z(SUM[4]) );
  NAND2_X1 U41 ( .A1(n24), .A2(B[4]), .ZN(n31) );
  NAND2_X1 U42 ( .A1(carry[4]), .A2(A[4]), .ZN(n32) );
  NAND2_X1 U43 ( .A1(B[4]), .A2(A[4]), .ZN(n33) );
  NAND3_X1 U44 ( .A1(n31), .A2(n32), .A3(n33), .ZN(carry[5]) );
  NAND3_X1 U45 ( .A1(n39), .A2(n38), .A3(n40), .ZN(n34) );
  NAND3_X1 U46 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n35) );
  NAND3_X1 U47 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n36) );
  XOR2_X1 U48 ( .A(B[11]), .B(A[11]), .Z(n37) );
  XOR2_X1 U49 ( .A(n19), .B(n37), .Z(SUM[11]) );
  NAND2_X1 U50 ( .A1(n18), .A2(B[11]), .ZN(n38) );
  NAND2_X1 U51 ( .A1(n19), .A2(A[11]), .ZN(n39) );
  NAND2_X1 U52 ( .A1(B[11]), .A2(A[11]), .ZN(n40) );
  NAND3_X1 U53 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[12]) );
  XOR2_X1 U54 ( .A(B[5]), .B(A[5]), .Z(n41) );
  XOR2_X1 U55 ( .A(n29), .B(n41), .Z(SUM[5]) );
  NAND2_X1 U56 ( .A1(n29), .A2(B[5]), .ZN(n42) );
  NAND2_X1 U57 ( .A1(carry[5]), .A2(A[5]), .ZN(n43) );
  NAND2_X1 U58 ( .A1(B[5]), .A2(A[5]), .ZN(n44) );
  NAND3_X1 U59 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[6]) );
  NAND3_X1 U60 ( .A1(n48), .A2(n47), .A3(n49), .ZN(n45) );
  XOR2_X1 U61 ( .A(B[12]), .B(A[12]), .Z(n46) );
  XOR2_X1 U62 ( .A(n35), .B(n46), .Z(SUM[12]) );
  NAND2_X1 U63 ( .A1(n34), .A2(B[12]), .ZN(n47) );
  NAND2_X1 U64 ( .A1(carry[12]), .A2(A[12]), .ZN(n48) );
  NAND2_X1 U65 ( .A1(B[12]), .A2(A[12]), .ZN(n49) );
  NAND3_X1 U66 ( .A1(n47), .A2(n48), .A3(n49), .ZN(carry[13]) );
  NAND3_X1 U67 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n50) );
  NAND3_X1 U68 ( .A1(n67), .A2(n66), .A3(n68), .ZN(n51) );
  NAND3_X1 U69 ( .A1(n74), .A2(n75), .A3(n76), .ZN(n52) );
  XOR2_X1 U70 ( .A(B[8]), .B(A[8]), .Z(n53) );
  XOR2_X1 U71 ( .A(n52), .B(n53), .Z(SUM[8]) );
  NAND2_X1 U72 ( .A1(n52), .A2(B[8]), .ZN(n54) );
  NAND2_X1 U73 ( .A1(carry[8]), .A2(A[8]), .ZN(n55) );
  NAND2_X1 U74 ( .A1(B[8]), .A2(A[8]), .ZN(n56) );
  NAND3_X1 U75 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[9]) );
  XOR2_X1 U76 ( .A(B[1]), .B(A[1]), .Z(n57) );
  XOR2_X1 U77 ( .A(n5), .B(n57), .Z(SUM[1]) );
  NAND2_X1 U78 ( .A1(n4), .A2(B[1]), .ZN(n58) );
  NAND2_X1 U79 ( .A1(n77), .A2(A[1]), .ZN(n59) );
  NAND2_X1 U80 ( .A1(B[1]), .A2(A[1]), .ZN(n60) );
  NAND3_X1 U81 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[2]) );
  XOR2_X1 U82 ( .A(B[13]), .B(A[13]), .Z(n61) );
  XOR2_X1 U83 ( .A(n45), .B(n61), .Z(SUM[13]) );
  NAND2_X1 U84 ( .A1(n45), .A2(B[13]), .ZN(n62) );
  NAND2_X1 U85 ( .A1(carry[13]), .A2(A[13]), .ZN(n63) );
  NAND2_X1 U86 ( .A1(B[13]), .A2(A[13]), .ZN(n64) );
  NAND3_X1 U87 ( .A1(n62), .A2(n63), .A3(n64), .ZN(carry[14]) );
  XOR2_X1 U88 ( .A(B[6]), .B(A[6]), .Z(n65) );
  XOR2_X1 U89 ( .A(carry[6]), .B(n65), .Z(SUM[6]) );
  NAND2_X1 U90 ( .A1(n36), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U91 ( .A1(carry[6]), .A2(A[6]), .ZN(n67) );
  NAND2_X1 U92 ( .A1(B[6]), .A2(A[6]), .ZN(n68) );
  NAND3_X1 U93 ( .A1(n67), .A2(n66), .A3(n68), .ZN(carry[7]) );
  XOR2_X1 U94 ( .A(B[14]), .B(A[14]), .Z(n69) );
  XOR2_X1 U95 ( .A(n50), .B(n69), .Z(SUM[14]) );
  NAND2_X1 U96 ( .A1(n50), .A2(B[14]), .ZN(n70) );
  NAND2_X1 U97 ( .A1(carry[14]), .A2(A[14]), .ZN(n71) );
  NAND2_X1 U98 ( .A1(B[14]), .A2(A[14]), .ZN(n72) );
  NAND3_X1 U99 ( .A1(n70), .A2(n71), .A3(n72), .ZN(carry[15]) );
  XOR2_X1 U100 ( .A(B[7]), .B(A[7]), .Z(n73) );
  XOR2_X1 U101 ( .A(n51), .B(n73), .Z(SUM[7]) );
  NAND2_X1 U102 ( .A1(n51), .A2(B[7]), .ZN(n74) );
  NAND2_X1 U103 ( .A1(carry[7]), .A2(A[7]), .ZN(n75) );
  NAND2_X1 U104 ( .A1(B[7]), .A2(A[7]), .ZN(n76) );
  NAND3_X1 U105 ( .A1(n74), .A2(n75), .A3(n76), .ZN(carry[8]) );
  XOR2_X1 U106 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_23_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n311), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n310), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n314), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n313), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n316), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n88), .B(n101), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n102), .B(n95), .CO(n55), .S(n56) );
  NAND3_X1 U157 ( .A1(n299), .A2(n300), .A3(n301), .ZN(n49) );
  NAND2_X1 U158 ( .A1(n279), .A2(n17), .ZN(n206) );
  CLKBUF_X1 U159 ( .A(n365), .Z(n207) );
  NAND2_X1 U160 ( .A1(n255), .A2(n34), .ZN(n208) );
  XOR2_X1 U161 ( .A(n102), .B(n95), .Z(n209) );
  CLKBUF_X1 U162 ( .A(n209), .Z(n210) );
  CLKBUF_X1 U163 ( .A(n267), .Z(n211) );
  INV_X1 U164 ( .A(n305), .ZN(n212) );
  XOR2_X1 U165 ( .A(a[3]), .B(a[2]), .Z(n362) );
  NAND2_X2 U166 ( .A1(n285), .A2(n286), .ZN(n213) );
  NAND2_X1 U167 ( .A1(n285), .A2(n286), .ZN(n324) );
  INV_X1 U168 ( .A(n315), .ZN(n214) );
  BUF_X2 U169 ( .A(a[1]), .Z(n289) );
  XNOR2_X1 U170 ( .A(n221), .B(n215), .ZN(product[14]) );
  XNOR2_X1 U171 ( .A(n308), .B(n15), .ZN(n215) );
  AND3_X1 U172 ( .A1(n223), .A2(n222), .A3(n224), .ZN(product[15]) );
  INV_X1 U173 ( .A(n306), .ZN(n217) );
  INV_X1 U174 ( .A(n306), .ZN(n305) );
  AND2_X1 U175 ( .A1(n104), .A2(n72), .ZN(n218) );
  NAND2_X1 U176 ( .A1(n239), .A2(n33), .ZN(n219) );
  NAND3_X1 U177 ( .A1(n206), .A2(n294), .A3(n296), .ZN(n220) );
  NAND3_X1 U178 ( .A1(n294), .A2(n206), .A3(n296), .ZN(n221) );
  CLKBUF_X1 U179 ( .A(b[1]), .Z(n265) );
  NAND2_X1 U180 ( .A1(n2), .A2(n308), .ZN(n222) );
  NAND2_X1 U181 ( .A1(n220), .A2(n15), .ZN(n223) );
  NAND2_X1 U182 ( .A1(n308), .A2(n15), .ZN(n224) );
  NAND2_X2 U183 ( .A1(n345), .A2(n364), .ZN(n347) );
  XOR2_X2 U184 ( .A(a[6]), .B(n312), .Z(n345) );
  NAND2_X1 U185 ( .A1(n7), .A2(n28), .ZN(n225) );
  NAND3_X1 U186 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n226) );
  NAND3_X1 U187 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n227) );
  NAND3_X1 U188 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n228) );
  NAND3_X1 U189 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n229) );
  CLKBUF_X1 U190 ( .A(n260), .Z(n230) );
  CLKBUF_X1 U191 ( .A(n228), .Z(n231) );
  NAND3_X1 U192 ( .A1(n219), .A2(n225), .A3(n244), .ZN(n232) );
  NAND3_X1 U193 ( .A1(n219), .A2(n225), .A3(n244), .ZN(n233) );
  CLKBUF_X1 U194 ( .A(n268), .Z(n234) );
  XOR2_X1 U195 ( .A(n27), .B(n24), .Z(n235) );
  XOR2_X1 U196 ( .A(n233), .B(n235), .Z(product[10]) );
  NAND2_X1 U197 ( .A1(n232), .A2(n27), .ZN(n236) );
  NAND2_X1 U198 ( .A1(n6), .A2(n24), .ZN(n237) );
  NAND2_X1 U199 ( .A1(n27), .A2(n24), .ZN(n238) );
  NAND3_X1 U200 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n5) );
  NAND3_X1 U201 ( .A1(n208), .A2(n260), .A3(n261), .ZN(n239) );
  NAND3_X1 U202 ( .A1(n208), .A2(n230), .A3(n261), .ZN(n240) );
  XOR2_X1 U203 ( .A(n33), .B(n28), .Z(n241) );
  XOR2_X1 U204 ( .A(n240), .B(n241), .Z(product[9]) );
  NAND2_X1 U205 ( .A1(n239), .A2(n33), .ZN(n242) );
  NAND2_X1 U206 ( .A1(n7), .A2(n28), .ZN(n243) );
  NAND2_X1 U207 ( .A1(n33), .A2(n28), .ZN(n244) );
  NAND3_X1 U208 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n6) );
  NAND3_X1 U209 ( .A1(n302), .A2(n304), .A3(n303), .ZN(n245) );
  NAND3_X1 U210 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n246) );
  XOR2_X1 U211 ( .A(n103), .B(n96), .Z(n247) );
  XOR2_X1 U212 ( .A(n218), .B(n247), .Z(product[2]) );
  NAND2_X1 U213 ( .A1(n218), .A2(n103), .ZN(n248) );
  NAND2_X1 U214 ( .A1(n14), .A2(n96), .ZN(n249) );
  NAND2_X1 U215 ( .A1(n103), .A2(n96), .ZN(n250) );
  NAND3_X1 U216 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n13) );
  XOR2_X1 U217 ( .A(n210), .B(n71), .Z(n251) );
  XOR2_X1 U218 ( .A(n227), .B(n251), .Z(product[3]) );
  NAND2_X1 U219 ( .A1(n227), .A2(n209), .ZN(n252) );
  NAND2_X1 U220 ( .A1(n13), .A2(n71), .ZN(n253) );
  NAND2_X1 U221 ( .A1(n56), .A2(n71), .ZN(n254) );
  NAND3_X1 U222 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n12) );
  NAND3_X1 U223 ( .A1(n267), .A2(n268), .A3(n269), .ZN(n255) );
  NAND3_X1 U224 ( .A1(n211), .A2(n234), .A3(n269), .ZN(n256) );
  NAND3_X1 U225 ( .A1(n281), .A2(n282), .A3(n283), .ZN(n257) );
  XOR2_X1 U226 ( .A(n34), .B(n39), .Z(n258) );
  XOR2_X1 U227 ( .A(n256), .B(n258), .Z(product[8]) );
  NAND2_X1 U228 ( .A1(n255), .A2(n34), .ZN(n259) );
  NAND2_X1 U229 ( .A1(n8), .A2(n39), .ZN(n260) );
  NAND2_X1 U230 ( .A1(n34), .A2(n39), .ZN(n261) );
  NAND3_X1 U231 ( .A1(n260), .A2(n259), .A3(n261), .ZN(n7) );
  CLKBUF_X1 U232 ( .A(n226), .Z(n262) );
  NAND3_X1 U233 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n263) );
  NAND3_X1 U234 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n264) );
  XOR2_X1 U235 ( .A(n40), .B(n45), .Z(n266) );
  XOR2_X1 U236 ( .A(n262), .B(n266), .Z(product[7]) );
  NAND2_X1 U237 ( .A1(n226), .A2(n40), .ZN(n267) );
  NAND2_X1 U238 ( .A1(n246), .A2(n45), .ZN(n268) );
  NAND2_X1 U239 ( .A1(n40), .A2(n45), .ZN(n269) );
  NAND3_X1 U240 ( .A1(n267), .A2(n268), .A3(n269), .ZN(n8) );
  XOR2_X1 U241 ( .A(n54), .B(n55), .Z(n270) );
  XOR2_X1 U242 ( .A(n12), .B(n270), .Z(product[4]) );
  NAND2_X1 U243 ( .A1(n54), .A2(n229), .ZN(n271) );
  NAND2_X1 U244 ( .A1(n12), .A2(n55), .ZN(n272) );
  NAND2_X1 U245 ( .A1(n54), .A2(n55), .ZN(n273) );
  NAND3_X1 U246 ( .A1(n272), .A2(n271), .A3(n273), .ZN(n11) );
  CLKBUF_X1 U247 ( .A(n245), .Z(n274) );
  XOR2_X1 U248 ( .A(n46), .B(n49), .Z(n275) );
  XOR2_X1 U249 ( .A(n274), .B(n275), .Z(product[6]) );
  NAND2_X1 U250 ( .A1(n245), .A2(n46), .ZN(n276) );
  NAND2_X1 U251 ( .A1(n10), .A2(n49), .ZN(n277) );
  NAND2_X1 U252 ( .A1(n46), .A2(n49), .ZN(n278) );
  NAND3_X1 U253 ( .A1(n293), .A2(n292), .A3(n291), .ZN(n279) );
  XNOR2_X2 U254 ( .A(a[4]), .B(a[3]), .ZN(n334) );
  XOR2_X1 U255 ( .A(n23), .B(n20), .Z(n280) );
  XOR2_X1 U256 ( .A(n231), .B(n280), .Z(product[11]) );
  NAND2_X1 U257 ( .A1(n228), .A2(n23), .ZN(n281) );
  NAND2_X1 U258 ( .A1(n5), .A2(n20), .ZN(n282) );
  NAND2_X1 U259 ( .A1(n23), .A2(n20), .ZN(n283) );
  NAND3_X1 U260 ( .A1(n281), .A2(n282), .A3(n283), .ZN(n4) );
  NAND2_X1 U261 ( .A1(a[2]), .A2(n289), .ZN(n285) );
  NAND2_X1 U262 ( .A1(n284), .A2(n317), .ZN(n286) );
  INV_X1 U263 ( .A(a[2]), .ZN(n284) );
  NAND2_X2 U264 ( .A1(n324), .A2(n362), .ZN(n326) );
  XOR2_X1 U265 ( .A(n297), .B(n52), .Z(n50) );
  XNOR2_X1 U266 ( .A(n287), .B(n288), .ZN(product[13]) );
  XNOR2_X1 U267 ( .A(n17), .B(n307), .ZN(n287) );
  INV_X1 U268 ( .A(n15), .ZN(n307) );
  INV_X1 U269 ( .A(n332), .ZN(n314) );
  INV_X1 U270 ( .A(n343), .ZN(n311) );
  INV_X1 U271 ( .A(n21), .ZN(n310) );
  INV_X1 U272 ( .A(n323), .ZN(n316) );
  INV_X1 U273 ( .A(n31), .ZN(n313) );
  INV_X1 U274 ( .A(b[0]), .ZN(n306) );
  INV_X1 U275 ( .A(n354), .ZN(n308) );
  INV_X1 U276 ( .A(a[0]), .ZN(n318) );
  INV_X1 U277 ( .A(a[3]), .ZN(n315) );
  INV_X1 U278 ( .A(a[5]), .ZN(n312) );
  INV_X1 U279 ( .A(a[7]), .ZN(n309) );
  NAND3_X1 U280 ( .A1(n293), .A2(n292), .A3(n291), .ZN(n288) );
  XOR2_X1 U281 ( .A(n19), .B(n18), .Z(n290) );
  XOR2_X1 U282 ( .A(n290), .B(n257), .Z(product[12]) );
  NAND2_X1 U283 ( .A1(n19), .A2(n18), .ZN(n291) );
  NAND2_X1 U284 ( .A1(n19), .A2(n4), .ZN(n292) );
  NAND2_X1 U285 ( .A1(n18), .A2(n4), .ZN(n293) );
  NAND3_X1 U286 ( .A1(n293), .A2(n292), .A3(n291), .ZN(n3) );
  NAND2_X1 U287 ( .A1(n17), .A2(n307), .ZN(n294) );
  NAND2_X1 U288 ( .A1(n279), .A2(n17), .ZN(n295) );
  NAND2_X1 U289 ( .A1(n307), .A2(n3), .ZN(n296) );
  NAND3_X1 U290 ( .A1(n296), .A2(n295), .A3(n294), .ZN(n2) );
  XOR2_X1 U291 ( .A(n93), .B(n100), .Z(n297) );
  XOR2_X1 U292 ( .A(n53), .B(n264), .Z(n298) );
  XOR2_X1 U293 ( .A(n298), .B(n50), .Z(product[5]) );
  NAND2_X1 U294 ( .A1(n93), .A2(n100), .ZN(n299) );
  NAND2_X1 U295 ( .A1(n93), .A2(n52), .ZN(n300) );
  NAND2_X1 U296 ( .A1(n100), .A2(n52), .ZN(n301) );
  NAND2_X1 U297 ( .A1(n53), .A2(n263), .ZN(n302) );
  NAND2_X1 U298 ( .A1(n53), .A2(n50), .ZN(n303) );
  NAND2_X1 U299 ( .A1(n11), .A2(n50), .ZN(n304) );
  NAND3_X1 U300 ( .A1(n302), .A2(n303), .A3(n304), .ZN(n10) );
  INV_X1 U301 ( .A(a[1]), .ZN(n317) );
  NOR2_X1 U302 ( .A1(n318), .A2(n212), .ZN(product[0]) );
  OAI22_X1 U303 ( .A1(n319), .A2(n320), .B1(n321), .B2(n318), .ZN(n99) );
  OAI22_X1 U304 ( .A1(n321), .A2(n320), .B1(n322), .B2(n318), .ZN(n98) );
  XNOR2_X1 U305 ( .A(b[6]), .B(n289), .ZN(n321) );
  OAI22_X1 U306 ( .A1(n318), .A2(n322), .B1(n320), .B2(n322), .ZN(n323) );
  XNOR2_X1 U307 ( .A(b[7]), .B(n289), .ZN(n322) );
  NOR2_X1 U308 ( .A1(n213), .A2(n306), .ZN(n96) );
  OAI22_X1 U309 ( .A1(n325), .A2(n326), .B1(n213), .B2(n327), .ZN(n95) );
  XNOR2_X1 U310 ( .A(a[3]), .B(n305), .ZN(n325) );
  OAI22_X1 U311 ( .A1(n327), .A2(n326), .B1(n213), .B2(n328), .ZN(n94) );
  XNOR2_X1 U312 ( .A(b[1]), .B(a[3]), .ZN(n327) );
  OAI22_X1 U313 ( .A1(n328), .A2(n326), .B1(n213), .B2(n329), .ZN(n93) );
  XNOR2_X1 U314 ( .A(b[2]), .B(a[3]), .ZN(n328) );
  OAI22_X1 U315 ( .A1(n329), .A2(n326), .B1(n213), .B2(n330), .ZN(n92) );
  XNOR2_X1 U316 ( .A(b[3]), .B(n214), .ZN(n329) );
  OAI22_X1 U317 ( .A1(n330), .A2(n326), .B1(n213), .B2(n331), .ZN(n91) );
  XNOR2_X1 U318 ( .A(b[4]), .B(a[3]), .ZN(n330) );
  OAI22_X1 U319 ( .A1(n333), .A2(n213), .B1(n326), .B2(n333), .ZN(n332) );
  NOR2_X1 U320 ( .A1(n334), .A2(n212), .ZN(n88) );
  OAI22_X1 U321 ( .A1(n335), .A2(n336), .B1(n334), .B2(n337), .ZN(n87) );
  XNOR2_X1 U322 ( .A(a[5]), .B(n217), .ZN(n335) );
  OAI22_X1 U323 ( .A1(n337), .A2(n336), .B1(n334), .B2(n338), .ZN(n86) );
  XNOR2_X1 U324 ( .A(n265), .B(a[5]), .ZN(n337) );
  OAI22_X1 U325 ( .A1(n338), .A2(n336), .B1(n334), .B2(n339), .ZN(n85) );
  XNOR2_X1 U326 ( .A(b[2]), .B(a[5]), .ZN(n338) );
  OAI22_X1 U327 ( .A1(n339), .A2(n336), .B1(n334), .B2(n340), .ZN(n84) );
  XNOR2_X1 U328 ( .A(b[3]), .B(a[5]), .ZN(n339) );
  OAI22_X1 U329 ( .A1(n340), .A2(n336), .B1(n334), .B2(n341), .ZN(n83) );
  XNOR2_X1 U330 ( .A(b[4]), .B(a[5]), .ZN(n340) );
  OAI22_X1 U331 ( .A1(n341), .A2(n336), .B1(n334), .B2(n342), .ZN(n82) );
  XNOR2_X1 U332 ( .A(b[5]), .B(a[5]), .ZN(n341) );
  OAI22_X1 U333 ( .A1(n344), .A2(n334), .B1(n336), .B2(n344), .ZN(n343) );
  NOR2_X1 U334 ( .A1(n345), .A2(n212), .ZN(n80) );
  OAI22_X1 U335 ( .A1(n346), .A2(n347), .B1(n345), .B2(n348), .ZN(n79) );
  XNOR2_X1 U336 ( .A(a[7]), .B(n217), .ZN(n346) );
  OAI22_X1 U337 ( .A1(n349), .A2(n347), .B1(n345), .B2(n350), .ZN(n77) );
  OAI22_X1 U338 ( .A1(n350), .A2(n347), .B1(n345), .B2(n351), .ZN(n76) );
  XNOR2_X1 U339 ( .A(b[3]), .B(a[7]), .ZN(n350) );
  OAI22_X1 U340 ( .A1(n351), .A2(n347), .B1(n345), .B2(n352), .ZN(n75) );
  XNOR2_X1 U341 ( .A(b[4]), .B(a[7]), .ZN(n351) );
  OAI22_X1 U342 ( .A1(n352), .A2(n347), .B1(n345), .B2(n353), .ZN(n74) );
  XNOR2_X1 U343 ( .A(b[5]), .B(a[7]), .ZN(n352) );
  OAI22_X1 U344 ( .A1(n355), .A2(n345), .B1(n347), .B2(n355), .ZN(n354) );
  OAI21_X1 U345 ( .B1(n305), .B2(n317), .A(n320), .ZN(n72) );
  OAI21_X1 U346 ( .B1(n315), .B2(n326), .A(n356), .ZN(n71) );
  OR3_X1 U347 ( .A1(n213), .A2(n217), .A3(n315), .ZN(n356) );
  OAI21_X1 U348 ( .B1(n312), .B2(n336), .A(n357), .ZN(n70) );
  OR3_X1 U349 ( .A1(n334), .A2(n217), .A3(n312), .ZN(n357) );
  OAI21_X1 U350 ( .B1(n309), .B2(n347), .A(n358), .ZN(n69) );
  OR3_X1 U351 ( .A1(n345), .A2(n217), .A3(n309), .ZN(n358) );
  XNOR2_X1 U352 ( .A(n359), .B(n360), .ZN(n38) );
  OR2_X1 U353 ( .A1(n359), .A2(n360), .ZN(n37) );
  OAI22_X1 U354 ( .A1(n331), .A2(n326), .B1(n213), .B2(n361), .ZN(n360) );
  XNOR2_X1 U355 ( .A(b[5]), .B(n214), .ZN(n331) );
  OAI22_X1 U356 ( .A1(n348), .A2(n347), .B1(n345), .B2(n349), .ZN(n359) );
  XNOR2_X1 U357 ( .A(b[2]), .B(a[7]), .ZN(n349) );
  XNOR2_X1 U358 ( .A(n265), .B(a[7]), .ZN(n348) );
  OAI22_X1 U359 ( .A1(n361), .A2(n326), .B1(n213), .B2(n333), .ZN(n31) );
  XNOR2_X1 U360 ( .A(b[7]), .B(n214), .ZN(n333) );
  XNOR2_X1 U361 ( .A(b[6]), .B(n214), .ZN(n361) );
  OAI22_X1 U362 ( .A1(n342), .A2(n336), .B1(n334), .B2(n344), .ZN(n21) );
  XNOR2_X1 U363 ( .A(b[7]), .B(a[5]), .ZN(n344) );
  NAND2_X1 U364 ( .A1(n334), .A2(n363), .ZN(n336) );
  XNOR2_X1 U365 ( .A(n312), .B(a[4]), .ZN(n363) );
  XNOR2_X1 U366 ( .A(b[6]), .B(a[5]), .ZN(n342) );
  OAI22_X1 U367 ( .A1(n353), .A2(n347), .B1(n345), .B2(n355), .ZN(n15) );
  XNOR2_X1 U368 ( .A(b[7]), .B(a[7]), .ZN(n355) );
  XNOR2_X1 U369 ( .A(n309), .B(a[6]), .ZN(n364) );
  XNOR2_X1 U370 ( .A(b[6]), .B(a[7]), .ZN(n353) );
  OAI22_X1 U371 ( .A1(n217), .A2(n320), .B1(n365), .B2(n318), .ZN(n104) );
  OAI22_X1 U372 ( .A1(n207), .A2(n320), .B1(n366), .B2(n318), .ZN(n103) );
  XNOR2_X1 U373 ( .A(b[1]), .B(n289), .ZN(n365) );
  OAI22_X1 U374 ( .A1(n366), .A2(n320), .B1(n367), .B2(n318), .ZN(n102) );
  XNOR2_X1 U375 ( .A(b[2]), .B(n289), .ZN(n366) );
  OAI22_X1 U376 ( .A1(n367), .A2(n320), .B1(n368), .B2(n318), .ZN(n101) );
  XNOR2_X1 U377 ( .A(b[3]), .B(n289), .ZN(n367) );
  OAI22_X1 U378 ( .A1(n368), .A2(n320), .B1(n319), .B2(n318), .ZN(n100) );
  XNOR2_X1 U379 ( .A(b[5]), .B(n289), .ZN(n319) );
  NAND2_X1 U380 ( .A1(n289), .A2(n318), .ZN(n320) );
  XNOR2_X1 U381 ( .A(b[4]), .B(n289), .ZN(n368) );
endmodule


module mac_23 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_23_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_23_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X2 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_22_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74;
  wire   [15:1] carry;

  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n74) );
  XOR2_X1 U2 ( .A(B[15]), .B(A[15]), .Z(n1) );
  XOR2_X1 U3 ( .A(carry[15]), .B(n1), .Z(SUM[15]) );
  NAND3_X1 U4 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n2) );
  NAND3_X1 U5 ( .A1(n9), .A2(n10), .A3(n11), .ZN(n3) );
  XOR2_X1 U6 ( .A(B[4]), .B(A[4]), .Z(n4) );
  XOR2_X1 U7 ( .A(carry[4]), .B(n4), .Z(SUM[4]) );
  NAND2_X1 U8 ( .A1(carry[4]), .A2(B[4]), .ZN(n5) );
  NAND2_X1 U9 ( .A1(carry[4]), .A2(A[4]), .ZN(n6) );
  NAND2_X1 U10 ( .A1(B[4]), .A2(A[4]), .ZN(n7) );
  NAND3_X1 U11 ( .A1(n5), .A2(n6), .A3(n7), .ZN(carry[5]) );
  XOR2_X1 U12 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR2_X1 U13 ( .A(carry[5]), .B(n8), .Z(SUM[5]) );
  NAND2_X1 U14 ( .A1(carry[5]), .A2(B[5]), .ZN(n9) );
  NAND2_X1 U15 ( .A1(carry[5]), .A2(A[5]), .ZN(n10) );
  NAND2_X1 U16 ( .A1(B[5]), .A2(A[5]), .ZN(n11) );
  NAND3_X1 U17 ( .A1(n9), .A2(n10), .A3(n11), .ZN(carry[6]) );
  NAND3_X1 U18 ( .A1(n71), .A2(n72), .A3(n73), .ZN(n12) );
  XOR2_X1 U19 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR2_X1 U20 ( .A(n12), .B(n13), .Z(SUM[3]) );
  NAND2_X1 U21 ( .A1(n12), .A2(B[3]), .ZN(n14) );
  NAND2_X1 U22 ( .A1(carry[3]), .A2(A[3]), .ZN(n15) );
  NAND2_X1 U23 ( .A1(B[3]), .A2(A[3]), .ZN(n16) );
  NAND3_X1 U24 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[4]) );
  NAND3_X1 U25 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n17) );
  XOR2_X1 U26 ( .A(B[6]), .B(A[6]), .Z(n18) );
  XOR2_X1 U27 ( .A(n3), .B(n18), .Z(SUM[6]) );
  NAND2_X1 U28 ( .A1(n3), .A2(B[6]), .ZN(n19) );
  NAND2_X1 U29 ( .A1(carry[6]), .A2(A[6]), .ZN(n20) );
  NAND2_X1 U30 ( .A1(B[6]), .A2(A[6]), .ZN(n21) );
  NAND3_X1 U31 ( .A1(n19), .A2(n20), .A3(n21), .ZN(carry[7]) );
  NAND3_X1 U32 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n22) );
  NAND3_X1 U33 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n23) );
  NAND3_X1 U34 ( .A1(n32), .A2(n33), .A3(n34), .ZN(n24) );
  NAND3_X1 U35 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n25) );
  NAND3_X1 U36 ( .A1(n48), .A2(n47), .A3(n49), .ZN(n26) );
  XOR2_X1 U37 ( .A(B[7]), .B(A[7]), .Z(n27) );
  XOR2_X1 U38 ( .A(n2), .B(n27), .Z(SUM[7]) );
  NAND2_X1 U39 ( .A1(n2), .A2(B[7]), .ZN(n28) );
  NAND2_X1 U40 ( .A1(carry[7]), .A2(A[7]), .ZN(n29) );
  NAND2_X1 U41 ( .A1(B[7]), .A2(A[7]), .ZN(n30) );
  NAND3_X1 U42 ( .A1(n29), .A2(n28), .A3(n30), .ZN(carry[8]) );
  XOR2_X1 U43 ( .A(B[13]), .B(A[13]), .Z(n31) );
  XOR2_X1 U44 ( .A(n23), .B(n31), .Z(SUM[13]) );
  NAND2_X1 U45 ( .A1(n22), .A2(B[13]), .ZN(n32) );
  NAND2_X1 U46 ( .A1(carry[13]), .A2(A[13]), .ZN(n33) );
  NAND2_X1 U47 ( .A1(B[13]), .A2(A[13]), .ZN(n34) );
  NAND3_X1 U48 ( .A1(n33), .A2(n32), .A3(n34), .ZN(carry[14]) );
  NAND3_X1 U49 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n35) );
  XOR2_X1 U50 ( .A(B[12]), .B(A[12]), .Z(n36) );
  XOR2_X1 U51 ( .A(n35), .B(n36), .Z(SUM[12]) );
  NAND2_X1 U52 ( .A1(n17), .A2(B[12]), .ZN(n37) );
  NAND2_X1 U53 ( .A1(carry[12]), .A2(A[12]), .ZN(n38) );
  NAND2_X1 U54 ( .A1(B[12]), .A2(A[12]), .ZN(n39) );
  NAND3_X1 U55 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[13]) );
  XOR2_X1 U56 ( .A(B[14]), .B(A[14]), .Z(n40) );
  XOR2_X1 U57 ( .A(n24), .B(n40), .Z(SUM[14]) );
  NAND2_X1 U58 ( .A1(n24), .A2(B[14]), .ZN(n41) );
  NAND2_X1 U59 ( .A1(carry[14]), .A2(A[14]), .ZN(n42) );
  NAND2_X1 U60 ( .A1(B[14]), .A2(A[14]), .ZN(n43) );
  NAND3_X1 U61 ( .A1(n41), .A2(n42), .A3(n43), .ZN(carry[15]) );
  NAND3_X1 U62 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n44) );
  NAND3_X1 U63 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n45) );
  XOR2_X1 U64 ( .A(B[10]), .B(A[10]), .Z(n46) );
  XOR2_X1 U65 ( .A(n45), .B(n46), .Z(SUM[10]) );
  NAND2_X1 U66 ( .A1(n44), .A2(B[10]), .ZN(n47) );
  NAND2_X1 U67 ( .A1(n44), .A2(A[10]), .ZN(n48) );
  NAND2_X1 U68 ( .A1(B[10]), .A2(A[10]), .ZN(n49) );
  NAND3_X1 U69 ( .A1(n47), .A2(n48), .A3(n49), .ZN(carry[11]) );
  XOR2_X1 U70 ( .A(B[11]), .B(A[11]), .Z(n50) );
  XOR2_X1 U71 ( .A(n26), .B(n50), .Z(SUM[11]) );
  NAND2_X1 U72 ( .A1(n26), .A2(B[11]), .ZN(n51) );
  NAND2_X1 U73 ( .A1(carry[11]), .A2(A[11]), .ZN(n52) );
  NAND2_X1 U74 ( .A1(B[11]), .A2(A[11]), .ZN(n53) );
  NAND3_X1 U75 ( .A1(n51), .A2(n52), .A3(n53), .ZN(carry[12]) );
  NAND3_X1 U76 ( .A1(n67), .A2(n68), .A3(n69), .ZN(n54) );
  NAND3_X1 U77 ( .A1(n67), .A2(n68), .A3(n69), .ZN(n55) );
  NAND3_X1 U78 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n56) );
  NAND3_X1 U79 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n57) );
  XOR2_X1 U80 ( .A(B[8]), .B(A[8]), .Z(n58) );
  XOR2_X1 U81 ( .A(n25), .B(n58), .Z(SUM[8]) );
  NAND2_X1 U82 ( .A1(n25), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U83 ( .A1(carry[8]), .A2(A[8]), .ZN(n60) );
  NAND2_X1 U84 ( .A1(B[8]), .A2(A[8]), .ZN(n61) );
  NAND3_X1 U85 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[9]) );
  XOR2_X1 U86 ( .A(B[9]), .B(A[9]), .Z(n62) );
  XOR2_X1 U87 ( .A(n57), .B(n62), .Z(SUM[9]) );
  NAND2_X1 U88 ( .A1(n56), .A2(B[9]), .ZN(n63) );
  NAND2_X1 U89 ( .A1(carry[9]), .A2(A[9]), .ZN(n64) );
  NAND2_X1 U90 ( .A1(B[9]), .A2(A[9]), .ZN(n65) );
  XOR2_X1 U91 ( .A(B[1]), .B(A[1]), .Z(n66) );
  XOR2_X1 U92 ( .A(n74), .B(n66), .Z(SUM[1]) );
  NAND2_X1 U93 ( .A1(n74), .A2(B[1]), .ZN(n67) );
  NAND2_X1 U94 ( .A1(n74), .A2(A[1]), .ZN(n68) );
  NAND2_X1 U95 ( .A1(B[1]), .A2(A[1]), .ZN(n69) );
  NAND3_X1 U96 ( .A1(n67), .A2(n68), .A3(n69), .ZN(carry[2]) );
  XOR2_X1 U97 ( .A(B[2]), .B(A[2]), .Z(n70) );
  XOR2_X1 U98 ( .A(n55), .B(n70), .Z(SUM[2]) );
  NAND2_X1 U99 ( .A1(n54), .A2(B[2]), .ZN(n71) );
  NAND2_X1 U100 ( .A1(carry[2]), .A2(A[2]), .ZN(n72) );
  NAND2_X1 U101 ( .A1(B[2]), .A2(A[2]), .ZN(n73) );
  NAND3_X1 U102 ( .A1(n71), .A2(n72), .A3(n73), .ZN(carry[3]) );
  XOR2_X1 U103 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_22_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n302), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n301), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n305), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n304), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n307), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  NAND3_X1 U157 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n206) );
  NAND3_X1 U158 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n207) );
  NAND2_X1 U159 ( .A1(n325), .A2(n354), .ZN(n327) );
  AND2_X1 U160 ( .A1(n235), .A2(n102), .ZN(n208) );
  NAND3_X1 U161 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n209) );
  XOR2_X1 U162 ( .A(a[5]), .B(a[4]), .Z(n354) );
  NAND3_X1 U163 ( .A1(n274), .A2(n273), .A3(n275), .ZN(n210) );
  NAND3_X1 U164 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n211) );
  CLKBUF_X1 U165 ( .A(n209), .Z(n212) );
  NAND3_X1 U166 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n213) );
  NAND3_X1 U167 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n214) );
  XOR2_X1 U168 ( .A(a[3]), .B(n297), .Z(n316) );
  BUF_X1 U169 ( .A(b[0]), .Z(n288) );
  NAND3_X1 U170 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n215) );
  CLKBUF_X1 U171 ( .A(n287), .Z(n216) );
  NAND2_X1 U172 ( .A1(n14), .A2(n96), .ZN(n217) );
  NAND2_X1 U173 ( .A1(n14), .A2(n96), .ZN(n218) );
  CLKBUF_X1 U174 ( .A(n211), .Z(n219) );
  CLKBUF_X1 U175 ( .A(n241), .Z(n220) );
  NAND3_X1 U176 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n221) );
  XOR2_X1 U177 ( .A(n46), .B(n49), .Z(n222) );
  XOR2_X1 U178 ( .A(n10), .B(n222), .Z(product[6]) );
  NAND2_X1 U179 ( .A1(n207), .A2(n46), .ZN(n223) );
  NAND2_X1 U180 ( .A1(n206), .A2(n49), .ZN(n224) );
  NAND2_X1 U181 ( .A1(n46), .A2(n49), .ZN(n225) );
  NAND3_X1 U182 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n9) );
  CLKBUF_X1 U183 ( .A(n254), .Z(n226) );
  XOR2_X1 U184 ( .A(n40), .B(n45), .Z(n227) );
  XOR2_X1 U185 ( .A(n212), .B(n227), .Z(product[7]) );
  NAND2_X1 U186 ( .A1(n209), .A2(n40), .ZN(n228) );
  NAND2_X1 U187 ( .A1(n9), .A2(n45), .ZN(n229) );
  NAND2_X1 U188 ( .A1(n40), .A2(n45), .ZN(n230) );
  NAND3_X1 U189 ( .A1(n229), .A2(n228), .A3(n230), .ZN(n8) );
  XOR2_X1 U190 ( .A(n34), .B(n39), .Z(n231) );
  XOR2_X1 U191 ( .A(n219), .B(n231), .Z(product[8]) );
  NAND2_X1 U192 ( .A1(n211), .A2(n34), .ZN(n232) );
  NAND2_X1 U193 ( .A1(n8), .A2(n39), .ZN(n233) );
  NAND2_X1 U194 ( .A1(n34), .A2(n39), .ZN(n234) );
  NAND3_X1 U195 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n7) );
  OAI22_X1 U196 ( .A1(n316), .A2(n317), .B1(n276), .B2(n318), .ZN(n235) );
  NAND3_X1 U197 ( .A1(n241), .A2(n240), .A3(n242), .ZN(n236) );
  XOR2_X1 U198 ( .A(n95), .B(n102), .Z(n56) );
  CLKBUF_X1 U199 ( .A(b[1]), .Z(n237) );
  CLKBUF_X1 U200 ( .A(n273), .Z(n238) );
  XOR2_X1 U201 ( .A(n33), .B(n28), .Z(n239) );
  XOR2_X1 U202 ( .A(n214), .B(n239), .Z(product[9]) );
  NAND2_X1 U203 ( .A1(n213), .A2(n33), .ZN(n240) );
  NAND2_X1 U204 ( .A1(n7), .A2(n28), .ZN(n241) );
  NAND2_X1 U205 ( .A1(n33), .A2(n28), .ZN(n242) );
  NAND3_X1 U206 ( .A1(n240), .A2(n220), .A3(n242), .ZN(n6) );
  NAND3_X1 U207 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n243) );
  NAND3_X1 U208 ( .A1(n251), .A2(n218), .A3(n253), .ZN(n244) );
  AND2_X1 U209 ( .A1(n104), .A2(n72), .ZN(n245) );
  XNOR2_X1 U210 ( .A(a[4]), .B(a[3]), .ZN(n246) );
  XNOR2_X1 U211 ( .A(a[4]), .B(a[3]), .ZN(n325) );
  CLKBUF_X1 U212 ( .A(n264), .Z(n247) );
  AND3_X1 U213 ( .A1(n286), .A2(n285), .A3(n284), .ZN(product[15]) );
  XNOR2_X1 U214 ( .A(n249), .B(n279), .ZN(product[14]) );
  XNOR2_X1 U215 ( .A(n299), .B(n15), .ZN(n249) );
  XOR2_X1 U216 ( .A(n103), .B(n96), .Z(n250) );
  XOR2_X1 U217 ( .A(n245), .B(n250), .Z(product[2]) );
  NAND2_X1 U218 ( .A1(n245), .A2(n103), .ZN(n251) );
  NAND2_X1 U219 ( .A1(n14), .A2(n96), .ZN(n252) );
  NAND2_X1 U220 ( .A1(n103), .A2(n96), .ZN(n253) );
  NAND3_X1 U221 ( .A1(n251), .A2(n217), .A3(n253), .ZN(n13) );
  NAND3_X1 U222 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n254) );
  XOR2_X1 U223 ( .A(n27), .B(n24), .Z(n255) );
  XOR2_X1 U224 ( .A(n6), .B(n255), .Z(product[10]) );
  NAND2_X1 U225 ( .A1(n236), .A2(n27), .ZN(n256) );
  NAND2_X1 U226 ( .A1(n215), .A2(n24), .ZN(n257) );
  NAND2_X1 U227 ( .A1(n27), .A2(n24), .ZN(n258) );
  NAND3_X1 U228 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n5) );
  NAND3_X1 U229 ( .A1(n268), .A2(n269), .A3(n270), .ZN(n259) );
  NAND3_X1 U230 ( .A1(n268), .A2(n269), .A3(n270), .ZN(n260) );
  NAND3_X1 U231 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n261) );
  NAND3_X1 U232 ( .A1(n247), .A2(n265), .A3(n266), .ZN(n262) );
  XOR2_X1 U233 ( .A(n23), .B(n20), .Z(n263) );
  XOR2_X1 U234 ( .A(n226), .B(n263), .Z(product[11]) );
  NAND2_X1 U235 ( .A1(n254), .A2(n23), .ZN(n264) );
  NAND2_X1 U236 ( .A1(n5), .A2(n20), .ZN(n265) );
  NAND2_X1 U237 ( .A1(n23), .A2(n20), .ZN(n266) );
  XOR2_X1 U238 ( .A(n56), .B(n71), .Z(n267) );
  XOR2_X1 U239 ( .A(n244), .B(n267), .Z(product[3]) );
  NAND2_X1 U240 ( .A1(n13), .A2(n56), .ZN(n268) );
  NAND2_X1 U241 ( .A1(n243), .A2(n71), .ZN(n269) );
  NAND2_X1 U242 ( .A1(n56), .A2(n71), .ZN(n270) );
  NAND3_X1 U243 ( .A1(n268), .A2(n269), .A3(n270), .ZN(n12) );
  NAND3_X1 U244 ( .A1(n238), .A2(n274), .A3(n275), .ZN(n271) );
  XOR2_X1 U245 ( .A(n18), .B(n19), .Z(n272) );
  XOR2_X1 U246 ( .A(n262), .B(n272), .Z(product[12]) );
  NAND2_X1 U247 ( .A1(n261), .A2(n18), .ZN(n273) );
  NAND2_X1 U248 ( .A1(n221), .A2(n19), .ZN(n274) );
  NAND2_X1 U249 ( .A1(n18), .A2(n19), .ZN(n275) );
  NAND3_X1 U250 ( .A1(n274), .A2(n273), .A3(n275), .ZN(n3) );
  XNOR2_X1 U251 ( .A(a[2]), .B(a[1]), .ZN(n276) );
  XNOR2_X1 U252 ( .A(a[2]), .B(a[1]), .ZN(n277) );
  XNOR2_X1 U253 ( .A(a[2]), .B(a[1]), .ZN(n315) );
  NAND3_X1 U254 ( .A1(n282), .A2(n283), .A3(n281), .ZN(n278) );
  NAND3_X1 U255 ( .A1(n282), .A2(n283), .A3(n281), .ZN(n279) );
  XOR2_X1 U256 ( .A(n17), .B(n298), .Z(n280) );
  XOR2_X1 U257 ( .A(n280), .B(n271), .Z(product[13]) );
  NAND2_X1 U258 ( .A1(n17), .A2(n298), .ZN(n281) );
  NAND2_X1 U259 ( .A1(n17), .A2(n210), .ZN(n282) );
  NAND2_X1 U260 ( .A1(n3), .A2(n298), .ZN(n283) );
  NAND3_X1 U261 ( .A1(n282), .A2(n283), .A3(n281), .ZN(n2) );
  NAND2_X1 U262 ( .A1(n299), .A2(n15), .ZN(n284) );
  NAND2_X1 U263 ( .A1(n2), .A2(n299), .ZN(n285) );
  NAND2_X1 U264 ( .A1(n278), .A2(n15), .ZN(n286) );
  NAND3_X1 U265 ( .A1(n290), .A2(n291), .A3(n292), .ZN(n287) );
  INV_X1 U266 ( .A(n15), .ZN(n298) );
  INV_X1 U267 ( .A(n21), .ZN(n301) );
  INV_X1 U268 ( .A(n334), .ZN(n302) );
  INV_X1 U269 ( .A(n314), .ZN(n307) );
  INV_X1 U270 ( .A(n323), .ZN(n305) );
  INV_X1 U271 ( .A(b[0]), .ZN(n297) );
  INV_X1 U272 ( .A(n345), .ZN(n299) );
  INV_X1 U273 ( .A(n31), .ZN(n304) );
  INV_X1 U274 ( .A(a[0]), .ZN(n309) );
  INV_X1 U275 ( .A(a[5]), .ZN(n303) );
  INV_X1 U276 ( .A(a[7]), .ZN(n300) );
  XOR2_X1 U277 ( .A(n54), .B(n208), .Z(n289) );
  XOR2_X1 U278 ( .A(n260), .B(n289), .Z(product[4]) );
  NAND2_X1 U279 ( .A1(n259), .A2(n54), .ZN(n290) );
  NAND2_X1 U280 ( .A1(n12), .A2(n208), .ZN(n291) );
  NAND2_X1 U281 ( .A1(n54), .A2(n208), .ZN(n292) );
  NAND3_X1 U282 ( .A1(n291), .A2(n290), .A3(n292), .ZN(n11) );
  XOR2_X1 U283 ( .A(n50), .B(n53), .Z(n293) );
  XOR2_X1 U284 ( .A(n216), .B(n293), .Z(product[5]) );
  NAND2_X1 U285 ( .A1(n287), .A2(n50), .ZN(n294) );
  NAND2_X1 U286 ( .A1(n11), .A2(n53), .ZN(n295) );
  NAND2_X1 U287 ( .A1(n50), .A2(n53), .ZN(n296) );
  NAND3_X1 U288 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n10) );
  INV_X1 U289 ( .A(a[3]), .ZN(n306) );
  INV_X1 U290 ( .A(a[1]), .ZN(n308) );
  NAND2_X2 U291 ( .A1(n315), .A2(n353), .ZN(n317) );
  XOR2_X2 U292 ( .A(a[6]), .B(n303), .Z(n336) );
  NOR2_X1 U293 ( .A1(n309), .A2(n297), .ZN(product[0]) );
  OAI22_X1 U294 ( .A1(n310), .A2(n311), .B1(n312), .B2(n309), .ZN(n99) );
  OAI22_X1 U295 ( .A1(n312), .A2(n311), .B1(n313), .B2(n309), .ZN(n98) );
  XNOR2_X1 U296 ( .A(b[6]), .B(a[1]), .ZN(n312) );
  OAI22_X1 U297 ( .A1(n309), .A2(n313), .B1(n311), .B2(n313), .ZN(n314) );
  XNOR2_X1 U298 ( .A(b[7]), .B(a[1]), .ZN(n313) );
  NOR2_X1 U299 ( .A1(n277), .A2(n297), .ZN(n96) );
  OAI22_X1 U300 ( .A1(n316), .A2(n317), .B1(n276), .B2(n318), .ZN(n95) );
  OAI22_X1 U301 ( .A1(n318), .A2(n317), .B1(n276), .B2(n319), .ZN(n94) );
  XNOR2_X1 U302 ( .A(b[1]), .B(a[3]), .ZN(n318) );
  OAI22_X1 U303 ( .A1(n319), .A2(n317), .B1(n276), .B2(n320), .ZN(n93) );
  XNOR2_X1 U304 ( .A(b[2]), .B(a[3]), .ZN(n319) );
  OAI22_X1 U305 ( .A1(n320), .A2(n317), .B1(n277), .B2(n321), .ZN(n92) );
  XNOR2_X1 U306 ( .A(b[3]), .B(a[3]), .ZN(n320) );
  OAI22_X1 U307 ( .A1(n321), .A2(n317), .B1(n277), .B2(n322), .ZN(n91) );
  XNOR2_X1 U308 ( .A(b[4]), .B(a[3]), .ZN(n321) );
  OAI22_X1 U309 ( .A1(n324), .A2(n276), .B1(n317), .B2(n324), .ZN(n323) );
  NOR2_X1 U310 ( .A1(n246), .A2(n297), .ZN(n88) );
  OAI22_X1 U311 ( .A1(n326), .A2(n327), .B1(n246), .B2(n328), .ZN(n87) );
  XNOR2_X1 U312 ( .A(a[5]), .B(n288), .ZN(n326) );
  OAI22_X1 U313 ( .A1(n328), .A2(n327), .B1(n246), .B2(n329), .ZN(n86) );
  XNOR2_X1 U314 ( .A(n237), .B(a[5]), .ZN(n328) );
  OAI22_X1 U315 ( .A1(n329), .A2(n327), .B1(n246), .B2(n330), .ZN(n85) );
  XNOR2_X1 U316 ( .A(b[2]), .B(a[5]), .ZN(n329) );
  OAI22_X1 U317 ( .A1(n330), .A2(n327), .B1(n246), .B2(n331), .ZN(n84) );
  XNOR2_X1 U318 ( .A(b[3]), .B(a[5]), .ZN(n330) );
  OAI22_X1 U319 ( .A1(n331), .A2(n327), .B1(n246), .B2(n332), .ZN(n83) );
  XNOR2_X1 U320 ( .A(b[4]), .B(a[5]), .ZN(n331) );
  OAI22_X1 U321 ( .A1(n332), .A2(n327), .B1(n246), .B2(n333), .ZN(n82) );
  XNOR2_X1 U322 ( .A(b[5]), .B(a[5]), .ZN(n332) );
  OAI22_X1 U323 ( .A1(n335), .A2(n246), .B1(n327), .B2(n335), .ZN(n334) );
  NOR2_X1 U324 ( .A1(n336), .A2(n297), .ZN(n80) );
  OAI22_X1 U325 ( .A1(n337), .A2(n338), .B1(n336), .B2(n339), .ZN(n79) );
  XNOR2_X1 U326 ( .A(a[7]), .B(n288), .ZN(n337) );
  OAI22_X1 U327 ( .A1(n340), .A2(n338), .B1(n336), .B2(n341), .ZN(n77) );
  OAI22_X1 U328 ( .A1(n341), .A2(n338), .B1(n336), .B2(n342), .ZN(n76) );
  XNOR2_X1 U329 ( .A(b[3]), .B(a[7]), .ZN(n341) );
  OAI22_X1 U330 ( .A1(n342), .A2(n338), .B1(n336), .B2(n343), .ZN(n75) );
  XNOR2_X1 U331 ( .A(b[4]), .B(a[7]), .ZN(n342) );
  OAI22_X1 U332 ( .A1(n343), .A2(n338), .B1(n336), .B2(n344), .ZN(n74) );
  XNOR2_X1 U333 ( .A(b[5]), .B(a[7]), .ZN(n343) );
  OAI22_X1 U334 ( .A1(n346), .A2(n336), .B1(n338), .B2(n346), .ZN(n345) );
  OAI21_X1 U335 ( .B1(n288), .B2(n308), .A(n311), .ZN(n72) );
  OAI21_X1 U336 ( .B1(n306), .B2(n317), .A(n347), .ZN(n71) );
  OR3_X1 U337 ( .A1(n277), .A2(n288), .A3(n306), .ZN(n347) );
  OAI21_X1 U338 ( .B1(n303), .B2(n327), .A(n348), .ZN(n70) );
  OR3_X1 U339 ( .A1(n246), .A2(n288), .A3(n303), .ZN(n348) );
  OAI21_X1 U340 ( .B1(n300), .B2(n338), .A(n349), .ZN(n69) );
  OR3_X1 U341 ( .A1(n336), .A2(n288), .A3(n300), .ZN(n349) );
  XNOR2_X1 U342 ( .A(n350), .B(n351), .ZN(n38) );
  OR2_X1 U343 ( .A1(n350), .A2(n351), .ZN(n37) );
  OAI22_X1 U344 ( .A1(n322), .A2(n317), .B1(n276), .B2(n352), .ZN(n351) );
  XNOR2_X1 U345 ( .A(b[5]), .B(a[3]), .ZN(n322) );
  OAI22_X1 U346 ( .A1(n339), .A2(n338), .B1(n336), .B2(n340), .ZN(n350) );
  XNOR2_X1 U347 ( .A(b[2]), .B(a[7]), .ZN(n340) );
  XNOR2_X1 U348 ( .A(n237), .B(a[7]), .ZN(n339) );
  OAI22_X1 U349 ( .A1(n352), .A2(n317), .B1(n277), .B2(n324), .ZN(n31) );
  XNOR2_X1 U350 ( .A(b[7]), .B(a[3]), .ZN(n324) );
  XNOR2_X1 U351 ( .A(n306), .B(a[2]), .ZN(n353) );
  XNOR2_X1 U352 ( .A(b[6]), .B(a[3]), .ZN(n352) );
  OAI22_X1 U353 ( .A1(n333), .A2(n327), .B1(n246), .B2(n335), .ZN(n21) );
  XNOR2_X1 U354 ( .A(b[7]), .B(a[5]), .ZN(n335) );
  XNOR2_X1 U355 ( .A(b[6]), .B(a[5]), .ZN(n333) );
  OAI22_X1 U356 ( .A1(n344), .A2(n338), .B1(n336), .B2(n346), .ZN(n15) );
  XNOR2_X1 U357 ( .A(b[7]), .B(a[7]), .ZN(n346) );
  NAND2_X1 U358 ( .A1(n336), .A2(n355), .ZN(n338) );
  XNOR2_X1 U359 ( .A(n300), .B(a[6]), .ZN(n355) );
  XNOR2_X1 U360 ( .A(b[6]), .B(a[7]), .ZN(n344) );
  OAI22_X1 U361 ( .A1(n288), .A2(n311), .B1(n356), .B2(n309), .ZN(n104) );
  OAI22_X1 U362 ( .A1(n356), .A2(n311), .B1(n309), .B2(n357), .ZN(n103) );
  XNOR2_X1 U363 ( .A(b[1]), .B(a[1]), .ZN(n356) );
  OAI22_X1 U364 ( .A1(n357), .A2(n311), .B1(n358), .B2(n309), .ZN(n102) );
  XNOR2_X1 U365 ( .A(b[2]), .B(a[1]), .ZN(n357) );
  OAI22_X1 U366 ( .A1(n358), .A2(n311), .B1(n359), .B2(n309), .ZN(n101) );
  XNOR2_X1 U367 ( .A(b[3]), .B(a[1]), .ZN(n358) );
  OAI22_X1 U368 ( .A1(n359), .A2(n311), .B1(n310), .B2(n309), .ZN(n100) );
  XNOR2_X1 U369 ( .A(b[5]), .B(a[1]), .ZN(n310) );
  NAND2_X1 U370 ( .A1(a[1]), .A2(n309), .ZN(n311) );
  XNOR2_X1 U371 ( .A(b[4]), .B(a[1]), .ZN(n359) );
endmodule


module mac_22 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  mac_22_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_22_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_21_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65;
  wire   [15:1] carry;

  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CLKBUF_X1 U1 ( .A(carry[10]), .Z(n1) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n65) );
  NAND3_X1 U3 ( .A1(n8), .A2(n9), .A3(n10), .ZN(n2) );
  NAND3_X1 U4 ( .A1(n8), .A2(n9), .A3(n10), .ZN(n3) );
  XOR2_X1 U5 ( .A(B[15]), .B(A[15]), .Z(n4) );
  XOR2_X1 U6 ( .A(carry[15]), .B(n4), .Z(SUM[15]) );
  CLKBUF_X1 U7 ( .A(n62), .Z(n5) );
  CLKBUF_X1 U8 ( .A(n37), .Z(n6) );
  XOR2_X1 U9 ( .A(B[10]), .B(A[10]), .Z(n7) );
  XOR2_X1 U10 ( .A(n1), .B(n7), .Z(SUM[10]) );
  NAND2_X1 U11 ( .A1(carry[10]), .A2(B[10]), .ZN(n8) );
  NAND2_X1 U12 ( .A1(carry[10]), .A2(A[10]), .ZN(n9) );
  NAND2_X1 U13 ( .A1(B[10]), .A2(A[10]), .ZN(n10) );
  NAND3_X1 U14 ( .A1(n8), .A2(n9), .A3(n10), .ZN(carry[11]) );
  NAND3_X1 U15 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n11) );
  NAND3_X1 U16 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n12) );
  NAND3_X1 U17 ( .A1(n5), .A2(n63), .A3(n64), .ZN(n13) );
  NAND3_X1 U18 ( .A1(n18), .A2(n17), .A3(n19), .ZN(n14) );
  NAND3_X1 U19 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n15) );
  XOR2_X1 U20 ( .A(B[1]), .B(A[1]), .Z(n16) );
  XOR2_X1 U21 ( .A(n65), .B(n16), .Z(SUM[1]) );
  NAND2_X1 U22 ( .A1(n65), .A2(B[1]), .ZN(n17) );
  NAND2_X1 U23 ( .A1(n65), .A2(A[1]), .ZN(n18) );
  NAND2_X1 U24 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  NAND3_X1 U25 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[2]) );
  XOR2_X1 U26 ( .A(B[2]), .B(A[2]), .Z(n20) );
  XOR2_X1 U27 ( .A(carry[2]), .B(n20), .Z(SUM[2]) );
  NAND2_X1 U28 ( .A1(n14), .A2(B[2]), .ZN(n21) );
  NAND2_X1 U29 ( .A1(carry[2]), .A2(A[2]), .ZN(n22) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(n23) );
  NAND3_X1 U31 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[3]) );
  XOR2_X1 U32 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR2_X1 U33 ( .A(n13), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U34 ( .A1(n12), .A2(B[8]), .ZN(n25) );
  NAND2_X1 U35 ( .A1(carry[8]), .A2(A[8]), .ZN(n26) );
  NAND2_X1 U36 ( .A1(B[8]), .A2(A[8]), .ZN(n27) );
  NAND3_X1 U37 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[9]) );
  CLKBUF_X1 U38 ( .A(n48), .Z(n28) );
  XOR2_X1 U39 ( .A(B[11]), .B(A[11]), .Z(n29) );
  XOR2_X1 U40 ( .A(n3), .B(n29), .Z(SUM[11]) );
  NAND2_X1 U41 ( .A1(n2), .A2(B[11]), .ZN(n30) );
  NAND2_X1 U42 ( .A1(carry[11]), .A2(A[11]), .ZN(n31) );
  NAND2_X1 U43 ( .A1(B[11]), .A2(A[11]), .ZN(n32) );
  NAND3_X1 U44 ( .A1(n30), .A2(n31), .A3(n32), .ZN(carry[12]) );
  XOR2_X1 U45 ( .A(B[4]), .B(A[4]), .Z(n33) );
  XOR2_X1 U46 ( .A(carry[4]), .B(n33), .Z(SUM[4]) );
  NAND2_X1 U47 ( .A1(carry[4]), .A2(B[4]), .ZN(n34) );
  NAND2_X1 U48 ( .A1(carry[4]), .A2(A[4]), .ZN(n35) );
  NAND2_X1 U49 ( .A1(B[4]), .A2(A[4]), .ZN(n36) );
  NAND3_X1 U50 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[5]) );
  NAND3_X1 U51 ( .A1(n40), .A2(n41), .A3(n42), .ZN(n37) );
  NAND3_X1 U52 ( .A1(n44), .A2(n45), .A3(n46), .ZN(n38) );
  XOR2_X1 U53 ( .A(B[12]), .B(A[12]), .Z(n39) );
  XOR2_X1 U54 ( .A(n11), .B(n39), .Z(SUM[12]) );
  NAND2_X1 U55 ( .A1(n11), .A2(B[12]), .ZN(n40) );
  NAND2_X1 U56 ( .A1(carry[12]), .A2(A[12]), .ZN(n41) );
  NAND2_X1 U57 ( .A1(B[12]), .A2(A[12]), .ZN(n42) );
  NAND3_X1 U58 ( .A1(n40), .A2(n41), .A3(n42), .ZN(carry[13]) );
  XOR2_X1 U59 ( .A(B[5]), .B(A[5]), .Z(n43) );
  XOR2_X1 U60 ( .A(carry[5]), .B(n43), .Z(SUM[5]) );
  NAND2_X1 U61 ( .A1(n15), .A2(B[5]), .ZN(n44) );
  NAND2_X1 U62 ( .A1(n15), .A2(A[5]), .ZN(n45) );
  NAND2_X1 U63 ( .A1(B[5]), .A2(A[5]), .ZN(n46) );
  NAND3_X1 U64 ( .A1(n44), .A2(n45), .A3(n46), .ZN(carry[6]) );
  NAND3_X1 U65 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n47) );
  NAND3_X1 U66 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n48) );
  XOR2_X1 U67 ( .A(B[13]), .B(A[13]), .Z(n49) );
  XOR2_X1 U68 ( .A(n6), .B(n49), .Z(SUM[13]) );
  NAND2_X1 U69 ( .A1(n37), .A2(B[13]), .ZN(n50) );
  NAND2_X1 U70 ( .A1(carry[13]), .A2(A[13]), .ZN(n51) );
  NAND2_X1 U71 ( .A1(B[13]), .A2(A[13]), .ZN(n52) );
  NAND3_X1 U72 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[14]) );
  XOR2_X1 U73 ( .A(B[6]), .B(A[6]), .Z(n53) );
  XOR2_X1 U74 ( .A(carry[6]), .B(n53), .Z(SUM[6]) );
  NAND2_X1 U75 ( .A1(n38), .A2(B[6]), .ZN(n54) );
  NAND2_X1 U76 ( .A1(n38), .A2(A[6]), .ZN(n55) );
  NAND2_X1 U77 ( .A1(B[6]), .A2(A[6]), .ZN(n56) );
  NAND3_X1 U78 ( .A1(n55), .A2(n54), .A3(n56), .ZN(carry[7]) );
  XOR2_X1 U79 ( .A(B[14]), .B(A[14]), .Z(n57) );
  XOR2_X1 U80 ( .A(carry[14]), .B(n57), .Z(SUM[14]) );
  NAND2_X1 U81 ( .A1(n47), .A2(B[14]), .ZN(n58) );
  NAND2_X1 U82 ( .A1(n47), .A2(A[14]), .ZN(n59) );
  NAND2_X1 U83 ( .A1(B[14]), .A2(A[14]), .ZN(n60) );
  NAND3_X1 U84 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[15]) );
  XOR2_X1 U85 ( .A(B[7]), .B(A[7]), .Z(n61) );
  XOR2_X1 U86 ( .A(n28), .B(n61), .Z(SUM[7]) );
  NAND2_X1 U87 ( .A1(n48), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U88 ( .A1(carry[7]), .A2(A[7]), .ZN(n63) );
  NAND2_X1 U89 ( .A1(B[7]), .A2(A[7]), .ZN(n64) );
  NAND3_X1 U90 ( .A1(n62), .A2(n63), .A3(n64), .ZN(carry[8]) );
  XOR2_X1 U91 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_21_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n309), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n308), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n312), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n311), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n314), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  BUF_X2 U157 ( .A(n322), .Z(n221) );
  NAND3_X1 U158 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n49) );
  INV_X1 U159 ( .A(n15), .ZN(n305) );
  AND2_X1 U160 ( .A1(n95), .A2(n102), .ZN(n206) );
  CLKBUF_X1 U161 ( .A(n222), .Z(n207) );
  NAND2_X1 U162 ( .A1(n253), .A2(n50), .ZN(n208) );
  CLKBUF_X1 U163 ( .A(n253), .Z(n209) );
  CLKBUF_X1 U164 ( .A(n232), .Z(n210) );
  INV_X1 U165 ( .A(n315), .ZN(n211) );
  CLKBUF_X1 U166 ( .A(n262), .Z(n212) );
  CLKBUF_X1 U167 ( .A(n258), .Z(n213) );
  CLKBUF_X1 U168 ( .A(n250), .Z(n214) );
  CLKBUF_X1 U169 ( .A(n263), .Z(n215) );
  INV_X1 U170 ( .A(n304), .ZN(n216) );
  INV_X1 U171 ( .A(n304), .ZN(n217) );
  INV_X1 U172 ( .A(n304), .ZN(n303) );
  CLKBUF_X1 U173 ( .A(n14), .Z(n218) );
  CLKBUF_X1 U174 ( .A(n208), .Z(n219) );
  NAND2_X1 U175 ( .A1(n5), .A2(n20), .ZN(n220) );
  XNOR2_X1 U176 ( .A(a[2]), .B(a[1]), .ZN(n322) );
  NAND2_X1 U177 ( .A1(n265), .A2(n19), .ZN(n222) );
  NAND3_X1 U178 ( .A1(n208), .A2(n284), .A3(n285), .ZN(n223) );
  NAND3_X1 U179 ( .A1(n219), .A2(n284), .A3(n285), .ZN(n224) );
  NAND3_X1 U180 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n225) );
  NAND3_X1 U181 ( .A1(n261), .A2(n212), .A3(n215), .ZN(n226) );
  NAND3_X1 U182 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n227) );
  XOR2_X1 U183 ( .A(n46), .B(n49), .Z(n228) );
  XOR2_X1 U184 ( .A(n224), .B(n228), .Z(product[6]) );
  NAND2_X1 U185 ( .A1(n223), .A2(n46), .ZN(n229) );
  NAND2_X1 U186 ( .A1(n10), .A2(n49), .ZN(n230) );
  NAND2_X1 U187 ( .A1(n46), .A2(n49), .ZN(n231) );
  NAND3_X1 U188 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n9) );
  NAND3_X1 U189 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n232) );
  NAND3_X1 U190 ( .A1(n259), .A2(n258), .A3(n257), .ZN(n233) );
  NAND3_X1 U191 ( .A1(n257), .A2(n213), .A3(n259), .ZN(n234) );
  XOR2_X1 U192 ( .A(n40), .B(n45), .Z(n235) );
  XOR2_X1 U193 ( .A(n9), .B(n235), .Z(product[7]) );
  NAND2_X1 U194 ( .A1(n227), .A2(n40), .ZN(n236) );
  NAND2_X1 U195 ( .A1(n9), .A2(n45), .ZN(n237) );
  NAND2_X1 U196 ( .A1(n40), .A2(n45), .ZN(n238) );
  NAND3_X1 U197 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n8) );
  XOR2_X1 U198 ( .A(n93), .B(n100), .Z(n239) );
  XOR2_X1 U199 ( .A(n52), .B(n239), .Z(n50) );
  NAND2_X1 U200 ( .A1(n52), .A2(n93), .ZN(n240) );
  NAND2_X1 U201 ( .A1(n52), .A2(n100), .ZN(n241) );
  NAND2_X1 U202 ( .A1(n93), .A2(n100), .ZN(n242) );
  NAND3_X1 U203 ( .A1(n287), .A2(n288), .A3(n289), .ZN(n243) );
  CLKBUF_X1 U204 ( .A(n220), .Z(n244) );
  NAND3_X1 U205 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n245) );
  NAND3_X1 U206 ( .A1(n214), .A2(n251), .A3(n252), .ZN(n246) );
  NAND3_X1 U207 ( .A1(n222), .A2(n301), .A3(n302), .ZN(n247) );
  CLKBUF_X1 U208 ( .A(n5), .Z(n248) );
  XOR2_X1 U209 ( .A(n34), .B(n39), .Z(n249) );
  XOR2_X1 U210 ( .A(n210), .B(n249), .Z(product[8]) );
  NAND2_X1 U211 ( .A1(n232), .A2(n34), .ZN(n250) );
  NAND2_X1 U212 ( .A1(n8), .A2(n39), .ZN(n251) );
  NAND2_X1 U213 ( .A1(n34), .A2(n39), .ZN(n252) );
  NAND3_X1 U214 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n7) );
  NAND3_X1 U215 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n253) );
  NAND3_X1 U216 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n254) );
  XNOR2_X1 U217 ( .A(b[1]), .B(n211), .ZN(n255) );
  NAND2_X2 U218 ( .A1(n332), .A2(n361), .ZN(n334) );
  XOR2_X1 U219 ( .A(n103), .B(n96), .Z(n256) );
  XOR2_X1 U220 ( .A(n256), .B(n218), .Z(product[2]) );
  NAND2_X1 U221 ( .A1(n103), .A2(n96), .ZN(n257) );
  NAND2_X1 U222 ( .A1(n103), .A2(n14), .ZN(n258) );
  NAND2_X1 U223 ( .A1(n96), .A2(n14), .ZN(n259) );
  NAND3_X1 U224 ( .A1(n259), .A2(n258), .A3(n257), .ZN(n13) );
  XOR2_X1 U225 ( .A(n56), .B(n71), .Z(n260) );
  XOR2_X1 U226 ( .A(n260), .B(n234), .Z(product[3]) );
  NAND2_X1 U227 ( .A1(n56), .A2(n71), .ZN(n261) );
  NAND2_X1 U228 ( .A1(n56), .A2(n233), .ZN(n262) );
  NAND2_X1 U229 ( .A1(n71), .A2(n13), .ZN(n263) );
  NAND3_X1 U230 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n12) );
  CLKBUF_X1 U231 ( .A(n301), .Z(n264) );
  NAND3_X1 U232 ( .A1(n220), .A2(n271), .A3(n272), .ZN(n265) );
  NAND3_X1 U233 ( .A1(n271), .A2(n244), .A3(n272), .ZN(n266) );
  NAND3_X1 U234 ( .A1(n301), .A2(n300), .A3(n302), .ZN(n267) );
  NAND3_X1 U235 ( .A1(n291), .A2(n292), .A3(n293), .ZN(n268) );
  NAND3_X1 U236 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n269) );
  XOR2_X1 U237 ( .A(n23), .B(n20), .Z(n270) );
  XOR2_X1 U238 ( .A(n248), .B(n270), .Z(product[11]) );
  NAND2_X1 U239 ( .A1(n268), .A2(n23), .ZN(n271) );
  NAND2_X1 U240 ( .A1(n23), .A2(n20), .ZN(n272) );
  NAND3_X1 U241 ( .A1(n220), .A2(n271), .A3(n272), .ZN(n4) );
  XOR2_X1 U242 ( .A(n17), .B(n305), .Z(n273) );
  XOR2_X1 U243 ( .A(n3), .B(n273), .Z(product[13]) );
  NAND2_X1 U244 ( .A1(n247), .A2(n17), .ZN(n274) );
  NAND2_X1 U245 ( .A1(n267), .A2(n305), .ZN(n275) );
  NAND2_X1 U246 ( .A1(n17), .A2(n305), .ZN(n276) );
  XOR2_X1 U247 ( .A(n54), .B(n206), .Z(n277) );
  XOR2_X1 U248 ( .A(n226), .B(n277), .Z(product[4]) );
  NAND2_X1 U249 ( .A1(n225), .A2(n54), .ZN(n278) );
  NAND2_X1 U250 ( .A1(n12), .A2(n206), .ZN(n279) );
  NAND2_X1 U251 ( .A1(n54), .A2(n206), .ZN(n280) );
  NAND3_X1 U252 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n11) );
  NAND3_X1 U253 ( .A1(n288), .A2(n287), .A3(n289), .ZN(n281) );
  XOR2_X1 U254 ( .A(n50), .B(n53), .Z(n282) );
  XOR2_X1 U255 ( .A(n209), .B(n282), .Z(product[5]) );
  NAND2_X1 U256 ( .A1(n253), .A2(n50), .ZN(n283) );
  NAND2_X1 U257 ( .A1(n11), .A2(n53), .ZN(n284) );
  NAND2_X1 U258 ( .A1(n50), .A2(n53), .ZN(n285) );
  NAND3_X1 U259 ( .A1(n283), .A2(n284), .A3(n285), .ZN(n10) );
  XOR2_X1 U260 ( .A(n33), .B(n28), .Z(n286) );
  XOR2_X1 U261 ( .A(n246), .B(n286), .Z(product[9]) );
  NAND2_X1 U262 ( .A1(n245), .A2(n33), .ZN(n287) );
  NAND2_X1 U263 ( .A1(n7), .A2(n28), .ZN(n288) );
  NAND2_X1 U264 ( .A1(n33), .A2(n28), .ZN(n289) );
  NAND3_X1 U265 ( .A1(n287), .A2(n288), .A3(n289), .ZN(n6) );
  XOR2_X1 U266 ( .A(n95), .B(n102), .Z(n56) );
  XOR2_X1 U267 ( .A(n27), .B(n24), .Z(n290) );
  XOR2_X1 U268 ( .A(n243), .B(n290), .Z(product[10]) );
  NAND2_X1 U269 ( .A1(n281), .A2(n27), .ZN(n291) );
  NAND2_X1 U270 ( .A1(n6), .A2(n24), .ZN(n292) );
  NAND2_X1 U271 ( .A1(n27), .A2(n24), .ZN(n293) );
  NAND3_X1 U272 ( .A1(n292), .A2(n291), .A3(n293), .ZN(n5) );
  XNOR2_X1 U273 ( .A(n269), .B(n294), .ZN(product[14]) );
  XNOR2_X1 U274 ( .A(n306), .B(n15), .ZN(n294) );
  XNOR2_X2 U275 ( .A(a[4]), .B(a[3]), .ZN(n332) );
  AND3_X1 U276 ( .A1(n297), .A2(n296), .A3(n298), .ZN(product[15]) );
  INV_X1 U277 ( .A(n330), .ZN(n312) );
  OAI22_X1 U278 ( .A1(n351), .A2(n345), .B1(n343), .B2(n353), .ZN(n15) );
  INV_X1 U279 ( .A(n341), .ZN(n309) );
  INV_X1 U280 ( .A(n21), .ZN(n308) );
  INV_X1 U281 ( .A(n321), .ZN(n314) );
  INV_X1 U282 ( .A(n31), .ZN(n311) );
  INV_X1 U283 ( .A(b[0]), .ZN(n304) );
  INV_X1 U284 ( .A(a[0]), .ZN(n316) );
  INV_X1 U285 ( .A(a[3]), .ZN(n313) );
  INV_X1 U286 ( .A(a[5]), .ZN(n310) );
  INV_X1 U287 ( .A(a[7]), .ZN(n307) );
  NAND2_X1 U288 ( .A1(n254), .A2(n306), .ZN(n296) );
  NAND2_X1 U289 ( .A1(n254), .A2(n15), .ZN(n297) );
  NAND2_X1 U290 ( .A1(n306), .A2(n15), .ZN(n298) );
  XOR2_X1 U291 ( .A(n19), .B(n18), .Z(n299) );
  XOR2_X1 U292 ( .A(n266), .B(n299), .Z(product[12]) );
  NAND2_X1 U293 ( .A1(n265), .A2(n19), .ZN(n300) );
  NAND2_X1 U294 ( .A1(n4), .A2(n18), .ZN(n301) );
  NAND2_X1 U295 ( .A1(n19), .A2(n18), .ZN(n302) );
  NAND3_X1 U296 ( .A1(n264), .A2(n207), .A3(n302), .ZN(n3) );
  INV_X1 U297 ( .A(n352), .ZN(n306) );
  INV_X1 U298 ( .A(a[1]), .ZN(n315) );
  NAND2_X2 U299 ( .A1(n360), .A2(n322), .ZN(n324) );
  XOR2_X2 U300 ( .A(a[6]), .B(n310), .Z(n343) );
  NOR2_X1 U301 ( .A1(n316), .A2(n304), .ZN(product[0]) );
  OAI22_X1 U302 ( .A1(n317), .A2(n318), .B1(n319), .B2(n316), .ZN(n99) );
  OAI22_X1 U303 ( .A1(n319), .A2(n318), .B1(n320), .B2(n316), .ZN(n98) );
  XNOR2_X1 U304 ( .A(b[6]), .B(n211), .ZN(n319) );
  OAI22_X1 U305 ( .A1(n316), .A2(n320), .B1(n318), .B2(n320), .ZN(n321) );
  XNOR2_X1 U306 ( .A(b[7]), .B(n211), .ZN(n320) );
  NOR2_X1 U307 ( .A1(n221), .A2(n304), .ZN(n96) );
  OAI22_X1 U308 ( .A1(n323), .A2(n324), .B1(n221), .B2(n325), .ZN(n95) );
  XNOR2_X1 U309 ( .A(a[3]), .B(n303), .ZN(n323) );
  OAI22_X1 U310 ( .A1(n325), .A2(n324), .B1(n221), .B2(n326), .ZN(n94) );
  XNOR2_X1 U311 ( .A(b[1]), .B(a[3]), .ZN(n325) );
  OAI22_X1 U312 ( .A1(n326), .A2(n324), .B1(n221), .B2(n327), .ZN(n93) );
  XNOR2_X1 U313 ( .A(b[2]), .B(a[3]), .ZN(n326) );
  OAI22_X1 U314 ( .A1(n327), .A2(n324), .B1(n221), .B2(n328), .ZN(n92) );
  XNOR2_X1 U315 ( .A(b[3]), .B(a[3]), .ZN(n327) );
  OAI22_X1 U316 ( .A1(n328), .A2(n324), .B1(n221), .B2(n329), .ZN(n91) );
  XNOR2_X1 U317 ( .A(b[4]), .B(a[3]), .ZN(n328) );
  OAI22_X1 U318 ( .A1(n331), .A2(n221), .B1(n324), .B2(n331), .ZN(n330) );
  NOR2_X1 U319 ( .A1(n332), .A2(n304), .ZN(n88) );
  OAI22_X1 U320 ( .A1(n333), .A2(n334), .B1(n332), .B2(n335), .ZN(n87) );
  XNOR2_X1 U321 ( .A(a[5]), .B(n216), .ZN(n333) );
  OAI22_X1 U322 ( .A1(n335), .A2(n334), .B1(n332), .B2(n336), .ZN(n86) );
  XNOR2_X1 U323 ( .A(b[1]), .B(a[5]), .ZN(n335) );
  OAI22_X1 U324 ( .A1(n336), .A2(n334), .B1(n332), .B2(n337), .ZN(n85) );
  XNOR2_X1 U325 ( .A(b[2]), .B(a[5]), .ZN(n336) );
  OAI22_X1 U326 ( .A1(n337), .A2(n334), .B1(n332), .B2(n338), .ZN(n84) );
  XNOR2_X1 U327 ( .A(b[3]), .B(a[5]), .ZN(n337) );
  OAI22_X1 U328 ( .A1(n338), .A2(n334), .B1(n332), .B2(n339), .ZN(n83) );
  XNOR2_X1 U329 ( .A(b[4]), .B(a[5]), .ZN(n338) );
  OAI22_X1 U330 ( .A1(n339), .A2(n334), .B1(n332), .B2(n340), .ZN(n82) );
  XNOR2_X1 U331 ( .A(b[5]), .B(a[5]), .ZN(n339) );
  OAI22_X1 U332 ( .A1(n342), .A2(n332), .B1(n334), .B2(n342), .ZN(n341) );
  NOR2_X1 U333 ( .A1(n343), .A2(n304), .ZN(n80) );
  OAI22_X1 U334 ( .A1(n344), .A2(n345), .B1(n343), .B2(n346), .ZN(n79) );
  XNOR2_X1 U335 ( .A(a[7]), .B(n216), .ZN(n344) );
  OAI22_X1 U336 ( .A1(n347), .A2(n345), .B1(n343), .B2(n348), .ZN(n77) );
  OAI22_X1 U337 ( .A1(n348), .A2(n345), .B1(n343), .B2(n349), .ZN(n76) );
  XNOR2_X1 U338 ( .A(b[3]), .B(a[7]), .ZN(n348) );
  OAI22_X1 U339 ( .A1(n349), .A2(n345), .B1(n343), .B2(n350), .ZN(n75) );
  XNOR2_X1 U340 ( .A(b[4]), .B(a[7]), .ZN(n349) );
  OAI22_X1 U341 ( .A1(n350), .A2(n345), .B1(n343), .B2(n351), .ZN(n74) );
  XNOR2_X1 U342 ( .A(b[5]), .B(a[7]), .ZN(n350) );
  OAI22_X1 U343 ( .A1(n353), .A2(n343), .B1(n345), .B2(n353), .ZN(n352) );
  OAI21_X1 U344 ( .B1(n303), .B2(n315), .A(n318), .ZN(n72) );
  OAI21_X1 U345 ( .B1(n313), .B2(n324), .A(n354), .ZN(n71) );
  OR3_X1 U346 ( .A1(n221), .A2(n217), .A3(n313), .ZN(n354) );
  OAI21_X1 U347 ( .B1(n310), .B2(n334), .A(n355), .ZN(n70) );
  OR3_X1 U348 ( .A1(n332), .A2(n217), .A3(n310), .ZN(n355) );
  OAI21_X1 U349 ( .B1(n307), .B2(n345), .A(n356), .ZN(n69) );
  OR3_X1 U350 ( .A1(n343), .A2(n217), .A3(n307), .ZN(n356) );
  XNOR2_X1 U351 ( .A(n357), .B(n358), .ZN(n38) );
  OR2_X1 U352 ( .A1(n357), .A2(n358), .ZN(n37) );
  OAI22_X1 U353 ( .A1(n329), .A2(n324), .B1(n221), .B2(n359), .ZN(n358) );
  XNOR2_X1 U354 ( .A(b[5]), .B(a[3]), .ZN(n329) );
  OAI22_X1 U355 ( .A1(n346), .A2(n345), .B1(n343), .B2(n347), .ZN(n357) );
  XNOR2_X1 U356 ( .A(b[2]), .B(a[7]), .ZN(n347) );
  XNOR2_X1 U357 ( .A(b[1]), .B(a[7]), .ZN(n346) );
  OAI22_X1 U358 ( .A1(n359), .A2(n324), .B1(n221), .B2(n331), .ZN(n31) );
  XNOR2_X1 U359 ( .A(b[7]), .B(a[3]), .ZN(n331) );
  XNOR2_X1 U360 ( .A(n313), .B(a[2]), .ZN(n360) );
  XNOR2_X1 U361 ( .A(b[6]), .B(a[3]), .ZN(n359) );
  OAI22_X1 U362 ( .A1(n340), .A2(n334), .B1(n332), .B2(n342), .ZN(n21) );
  XNOR2_X1 U363 ( .A(b[7]), .B(a[5]), .ZN(n342) );
  XNOR2_X1 U364 ( .A(n310), .B(a[4]), .ZN(n361) );
  XNOR2_X1 U365 ( .A(b[6]), .B(a[5]), .ZN(n340) );
  XNOR2_X1 U366 ( .A(b[7]), .B(a[7]), .ZN(n353) );
  NAND2_X1 U367 ( .A1(n343), .A2(n362), .ZN(n345) );
  XNOR2_X1 U368 ( .A(n307), .B(a[6]), .ZN(n362) );
  XNOR2_X1 U369 ( .A(b[6]), .B(a[7]), .ZN(n351) );
  OAI22_X1 U370 ( .A1(n217), .A2(n318), .B1(n363), .B2(n316), .ZN(n104) );
  OAI22_X1 U371 ( .A1(n255), .A2(n318), .B1(n364), .B2(n316), .ZN(n103) );
  XNOR2_X1 U372 ( .A(b[1]), .B(a[1]), .ZN(n363) );
  OAI22_X1 U373 ( .A1(n364), .A2(n318), .B1(n365), .B2(n316), .ZN(n102) );
  XNOR2_X1 U374 ( .A(b[2]), .B(a[1]), .ZN(n364) );
  OAI22_X1 U375 ( .A1(n365), .A2(n318), .B1(n366), .B2(n316), .ZN(n101) );
  XNOR2_X1 U376 ( .A(b[3]), .B(a[1]), .ZN(n365) );
  OAI22_X1 U377 ( .A1(n366), .A2(n318), .B1(n317), .B2(n316), .ZN(n100) );
  XNOR2_X1 U378 ( .A(b[5]), .B(n211), .ZN(n317) );
  NAND2_X1 U379 ( .A1(a[1]), .A2(n316), .ZN(n318) );
  XNOR2_X1 U380 ( .A(b[4]), .B(a[1]), .ZN(n366) );
endmodule


module mac_21 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   n6, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, n2, n4;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(n6), .QN(n2) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_21_DW01_add_0 add_356 ( .A(pipeline), .B({mac_out[15:1], n6}), .CI(1'b0), 
        .SUM(sum) );
  mac_21_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n4), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n4), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n4), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n4), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n4), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n4), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n4), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n4), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n4), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n4), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n4), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n4), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n4), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n4), .ZN(N6) );
  INV_X1 U18 ( .A(n2), .ZN(mac_out[0]) );
  AND2_X1 U19 ( .A1(sum[0]), .A2(n4), .ZN(N3) );
  AND2_X1 U20 ( .A1(sum[15]), .A2(n4), .ZN(N18) );
  INV_X1 U21 ( .A(clear_acc), .ZN(n4) );
endmodule


module mac_20_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73;
  wire   [15:1] carry;

  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n73) );
  XOR2_X1 U2 ( .A(B[15]), .B(A[15]), .Z(n1) );
  XOR2_X1 U3 ( .A(carry[15]), .B(n1), .Z(SUM[15]) );
  XOR2_X1 U4 ( .A(B[4]), .B(A[4]), .Z(n2) );
  XOR2_X1 U5 ( .A(carry[4]), .B(n2), .Z(SUM[4]) );
  NAND2_X1 U6 ( .A1(carry[4]), .A2(B[4]), .ZN(n3) );
  NAND2_X1 U7 ( .A1(carry[4]), .A2(A[4]), .ZN(n4) );
  NAND2_X1 U8 ( .A1(B[4]), .A2(A[4]), .ZN(n5) );
  NAND3_X1 U9 ( .A1(n3), .A2(n4), .A3(n5), .ZN(carry[5]) );
  NAND2_X1 U10 ( .A1(n32), .A2(B[13]), .ZN(n6) );
  NAND3_X1 U11 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n7) );
  NAND3_X1 U12 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n8) );
  NAND3_X1 U13 ( .A1(n12), .A2(n13), .A3(n14), .ZN(n9) );
  NAND3_X1 U14 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n10) );
  XOR2_X1 U15 ( .A(B[10]), .B(A[10]), .Z(n11) );
  XOR2_X1 U16 ( .A(n7), .B(n11), .Z(SUM[10]) );
  NAND2_X1 U17 ( .A1(n7), .A2(B[10]), .ZN(n12) );
  NAND2_X1 U18 ( .A1(carry[10]), .A2(A[10]), .ZN(n13) );
  NAND2_X1 U19 ( .A1(B[10]), .A2(A[10]), .ZN(n14) );
  NAND3_X1 U20 ( .A1(n12), .A2(n13), .A3(n14), .ZN(carry[11]) );
  NAND3_X1 U21 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n15) );
  NAND3_X1 U22 ( .A1(n70), .A2(n71), .A3(n72), .ZN(n16) );
  NAND3_X1 U23 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n17) );
  NAND3_X1 U24 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n18) );
  XOR2_X1 U25 ( .A(B[3]), .B(A[3]), .Z(n19) );
  XOR2_X1 U26 ( .A(n16), .B(n19), .Z(SUM[3]) );
  NAND2_X1 U27 ( .A1(n16), .A2(B[3]), .ZN(n20) );
  NAND2_X1 U28 ( .A1(carry[3]), .A2(A[3]), .ZN(n21) );
  NAND2_X1 U29 ( .A1(B[3]), .A2(A[3]), .ZN(n22) );
  NAND3_X1 U30 ( .A1(n20), .A2(n21), .A3(n22), .ZN(carry[4]) );
  NAND3_X1 U31 ( .A1(n6), .A2(n45), .A3(n46), .ZN(n23) );
  XOR2_X1 U32 ( .A(B[11]), .B(A[11]), .Z(n24) );
  XOR2_X1 U33 ( .A(n9), .B(n24), .Z(SUM[11]) );
  NAND2_X1 U34 ( .A1(n9), .A2(B[11]), .ZN(n25) );
  NAND2_X1 U35 ( .A1(carry[11]), .A2(A[11]), .ZN(n26) );
  NAND2_X1 U36 ( .A1(B[11]), .A2(A[11]), .ZN(n27) );
  NAND3_X1 U37 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[12]) );
  XOR2_X1 U38 ( .A(B[5]), .B(A[5]), .Z(n28) );
  XOR2_X1 U39 ( .A(carry[5]), .B(n28), .Z(SUM[5]) );
  NAND2_X1 U40 ( .A1(carry[5]), .A2(B[5]), .ZN(n29) );
  NAND2_X1 U41 ( .A1(carry[5]), .A2(A[5]), .ZN(n30) );
  NAND2_X1 U42 ( .A1(B[5]), .A2(A[5]), .ZN(n31) );
  NAND3_X1 U43 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[6]) );
  NAND3_X1 U44 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n32) );
  XOR2_X1 U45 ( .A(B[12]), .B(A[12]), .Z(n33) );
  XOR2_X1 U46 ( .A(n8), .B(n33), .Z(SUM[12]) );
  NAND2_X1 U47 ( .A1(n8), .A2(B[12]), .ZN(n34) );
  NAND2_X1 U48 ( .A1(carry[12]), .A2(A[12]), .ZN(n35) );
  NAND2_X1 U49 ( .A1(B[12]), .A2(A[12]), .ZN(n36) );
  NAND3_X1 U50 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[13]) );
  XOR2_X1 U51 ( .A(B[6]), .B(A[6]), .Z(n37) );
  XOR2_X1 U52 ( .A(n18), .B(n37), .Z(SUM[6]) );
  NAND2_X1 U53 ( .A1(n17), .A2(B[6]), .ZN(n38) );
  NAND2_X1 U54 ( .A1(carry[6]), .A2(A[6]), .ZN(n39) );
  NAND2_X1 U55 ( .A1(B[6]), .A2(A[6]), .ZN(n40) );
  NAND3_X1 U56 ( .A1(n39), .A2(n38), .A3(n40), .ZN(carry[7]) );
  NAND3_X1 U57 ( .A1(n6), .A2(n45), .A3(n46), .ZN(n41) );
  NAND3_X1 U58 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n42) );
  XOR2_X1 U59 ( .A(B[13]), .B(A[13]), .Z(n43) );
  XOR2_X1 U60 ( .A(n32), .B(n43), .Z(SUM[13]) );
  NAND2_X1 U61 ( .A1(n32), .A2(B[13]), .ZN(n44) );
  NAND2_X1 U62 ( .A1(carry[13]), .A2(A[13]), .ZN(n45) );
  NAND2_X1 U63 ( .A1(B[13]), .A2(A[13]), .ZN(n46) );
  NAND3_X1 U64 ( .A1(n44), .A2(n45), .A3(n46), .ZN(carry[14]) );
  XOR2_X1 U65 ( .A(B[7]), .B(A[7]), .Z(n47) );
  XOR2_X1 U66 ( .A(n15), .B(n47), .Z(SUM[7]) );
  NAND2_X1 U67 ( .A1(n15), .A2(B[7]), .ZN(n48) );
  NAND2_X1 U68 ( .A1(carry[7]), .A2(A[7]), .ZN(n49) );
  NAND2_X1 U69 ( .A1(B[7]), .A2(A[7]), .ZN(n50) );
  NAND3_X1 U70 ( .A1(n48), .A2(n49), .A3(n50), .ZN(carry[8]) );
  NAND3_X1 U71 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n51) );
  NAND3_X1 U72 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n52) );
  XOR2_X1 U73 ( .A(B[14]), .B(A[14]), .Z(n53) );
  XOR2_X1 U74 ( .A(n23), .B(n53), .Z(SUM[14]) );
  NAND2_X1 U75 ( .A1(n41), .A2(B[14]), .ZN(n54) );
  NAND2_X1 U76 ( .A1(carry[14]), .A2(A[14]), .ZN(n55) );
  NAND2_X1 U77 ( .A1(B[14]), .A2(A[14]), .ZN(n56) );
  NAND3_X1 U78 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[15]) );
  XOR2_X1 U79 ( .A(B[8]), .B(A[8]), .Z(n57) );
  XOR2_X1 U80 ( .A(n42), .B(n57), .Z(SUM[8]) );
  NAND2_X1 U81 ( .A1(n42), .A2(B[8]), .ZN(n58) );
  NAND2_X1 U82 ( .A1(carry[8]), .A2(A[8]), .ZN(n59) );
  NAND2_X1 U83 ( .A1(B[8]), .A2(A[8]), .ZN(n60) );
  NAND3_X1 U84 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[9]) );
  XOR2_X1 U85 ( .A(B[9]), .B(A[9]), .Z(n61) );
  XOR2_X1 U86 ( .A(n10), .B(n61), .Z(SUM[9]) );
  NAND2_X1 U87 ( .A1(n10), .A2(B[9]), .ZN(n62) );
  NAND2_X1 U88 ( .A1(carry[9]), .A2(A[9]), .ZN(n63) );
  NAND2_X1 U89 ( .A1(B[9]), .A2(A[9]), .ZN(n64) );
  NAND3_X1 U90 ( .A1(n62), .A2(n63), .A3(n64), .ZN(carry[10]) );
  XOR2_X1 U91 ( .A(B[1]), .B(A[1]), .Z(n65) );
  XOR2_X1 U92 ( .A(n73), .B(n65), .Z(SUM[1]) );
  NAND2_X1 U93 ( .A1(n73), .A2(B[1]), .ZN(n66) );
  NAND2_X1 U94 ( .A1(n73), .A2(A[1]), .ZN(n67) );
  NAND2_X1 U95 ( .A1(B[1]), .A2(A[1]), .ZN(n68) );
  NAND3_X1 U96 ( .A1(n66), .A2(n67), .A3(n68), .ZN(carry[2]) );
  XOR2_X1 U97 ( .A(B[2]), .B(A[2]), .Z(n69) );
  XOR2_X1 U98 ( .A(n52), .B(n69), .Z(SUM[2]) );
  NAND2_X1 U99 ( .A1(n51), .A2(B[2]), .ZN(n70) );
  NAND2_X1 U100 ( .A1(carry[2]), .A2(A[2]), .ZN(n71) );
  NAND2_X1 U101 ( .A1(B[2]), .A2(A[2]), .ZN(n72) );
  NAND3_X1 U102 ( .A1(n70), .A2(n71), .A3(n72), .ZN(carry[3]) );
  XOR2_X1 U103 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_20_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n306), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n305), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n309), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n308), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n310), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  BUF_X1 U157 ( .A(n301), .Z(n256) );
  CLKBUF_X1 U158 ( .A(n212), .Z(n206) );
  BUF_X2 U159 ( .A(a[1]), .Z(n216) );
  XOR2_X1 U160 ( .A(n301), .B(a[3]), .Z(n319) );
  NAND3_X1 U161 ( .A1(n269), .A2(n268), .A3(n270), .ZN(n207) );
  INV_X1 U162 ( .A(n301), .ZN(n300) );
  AND2_X1 U163 ( .A1(n104), .A2(n72), .ZN(n208) );
  AND2_X1 U164 ( .A1(n104), .A2(n72), .ZN(n209) );
  CLKBUF_X1 U165 ( .A(a[3]), .Z(n210) );
  AND2_X1 U166 ( .A1(n228), .A2(n102), .ZN(n211) );
  NAND2_X1 U167 ( .A1(n215), .A2(n34), .ZN(n212) );
  CLKBUF_X1 U168 ( .A(n227), .Z(n213) );
  NAND2_X2 U169 ( .A1(n235), .A2(n236), .ZN(n214) );
  NAND2_X1 U170 ( .A1(n235), .A2(n236), .ZN(n328) );
  NAND3_X1 U171 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n215) );
  CLKBUF_X1 U172 ( .A(b[1]), .Z(n217) );
  CLKBUF_X1 U173 ( .A(n3), .Z(n218) );
  NAND3_X1 U174 ( .A1(n239), .A2(n238), .A3(n240), .ZN(n219) );
  NAND3_X1 U175 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n220) );
  NAND3_X1 U176 ( .A1(n212), .A2(n250), .A3(n251), .ZN(n221) );
  NAND3_X1 U177 ( .A1(n206), .A2(n250), .A3(n251), .ZN(n222) );
  XOR2_X2 U178 ( .A(a[6]), .B(n307), .Z(n339) );
  NAND3_X1 U179 ( .A1(n277), .A2(n276), .A3(n278), .ZN(n223) );
  NAND3_X1 U180 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n224) );
  NAND3_X1 U181 ( .A1(n285), .A2(n286), .A3(n287), .ZN(n225) );
  NAND3_X1 U182 ( .A1(n285), .A2(n286), .A3(n287), .ZN(n226) );
  NAND3_X1 U183 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n227) );
  XOR2_X1 U184 ( .A(n102), .B(n95), .Z(n56) );
  OAI22_X1 U185 ( .A1(n319), .A2(n320), .B1(n290), .B2(n321), .ZN(n228) );
  CLKBUF_X1 U186 ( .A(n265), .Z(n229) );
  CLKBUF_X1 U187 ( .A(n6), .Z(n230) );
  CLKBUF_X1 U188 ( .A(n223), .Z(n231) );
  NAND3_X1 U189 ( .A1(n298), .A2(n297), .A3(n299), .ZN(n232) );
  NAND2_X1 U190 ( .A1(a[4]), .A2(a[3]), .ZN(n235) );
  NAND2_X1 U191 ( .A1(n233), .A2(n234), .ZN(n236) );
  INV_X1 U192 ( .A(a[4]), .ZN(n233) );
  INV_X1 U193 ( .A(a[3]), .ZN(n234) );
  XOR2_X1 U194 ( .A(n33), .B(n28), .Z(n237) );
  XOR2_X1 U195 ( .A(n222), .B(n237), .Z(product[9]) );
  NAND2_X1 U196 ( .A1(n221), .A2(n33), .ZN(n238) );
  NAND2_X1 U197 ( .A1(n7), .A2(n28), .ZN(n239) );
  NAND2_X1 U198 ( .A1(n33), .A2(n28), .ZN(n240) );
  NAND3_X1 U199 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n6) );
  XOR2_X1 U200 ( .A(n103), .B(n96), .Z(n241) );
  XOR2_X1 U201 ( .A(n14), .B(n241), .Z(product[2]) );
  NAND2_X1 U202 ( .A1(n209), .A2(n103), .ZN(n242) );
  NAND2_X1 U203 ( .A1(n208), .A2(n96), .ZN(n243) );
  NAND2_X1 U204 ( .A1(n103), .A2(n96), .ZN(n244) );
  NAND3_X1 U205 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n13) );
  CLKBUF_X1 U206 ( .A(n215), .Z(n245) );
  NAND3_X1 U207 ( .A1(n269), .A2(n268), .A3(n270), .ZN(n246) );
  NAND3_X1 U208 ( .A1(n269), .A2(n268), .A3(n270), .ZN(n247) );
  XOR2_X1 U209 ( .A(n34), .B(n39), .Z(n248) );
  XOR2_X1 U210 ( .A(n245), .B(n248), .Z(product[8]) );
  NAND2_X1 U211 ( .A1(n215), .A2(n34), .ZN(n249) );
  NAND2_X1 U212 ( .A1(n8), .A2(n39), .ZN(n250) );
  NAND2_X1 U213 ( .A1(n34), .A2(n39), .ZN(n251) );
  NAND3_X1 U214 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n7) );
  XOR2_X1 U215 ( .A(n46), .B(n49), .Z(n252) );
  XOR2_X1 U216 ( .A(n226), .B(n252), .Z(product[6]) );
  NAND2_X1 U217 ( .A1(n225), .A2(n46), .ZN(n253) );
  NAND2_X1 U218 ( .A1(n10), .A2(n49), .ZN(n254) );
  NAND2_X1 U219 ( .A1(n46), .A2(n49), .ZN(n255) );
  NAND3_X1 U220 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n9) );
  XOR2_X1 U221 ( .A(n40), .B(n45), .Z(n257) );
  XOR2_X1 U222 ( .A(n213), .B(n257), .Z(product[7]) );
  NAND2_X1 U223 ( .A1(n227), .A2(n40), .ZN(n258) );
  NAND2_X1 U224 ( .A1(n9), .A2(n45), .ZN(n259) );
  NAND2_X1 U225 ( .A1(n40), .A2(n45), .ZN(n260) );
  NAND3_X1 U226 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n8) );
  XOR2_X1 U227 ( .A(n20), .B(n23), .Z(n261) );
  XOR2_X1 U228 ( .A(n231), .B(n261), .Z(product[11]) );
  NAND2_X1 U229 ( .A1(n223), .A2(n20), .ZN(n262) );
  NAND2_X1 U230 ( .A1(n5), .A2(n23), .ZN(n263) );
  NAND2_X1 U231 ( .A1(n20), .A2(n23), .ZN(n264) );
  NAND3_X1 U232 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n4) );
  NAND3_X1 U233 ( .A1(n272), .A2(n274), .A3(n273), .ZN(n265) );
  NAND3_X1 U234 ( .A1(n281), .A2(n282), .A3(n283), .ZN(n266) );
  XOR2_X1 U235 ( .A(n302), .B(n17), .Z(n267) );
  XOR2_X1 U236 ( .A(n218), .B(n267), .Z(product[13]) );
  NAND2_X1 U237 ( .A1(n232), .A2(n302), .ZN(n268) );
  NAND2_X1 U238 ( .A1(n3), .A2(n17), .ZN(n269) );
  NAND2_X1 U239 ( .A1(n302), .A2(n17), .ZN(n270) );
  XOR2_X1 U240 ( .A(n56), .B(n71), .Z(n271) );
  XOR2_X1 U241 ( .A(n220), .B(n271), .Z(product[3]) );
  NAND2_X1 U242 ( .A1(n220), .A2(n56), .ZN(n272) );
  NAND2_X1 U243 ( .A1(n13), .A2(n71), .ZN(n273) );
  NAND2_X1 U244 ( .A1(n56), .A2(n71), .ZN(n274) );
  NAND3_X1 U245 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n12) );
  XOR2_X1 U246 ( .A(n27), .B(n24), .Z(n275) );
  XOR2_X1 U247 ( .A(n230), .B(n275), .Z(product[10]) );
  NAND2_X1 U248 ( .A1(n6), .A2(n27), .ZN(n276) );
  NAND2_X1 U249 ( .A1(n219), .A2(n24), .ZN(n277) );
  NAND2_X1 U250 ( .A1(n27), .A2(n24), .ZN(n278) );
  NAND3_X1 U251 ( .A1(n277), .A2(n276), .A3(n278), .ZN(n5) );
  CLKBUF_X1 U252 ( .A(n266), .Z(n279) );
  XOR2_X1 U253 ( .A(n54), .B(n211), .Z(n280) );
  XOR2_X1 U254 ( .A(n229), .B(n280), .Z(product[4]) );
  NAND2_X1 U255 ( .A1(n265), .A2(n54), .ZN(n281) );
  NAND2_X1 U256 ( .A1(n12), .A2(n211), .ZN(n282) );
  NAND2_X1 U257 ( .A1(n54), .A2(n211), .ZN(n283) );
  NAND3_X1 U258 ( .A1(n281), .A2(n282), .A3(n283), .ZN(n11) );
  XOR2_X1 U259 ( .A(n50), .B(n53), .Z(n284) );
  XOR2_X1 U260 ( .A(n279), .B(n284), .Z(product[5]) );
  NAND2_X1 U261 ( .A1(n266), .A2(n50), .ZN(n285) );
  NAND2_X1 U262 ( .A1(n11), .A2(n53), .ZN(n286) );
  NAND2_X1 U263 ( .A1(n50), .A2(n53), .ZN(n287) );
  NAND3_X1 U264 ( .A1(n285), .A2(n286), .A3(n287), .ZN(n10) );
  XNOR2_X1 U265 ( .A(n217), .B(n216), .ZN(n288) );
  NAND2_X2 U266 ( .A1(n318), .A2(n356), .ZN(n320) );
  NAND2_X2 U267 ( .A1(n328), .A2(n357), .ZN(n330) );
  XOR2_X1 U268 ( .A(a[2]), .B(n311), .Z(n289) );
  XOR2_X1 U269 ( .A(a[2]), .B(n311), .Z(n290) );
  INV_X1 U270 ( .A(n15), .ZN(n302) );
  XNOR2_X1 U271 ( .A(n224), .B(n291), .ZN(product[12]) );
  XNOR2_X1 U272 ( .A(n19), .B(n18), .ZN(n291) );
  XNOR2_X1 U273 ( .A(n247), .B(n292), .ZN(product[14]) );
  XNOR2_X1 U274 ( .A(n303), .B(n15), .ZN(n292) );
  AND3_X1 U275 ( .A1(n295), .A2(n294), .A3(n296), .ZN(product[15]) );
  OAI22_X1 U276 ( .A1(n347), .A2(n341), .B1(n339), .B2(n349), .ZN(n15) );
  INV_X1 U277 ( .A(n337), .ZN(n306) );
  INV_X1 U278 ( .A(n21), .ZN(n305) );
  INV_X1 U279 ( .A(n317), .ZN(n310) );
  INV_X1 U280 ( .A(n326), .ZN(n309) );
  INV_X1 U281 ( .A(n31), .ZN(n308) );
  INV_X1 U282 ( .A(b[0]), .ZN(n301) );
  XOR2_X1 U283 ( .A(a[2]), .B(n311), .Z(n318) );
  INV_X1 U284 ( .A(a[0]), .ZN(n312) );
  INV_X1 U285 ( .A(a[5]), .ZN(n307) );
  INV_X1 U286 ( .A(a[7]), .ZN(n304) );
  NAND2_X1 U287 ( .A1(n246), .A2(n303), .ZN(n294) );
  NAND2_X1 U288 ( .A1(n207), .A2(n15), .ZN(n295) );
  NAND2_X1 U289 ( .A1(n303), .A2(n15), .ZN(n296) );
  NAND2_X1 U290 ( .A1(n4), .A2(n19), .ZN(n297) );
  NAND2_X1 U291 ( .A1(n224), .A2(n18), .ZN(n298) );
  NAND2_X1 U292 ( .A1(n19), .A2(n18), .ZN(n299) );
  NAND3_X1 U293 ( .A1(n298), .A2(n297), .A3(n299), .ZN(n3) );
  INV_X1 U294 ( .A(n348), .ZN(n303) );
  INV_X1 U295 ( .A(a[1]), .ZN(n311) );
  NOR2_X1 U296 ( .A1(n312), .A2(n256), .ZN(product[0]) );
  OAI22_X1 U297 ( .A1(n313), .A2(n314), .B1(n315), .B2(n312), .ZN(n99) );
  OAI22_X1 U298 ( .A1(n315), .A2(n314), .B1(n316), .B2(n312), .ZN(n98) );
  XNOR2_X1 U299 ( .A(b[6]), .B(n216), .ZN(n315) );
  OAI22_X1 U300 ( .A1(n312), .A2(n316), .B1(n314), .B2(n316), .ZN(n317) );
  XNOR2_X1 U301 ( .A(b[7]), .B(n216), .ZN(n316) );
  NOR2_X1 U302 ( .A1(n289), .A2(n256), .ZN(n96) );
  OAI22_X1 U303 ( .A1(n319), .A2(n320), .B1(n290), .B2(n321), .ZN(n95) );
  OAI22_X1 U304 ( .A1(n321), .A2(n320), .B1(n290), .B2(n322), .ZN(n94) );
  XNOR2_X1 U305 ( .A(b[1]), .B(a[3]), .ZN(n321) );
  OAI22_X1 U306 ( .A1(n322), .A2(n320), .B1(n289), .B2(n323), .ZN(n93) );
  XNOR2_X1 U307 ( .A(b[2]), .B(a[3]), .ZN(n322) );
  OAI22_X1 U308 ( .A1(n323), .A2(n320), .B1(n290), .B2(n324), .ZN(n92) );
  XNOR2_X1 U309 ( .A(b[3]), .B(n210), .ZN(n323) );
  OAI22_X1 U310 ( .A1(n324), .A2(n320), .B1(n290), .B2(n325), .ZN(n91) );
  XNOR2_X1 U311 ( .A(b[4]), .B(a[3]), .ZN(n324) );
  OAI22_X1 U312 ( .A1(n327), .A2(n289), .B1(n320), .B2(n327), .ZN(n326) );
  NOR2_X1 U313 ( .A1(n214), .A2(n256), .ZN(n88) );
  OAI22_X1 U314 ( .A1(n329), .A2(n330), .B1(n214), .B2(n331), .ZN(n87) );
  XNOR2_X1 U315 ( .A(a[5]), .B(n300), .ZN(n329) );
  OAI22_X1 U316 ( .A1(n331), .A2(n330), .B1(n214), .B2(n332), .ZN(n86) );
  XNOR2_X1 U317 ( .A(b[1]), .B(a[5]), .ZN(n331) );
  OAI22_X1 U318 ( .A1(n332), .A2(n330), .B1(n214), .B2(n333), .ZN(n85) );
  XNOR2_X1 U319 ( .A(b[2]), .B(a[5]), .ZN(n332) );
  OAI22_X1 U320 ( .A1(n333), .A2(n330), .B1(n214), .B2(n334), .ZN(n84) );
  XNOR2_X1 U321 ( .A(b[3]), .B(a[5]), .ZN(n333) );
  OAI22_X1 U322 ( .A1(n334), .A2(n330), .B1(n214), .B2(n335), .ZN(n83) );
  XNOR2_X1 U323 ( .A(b[4]), .B(a[5]), .ZN(n334) );
  OAI22_X1 U324 ( .A1(n335), .A2(n330), .B1(n214), .B2(n336), .ZN(n82) );
  XNOR2_X1 U325 ( .A(b[5]), .B(a[5]), .ZN(n335) );
  OAI22_X1 U326 ( .A1(n338), .A2(n214), .B1(n330), .B2(n338), .ZN(n337) );
  NOR2_X1 U327 ( .A1(n339), .A2(n256), .ZN(n80) );
  OAI22_X1 U328 ( .A1(n340), .A2(n341), .B1(n339), .B2(n342), .ZN(n79) );
  XNOR2_X1 U329 ( .A(a[7]), .B(n300), .ZN(n340) );
  OAI22_X1 U330 ( .A1(n343), .A2(n341), .B1(n339), .B2(n344), .ZN(n77) );
  OAI22_X1 U331 ( .A1(n344), .A2(n341), .B1(n339), .B2(n345), .ZN(n76) );
  XNOR2_X1 U332 ( .A(b[3]), .B(a[7]), .ZN(n344) );
  OAI22_X1 U333 ( .A1(n345), .A2(n341), .B1(n339), .B2(n346), .ZN(n75) );
  XNOR2_X1 U334 ( .A(b[4]), .B(a[7]), .ZN(n345) );
  OAI22_X1 U335 ( .A1(n346), .A2(n341), .B1(n339), .B2(n347), .ZN(n74) );
  XNOR2_X1 U336 ( .A(b[5]), .B(a[7]), .ZN(n346) );
  OAI22_X1 U337 ( .A1(n349), .A2(n339), .B1(n341), .B2(n349), .ZN(n348) );
  OAI21_X1 U338 ( .B1(n300), .B2(n311), .A(n314), .ZN(n72) );
  OAI21_X1 U339 ( .B1(n234), .B2(n320), .A(n350), .ZN(n71) );
  OR3_X1 U340 ( .A1(n289), .A2(n300), .A3(n234), .ZN(n350) );
  OAI21_X1 U341 ( .B1(n307), .B2(n330), .A(n351), .ZN(n70) );
  OR3_X1 U342 ( .A1(n328), .A2(n300), .A3(n307), .ZN(n351) );
  OAI21_X1 U343 ( .B1(n304), .B2(n341), .A(n352), .ZN(n69) );
  OR3_X1 U344 ( .A1(n339), .A2(n300), .A3(n304), .ZN(n352) );
  XNOR2_X1 U345 ( .A(n353), .B(n354), .ZN(n38) );
  OR2_X1 U346 ( .A1(n353), .A2(n354), .ZN(n37) );
  OAI22_X1 U347 ( .A1(n325), .A2(n320), .B1(n289), .B2(n355), .ZN(n354) );
  XNOR2_X1 U348 ( .A(b[5]), .B(n210), .ZN(n325) );
  OAI22_X1 U349 ( .A1(n342), .A2(n341), .B1(n339), .B2(n343), .ZN(n353) );
  XNOR2_X1 U350 ( .A(b[2]), .B(a[7]), .ZN(n343) );
  XNOR2_X1 U351 ( .A(n217), .B(a[7]), .ZN(n342) );
  OAI22_X1 U352 ( .A1(n355), .A2(n320), .B1(n290), .B2(n327), .ZN(n31) );
  XNOR2_X1 U353 ( .A(b[7]), .B(n210), .ZN(n327) );
  XNOR2_X1 U354 ( .A(n234), .B(a[2]), .ZN(n356) );
  XNOR2_X1 U355 ( .A(b[6]), .B(n210), .ZN(n355) );
  OAI22_X1 U356 ( .A1(n336), .A2(n330), .B1(n214), .B2(n338), .ZN(n21) );
  XNOR2_X1 U357 ( .A(b[7]), .B(a[5]), .ZN(n338) );
  XNOR2_X1 U358 ( .A(n307), .B(a[4]), .ZN(n357) );
  XNOR2_X1 U359 ( .A(b[6]), .B(a[5]), .ZN(n336) );
  XNOR2_X1 U360 ( .A(b[7]), .B(a[7]), .ZN(n349) );
  NAND2_X1 U361 ( .A1(n339), .A2(n358), .ZN(n341) );
  XNOR2_X1 U362 ( .A(n304), .B(a[6]), .ZN(n358) );
  XNOR2_X1 U363 ( .A(b[6]), .B(a[7]), .ZN(n347) );
  OAI22_X1 U364 ( .A1(n300), .A2(n314), .B1(n359), .B2(n312), .ZN(n104) );
  OAI22_X1 U365 ( .A1(n288), .A2(n314), .B1(n360), .B2(n312), .ZN(n103) );
  XNOR2_X1 U366 ( .A(b[1]), .B(a[1]), .ZN(n359) );
  OAI22_X1 U367 ( .A1(n360), .A2(n314), .B1(n361), .B2(n312), .ZN(n102) );
  XNOR2_X1 U368 ( .A(b[2]), .B(a[1]), .ZN(n360) );
  OAI22_X1 U369 ( .A1(n361), .A2(n314), .B1(n362), .B2(n312), .ZN(n101) );
  XNOR2_X1 U370 ( .A(b[3]), .B(n216), .ZN(n361) );
  OAI22_X1 U371 ( .A1(n362), .A2(n314), .B1(n313), .B2(n312), .ZN(n100) );
  XNOR2_X1 U372 ( .A(b[5]), .B(n216), .ZN(n313) );
  NAND2_X1 U373 ( .A1(a[1]), .A2(n312), .ZN(n314) );
  XNOR2_X1 U374 ( .A(b[4]), .B(n216), .ZN(n362) );
endmodule


module mac_20 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  mac_20_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_20_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_19_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;
  wire   [15:1] carry;

  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n77) );
  XOR2_X1 U2 ( .A(B[15]), .B(A[15]), .Z(n1) );
  XOR2_X1 U3 ( .A(carry[15]), .B(n1), .Z(SUM[15]) );
  NAND2_X1 U4 ( .A1(carry[10]), .A2(A[10]), .ZN(n2) );
  NAND3_X1 U5 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n3) );
  NAND3_X1 U6 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n4) );
  XOR2_X1 U7 ( .A(B[2]), .B(A[2]), .Z(n5) );
  XOR2_X1 U8 ( .A(n4), .B(n5), .Z(SUM[2]) );
  NAND2_X1 U9 ( .A1(n3), .A2(B[2]), .ZN(n6) );
  NAND2_X1 U10 ( .A1(carry[2]), .A2(A[2]), .ZN(n7) );
  NAND2_X1 U11 ( .A1(B[2]), .A2(A[2]), .ZN(n8) );
  NAND3_X1 U12 ( .A1(n6), .A2(n7), .A3(n8), .ZN(carry[3]) );
  XOR2_X1 U13 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U14 ( .A(carry[3]), .B(n9), .Z(SUM[3]) );
  NAND2_X1 U15 ( .A1(carry[3]), .A2(B[3]), .ZN(n10) );
  NAND2_X1 U16 ( .A1(carry[3]), .A2(A[3]), .ZN(n11) );
  NAND2_X1 U17 ( .A1(B[3]), .A2(A[3]), .ZN(n12) );
  NAND3_X1 U18 ( .A1(n10), .A2(n11), .A3(n12), .ZN(carry[4]) );
  NAND3_X1 U19 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n13) );
  NAND2_X1 U20 ( .A1(n29), .A2(B[6]), .ZN(n14) );
  NAND3_X1 U21 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n15) );
  NAND3_X1 U22 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n16) );
  XOR2_X1 U23 ( .A(B[4]), .B(A[4]), .Z(n17) );
  XOR2_X1 U24 ( .A(carry[4]), .B(n17), .Z(SUM[4]) );
  NAND2_X1 U25 ( .A1(carry[4]), .A2(B[4]), .ZN(n18) );
  NAND2_X1 U26 ( .A1(carry[4]), .A2(A[4]), .ZN(n19) );
  NAND2_X1 U27 ( .A1(B[4]), .A2(A[4]), .ZN(n20) );
  NAND3_X1 U28 ( .A1(n18), .A2(n19), .A3(n20), .ZN(carry[5]) );
  NAND3_X1 U29 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n21) );
  NAND3_X1 U30 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n22) );
  NAND3_X1 U31 ( .A1(n26), .A2(n2), .A3(n28), .ZN(n23) );
  NAND3_X1 U32 ( .A1(n26), .A2(n2), .A3(n28), .ZN(n24) );
  XOR2_X1 U33 ( .A(B[10]), .B(A[10]), .Z(n25) );
  XOR2_X1 U34 ( .A(n22), .B(n25), .Z(SUM[10]) );
  NAND2_X1 U35 ( .A1(n21), .A2(B[10]), .ZN(n26) );
  NAND2_X1 U36 ( .A1(carry[10]), .A2(A[10]), .ZN(n27) );
  NAND2_X1 U37 ( .A1(B[10]), .A2(A[10]), .ZN(n28) );
  NAND3_X1 U38 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[11]) );
  NAND3_X1 U39 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n29) );
  NAND3_X1 U40 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n30) );
  NAND3_X1 U41 ( .A1(n74), .A2(n75), .A3(n76), .ZN(n31) );
  XOR2_X1 U42 ( .A(B[11]), .B(A[11]), .Z(n32) );
  XOR2_X1 U43 ( .A(n24), .B(n32), .Z(SUM[11]) );
  NAND2_X1 U44 ( .A1(n23), .A2(B[11]), .ZN(n33) );
  NAND2_X1 U45 ( .A1(carry[11]), .A2(A[11]), .ZN(n34) );
  NAND2_X1 U46 ( .A1(B[11]), .A2(A[11]), .ZN(n35) );
  NAND3_X1 U47 ( .A1(n34), .A2(n33), .A3(n35), .ZN(carry[12]) );
  XOR2_X1 U48 ( .A(B[5]), .B(A[5]), .Z(n36) );
  XOR2_X1 U49 ( .A(n15), .B(n36), .Z(SUM[5]) );
  NAND2_X1 U50 ( .A1(n15), .A2(B[5]), .ZN(n37) );
  NAND2_X1 U51 ( .A1(carry[5]), .A2(A[5]), .ZN(n38) );
  NAND2_X1 U52 ( .A1(B[5]), .A2(A[5]), .ZN(n39) );
  NAND3_X1 U53 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[6]) );
  NAND3_X1 U54 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n40) );
  XOR2_X1 U55 ( .A(B[12]), .B(A[12]), .Z(n41) );
  XOR2_X1 U56 ( .A(n16), .B(n41), .Z(SUM[12]) );
  NAND2_X1 U57 ( .A1(n16), .A2(B[12]), .ZN(n42) );
  NAND2_X1 U58 ( .A1(carry[12]), .A2(A[12]), .ZN(n43) );
  NAND2_X1 U59 ( .A1(B[12]), .A2(A[12]), .ZN(n44) );
  NAND3_X1 U60 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[13]) );
  NAND3_X1 U61 ( .A1(n14), .A2(n67), .A3(n68), .ZN(n45) );
  NAND3_X1 U62 ( .A1(n14), .A2(n67), .A3(n68), .ZN(n46) );
  NAND3_X1 U63 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n47) );
  XOR2_X1 U64 ( .A(B[9]), .B(A[9]), .Z(n48) );
  XOR2_X1 U65 ( .A(n47), .B(n48), .Z(SUM[9]) );
  NAND2_X1 U66 ( .A1(n47), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U67 ( .A1(carry[9]), .A2(A[9]), .ZN(n50) );
  NAND2_X1 U68 ( .A1(B[9]), .A2(A[9]), .ZN(n51) );
  NAND3_X1 U69 ( .A1(n49), .A2(n50), .A3(n51), .ZN(carry[10]) );
  NAND3_X1 U70 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n52) );
  XOR2_X1 U71 ( .A(B[8]), .B(A[8]), .Z(n53) );
  XOR2_X1 U72 ( .A(n31), .B(n53), .Z(SUM[8]) );
  NAND2_X1 U73 ( .A1(n31), .A2(B[8]), .ZN(n54) );
  NAND2_X1 U74 ( .A1(carry[8]), .A2(A[8]), .ZN(n55) );
  NAND2_X1 U75 ( .A1(B[8]), .A2(A[8]), .ZN(n56) );
  NAND3_X1 U76 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[9]) );
  XOR2_X1 U77 ( .A(B[1]), .B(A[1]), .Z(n57) );
  XOR2_X1 U78 ( .A(n77), .B(n57), .Z(SUM[1]) );
  NAND2_X1 U79 ( .A1(n77), .A2(B[1]), .ZN(n58) );
  NAND2_X1 U80 ( .A1(n77), .A2(A[1]), .ZN(n59) );
  NAND2_X1 U81 ( .A1(B[1]), .A2(A[1]), .ZN(n60) );
  NAND3_X1 U82 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[2]) );
  XOR2_X1 U83 ( .A(B[13]), .B(A[13]), .Z(n61) );
  XOR2_X1 U84 ( .A(n13), .B(n61), .Z(SUM[13]) );
  NAND2_X1 U85 ( .A1(carry[13]), .A2(B[13]), .ZN(n62) );
  NAND2_X1 U86 ( .A1(n40), .A2(A[13]), .ZN(n63) );
  NAND2_X1 U87 ( .A1(B[13]), .A2(A[13]), .ZN(n64) );
  XOR2_X1 U88 ( .A(B[6]), .B(A[6]), .Z(n65) );
  XOR2_X1 U89 ( .A(n29), .B(n65), .Z(SUM[6]) );
  NAND2_X1 U90 ( .A1(n29), .A2(B[6]), .ZN(n66) );
  NAND2_X1 U91 ( .A1(carry[6]), .A2(A[6]), .ZN(n67) );
  NAND2_X1 U92 ( .A1(B[6]), .A2(A[6]), .ZN(n68) );
  NAND3_X1 U93 ( .A1(n66), .A2(n67), .A3(n68), .ZN(carry[7]) );
  XOR2_X1 U94 ( .A(B[14]), .B(A[14]), .Z(n69) );
  XOR2_X1 U95 ( .A(n30), .B(n69), .Z(SUM[14]) );
  NAND2_X1 U96 ( .A1(n52), .A2(B[14]), .ZN(n70) );
  NAND2_X1 U97 ( .A1(n52), .A2(A[14]), .ZN(n71) );
  NAND2_X1 U98 ( .A1(B[14]), .A2(A[14]), .ZN(n72) );
  NAND3_X1 U99 ( .A1(n70), .A2(n71), .A3(n72), .ZN(carry[15]) );
  XOR2_X1 U100 ( .A(B[7]), .B(A[7]), .Z(n73) );
  XOR2_X1 U101 ( .A(n46), .B(n73), .Z(SUM[7]) );
  NAND2_X1 U102 ( .A1(n45), .A2(B[7]), .ZN(n74) );
  NAND2_X1 U103 ( .A1(carry[7]), .A2(A[7]), .ZN(n75) );
  NAND2_X1 U104 ( .A1(B[7]), .A2(A[7]), .ZN(n76) );
  NAND3_X1 U105 ( .A1(n74), .A2(n75), .A3(n76), .ZN(carry[8]) );
  XOR2_X1 U106 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_19_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n307), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n306), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n310), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n309), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n312), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  BUF_X1 U157 ( .A(n302), .Z(n229) );
  AND2_X1 U158 ( .A1(n95), .A2(n102), .ZN(n206) );
  XOR2_X1 U159 ( .A(a[5]), .B(a[4]), .Z(n359) );
  NAND2_X1 U160 ( .A1(n237), .A2(n34), .ZN(n207) );
  NAND3_X1 U161 ( .A1(n217), .A2(n218), .A3(n219), .ZN(n208) );
  NAND3_X1 U162 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n209) );
  NAND3_X1 U163 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n210) );
  CLKBUF_X1 U164 ( .A(n208), .Z(n211) );
  CLKBUF_X3 U165 ( .A(a[3]), .Z(n212) );
  CLKBUF_X1 U166 ( .A(n322), .Z(n213) );
  CLKBUF_X1 U167 ( .A(n230), .Z(n214) );
  CLKBUF_X1 U168 ( .A(n207), .Z(n215) );
  XOR2_X1 U169 ( .A(n27), .B(n24), .Z(n216) );
  XOR2_X1 U170 ( .A(n210), .B(n216), .Z(product[10]) );
  NAND2_X1 U171 ( .A1(n209), .A2(n27), .ZN(n217) );
  NAND2_X1 U172 ( .A1(n6), .A2(n24), .ZN(n218) );
  NAND2_X1 U173 ( .A1(n27), .A2(n24), .ZN(n219) );
  NAND3_X1 U174 ( .A1(n217), .A2(n218), .A3(n219), .ZN(n5) );
  CLKBUF_X1 U175 ( .A(n295), .Z(n220) );
  CLKBUF_X1 U176 ( .A(b[1]), .Z(n221) );
  NAND2_X2 U177 ( .A1(n341), .A2(n360), .ZN(n343) );
  XOR2_X2 U178 ( .A(a[6]), .B(n308), .Z(n341) );
  AND2_X1 U179 ( .A1(n104), .A2(n72), .ZN(n222) );
  NAND3_X1 U180 ( .A1(n207), .A2(n270), .A3(n271), .ZN(n223) );
  NAND3_X1 U181 ( .A1(n215), .A2(n270), .A3(n271), .ZN(n224) );
  NAND3_X1 U182 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n225) );
  NAND3_X1 U183 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n226) );
  INV_X1 U184 ( .A(n302), .ZN(n227) );
  INV_X1 U185 ( .A(n302), .ZN(n228) );
  NAND3_X1 U186 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n230) );
  NAND2_X1 U187 ( .A1(a[4]), .A2(a[3]), .ZN(n233) );
  NAND2_X1 U188 ( .A1(n231), .A2(n232), .ZN(n234) );
  NAND2_X2 U189 ( .A1(n233), .A2(n234), .ZN(n330) );
  INV_X1 U190 ( .A(a[4]), .ZN(n231) );
  INV_X1 U191 ( .A(a[3]), .ZN(n232) );
  NAND3_X1 U192 ( .A1(n291), .A2(n290), .A3(n292), .ZN(n235) );
  NAND3_X1 U193 ( .A1(n265), .A2(n266), .A3(n267), .ZN(n236) );
  NAND3_X1 U194 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n237) );
  CLKBUF_X1 U195 ( .A(n287), .Z(n238) );
  XOR2_X1 U196 ( .A(n33), .B(n28), .Z(n239) );
  XOR2_X1 U197 ( .A(n224), .B(n239), .Z(product[9]) );
  NAND2_X1 U198 ( .A1(n223), .A2(n33), .ZN(n240) );
  NAND2_X1 U199 ( .A1(n7), .A2(n28), .ZN(n241) );
  NAND2_X1 U200 ( .A1(n33), .A2(n28), .ZN(n242) );
  NAND3_X1 U201 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n6) );
  NAND2_X1 U202 ( .A1(n10), .A2(n49), .ZN(n243) );
  CLKBUF_X1 U203 ( .A(n243), .Z(n244) );
  CLKBUF_X1 U204 ( .A(n300), .Z(n245) );
  XOR2_X1 U205 ( .A(n103), .B(n96), .Z(n246) );
  XOR2_X1 U206 ( .A(n222), .B(n246), .Z(product[2]) );
  NAND2_X1 U207 ( .A1(n222), .A2(n103), .ZN(n247) );
  NAND2_X1 U208 ( .A1(n14), .A2(n96), .ZN(n248) );
  NAND2_X1 U209 ( .A1(n103), .A2(n96), .ZN(n249) );
  NAND3_X1 U210 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n13) );
  CLKBUF_X1 U211 ( .A(n236), .Z(n250) );
  CLKBUF_X1 U212 ( .A(n237), .Z(n251) );
  NAND3_X1 U213 ( .A1(n299), .A2(n300), .A3(n301), .ZN(n252) );
  NAND3_X1 U214 ( .A1(n299), .A2(n245), .A3(n301), .ZN(n253) );
  NAND3_X1 U215 ( .A1(n257), .A2(n243), .A3(n259), .ZN(n254) );
  NAND3_X1 U216 ( .A1(n257), .A2(n244), .A3(n259), .ZN(n255) );
  XOR2_X1 U217 ( .A(n46), .B(n49), .Z(n256) );
  XOR2_X1 U218 ( .A(n253), .B(n256), .Z(product[6]) );
  NAND2_X1 U219 ( .A1(n252), .A2(n46), .ZN(n257) );
  NAND2_X1 U220 ( .A1(n10), .A2(n49), .ZN(n258) );
  NAND2_X1 U221 ( .A1(n46), .A2(n49), .ZN(n259) );
  NAND3_X1 U222 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n9) );
  XOR2_X1 U223 ( .A(n40), .B(n45), .Z(n260) );
  XOR2_X1 U224 ( .A(n255), .B(n260), .Z(product[7]) );
  NAND2_X1 U225 ( .A1(n254), .A2(n40), .ZN(n261) );
  NAND2_X1 U226 ( .A1(n9), .A2(n45), .ZN(n262) );
  NAND2_X1 U227 ( .A1(n40), .A2(n45), .ZN(n263) );
  NAND3_X1 U228 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n8) );
  XOR2_X1 U229 ( .A(n56), .B(n71), .Z(n264) );
  XOR2_X1 U230 ( .A(n214), .B(n264), .Z(product[3]) );
  NAND2_X1 U231 ( .A1(n230), .A2(n56), .ZN(n265) );
  NAND2_X1 U232 ( .A1(n13), .A2(n71), .ZN(n266) );
  NAND2_X1 U233 ( .A1(n56), .A2(n71), .ZN(n267) );
  NAND3_X1 U234 ( .A1(n265), .A2(n266), .A3(n267), .ZN(n12) );
  XOR2_X1 U235 ( .A(n34), .B(n39), .Z(n268) );
  XOR2_X1 U236 ( .A(n251), .B(n268), .Z(product[8]) );
  NAND2_X1 U237 ( .A1(n237), .A2(n34), .ZN(n269) );
  NAND2_X1 U238 ( .A1(n8), .A2(n39), .ZN(n270) );
  NAND2_X1 U239 ( .A1(n34), .A2(n39), .ZN(n271) );
  NAND3_X1 U240 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n7) );
  NAND3_X1 U241 ( .A1(n295), .A2(n296), .A3(n297), .ZN(n272) );
  XOR2_X1 U242 ( .A(n20), .B(n23), .Z(n273) );
  XOR2_X1 U243 ( .A(n211), .B(n273), .Z(product[11]) );
  NAND2_X1 U244 ( .A1(n208), .A2(n20), .ZN(n274) );
  NAND2_X1 U245 ( .A1(n5), .A2(n23), .ZN(n275) );
  NAND2_X1 U246 ( .A1(n20), .A2(n23), .ZN(n276) );
  NAND3_X1 U247 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n4) );
  XOR2_X1 U248 ( .A(n95), .B(n102), .Z(n56) );
  NAND3_X1 U249 ( .A1(n288), .A2(n287), .A3(n286), .ZN(n277) );
  NAND3_X1 U250 ( .A1(n288), .A2(n238), .A3(n286), .ZN(n278) );
  NAND2_X2 U251 ( .A1(n330), .A2(n359), .ZN(n332) );
  CLKBUF_X1 U252 ( .A(n320), .Z(n279) );
  XOR2_X2 U253 ( .A(a[2]), .B(n313), .Z(n320) );
  XNOR2_X1 U254 ( .A(n235), .B(n280), .ZN(product[14]) );
  XNOR2_X1 U255 ( .A(n304), .B(n15), .ZN(n280) );
  INV_X1 U256 ( .A(n15), .ZN(n303) );
  AND3_X1 U257 ( .A1(n282), .A2(n283), .A3(n284), .ZN(product[15]) );
  INV_X1 U258 ( .A(n339), .ZN(n307) );
  INV_X1 U259 ( .A(n21), .ZN(n306) );
  INV_X1 U260 ( .A(n319), .ZN(n312) );
  INV_X1 U261 ( .A(n328), .ZN(n310) );
  INV_X1 U262 ( .A(n31), .ZN(n309) );
  INV_X1 U263 ( .A(b[0]), .ZN(n302) );
  NAND2_X1 U264 ( .A1(n320), .A2(n358), .ZN(n322) );
  INV_X1 U265 ( .A(a[0]), .ZN(n314) );
  BUF_X1 U266 ( .A(a[1]), .Z(n293) );
  INV_X1 U267 ( .A(a[5]), .ZN(n308) );
  INV_X1 U268 ( .A(a[7]), .ZN(n305) );
  NAND2_X1 U269 ( .A1(n235), .A2(n304), .ZN(n282) );
  NAND2_X1 U270 ( .A1(n2), .A2(n15), .ZN(n283) );
  NAND2_X1 U271 ( .A1(n304), .A2(n15), .ZN(n284) );
  XOR2_X1 U272 ( .A(n19), .B(n18), .Z(n285) );
  XOR2_X1 U273 ( .A(n285), .B(n226), .Z(product[12]) );
  NAND2_X1 U274 ( .A1(n19), .A2(n18), .ZN(n286) );
  NAND2_X1 U275 ( .A1(n19), .A2(n4), .ZN(n287) );
  NAND2_X1 U276 ( .A1(n18), .A2(n225), .ZN(n288) );
  NAND3_X1 U277 ( .A1(n288), .A2(n287), .A3(n286), .ZN(n3) );
  XOR2_X1 U278 ( .A(n17), .B(n303), .Z(n289) );
  XOR2_X1 U279 ( .A(n289), .B(n278), .Z(product[13]) );
  NAND2_X1 U280 ( .A1(n17), .A2(n303), .ZN(n290) );
  NAND2_X1 U281 ( .A1(n17), .A2(n277), .ZN(n291) );
  NAND2_X1 U282 ( .A1(n3), .A2(n303), .ZN(n292) );
  NAND3_X1 U283 ( .A1(n290), .A2(n291), .A3(n292), .ZN(n2) );
  INV_X1 U284 ( .A(n350), .ZN(n304) );
  XOR2_X1 U285 ( .A(n54), .B(n206), .Z(n294) );
  XOR2_X1 U286 ( .A(n250), .B(n294), .Z(product[4]) );
  NAND2_X1 U287 ( .A1(n236), .A2(n54), .ZN(n295) );
  NAND2_X1 U288 ( .A1(n12), .A2(n206), .ZN(n296) );
  NAND2_X1 U289 ( .A1(n54), .A2(n206), .ZN(n297) );
  NAND3_X1 U290 ( .A1(n220), .A2(n296), .A3(n297), .ZN(n11) );
  XOR2_X1 U291 ( .A(n50), .B(n53), .Z(n298) );
  XOR2_X1 U292 ( .A(n11), .B(n298), .Z(product[5]) );
  NAND2_X1 U293 ( .A1(n272), .A2(n50), .ZN(n299) );
  NAND2_X1 U294 ( .A1(n272), .A2(n53), .ZN(n300) );
  NAND2_X1 U295 ( .A1(n50), .A2(n53), .ZN(n301) );
  NAND3_X1 U296 ( .A1(n299), .A2(n300), .A3(n301), .ZN(n10) );
  INV_X1 U297 ( .A(a[3]), .ZN(n311) );
  INV_X1 U298 ( .A(a[1]), .ZN(n313) );
  NOR2_X1 U299 ( .A1(n314), .A2(n229), .ZN(product[0]) );
  OAI22_X1 U300 ( .A1(n315), .A2(n316), .B1(n317), .B2(n314), .ZN(n99) );
  OAI22_X1 U301 ( .A1(n317), .A2(n316), .B1(n318), .B2(n314), .ZN(n98) );
  XNOR2_X1 U302 ( .A(b[6]), .B(n293), .ZN(n317) );
  OAI22_X1 U303 ( .A1(n314), .A2(n318), .B1(n316), .B2(n318), .ZN(n319) );
  XNOR2_X1 U304 ( .A(b[7]), .B(n293), .ZN(n318) );
  NOR2_X1 U305 ( .A1(n320), .A2(n229), .ZN(n96) );
  OAI22_X1 U306 ( .A1(n321), .A2(n322), .B1(n320), .B2(n323), .ZN(n95) );
  XNOR2_X1 U307 ( .A(n212), .B(n228), .ZN(n321) );
  OAI22_X1 U308 ( .A1(n323), .A2(n322), .B1(n320), .B2(n324), .ZN(n94) );
  XNOR2_X1 U309 ( .A(n221), .B(n212), .ZN(n323) );
  OAI22_X1 U310 ( .A1(n324), .A2(n322), .B1(n279), .B2(n325), .ZN(n93) );
  XNOR2_X1 U311 ( .A(b[2]), .B(n212), .ZN(n324) );
  OAI22_X1 U312 ( .A1(n325), .A2(n322), .B1(n279), .B2(n326), .ZN(n92) );
  XNOR2_X1 U313 ( .A(b[3]), .B(n212), .ZN(n325) );
  OAI22_X1 U314 ( .A1(n326), .A2(n213), .B1(n279), .B2(n327), .ZN(n91) );
  XNOR2_X1 U315 ( .A(b[4]), .B(n212), .ZN(n326) );
  OAI22_X1 U316 ( .A1(n329), .A2(n279), .B1(n213), .B2(n329), .ZN(n328) );
  NOR2_X1 U317 ( .A1(n330), .A2(n229), .ZN(n88) );
  OAI22_X1 U318 ( .A1(n331), .A2(n332), .B1(n330), .B2(n333), .ZN(n87) );
  XNOR2_X1 U319 ( .A(a[5]), .B(n227), .ZN(n331) );
  OAI22_X1 U320 ( .A1(n333), .A2(n332), .B1(n330), .B2(n334), .ZN(n86) );
  XNOR2_X1 U321 ( .A(b[1]), .B(a[5]), .ZN(n333) );
  OAI22_X1 U322 ( .A1(n334), .A2(n332), .B1(n330), .B2(n335), .ZN(n85) );
  XNOR2_X1 U323 ( .A(b[2]), .B(a[5]), .ZN(n334) );
  OAI22_X1 U324 ( .A1(n335), .A2(n332), .B1(n330), .B2(n336), .ZN(n84) );
  XNOR2_X1 U325 ( .A(b[3]), .B(a[5]), .ZN(n335) );
  OAI22_X1 U326 ( .A1(n336), .A2(n332), .B1(n330), .B2(n337), .ZN(n83) );
  XNOR2_X1 U327 ( .A(b[4]), .B(a[5]), .ZN(n336) );
  OAI22_X1 U328 ( .A1(n337), .A2(n332), .B1(n330), .B2(n338), .ZN(n82) );
  XNOR2_X1 U329 ( .A(b[5]), .B(a[5]), .ZN(n337) );
  OAI22_X1 U330 ( .A1(n340), .A2(n330), .B1(n332), .B2(n340), .ZN(n339) );
  NOR2_X1 U331 ( .A1(n341), .A2(n229), .ZN(n80) );
  OAI22_X1 U332 ( .A1(n342), .A2(n343), .B1(n341), .B2(n344), .ZN(n79) );
  XNOR2_X1 U333 ( .A(a[7]), .B(n227), .ZN(n342) );
  OAI22_X1 U334 ( .A1(n345), .A2(n343), .B1(n341), .B2(n346), .ZN(n77) );
  OAI22_X1 U335 ( .A1(n346), .A2(n343), .B1(n341), .B2(n347), .ZN(n76) );
  XNOR2_X1 U336 ( .A(b[3]), .B(a[7]), .ZN(n346) );
  OAI22_X1 U337 ( .A1(n347), .A2(n343), .B1(n341), .B2(n348), .ZN(n75) );
  XNOR2_X1 U338 ( .A(b[4]), .B(a[7]), .ZN(n347) );
  OAI22_X1 U339 ( .A1(n348), .A2(n343), .B1(n341), .B2(n349), .ZN(n74) );
  XNOR2_X1 U340 ( .A(b[5]), .B(a[7]), .ZN(n348) );
  OAI22_X1 U341 ( .A1(n351), .A2(n341), .B1(n343), .B2(n351), .ZN(n350) );
  OAI21_X1 U342 ( .B1(n228), .B2(n313), .A(n316), .ZN(n72) );
  OAI21_X1 U343 ( .B1(n311), .B2(n322), .A(n352), .ZN(n71) );
  OR3_X1 U344 ( .A1(n320), .A2(n228), .A3(n311), .ZN(n352) );
  OAI21_X1 U345 ( .B1(n308), .B2(n332), .A(n353), .ZN(n70) );
  OR3_X1 U346 ( .A1(n330), .A2(b[0]), .A3(n308), .ZN(n353) );
  OAI21_X1 U347 ( .B1(n305), .B2(n343), .A(n354), .ZN(n69) );
  OR3_X1 U348 ( .A1(n341), .A2(n228), .A3(n305), .ZN(n354) );
  XNOR2_X1 U349 ( .A(n355), .B(n356), .ZN(n38) );
  OR2_X1 U350 ( .A1(n355), .A2(n356), .ZN(n37) );
  OAI22_X1 U351 ( .A1(n327), .A2(n213), .B1(n279), .B2(n357), .ZN(n356) );
  XNOR2_X1 U352 ( .A(b[5]), .B(n212), .ZN(n327) );
  OAI22_X1 U353 ( .A1(n344), .A2(n343), .B1(n341), .B2(n345), .ZN(n355) );
  XNOR2_X1 U354 ( .A(b[2]), .B(a[7]), .ZN(n345) );
  XNOR2_X1 U355 ( .A(b[1]), .B(a[7]), .ZN(n344) );
  OAI22_X1 U356 ( .A1(n357), .A2(n213), .B1(n279), .B2(n329), .ZN(n31) );
  XNOR2_X1 U357 ( .A(b[7]), .B(n212), .ZN(n329) );
  XNOR2_X1 U358 ( .A(n311), .B(a[2]), .ZN(n358) );
  XNOR2_X1 U359 ( .A(b[6]), .B(n212), .ZN(n357) );
  OAI22_X1 U360 ( .A1(n338), .A2(n332), .B1(n330), .B2(n340), .ZN(n21) );
  XNOR2_X1 U361 ( .A(b[7]), .B(a[5]), .ZN(n340) );
  XNOR2_X1 U362 ( .A(b[6]), .B(a[5]), .ZN(n338) );
  OAI22_X1 U363 ( .A1(n349), .A2(n343), .B1(n341), .B2(n351), .ZN(n15) );
  XNOR2_X1 U364 ( .A(b[7]), .B(a[7]), .ZN(n351) );
  XNOR2_X1 U365 ( .A(n305), .B(a[6]), .ZN(n360) );
  XNOR2_X1 U366 ( .A(b[6]), .B(a[7]), .ZN(n349) );
  OAI22_X1 U367 ( .A1(n227), .A2(n316), .B1(n361), .B2(n314), .ZN(n104) );
  OAI22_X1 U368 ( .A1(n316), .A2(n361), .B1(n362), .B2(n314), .ZN(n103) );
  XNOR2_X1 U369 ( .A(b[1]), .B(n293), .ZN(n361) );
  OAI22_X1 U370 ( .A1(n362), .A2(n316), .B1(n363), .B2(n314), .ZN(n102) );
  XNOR2_X1 U371 ( .A(b[2]), .B(n293), .ZN(n362) );
  OAI22_X1 U372 ( .A1(n363), .A2(n316), .B1(n364), .B2(n314), .ZN(n101) );
  XNOR2_X1 U373 ( .A(b[3]), .B(n293), .ZN(n363) );
  OAI22_X1 U374 ( .A1(n364), .A2(n316), .B1(n315), .B2(n314), .ZN(n100) );
  XNOR2_X1 U375 ( .A(b[5]), .B(n293), .ZN(n315) );
  NAND2_X1 U376 ( .A1(a[1]), .A2(n314), .ZN(n316) );
  XNOR2_X1 U377 ( .A(b[4]), .B(n293), .ZN(n364) );
endmodule


module mac_19 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_19_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_19_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_18_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88;
  wire   [15:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .S(SUM[15]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n88) );
  CLKBUF_X1 U2 ( .A(n27), .Z(n1) );
  CLKBUF_X1 U3 ( .A(n55), .Z(n2) );
  NAND2_X1 U4 ( .A1(n9), .A2(A[8]), .ZN(n3) );
  CLKBUF_X1 U5 ( .A(n51), .Z(n4) );
  CLKBUF_X1 U6 ( .A(n82), .Z(n5) );
  CLKBUF_X1 U7 ( .A(n73), .Z(n6) );
  CLKBUF_X1 U8 ( .A(carry[14]), .Z(n7) );
  CLKBUF_X1 U9 ( .A(carry[10]), .Z(n8) );
  NAND3_X1 U10 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n9) );
  NAND3_X1 U11 ( .A1(n23), .A2(n22), .A3(n24), .ZN(n10) );
  XOR2_X1 U12 ( .A(B[14]), .B(A[14]), .Z(n11) );
  XOR2_X1 U13 ( .A(n7), .B(n11), .Z(SUM[14]) );
  NAND2_X1 U14 ( .A1(n10), .A2(B[14]), .ZN(n12) );
  NAND2_X1 U15 ( .A1(carry[14]), .A2(A[14]), .ZN(n13) );
  NAND2_X1 U16 ( .A1(B[14]), .A2(A[14]), .ZN(n14) );
  NAND3_X1 U17 ( .A1(n12), .A2(n13), .A3(n14), .ZN(carry[15]) );
  NAND3_X1 U18 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n15) );
  NAND3_X1 U19 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n16) );
  NAND3_X1 U20 ( .A1(n4), .A2(n52), .A3(n53), .ZN(n17) );
  NAND3_X1 U21 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n18) );
  NAND3_X1 U22 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n19) );
  NAND3_X1 U23 ( .A1(n1), .A2(n28), .A3(n29), .ZN(n20) );
  XOR2_X1 U24 ( .A(B[13]), .B(A[13]), .Z(n21) );
  XOR2_X1 U25 ( .A(n17), .B(n21), .Z(SUM[13]) );
  NAND2_X1 U26 ( .A1(n16), .A2(B[13]), .ZN(n22) );
  NAND2_X1 U27 ( .A1(carry[13]), .A2(A[13]), .ZN(n23) );
  NAND2_X1 U28 ( .A1(B[13]), .A2(A[13]), .ZN(n24) );
  NAND3_X1 U29 ( .A1(n22), .A2(n23), .A3(n24), .ZN(carry[14]) );
  CLKBUF_X1 U30 ( .A(n48), .Z(n25) );
  XOR2_X1 U31 ( .A(B[5]), .B(A[5]), .Z(n26) );
  XOR2_X1 U32 ( .A(n18), .B(n26), .Z(SUM[5]) );
  NAND2_X1 U33 ( .A1(n18), .A2(B[5]), .ZN(n27) );
  NAND2_X1 U34 ( .A1(carry[5]), .A2(A[5]), .ZN(n28) );
  NAND2_X1 U35 ( .A1(B[5]), .A2(A[5]), .ZN(n29) );
  NAND3_X1 U36 ( .A1(n27), .A2(n28), .A3(n29), .ZN(carry[6]) );
  CLKBUF_X1 U37 ( .A(n15), .Z(n30) );
  NAND3_X1 U38 ( .A1(n85), .A2(n86), .A3(n87), .ZN(n31) );
  NAND3_X1 U39 ( .A1(n35), .A2(n36), .A3(n37), .ZN(n32) );
  NAND3_X1 U40 ( .A1(n35), .A2(n36), .A3(n37), .ZN(n33) );
  XOR2_X1 U41 ( .A(B[3]), .B(A[3]), .Z(n34) );
  XOR2_X1 U42 ( .A(n31), .B(n34), .Z(SUM[3]) );
  NAND2_X1 U43 ( .A1(n31), .A2(B[3]), .ZN(n35) );
  NAND2_X1 U44 ( .A1(carry[3]), .A2(A[3]), .ZN(n36) );
  NAND2_X1 U45 ( .A1(B[3]), .A2(A[3]), .ZN(n37) );
  NAND3_X1 U46 ( .A1(n35), .A2(n36), .A3(n37), .ZN(carry[4]) );
  XOR2_X1 U47 ( .A(B[4]), .B(A[4]), .Z(n38) );
  XOR2_X1 U48 ( .A(n33), .B(n38), .Z(SUM[4]) );
  NAND2_X1 U49 ( .A1(n32), .A2(B[4]), .ZN(n39) );
  NAND2_X1 U50 ( .A1(carry[4]), .A2(A[4]), .ZN(n40) );
  NAND2_X1 U51 ( .A1(B[4]), .A2(A[4]), .ZN(n41) );
  NAND3_X1 U52 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[5]) );
  CLKBUF_X1 U53 ( .A(n3), .Z(n42) );
  NAND3_X1 U54 ( .A1(n62), .A2(n61), .A3(n63), .ZN(n43) );
  XOR2_X1 U55 ( .A(B[6]), .B(A[6]), .Z(n44) );
  XOR2_X1 U56 ( .A(n20), .B(n44), .Z(SUM[6]) );
  NAND2_X1 U57 ( .A1(n19), .A2(B[6]), .ZN(n45) );
  NAND2_X1 U58 ( .A1(carry[6]), .A2(A[6]), .ZN(n46) );
  NAND2_X1 U59 ( .A1(B[6]), .A2(A[6]), .ZN(n47) );
  NAND3_X1 U60 ( .A1(n45), .A2(n46), .A3(n47), .ZN(carry[7]) );
  NAND3_X1 U61 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n48) );
  NAND3_X1 U62 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n49) );
  XOR2_X1 U63 ( .A(B[12]), .B(A[12]), .Z(n50) );
  XOR2_X1 U64 ( .A(n25), .B(n50), .Z(SUM[12]) );
  NAND2_X1 U65 ( .A1(n48), .A2(B[12]), .ZN(n51) );
  NAND2_X1 U66 ( .A1(carry[12]), .A2(A[12]), .ZN(n52) );
  NAND2_X1 U67 ( .A1(B[12]), .A2(A[12]), .ZN(n53) );
  NAND3_X1 U68 ( .A1(n51), .A2(n52), .A3(n53), .ZN(carry[13]) );
  XOR2_X1 U69 ( .A(B[7]), .B(A[7]), .Z(n54) );
  XOR2_X1 U70 ( .A(n30), .B(n54), .Z(SUM[7]) );
  NAND2_X1 U71 ( .A1(n15), .A2(B[7]), .ZN(n55) );
  NAND2_X1 U72 ( .A1(carry[7]), .A2(A[7]), .ZN(n56) );
  NAND2_X1 U73 ( .A1(B[7]), .A2(A[7]), .ZN(n57) );
  NAND3_X1 U74 ( .A1(n2), .A2(n56), .A3(n57), .ZN(carry[8]) );
  CLKBUF_X1 U75 ( .A(n43), .Z(n58) );
  NAND3_X1 U76 ( .A1(n78), .A2(n77), .A3(n79), .ZN(n59) );
  XOR2_X1 U77 ( .A(B[10]), .B(A[10]), .Z(n60) );
  XOR2_X1 U78 ( .A(n8), .B(n60), .Z(SUM[10]) );
  NAND2_X1 U79 ( .A1(n59), .A2(B[10]), .ZN(n61) );
  NAND2_X1 U80 ( .A1(carry[10]), .A2(A[10]), .ZN(n62) );
  NAND2_X1 U81 ( .A1(B[10]), .A2(A[10]), .ZN(n63) );
  NAND3_X1 U82 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[11]) );
  XOR2_X1 U83 ( .A(B[11]), .B(A[11]), .Z(n64) );
  XOR2_X1 U84 ( .A(n58), .B(n64), .Z(SUM[11]) );
  NAND2_X1 U85 ( .A1(n43), .A2(B[11]), .ZN(n65) );
  NAND2_X1 U86 ( .A1(carry[11]), .A2(A[11]), .ZN(n66) );
  NAND2_X1 U87 ( .A1(B[11]), .A2(A[11]), .ZN(n67) );
  NAND3_X1 U88 ( .A1(n65), .A2(n66), .A3(n67), .ZN(carry[12]) );
  NAND3_X1 U89 ( .A1(n81), .A2(n82), .A3(n83), .ZN(n68) );
  NAND3_X1 U90 ( .A1(n81), .A2(n5), .A3(n83), .ZN(n69) );
  NAND3_X1 U91 ( .A1(n3), .A2(n73), .A3(n75), .ZN(n70) );
  NAND3_X1 U92 ( .A1(n6), .A2(n42), .A3(n75), .ZN(n71) );
  XOR2_X1 U93 ( .A(B[8]), .B(A[8]), .Z(n72) );
  XOR2_X1 U94 ( .A(carry[8]), .B(n72), .Z(SUM[8]) );
  NAND2_X1 U95 ( .A1(n49), .A2(B[8]), .ZN(n73) );
  NAND2_X1 U96 ( .A1(n9), .A2(A[8]), .ZN(n74) );
  NAND2_X1 U97 ( .A1(B[8]), .A2(A[8]), .ZN(n75) );
  NAND3_X1 U98 ( .A1(n73), .A2(n74), .A3(n75), .ZN(carry[9]) );
  XOR2_X1 U99 ( .A(B[9]), .B(A[9]), .Z(n76) );
  XOR2_X1 U100 ( .A(n71), .B(n76), .Z(SUM[9]) );
  NAND2_X1 U101 ( .A1(n70), .A2(B[9]), .ZN(n77) );
  NAND2_X1 U102 ( .A1(carry[9]), .A2(A[9]), .ZN(n78) );
  NAND2_X1 U103 ( .A1(B[9]), .A2(A[9]), .ZN(n79) );
  NAND3_X1 U104 ( .A1(n77), .A2(n78), .A3(n79), .ZN(carry[10]) );
  XOR2_X1 U105 ( .A(B[1]), .B(A[1]), .Z(n80) );
  XOR2_X1 U106 ( .A(n88), .B(n80), .Z(SUM[1]) );
  NAND2_X1 U107 ( .A1(n88), .A2(B[1]), .ZN(n81) );
  NAND2_X1 U108 ( .A1(n88), .A2(A[1]), .ZN(n82) );
  NAND2_X1 U109 ( .A1(B[1]), .A2(A[1]), .ZN(n83) );
  NAND3_X1 U110 ( .A1(n81), .A2(n82), .A3(n83), .ZN(carry[2]) );
  XOR2_X1 U111 ( .A(B[2]), .B(A[2]), .Z(n84) );
  XOR2_X1 U112 ( .A(n69), .B(n84), .Z(SUM[2]) );
  NAND2_X1 U113 ( .A1(n68), .A2(B[2]), .ZN(n85) );
  NAND2_X1 U114 ( .A1(carry[2]), .A2(A[2]), .ZN(n86) );
  NAND2_X1 U115 ( .A1(B[2]), .A2(A[2]), .ZN(n87) );
  NAND3_X1 U116 ( .A1(n85), .A2(n86), .A3(n87), .ZN(carry[3]) );
  XOR2_X1 U117 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_18_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n300), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n299), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n303), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n302), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n305), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  BUF_X1 U157 ( .A(b[2]), .Z(n220) );
  INV_X1 U158 ( .A(n295), .ZN(n294) );
  NAND2_X1 U159 ( .A1(n313), .A2(n351), .ZN(n315) );
  NOR2_X1 U160 ( .A1(n276), .A2(n275), .ZN(n96) );
  AND2_X1 U161 ( .A1(n95), .A2(n102), .ZN(n206) );
  NAND3_X1 U162 ( .A1(n216), .A2(n217), .A3(n218), .ZN(n207) );
  NAND3_X1 U163 ( .A1(n216), .A2(n217), .A3(n218), .ZN(n208) );
  NAND3_X1 U164 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n209) );
  NAND3_X1 U165 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n210) );
  NAND3_X1 U166 ( .A1(n291), .A2(n292), .A3(n293), .ZN(n211) );
  NAND3_X1 U167 ( .A1(n291), .A2(n292), .A3(n293), .ZN(n212) );
  XNOR2_X1 U168 ( .A(a[6]), .B(a[5]), .ZN(n334) );
  XNOR2_X1 U169 ( .A(a[6]), .B(a[5]), .ZN(n213) );
  NAND3_X1 U170 ( .A1(n230), .A2(n231), .A3(n232), .ZN(n214) );
  XOR2_X1 U171 ( .A(n56), .B(n71), .Z(n215) );
  XOR2_X1 U172 ( .A(n210), .B(n215), .Z(product[3]) );
  NAND2_X1 U173 ( .A1(n209), .A2(n56), .ZN(n216) );
  NAND2_X1 U174 ( .A1(n13), .A2(n71), .ZN(n217) );
  NAND2_X1 U175 ( .A1(n56), .A2(n71), .ZN(n218) );
  NAND3_X1 U176 ( .A1(n216), .A2(n217), .A3(n218), .ZN(n12) );
  NAND2_X1 U177 ( .A1(n323), .A2(n352), .ZN(n219) );
  NAND2_X1 U178 ( .A1(n323), .A2(n352), .ZN(n325) );
  CLKBUF_X1 U179 ( .A(b[3]), .Z(n221) );
  AND2_X1 U180 ( .A1(n104), .A2(n72), .ZN(n222) );
  XOR2_X1 U181 ( .A(a[3]), .B(a[2]), .Z(n351) );
  XOR2_X1 U182 ( .A(n103), .B(n96), .Z(n223) );
  XOR2_X1 U183 ( .A(n222), .B(n223), .Z(product[2]) );
  NAND2_X1 U184 ( .A1(n222), .A2(n103), .ZN(n224) );
  NAND2_X1 U185 ( .A1(n14), .A2(n96), .ZN(n225) );
  NAND2_X1 U186 ( .A1(n103), .A2(n96), .ZN(n226) );
  NAND3_X1 U187 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n13) );
  NAND3_X1 U188 ( .A1(n230), .A2(n231), .A3(n232), .ZN(n227) );
  NAND3_X1 U189 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n228) );
  XOR2_X1 U190 ( .A(n54), .B(n206), .Z(n229) );
  XOR2_X1 U191 ( .A(n208), .B(n229), .Z(product[4]) );
  NAND2_X1 U192 ( .A1(n12), .A2(n54), .ZN(n230) );
  NAND2_X1 U193 ( .A1(n207), .A2(n206), .ZN(n231) );
  NAND2_X1 U194 ( .A1(n54), .A2(n206), .ZN(n232) );
  NAND3_X1 U195 ( .A1(n230), .A2(n231), .A3(n232), .ZN(n11) );
  CLKBUF_X1 U196 ( .A(n7), .Z(n233) );
  NAND3_X1 U197 ( .A1(n266), .A2(n265), .A3(n267), .ZN(n234) );
  CLKBUF_X1 U198 ( .A(n270), .Z(n235) );
  XOR2_X1 U199 ( .A(n34), .B(n39), .Z(n236) );
  XOR2_X1 U200 ( .A(n212), .B(n236), .Z(product[8]) );
  NAND2_X1 U201 ( .A1(n211), .A2(n34), .ZN(n237) );
  NAND2_X1 U202 ( .A1(n8), .A2(n39), .ZN(n238) );
  NAND2_X1 U203 ( .A1(n34), .A2(n39), .ZN(n239) );
  NAND3_X1 U204 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n7) );
  CLKBUF_X1 U205 ( .A(n6), .Z(n240) );
  CLKBUF_X1 U206 ( .A(n244), .Z(n241) );
  NAND3_X1 U207 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n242) );
  CLKBUF_X1 U208 ( .A(n234), .Z(n243) );
  NAND3_X1 U209 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n244) );
  NAND3_X1 U210 ( .A1(n287), .A2(n288), .A3(n289), .ZN(n245) );
  XOR2_X1 U211 ( .A(n50), .B(n53), .Z(n246) );
  XOR2_X1 U212 ( .A(n11), .B(n246), .Z(product[5]) );
  NAND2_X1 U213 ( .A1(n214), .A2(n50), .ZN(n247) );
  NAND2_X1 U214 ( .A1(n227), .A2(n53), .ZN(n248) );
  NAND2_X1 U215 ( .A1(n50), .A2(n53), .ZN(n249) );
  NAND3_X1 U216 ( .A1(n248), .A2(n247), .A3(n249), .ZN(n10) );
  CLKBUF_X1 U217 ( .A(b[1]), .Z(n250) );
  CLKBUF_X1 U218 ( .A(n242), .Z(n251) );
  XOR2_X1 U219 ( .A(n33), .B(n28), .Z(n252) );
  XOR2_X1 U220 ( .A(n233), .B(n252), .Z(product[9]) );
  NAND2_X1 U221 ( .A1(n7), .A2(n33), .ZN(n253) );
  NAND2_X1 U222 ( .A1(n7), .A2(n28), .ZN(n254) );
  NAND2_X1 U223 ( .A1(n33), .A2(n28), .ZN(n255) );
  NAND3_X1 U224 ( .A1(n254), .A2(n253), .A3(n255), .ZN(n6) );
  XOR2_X1 U225 ( .A(n20), .B(n23), .Z(n256) );
  XOR2_X1 U226 ( .A(n243), .B(n256), .Z(product[11]) );
  NAND2_X1 U227 ( .A1(n234), .A2(n20), .ZN(n257) );
  NAND2_X1 U228 ( .A1(n5), .A2(n23), .ZN(n258) );
  NAND2_X1 U229 ( .A1(n20), .A2(n23), .ZN(n259) );
  NAND3_X1 U230 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n4) );
  XNOR2_X1 U231 ( .A(b[1]), .B(a[1]), .ZN(n260) );
  NAND3_X1 U232 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n261) );
  NAND3_X1 U233 ( .A1(n235), .A2(n271), .A3(n272), .ZN(n262) );
  NAND3_X1 U234 ( .A1(n281), .A2(n282), .A3(n280), .ZN(n263) );
  XOR2_X1 U235 ( .A(n27), .B(n24), .Z(n264) );
  XOR2_X1 U236 ( .A(n240), .B(n264), .Z(product[10]) );
  NAND2_X1 U237 ( .A1(n228), .A2(n27), .ZN(n265) );
  NAND2_X1 U238 ( .A1(n6), .A2(n24), .ZN(n266) );
  NAND2_X1 U239 ( .A1(n27), .A2(n24), .ZN(n267) );
  NAND3_X1 U240 ( .A1(n266), .A2(n265), .A3(n267), .ZN(n5) );
  XNOR2_X1 U241 ( .A(a[2]), .B(a[1]), .ZN(n313) );
  XNOR2_X1 U242 ( .A(n268), .B(n263), .ZN(product[14]) );
  XNOR2_X1 U243 ( .A(n297), .B(n15), .ZN(n268) );
  XOR2_X1 U244 ( .A(n18), .B(n19), .Z(n269) );
  XOR2_X1 U245 ( .A(n251), .B(n269), .Z(product[12]) );
  NAND2_X1 U246 ( .A1(n242), .A2(n18), .ZN(n270) );
  NAND2_X1 U247 ( .A1(n4), .A2(n19), .ZN(n271) );
  NAND2_X1 U248 ( .A1(n18), .A2(n19), .ZN(n272) );
  NAND3_X1 U249 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n3) );
  CLKBUF_X1 U250 ( .A(n245), .Z(n273) );
  INV_X1 U251 ( .A(n295), .ZN(n274) );
  INV_X1 U252 ( .A(n274), .ZN(n275) );
  XOR2_X1 U253 ( .A(n95), .B(n102), .Z(n56) );
  XNOR2_X2 U254 ( .A(a[4]), .B(a[3]), .ZN(n323) );
  XOR2_X1 U255 ( .A(a[2]), .B(n306), .Z(n276) );
  XOR2_X1 U256 ( .A(a[2]), .B(n306), .Z(n277) );
  INV_X1 U257 ( .A(n15), .ZN(n296) );
  AND3_X1 U258 ( .A1(n285), .A2(n284), .A3(n283), .ZN(product[15]) );
  INV_X1 U259 ( .A(n343), .ZN(n297) );
  INV_X1 U260 ( .A(n21), .ZN(n299) );
  INV_X1 U261 ( .A(n332), .ZN(n300) );
  INV_X1 U262 ( .A(n312), .ZN(n305) );
  INV_X1 U263 ( .A(n321), .ZN(n303) );
  INV_X1 U264 ( .A(n31), .ZN(n302) );
  INV_X1 U265 ( .A(b[0]), .ZN(n295) );
  INV_X1 U266 ( .A(a[0]), .ZN(n307) );
  INV_X1 U267 ( .A(a[5]), .ZN(n301) );
  INV_X1 U268 ( .A(a[7]), .ZN(n298) );
  XOR2_X1 U269 ( .A(n17), .B(n296), .Z(n279) );
  XOR2_X1 U270 ( .A(n279), .B(n262), .Z(product[13]) );
  NAND2_X1 U271 ( .A1(n17), .A2(n296), .ZN(n280) );
  NAND2_X1 U272 ( .A1(n17), .A2(n3), .ZN(n281) );
  NAND2_X1 U273 ( .A1(n261), .A2(n296), .ZN(n282) );
  NAND3_X1 U274 ( .A1(n281), .A2(n282), .A3(n280), .ZN(n2) );
  NAND2_X1 U275 ( .A1(n297), .A2(n15), .ZN(n283) );
  NAND2_X1 U276 ( .A1(n297), .A2(n2), .ZN(n284) );
  NAND2_X1 U277 ( .A1(n263), .A2(n15), .ZN(n285) );
  INV_X1 U278 ( .A(a[3]), .ZN(n304) );
  XOR2_X1 U279 ( .A(n46), .B(n49), .Z(n286) );
  XOR2_X1 U280 ( .A(n241), .B(n286), .Z(product[6]) );
  NAND2_X1 U281 ( .A1(n244), .A2(n46), .ZN(n287) );
  NAND2_X1 U282 ( .A1(n10), .A2(n49), .ZN(n288) );
  NAND2_X1 U283 ( .A1(n46), .A2(n49), .ZN(n289) );
  NAND3_X1 U284 ( .A1(n287), .A2(n288), .A3(n289), .ZN(n9) );
  XOR2_X1 U285 ( .A(n40), .B(n45), .Z(n290) );
  XOR2_X1 U286 ( .A(n273), .B(n290), .Z(product[7]) );
  NAND2_X1 U287 ( .A1(n245), .A2(n40), .ZN(n291) );
  NAND2_X1 U288 ( .A1(n9), .A2(n45), .ZN(n292) );
  NAND2_X1 U289 ( .A1(n40), .A2(n45), .ZN(n293) );
  NAND3_X1 U290 ( .A1(n291), .A2(n292), .A3(n293), .ZN(n8) );
  INV_X1 U291 ( .A(a[1]), .ZN(n306) );
  NOR2_X1 U292 ( .A1(n307), .A2(n275), .ZN(product[0]) );
  OAI22_X1 U293 ( .A1(n308), .A2(n309), .B1(n310), .B2(n307), .ZN(n99) );
  OAI22_X1 U294 ( .A1(n310), .A2(n309), .B1(n311), .B2(n307), .ZN(n98) );
  XNOR2_X1 U295 ( .A(b[6]), .B(a[1]), .ZN(n310) );
  OAI22_X1 U296 ( .A1(n307), .A2(n311), .B1(n309), .B2(n311), .ZN(n312) );
  XNOR2_X1 U297 ( .A(b[7]), .B(a[1]), .ZN(n311) );
  OAI22_X1 U298 ( .A1(n314), .A2(n315), .B1(n277), .B2(n316), .ZN(n95) );
  XNOR2_X1 U299 ( .A(a[3]), .B(n294), .ZN(n314) );
  OAI22_X1 U300 ( .A1(n316), .A2(n315), .B1(n277), .B2(n317), .ZN(n94) );
  XNOR2_X1 U301 ( .A(b[1]), .B(a[3]), .ZN(n316) );
  OAI22_X1 U302 ( .A1(n317), .A2(n315), .B1(n277), .B2(n318), .ZN(n93) );
  XNOR2_X1 U303 ( .A(n220), .B(a[3]), .ZN(n317) );
  OAI22_X1 U304 ( .A1(n318), .A2(n315), .B1(n276), .B2(n319), .ZN(n92) );
  XNOR2_X1 U305 ( .A(b[3]), .B(a[3]), .ZN(n318) );
  OAI22_X1 U306 ( .A1(n319), .A2(n315), .B1(n277), .B2(n320), .ZN(n91) );
  XNOR2_X1 U307 ( .A(b[4]), .B(a[3]), .ZN(n319) );
  OAI22_X1 U308 ( .A1(n322), .A2(n276), .B1(n315), .B2(n322), .ZN(n321) );
  NOR2_X1 U309 ( .A1(n323), .A2(n275), .ZN(n88) );
  OAI22_X1 U310 ( .A1(n324), .A2(n325), .B1(n323), .B2(n326), .ZN(n87) );
  XNOR2_X1 U311 ( .A(a[5]), .B(n274), .ZN(n324) );
  OAI22_X1 U312 ( .A1(n326), .A2(n219), .B1(n323), .B2(n327), .ZN(n86) );
  XNOR2_X1 U313 ( .A(a[5]), .B(b[1]), .ZN(n326) );
  OAI22_X1 U314 ( .A1(n327), .A2(n219), .B1(n323), .B2(n328), .ZN(n85) );
  XNOR2_X1 U315 ( .A(n220), .B(a[5]), .ZN(n327) );
  OAI22_X1 U316 ( .A1(n328), .A2(n219), .B1(n323), .B2(n329), .ZN(n84) );
  XNOR2_X1 U317 ( .A(n221), .B(a[5]), .ZN(n328) );
  OAI22_X1 U318 ( .A1(n329), .A2(n219), .B1(n323), .B2(n330), .ZN(n83) );
  XNOR2_X1 U319 ( .A(b[4]), .B(a[5]), .ZN(n329) );
  OAI22_X1 U320 ( .A1(n330), .A2(n219), .B1(n323), .B2(n331), .ZN(n82) );
  XNOR2_X1 U321 ( .A(b[5]), .B(a[5]), .ZN(n330) );
  OAI22_X1 U322 ( .A1(n333), .A2(n323), .B1(n219), .B2(n333), .ZN(n332) );
  NOR2_X1 U323 ( .A1(n334), .A2(n275), .ZN(n80) );
  OAI22_X1 U324 ( .A1(n335), .A2(n336), .B1(n213), .B2(n337), .ZN(n79) );
  XNOR2_X1 U325 ( .A(a[7]), .B(n294), .ZN(n335) );
  OAI22_X1 U326 ( .A1(n338), .A2(n336), .B1(n213), .B2(n339), .ZN(n77) );
  OAI22_X1 U327 ( .A1(n339), .A2(n336), .B1(n213), .B2(n340), .ZN(n76) );
  XNOR2_X1 U328 ( .A(n221), .B(a[7]), .ZN(n339) );
  OAI22_X1 U329 ( .A1(n340), .A2(n336), .B1(n213), .B2(n341), .ZN(n75) );
  XNOR2_X1 U330 ( .A(b[4]), .B(a[7]), .ZN(n340) );
  OAI22_X1 U331 ( .A1(n341), .A2(n336), .B1(n213), .B2(n342), .ZN(n74) );
  XNOR2_X1 U332 ( .A(b[5]), .B(a[7]), .ZN(n341) );
  OAI22_X1 U333 ( .A1(n344), .A2(n213), .B1(n336), .B2(n344), .ZN(n343) );
  OAI21_X1 U334 ( .B1(n294), .B2(n306), .A(n309), .ZN(n72) );
  OAI21_X1 U335 ( .B1(n304), .B2(n315), .A(n345), .ZN(n71) );
  OR3_X1 U336 ( .A1(n276), .A2(n294), .A3(n304), .ZN(n345) );
  OAI21_X1 U337 ( .B1(n301), .B2(n325), .A(n346), .ZN(n70) );
  OR3_X1 U338 ( .A1(n323), .A2(n294), .A3(n301), .ZN(n346) );
  OAI21_X1 U339 ( .B1(n298), .B2(n336), .A(n347), .ZN(n69) );
  OR3_X1 U340 ( .A1(n213), .A2(n274), .A3(n298), .ZN(n347) );
  XNOR2_X1 U341 ( .A(n348), .B(n349), .ZN(n38) );
  OR2_X1 U342 ( .A1(n348), .A2(n349), .ZN(n37) );
  OAI22_X1 U343 ( .A1(n320), .A2(n315), .B1(n276), .B2(n350), .ZN(n349) );
  XNOR2_X1 U344 ( .A(b[5]), .B(a[3]), .ZN(n320) );
  OAI22_X1 U345 ( .A1(n337), .A2(n336), .B1(n213), .B2(n338), .ZN(n348) );
  XNOR2_X1 U346 ( .A(n220), .B(a[7]), .ZN(n338) );
  XNOR2_X1 U347 ( .A(n250), .B(a[7]), .ZN(n337) );
  OAI22_X1 U348 ( .A1(n350), .A2(n315), .B1(n277), .B2(n322), .ZN(n31) );
  XNOR2_X1 U349 ( .A(b[7]), .B(a[3]), .ZN(n322) );
  XNOR2_X1 U350 ( .A(b[6]), .B(a[3]), .ZN(n350) );
  OAI22_X1 U351 ( .A1(n331), .A2(n219), .B1(n323), .B2(n333), .ZN(n21) );
  XNOR2_X1 U352 ( .A(b[7]), .B(a[5]), .ZN(n333) );
  XNOR2_X1 U353 ( .A(n301), .B(a[4]), .ZN(n352) );
  XNOR2_X1 U354 ( .A(b[6]), .B(a[5]), .ZN(n331) );
  OAI22_X1 U355 ( .A1(n342), .A2(n336), .B1(n213), .B2(n344), .ZN(n15) );
  XNOR2_X1 U356 ( .A(b[7]), .B(a[7]), .ZN(n344) );
  NAND2_X1 U357 ( .A1(n334), .A2(n353), .ZN(n336) );
  XNOR2_X1 U358 ( .A(n298), .B(a[6]), .ZN(n353) );
  XNOR2_X1 U359 ( .A(b[6]), .B(a[7]), .ZN(n342) );
  OAI22_X1 U360 ( .A1(n274), .A2(n309), .B1(n354), .B2(n307), .ZN(n104) );
  OAI22_X1 U361 ( .A1(n260), .A2(n309), .B1(n355), .B2(n307), .ZN(n103) );
  XNOR2_X1 U362 ( .A(b[1]), .B(a[1]), .ZN(n354) );
  OAI22_X1 U363 ( .A1(n355), .A2(n309), .B1(n356), .B2(n307), .ZN(n102) );
  XNOR2_X1 U364 ( .A(b[2]), .B(a[1]), .ZN(n355) );
  OAI22_X1 U365 ( .A1(n356), .A2(n309), .B1(n357), .B2(n307), .ZN(n101) );
  XNOR2_X1 U366 ( .A(b[3]), .B(a[1]), .ZN(n356) );
  OAI22_X1 U367 ( .A1(n357), .A2(n309), .B1(n308), .B2(n307), .ZN(n100) );
  XNOR2_X1 U368 ( .A(b[5]), .B(a[1]), .ZN(n308) );
  NAND2_X1 U369 ( .A1(a[1]), .A2(n307), .ZN(n309) );
  XNOR2_X1 U370 ( .A(b[4]), .B(a[1]), .ZN(n357) );
endmodule


module mac_18 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  mac_18_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_18_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_17_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66;
  wire   [15:1] carry;

  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n66), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(carry[9]), .Z(n1) );
  XNOR2_X1 U2 ( .A(B[15]), .B(A[15]), .ZN(n2) );
  NAND3_X1 U3 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n3) );
  NAND3_X1 U4 ( .A1(n20), .A2(n21), .A3(n22), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(carry[10]), .Z(n5) );
  NAND3_X1 U6 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n6) );
  NAND3_X1 U7 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n7) );
  CLKBUF_X1 U8 ( .A(n4), .Z(n8) );
  CLKBUF_X1 U9 ( .A(n3), .Z(n9) );
  XOR2_X1 U10 ( .A(B[8]), .B(A[8]), .Z(n10) );
  XOR2_X1 U11 ( .A(carry[8]), .B(n10), .Z(SUM[8]) );
  NAND2_X1 U12 ( .A1(carry[8]), .A2(B[8]), .ZN(n11) );
  NAND2_X1 U13 ( .A1(carry[8]), .A2(A[8]), .ZN(n12) );
  NAND2_X1 U14 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND3_X1 U15 ( .A1(n11), .A2(n12), .A3(n13), .ZN(carry[9]) );
  CLKBUF_X1 U16 ( .A(n49), .Z(n14) );
  XOR2_X1 U17 ( .A(B[9]), .B(A[9]), .Z(n15) );
  XOR2_X1 U18 ( .A(n1), .B(n15), .Z(SUM[9]) );
  NAND2_X1 U19 ( .A1(carry[9]), .A2(B[9]), .ZN(n16) );
  NAND2_X1 U20 ( .A1(carry[9]), .A2(A[9]), .ZN(n17) );
  NAND2_X1 U21 ( .A1(B[9]), .A2(A[9]), .ZN(n18) );
  NAND3_X1 U22 ( .A1(n16), .A2(n17), .A3(n18), .ZN(carry[10]) );
  XOR2_X1 U23 ( .A(B[10]), .B(A[10]), .Z(n19) );
  XOR2_X1 U24 ( .A(n5), .B(n19), .Z(SUM[10]) );
  NAND2_X1 U25 ( .A1(carry[10]), .A2(B[10]), .ZN(n20) );
  NAND2_X1 U26 ( .A1(carry[10]), .A2(A[10]), .ZN(n21) );
  NAND2_X1 U27 ( .A1(B[10]), .A2(A[10]), .ZN(n22) );
  NAND3_X1 U28 ( .A1(n20), .A2(n21), .A3(n22), .ZN(carry[11]) );
  XOR2_X1 U29 ( .A(B[3]), .B(A[3]), .Z(n23) );
  XOR2_X1 U30 ( .A(carry[3]), .B(n23), .Z(SUM[3]) );
  NAND2_X1 U31 ( .A1(carry[3]), .A2(B[3]), .ZN(n24) );
  NAND2_X1 U32 ( .A1(carry[3]), .A2(A[3]), .ZN(n25) );
  NAND2_X1 U33 ( .A1(B[3]), .A2(A[3]), .ZN(n26) );
  NAND3_X1 U34 ( .A1(n24), .A2(n25), .A3(n26), .ZN(carry[4]) );
  NAND3_X1 U35 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n27) );
  NAND3_X1 U36 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n28) );
  XOR2_X1 U37 ( .A(B[11]), .B(A[11]), .Z(n29) );
  XOR2_X1 U38 ( .A(n8), .B(n29), .Z(SUM[11]) );
  NAND2_X1 U39 ( .A1(n4), .A2(B[11]), .ZN(n30) );
  NAND2_X1 U40 ( .A1(carry[11]), .A2(A[11]), .ZN(n31) );
  NAND2_X1 U41 ( .A1(B[11]), .A2(A[11]), .ZN(n32) );
  XOR2_X1 U42 ( .A(B[4]), .B(A[4]), .Z(n33) );
  XOR2_X1 U43 ( .A(n7), .B(n33), .Z(SUM[4]) );
  NAND2_X1 U44 ( .A1(n6), .A2(B[4]), .ZN(n34) );
  NAND2_X1 U45 ( .A1(carry[4]), .A2(A[4]), .ZN(n35) );
  NAND2_X1 U46 ( .A1(B[4]), .A2(A[4]), .ZN(n36) );
  NAND3_X1 U47 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[5]) );
  NAND3_X1 U48 ( .A1(n40), .A2(n41), .A3(n42), .ZN(n37) );
  NAND3_X1 U49 ( .A1(n44), .A2(n45), .A3(n46), .ZN(n38) );
  XOR2_X1 U50 ( .A(B[12]), .B(A[12]), .Z(n39) );
  XOR2_X1 U51 ( .A(n9), .B(n39), .Z(SUM[12]) );
  NAND2_X1 U52 ( .A1(n3), .A2(B[12]), .ZN(n40) );
  NAND2_X1 U53 ( .A1(n27), .A2(A[12]), .ZN(n41) );
  NAND2_X1 U54 ( .A1(B[12]), .A2(A[12]), .ZN(n42) );
  NAND3_X1 U55 ( .A1(n40), .A2(n41), .A3(n42), .ZN(carry[13]) );
  XOR2_X1 U56 ( .A(B[5]), .B(A[5]), .Z(n43) );
  XOR2_X1 U57 ( .A(n28), .B(n43), .Z(SUM[5]) );
  NAND2_X1 U58 ( .A1(n28), .A2(B[5]), .ZN(n44) );
  NAND2_X1 U59 ( .A1(carry[5]), .A2(A[5]), .ZN(n45) );
  NAND2_X1 U60 ( .A1(B[5]), .A2(A[5]), .ZN(n46) );
  NAND3_X1 U61 ( .A1(n44), .A2(n45), .A3(n46), .ZN(carry[6]) );
  XNOR2_X1 U62 ( .A(carry[15]), .B(n2), .ZN(SUM[15]) );
  NAND3_X1 U63 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n47) );
  NAND3_X1 U64 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n48) );
  NAND3_X1 U65 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n49) );
  XOR2_X1 U66 ( .A(B[13]), .B(A[13]), .Z(n50) );
  XOR2_X1 U67 ( .A(carry[13]), .B(n50), .Z(SUM[13]) );
  NAND2_X1 U68 ( .A1(n37), .A2(B[13]), .ZN(n51) );
  NAND2_X1 U69 ( .A1(carry[13]), .A2(A[13]), .ZN(n52) );
  NAND2_X1 U70 ( .A1(B[13]), .A2(A[13]), .ZN(n53) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(n54) );
  XOR2_X1 U72 ( .A(carry[6]), .B(n54), .Z(SUM[6]) );
  NAND2_X1 U73 ( .A1(n38), .A2(B[6]), .ZN(n55) );
  NAND2_X1 U74 ( .A1(carry[6]), .A2(A[6]), .ZN(n56) );
  NAND2_X1 U75 ( .A1(B[6]), .A2(A[6]), .ZN(n57) );
  NAND3_X1 U76 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[7]) );
  XOR2_X1 U77 ( .A(B[14]), .B(A[14]), .Z(n58) );
  XOR2_X1 U78 ( .A(n48), .B(n58), .Z(SUM[14]) );
  NAND2_X1 U79 ( .A1(n47), .A2(B[14]), .ZN(n59) );
  NAND2_X1 U80 ( .A1(n47), .A2(A[14]), .ZN(n60) );
  NAND2_X1 U81 ( .A1(B[14]), .A2(A[14]), .ZN(n61) );
  NAND3_X1 U82 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[15]) );
  XOR2_X1 U83 ( .A(B[7]), .B(A[7]), .Z(n62) );
  XOR2_X1 U84 ( .A(n14), .B(n62), .Z(SUM[7]) );
  NAND2_X1 U85 ( .A1(n49), .A2(B[7]), .ZN(n63) );
  NAND2_X1 U86 ( .A1(carry[7]), .A2(A[7]), .ZN(n64) );
  NAND2_X1 U87 ( .A1(B[7]), .A2(A[7]), .ZN(n65) );
  NAND3_X1 U88 ( .A1(n63), .A2(n64), .A3(n65), .ZN(carry[8]) );
  AND2_X1 U89 ( .A1(B[0]), .A2(A[0]), .ZN(n66) );
  XOR2_X1 U90 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_17_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n313), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n312), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n316), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n315), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n318), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  BUF_X1 U157 ( .A(n326), .Z(n284) );
  NAND2_X1 U158 ( .A1(n336), .A2(n365), .ZN(n338) );
  NAND2_X1 U159 ( .A1(n4), .A2(n19), .ZN(n206) );
  AND2_X1 U160 ( .A1(n95), .A2(n102), .ZN(n207) );
  NAND2_X2 U161 ( .A1(n233), .A2(n234), .ZN(n208) );
  INV_X1 U162 ( .A(n317), .ZN(n209) );
  NAND2_X1 U163 ( .A1(n233), .A2(n234), .ZN(n336) );
  NAND2_X1 U164 ( .A1(n223), .A2(n34), .ZN(n210) );
  CLKBUF_X1 U165 ( .A(b[1]), .Z(n211) );
  INV_X1 U166 ( .A(n308), .ZN(n212) );
  INV_X1 U167 ( .A(n308), .ZN(n213) );
  INV_X1 U168 ( .A(n308), .ZN(n307) );
  NAND2_X2 U169 ( .A1(n326), .A2(n364), .ZN(n328) );
  XNOR2_X1 U170 ( .A(n211), .B(n298), .ZN(n214) );
  CLKBUF_X3 U171 ( .A(a[1]), .Z(n298) );
  XNOR2_X1 U172 ( .A(a[6]), .B(a[5]), .ZN(n347) );
  XNOR2_X1 U173 ( .A(a[6]), .B(a[5]), .ZN(n215) );
  CLKBUF_X1 U174 ( .A(n223), .Z(n216) );
  NAND3_X1 U175 ( .A1(n297), .A2(n296), .A3(n295), .ZN(n217) );
  CLKBUF_X1 U176 ( .A(n293), .Z(n218) );
  NAND3_X1 U177 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n219) );
  CLKBUF_X1 U178 ( .A(n306), .Z(n220) );
  CLKBUF_X1 U179 ( .A(n210), .Z(n221) );
  XNOR2_X1 U180 ( .A(n222), .B(n42), .ZN(n40) );
  XNOR2_X1 U181 ( .A(n47), .B(n44), .ZN(n222) );
  NAND3_X1 U182 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n223) );
  CLKBUF_X1 U183 ( .A(n219), .Z(n224) );
  XOR2_X1 U184 ( .A(n45), .B(n224), .Z(n225) );
  XOR2_X1 U185 ( .A(n225), .B(n40), .Z(product[7]) );
  NAND2_X1 U186 ( .A1(n47), .A2(n44), .ZN(n226) );
  NAND2_X1 U187 ( .A1(n47), .A2(n42), .ZN(n227) );
  NAND2_X1 U188 ( .A1(n44), .A2(n42), .ZN(n228) );
  NAND3_X1 U189 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n39) );
  NAND2_X1 U190 ( .A1(n219), .A2(n45), .ZN(n229) );
  NAND2_X1 U191 ( .A1(n45), .A2(n40), .ZN(n230) );
  NAND2_X1 U192 ( .A1(n9), .A2(n40), .ZN(n231) );
  NAND3_X1 U193 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n8) );
  NAND2_X1 U194 ( .A1(a[4]), .A2(a[3]), .ZN(n233) );
  NAND2_X1 U195 ( .A1(n232), .A2(n317), .ZN(n234) );
  INV_X1 U196 ( .A(a[4]), .ZN(n232) );
  CLKBUF_X1 U197 ( .A(n4), .Z(n235) );
  CLKBUF_X1 U198 ( .A(n257), .Z(n236) );
  NAND3_X1 U199 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n237) );
  NAND3_X1 U200 ( .A1(n221), .A2(n243), .A3(n244), .ZN(n238) );
  CLKBUF_X1 U201 ( .A(n206), .Z(n239) );
  NAND3_X1 U202 ( .A1(n277), .A2(n278), .A3(n279), .ZN(n240) );
  XOR2_X1 U203 ( .A(n34), .B(n39), .Z(n241) );
  XOR2_X1 U204 ( .A(n216), .B(n241), .Z(product[8]) );
  NAND2_X1 U205 ( .A1(n223), .A2(n34), .ZN(n242) );
  NAND2_X1 U206 ( .A1(n8), .A2(n39), .ZN(n243) );
  NAND2_X1 U207 ( .A1(n34), .A2(n39), .ZN(n244) );
  NAND3_X1 U208 ( .A1(n210), .A2(n243), .A3(n244), .ZN(n7) );
  NAND3_X1 U209 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n245) );
  NAND3_X1 U210 ( .A1(n256), .A2(n236), .A3(n258), .ZN(n246) );
  NAND3_X1 U211 ( .A1(n306), .A2(n305), .A3(n304), .ZN(n247) );
  NAND3_X1 U212 ( .A1(n304), .A2(n305), .A3(n220), .ZN(n248) );
  XOR2_X1 U213 ( .A(n46), .B(n49), .Z(n249) );
  XOR2_X1 U214 ( .A(n248), .B(n249), .Z(product[6]) );
  NAND2_X1 U215 ( .A1(n247), .A2(n46), .ZN(n250) );
  NAND2_X1 U216 ( .A1(n10), .A2(n49), .ZN(n251) );
  NAND2_X1 U217 ( .A1(n46), .A2(n49), .ZN(n252) );
  NAND3_X1 U218 ( .A1(n251), .A2(n250), .A3(n252), .ZN(n9) );
  CLKBUF_X1 U219 ( .A(n259), .Z(n253) );
  CLKBUF_X1 U220 ( .A(n275), .Z(n254) );
  XOR2_X1 U221 ( .A(n103), .B(n96), .Z(n255) );
  XOR2_X1 U222 ( .A(n14), .B(n255), .Z(product[2]) );
  NAND2_X1 U223 ( .A1(n14), .A2(n103), .ZN(n256) );
  NAND2_X1 U224 ( .A1(n14), .A2(n96), .ZN(n257) );
  NAND2_X1 U225 ( .A1(n103), .A2(n96), .ZN(n258) );
  NAND3_X1 U226 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n13) );
  NAND3_X1 U227 ( .A1(n262), .A2(n261), .A3(n263), .ZN(n259) );
  XOR2_X1 U228 ( .A(n33), .B(n28), .Z(n260) );
  XOR2_X1 U229 ( .A(n238), .B(n260), .Z(product[9]) );
  NAND2_X1 U230 ( .A1(n237), .A2(n33), .ZN(n261) );
  NAND2_X1 U231 ( .A1(n7), .A2(n28), .ZN(n262) );
  NAND2_X1 U232 ( .A1(n33), .A2(n28), .ZN(n263) );
  NAND3_X1 U233 ( .A1(n262), .A2(n261), .A3(n263), .ZN(n6) );
  CLKBUF_X1 U234 ( .A(n240), .Z(n264) );
  NAND3_X1 U235 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n265) );
  NAND3_X1 U236 ( .A1(n273), .A2(n275), .A3(n274), .ZN(n266) );
  NAND3_X1 U237 ( .A1(n273), .A2(n274), .A3(n254), .ZN(n267) );
  XOR2_X1 U238 ( .A(n20), .B(n23), .Z(n268) );
  XOR2_X1 U239 ( .A(n264), .B(n268), .Z(product[11]) );
  NAND2_X1 U240 ( .A1(n240), .A2(n20), .ZN(n269) );
  NAND2_X1 U241 ( .A1(n5), .A2(n23), .ZN(n270) );
  NAND2_X1 U242 ( .A1(n20), .A2(n23), .ZN(n271) );
  NAND3_X1 U243 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n4) );
  XOR2_X1 U244 ( .A(n246), .B(n71), .Z(n272) );
  XOR2_X1 U245 ( .A(n56), .B(n272), .Z(product[3]) );
  NAND2_X1 U246 ( .A1(n245), .A2(n56), .ZN(n273) );
  NAND2_X1 U247 ( .A1(n56), .A2(n71), .ZN(n274) );
  NAND2_X1 U248 ( .A1(n13), .A2(n71), .ZN(n275) );
  NAND3_X1 U249 ( .A1(n273), .A2(n275), .A3(n274), .ZN(n12) );
  XOR2_X1 U250 ( .A(n27), .B(n24), .Z(n276) );
  XOR2_X1 U251 ( .A(n253), .B(n276), .Z(product[10]) );
  NAND2_X1 U252 ( .A1(n259), .A2(n27), .ZN(n277) );
  NAND2_X1 U253 ( .A1(n6), .A2(n24), .ZN(n278) );
  NAND2_X1 U254 ( .A1(n27), .A2(n24), .ZN(n279) );
  NAND3_X1 U255 ( .A1(n277), .A2(n278), .A3(n279), .ZN(n5) );
  NAND3_X1 U256 ( .A1(n300), .A2(n301), .A3(n302), .ZN(n280) );
  INV_X1 U257 ( .A(n212), .ZN(n281) );
  NAND3_X1 U258 ( .A1(n292), .A2(n291), .A3(n293), .ZN(n282) );
  NAND3_X1 U259 ( .A1(n291), .A2(n239), .A3(n218), .ZN(n283) );
  XOR2_X1 U260 ( .A(n95), .B(n102), .Z(n56) );
  XNOR2_X1 U261 ( .A(n217), .B(n285), .ZN(product[14]) );
  XNOR2_X1 U262 ( .A(n310), .B(n15), .ZN(n285) );
  INV_X1 U263 ( .A(n15), .ZN(n309) );
  AND3_X1 U264 ( .A1(n287), .A2(n288), .A3(n289), .ZN(product[15]) );
  INV_X1 U265 ( .A(n334), .ZN(n316) );
  INV_X1 U266 ( .A(n345), .ZN(n313) );
  INV_X1 U267 ( .A(n21), .ZN(n312) );
  INV_X1 U268 ( .A(n325), .ZN(n318) );
  INV_X1 U269 ( .A(n31), .ZN(n315) );
  INV_X1 U270 ( .A(b[0]), .ZN(n308) );
  XOR2_X1 U271 ( .A(a[2]), .B(n319), .Z(n326) );
  INV_X1 U272 ( .A(a[0]), .ZN(n320) );
  INV_X1 U273 ( .A(a[3]), .ZN(n317) );
  INV_X1 U274 ( .A(a[5]), .ZN(n314) );
  INV_X1 U275 ( .A(a[7]), .ZN(n311) );
  NAND2_X1 U276 ( .A1(n217), .A2(n310), .ZN(n287) );
  NAND2_X1 U277 ( .A1(n2), .A2(n15), .ZN(n288) );
  NAND2_X1 U278 ( .A1(n310), .A2(n15), .ZN(n289) );
  XOR2_X1 U279 ( .A(n19), .B(n18), .Z(n290) );
  XOR2_X1 U280 ( .A(n290), .B(n235), .Z(product[12]) );
  NAND2_X1 U281 ( .A1(n19), .A2(n18), .ZN(n291) );
  NAND2_X1 U282 ( .A1(n4), .A2(n19), .ZN(n292) );
  NAND2_X1 U283 ( .A1(n18), .A2(n265), .ZN(n293) );
  NAND3_X1 U284 ( .A1(n206), .A2(n293), .A3(n291), .ZN(n3) );
  XOR2_X1 U285 ( .A(n17), .B(n309), .Z(n294) );
  XOR2_X1 U286 ( .A(n294), .B(n283), .Z(product[13]) );
  NAND2_X1 U287 ( .A1(n17), .A2(n309), .ZN(n295) );
  NAND2_X1 U288 ( .A1(n17), .A2(n282), .ZN(n296) );
  NAND2_X1 U289 ( .A1(n309), .A2(n3), .ZN(n297) );
  NAND3_X1 U290 ( .A1(n297), .A2(n295), .A3(n296), .ZN(n2) );
  INV_X1 U291 ( .A(n356), .ZN(n310) );
  XOR2_X1 U292 ( .A(n54), .B(n207), .Z(n299) );
  XOR2_X1 U293 ( .A(n299), .B(n267), .Z(product[4]) );
  NAND2_X1 U294 ( .A1(n54), .A2(n207), .ZN(n300) );
  NAND2_X1 U295 ( .A1(n54), .A2(n266), .ZN(n301) );
  NAND2_X1 U296 ( .A1(n207), .A2(n12), .ZN(n302) );
  NAND3_X1 U297 ( .A1(n300), .A2(n301), .A3(n302), .ZN(n11) );
  XOR2_X1 U298 ( .A(n50), .B(n53), .Z(n303) );
  XOR2_X1 U299 ( .A(n303), .B(n11), .Z(product[5]) );
  NAND2_X1 U300 ( .A1(n50), .A2(n53), .ZN(n304) );
  NAND2_X1 U301 ( .A1(n50), .A2(n280), .ZN(n305) );
  NAND2_X1 U302 ( .A1(n53), .A2(n11), .ZN(n306) );
  NAND3_X1 U303 ( .A1(n306), .A2(n305), .A3(n304), .ZN(n10) );
  INV_X1 U304 ( .A(a[1]), .ZN(n319) );
  NOR2_X1 U305 ( .A1(n320), .A2(n281), .ZN(product[0]) );
  OAI22_X1 U306 ( .A1(n321), .A2(n322), .B1(n323), .B2(n320), .ZN(n99) );
  OAI22_X1 U307 ( .A1(n323), .A2(n322), .B1(n324), .B2(n320), .ZN(n98) );
  XNOR2_X1 U308 ( .A(b[6]), .B(n298), .ZN(n323) );
  OAI22_X1 U309 ( .A1(n320), .A2(n324), .B1(n322), .B2(n324), .ZN(n325) );
  XNOR2_X1 U310 ( .A(b[7]), .B(n298), .ZN(n324) );
  NOR2_X1 U311 ( .A1(n326), .A2(n308), .ZN(n96) );
  OAI22_X1 U312 ( .A1(n327), .A2(n328), .B1(n326), .B2(n329), .ZN(n95) );
  XNOR2_X1 U313 ( .A(a[3]), .B(n307), .ZN(n327) );
  OAI22_X1 U314 ( .A1(n329), .A2(n328), .B1(n284), .B2(n330), .ZN(n94) );
  XNOR2_X1 U315 ( .A(b[1]), .B(a[3]), .ZN(n329) );
  OAI22_X1 U316 ( .A1(n330), .A2(n328), .B1(n284), .B2(n331), .ZN(n93) );
  XNOR2_X1 U317 ( .A(b[2]), .B(a[3]), .ZN(n330) );
  OAI22_X1 U318 ( .A1(n331), .A2(n328), .B1(n284), .B2(n332), .ZN(n92) );
  XNOR2_X1 U319 ( .A(b[3]), .B(n209), .ZN(n331) );
  OAI22_X1 U320 ( .A1(n332), .A2(n328), .B1(n284), .B2(n333), .ZN(n91) );
  XNOR2_X1 U321 ( .A(b[4]), .B(a[3]), .ZN(n332) );
  OAI22_X1 U322 ( .A1(n335), .A2(n284), .B1(n328), .B2(n335), .ZN(n334) );
  NOR2_X1 U323 ( .A1(n208), .A2(n281), .ZN(n88) );
  OAI22_X1 U324 ( .A1(n337), .A2(n338), .B1(n208), .B2(n339), .ZN(n87) );
  XNOR2_X1 U325 ( .A(a[5]), .B(n213), .ZN(n337) );
  OAI22_X1 U326 ( .A1(n339), .A2(n338), .B1(n208), .B2(n340), .ZN(n86) );
  XNOR2_X1 U327 ( .A(n211), .B(a[5]), .ZN(n339) );
  OAI22_X1 U328 ( .A1(n340), .A2(n338), .B1(n208), .B2(n341), .ZN(n85) );
  XNOR2_X1 U329 ( .A(b[2]), .B(a[5]), .ZN(n340) );
  OAI22_X1 U330 ( .A1(n341), .A2(n338), .B1(n208), .B2(n342), .ZN(n84) );
  XNOR2_X1 U331 ( .A(b[3]), .B(a[5]), .ZN(n341) );
  OAI22_X1 U332 ( .A1(n342), .A2(n338), .B1(n208), .B2(n343), .ZN(n83) );
  XNOR2_X1 U333 ( .A(b[4]), .B(a[5]), .ZN(n342) );
  OAI22_X1 U334 ( .A1(n343), .A2(n338), .B1(n208), .B2(n344), .ZN(n82) );
  XNOR2_X1 U335 ( .A(b[5]), .B(a[5]), .ZN(n343) );
  OAI22_X1 U336 ( .A1(n346), .A2(n208), .B1(n338), .B2(n346), .ZN(n345) );
  NOR2_X1 U337 ( .A1(n347), .A2(n281), .ZN(n80) );
  OAI22_X1 U338 ( .A1(n348), .A2(n349), .B1(n215), .B2(n350), .ZN(n79) );
  XNOR2_X1 U339 ( .A(a[7]), .B(n212), .ZN(n348) );
  OAI22_X1 U340 ( .A1(n351), .A2(n349), .B1(n215), .B2(n352), .ZN(n77) );
  OAI22_X1 U341 ( .A1(n352), .A2(n349), .B1(n215), .B2(n353), .ZN(n76) );
  XNOR2_X1 U342 ( .A(b[3]), .B(a[7]), .ZN(n352) );
  OAI22_X1 U343 ( .A1(n353), .A2(n349), .B1(n215), .B2(n354), .ZN(n75) );
  XNOR2_X1 U344 ( .A(b[4]), .B(a[7]), .ZN(n353) );
  OAI22_X1 U345 ( .A1(n354), .A2(n349), .B1(n215), .B2(n355), .ZN(n74) );
  XNOR2_X1 U346 ( .A(b[5]), .B(a[7]), .ZN(n354) );
  OAI22_X1 U347 ( .A1(n357), .A2(n215), .B1(n349), .B2(n357), .ZN(n356) );
  OAI21_X1 U348 ( .B1(n212), .B2(n319), .A(n322), .ZN(n72) );
  OAI21_X1 U349 ( .B1(n317), .B2(n328), .A(n358), .ZN(n71) );
  OR3_X1 U350 ( .A1(n284), .A2(n213), .A3(n317), .ZN(n358) );
  OAI21_X1 U351 ( .B1(n314), .B2(n338), .A(n359), .ZN(n70) );
  OR3_X1 U352 ( .A1(n336), .A2(n307), .A3(n314), .ZN(n359) );
  OAI21_X1 U353 ( .B1(n311), .B2(n349), .A(n360), .ZN(n69) );
  OR3_X1 U354 ( .A1(n215), .A2(n213), .A3(n311), .ZN(n360) );
  XNOR2_X1 U355 ( .A(n361), .B(n362), .ZN(n38) );
  OR2_X1 U356 ( .A1(n361), .A2(n362), .ZN(n37) );
  OAI22_X1 U357 ( .A1(n333), .A2(n328), .B1(n284), .B2(n363), .ZN(n362) );
  XNOR2_X1 U358 ( .A(b[5]), .B(n209), .ZN(n333) );
  OAI22_X1 U359 ( .A1(n350), .A2(n349), .B1(n215), .B2(n351), .ZN(n361) );
  XNOR2_X1 U360 ( .A(b[2]), .B(a[7]), .ZN(n351) );
  XNOR2_X1 U361 ( .A(b[1]), .B(a[7]), .ZN(n350) );
  OAI22_X1 U362 ( .A1(n363), .A2(n328), .B1(n284), .B2(n335), .ZN(n31) );
  XNOR2_X1 U363 ( .A(b[7]), .B(n209), .ZN(n335) );
  XNOR2_X1 U364 ( .A(n317), .B(a[2]), .ZN(n364) );
  XNOR2_X1 U365 ( .A(b[6]), .B(n209), .ZN(n363) );
  OAI22_X1 U366 ( .A1(n344), .A2(n338), .B1(n208), .B2(n346), .ZN(n21) );
  XNOR2_X1 U367 ( .A(b[7]), .B(a[5]), .ZN(n346) );
  XNOR2_X1 U368 ( .A(n314), .B(a[4]), .ZN(n365) );
  XNOR2_X1 U369 ( .A(b[6]), .B(a[5]), .ZN(n344) );
  OAI22_X1 U370 ( .A1(n355), .A2(n349), .B1(n215), .B2(n357), .ZN(n15) );
  XNOR2_X1 U371 ( .A(b[7]), .B(a[7]), .ZN(n357) );
  NAND2_X1 U372 ( .A1(n347), .A2(n366), .ZN(n349) );
  XNOR2_X1 U373 ( .A(n311), .B(a[6]), .ZN(n366) );
  XNOR2_X1 U374 ( .A(b[6]), .B(a[7]), .ZN(n355) );
  OAI22_X1 U375 ( .A1(n213), .A2(n322), .B1(n367), .B2(n320), .ZN(n104) );
  OAI22_X1 U376 ( .A1(n214), .A2(n322), .B1(n368), .B2(n320), .ZN(n103) );
  XNOR2_X1 U377 ( .A(b[1]), .B(n298), .ZN(n367) );
  OAI22_X1 U378 ( .A1(n368), .A2(n322), .B1(n369), .B2(n320), .ZN(n102) );
  XNOR2_X1 U379 ( .A(b[2]), .B(n298), .ZN(n368) );
  OAI22_X1 U380 ( .A1(n369), .A2(n322), .B1(n370), .B2(n320), .ZN(n101) );
  XNOR2_X1 U381 ( .A(b[3]), .B(n298), .ZN(n369) );
  OAI22_X1 U382 ( .A1(n370), .A2(n322), .B1(n321), .B2(n320), .ZN(n100) );
  XNOR2_X1 U383 ( .A(b[5]), .B(n298), .ZN(n321) );
  NAND2_X1 U384 ( .A1(a[1]), .A2(n320), .ZN(n322) );
  XNOR2_X1 U385 ( .A(b[4]), .B(n298), .ZN(n370) );
endmodule


module mac_17 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_17_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_17_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_16_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88;
  wire   [15:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .S(SUM[15]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n88) );
  CLKBUF_X1 U2 ( .A(n38), .Z(n1) );
  NAND2_X1 U3 ( .A1(n51), .A2(B[10]), .ZN(n2) );
  NAND3_X1 U4 ( .A1(n85), .A2(n86), .A3(n87), .ZN(n3) );
  NAND3_X1 U5 ( .A1(n85), .A2(n86), .A3(n87), .ZN(n4) );
  NAND3_X1 U6 ( .A1(n9), .A2(n10), .A3(n11), .ZN(n5) );
  NAND3_X1 U7 ( .A1(n9), .A2(n10), .A3(n11), .ZN(n6) );
  CLKBUF_X1 U8 ( .A(n82), .Z(n7) );
  XOR2_X1 U9 ( .A(B[3]), .B(A[3]), .Z(n8) );
  XOR2_X1 U10 ( .A(n4), .B(n8), .Z(SUM[3]) );
  NAND2_X1 U11 ( .A1(n3), .A2(B[3]), .ZN(n9) );
  NAND2_X1 U12 ( .A1(carry[3]), .A2(A[3]), .ZN(n10) );
  NAND2_X1 U13 ( .A1(B[3]), .A2(A[3]), .ZN(n11) );
  NAND3_X1 U14 ( .A1(n9), .A2(n10), .A3(n11), .ZN(carry[4]) );
  CLKBUF_X1 U15 ( .A(n55), .Z(n12) );
  NAND3_X1 U16 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n13) );
  NAND3_X1 U17 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n14) );
  NAND3_X1 U18 ( .A1(n37), .A2(n1), .A3(n39), .ZN(n15) );
  NAND3_X1 U19 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n16) );
  NAND3_X1 U20 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n17) );
  NAND3_X1 U21 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n18) );
  NAND3_X1 U22 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n19) );
  NAND3_X1 U23 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n20) );
  XOR2_X1 U24 ( .A(B[5]), .B(A[5]), .Z(n21) );
  XOR2_X1 U25 ( .A(n17), .B(n21), .Z(SUM[5]) );
  NAND2_X1 U26 ( .A1(n16), .A2(B[5]), .ZN(n22) );
  NAND2_X1 U27 ( .A1(carry[5]), .A2(A[5]), .ZN(n23) );
  NAND2_X1 U28 ( .A1(B[5]), .A2(A[5]), .ZN(n24) );
  NAND3_X1 U29 ( .A1(n22), .A2(n23), .A3(n24), .ZN(carry[6]) );
  CLKBUF_X1 U30 ( .A(n13), .Z(n25) );
  NAND3_X1 U31 ( .A1(n2), .A2(n55), .A3(n56), .ZN(n26) );
  NAND3_X1 U32 ( .A1(n2), .A2(n12), .A3(n56), .ZN(n27) );
  XOR2_X1 U33 ( .A(B[4]), .B(A[4]), .Z(n28) );
  XOR2_X1 U34 ( .A(n6), .B(n28), .Z(SUM[4]) );
  NAND2_X1 U35 ( .A1(n5), .A2(B[4]), .ZN(n29) );
  NAND2_X1 U36 ( .A1(carry[4]), .A2(A[4]), .ZN(n30) );
  NAND2_X1 U37 ( .A1(B[4]), .A2(A[4]), .ZN(n31) );
  NAND3_X1 U38 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[5]) );
  CLKBUF_X1 U39 ( .A(n63), .Z(n32) );
  CLKBUF_X1 U40 ( .A(n44), .Z(n33) );
  CLKBUF_X1 U41 ( .A(n78), .Z(n34) );
  NAND3_X1 U42 ( .A1(n74), .A2(n73), .A3(n75), .ZN(n35) );
  XOR2_X1 U43 ( .A(B[6]), .B(A[6]), .Z(n36) );
  XOR2_X1 U44 ( .A(n19), .B(n36), .Z(SUM[6]) );
  NAND2_X1 U45 ( .A1(n18), .A2(B[6]), .ZN(n37) );
  NAND2_X1 U46 ( .A1(carry[6]), .A2(A[6]), .ZN(n38) );
  NAND2_X1 U47 ( .A1(B[6]), .A2(A[6]), .ZN(n39) );
  NAND3_X1 U48 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[7]) );
  XOR2_X1 U49 ( .A(B[11]), .B(A[11]), .Z(n40) );
  XOR2_X1 U50 ( .A(n27), .B(n40), .Z(SUM[11]) );
  NAND2_X1 U51 ( .A1(n26), .A2(B[11]), .ZN(n41) );
  NAND2_X1 U52 ( .A1(carry[11]), .A2(A[11]), .ZN(n42) );
  NAND2_X1 U53 ( .A1(B[11]), .A2(A[11]), .ZN(n43) );
  NAND3_X1 U54 ( .A1(n41), .A2(n42), .A3(n43), .ZN(carry[12]) );
  NAND3_X1 U55 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n44) );
  XOR2_X1 U56 ( .A(B[12]), .B(A[12]), .Z(n45) );
  XOR2_X1 U57 ( .A(n25), .B(n45), .Z(SUM[12]) );
  NAND2_X1 U58 ( .A1(n13), .A2(B[12]), .ZN(n46) );
  NAND2_X1 U59 ( .A1(carry[12]), .A2(A[12]), .ZN(n47) );
  NAND2_X1 U60 ( .A1(B[12]), .A2(A[12]), .ZN(n48) );
  NAND3_X1 U61 ( .A1(n47), .A2(n46), .A3(n48), .ZN(carry[13]) );
  CLKBUF_X1 U62 ( .A(n20), .Z(n49) );
  NAND3_X1 U63 ( .A1(n62), .A2(n32), .A3(n64), .ZN(n50) );
  NAND3_X1 U64 ( .A1(n78), .A2(n77), .A3(n79), .ZN(n51) );
  NAND3_X1 U65 ( .A1(n77), .A2(n34), .A3(n79), .ZN(n52) );
  XOR2_X1 U66 ( .A(B[10]), .B(A[10]), .Z(n53) );
  XOR2_X1 U67 ( .A(n52), .B(n53), .Z(SUM[10]) );
  NAND2_X1 U68 ( .A1(n51), .A2(B[10]), .ZN(n54) );
  NAND2_X1 U69 ( .A1(carry[10]), .A2(A[10]), .ZN(n55) );
  NAND2_X1 U70 ( .A1(B[10]), .A2(A[10]), .ZN(n56) );
  NAND3_X1 U71 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[11]) );
  XOR2_X1 U72 ( .A(B[13]), .B(A[13]), .Z(n57) );
  XOR2_X1 U73 ( .A(n33), .B(n57), .Z(SUM[13]) );
  NAND2_X1 U74 ( .A1(n44), .A2(B[13]), .ZN(n58) );
  NAND2_X1 U75 ( .A1(carry[13]), .A2(A[13]), .ZN(n59) );
  NAND2_X1 U76 ( .A1(B[13]), .A2(A[13]), .ZN(n60) );
  NAND3_X1 U77 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[14]) );
  XOR2_X1 U78 ( .A(B[7]), .B(A[7]), .Z(n61) );
  XOR2_X1 U79 ( .A(n15), .B(n61), .Z(SUM[7]) );
  NAND2_X1 U80 ( .A1(n14), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U81 ( .A1(carry[7]), .A2(A[7]), .ZN(n63) );
  NAND2_X1 U82 ( .A1(B[7]), .A2(A[7]), .ZN(n64) );
  NAND3_X1 U83 ( .A1(n62), .A2(n63), .A3(n64), .ZN(carry[8]) );
  NAND3_X1 U84 ( .A1(n81), .A2(n82), .A3(n83), .ZN(n65) );
  NAND3_X1 U85 ( .A1(n81), .A2(n7), .A3(n83), .ZN(n66) );
  XOR2_X1 U86 ( .A(B[14]), .B(A[14]), .Z(n67) );
  XOR2_X1 U87 ( .A(n49), .B(n67), .Z(SUM[14]) );
  NAND2_X1 U88 ( .A1(n20), .A2(B[14]), .ZN(n68) );
  NAND2_X1 U89 ( .A1(carry[14]), .A2(A[14]), .ZN(n69) );
  NAND2_X1 U90 ( .A1(B[14]), .A2(A[14]), .ZN(n70) );
  NAND3_X1 U91 ( .A1(n68), .A2(n69), .A3(n70), .ZN(carry[15]) );
  CLKBUF_X1 U92 ( .A(carry[9]), .Z(n71) );
  XOR2_X1 U93 ( .A(B[8]), .B(A[8]), .Z(n72) );
  XOR2_X1 U94 ( .A(n50), .B(n72), .Z(SUM[8]) );
  NAND2_X1 U95 ( .A1(carry[8]), .A2(B[8]), .ZN(n73) );
  NAND2_X1 U96 ( .A1(carry[8]), .A2(A[8]), .ZN(n74) );
  NAND2_X1 U97 ( .A1(B[8]), .A2(A[8]), .ZN(n75) );
  NAND3_X1 U98 ( .A1(n73), .A2(n74), .A3(n75), .ZN(carry[9]) );
  XOR2_X1 U99 ( .A(B[9]), .B(A[9]), .Z(n76) );
  XOR2_X1 U100 ( .A(n71), .B(n76), .Z(SUM[9]) );
  NAND2_X1 U101 ( .A1(n35), .A2(B[9]), .ZN(n77) );
  NAND2_X1 U102 ( .A1(carry[9]), .A2(A[9]), .ZN(n78) );
  NAND2_X1 U103 ( .A1(B[9]), .A2(A[9]), .ZN(n79) );
  NAND3_X1 U104 ( .A1(n78), .A2(n77), .A3(n79), .ZN(carry[10]) );
  XOR2_X1 U105 ( .A(B[1]), .B(A[1]), .Z(n80) );
  XOR2_X1 U106 ( .A(n88), .B(n80), .Z(SUM[1]) );
  NAND2_X1 U107 ( .A1(n88), .A2(B[1]), .ZN(n81) );
  NAND2_X1 U108 ( .A1(n88), .A2(A[1]), .ZN(n82) );
  NAND2_X1 U109 ( .A1(B[1]), .A2(A[1]), .ZN(n83) );
  NAND3_X1 U110 ( .A1(n81), .A2(n82), .A3(n83), .ZN(carry[2]) );
  XOR2_X1 U111 ( .A(B[2]), .B(A[2]), .Z(n84) );
  XOR2_X1 U112 ( .A(n66), .B(n84), .Z(SUM[2]) );
  NAND2_X1 U113 ( .A1(n65), .A2(B[2]), .ZN(n85) );
  NAND2_X1 U114 ( .A1(carry[2]), .A2(A[2]), .ZN(n86) );
  NAND2_X1 U115 ( .A1(B[2]), .A2(A[2]), .ZN(n87) );
  NAND3_X1 U116 ( .A1(n85), .A2(n86), .A3(n87), .ZN(carry[3]) );
  XOR2_X1 U117 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_16_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n313), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n312), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n316), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n315), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n318), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n94), .B(n88), .CI(n101), .CO(n53), .S(n54) );
  INV_X1 U157 ( .A(n308), .ZN(n307) );
  NAND3_X1 U158 ( .A1(n301), .A2(n302), .A3(n303), .ZN(n49) );
  CLKBUF_X1 U159 ( .A(n326), .Z(n206) );
  XNOR2_X1 U160 ( .A(a[2]), .B(a[1]), .ZN(n326) );
  CLKBUF_X1 U161 ( .A(n367), .Z(n207) );
  AND2_X1 U162 ( .A1(n102), .A2(n95), .ZN(n208) );
  AND3_X1 U163 ( .A1(n216), .A2(n215), .A3(n217), .ZN(product[15]) );
  NAND2_X1 U164 ( .A1(n326), .A2(n364), .ZN(n210) );
  NAND2_X1 U165 ( .A1(n326), .A2(n364), .ZN(n328) );
  XOR2_X1 U166 ( .A(n102), .B(n95), .Z(n56) );
  NAND3_X1 U167 ( .A1(n297), .A2(n298), .A3(n296), .ZN(n211) );
  NAND3_X1 U168 ( .A1(n297), .A2(n298), .A3(n296), .ZN(n212) );
  CLKBUF_X1 U169 ( .A(n56), .Z(n213) );
  XOR2_X1 U170 ( .A(n310), .B(n15), .Z(n214) );
  XOR2_X1 U171 ( .A(n212), .B(n214), .Z(product[14]) );
  NAND2_X1 U172 ( .A1(n211), .A2(n310), .ZN(n215) );
  NAND2_X1 U173 ( .A1(n2), .A2(n15), .ZN(n216) );
  NAND2_X1 U174 ( .A1(n310), .A2(n15), .ZN(n217) );
  NAND2_X1 U175 ( .A1(n11), .A2(n50), .ZN(n218) );
  CLKBUF_X1 U176 ( .A(b[4]), .Z(n219) );
  NAND2_X1 U177 ( .A1(n236), .A2(n23), .ZN(n220) );
  CLKBUF_X1 U178 ( .A(n293), .Z(n221) );
  CLKBUF_X1 U179 ( .A(b[1]), .Z(n267) );
  CLKBUF_X1 U180 ( .A(n220), .Z(n222) );
  CLKBUF_X1 U181 ( .A(n253), .Z(n223) );
  CLKBUF_X1 U182 ( .A(n240), .Z(n224) );
  CLKBUF_X1 U183 ( .A(n266), .Z(n225) );
  NAND3_X1 U184 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n226) );
  NAND3_X1 U185 ( .A1(n239), .A2(n224), .A3(n241), .ZN(n227) );
  NAND3_X1 U186 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n228) );
  NAND3_X1 U187 ( .A1(n223), .A2(n254), .A3(n255), .ZN(n229) );
  NAND3_X1 U188 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n230) );
  NAND3_X1 U189 ( .A1(n222), .A2(n258), .A3(n259), .ZN(n231) );
  CLKBUF_X1 U190 ( .A(n236), .Z(n232) );
  CLKBUF_X1 U191 ( .A(n251), .Z(n233) );
  CLKBUF_X1 U192 ( .A(n304), .Z(n234) );
  XNOR2_X2 U193 ( .A(a[4]), .B(a[3]), .ZN(n336) );
  NAND3_X1 U194 ( .A1(n304), .A2(n218), .A3(n305), .ZN(n235) );
  NAND3_X1 U195 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n236) );
  CLKBUF_X1 U196 ( .A(n218), .Z(n237) );
  XOR2_X1 U197 ( .A(n103), .B(n96), .Z(n238) );
  XOR2_X1 U198 ( .A(n14), .B(n238), .Z(product[2]) );
  NAND2_X1 U199 ( .A1(n14), .A2(n103), .ZN(n239) );
  NAND2_X1 U200 ( .A1(n14), .A2(n96), .ZN(n240) );
  NAND2_X1 U201 ( .A1(n103), .A2(n96), .ZN(n241) );
  NAND3_X1 U202 ( .A1(n240), .A2(n239), .A3(n241), .ZN(n13) );
  CLKBUF_X1 U203 ( .A(n263), .Z(n242) );
  CLKBUF_X1 U204 ( .A(n264), .Z(n243) );
  NAND3_X1 U205 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n244) );
  NAND3_X1 U206 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n245) );
  CLKBUF_X1 U207 ( .A(n277), .Z(n246) );
  XOR2_X1 U208 ( .A(n213), .B(n71), .Z(n247) );
  XOR2_X1 U209 ( .A(n227), .B(n247), .Z(product[3]) );
  NAND2_X1 U210 ( .A1(n13), .A2(n56), .ZN(n248) );
  NAND2_X1 U211 ( .A1(n226), .A2(n71), .ZN(n249) );
  NAND2_X1 U212 ( .A1(n56), .A2(n71), .ZN(n250) );
  NAND3_X1 U213 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n12) );
  NAND3_X1 U214 ( .A1(n283), .A2(n284), .A3(n285), .ZN(n251) );
  NAND2_X2 U215 ( .A1(n336), .A2(n365), .ZN(n338) );
  XOR2_X1 U216 ( .A(n34), .B(n39), .Z(n252) );
  XOR2_X1 U217 ( .A(n233), .B(n252), .Z(product[8]) );
  NAND2_X1 U218 ( .A1(n251), .A2(n34), .ZN(n253) );
  NAND2_X1 U219 ( .A1(n8), .A2(n39), .ZN(n254) );
  NAND2_X1 U220 ( .A1(n34), .A2(n39), .ZN(n255) );
  NAND3_X1 U221 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n7) );
  XOR2_X1 U222 ( .A(n23), .B(n20), .Z(n256) );
  XOR2_X1 U223 ( .A(n232), .B(n256), .Z(product[11]) );
  NAND2_X1 U224 ( .A1(n236), .A2(n23), .ZN(n257) );
  NAND2_X1 U225 ( .A1(n5), .A2(n20), .ZN(n258) );
  NAND2_X1 U226 ( .A1(n23), .A2(n20), .ZN(n259) );
  NAND3_X1 U227 ( .A1(n220), .A2(n258), .A3(n259), .ZN(n4) );
  NAND3_X1 U228 ( .A1(n264), .A2(n263), .A3(n265), .ZN(n260) );
  NAND3_X1 U229 ( .A1(n242), .A2(n243), .A3(n265), .ZN(n261) );
  XOR2_X1 U230 ( .A(n54), .B(n208), .Z(n262) );
  XOR2_X1 U231 ( .A(n245), .B(n262), .Z(product[4]) );
  NAND2_X1 U232 ( .A1(n12), .A2(n54), .ZN(n263) );
  NAND2_X1 U233 ( .A1(n244), .A2(n208), .ZN(n264) );
  NAND2_X1 U234 ( .A1(n54), .A2(n208), .ZN(n265) );
  NAND3_X1 U235 ( .A1(n263), .A2(n264), .A3(n265), .ZN(n11) );
  NAND3_X1 U236 ( .A1(n270), .A2(n269), .A3(n271), .ZN(n266) );
  XOR2_X1 U237 ( .A(n33), .B(n28), .Z(n268) );
  XOR2_X1 U238 ( .A(n229), .B(n268), .Z(product[9]) );
  NAND2_X1 U239 ( .A1(n7), .A2(n33), .ZN(n269) );
  NAND2_X1 U240 ( .A1(n228), .A2(n28), .ZN(n270) );
  NAND2_X1 U241 ( .A1(n33), .A2(n28), .ZN(n271) );
  NAND3_X1 U242 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n6) );
  NAND3_X1 U243 ( .A1(n304), .A2(n306), .A3(n305), .ZN(n272) );
  XOR2_X1 U244 ( .A(n24), .B(n27), .Z(n273) );
  XOR2_X1 U245 ( .A(n225), .B(n273), .Z(product[10]) );
  NAND2_X1 U246 ( .A1(n266), .A2(n24), .ZN(n274) );
  NAND2_X1 U247 ( .A1(n6), .A2(n27), .ZN(n275) );
  NAND2_X1 U248 ( .A1(n24), .A2(n27), .ZN(n276) );
  NAND3_X1 U249 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n5) );
  NAND3_X1 U250 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n277) );
  XOR2_X1 U251 ( .A(n46), .B(n49), .Z(n278) );
  XOR2_X1 U252 ( .A(n10), .B(n278), .Z(product[6]) );
  NAND2_X1 U253 ( .A1(n235), .A2(n46), .ZN(n279) );
  NAND2_X1 U254 ( .A1(n272), .A2(n49), .ZN(n280) );
  NAND2_X1 U255 ( .A1(n46), .A2(n49), .ZN(n281) );
  NAND3_X1 U256 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n9) );
  XOR2_X1 U257 ( .A(n40), .B(n45), .Z(n282) );
  XOR2_X1 U258 ( .A(n246), .B(n282), .Z(product[7]) );
  NAND2_X1 U259 ( .A1(n277), .A2(n40), .ZN(n283) );
  NAND2_X1 U260 ( .A1(n9), .A2(n45), .ZN(n284) );
  NAND2_X1 U261 ( .A1(n40), .A2(n45), .ZN(n285) );
  NAND3_X1 U262 ( .A1(n283), .A2(n284), .A3(n285), .ZN(n8) );
  INV_X1 U263 ( .A(n308), .ZN(n286) );
  INV_X1 U264 ( .A(n286), .ZN(n287) );
  NAND3_X1 U265 ( .A1(n293), .A2(n294), .A3(n292), .ZN(n288) );
  NAND3_X1 U266 ( .A1(n221), .A2(n292), .A3(n294), .ZN(n289) );
  XNOR2_X1 U267 ( .A(b[2]), .B(a[1]), .ZN(n290) );
  XOR2_X1 U268 ( .A(n299), .B(n52), .Z(n50) );
  INV_X1 U269 ( .A(n15), .ZN(n309) );
  INV_X1 U270 ( .A(n345), .ZN(n313) );
  INV_X1 U271 ( .A(n21), .ZN(n312) );
  INV_X1 U272 ( .A(n325), .ZN(n318) );
  INV_X1 U273 ( .A(n334), .ZN(n316) );
  INV_X1 U274 ( .A(b[0]), .ZN(n308) );
  INV_X1 U275 ( .A(n356), .ZN(n310) );
  INV_X1 U276 ( .A(n31), .ZN(n315) );
  INV_X1 U277 ( .A(a[0]), .ZN(n320) );
  INV_X1 U278 ( .A(a[5]), .ZN(n314) );
  INV_X1 U279 ( .A(a[7]), .ZN(n311) );
  XOR2_X1 U280 ( .A(n19), .B(n18), .Z(n291) );
  XOR2_X1 U281 ( .A(n291), .B(n231), .Z(product[12]) );
  NAND2_X1 U282 ( .A1(n19), .A2(n18), .ZN(n292) );
  NAND2_X1 U283 ( .A1(n4), .A2(n19), .ZN(n293) );
  NAND2_X1 U284 ( .A1(n18), .A2(n230), .ZN(n294) );
  NAND3_X1 U285 ( .A1(n294), .A2(n293), .A3(n292), .ZN(n3) );
  XOR2_X1 U286 ( .A(n17), .B(n309), .Z(n295) );
  XOR2_X1 U287 ( .A(n295), .B(n289), .Z(product[13]) );
  NAND2_X1 U288 ( .A1(n17), .A2(n309), .ZN(n296) );
  NAND2_X1 U289 ( .A1(n288), .A2(n17), .ZN(n297) );
  NAND2_X1 U290 ( .A1(n3), .A2(n309), .ZN(n298) );
  NAND3_X1 U291 ( .A1(n297), .A2(n298), .A3(n296), .ZN(n2) );
  XOR2_X1 U292 ( .A(n93), .B(n100), .Z(n299) );
  XOR2_X1 U293 ( .A(n53), .B(n261), .Z(n300) );
  XOR2_X1 U294 ( .A(n300), .B(n50), .Z(product[5]) );
  NAND2_X1 U295 ( .A1(n93), .A2(n100), .ZN(n301) );
  NAND2_X1 U296 ( .A1(n93), .A2(n52), .ZN(n302) );
  NAND2_X1 U297 ( .A1(n52), .A2(n100), .ZN(n303) );
  NAND2_X1 U298 ( .A1(n53), .A2(n260), .ZN(n304) );
  NAND2_X1 U299 ( .A1(n50), .A2(n53), .ZN(n305) );
  NAND2_X1 U300 ( .A1(n11), .A2(n50), .ZN(n306) );
  NAND3_X1 U301 ( .A1(n234), .A2(n305), .A3(n237), .ZN(n10) );
  INV_X1 U302 ( .A(a[3]), .ZN(n317) );
  INV_X1 U303 ( .A(a[1]), .ZN(n319) );
  XOR2_X2 U304 ( .A(a[6]), .B(n314), .Z(n347) );
  NOR2_X1 U305 ( .A1(n320), .A2(n287), .ZN(product[0]) );
  OAI22_X1 U306 ( .A1(n321), .A2(n322), .B1(n323), .B2(n320), .ZN(n99) );
  OAI22_X1 U307 ( .A1(n323), .A2(n322), .B1(n324), .B2(n320), .ZN(n98) );
  XNOR2_X1 U308 ( .A(b[6]), .B(a[1]), .ZN(n323) );
  OAI22_X1 U309 ( .A1(n320), .A2(n324), .B1(n322), .B2(n324), .ZN(n325) );
  XNOR2_X1 U310 ( .A(b[7]), .B(a[1]), .ZN(n324) );
  NOR2_X1 U311 ( .A1(n326), .A2(n287), .ZN(n96) );
  OAI22_X1 U312 ( .A1(n327), .A2(n328), .B1(n326), .B2(n329), .ZN(n95) );
  XNOR2_X1 U313 ( .A(a[3]), .B(n307), .ZN(n327) );
  OAI22_X1 U314 ( .A1(n329), .A2(n328), .B1(n326), .B2(n330), .ZN(n94) );
  XNOR2_X1 U315 ( .A(b[1]), .B(a[3]), .ZN(n329) );
  OAI22_X1 U316 ( .A1(n330), .A2(n210), .B1(n206), .B2(n331), .ZN(n93) );
  XNOR2_X1 U317 ( .A(b[2]), .B(a[3]), .ZN(n330) );
  OAI22_X1 U318 ( .A1(n331), .A2(n210), .B1(n326), .B2(n332), .ZN(n92) );
  XNOR2_X1 U319 ( .A(b[3]), .B(a[3]), .ZN(n331) );
  OAI22_X1 U320 ( .A1(n332), .A2(n210), .B1(n206), .B2(n333), .ZN(n91) );
  XNOR2_X1 U321 ( .A(b[4]), .B(a[3]), .ZN(n332) );
  OAI22_X1 U322 ( .A1(n335), .A2(n206), .B1(n210), .B2(n335), .ZN(n334) );
  NOR2_X1 U323 ( .A1(n336), .A2(n287), .ZN(n88) );
  OAI22_X1 U324 ( .A1(n337), .A2(n338), .B1(n336), .B2(n339), .ZN(n87) );
  XNOR2_X1 U325 ( .A(a[5]), .B(n286), .ZN(n337) );
  OAI22_X1 U326 ( .A1(n339), .A2(n338), .B1(n336), .B2(n340), .ZN(n86) );
  XNOR2_X1 U327 ( .A(n267), .B(a[5]), .ZN(n339) );
  OAI22_X1 U328 ( .A1(n340), .A2(n338), .B1(n336), .B2(n341), .ZN(n85) );
  XNOR2_X1 U329 ( .A(b[2]), .B(a[5]), .ZN(n340) );
  OAI22_X1 U330 ( .A1(n341), .A2(n338), .B1(n336), .B2(n342), .ZN(n84) );
  XNOR2_X1 U331 ( .A(b[3]), .B(a[5]), .ZN(n341) );
  OAI22_X1 U332 ( .A1(n342), .A2(n338), .B1(n336), .B2(n343), .ZN(n83) );
  XNOR2_X1 U333 ( .A(n219), .B(a[5]), .ZN(n342) );
  OAI22_X1 U334 ( .A1(n343), .A2(n338), .B1(n336), .B2(n344), .ZN(n82) );
  XNOR2_X1 U335 ( .A(b[5]), .B(a[5]), .ZN(n343) );
  OAI22_X1 U336 ( .A1(n346), .A2(n336), .B1(n338), .B2(n346), .ZN(n345) );
  NOR2_X1 U337 ( .A1(n347), .A2(n287), .ZN(n80) );
  OAI22_X1 U338 ( .A1(n348), .A2(n349), .B1(n347), .B2(n350), .ZN(n79) );
  XNOR2_X1 U339 ( .A(a[7]), .B(n307), .ZN(n348) );
  OAI22_X1 U340 ( .A1(n351), .A2(n349), .B1(n347), .B2(n352), .ZN(n77) );
  OAI22_X1 U341 ( .A1(n352), .A2(n349), .B1(n347), .B2(n353), .ZN(n76) );
  XNOR2_X1 U342 ( .A(b[3]), .B(a[7]), .ZN(n352) );
  OAI22_X1 U343 ( .A1(n353), .A2(n349), .B1(n347), .B2(n354), .ZN(n75) );
  XNOR2_X1 U344 ( .A(n219), .B(a[7]), .ZN(n353) );
  OAI22_X1 U345 ( .A1(n354), .A2(n349), .B1(n347), .B2(n355), .ZN(n74) );
  XNOR2_X1 U346 ( .A(b[5]), .B(a[7]), .ZN(n354) );
  OAI22_X1 U347 ( .A1(n357), .A2(n347), .B1(n349), .B2(n357), .ZN(n356) );
  OAI21_X1 U348 ( .B1(n286), .B2(n319), .A(n322), .ZN(n72) );
  OAI21_X1 U349 ( .B1(n317), .B2(n210), .A(n358), .ZN(n71) );
  OR3_X1 U350 ( .A1(n326), .A2(n307), .A3(n317), .ZN(n358) );
  OAI21_X1 U351 ( .B1(n314), .B2(n338), .A(n359), .ZN(n70) );
  OR3_X1 U352 ( .A1(n336), .A2(n307), .A3(n314), .ZN(n359) );
  OAI21_X1 U353 ( .B1(n311), .B2(n349), .A(n360), .ZN(n69) );
  OR3_X1 U354 ( .A1(n347), .A2(n286), .A3(n311), .ZN(n360) );
  XNOR2_X1 U355 ( .A(n361), .B(n362), .ZN(n38) );
  OR2_X1 U356 ( .A1(n361), .A2(n362), .ZN(n37) );
  OAI22_X1 U357 ( .A1(n333), .A2(n210), .B1(n206), .B2(n363), .ZN(n362) );
  XNOR2_X1 U358 ( .A(b[5]), .B(a[3]), .ZN(n333) );
  OAI22_X1 U359 ( .A1(n350), .A2(n349), .B1(n347), .B2(n351), .ZN(n361) );
  XNOR2_X1 U360 ( .A(b[2]), .B(a[7]), .ZN(n351) );
  XNOR2_X1 U361 ( .A(n267), .B(a[7]), .ZN(n350) );
  OAI22_X1 U362 ( .A1(n363), .A2(n210), .B1(n206), .B2(n335), .ZN(n31) );
  XNOR2_X1 U363 ( .A(b[7]), .B(a[3]), .ZN(n335) );
  XNOR2_X1 U364 ( .A(n317), .B(a[2]), .ZN(n364) );
  XNOR2_X1 U365 ( .A(b[6]), .B(a[3]), .ZN(n363) );
  OAI22_X1 U366 ( .A1(n344), .A2(n338), .B1(n336), .B2(n346), .ZN(n21) );
  XNOR2_X1 U367 ( .A(b[7]), .B(a[5]), .ZN(n346) );
  XNOR2_X1 U368 ( .A(n314), .B(a[4]), .ZN(n365) );
  XNOR2_X1 U369 ( .A(b[6]), .B(a[5]), .ZN(n344) );
  OAI22_X1 U370 ( .A1(n355), .A2(n349), .B1(n347), .B2(n357), .ZN(n15) );
  XNOR2_X1 U371 ( .A(b[7]), .B(a[7]), .ZN(n357) );
  NAND2_X1 U372 ( .A1(n347), .A2(n366), .ZN(n349) );
  XNOR2_X1 U373 ( .A(n311), .B(a[6]), .ZN(n366) );
  XNOR2_X1 U374 ( .A(b[6]), .B(a[7]), .ZN(n355) );
  OAI22_X1 U375 ( .A1(n307), .A2(n322), .B1(n367), .B2(n320), .ZN(n104) );
  OAI22_X1 U376 ( .A1(n207), .A2(n322), .B1(n368), .B2(n320), .ZN(n103) );
  XNOR2_X1 U377 ( .A(b[1]), .B(a[1]), .ZN(n367) );
  OAI22_X1 U378 ( .A1(n290), .A2(n322), .B1(n369), .B2(n320), .ZN(n102) );
  XNOR2_X1 U379 ( .A(b[2]), .B(a[1]), .ZN(n368) );
  OAI22_X1 U380 ( .A1(n369), .A2(n322), .B1(n370), .B2(n320), .ZN(n101) );
  XNOR2_X1 U381 ( .A(b[3]), .B(a[1]), .ZN(n369) );
  OAI22_X1 U382 ( .A1(n370), .A2(n322), .B1(n321), .B2(n320), .ZN(n100) );
  XNOR2_X1 U383 ( .A(b[5]), .B(a[1]), .ZN(n321) );
  NAND2_X1 U384 ( .A1(a[1]), .A2(n320), .ZN(n322) );
  XNOR2_X1 U385 ( .A(b[4]), .B(a[1]), .ZN(n370) );
endmodule


module mac_16 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   n6, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, n2, n4;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(n6), .QN(n2) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  mac_16_DW01_add_0 add_356 ( .A(pipeline), .B({mac_out[15:1], n6}), .CI(1'b0), 
        .SUM(sum) );
  mac_16_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n4), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n4), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n4), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n4), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n4), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n4), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n4), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n4), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n4), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n4), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n4), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n4), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n4), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n4), .ZN(N6) );
  INV_X1 U18 ( .A(n2), .ZN(mac_out[0]) );
  AND2_X1 U19 ( .A1(sum[0]), .A2(n4), .ZN(N3) );
  AND2_X1 U20 ( .A1(sum[15]), .A2(n4), .ZN(N18) );
  INV_X1 U21 ( .A(clear_acc), .ZN(n4) );
endmodule


module mac_15_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74;
  wire   [15:1] carry;

  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n74) );
  XOR2_X1 U2 ( .A(B[15]), .B(A[15]), .Z(n1) );
  XOR2_X1 U3 ( .A(carry[15]), .B(n1), .Z(SUM[15]) );
  NAND3_X1 U4 ( .A1(n9), .A2(n10), .A3(n11), .ZN(n2) );
  NAND3_X1 U5 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n3) );
  NAND3_X1 U6 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n4) );
  NAND3_X1 U7 ( .A1(n13), .A2(n14), .A3(n15), .ZN(n5) );
  NAND3_X1 U8 ( .A1(n13), .A2(n14), .A3(n15), .ZN(n6) );
  NAND3_X1 U9 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n7) );
  XOR2_X1 U10 ( .A(B[9]), .B(A[9]), .Z(n8) );
  XOR2_X1 U11 ( .A(carry[9]), .B(n8), .Z(SUM[9]) );
  NAND2_X1 U12 ( .A1(carry[9]), .A2(B[9]), .ZN(n9) );
  NAND2_X1 U13 ( .A1(carry[9]), .A2(A[9]), .ZN(n10) );
  NAND2_X1 U14 ( .A1(B[9]), .A2(A[9]), .ZN(n11) );
  NAND3_X1 U15 ( .A1(n9), .A2(n10), .A3(n11), .ZN(carry[10]) );
  XOR2_X1 U16 ( .A(B[2]), .B(A[2]), .Z(n12) );
  XOR2_X1 U17 ( .A(n4), .B(n12), .Z(SUM[2]) );
  NAND2_X1 U18 ( .A1(n3), .A2(B[2]), .ZN(n13) );
  NAND2_X1 U19 ( .A1(carry[2]), .A2(A[2]), .ZN(n14) );
  NAND2_X1 U20 ( .A1(B[2]), .A2(A[2]), .ZN(n15) );
  NAND3_X1 U21 ( .A1(n13), .A2(n14), .A3(n15), .ZN(carry[3]) );
  NAND3_X1 U22 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n16) );
  XOR2_X1 U23 ( .A(B[10]), .B(A[10]), .Z(n17) );
  XOR2_X1 U24 ( .A(n2), .B(n17), .Z(SUM[10]) );
  NAND2_X1 U25 ( .A1(n2), .A2(B[10]), .ZN(n18) );
  NAND2_X1 U26 ( .A1(carry[10]), .A2(A[10]), .ZN(n19) );
  NAND2_X1 U27 ( .A1(B[10]), .A2(A[10]), .ZN(n20) );
  NAND3_X1 U28 ( .A1(n19), .A2(n18), .A3(n20), .ZN(carry[11]) );
  NAND3_X1 U29 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n21) );
  NAND3_X1 U30 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n22) );
  XOR2_X1 U31 ( .A(B[3]), .B(A[3]), .Z(n23) );
  XOR2_X1 U32 ( .A(n6), .B(n23), .Z(SUM[3]) );
  NAND2_X1 U33 ( .A1(n5), .A2(B[3]), .ZN(n24) );
  NAND2_X1 U34 ( .A1(carry[3]), .A2(A[3]), .ZN(n25) );
  NAND2_X1 U35 ( .A1(B[3]), .A2(A[3]), .ZN(n26) );
  NAND3_X1 U36 ( .A1(n24), .A2(n25), .A3(n26), .ZN(carry[4]) );
  NAND3_X1 U37 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n27) );
  NAND3_X1 U38 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n28) );
  XOR2_X1 U39 ( .A(B[11]), .B(A[11]), .Z(n29) );
  XOR2_X1 U40 ( .A(n7), .B(n29), .Z(SUM[11]) );
  NAND2_X1 U41 ( .A1(n7), .A2(B[11]), .ZN(n30) );
  NAND2_X1 U42 ( .A1(carry[11]), .A2(A[11]), .ZN(n31) );
  NAND2_X1 U43 ( .A1(B[11]), .A2(A[11]), .ZN(n32) );
  NAND3_X1 U44 ( .A1(n30), .A2(n31), .A3(n32), .ZN(carry[12]) );
  XOR2_X1 U45 ( .A(B[4]), .B(A[4]), .Z(n33) );
  XOR2_X1 U46 ( .A(n22), .B(n33), .Z(SUM[4]) );
  NAND2_X1 U47 ( .A1(n21), .A2(B[4]), .ZN(n34) );
  NAND2_X1 U48 ( .A1(carry[4]), .A2(A[4]), .ZN(n35) );
  NAND2_X1 U49 ( .A1(B[4]), .A2(A[4]), .ZN(n36) );
  NAND3_X1 U50 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[5]) );
  NAND3_X1 U51 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n37) );
  XOR2_X1 U52 ( .A(B[5]), .B(A[5]), .Z(n38) );
  XOR2_X1 U53 ( .A(n28), .B(n38), .Z(SUM[5]) );
  NAND2_X1 U54 ( .A1(n28), .A2(B[5]), .ZN(n39) );
  NAND2_X1 U55 ( .A1(carry[5]), .A2(A[5]), .ZN(n40) );
  NAND2_X1 U56 ( .A1(B[5]), .A2(A[5]), .ZN(n41) );
  NAND3_X1 U57 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[6]) );
  NAND3_X1 U58 ( .A1(n44), .A2(n45), .A3(n46), .ZN(n42) );
  XOR2_X1 U59 ( .A(B[12]), .B(A[12]), .Z(n43) );
  XOR2_X1 U60 ( .A(n27), .B(n43), .Z(SUM[12]) );
  NAND2_X1 U61 ( .A1(n27), .A2(B[12]), .ZN(n44) );
  NAND2_X1 U62 ( .A1(carry[12]), .A2(A[12]), .ZN(n45) );
  NAND2_X1 U63 ( .A1(B[12]), .A2(A[12]), .ZN(n46) );
  NAND3_X1 U64 ( .A1(n44), .A2(n45), .A3(n46), .ZN(carry[13]) );
  NAND3_X1 U65 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n47) );
  NAND3_X1 U66 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n48) );
  NAND3_X1 U67 ( .A1(n71), .A2(n72), .A3(n73), .ZN(n49) );
  XOR2_X1 U68 ( .A(B[8]), .B(A[8]), .Z(n50) );
  XOR2_X1 U69 ( .A(n49), .B(n50), .Z(SUM[8]) );
  NAND2_X1 U70 ( .A1(n49), .A2(B[8]), .ZN(n51) );
  NAND2_X1 U71 ( .A1(carry[8]), .A2(A[8]), .ZN(n52) );
  NAND2_X1 U72 ( .A1(B[8]), .A2(A[8]), .ZN(n53) );
  NAND3_X1 U73 ( .A1(n51), .A2(n52), .A3(n53), .ZN(carry[9]) );
  XOR2_X1 U74 ( .A(B[1]), .B(A[1]), .Z(n54) );
  XOR2_X1 U75 ( .A(n74), .B(n54), .Z(SUM[1]) );
  NAND2_X1 U76 ( .A1(n74), .A2(B[1]), .ZN(n55) );
  NAND2_X1 U77 ( .A1(n74), .A2(A[1]), .ZN(n56) );
  NAND2_X1 U78 ( .A1(B[1]), .A2(A[1]), .ZN(n57) );
  NAND3_X1 U79 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[2]) );
  XOR2_X1 U80 ( .A(B[13]), .B(A[13]), .Z(n58) );
  XOR2_X1 U81 ( .A(n42), .B(n58), .Z(SUM[13]) );
  NAND2_X1 U82 ( .A1(n42), .A2(B[13]), .ZN(n59) );
  NAND2_X1 U83 ( .A1(carry[13]), .A2(A[13]), .ZN(n60) );
  NAND2_X1 U84 ( .A1(B[13]), .A2(A[13]), .ZN(n61) );
  NAND3_X1 U85 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[14]) );
  XOR2_X1 U86 ( .A(B[6]), .B(A[6]), .Z(n62) );
  XOR2_X1 U87 ( .A(carry[6]), .B(n62), .Z(SUM[6]) );
  NAND2_X1 U88 ( .A1(n37), .A2(B[6]), .ZN(n63) );
  NAND2_X1 U89 ( .A1(carry[6]), .A2(A[6]), .ZN(n64) );
  NAND2_X1 U90 ( .A1(B[6]), .A2(A[6]), .ZN(n65) );
  NAND3_X1 U91 ( .A1(n63), .A2(n64), .A3(n65), .ZN(carry[7]) );
  XOR2_X1 U92 ( .A(B[14]), .B(A[14]), .Z(n66) );
  XOR2_X1 U93 ( .A(n16), .B(n66), .Z(SUM[14]) );
  NAND2_X1 U94 ( .A1(n16), .A2(B[14]), .ZN(n67) );
  NAND2_X1 U95 ( .A1(carry[14]), .A2(A[14]), .ZN(n68) );
  NAND2_X1 U96 ( .A1(B[14]), .A2(A[14]), .ZN(n69) );
  NAND3_X1 U97 ( .A1(n67), .A2(n68), .A3(n69), .ZN(carry[15]) );
  XOR2_X1 U98 ( .A(B[7]), .B(A[7]), .Z(n70) );
  XOR2_X1 U99 ( .A(n48), .B(n70), .Z(SUM[7]) );
  NAND2_X1 U100 ( .A1(n47), .A2(B[7]), .ZN(n71) );
  NAND2_X1 U101 ( .A1(carry[7]), .A2(A[7]), .ZN(n72) );
  NAND2_X1 U102 ( .A1(B[7]), .A2(A[7]), .ZN(n73) );
  NAND3_X1 U103 ( .A1(n72), .A2(n71), .A3(n73), .ZN(carry[8]) );
  XOR2_X1 U104 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_15_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n302), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n301), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n305), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n304), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n307), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  INV_X1 U157 ( .A(n297), .ZN(n296) );
  CLKBUF_X1 U158 ( .A(n257), .Z(n206) );
  AND2_X1 U159 ( .A1(n208), .A2(n102), .ZN(n207) );
  OAI22_X1 U160 ( .A1(n316), .A2(n317), .B1(n286), .B2(n318), .ZN(n208) );
  BUF_X1 U161 ( .A(n325), .Z(n209) );
  BUF_X1 U162 ( .A(n325), .Z(n210) );
  XNOR2_X1 U163 ( .A(a[4]), .B(a[3]), .ZN(n325) );
  CLKBUF_X1 U164 ( .A(a[1]), .Z(n211) );
  CLKBUF_X1 U165 ( .A(n297), .Z(n212) );
  CLKBUF_X1 U166 ( .A(b[1]), .Z(n213) );
  XNOR2_X1 U167 ( .A(a[6]), .B(a[5]), .ZN(n336) );
  CLKBUF_X1 U168 ( .A(n219), .Z(n214) );
  NAND3_X1 U169 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n215) );
  CLKBUF_X1 U170 ( .A(n56), .Z(n216) );
  AND2_X1 U171 ( .A1(n104), .A2(n72), .ZN(n217) );
  CLKBUF_X1 U172 ( .A(n3), .Z(n218) );
  NAND3_X1 U173 ( .A1(n282), .A2(n283), .A3(n284), .ZN(n219) );
  NAND3_X1 U174 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n220) );
  CLKBUF_X1 U175 ( .A(n255), .Z(n221) );
  NAND3_X1 U176 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n222) );
  NAND3_X1 U177 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n223) );
  NAND3_X1 U178 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n224) );
  NAND3_X1 U179 ( .A1(n254), .A2(n221), .A3(n256), .ZN(n225) );
  CLKBUF_X1 U180 ( .A(n258), .Z(n226) );
  NAND3_X1 U181 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n227) );
  XOR2_X1 U182 ( .A(n46), .B(n49), .Z(n228) );
  XOR2_X1 U183 ( .A(n214), .B(n228), .Z(product[6]) );
  NAND2_X1 U184 ( .A1(n219), .A2(n46), .ZN(n229) );
  NAND2_X1 U185 ( .A1(n10), .A2(n49), .ZN(n230) );
  NAND2_X1 U186 ( .A1(n46), .A2(n49), .ZN(n231) );
  NAND3_X1 U187 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n9) );
  CLKBUF_X1 U188 ( .A(n213), .Z(n232) );
  CLKBUF_X1 U189 ( .A(n274), .Z(n233) );
  NAND3_X1 U190 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n234) );
  NAND2_X1 U191 ( .A1(n210), .A2(n354), .ZN(n235) );
  NAND2_X1 U192 ( .A1(n209), .A2(n354), .ZN(n236) );
  NAND2_X1 U193 ( .A1(n325), .A2(n354), .ZN(n327) );
  NAND3_X1 U194 ( .A1(n294), .A2(n293), .A3(n295), .ZN(n237) );
  CLKBUF_X1 U195 ( .A(n6), .Z(n238) );
  XOR2_X1 U196 ( .A(n33), .B(n28), .Z(n239) );
  XOR2_X1 U197 ( .A(n225), .B(n239), .Z(product[9]) );
  NAND2_X1 U198 ( .A1(n224), .A2(n33), .ZN(n240) );
  NAND2_X1 U199 ( .A1(n7), .A2(n28), .ZN(n241) );
  NAND2_X1 U200 ( .A1(n33), .A2(n28), .ZN(n242) );
  NAND3_X1 U201 ( .A1(n241), .A2(n240), .A3(n242), .ZN(n6) );
  CLKBUF_X1 U202 ( .A(n8), .Z(n243) );
  XOR2_X1 U203 ( .A(n40), .B(n45), .Z(n244) );
  XOR2_X1 U204 ( .A(n9), .B(n244), .Z(product[7]) );
  NAND2_X1 U205 ( .A1(n215), .A2(n40), .ZN(n245) );
  NAND2_X1 U206 ( .A1(n215), .A2(n45), .ZN(n246) );
  NAND2_X1 U207 ( .A1(n40), .A2(n45), .ZN(n247) );
  NAND3_X1 U208 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n8) );
  XOR2_X1 U209 ( .A(n103), .B(n96), .Z(n248) );
  XOR2_X1 U210 ( .A(n217), .B(n248), .Z(product[2]) );
  NAND2_X1 U211 ( .A1(n217), .A2(n103), .ZN(n249) );
  NAND2_X1 U212 ( .A1(n14), .A2(n96), .ZN(n250) );
  NAND2_X1 U213 ( .A1(n103), .A2(n96), .ZN(n251) );
  NAND3_X1 U214 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n13) );
  NAND3_X1 U215 ( .A1(n274), .A2(n273), .A3(n275), .ZN(n252) );
  XOR2_X1 U216 ( .A(n34), .B(n39), .Z(n253) );
  XOR2_X1 U217 ( .A(n243), .B(n253), .Z(product[8]) );
  NAND2_X1 U218 ( .A1(n227), .A2(n34), .ZN(n254) );
  NAND2_X1 U219 ( .A1(n8), .A2(n39), .ZN(n255) );
  NAND2_X1 U220 ( .A1(n34), .A2(n39), .ZN(n256) );
  NAND3_X1 U221 ( .A1(n255), .A2(n254), .A3(n256), .ZN(n7) );
  NAND3_X1 U222 ( .A1(n265), .A2(n267), .A3(n266), .ZN(n257) );
  NAND3_X1 U223 ( .A1(n262), .A2(n261), .A3(n263), .ZN(n258) );
  NAND3_X1 U224 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n259) );
  XOR2_X1 U225 ( .A(n20), .B(n23), .Z(n260) );
  XOR2_X1 U226 ( .A(n5), .B(n260), .Z(product[11]) );
  NAND2_X1 U227 ( .A1(n252), .A2(n20), .ZN(n261) );
  NAND2_X1 U228 ( .A1(n220), .A2(n23), .ZN(n262) );
  NAND2_X1 U229 ( .A1(n20), .A2(n23), .ZN(n263) );
  NAND3_X1 U230 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n4) );
  XOR2_X1 U231 ( .A(n216), .B(n71), .Z(n264) );
  XOR2_X1 U232 ( .A(n223), .B(n264), .Z(product[3]) );
  NAND2_X1 U233 ( .A1(n223), .A2(n56), .ZN(n265) );
  NAND2_X1 U234 ( .A1(n13), .A2(n71), .ZN(n266) );
  NAND2_X1 U235 ( .A1(n56), .A2(n71), .ZN(n267) );
  NAND3_X1 U236 ( .A1(n265), .A2(n266), .A3(n267), .ZN(n12) );
  XOR2_X1 U237 ( .A(n298), .B(n17), .Z(n268) );
  XOR2_X1 U238 ( .A(n218), .B(n268), .Z(product[13]) );
  NAND2_X1 U239 ( .A1(n3), .A2(n298), .ZN(n269) );
  NAND2_X1 U240 ( .A1(n237), .A2(n17), .ZN(n270) );
  NAND2_X1 U241 ( .A1(n298), .A2(n17), .ZN(n271) );
  NAND3_X1 U242 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n2) );
  XOR2_X1 U243 ( .A(n208), .B(n102), .Z(n56) );
  XOR2_X1 U244 ( .A(n27), .B(n24), .Z(n272) );
  XOR2_X1 U245 ( .A(n238), .B(n272), .Z(product[10]) );
  NAND2_X1 U246 ( .A1(n222), .A2(n27), .ZN(n273) );
  NAND2_X1 U247 ( .A1(n6), .A2(n24), .ZN(n274) );
  NAND2_X1 U248 ( .A1(n27), .A2(n24), .ZN(n275) );
  NAND3_X1 U249 ( .A1(n273), .A2(n233), .A3(n275), .ZN(n5) );
  CLKBUF_X1 U250 ( .A(n259), .Z(n276) );
  XOR2_X1 U251 ( .A(n54), .B(n207), .Z(n277) );
  XOR2_X1 U252 ( .A(n206), .B(n277), .Z(product[4]) );
  NAND2_X1 U253 ( .A1(n257), .A2(n54), .ZN(n278) );
  NAND2_X1 U254 ( .A1(n12), .A2(n207), .ZN(n279) );
  NAND2_X1 U255 ( .A1(n54), .A2(n207), .ZN(n280) );
  NAND3_X1 U256 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n11) );
  XOR2_X1 U257 ( .A(n50), .B(n53), .Z(n281) );
  XOR2_X1 U258 ( .A(n276), .B(n281), .Z(product[5]) );
  NAND2_X1 U259 ( .A1(n259), .A2(n50), .ZN(n282) );
  NAND2_X1 U260 ( .A1(n11), .A2(n53), .ZN(n283) );
  NAND2_X1 U261 ( .A1(n50), .A2(n53), .ZN(n284) );
  NAND3_X1 U262 ( .A1(n282), .A2(n283), .A3(n284), .ZN(n10) );
  NAND2_X2 U263 ( .A1(n315), .A2(n353), .ZN(n317) );
  XOR2_X1 U264 ( .A(a[2]), .B(n308), .Z(n285) );
  XOR2_X1 U265 ( .A(a[2]), .B(n308), .Z(n286) );
  INV_X1 U266 ( .A(n15), .ZN(n298) );
  XNOR2_X1 U267 ( .A(n226), .B(n287), .ZN(product[12]) );
  XNOR2_X1 U268 ( .A(n19), .B(n18), .ZN(n287) );
  XNOR2_X1 U269 ( .A(n234), .B(n288), .ZN(product[14]) );
  XNOR2_X1 U270 ( .A(n299), .B(n15), .ZN(n288) );
  AND3_X1 U271 ( .A1(n291), .A2(n290), .A3(n292), .ZN(product[15]) );
  OAI22_X1 U272 ( .A1(n344), .A2(n338), .B1(n336), .B2(n346), .ZN(n15) );
  INV_X1 U273 ( .A(n323), .ZN(n305) );
  INV_X1 U274 ( .A(n334), .ZN(n302) );
  INV_X1 U275 ( .A(n21), .ZN(n301) );
  INV_X1 U276 ( .A(n314), .ZN(n307) );
  INV_X1 U277 ( .A(b[0]), .ZN(n297) );
  INV_X1 U278 ( .A(n31), .ZN(n304) );
  XOR2_X1 U279 ( .A(a[2]), .B(n308), .Z(n315) );
  INV_X1 U280 ( .A(a[0]), .ZN(n309) );
  INV_X1 U281 ( .A(a[5]), .ZN(n303) );
  INV_X1 U282 ( .A(a[7]), .ZN(n300) );
  NAND2_X1 U283 ( .A1(n2), .A2(n299), .ZN(n290) );
  NAND2_X1 U284 ( .A1(n2), .A2(n15), .ZN(n291) );
  NAND2_X1 U285 ( .A1(n299), .A2(n15), .ZN(n292) );
  NAND2_X1 U286 ( .A1(n4), .A2(n19), .ZN(n293) );
  NAND2_X1 U287 ( .A1(n258), .A2(n18), .ZN(n294) );
  NAND2_X1 U288 ( .A1(n19), .A2(n18), .ZN(n295) );
  NAND3_X1 U289 ( .A1(n294), .A2(n293), .A3(n295), .ZN(n3) );
  INV_X1 U290 ( .A(n345), .ZN(n299) );
  INV_X1 U291 ( .A(a[3]), .ZN(n306) );
  INV_X1 U292 ( .A(a[1]), .ZN(n308) );
  NOR2_X1 U293 ( .A1(n309), .A2(n212), .ZN(product[0]) );
  OAI22_X1 U294 ( .A1(n310), .A2(n311), .B1(n312), .B2(n309), .ZN(n99) );
  OAI22_X1 U295 ( .A1(n312), .A2(n311), .B1(n313), .B2(n309), .ZN(n98) );
  XNOR2_X1 U296 ( .A(b[6]), .B(n211), .ZN(n312) );
  OAI22_X1 U297 ( .A1(n309), .A2(n313), .B1(n311), .B2(n313), .ZN(n314) );
  XNOR2_X1 U298 ( .A(b[7]), .B(n211), .ZN(n313) );
  NOR2_X1 U299 ( .A1(n285), .A2(n212), .ZN(n96) );
  XNOR2_X1 U300 ( .A(a[3]), .B(n296), .ZN(n316) );
  OAI22_X1 U301 ( .A1(n318), .A2(n317), .B1(n286), .B2(n319), .ZN(n94) );
  XNOR2_X1 U302 ( .A(n213), .B(a[3]), .ZN(n318) );
  OAI22_X1 U303 ( .A1(n319), .A2(n317), .B1(n285), .B2(n320), .ZN(n93) );
  XNOR2_X1 U304 ( .A(b[2]), .B(a[3]), .ZN(n319) );
  OAI22_X1 U305 ( .A1(n320), .A2(n317), .B1(n286), .B2(n321), .ZN(n92) );
  XNOR2_X1 U306 ( .A(b[3]), .B(a[3]), .ZN(n320) );
  OAI22_X1 U307 ( .A1(n321), .A2(n317), .B1(n286), .B2(n322), .ZN(n91) );
  XNOR2_X1 U308 ( .A(b[4]), .B(a[3]), .ZN(n321) );
  OAI22_X1 U309 ( .A1(n324), .A2(n285), .B1(n317), .B2(n324), .ZN(n323) );
  NOR2_X1 U310 ( .A1(n210), .A2(n212), .ZN(n88) );
  OAI22_X1 U311 ( .A1(n326), .A2(n327), .B1(n209), .B2(n328), .ZN(n87) );
  XNOR2_X1 U312 ( .A(a[5]), .B(n296), .ZN(n326) );
  OAI22_X1 U313 ( .A1(n328), .A2(n235), .B1(n210), .B2(n329), .ZN(n86) );
  XNOR2_X1 U314 ( .A(n213), .B(a[5]), .ZN(n328) );
  OAI22_X1 U315 ( .A1(n329), .A2(n236), .B1(n209), .B2(n330), .ZN(n85) );
  XNOR2_X1 U316 ( .A(b[2]), .B(a[5]), .ZN(n329) );
  OAI22_X1 U317 ( .A1(n330), .A2(n236), .B1(n209), .B2(n331), .ZN(n84) );
  XNOR2_X1 U318 ( .A(b[3]), .B(a[5]), .ZN(n330) );
  OAI22_X1 U319 ( .A1(n331), .A2(n235), .B1(n210), .B2(n332), .ZN(n83) );
  XNOR2_X1 U320 ( .A(b[4]), .B(a[5]), .ZN(n331) );
  OAI22_X1 U321 ( .A1(n332), .A2(n236), .B1(n209), .B2(n333), .ZN(n82) );
  XNOR2_X1 U322 ( .A(b[5]), .B(a[5]), .ZN(n332) );
  OAI22_X1 U323 ( .A1(n335), .A2(n209), .B1(n235), .B2(n335), .ZN(n334) );
  NOR2_X1 U324 ( .A1(n336), .A2(n212), .ZN(n80) );
  OAI22_X1 U325 ( .A1(n337), .A2(n338), .B1(n336), .B2(n339), .ZN(n79) );
  XNOR2_X1 U326 ( .A(a[7]), .B(n296), .ZN(n337) );
  OAI22_X1 U327 ( .A1(n340), .A2(n338), .B1(n336), .B2(n341), .ZN(n77) );
  OAI22_X1 U328 ( .A1(n341), .A2(n338), .B1(n336), .B2(n342), .ZN(n76) );
  XNOR2_X1 U329 ( .A(b[3]), .B(a[7]), .ZN(n341) );
  OAI22_X1 U330 ( .A1(n342), .A2(n338), .B1(n336), .B2(n343), .ZN(n75) );
  XNOR2_X1 U331 ( .A(b[4]), .B(a[7]), .ZN(n342) );
  OAI22_X1 U332 ( .A1(n343), .A2(n338), .B1(n336), .B2(n344), .ZN(n74) );
  XNOR2_X1 U333 ( .A(b[5]), .B(a[7]), .ZN(n343) );
  OAI22_X1 U334 ( .A1(n346), .A2(n336), .B1(n338), .B2(n346), .ZN(n345) );
  OAI21_X1 U335 ( .B1(n296), .B2(n308), .A(n311), .ZN(n72) );
  OAI21_X1 U336 ( .B1(n306), .B2(n317), .A(n347), .ZN(n71) );
  OR3_X1 U337 ( .A1(n285), .A2(n296), .A3(n306), .ZN(n347) );
  OAI21_X1 U338 ( .B1(n303), .B2(n327), .A(n348), .ZN(n70) );
  OR3_X1 U339 ( .A1(n210), .A2(n296), .A3(n303), .ZN(n348) );
  OAI21_X1 U340 ( .B1(n300), .B2(n338), .A(n349), .ZN(n69) );
  OR3_X1 U341 ( .A1(n336), .A2(n296), .A3(n300), .ZN(n349) );
  XNOR2_X1 U342 ( .A(n350), .B(n351), .ZN(n38) );
  OR2_X1 U343 ( .A1(n350), .A2(n351), .ZN(n37) );
  OAI22_X1 U344 ( .A1(n322), .A2(n317), .B1(n285), .B2(n352), .ZN(n351) );
  XNOR2_X1 U345 ( .A(b[5]), .B(a[3]), .ZN(n322) );
  OAI22_X1 U346 ( .A1(n339), .A2(n338), .B1(n336), .B2(n340), .ZN(n350) );
  XNOR2_X1 U347 ( .A(b[2]), .B(a[7]), .ZN(n340) );
  XNOR2_X1 U348 ( .A(n232), .B(a[7]), .ZN(n339) );
  OAI22_X1 U349 ( .A1(n352), .A2(n317), .B1(n286), .B2(n324), .ZN(n31) );
  XNOR2_X1 U350 ( .A(b[7]), .B(a[3]), .ZN(n324) );
  XNOR2_X1 U351 ( .A(n306), .B(a[2]), .ZN(n353) );
  XNOR2_X1 U352 ( .A(b[6]), .B(a[3]), .ZN(n352) );
  OAI22_X1 U353 ( .A1(n333), .A2(n236), .B1(n210), .B2(n335), .ZN(n21) );
  XNOR2_X1 U354 ( .A(b[7]), .B(a[5]), .ZN(n335) );
  XNOR2_X1 U355 ( .A(n303), .B(a[4]), .ZN(n354) );
  XNOR2_X1 U356 ( .A(b[6]), .B(a[5]), .ZN(n333) );
  XNOR2_X1 U357 ( .A(b[7]), .B(a[7]), .ZN(n346) );
  NAND2_X1 U358 ( .A1(n336), .A2(n355), .ZN(n338) );
  XNOR2_X1 U359 ( .A(n300), .B(a[6]), .ZN(n355) );
  XNOR2_X1 U360 ( .A(b[6]), .B(a[7]), .ZN(n344) );
  OAI22_X1 U361 ( .A1(n296), .A2(n311), .B1(n356), .B2(n309), .ZN(n104) );
  OAI22_X1 U362 ( .A1(n356), .A2(n311), .B1(n357), .B2(n309), .ZN(n103) );
  XNOR2_X1 U363 ( .A(b[1]), .B(a[1]), .ZN(n356) );
  OAI22_X1 U364 ( .A1(n357), .A2(n311), .B1(n358), .B2(n309), .ZN(n102) );
  XNOR2_X1 U365 ( .A(b[2]), .B(a[1]), .ZN(n357) );
  OAI22_X1 U366 ( .A1(n358), .A2(n311), .B1(n359), .B2(n309), .ZN(n101) );
  XNOR2_X1 U367 ( .A(b[3]), .B(a[1]), .ZN(n358) );
  OAI22_X1 U368 ( .A1(n359), .A2(n311), .B1(n310), .B2(n309), .ZN(n100) );
  XNOR2_X1 U369 ( .A(b[5]), .B(n211), .ZN(n310) );
  NAND2_X1 U370 ( .A1(a[1]), .A2(n309), .ZN(n311) );
  XNOR2_X1 U371 ( .A(b[4]), .B(n211), .ZN(n359) );
endmodule


module mac_15 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_15_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_15_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_14_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74;
  wire   [15:1] carry;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n1) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
  XOR2_X1 U3 ( .A(B[15]), .B(A[15]), .Z(n3) );
  XOR2_X1 U4 ( .A(carry[15]), .B(n3), .Z(SUM[15]) );
  AND2_X1 U5 ( .A1(B[0]), .A2(A[0]), .ZN(n74) );
  NAND2_X1 U6 ( .A1(carry[12]), .A2(A[12]), .ZN(n4) );
  NAND3_X1 U7 ( .A1(n9), .A2(n10), .A3(n11), .ZN(n5) );
  NAND3_X1 U8 ( .A1(n9), .A2(n10), .A3(n11), .ZN(n6) );
  NAND3_X1 U9 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n7) );
  XOR2_X1 U10 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR2_X1 U11 ( .A(carry[5]), .B(n8), .Z(SUM[5]) );
  NAND2_X1 U12 ( .A1(carry[5]), .A2(B[5]), .ZN(n9) );
  NAND2_X1 U13 ( .A1(carry[5]), .A2(A[5]), .ZN(n10) );
  NAND2_X1 U14 ( .A1(B[5]), .A2(A[5]), .ZN(n11) );
  NAND3_X1 U15 ( .A1(n9), .A2(n10), .A3(n11), .ZN(carry[6]) );
  NAND3_X1 U16 ( .A1(n15), .A2(n14), .A3(n16), .ZN(n12) );
  XOR2_X1 U17 ( .A(B[6]), .B(A[6]), .Z(n13) );
  XOR2_X1 U18 ( .A(n6), .B(n13), .Z(SUM[6]) );
  NAND2_X1 U19 ( .A1(n5), .A2(B[6]), .ZN(n14) );
  NAND2_X1 U20 ( .A1(carry[6]), .A2(A[6]), .ZN(n15) );
  NAND2_X1 U21 ( .A1(B[6]), .A2(A[6]), .ZN(n16) );
  NAND3_X1 U22 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[7]) );
  NAND3_X1 U23 ( .A1(n38), .A2(n4), .A3(n40), .ZN(n17) );
  NAND3_X1 U24 ( .A1(n38), .A2(n4), .A3(n40), .ZN(n18) );
  NAND3_X1 U25 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n19) );
  NAND3_X1 U26 ( .A1(n25), .A2(n24), .A3(n26), .ZN(n20) );
  NAND3_X1 U27 ( .A1(n72), .A2(n71), .A3(n73), .ZN(n21) );
  NAND3_X1 U28 ( .A1(n49), .A2(n48), .A3(n50), .ZN(n22) );
  XOR2_X1 U29 ( .A(B[7]), .B(A[7]), .Z(n23) );
  XOR2_X1 U30 ( .A(carry[7]), .B(n23), .Z(SUM[7]) );
  NAND2_X1 U31 ( .A1(n12), .A2(B[7]), .ZN(n24) );
  NAND2_X1 U32 ( .A1(carry[7]), .A2(A[7]), .ZN(n25) );
  NAND2_X1 U33 ( .A1(B[7]), .A2(A[7]), .ZN(n26) );
  NAND3_X1 U34 ( .A1(n25), .A2(n24), .A3(n26), .ZN(carry[8]) );
  XOR2_X1 U35 ( .A(B[13]), .B(A[13]), .Z(n27) );
  XOR2_X1 U36 ( .A(n18), .B(n27), .Z(SUM[13]) );
  NAND2_X1 U37 ( .A1(n17), .A2(B[13]), .ZN(n28) );
  NAND2_X1 U38 ( .A1(carry[13]), .A2(A[13]), .ZN(n29) );
  NAND2_X1 U39 ( .A1(B[13]), .A2(A[13]), .ZN(n30) );
  NAND3_X1 U40 ( .A1(n28), .A2(n29), .A3(n30), .ZN(carry[14]) );
  XOR2_X1 U41 ( .A(B[3]), .B(A[3]), .Z(n31) );
  XOR2_X1 U42 ( .A(n21), .B(n31), .Z(SUM[3]) );
  NAND2_X1 U43 ( .A1(n21), .A2(B[3]), .ZN(n32) );
  NAND2_X1 U44 ( .A1(carry[3]), .A2(A[3]), .ZN(n33) );
  NAND2_X1 U45 ( .A1(B[3]), .A2(A[3]), .ZN(n34) );
  NAND3_X1 U46 ( .A1(n32), .A2(n33), .A3(n34), .ZN(carry[4]) );
  NAND3_X1 U47 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n35) );
  NAND3_X1 U48 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n36) );
  XOR2_X1 U49 ( .A(B[12]), .B(A[12]), .Z(n37) );
  XOR2_X1 U50 ( .A(n36), .B(n37), .Z(SUM[12]) );
  NAND2_X1 U51 ( .A1(n35), .A2(B[12]), .ZN(n38) );
  NAND2_X1 U52 ( .A1(carry[12]), .A2(A[12]), .ZN(n39) );
  NAND2_X1 U53 ( .A1(B[12]), .A2(A[12]), .ZN(n40) );
  NAND3_X1 U54 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[13]) );
  XOR2_X1 U55 ( .A(B[14]), .B(A[14]), .Z(n41) );
  XOR2_X1 U56 ( .A(n19), .B(n41), .Z(SUM[14]) );
  NAND2_X1 U57 ( .A1(n19), .A2(B[14]), .ZN(n42) );
  NAND2_X1 U58 ( .A1(carry[14]), .A2(A[14]), .ZN(n43) );
  NAND2_X1 U59 ( .A1(B[14]), .A2(A[14]), .ZN(n44) );
  NAND3_X1 U60 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[15]) );
  NAND3_X1 U61 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n45) );
  NAND3_X1 U62 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n46) );
  XOR2_X1 U63 ( .A(B[10]), .B(A[10]), .Z(n47) );
  XOR2_X1 U64 ( .A(n46), .B(n47), .Z(SUM[10]) );
  NAND2_X1 U65 ( .A1(n45), .A2(B[10]), .ZN(n48) );
  NAND2_X1 U66 ( .A1(carry[10]), .A2(A[10]), .ZN(n49) );
  NAND2_X1 U67 ( .A1(B[10]), .A2(A[10]), .ZN(n50) );
  XOR2_X1 U68 ( .A(B[11]), .B(A[11]), .Z(n51) );
  XOR2_X1 U69 ( .A(n7), .B(n51), .Z(SUM[11]) );
  NAND2_X1 U70 ( .A1(n7), .A2(B[11]), .ZN(n52) );
  NAND2_X1 U71 ( .A1(n22), .A2(A[11]), .ZN(n53) );
  NAND2_X1 U72 ( .A1(B[11]), .A2(A[11]), .ZN(n54) );
  NAND3_X1 U73 ( .A1(n52), .A2(n53), .A3(n54), .ZN(carry[12]) );
  NAND3_X1 U74 ( .A1(n67), .A2(n68), .A3(n69), .ZN(n55) );
  NAND3_X1 U75 ( .A1(n67), .A2(n68), .A3(n69), .ZN(n56) );
  NAND3_X1 U76 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n57) );
  XOR2_X1 U77 ( .A(B[8]), .B(A[8]), .Z(n58) );
  XOR2_X1 U78 ( .A(n20), .B(n58), .Z(SUM[8]) );
  NAND2_X1 U79 ( .A1(n20), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U80 ( .A1(carry[8]), .A2(A[8]), .ZN(n60) );
  NAND2_X1 U81 ( .A1(B[8]), .A2(A[8]), .ZN(n61) );
  NAND3_X1 U82 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[9]) );
  XOR2_X1 U83 ( .A(B[9]), .B(A[9]), .Z(n62) );
  XOR2_X1 U84 ( .A(n57), .B(n62), .Z(SUM[9]) );
  NAND2_X1 U85 ( .A1(n57), .A2(B[9]), .ZN(n63) );
  NAND2_X1 U86 ( .A1(carry[9]), .A2(A[9]), .ZN(n64) );
  NAND2_X1 U87 ( .A1(B[9]), .A2(A[9]), .ZN(n65) );
  NAND3_X1 U88 ( .A1(n63), .A2(n64), .A3(n65), .ZN(carry[10]) );
  XOR2_X1 U89 ( .A(B[1]), .B(A[1]), .Z(n66) );
  XOR2_X1 U90 ( .A(n2), .B(n66), .Z(SUM[1]) );
  NAND2_X1 U91 ( .A1(n1), .A2(B[1]), .ZN(n67) );
  NAND2_X1 U92 ( .A1(n74), .A2(A[1]), .ZN(n68) );
  NAND2_X1 U93 ( .A1(B[1]), .A2(A[1]), .ZN(n69) );
  NAND3_X1 U94 ( .A1(n67), .A2(n68), .A3(n69), .ZN(carry[2]) );
  XOR2_X1 U95 ( .A(B[2]), .B(A[2]), .Z(n70) );
  XOR2_X1 U96 ( .A(n56), .B(n70), .Z(SUM[2]) );
  NAND2_X1 U97 ( .A1(n55), .A2(B[2]), .ZN(n71) );
  NAND2_X1 U98 ( .A1(carry[2]), .A2(A[2]), .ZN(n72) );
  NAND2_X1 U99 ( .A1(B[2]), .A2(A[2]), .ZN(n73) );
  NAND3_X1 U100 ( .A1(n71), .A2(n72), .A3(n73), .ZN(carry[3]) );
  XOR2_X1 U101 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_14_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n305), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n304), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n308), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n307), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n310), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  INV_X2 U157 ( .A(n300), .ZN(n299) );
  AND2_X1 U158 ( .A1(n207), .A2(n102), .ZN(n206) );
  CLKBUF_X1 U159 ( .A(n216), .Z(n207) );
  XOR2_X1 U160 ( .A(a[3]), .B(a[2]), .Z(n356) );
  CLKBUF_X1 U161 ( .A(a[1]), .Z(n208) );
  NAND2_X1 U162 ( .A1(n7), .A2(n28), .ZN(n209) );
  CLKBUF_X1 U163 ( .A(n11), .Z(n210) );
  AND2_X1 U164 ( .A1(n104), .A2(n72), .ZN(n211) );
  BUF_X1 U165 ( .A(n328), .Z(n212) );
  BUF_X2 U166 ( .A(n328), .Z(n213) );
  XNOR2_X1 U167 ( .A(a[4]), .B(a[3]), .ZN(n328) );
  NAND3_X1 U168 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n214) );
  CLKBUF_X1 U169 ( .A(n209), .Z(n215) );
  XOR2_X1 U170 ( .A(n216), .B(n102), .Z(n56) );
  OAI22_X1 U171 ( .A1(n319), .A2(n320), .B1(n289), .B2(n321), .ZN(n216) );
  XOR2_X2 U172 ( .A(a[6]), .B(n306), .Z(n339) );
  CLKBUF_X1 U173 ( .A(n50), .Z(n217) );
  NAND3_X1 U174 ( .A1(n209), .A2(n275), .A3(n277), .ZN(n218) );
  NAND3_X1 U175 ( .A1(n285), .A2(n284), .A3(n283), .ZN(n219) );
  NAND3_X1 U176 ( .A1(n230), .A2(n229), .A3(n231), .ZN(n220) );
  CLKBUF_X1 U177 ( .A(n271), .Z(n221) );
  CLKBUF_X1 U178 ( .A(n254), .Z(n222) );
  CLKBUF_X1 U179 ( .A(n238), .Z(n223) );
  CLKBUF_X1 U180 ( .A(n285), .Z(n224) );
  NAND3_X1 U181 ( .A1(n248), .A2(n247), .A3(n249), .ZN(n225) );
  NAND3_X1 U182 ( .A1(n276), .A2(n275), .A3(n277), .ZN(n226) );
  CLKBUF_X1 U183 ( .A(n56), .Z(n227) );
  XOR2_X1 U184 ( .A(n27), .B(n24), .Z(n228) );
  XOR2_X1 U185 ( .A(n6), .B(n228), .Z(product[10]) );
  NAND2_X1 U186 ( .A1(n226), .A2(n27), .ZN(n229) );
  NAND2_X1 U187 ( .A1(n218), .A2(n24), .ZN(n230) );
  NAND2_X1 U188 ( .A1(n27), .A2(n24), .ZN(n231) );
  NAND3_X1 U189 ( .A1(n230), .A2(n229), .A3(n231), .ZN(n5) );
  NAND3_X1 U190 ( .A1(n267), .A2(n268), .A3(n269), .ZN(n232) );
  XNOR2_X1 U191 ( .A(b[1]), .B(n208), .ZN(n233) );
  NAND3_X1 U192 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n234) );
  CLKBUF_X1 U193 ( .A(n284), .Z(n235) );
  NAND3_X1 U194 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n236) );
  NAND3_X1 U195 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n237) );
  NAND3_X1 U196 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n238) );
  CLKBUF_X1 U197 ( .A(n7), .Z(n239) );
  NAND3_X1 U198 ( .A1(n244), .A2(n245), .A3(n243), .ZN(n240) );
  NAND3_X1 U199 ( .A1(n224), .A2(n235), .A3(n283), .ZN(n241) );
  XOR2_X1 U200 ( .A(n103), .B(n96), .Z(n242) );
  XOR2_X1 U201 ( .A(n242), .B(n211), .Z(product[2]) );
  NAND2_X1 U202 ( .A1(n103), .A2(n96), .ZN(n243) );
  NAND2_X1 U203 ( .A1(n103), .A2(n14), .ZN(n244) );
  NAND2_X1 U204 ( .A1(n96), .A2(n211), .ZN(n245) );
  NAND3_X1 U205 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n13) );
  XOR2_X1 U206 ( .A(n227), .B(n71), .Z(n246) );
  XOR2_X1 U207 ( .A(n246), .B(n240), .Z(product[3]) );
  NAND2_X1 U208 ( .A1(n56), .A2(n71), .ZN(n247) );
  NAND2_X1 U209 ( .A1(n56), .A2(n240), .ZN(n248) );
  NAND2_X1 U210 ( .A1(n71), .A2(n13), .ZN(n249) );
  NAND3_X1 U211 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n12) );
  XOR2_X1 U212 ( .A(n54), .B(n206), .Z(n250) );
  XOR2_X1 U213 ( .A(n12), .B(n250), .Z(product[4]) );
  NAND2_X1 U214 ( .A1(n225), .A2(n54), .ZN(n251) );
  NAND2_X1 U215 ( .A1(n225), .A2(n206), .ZN(n252) );
  NAND2_X1 U216 ( .A1(n54), .A2(n206), .ZN(n253) );
  NAND3_X1 U217 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n11) );
  NAND3_X1 U218 ( .A1(n256), .A2(n258), .A3(n257), .ZN(n254) );
  XOR2_X1 U219 ( .A(n217), .B(n53), .Z(n255) );
  XOR2_X1 U220 ( .A(n210), .B(n255), .Z(product[5]) );
  NAND2_X1 U221 ( .A1(n11), .A2(n50), .ZN(n256) );
  NAND2_X1 U222 ( .A1(n237), .A2(n53), .ZN(n257) );
  NAND2_X1 U223 ( .A1(n50), .A2(n53), .ZN(n258) );
  NAND3_X1 U224 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n10) );
  CLKBUF_X1 U225 ( .A(b[1]), .Z(n259) );
  XOR2_X1 U226 ( .A(n34), .B(n39), .Z(n260) );
  XOR2_X1 U227 ( .A(n8), .B(n260), .Z(product[8]) );
  NAND2_X1 U228 ( .A1(n236), .A2(n34), .ZN(n261) );
  NAND2_X1 U229 ( .A1(n214), .A2(n39), .ZN(n262) );
  NAND2_X1 U230 ( .A1(n34), .A2(n39), .ZN(n263) );
  NAND3_X1 U231 ( .A1(n262), .A2(n261), .A3(n263), .ZN(n7) );
  CLKBUF_X1 U232 ( .A(n220), .Z(n264) );
  CLKBUF_X1 U233 ( .A(n232), .Z(n265) );
  XOR2_X1 U234 ( .A(n46), .B(n49), .Z(n266) );
  XOR2_X1 U235 ( .A(n222), .B(n266), .Z(product[6]) );
  NAND2_X1 U236 ( .A1(n254), .A2(n46), .ZN(n267) );
  NAND2_X1 U237 ( .A1(n10), .A2(n49), .ZN(n268) );
  NAND2_X1 U238 ( .A1(n46), .A2(n49), .ZN(n269) );
  NAND3_X1 U239 ( .A1(n267), .A2(n268), .A3(n269), .ZN(n9) );
  XOR2_X1 U240 ( .A(n40), .B(n45), .Z(n270) );
  XOR2_X1 U241 ( .A(n265), .B(n270), .Z(product[7]) );
  NAND2_X1 U242 ( .A1(n232), .A2(n40), .ZN(n271) );
  NAND2_X1 U243 ( .A1(n9), .A2(n45), .ZN(n272) );
  NAND2_X1 U244 ( .A1(n40), .A2(n45), .ZN(n273) );
  NAND3_X1 U245 ( .A1(n221), .A2(n272), .A3(n273), .ZN(n8) );
  XOR2_X1 U246 ( .A(n33), .B(n28), .Z(n274) );
  XOR2_X1 U247 ( .A(n239), .B(n274), .Z(product[9]) );
  NAND2_X1 U248 ( .A1(n234), .A2(n33), .ZN(n275) );
  NAND2_X1 U249 ( .A1(n7), .A2(n28), .ZN(n276) );
  NAND2_X1 U250 ( .A1(n33), .A2(n28), .ZN(n277) );
  NAND3_X1 U251 ( .A1(n275), .A2(n215), .A3(n277), .ZN(n6) );
  XOR2_X1 U252 ( .A(n20), .B(n23), .Z(n278) );
  XOR2_X1 U253 ( .A(n278), .B(n264), .Z(product[11]) );
  NAND2_X1 U254 ( .A1(n20), .A2(n23), .ZN(n279) );
  NAND2_X1 U255 ( .A1(n20), .A2(n220), .ZN(n280) );
  NAND2_X1 U256 ( .A1(n23), .A2(n5), .ZN(n281) );
  NAND3_X1 U257 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n4) );
  XOR2_X1 U258 ( .A(n19), .B(n18), .Z(n282) );
  XOR2_X1 U259 ( .A(n282), .B(n223), .Z(product[12]) );
  NAND2_X1 U260 ( .A1(n19), .A2(n18), .ZN(n283) );
  NAND2_X1 U261 ( .A1(n19), .A2(n4), .ZN(n284) );
  NAND2_X1 U262 ( .A1(n238), .A2(n18), .ZN(n285) );
  NAND3_X1 U263 ( .A1(n285), .A2(n284), .A3(n283), .ZN(n3) );
  NAND2_X2 U264 ( .A1(n318), .A2(n356), .ZN(n320) );
  NAND2_X2 U265 ( .A1(n212), .A2(n357), .ZN(n330) );
  NAND3_X1 U266 ( .A1(n293), .A2(n294), .A3(n292), .ZN(n286) );
  NAND3_X1 U267 ( .A1(n293), .A2(n292), .A3(n294), .ZN(n287) );
  XOR2_X1 U268 ( .A(a[2]), .B(n311), .Z(n288) );
  XOR2_X1 U269 ( .A(a[2]), .B(n311), .Z(n289) );
  INV_X1 U270 ( .A(n15), .ZN(n301) );
  AND3_X1 U271 ( .A1(n296), .A2(n297), .A3(n298), .ZN(product[15]) );
  INV_X1 U272 ( .A(n348), .ZN(n302) );
  INV_X1 U273 ( .A(n21), .ZN(n304) );
  INV_X1 U274 ( .A(n337), .ZN(n305) );
  INV_X1 U275 ( .A(n317), .ZN(n310) );
  INV_X1 U276 ( .A(n326), .ZN(n308) );
  INV_X1 U277 ( .A(n31), .ZN(n307) );
  INV_X1 U278 ( .A(b[0]), .ZN(n300) );
  XOR2_X1 U279 ( .A(a[2]), .B(n311), .Z(n318) );
  INV_X1 U280 ( .A(a[0]), .ZN(n312) );
  INV_X1 U281 ( .A(a[5]), .ZN(n306) );
  INV_X1 U282 ( .A(a[7]), .ZN(n303) );
  INV_X1 U283 ( .A(a[3]), .ZN(n309) );
  XOR2_X1 U284 ( .A(n17), .B(n301), .Z(n291) );
  XOR2_X1 U285 ( .A(n291), .B(n241), .Z(product[13]) );
  NAND2_X1 U286 ( .A1(n17), .A2(n301), .ZN(n292) );
  NAND2_X1 U287 ( .A1(n17), .A2(n3), .ZN(n293) );
  NAND2_X1 U288 ( .A1(n301), .A2(n219), .ZN(n294) );
  XOR2_X1 U289 ( .A(n302), .B(n15), .Z(n295) );
  XOR2_X1 U290 ( .A(n295), .B(n287), .Z(product[14]) );
  NAND2_X1 U291 ( .A1(n302), .A2(n15), .ZN(n296) );
  NAND2_X1 U292 ( .A1(n286), .A2(n302), .ZN(n297) );
  NAND2_X1 U293 ( .A1(n286), .A2(n15), .ZN(n298) );
  INV_X1 U294 ( .A(a[1]), .ZN(n311) );
  NOR2_X1 U295 ( .A1(n312), .A2(n300), .ZN(product[0]) );
  OAI22_X1 U296 ( .A1(n313), .A2(n314), .B1(n315), .B2(n312), .ZN(n99) );
  OAI22_X1 U297 ( .A1(n315), .A2(n314), .B1(n316), .B2(n312), .ZN(n98) );
  XNOR2_X1 U298 ( .A(b[6]), .B(n208), .ZN(n315) );
  OAI22_X1 U299 ( .A1(n312), .A2(n316), .B1(n314), .B2(n316), .ZN(n317) );
  XNOR2_X1 U300 ( .A(b[7]), .B(n208), .ZN(n316) );
  NOR2_X1 U301 ( .A1(n288), .A2(n300), .ZN(n96) );
  XNOR2_X1 U302 ( .A(a[3]), .B(n299), .ZN(n319) );
  OAI22_X1 U303 ( .A1(n321), .A2(n320), .B1(n289), .B2(n322), .ZN(n94) );
  XNOR2_X1 U304 ( .A(b[1]), .B(a[3]), .ZN(n321) );
  OAI22_X1 U305 ( .A1(n322), .A2(n320), .B1(n288), .B2(n323), .ZN(n93) );
  XNOR2_X1 U306 ( .A(b[2]), .B(a[3]), .ZN(n322) );
  OAI22_X1 U307 ( .A1(n323), .A2(n320), .B1(n289), .B2(n324), .ZN(n92) );
  XNOR2_X1 U308 ( .A(b[3]), .B(a[3]), .ZN(n323) );
  OAI22_X1 U309 ( .A1(n324), .A2(n320), .B1(n289), .B2(n325), .ZN(n91) );
  XNOR2_X1 U310 ( .A(b[4]), .B(a[3]), .ZN(n324) );
  OAI22_X1 U311 ( .A1(n327), .A2(n288), .B1(n320), .B2(n327), .ZN(n326) );
  NOR2_X1 U312 ( .A1(n213), .A2(n300), .ZN(n88) );
  OAI22_X1 U313 ( .A1(n329), .A2(n330), .B1(n213), .B2(n331), .ZN(n87) );
  XNOR2_X1 U314 ( .A(a[5]), .B(n299), .ZN(n329) );
  OAI22_X1 U315 ( .A1(n331), .A2(n330), .B1(n213), .B2(n332), .ZN(n86) );
  XNOR2_X1 U316 ( .A(b[1]), .B(a[5]), .ZN(n331) );
  OAI22_X1 U317 ( .A1(n332), .A2(n330), .B1(n213), .B2(n333), .ZN(n85) );
  XNOR2_X1 U318 ( .A(b[2]), .B(a[5]), .ZN(n332) );
  OAI22_X1 U319 ( .A1(n333), .A2(n330), .B1(n213), .B2(n334), .ZN(n84) );
  XNOR2_X1 U320 ( .A(b[3]), .B(a[5]), .ZN(n333) );
  OAI22_X1 U321 ( .A1(n334), .A2(n330), .B1(n213), .B2(n335), .ZN(n83) );
  XNOR2_X1 U322 ( .A(b[4]), .B(a[5]), .ZN(n334) );
  OAI22_X1 U323 ( .A1(n335), .A2(n330), .B1(n213), .B2(n336), .ZN(n82) );
  XNOR2_X1 U324 ( .A(b[5]), .B(a[5]), .ZN(n335) );
  OAI22_X1 U325 ( .A1(n338), .A2(n213), .B1(n330), .B2(n338), .ZN(n337) );
  NOR2_X1 U326 ( .A1(n339), .A2(n300), .ZN(n80) );
  OAI22_X1 U327 ( .A1(n340), .A2(n341), .B1(n339), .B2(n342), .ZN(n79) );
  XNOR2_X1 U328 ( .A(a[7]), .B(n299), .ZN(n340) );
  OAI22_X1 U329 ( .A1(n343), .A2(n341), .B1(n339), .B2(n344), .ZN(n77) );
  OAI22_X1 U330 ( .A1(n344), .A2(n341), .B1(n339), .B2(n345), .ZN(n76) );
  XNOR2_X1 U331 ( .A(b[3]), .B(a[7]), .ZN(n344) );
  OAI22_X1 U332 ( .A1(n345), .A2(n341), .B1(n339), .B2(n346), .ZN(n75) );
  XNOR2_X1 U333 ( .A(b[4]), .B(a[7]), .ZN(n345) );
  OAI22_X1 U334 ( .A1(n346), .A2(n341), .B1(n339), .B2(n347), .ZN(n74) );
  XNOR2_X1 U335 ( .A(b[5]), .B(a[7]), .ZN(n346) );
  OAI22_X1 U336 ( .A1(n349), .A2(n339), .B1(n341), .B2(n349), .ZN(n348) );
  OAI21_X1 U337 ( .B1(n299), .B2(n311), .A(n314), .ZN(n72) );
  OAI21_X1 U338 ( .B1(n309), .B2(n320), .A(n350), .ZN(n71) );
  OR3_X1 U339 ( .A1(n288), .A2(n299), .A3(n309), .ZN(n350) );
  OAI21_X1 U340 ( .B1(n306), .B2(n330), .A(n351), .ZN(n70) );
  OR3_X1 U341 ( .A1(n213), .A2(n299), .A3(n306), .ZN(n351) );
  OAI21_X1 U342 ( .B1(n303), .B2(n341), .A(n352), .ZN(n69) );
  OR3_X1 U343 ( .A1(n339), .A2(n299), .A3(n303), .ZN(n352) );
  XNOR2_X1 U344 ( .A(n353), .B(n354), .ZN(n38) );
  OR2_X1 U345 ( .A1(n353), .A2(n354), .ZN(n37) );
  OAI22_X1 U346 ( .A1(n325), .A2(n320), .B1(n288), .B2(n355), .ZN(n354) );
  XNOR2_X1 U347 ( .A(b[5]), .B(a[3]), .ZN(n325) );
  OAI22_X1 U348 ( .A1(n342), .A2(n341), .B1(n339), .B2(n343), .ZN(n353) );
  XNOR2_X1 U349 ( .A(b[2]), .B(a[7]), .ZN(n343) );
  XNOR2_X1 U350 ( .A(n259), .B(a[7]), .ZN(n342) );
  OAI22_X1 U351 ( .A1(n355), .A2(n320), .B1(n289), .B2(n327), .ZN(n31) );
  XNOR2_X1 U352 ( .A(b[7]), .B(a[3]), .ZN(n327) );
  XNOR2_X1 U353 ( .A(b[6]), .B(a[3]), .ZN(n355) );
  OAI22_X1 U354 ( .A1(n336), .A2(n330), .B1(n213), .B2(n338), .ZN(n21) );
  XNOR2_X1 U355 ( .A(b[7]), .B(a[5]), .ZN(n338) );
  XNOR2_X1 U356 ( .A(n306), .B(a[4]), .ZN(n357) );
  XNOR2_X1 U357 ( .A(b[6]), .B(a[5]), .ZN(n336) );
  OAI22_X1 U358 ( .A1(n347), .A2(n341), .B1(n339), .B2(n349), .ZN(n15) );
  XNOR2_X1 U359 ( .A(b[7]), .B(a[7]), .ZN(n349) );
  NAND2_X1 U360 ( .A1(n339), .A2(n358), .ZN(n341) );
  XNOR2_X1 U361 ( .A(n303), .B(a[6]), .ZN(n358) );
  XNOR2_X1 U362 ( .A(b[6]), .B(a[7]), .ZN(n347) );
  OAI22_X1 U363 ( .A1(n299), .A2(n314), .B1(n359), .B2(n312), .ZN(n104) );
  OAI22_X1 U364 ( .A1(n233), .A2(n314), .B1(n360), .B2(n312), .ZN(n103) );
  XNOR2_X1 U365 ( .A(b[1]), .B(a[1]), .ZN(n359) );
  OAI22_X1 U366 ( .A1(n360), .A2(n314), .B1(n361), .B2(n312), .ZN(n102) );
  XNOR2_X1 U367 ( .A(b[2]), .B(a[1]), .ZN(n360) );
  OAI22_X1 U368 ( .A1(n361), .A2(n314), .B1(n362), .B2(n312), .ZN(n101) );
  XNOR2_X1 U369 ( .A(b[3]), .B(a[1]), .ZN(n361) );
  OAI22_X1 U370 ( .A1(n362), .A2(n314), .B1(n313), .B2(n312), .ZN(n100) );
  XNOR2_X1 U371 ( .A(b[5]), .B(n208), .ZN(n313) );
  NAND2_X1 U372 ( .A1(a[1]), .A2(n312), .ZN(n314) );
  XNOR2_X1 U373 ( .A(b[4]), .B(n208), .ZN(n362) );
endmodule


module mac_14 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_14_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_14_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X2 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_13_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66;
  wire   [15:1] carry;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n66) );
  CLKBUF_X1 U2 ( .A(carry[11]), .Z(n1) );
  NAND3_X1 U3 ( .A1(n6), .A2(n7), .A3(n8), .ZN(n2) );
  XNOR2_X1 U4 ( .A(B[15]), .B(A[15]), .ZN(n3) );
  CLKBUF_X1 U5 ( .A(carry[12]), .Z(n4) );
  XNOR2_X1 U6 ( .A(carry[15]), .B(n3), .ZN(SUM[15]) );
  XOR2_X1 U7 ( .A(B[11]), .B(A[11]), .Z(n5) );
  XOR2_X1 U8 ( .A(n1), .B(n5), .Z(SUM[11]) );
  NAND2_X1 U9 ( .A1(carry[11]), .A2(B[11]), .ZN(n6) );
  NAND2_X1 U10 ( .A1(carry[11]), .A2(A[11]), .ZN(n7) );
  NAND2_X1 U11 ( .A1(B[11]), .A2(A[11]), .ZN(n8) );
  NAND3_X1 U12 ( .A1(n6), .A2(n7), .A3(n8), .ZN(carry[12]) );
  XOR2_X1 U13 ( .A(B[9]), .B(A[9]), .Z(n9) );
  XOR2_X1 U14 ( .A(carry[9]), .B(n9), .Z(SUM[9]) );
  NAND2_X1 U15 ( .A1(carry[9]), .A2(B[9]), .ZN(n10) );
  NAND2_X1 U16 ( .A1(carry[9]), .A2(A[9]), .ZN(n11) );
  NAND2_X1 U17 ( .A1(B[9]), .A2(A[9]), .ZN(n12) );
  NAND3_X1 U18 ( .A1(n10), .A2(n11), .A3(n12), .ZN(carry[10]) );
  NAND3_X1 U19 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n13) );
  NAND3_X1 U20 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n14) );
  NAND3_X1 U21 ( .A1(n23), .A2(n24), .A3(n25), .ZN(n15) );
  NAND3_X1 U22 ( .A1(n23), .A2(n24), .A3(n25), .ZN(n16) );
  NAND3_X1 U23 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n17) );
  XOR2_X1 U24 ( .A(B[3]), .B(A[3]), .Z(n18) );
  XOR2_X1 U25 ( .A(n17), .B(n18), .Z(SUM[3]) );
  NAND2_X1 U26 ( .A1(n17), .A2(B[3]), .ZN(n19) );
  NAND2_X1 U27 ( .A1(carry[3]), .A2(A[3]), .ZN(n20) );
  NAND2_X1 U28 ( .A1(B[3]), .A2(A[3]), .ZN(n21) );
  NAND3_X1 U29 ( .A1(n19), .A2(n20), .A3(n21), .ZN(carry[4]) );
  XOR2_X1 U30 ( .A(B[1]), .B(A[1]), .Z(n22) );
  XOR2_X1 U31 ( .A(n66), .B(n22), .Z(SUM[1]) );
  NAND2_X1 U32 ( .A1(n66), .A2(B[1]), .ZN(n23) );
  NAND2_X1 U33 ( .A1(n66), .A2(A[1]), .ZN(n24) );
  NAND2_X1 U34 ( .A1(B[1]), .A2(A[1]), .ZN(n25) );
  NAND3_X1 U35 ( .A1(n23), .A2(n24), .A3(n25), .ZN(carry[2]) );
  XOR2_X1 U36 ( .A(B[2]), .B(A[2]), .Z(n26) );
  XOR2_X1 U37 ( .A(n16), .B(n26), .Z(SUM[2]) );
  NAND2_X1 U38 ( .A1(n15), .A2(B[2]), .ZN(n27) );
  NAND2_X1 U39 ( .A1(carry[2]), .A2(A[2]), .ZN(n28) );
  NAND2_X1 U40 ( .A1(B[2]), .A2(A[2]), .ZN(n29) );
  NAND3_X1 U41 ( .A1(n27), .A2(n28), .A3(n29), .ZN(carry[3]) );
  NAND3_X1 U42 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n30) );
  NAND3_X1 U43 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n31) );
  XOR2_X1 U44 ( .A(B[8]), .B(A[8]), .Z(n32) );
  XOR2_X1 U45 ( .A(n31), .B(n32), .Z(SUM[8]) );
  NAND2_X1 U46 ( .A1(n30), .A2(B[8]), .ZN(n33) );
  NAND2_X1 U47 ( .A1(carry[8]), .A2(A[8]), .ZN(n34) );
  NAND2_X1 U48 ( .A1(B[8]), .A2(A[8]), .ZN(n35) );
  NAND3_X1 U49 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[9]) );
  XOR2_X1 U50 ( .A(B[10]), .B(A[10]), .Z(n36) );
  XOR2_X1 U51 ( .A(carry[10]), .B(n36), .Z(SUM[10]) );
  NAND2_X1 U52 ( .A1(carry[10]), .A2(B[10]), .ZN(n37) );
  NAND2_X1 U53 ( .A1(carry[10]), .A2(A[10]), .ZN(n38) );
  NAND2_X1 U54 ( .A1(B[10]), .A2(A[10]), .ZN(n39) );
  NAND3_X1 U55 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[11]) );
  XOR2_X1 U56 ( .A(B[12]), .B(A[12]), .Z(n40) );
  XOR2_X1 U57 ( .A(n4), .B(n40), .Z(SUM[12]) );
  NAND2_X1 U58 ( .A1(n2), .A2(B[12]), .ZN(n41) );
  NAND2_X1 U59 ( .A1(carry[12]), .A2(A[12]), .ZN(n42) );
  NAND2_X1 U60 ( .A1(B[12]), .A2(A[12]), .ZN(n43) );
  NAND3_X1 U61 ( .A1(n41), .A2(n42), .A3(n43), .ZN(carry[13]) );
  XOR2_X1 U62 ( .A(B[5]), .B(A[5]), .Z(n44) );
  XOR2_X1 U63 ( .A(carry[5]), .B(n44), .Z(SUM[5]) );
  NAND2_X1 U64 ( .A1(carry[5]), .A2(B[5]), .ZN(n45) );
  NAND2_X1 U65 ( .A1(carry[5]), .A2(A[5]), .ZN(n46) );
  NAND2_X1 U66 ( .A1(B[5]), .A2(A[5]), .ZN(n47) );
  NAND3_X1 U67 ( .A1(n45), .A2(n46), .A3(n47), .ZN(carry[6]) );
  NAND3_X1 U68 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n48) );
  NAND3_X1 U69 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n49) );
  XOR2_X1 U70 ( .A(B[13]), .B(A[13]), .Z(n50) );
  XOR2_X1 U71 ( .A(carry[13]), .B(n50), .Z(SUM[13]) );
  NAND2_X1 U72 ( .A1(n13), .A2(B[13]), .ZN(n51) );
  NAND2_X1 U73 ( .A1(carry[13]), .A2(A[13]), .ZN(n52) );
  NAND2_X1 U74 ( .A1(B[13]), .A2(A[13]), .ZN(n53) );
  NAND3_X1 U75 ( .A1(n51), .A2(n52), .A3(n53), .ZN(carry[14]) );
  XOR2_X1 U76 ( .A(B[6]), .B(A[6]), .Z(n54) );
  XOR2_X1 U77 ( .A(carry[6]), .B(n54), .Z(SUM[6]) );
  NAND2_X1 U78 ( .A1(carry[6]), .A2(B[6]), .ZN(n55) );
  NAND2_X1 U79 ( .A1(n14), .A2(A[6]), .ZN(n56) );
  NAND2_X1 U80 ( .A1(B[6]), .A2(A[6]), .ZN(n57) );
  NAND3_X1 U81 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[7]) );
  XOR2_X1 U82 ( .A(B[14]), .B(A[14]), .Z(n58) );
  XOR2_X1 U83 ( .A(carry[14]), .B(n58), .Z(SUM[14]) );
  NAND2_X1 U84 ( .A1(n48), .A2(B[14]), .ZN(n59) );
  NAND2_X1 U85 ( .A1(n48), .A2(A[14]), .ZN(n60) );
  NAND2_X1 U86 ( .A1(B[14]), .A2(A[14]), .ZN(n61) );
  NAND3_X1 U87 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[15]) );
  XOR2_X1 U88 ( .A(B[7]), .B(A[7]), .Z(n62) );
  XOR2_X1 U89 ( .A(carry[7]), .B(n62), .Z(SUM[7]) );
  NAND2_X1 U90 ( .A1(n49), .A2(B[7]), .ZN(n63) );
  NAND2_X1 U91 ( .A1(n49), .A2(A[7]), .ZN(n64) );
  NAND2_X1 U92 ( .A1(B[7]), .A2(A[7]), .ZN(n65) );
  NAND3_X1 U93 ( .A1(n63), .A2(n64), .A3(n65), .ZN(carry[8]) );
  XOR2_X1 U94 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_13_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18, n19,
         n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76, n77,
         n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94, n95,
         n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n308), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n307), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n311), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n310), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n313), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  INV_X1 U157 ( .A(n15), .ZN(n304) );
  INV_X2 U158 ( .A(n303), .ZN(n302) );
  CLKBUF_X1 U159 ( .A(n56), .Z(n206) );
  CLKBUF_X1 U160 ( .A(n289), .Z(n207) );
  AND2_X1 U161 ( .A1(n95), .A2(n102), .ZN(n208) );
  CLKBUF_X1 U162 ( .A(n251), .Z(n209) );
  CLKBUF_X1 U163 ( .A(n233), .Z(n210) );
  NAND2_X1 U164 ( .A1(n3), .A2(n17), .ZN(n211) );
  CLKBUF_X1 U165 ( .A(b[1]), .Z(n212) );
  CLKBUF_X1 U166 ( .A(b[1]), .Z(n213) );
  CLKBUF_X1 U167 ( .A(b[1]), .Z(n214) );
  NAND3_X1 U168 ( .A1(n266), .A2(n211), .A3(n267), .ZN(n215) );
  CLKBUF_X1 U169 ( .A(n299), .Z(n216) );
  NAND3_X1 U170 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n217) );
  NAND3_X1 U171 ( .A1(n216), .A2(n300), .A3(n301), .ZN(n218) );
  NAND2_X1 U172 ( .A1(n253), .A2(n27), .ZN(n219) );
  CLKBUF_X1 U173 ( .A(n253), .Z(n220) );
  NAND2_X1 U174 ( .A1(a[4]), .A2(a[3]), .ZN(n223) );
  NAND2_X1 U175 ( .A1(n221), .A2(n222), .ZN(n224) );
  NAND2_X2 U176 ( .A1(n223), .A2(n224), .ZN(n331) );
  INV_X1 U177 ( .A(a[4]), .ZN(n221) );
  INV_X1 U178 ( .A(a[3]), .ZN(n222) );
  CLKBUF_X1 U179 ( .A(n219), .Z(n225) );
  CLKBUF_X1 U180 ( .A(n279), .Z(n226) );
  NAND3_X1 U181 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n227) );
  NAND3_X1 U182 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n228) );
  NAND3_X1 U183 ( .A1(n219), .A2(n289), .A3(n290), .ZN(n229) );
  NAND3_X1 U184 ( .A1(n225), .A2(n207), .A3(n290), .ZN(n230) );
  NAND3_X1 U185 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n231) );
  NAND3_X1 U186 ( .A1(n226), .A2(n280), .A3(n281), .ZN(n232) );
  NAND3_X1 U187 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n233) );
  NAND3_X1 U188 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n234) );
  XOR2_X1 U189 ( .A(n40), .B(n45), .Z(n235) );
  XOR2_X1 U190 ( .A(n232), .B(n235), .Z(product[7]) );
  NAND2_X1 U191 ( .A1(n231), .A2(n40), .ZN(n236) );
  NAND2_X1 U192 ( .A1(n9), .A2(n45), .ZN(n237) );
  NAND2_X1 U193 ( .A1(n40), .A2(n45), .ZN(n238) );
  NAND3_X1 U194 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n8) );
  CLKBUF_X1 U195 ( .A(n228), .Z(n239) );
  NAND3_X1 U196 ( .A1(n259), .A2(n258), .A3(n257), .ZN(n240) );
  NAND3_X1 U197 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n241) );
  XOR2_X1 U198 ( .A(n23), .B(n20), .Z(n242) );
  XOR2_X1 U199 ( .A(n230), .B(n242), .Z(product[11]) );
  NAND2_X1 U200 ( .A1(n229), .A2(n23), .ZN(n243) );
  NAND2_X1 U201 ( .A1(n5), .A2(n20), .ZN(n244) );
  NAND2_X1 U202 ( .A1(n23), .A2(n20), .ZN(n245) );
  NAND3_X1 U203 ( .A1(n244), .A2(n243), .A3(n245), .ZN(n4) );
  XOR2_X1 U204 ( .A(n54), .B(n208), .Z(n246) );
  XOR2_X1 U205 ( .A(n227), .B(n246), .Z(product[4]) );
  NAND2_X1 U206 ( .A1(n227), .A2(n54), .ZN(n247) );
  NAND2_X1 U207 ( .A1(n12), .A2(n208), .ZN(n248) );
  NAND2_X1 U208 ( .A1(n54), .A2(n208), .ZN(n249) );
  NAND3_X1 U209 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n11) );
  NAND3_X1 U210 ( .A1(n299), .A2(n300), .A3(n301), .ZN(n250) );
  NAND3_X1 U211 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n251) );
  XNOR2_X1 U212 ( .A(n214), .B(n291), .ZN(n252) );
  NAND3_X1 U213 ( .A1(n284), .A2(n283), .A3(n285), .ZN(n253) );
  NAND3_X1 U214 ( .A1(n266), .A2(n265), .A3(n267), .ZN(n254) );
  NAND3_X1 U215 ( .A1(n211), .A2(n267), .A3(n266), .ZN(n255) );
  NAND2_X2 U216 ( .A1(n331), .A2(n360), .ZN(n333) );
  XOR2_X1 U217 ( .A(n103), .B(n96), .Z(n256) );
  XOR2_X1 U218 ( .A(n256), .B(n14), .Z(product[2]) );
  NAND2_X1 U219 ( .A1(n103), .A2(n96), .ZN(n257) );
  NAND2_X1 U220 ( .A1(n103), .A2(n14), .ZN(n258) );
  NAND2_X1 U221 ( .A1(n96), .A2(n14), .ZN(n259) );
  NAND3_X1 U222 ( .A1(n259), .A2(n258), .A3(n257), .ZN(n13) );
  XOR2_X1 U223 ( .A(n206), .B(n71), .Z(n260) );
  XOR2_X1 U224 ( .A(n260), .B(n241), .Z(product[3]) );
  NAND2_X1 U225 ( .A1(n56), .A2(n71), .ZN(n261) );
  NAND2_X1 U226 ( .A1(n56), .A2(n240), .ZN(n262) );
  NAND2_X1 U227 ( .A1(n71), .A2(n13), .ZN(n263) );
  NAND3_X1 U228 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n12) );
  XOR2_X1 U229 ( .A(n17), .B(n304), .Z(n264) );
  XOR2_X1 U230 ( .A(n218), .B(n264), .Z(product[13]) );
  NAND2_X1 U231 ( .A1(n3), .A2(n17), .ZN(n265) );
  NAND2_X1 U232 ( .A1(n250), .A2(n304), .ZN(n266) );
  NAND2_X1 U233 ( .A1(n17), .A2(n304), .ZN(n267) );
  CLKBUF_X1 U234 ( .A(n7), .Z(n268) );
  XOR2_X1 U235 ( .A(n34), .B(n39), .Z(n269) );
  XOR2_X1 U236 ( .A(n210), .B(n269), .Z(product[8]) );
  NAND2_X1 U237 ( .A1(n233), .A2(n34), .ZN(n270) );
  NAND2_X1 U238 ( .A1(n8), .A2(n39), .ZN(n271) );
  NAND2_X1 U239 ( .A1(n34), .A2(n39), .ZN(n272) );
  NAND3_X1 U240 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n7) );
  XOR2_X1 U241 ( .A(n50), .B(n53), .Z(n273) );
  XOR2_X1 U242 ( .A(n217), .B(n273), .Z(product[5]) );
  NAND2_X1 U243 ( .A1(n217), .A2(n50), .ZN(n274) );
  NAND2_X1 U244 ( .A1(n11), .A2(n53), .ZN(n275) );
  NAND2_X1 U245 ( .A1(n50), .A2(n53), .ZN(n276) );
  NAND3_X1 U246 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n10) );
  NAND3_X1 U247 ( .A1(n283), .A2(n284), .A3(n285), .ZN(n277) );
  XOR2_X1 U248 ( .A(n46), .B(n49), .Z(n278) );
  XOR2_X1 U249 ( .A(n209), .B(n278), .Z(product[6]) );
  NAND2_X1 U250 ( .A1(n251), .A2(n46), .ZN(n279) );
  NAND2_X1 U251 ( .A1(n10), .A2(n49), .ZN(n280) );
  NAND2_X1 U252 ( .A1(n46), .A2(n49), .ZN(n281) );
  NAND3_X1 U253 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n9) );
  XOR2_X1 U254 ( .A(n33), .B(n28), .Z(n282) );
  XOR2_X1 U255 ( .A(n268), .B(n282), .Z(product[9]) );
  NAND2_X1 U256 ( .A1(n234), .A2(n33), .ZN(n283) );
  NAND2_X1 U257 ( .A1(n7), .A2(n28), .ZN(n284) );
  NAND2_X1 U258 ( .A1(n33), .A2(n28), .ZN(n285) );
  INV_X1 U259 ( .A(n302), .ZN(n286) );
  XOR2_X1 U260 ( .A(n27), .B(n24), .Z(n287) );
  XOR2_X1 U261 ( .A(n220), .B(n287), .Z(product[10]) );
  NAND2_X1 U262 ( .A1(n253), .A2(n27), .ZN(n288) );
  NAND2_X1 U263 ( .A1(n277), .A2(n24), .ZN(n289) );
  NAND2_X1 U264 ( .A1(n27), .A2(n24), .ZN(n290) );
  NAND3_X1 U265 ( .A1(n288), .A2(n289), .A3(n290), .ZN(n5) );
  XOR2_X1 U266 ( .A(n95), .B(n102), .Z(n56) );
  BUF_X2 U267 ( .A(a[1]), .Z(n291) );
  XNOR2_X1 U268 ( .A(n215), .B(n292), .ZN(product[14]) );
  XNOR2_X1 U269 ( .A(n305), .B(n15), .ZN(n292) );
  XOR2_X2 U270 ( .A(a[2]), .B(n314), .Z(n293) );
  XOR2_X1 U271 ( .A(a[2]), .B(n314), .Z(n321) );
  AND3_X1 U272 ( .A1(n296), .A2(n295), .A3(n297), .ZN(product[15]) );
  INV_X1 U273 ( .A(n329), .ZN(n311) );
  OAI22_X1 U274 ( .A1(n350), .A2(n344), .B1(n342), .B2(n352), .ZN(n15) );
  INV_X1 U275 ( .A(n340), .ZN(n308) );
  INV_X1 U276 ( .A(n21), .ZN(n307) );
  INV_X1 U277 ( .A(n320), .ZN(n313) );
  INV_X1 U278 ( .A(n31), .ZN(n310) );
  INV_X1 U279 ( .A(b[0]), .ZN(n303) );
  INV_X1 U280 ( .A(a[0]), .ZN(n315) );
  INV_X1 U281 ( .A(a[3]), .ZN(n312) );
  INV_X1 U282 ( .A(a[5]), .ZN(n309) );
  INV_X1 U283 ( .A(a[7]), .ZN(n306) );
  NAND2_X1 U284 ( .A1(n254), .A2(n305), .ZN(n295) );
  NAND2_X1 U285 ( .A1(n255), .A2(n15), .ZN(n296) );
  NAND2_X1 U286 ( .A1(n305), .A2(n15), .ZN(n297) );
  XOR2_X1 U287 ( .A(n19), .B(n18), .Z(n298) );
  XOR2_X1 U288 ( .A(n239), .B(n298), .Z(product[12]) );
  NAND2_X1 U289 ( .A1(n228), .A2(n19), .ZN(n299) );
  NAND2_X1 U290 ( .A1(n4), .A2(n18), .ZN(n300) );
  NAND2_X1 U291 ( .A1(n19), .A2(n18), .ZN(n301) );
  NAND3_X1 U292 ( .A1(n299), .A2(n300), .A3(n301), .ZN(n3) );
  INV_X1 U293 ( .A(n351), .ZN(n305) );
  INV_X1 U294 ( .A(a[1]), .ZN(n314) );
  NAND2_X2 U295 ( .A1(n321), .A2(n359), .ZN(n323) );
  XOR2_X2 U296 ( .A(a[6]), .B(n309), .Z(n342) );
  NOR2_X1 U297 ( .A1(n315), .A2(n286), .ZN(product[0]) );
  OAI22_X1 U298 ( .A1(n316), .A2(n317), .B1(n318), .B2(n315), .ZN(n99) );
  OAI22_X1 U299 ( .A1(n318), .A2(n317), .B1(n319), .B2(n315), .ZN(n98) );
  XNOR2_X1 U300 ( .A(b[6]), .B(n291), .ZN(n318) );
  OAI22_X1 U301 ( .A1(n315), .A2(n319), .B1(n317), .B2(n319), .ZN(n320) );
  XNOR2_X1 U302 ( .A(b[7]), .B(n291), .ZN(n319) );
  NOR2_X1 U303 ( .A1(n293), .A2(n286), .ZN(n96) );
  OAI22_X1 U304 ( .A1(n322), .A2(n323), .B1(n293), .B2(n324), .ZN(n95) );
  XNOR2_X1 U305 ( .A(a[3]), .B(n302), .ZN(n322) );
  OAI22_X1 U306 ( .A1(n324), .A2(n323), .B1(n293), .B2(n325), .ZN(n94) );
  XNOR2_X1 U307 ( .A(n212), .B(a[3]), .ZN(n324) );
  OAI22_X1 U308 ( .A1(n325), .A2(n323), .B1(n293), .B2(n326), .ZN(n93) );
  XNOR2_X1 U309 ( .A(b[2]), .B(a[3]), .ZN(n325) );
  OAI22_X1 U310 ( .A1(n326), .A2(n323), .B1(n293), .B2(n327), .ZN(n92) );
  XNOR2_X1 U311 ( .A(b[3]), .B(a[3]), .ZN(n326) );
  OAI22_X1 U312 ( .A1(n327), .A2(n323), .B1(n293), .B2(n328), .ZN(n91) );
  XNOR2_X1 U313 ( .A(b[4]), .B(a[3]), .ZN(n327) );
  OAI22_X1 U314 ( .A1(n330), .A2(n293), .B1(n323), .B2(n330), .ZN(n329) );
  NOR2_X1 U315 ( .A1(n331), .A2(n286), .ZN(n88) );
  OAI22_X1 U316 ( .A1(n332), .A2(n333), .B1(n331), .B2(n334), .ZN(n87) );
  XNOR2_X1 U317 ( .A(a[5]), .B(n302), .ZN(n332) );
  OAI22_X1 U318 ( .A1(n334), .A2(n333), .B1(n331), .B2(n335), .ZN(n86) );
  XNOR2_X1 U319 ( .A(n213), .B(a[5]), .ZN(n334) );
  OAI22_X1 U320 ( .A1(n335), .A2(n333), .B1(n331), .B2(n336), .ZN(n85) );
  XNOR2_X1 U321 ( .A(b[2]), .B(a[5]), .ZN(n335) );
  OAI22_X1 U322 ( .A1(n336), .A2(n333), .B1(n331), .B2(n337), .ZN(n84) );
  XNOR2_X1 U323 ( .A(b[3]), .B(a[5]), .ZN(n336) );
  OAI22_X1 U324 ( .A1(n337), .A2(n333), .B1(n331), .B2(n338), .ZN(n83) );
  XNOR2_X1 U325 ( .A(b[4]), .B(a[5]), .ZN(n337) );
  OAI22_X1 U326 ( .A1(n338), .A2(n333), .B1(n331), .B2(n339), .ZN(n82) );
  XNOR2_X1 U327 ( .A(b[5]), .B(a[5]), .ZN(n338) );
  OAI22_X1 U328 ( .A1(n341), .A2(n331), .B1(n333), .B2(n341), .ZN(n340) );
  NOR2_X1 U329 ( .A1(n342), .A2(n286), .ZN(n80) );
  OAI22_X1 U330 ( .A1(n343), .A2(n344), .B1(n342), .B2(n345), .ZN(n79) );
  XNOR2_X1 U331 ( .A(a[7]), .B(n302), .ZN(n343) );
  OAI22_X1 U332 ( .A1(n346), .A2(n344), .B1(n342), .B2(n347), .ZN(n77) );
  OAI22_X1 U333 ( .A1(n347), .A2(n344), .B1(n342), .B2(n348), .ZN(n76) );
  XNOR2_X1 U334 ( .A(b[3]), .B(a[7]), .ZN(n347) );
  OAI22_X1 U335 ( .A1(n348), .A2(n344), .B1(n342), .B2(n349), .ZN(n75) );
  XNOR2_X1 U336 ( .A(b[4]), .B(a[7]), .ZN(n348) );
  OAI22_X1 U337 ( .A1(n349), .A2(n344), .B1(n342), .B2(n350), .ZN(n74) );
  XNOR2_X1 U338 ( .A(b[5]), .B(a[7]), .ZN(n349) );
  OAI22_X1 U339 ( .A1(n352), .A2(n342), .B1(n344), .B2(n352), .ZN(n351) );
  OAI21_X1 U340 ( .B1(n302), .B2(n314), .A(n317), .ZN(n72) );
  OAI21_X1 U341 ( .B1(n312), .B2(n323), .A(n353), .ZN(n71) );
  OR3_X1 U342 ( .A1(n293), .A2(n302), .A3(n312), .ZN(n353) );
  OAI21_X1 U343 ( .B1(n309), .B2(n333), .A(n354), .ZN(n70) );
  OR3_X1 U344 ( .A1(n331), .A2(n302), .A3(n309), .ZN(n354) );
  OAI21_X1 U345 ( .B1(n306), .B2(n344), .A(n355), .ZN(n69) );
  OR3_X1 U346 ( .A1(n342), .A2(n302), .A3(n306), .ZN(n355) );
  XNOR2_X1 U347 ( .A(n356), .B(n357), .ZN(n38) );
  OR2_X1 U348 ( .A1(n356), .A2(n357), .ZN(n37) );
  OAI22_X1 U349 ( .A1(n328), .A2(n323), .B1(n293), .B2(n358), .ZN(n357) );
  XNOR2_X1 U350 ( .A(b[5]), .B(a[3]), .ZN(n328) );
  OAI22_X1 U351 ( .A1(n345), .A2(n344), .B1(n342), .B2(n346), .ZN(n356) );
  XNOR2_X1 U352 ( .A(b[2]), .B(a[7]), .ZN(n346) );
  XNOR2_X1 U353 ( .A(n213), .B(a[7]), .ZN(n345) );
  OAI22_X1 U354 ( .A1(n358), .A2(n323), .B1(n293), .B2(n330), .ZN(n31) );
  XNOR2_X1 U355 ( .A(b[7]), .B(a[3]), .ZN(n330) );
  XNOR2_X1 U356 ( .A(n312), .B(a[2]), .ZN(n359) );
  XNOR2_X1 U357 ( .A(b[6]), .B(a[3]), .ZN(n358) );
  OAI22_X1 U358 ( .A1(n339), .A2(n333), .B1(n331), .B2(n341), .ZN(n21) );
  XNOR2_X1 U359 ( .A(b[7]), .B(a[5]), .ZN(n341) );
  XNOR2_X1 U360 ( .A(n309), .B(a[4]), .ZN(n360) );
  XNOR2_X1 U361 ( .A(b[6]), .B(a[5]), .ZN(n339) );
  XNOR2_X1 U362 ( .A(b[7]), .B(a[7]), .ZN(n352) );
  NAND2_X1 U363 ( .A1(n342), .A2(n361), .ZN(n344) );
  XNOR2_X1 U364 ( .A(n306), .B(a[6]), .ZN(n361) );
  XNOR2_X1 U365 ( .A(b[6]), .B(a[7]), .ZN(n350) );
  OAI22_X1 U366 ( .A1(n302), .A2(n317), .B1(n362), .B2(n315), .ZN(n104) );
  OAI22_X1 U367 ( .A1(n252), .A2(n317), .B1(n363), .B2(n315), .ZN(n103) );
  XNOR2_X1 U368 ( .A(b[1]), .B(n291), .ZN(n362) );
  OAI22_X1 U369 ( .A1(n363), .A2(n317), .B1(n364), .B2(n315), .ZN(n102) );
  XNOR2_X1 U370 ( .A(b[2]), .B(n291), .ZN(n363) );
  OAI22_X1 U371 ( .A1(n364), .A2(n317), .B1(n365), .B2(n315), .ZN(n101) );
  XNOR2_X1 U372 ( .A(b[3]), .B(n291), .ZN(n364) );
  OAI22_X1 U373 ( .A1(n365), .A2(n317), .B1(n316), .B2(n315), .ZN(n100) );
  XNOR2_X1 U374 ( .A(b[5]), .B(n291), .ZN(n316) );
  NAND2_X1 U375 ( .A1(n291), .A2(n315), .ZN(n317) );
  XNOR2_X1 U376 ( .A(b[4]), .B(n291), .ZN(n365) );
endmodule


module mac_13 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_13_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_13_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_12_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  wire   [15:1] carry;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CLKBUF_X1 U1 ( .A(carry[10]), .Z(n1) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n64) );
  XNOR2_X1 U3 ( .A(B[15]), .B(A[15]), .ZN(n2) );
  CLKBUF_X1 U4 ( .A(carry[11]), .Z(n3) );
  XOR2_X1 U5 ( .A(B[10]), .B(A[10]), .Z(n4) );
  XOR2_X1 U6 ( .A(n1), .B(n4), .Z(SUM[10]) );
  NAND2_X1 U7 ( .A1(carry[10]), .A2(B[10]), .ZN(n5) );
  NAND2_X1 U8 ( .A1(carry[10]), .A2(A[10]), .ZN(n6) );
  NAND2_X1 U9 ( .A1(B[10]), .A2(A[10]), .ZN(n7) );
  NAND3_X1 U10 ( .A1(n5), .A2(n6), .A3(n7), .ZN(carry[11]) );
  NAND3_X1 U11 ( .A1(n15), .A2(n16), .A3(n17), .ZN(n8) );
  NAND3_X1 U12 ( .A1(n11), .A2(n12), .A3(n13), .ZN(n9) );
  XOR2_X1 U13 ( .A(B[11]), .B(A[11]), .Z(n10) );
  XOR2_X1 U14 ( .A(n3), .B(n10), .Z(SUM[11]) );
  NAND2_X1 U15 ( .A1(carry[11]), .A2(B[11]), .ZN(n11) );
  NAND2_X1 U16 ( .A1(carry[11]), .A2(A[11]), .ZN(n12) );
  NAND2_X1 U17 ( .A1(B[11]), .A2(A[11]), .ZN(n13) );
  NAND3_X1 U18 ( .A1(n11), .A2(n12), .A3(n13), .ZN(carry[12]) );
  XOR2_X1 U19 ( .A(B[5]), .B(A[5]), .Z(n14) );
  XOR2_X1 U20 ( .A(carry[5]), .B(n14), .Z(SUM[5]) );
  NAND2_X1 U21 ( .A1(carry[5]), .A2(B[5]), .ZN(n15) );
  NAND2_X1 U22 ( .A1(carry[5]), .A2(A[5]), .ZN(n16) );
  NAND2_X1 U23 ( .A1(B[5]), .A2(A[5]), .ZN(n17) );
  NAND3_X1 U24 ( .A1(n15), .A2(n16), .A3(n17), .ZN(carry[6]) );
  NAND3_X1 U25 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n18) );
  NAND3_X1 U26 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n19) );
  NAND3_X1 U27 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n20) );
  XOR2_X1 U28 ( .A(B[12]), .B(A[12]), .Z(n21) );
  XOR2_X1 U29 ( .A(n9), .B(n21), .Z(SUM[12]) );
  NAND2_X1 U30 ( .A1(n9), .A2(B[12]), .ZN(n22) );
  NAND2_X1 U31 ( .A1(carry[12]), .A2(A[12]), .ZN(n23) );
  NAND2_X1 U32 ( .A1(B[12]), .A2(A[12]), .ZN(n24) );
  NAND3_X1 U33 ( .A1(n22), .A2(n23), .A3(n24), .ZN(carry[13]) );
  XOR2_X1 U34 ( .A(B[6]), .B(A[6]), .Z(n25) );
  XOR2_X1 U35 ( .A(n8), .B(n25), .Z(SUM[6]) );
  NAND2_X1 U36 ( .A1(n8), .A2(B[6]), .ZN(n26) );
  NAND2_X1 U37 ( .A1(carry[6]), .A2(A[6]), .ZN(n27) );
  NAND2_X1 U38 ( .A1(B[6]), .A2(A[6]), .ZN(n28) );
  NAND3_X1 U39 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[7]) );
  XNOR2_X1 U40 ( .A(carry[15]), .B(n2), .ZN(SUM[15]) );
  NAND3_X1 U41 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n29) );
  NAND3_X1 U42 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n30) );
  NAND3_X1 U43 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n31) );
  NAND3_X1 U44 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n32) );
  XOR2_X1 U45 ( .A(B[13]), .B(A[13]), .Z(n33) );
  XOR2_X1 U46 ( .A(n18), .B(n33), .Z(SUM[13]) );
  NAND2_X1 U47 ( .A1(n18), .A2(B[13]), .ZN(n34) );
  NAND2_X1 U48 ( .A1(carry[13]), .A2(A[13]), .ZN(n35) );
  NAND2_X1 U49 ( .A1(B[13]), .A2(A[13]), .ZN(n36) );
  XOR2_X1 U50 ( .A(B[7]), .B(A[7]), .Z(n37) );
  XOR2_X1 U51 ( .A(carry[7]), .B(n37), .Z(SUM[7]) );
  NAND2_X1 U52 ( .A1(n19), .A2(B[7]), .ZN(n38) );
  NAND2_X1 U53 ( .A1(carry[7]), .A2(A[7]), .ZN(n39) );
  NAND2_X1 U54 ( .A1(B[7]), .A2(A[7]), .ZN(n40) );
  NAND3_X1 U55 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[8]) );
  NAND3_X1 U56 ( .A1(n57), .A2(n58), .A3(n59), .ZN(n41) );
  NAND3_X1 U57 ( .A1(n57), .A2(n58), .A3(n59), .ZN(n42) );
  XOR2_X1 U58 ( .A(B[14]), .B(A[14]), .Z(n43) );
  XOR2_X1 U59 ( .A(n30), .B(n43), .Z(SUM[14]) );
  NAND2_X1 U60 ( .A1(n29), .A2(B[14]), .ZN(n44) );
  NAND2_X1 U61 ( .A1(n29), .A2(A[14]), .ZN(n45) );
  NAND2_X1 U62 ( .A1(B[14]), .A2(A[14]), .ZN(n46) );
  NAND3_X1 U63 ( .A1(n44), .A2(n45), .A3(n46), .ZN(carry[15]) );
  CLKBUF_X1 U64 ( .A(n20), .Z(n47) );
  XOR2_X1 U65 ( .A(B[8]), .B(A[8]), .Z(n48) );
  XOR2_X1 U66 ( .A(n32), .B(n48), .Z(SUM[8]) );
  NAND2_X1 U67 ( .A1(n31), .A2(B[8]), .ZN(n49) );
  NAND2_X1 U68 ( .A1(carry[8]), .A2(A[8]), .ZN(n50) );
  NAND2_X1 U69 ( .A1(B[8]), .A2(A[8]), .ZN(n51) );
  NAND3_X1 U70 ( .A1(n49), .A2(n50), .A3(n51), .ZN(carry[9]) );
  XOR2_X1 U71 ( .A(B[9]), .B(A[9]), .Z(n52) );
  XOR2_X1 U72 ( .A(n47), .B(n52), .Z(SUM[9]) );
  NAND2_X1 U73 ( .A1(n20), .A2(B[9]), .ZN(n53) );
  NAND2_X1 U74 ( .A1(carry[9]), .A2(A[9]), .ZN(n54) );
  NAND2_X1 U75 ( .A1(B[9]), .A2(A[9]), .ZN(n55) );
  NAND3_X1 U76 ( .A1(n53), .A2(n54), .A3(n55), .ZN(carry[10]) );
  XOR2_X1 U77 ( .A(B[1]), .B(A[1]), .Z(n56) );
  XOR2_X1 U78 ( .A(n64), .B(n56), .Z(SUM[1]) );
  NAND2_X1 U79 ( .A1(n64), .A2(B[1]), .ZN(n57) );
  NAND2_X1 U80 ( .A1(n64), .A2(A[1]), .ZN(n58) );
  NAND2_X1 U81 ( .A1(B[1]), .A2(A[1]), .ZN(n59) );
  NAND3_X1 U82 ( .A1(n57), .A2(n58), .A3(n59), .ZN(carry[2]) );
  XOR2_X1 U83 ( .A(B[2]), .B(A[2]), .Z(n60) );
  XOR2_X1 U84 ( .A(n42), .B(n60), .Z(SUM[2]) );
  NAND2_X1 U85 ( .A1(n41), .A2(B[2]), .ZN(n61) );
  NAND2_X1 U86 ( .A1(carry[2]), .A2(A[2]), .ZN(n62) );
  NAND2_X1 U87 ( .A1(B[2]), .A2(A[2]), .ZN(n63) );
  NAND3_X1 U88 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[3]) );
  XOR2_X1 U89 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_12_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74,
         n75, n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92,
         n93, n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n303), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n302), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n306), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n305), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n308), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  CLKBUF_X1 U157 ( .A(n50), .Z(n206) );
  CLKBUF_X1 U158 ( .A(n244), .Z(n207) );
  INV_X1 U159 ( .A(n297), .ZN(n208) );
  CLKBUF_X1 U160 ( .A(n294), .Z(n209) );
  CLKBUF_X1 U161 ( .A(b[1]), .Z(n210) );
  CLKBUF_X1 U162 ( .A(a[3]), .Z(n211) );
  INV_X1 U163 ( .A(n309), .ZN(n212) );
  NAND2_X2 U164 ( .A1(n226), .A2(n227), .ZN(n213) );
  NAND2_X1 U165 ( .A1(n226), .A2(n227), .ZN(n326) );
  NAND2_X1 U166 ( .A1(n241), .A2(n18), .ZN(n214) );
  CLKBUF_X1 U167 ( .A(n9), .Z(n215) );
  CLKBUF_X1 U168 ( .A(n259), .Z(n216) );
  NAND3_X1 U169 ( .A1(n207), .A2(n245), .A3(n246), .ZN(n217) );
  CLKBUF_X1 U170 ( .A(n269), .Z(n218) );
  AND2_X1 U171 ( .A1(n104), .A2(n72), .ZN(n219) );
  NAND3_X1 U172 ( .A1(n230), .A2(n229), .A3(n231), .ZN(n220) );
  NAND3_X1 U173 ( .A1(n267), .A2(n266), .A3(n268), .ZN(n221) );
  CLKBUF_X1 U174 ( .A(n220), .Z(n222) );
  NAND3_X1 U175 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n223) );
  NAND3_X1 U176 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n224) );
  NAND2_X1 U177 ( .A1(a[4]), .A2(a[3]), .ZN(n226) );
  NAND2_X1 U178 ( .A1(n225), .A2(n307), .ZN(n227) );
  INV_X1 U179 ( .A(a[4]), .ZN(n225) );
  XOR2_X1 U180 ( .A(n27), .B(n24), .Z(n228) );
  XOR2_X1 U181 ( .A(n224), .B(n228), .Z(product[10]) );
  NAND2_X1 U182 ( .A1(n6), .A2(n27), .ZN(n229) );
  NAND2_X1 U183 ( .A1(n223), .A2(n24), .ZN(n230) );
  NAND2_X1 U184 ( .A1(n27), .A2(n24), .ZN(n231) );
  NAND3_X1 U185 ( .A1(n230), .A2(n229), .A3(n231), .ZN(n5) );
  NAND3_X1 U186 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n232) );
  NAND3_X1 U187 ( .A1(n209), .A2(n295), .A3(n296), .ZN(n233) );
  NAND3_X1 U188 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n234) );
  CLKBUF_X1 U189 ( .A(n56), .Z(n235) );
  BUF_X2 U190 ( .A(n316), .Z(n236) );
  XNOR2_X1 U191 ( .A(a[2]), .B(a[1]), .ZN(n316) );
  XOR2_X1 U192 ( .A(n46), .B(n49), .Z(n237) );
  XOR2_X1 U193 ( .A(n233), .B(n237), .Z(product[6]) );
  NAND2_X1 U194 ( .A1(n232), .A2(n46), .ZN(n238) );
  NAND2_X1 U195 ( .A1(n10), .A2(n49), .ZN(n239) );
  NAND2_X1 U196 ( .A1(n46), .A2(n49), .ZN(n240) );
  NAND3_X1 U197 ( .A1(n239), .A2(n238), .A3(n240), .ZN(n9) );
  NAND3_X1 U198 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n241) );
  NAND3_X1 U199 ( .A1(n285), .A2(n214), .A3(n287), .ZN(n242) );
  XOR2_X1 U200 ( .A(n23), .B(n20), .Z(n243) );
  XOR2_X1 U201 ( .A(n222), .B(n243), .Z(product[11]) );
  NAND2_X1 U202 ( .A1(n220), .A2(n23), .ZN(n244) );
  NAND2_X1 U203 ( .A1(n5), .A2(n20), .ZN(n245) );
  NAND2_X1 U204 ( .A1(n23), .A2(n20), .ZN(n246) );
  NAND3_X1 U205 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n4) );
  AND3_X1 U206 ( .A1(n258), .A2(n257), .A3(n256), .ZN(product[15]) );
  NAND3_X1 U207 ( .A1(n285), .A2(n286), .A3(n287), .ZN(n248) );
  NAND3_X1 U208 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n249) );
  XNOR2_X1 U209 ( .A(b[1]), .B(a[1]), .ZN(n250) );
  XOR2_X1 U210 ( .A(n17), .B(n299), .Z(n251) );
  XOR2_X1 U211 ( .A(n251), .B(n242), .Z(product[13]) );
  NAND2_X1 U212 ( .A1(n17), .A2(n299), .ZN(n252) );
  NAND2_X1 U213 ( .A1(n17), .A2(n248), .ZN(n253) );
  NAND2_X1 U214 ( .A1(n299), .A2(n3), .ZN(n254) );
  NAND3_X1 U215 ( .A1(n254), .A2(n253), .A3(n252), .ZN(n2) );
  XOR2_X1 U216 ( .A(n300), .B(n15), .Z(n255) );
  XOR2_X1 U217 ( .A(n255), .B(n249), .Z(product[14]) );
  NAND2_X1 U218 ( .A1(n300), .A2(n15), .ZN(n256) );
  NAND2_X1 U219 ( .A1(n300), .A2(n2), .ZN(n257) );
  NAND2_X1 U220 ( .A1(n15), .A2(n2), .ZN(n258) );
  NAND3_X1 U221 ( .A1(n263), .A2(n262), .A3(n264), .ZN(n259) );
  INV_X1 U222 ( .A(n298), .ZN(n260) );
  INV_X1 U223 ( .A(n298), .ZN(n297) );
  XOR2_X1 U224 ( .A(n40), .B(n45), .Z(n261) );
  XOR2_X1 U225 ( .A(n215), .B(n261), .Z(product[7]) );
  NAND2_X1 U226 ( .A1(n234), .A2(n40), .ZN(n262) );
  NAND2_X1 U227 ( .A1(n9), .A2(n45), .ZN(n263) );
  NAND2_X1 U228 ( .A1(n40), .A2(n45), .ZN(n264) );
  NAND3_X1 U229 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n8) );
  XOR2_X1 U230 ( .A(n103), .B(n96), .Z(n265) );
  XOR2_X1 U231 ( .A(n219), .B(n265), .Z(product[2]) );
  NAND2_X1 U232 ( .A1(n219), .A2(n103), .ZN(n266) );
  NAND2_X1 U233 ( .A1(n14), .A2(n96), .ZN(n267) );
  NAND2_X1 U234 ( .A1(n103), .A2(n96), .ZN(n268) );
  NAND3_X1 U235 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n13) );
  NAND3_X1 U236 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n269) );
  XOR2_X1 U237 ( .A(n34), .B(n39), .Z(n270) );
  XOR2_X1 U238 ( .A(n216), .B(n270), .Z(product[8]) );
  NAND2_X1 U239 ( .A1(n259), .A2(n34), .ZN(n271) );
  NAND2_X1 U240 ( .A1(n8), .A2(n39), .ZN(n272) );
  NAND2_X1 U241 ( .A1(n34), .A2(n39), .ZN(n273) );
  NAND3_X1 U242 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n7) );
  NAND3_X1 U243 ( .A1(n281), .A2(n282), .A3(n283), .ZN(n274) );
  XOR2_X1 U244 ( .A(n33), .B(n28), .Z(n275) );
  XOR2_X1 U245 ( .A(n218), .B(n275), .Z(product[9]) );
  NAND2_X1 U246 ( .A1(n269), .A2(n33), .ZN(n276) );
  NAND2_X1 U247 ( .A1(n7), .A2(n28), .ZN(n277) );
  NAND2_X1 U248 ( .A1(n33), .A2(n28), .ZN(n278) );
  NAND3_X1 U249 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n6) );
  NAND3_X1 U250 ( .A1(n290), .A2(n291), .A3(n292), .ZN(n279) );
  XOR2_X1 U251 ( .A(n235), .B(n71), .Z(n280) );
  XOR2_X1 U252 ( .A(n221), .B(n280), .Z(product[3]) );
  NAND2_X1 U253 ( .A1(n221), .A2(n56), .ZN(n281) );
  NAND2_X1 U254 ( .A1(n13), .A2(n71), .ZN(n282) );
  NAND2_X1 U255 ( .A1(n56), .A2(n71), .ZN(n283) );
  NAND3_X1 U256 ( .A1(n281), .A2(n282), .A3(n283), .ZN(n12) );
  XOR2_X1 U257 ( .A(n19), .B(n18), .Z(n284) );
  XOR2_X1 U258 ( .A(n217), .B(n284), .Z(product[12]) );
  NAND2_X1 U259 ( .A1(n4), .A2(n19), .ZN(n285) );
  NAND2_X1 U260 ( .A1(n241), .A2(n18), .ZN(n286) );
  NAND2_X1 U261 ( .A1(n19), .A2(n18), .ZN(n287) );
  NAND3_X1 U262 ( .A1(n214), .A2(n285), .A3(n287), .ZN(n3) );
  CLKBUF_X1 U263 ( .A(n279), .Z(n288) );
  INV_X1 U264 ( .A(n15), .ZN(n299) );
  INV_X1 U265 ( .A(n21), .ZN(n302) );
  INV_X1 U266 ( .A(n335), .ZN(n303) );
  INV_X1 U267 ( .A(n315), .ZN(n308) );
  INV_X1 U268 ( .A(n324), .ZN(n306) );
  INV_X1 U269 ( .A(b[0]), .ZN(n298) );
  INV_X1 U270 ( .A(n346), .ZN(n300) );
  INV_X1 U271 ( .A(n31), .ZN(n305) );
  INV_X1 U272 ( .A(a[0]), .ZN(n310) );
  INV_X1 U273 ( .A(a[5]), .ZN(n304) );
  INV_X1 U274 ( .A(a[7]), .ZN(n301) );
  XOR2_X1 U275 ( .A(n54), .B(n55), .Z(n289) );
  XOR2_X1 U276 ( .A(n274), .B(n289), .Z(product[4]) );
  NAND2_X1 U277 ( .A1(n274), .A2(n54), .ZN(n290) );
  NAND2_X1 U278 ( .A1(n12), .A2(n55), .ZN(n291) );
  NAND2_X1 U279 ( .A1(n54), .A2(n55), .ZN(n292) );
  NAND3_X1 U280 ( .A1(n290), .A2(n291), .A3(n292), .ZN(n11) );
  XOR2_X1 U281 ( .A(n206), .B(n53), .Z(n293) );
  XOR2_X1 U282 ( .A(n288), .B(n293), .Z(product[5]) );
  NAND2_X1 U283 ( .A1(n279), .A2(n50), .ZN(n294) );
  NAND2_X1 U284 ( .A1(n11), .A2(n53), .ZN(n295) );
  NAND2_X1 U285 ( .A1(n50), .A2(n53), .ZN(n296) );
  NAND3_X1 U286 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n10) );
  NAND2_X2 U287 ( .A1(n326), .A2(n355), .ZN(n328) );
  INV_X1 U288 ( .A(a[3]), .ZN(n307) );
  INV_X1 U289 ( .A(a[1]), .ZN(n309) );
  NAND2_X2 U290 ( .A1(n316), .A2(n354), .ZN(n318) );
  XOR2_X2 U291 ( .A(a[6]), .B(n304), .Z(n337) );
  NOR2_X1 U292 ( .A1(n310), .A2(n208), .ZN(product[0]) );
  OAI22_X1 U293 ( .A1(n311), .A2(n312), .B1(n313), .B2(n310), .ZN(n99) );
  OAI22_X1 U294 ( .A1(n313), .A2(n312), .B1(n314), .B2(n310), .ZN(n98) );
  XNOR2_X1 U295 ( .A(b[6]), .B(n212), .ZN(n313) );
  OAI22_X1 U296 ( .A1(n310), .A2(n314), .B1(n312), .B2(n314), .ZN(n315) );
  XNOR2_X1 U297 ( .A(b[7]), .B(n212), .ZN(n314) );
  NOR2_X1 U298 ( .A1(n236), .A2(n298), .ZN(n96) );
  OAI22_X1 U299 ( .A1(n317), .A2(n318), .B1(n236), .B2(n319), .ZN(n95) );
  XNOR2_X1 U300 ( .A(a[3]), .B(n297), .ZN(n317) );
  OAI22_X1 U301 ( .A1(n319), .A2(n318), .B1(n236), .B2(n320), .ZN(n94) );
  XNOR2_X1 U302 ( .A(b[1]), .B(a[3]), .ZN(n319) );
  OAI22_X1 U303 ( .A1(n320), .A2(n318), .B1(n236), .B2(n321), .ZN(n93) );
  XNOR2_X1 U304 ( .A(b[2]), .B(a[3]), .ZN(n320) );
  OAI22_X1 U305 ( .A1(n321), .A2(n318), .B1(n236), .B2(n322), .ZN(n92) );
  XNOR2_X1 U306 ( .A(b[3]), .B(n211), .ZN(n321) );
  OAI22_X1 U307 ( .A1(n322), .A2(n318), .B1(n236), .B2(n323), .ZN(n91) );
  XNOR2_X1 U308 ( .A(b[4]), .B(a[3]), .ZN(n322) );
  OAI22_X1 U309 ( .A1(n325), .A2(n236), .B1(n318), .B2(n325), .ZN(n324) );
  NOR2_X1 U310 ( .A1(n213), .A2(n208), .ZN(n88) );
  OAI22_X1 U311 ( .A1(n327), .A2(n328), .B1(n213), .B2(n329), .ZN(n87) );
  XNOR2_X1 U312 ( .A(a[5]), .B(n260), .ZN(n327) );
  OAI22_X1 U313 ( .A1(n329), .A2(n328), .B1(n213), .B2(n330), .ZN(n86) );
  XNOR2_X1 U314 ( .A(b[1]), .B(a[5]), .ZN(n329) );
  OAI22_X1 U315 ( .A1(n330), .A2(n328), .B1(n213), .B2(n331), .ZN(n85) );
  XNOR2_X1 U316 ( .A(b[2]), .B(a[5]), .ZN(n330) );
  OAI22_X1 U317 ( .A1(n331), .A2(n328), .B1(n213), .B2(n332), .ZN(n84) );
  XNOR2_X1 U318 ( .A(b[3]), .B(a[5]), .ZN(n331) );
  OAI22_X1 U319 ( .A1(n332), .A2(n328), .B1(n213), .B2(n333), .ZN(n83) );
  XNOR2_X1 U320 ( .A(b[4]), .B(a[5]), .ZN(n332) );
  OAI22_X1 U321 ( .A1(n333), .A2(n328), .B1(n213), .B2(n334), .ZN(n82) );
  XNOR2_X1 U322 ( .A(b[5]), .B(a[5]), .ZN(n333) );
  OAI22_X1 U323 ( .A1(n336), .A2(n213), .B1(n328), .B2(n336), .ZN(n335) );
  NOR2_X1 U324 ( .A1(n337), .A2(n208), .ZN(n80) );
  OAI22_X1 U325 ( .A1(n338), .A2(n339), .B1(n337), .B2(n340), .ZN(n79) );
  XNOR2_X1 U326 ( .A(a[7]), .B(n260), .ZN(n338) );
  OAI22_X1 U327 ( .A1(n341), .A2(n339), .B1(n337), .B2(n342), .ZN(n77) );
  OAI22_X1 U328 ( .A1(n342), .A2(n339), .B1(n337), .B2(n343), .ZN(n76) );
  XNOR2_X1 U329 ( .A(b[3]), .B(a[7]), .ZN(n342) );
  OAI22_X1 U330 ( .A1(n343), .A2(n339), .B1(n337), .B2(n344), .ZN(n75) );
  XNOR2_X1 U331 ( .A(b[4]), .B(a[7]), .ZN(n343) );
  OAI22_X1 U332 ( .A1(n344), .A2(n339), .B1(n337), .B2(n345), .ZN(n74) );
  XNOR2_X1 U333 ( .A(b[5]), .B(a[7]), .ZN(n344) );
  OAI22_X1 U334 ( .A1(n347), .A2(n337), .B1(n339), .B2(n347), .ZN(n346) );
  OAI21_X1 U335 ( .B1(n297), .B2(n309), .A(n312), .ZN(n72) );
  OAI21_X1 U336 ( .B1(n307), .B2(n318), .A(n348), .ZN(n71) );
  OR3_X1 U337 ( .A1(n236), .A2(n260), .A3(n307), .ZN(n348) );
  OAI21_X1 U338 ( .B1(n304), .B2(n328), .A(n349), .ZN(n70) );
  OR3_X1 U339 ( .A1(n326), .A2(n297), .A3(n304), .ZN(n349) );
  OAI21_X1 U340 ( .B1(n301), .B2(n339), .A(n350), .ZN(n69) );
  OR3_X1 U341 ( .A1(n337), .A2(n260), .A3(n301), .ZN(n350) );
  XNOR2_X1 U342 ( .A(n351), .B(n352), .ZN(n38) );
  OR2_X1 U343 ( .A1(n351), .A2(n352), .ZN(n37) );
  OAI22_X1 U344 ( .A1(n323), .A2(n318), .B1(n236), .B2(n353), .ZN(n352) );
  XNOR2_X1 U345 ( .A(b[5]), .B(n211), .ZN(n323) );
  OAI22_X1 U346 ( .A1(n340), .A2(n339), .B1(n337), .B2(n341), .ZN(n351) );
  XNOR2_X1 U347 ( .A(b[2]), .B(a[7]), .ZN(n341) );
  XNOR2_X1 U348 ( .A(n210), .B(a[7]), .ZN(n340) );
  OAI22_X1 U349 ( .A1(n353), .A2(n318), .B1(n236), .B2(n325), .ZN(n31) );
  XNOR2_X1 U350 ( .A(b[7]), .B(n211), .ZN(n325) );
  XNOR2_X1 U351 ( .A(n307), .B(a[2]), .ZN(n354) );
  XNOR2_X1 U352 ( .A(b[6]), .B(n211), .ZN(n353) );
  OAI22_X1 U353 ( .A1(n334), .A2(n328), .B1(n213), .B2(n336), .ZN(n21) );
  XNOR2_X1 U354 ( .A(b[7]), .B(a[5]), .ZN(n336) );
  XNOR2_X1 U355 ( .A(n304), .B(a[4]), .ZN(n355) );
  XNOR2_X1 U356 ( .A(b[6]), .B(a[5]), .ZN(n334) );
  OAI22_X1 U357 ( .A1(n345), .A2(n339), .B1(n337), .B2(n347), .ZN(n15) );
  XNOR2_X1 U358 ( .A(b[7]), .B(a[7]), .ZN(n347) );
  NAND2_X1 U359 ( .A1(n337), .A2(n356), .ZN(n339) );
  XNOR2_X1 U360 ( .A(n301), .B(a[6]), .ZN(n356) );
  XNOR2_X1 U361 ( .A(b[6]), .B(a[7]), .ZN(n345) );
  OAI22_X1 U362 ( .A1(n260), .A2(n312), .B1(n357), .B2(n310), .ZN(n104) );
  OAI22_X1 U363 ( .A1(n250), .A2(n312), .B1(n358), .B2(n310), .ZN(n103) );
  XNOR2_X1 U364 ( .A(b[1]), .B(a[1]), .ZN(n357) );
  OAI22_X1 U365 ( .A1(n358), .A2(n312), .B1(n359), .B2(n310), .ZN(n102) );
  XNOR2_X1 U366 ( .A(b[2]), .B(a[1]), .ZN(n358) );
  OAI22_X1 U367 ( .A1(n359), .A2(n312), .B1(n360), .B2(n310), .ZN(n101) );
  XNOR2_X1 U368 ( .A(b[3]), .B(a[1]), .ZN(n359) );
  OAI22_X1 U369 ( .A1(n360), .A2(n312), .B1(n311), .B2(n310), .ZN(n100) );
  XNOR2_X1 U370 ( .A(b[5]), .B(n212), .ZN(n311) );
  NAND2_X1 U371 ( .A1(a[1]), .A2(n310), .ZN(n312) );
  XNOR2_X1 U372 ( .A(b[4]), .B(a[1]), .ZN(n360) );
endmodule


module mac_12 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  mac_12_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_12_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_11_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82;
  wire   [15:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .S(SUM[15]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  AND2_X2 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n82) );
  CLKBUF_X1 U2 ( .A(n54), .Z(n1) );
  CLKBUF_X1 U3 ( .A(n53), .Z(n2) );
  CLKBUF_X1 U4 ( .A(n16), .Z(n3) );
  NAND2_X1 U5 ( .A1(n32), .A2(B[8]), .ZN(n4) );
  CLKBUF_X1 U6 ( .A(n46), .Z(n5) );
  NAND3_X1 U7 ( .A1(n4), .A2(n60), .A3(n61), .ZN(n6) );
  CLKBUF_X1 U8 ( .A(n4), .Z(n7) );
  CLKBUF_X1 U9 ( .A(A[0]), .Z(n8) );
  CLKBUF_X1 U10 ( .A(carry[3]), .Z(n9) );
  NAND3_X1 U11 ( .A1(n15), .A2(n16), .A3(n17), .ZN(n10) );
  NAND3_X1 U12 ( .A1(n15), .A2(n3), .A3(n17), .ZN(n11) );
  NAND3_X1 U13 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n12) );
  NAND3_X1 U14 ( .A1(n27), .A2(n26), .A3(n28), .ZN(n13) );
  XOR2_X1 U15 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR2_X1 U16 ( .A(n9), .B(n14), .Z(SUM[3]) );
  NAND2_X1 U17 ( .A1(carry[3]), .A2(B[3]), .ZN(n15) );
  NAND2_X1 U18 ( .A1(carry[3]), .A2(A[3]), .ZN(n16) );
  NAND2_X1 U19 ( .A1(B[3]), .A2(A[3]), .ZN(n17) );
  NAND3_X1 U20 ( .A1(n15), .A2(n16), .A3(n17), .ZN(carry[4]) );
  NAND3_X1 U21 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n18) );
  NAND3_X1 U22 ( .A1(n2), .A2(n1), .A3(n55), .ZN(n19) );
  CLKBUF_X1 U23 ( .A(n45), .Z(n20) );
  CLKBUF_X1 U24 ( .A(n13), .Z(n21) );
  NAND3_X1 U25 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n22) );
  NAND3_X1 U26 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n23) );
  CLKBUF_X1 U27 ( .A(n67), .Z(n24) );
  XOR2_X1 U28 ( .A(B[10]), .B(A[10]), .Z(n25) );
  XOR2_X1 U29 ( .A(n19), .B(n25), .Z(SUM[10]) );
  NAND2_X1 U30 ( .A1(n18), .A2(B[10]), .ZN(n26) );
  NAND2_X1 U31 ( .A1(carry[10]), .A2(A[10]), .ZN(n27) );
  NAND2_X1 U32 ( .A1(B[10]), .A2(A[10]), .ZN(n28) );
  NAND3_X1 U33 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[11]) );
  CLKBUF_X1 U34 ( .A(n12), .Z(n29) );
  CLKBUF_X1 U35 ( .A(n23), .Z(n30) );
  NAND3_X1 U36 ( .A1(n24), .A2(n68), .A3(n69), .ZN(n31) );
  NAND3_X1 U37 ( .A1(n79), .A2(n80), .A3(n81), .ZN(n32) );
  XOR2_X1 U38 ( .A(B[4]), .B(A[4]), .Z(n33) );
  XOR2_X1 U39 ( .A(n11), .B(n33), .Z(SUM[4]) );
  NAND2_X1 U40 ( .A1(n10), .A2(B[4]), .ZN(n34) );
  NAND2_X1 U41 ( .A1(carry[4]), .A2(A[4]), .ZN(n35) );
  NAND2_X1 U42 ( .A1(B[4]), .A2(A[4]), .ZN(n36) );
  NAND3_X1 U43 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[5]) );
  XOR2_X1 U44 ( .A(B[11]), .B(A[11]), .Z(n37) );
  XOR2_X1 U45 ( .A(n21), .B(n37), .Z(SUM[11]) );
  NAND2_X1 U46 ( .A1(n13), .A2(B[11]), .ZN(n38) );
  NAND2_X1 U47 ( .A1(carry[11]), .A2(A[11]), .ZN(n39) );
  NAND2_X1 U48 ( .A1(B[11]), .A2(A[11]), .ZN(n40) );
  NAND3_X1 U49 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[12]) );
  XOR2_X1 U50 ( .A(B[5]), .B(A[5]), .Z(n41) );
  XOR2_X1 U51 ( .A(carry[5]), .B(n41), .Z(SUM[5]) );
  NAND2_X1 U52 ( .A1(n22), .A2(B[5]), .ZN(n42) );
  NAND2_X1 U53 ( .A1(n22), .A2(A[5]), .ZN(n43) );
  NAND2_X1 U54 ( .A1(B[5]), .A2(A[5]), .ZN(n44) );
  NAND3_X1 U55 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[6]) );
  NAND3_X1 U56 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n45) );
  NAND3_X1 U57 ( .A1(n71), .A2(n72), .A3(n73), .ZN(n46) );
  XOR2_X1 U58 ( .A(B[12]), .B(A[12]), .Z(n47) );
  XOR2_X1 U59 ( .A(n29), .B(n47), .Z(SUM[12]) );
  NAND2_X1 U60 ( .A1(n12), .A2(B[12]), .ZN(n48) );
  NAND2_X1 U61 ( .A1(carry[12]), .A2(A[12]), .ZN(n49) );
  NAND2_X1 U62 ( .A1(B[12]), .A2(A[12]), .ZN(n50) );
  NAND3_X1 U63 ( .A1(n48), .A2(n49), .A3(n50), .ZN(carry[13]) );
  NAND3_X1 U64 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n51) );
  XOR2_X1 U65 ( .A(B[9]), .B(A[9]), .Z(n52) );
  XOR2_X1 U66 ( .A(carry[9]), .B(n52), .Z(SUM[9]) );
  NAND2_X1 U67 ( .A1(n6), .A2(B[9]), .ZN(n53) );
  NAND2_X1 U68 ( .A1(n51), .A2(A[9]), .ZN(n54) );
  NAND2_X1 U69 ( .A1(B[9]), .A2(A[9]), .ZN(n55) );
  NAND3_X1 U70 ( .A1(n53), .A2(n54), .A3(n55), .ZN(carry[10]) );
  NAND3_X1 U71 ( .A1(n67), .A2(n68), .A3(n69), .ZN(n56) );
  CLKBUF_X1 U72 ( .A(n32), .Z(n57) );
  XOR2_X1 U73 ( .A(B[8]), .B(A[8]), .Z(n58) );
  XOR2_X1 U74 ( .A(n57), .B(n58), .Z(SUM[8]) );
  NAND2_X1 U75 ( .A1(n32), .A2(B[8]), .ZN(n59) );
  NAND2_X1 U76 ( .A1(carry[8]), .A2(A[8]), .ZN(n60) );
  NAND2_X1 U77 ( .A1(B[8]), .A2(A[8]), .ZN(n61) );
  NAND3_X1 U78 ( .A1(n7), .A2(n60), .A3(n61), .ZN(carry[9]) );
  XOR2_X1 U79 ( .A(B[1]), .B(A[1]), .Z(n62) );
  XOR2_X1 U80 ( .A(n82), .B(n62), .Z(SUM[1]) );
  NAND2_X1 U81 ( .A1(n82), .A2(B[1]), .ZN(n63) );
  NAND2_X1 U82 ( .A1(n82), .A2(A[1]), .ZN(n64) );
  NAND2_X1 U83 ( .A1(B[1]), .A2(A[1]), .ZN(n65) );
  NAND3_X1 U84 ( .A1(n63), .A2(n64), .A3(n65), .ZN(carry[2]) );
  XOR2_X1 U85 ( .A(B[13]), .B(A[13]), .Z(n66) );
  XOR2_X1 U86 ( .A(n20), .B(n66), .Z(SUM[13]) );
  NAND2_X1 U87 ( .A1(n45), .A2(B[13]), .ZN(n67) );
  NAND2_X1 U88 ( .A1(carry[13]), .A2(A[13]), .ZN(n68) );
  NAND2_X1 U89 ( .A1(B[13]), .A2(A[13]), .ZN(n69) );
  NAND3_X1 U90 ( .A1(n67), .A2(n68), .A3(n69), .ZN(carry[14]) );
  XOR2_X1 U91 ( .A(B[6]), .B(A[6]), .Z(n70) );
  XOR2_X1 U92 ( .A(n30), .B(n70), .Z(SUM[6]) );
  NAND2_X1 U93 ( .A1(n23), .A2(B[6]), .ZN(n71) );
  NAND2_X1 U94 ( .A1(carry[6]), .A2(A[6]), .ZN(n72) );
  NAND2_X1 U95 ( .A1(B[6]), .A2(A[6]), .ZN(n73) );
  NAND3_X1 U96 ( .A1(n71), .A2(n72), .A3(n73), .ZN(carry[7]) );
  XOR2_X1 U97 ( .A(B[14]), .B(A[14]), .Z(n74) );
  XOR2_X1 U98 ( .A(n31), .B(n74), .Z(SUM[14]) );
  NAND2_X1 U99 ( .A1(n56), .A2(B[14]), .ZN(n75) );
  NAND2_X1 U100 ( .A1(carry[14]), .A2(A[14]), .ZN(n76) );
  NAND2_X1 U101 ( .A1(B[14]), .A2(A[14]), .ZN(n77) );
  NAND3_X1 U102 ( .A1(n75), .A2(n76), .A3(n77), .ZN(carry[15]) );
  XOR2_X1 U103 ( .A(B[7]), .B(A[7]), .Z(n78) );
  XOR2_X1 U104 ( .A(n5), .B(n78), .Z(SUM[7]) );
  NAND2_X1 U105 ( .A1(n46), .A2(B[7]), .ZN(n79) );
  NAND2_X1 U106 ( .A1(carry[7]), .A2(A[7]), .ZN(n80) );
  NAND2_X1 U107 ( .A1(B[7]), .A2(A[7]), .ZN(n81) );
  NAND3_X1 U108 ( .A1(n79), .A2(n80), .A3(n81), .ZN(carry[8]) );
  XOR2_X1 U109 ( .A(B[0]), .B(n8), .Z(SUM[0]) );
endmodule


module mac_11_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n311), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n310), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n314), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n313), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n316), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n209), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  XOR2_X1 U157 ( .A(n70), .B(n87), .Z(n52) );
  XOR2_X1 U158 ( .A(n52), .B(n211), .Z(n50) );
  BUF_X1 U159 ( .A(n363), .Z(n206) );
  AND2_X1 U160 ( .A1(n104), .A2(n72), .ZN(n207) );
  AND2_X1 U161 ( .A1(n95), .A2(n215), .ZN(n208) );
  AND2_X1 U162 ( .A1(n70), .A2(n87), .ZN(n209) );
  CLKBUF_X1 U163 ( .A(n258), .Z(n210) );
  XOR2_X1 U164 ( .A(a[3]), .B(a[2]), .Z(n360) );
  XOR2_X2 U165 ( .A(a[6]), .B(n312), .Z(n343) );
  NAND2_X1 U166 ( .A1(n343), .A2(n362), .ZN(n345) );
  XOR2_X1 U167 ( .A(n100), .B(n93), .Z(n211) );
  NAND2_X1 U168 ( .A1(n52), .A2(n100), .ZN(n212) );
  NAND2_X1 U169 ( .A1(n52), .A2(n93), .ZN(n213) );
  NAND2_X1 U170 ( .A1(n100), .A2(n93), .ZN(n214) );
  NAND3_X1 U171 ( .A1(n212), .A2(n213), .A3(n214), .ZN(n49) );
  CLKBUF_X1 U172 ( .A(n102), .Z(n215) );
  CLKBUF_X1 U173 ( .A(n281), .Z(n216) );
  CLKBUF_X1 U174 ( .A(n273), .Z(n217) );
  NAND2_X1 U175 ( .A1(n207), .A2(n96), .ZN(n218) );
  NAND2_X1 U176 ( .A1(n207), .A2(n96), .ZN(n219) );
  CLKBUF_X1 U177 ( .A(b[1]), .Z(n220) );
  XNOR2_X2 U178 ( .A(a[2]), .B(a[1]), .ZN(n221) );
  XNOR2_X1 U179 ( .A(a[2]), .B(a[1]), .ZN(n324) );
  NAND3_X1 U180 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n222) );
  NAND3_X1 U181 ( .A1(n239), .A2(n219), .A3(n241), .ZN(n223) );
  NAND3_X1 U182 ( .A1(n277), .A2(n278), .A3(n279), .ZN(n224) );
  NAND3_X1 U183 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n225) );
  NAND3_X1 U184 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n226) );
  CLKBUF_X1 U185 ( .A(n242), .Z(n227) );
  CLKBUF_X1 U186 ( .A(n272), .Z(n228) );
  NAND3_X1 U187 ( .A1(n217), .A2(n228), .A3(n274), .ZN(n229) );
  CLKBUF_X1 U188 ( .A(n233), .Z(n230) );
  XNOR2_X1 U189 ( .A(a[4]), .B(a[3]), .ZN(n332) );
  AND2_X1 U190 ( .A1(n104), .A2(n72), .ZN(n231) );
  NAND2_X2 U191 ( .A1(n332), .A2(n361), .ZN(n334) );
  BUF_X2 U192 ( .A(n332), .Z(n286) );
  CLKBUF_X1 U193 ( .A(n255), .Z(n232) );
  NAND3_X1 U194 ( .A1(n300), .A2(n302), .A3(n301), .ZN(n233) );
  XNOR2_X1 U195 ( .A(a[3]), .B(n306), .ZN(n287) );
  XOR2_X1 U196 ( .A(n54), .B(n208), .Z(n234) );
  XOR2_X1 U197 ( .A(n230), .B(n234), .Z(product[4]) );
  NAND2_X1 U198 ( .A1(n233), .A2(n54), .ZN(n235) );
  NAND2_X1 U199 ( .A1(n12), .A2(n208), .ZN(n236) );
  NAND2_X1 U200 ( .A1(n54), .A2(n208), .ZN(n237) );
  NAND3_X1 U201 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n11) );
  XOR2_X1 U202 ( .A(n102), .B(n95), .Z(n56) );
  XOR2_X1 U203 ( .A(n103), .B(n96), .Z(n238) );
  XOR2_X1 U204 ( .A(n231), .B(n238), .Z(product[2]) );
  NAND2_X1 U205 ( .A1(n231), .A2(n103), .ZN(n239) );
  NAND2_X1 U206 ( .A1(n14), .A2(n96), .ZN(n240) );
  NAND2_X1 U207 ( .A1(n103), .A2(n96), .ZN(n241) );
  NAND3_X1 U208 ( .A1(n239), .A2(n218), .A3(n241), .ZN(n13) );
  NAND3_X1 U209 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n242) );
  AND3_X1 U210 ( .A1(n265), .A2(n266), .A3(n267), .ZN(product[15]) );
  XOR2_X1 U211 ( .A(n20), .B(n23), .Z(n244) );
  XOR2_X1 U212 ( .A(n229), .B(n244), .Z(product[11]) );
  NAND2_X1 U213 ( .A1(n5), .A2(n20), .ZN(n245) );
  NAND2_X1 U214 ( .A1(n5), .A2(n23), .ZN(n246) );
  NAND2_X1 U215 ( .A1(n20), .A2(n23), .ZN(n247) );
  NAND3_X1 U216 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n4) );
  NAND3_X1 U217 ( .A1(n251), .A2(n253), .A3(n252), .ZN(n248) );
  NAND3_X1 U218 ( .A1(n232), .A2(n256), .A3(n257), .ZN(n249) );
  XOR2_X1 U219 ( .A(n50), .B(n53), .Z(n250) );
  XOR2_X1 U220 ( .A(n11), .B(n250), .Z(product[5]) );
  NAND2_X1 U221 ( .A1(n11), .A2(n50), .ZN(n251) );
  NAND2_X1 U222 ( .A1(n226), .A2(n53), .ZN(n252) );
  NAND2_X1 U223 ( .A1(n50), .A2(n53), .ZN(n253) );
  NAND3_X1 U224 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n10) );
  XOR2_X1 U225 ( .A(n18), .B(n19), .Z(n254) );
  XOR2_X1 U226 ( .A(n227), .B(n254), .Z(product[12]) );
  NAND2_X1 U227 ( .A1(n242), .A2(n18), .ZN(n255) );
  NAND2_X1 U228 ( .A1(n4), .A2(n19), .ZN(n256) );
  NAND2_X1 U229 ( .A1(n18), .A2(n19), .ZN(n257) );
  NAND3_X1 U230 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n3) );
  NAND3_X1 U231 ( .A1(n290), .A2(n291), .A3(n292), .ZN(n258) );
  NAND3_X1 U232 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n259) );
  XOR2_X1 U233 ( .A(n17), .B(n307), .Z(n260) );
  XOR2_X1 U234 ( .A(n260), .B(n249), .Z(product[13]) );
  NAND2_X1 U235 ( .A1(n17), .A2(n307), .ZN(n261) );
  NAND2_X1 U236 ( .A1(n3), .A2(n17), .ZN(n262) );
  NAND2_X1 U237 ( .A1(n3), .A2(n307), .ZN(n263) );
  NAND3_X1 U238 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n2) );
  XOR2_X1 U239 ( .A(n308), .B(n15), .Z(n264) );
  XOR2_X1 U240 ( .A(n264), .B(n259), .Z(product[14]) );
  NAND2_X1 U241 ( .A1(n308), .A2(n15), .ZN(n265) );
  NAND2_X1 U242 ( .A1(n2), .A2(n308), .ZN(n266) );
  NAND2_X1 U243 ( .A1(n2), .A2(n15), .ZN(n267) );
  NAND3_X1 U244 ( .A1(n281), .A2(n282), .A3(n283), .ZN(n268) );
  NAND3_X1 U245 ( .A1(n216), .A2(n282), .A3(n283), .ZN(n269) );
  CLKBUF_X1 U246 ( .A(n225), .Z(n270) );
  XOR2_X1 U247 ( .A(n27), .B(n24), .Z(n271) );
  XOR2_X1 U248 ( .A(n269), .B(n271), .Z(product[10]) );
  NAND2_X1 U249 ( .A1(n268), .A2(n27), .ZN(n272) );
  NAND2_X1 U250 ( .A1(n6), .A2(n24), .ZN(n273) );
  NAND2_X1 U251 ( .A1(n27), .A2(n24), .ZN(n274) );
  NAND3_X1 U252 ( .A1(n273), .A2(n272), .A3(n274), .ZN(n5) );
  CLKBUF_X1 U253 ( .A(n7), .Z(n275) );
  XOR2_X1 U254 ( .A(n34), .B(n39), .Z(n276) );
  XOR2_X1 U255 ( .A(n270), .B(n276), .Z(product[8]) );
  NAND2_X1 U256 ( .A1(n225), .A2(n34), .ZN(n277) );
  NAND2_X1 U257 ( .A1(n8), .A2(n39), .ZN(n278) );
  NAND2_X1 U258 ( .A1(n34), .A2(n39), .ZN(n279) );
  NAND3_X1 U259 ( .A1(n277), .A2(n278), .A3(n279), .ZN(n7) );
  XOR2_X1 U260 ( .A(n33), .B(n28), .Z(n280) );
  XOR2_X1 U261 ( .A(n275), .B(n280), .Z(product[9]) );
  NAND2_X1 U262 ( .A1(n7), .A2(n33), .ZN(n281) );
  NAND2_X1 U263 ( .A1(n224), .A2(n28), .ZN(n282) );
  NAND2_X1 U264 ( .A1(n33), .A2(n28), .ZN(n283) );
  NAND3_X1 U265 ( .A1(n282), .A2(n281), .A3(n283), .ZN(n6) );
  INV_X1 U266 ( .A(n306), .ZN(n284) );
  CLKBUF_X1 U267 ( .A(n56), .Z(n285) );
  INV_X1 U268 ( .A(n15), .ZN(n307) );
  INV_X1 U269 ( .A(n21), .ZN(n310) );
  INV_X1 U270 ( .A(n341), .ZN(n311) );
  INV_X1 U271 ( .A(n323), .ZN(n316) );
  INV_X1 U272 ( .A(n330), .ZN(n314) );
  INV_X1 U273 ( .A(n31), .ZN(n313) );
  INV_X1 U274 ( .A(b[0]), .ZN(n306) );
  INV_X1 U275 ( .A(n352), .ZN(n308) );
  INV_X1 U276 ( .A(a[0]), .ZN(n318) );
  INV_X1 U277 ( .A(a[5]), .ZN(n312) );
  INV_X1 U278 ( .A(a[7]), .ZN(n309) );
  NAND2_X1 U279 ( .A1(n287), .A2(n288), .ZN(n303) );
  AND2_X1 U280 ( .A1(n324), .A2(n360), .ZN(n288) );
  XOR2_X1 U281 ( .A(n46), .B(n49), .Z(n289) );
  XOR2_X1 U282 ( .A(n10), .B(n289), .Z(product[6]) );
  NAND2_X1 U283 ( .A1(n248), .A2(n46), .ZN(n290) );
  NAND2_X1 U284 ( .A1(n248), .A2(n49), .ZN(n291) );
  NAND2_X1 U285 ( .A1(n46), .A2(n49), .ZN(n292) );
  NAND3_X1 U286 ( .A1(n290), .A2(n291), .A3(n292), .ZN(n9) );
  XOR2_X1 U287 ( .A(n40), .B(n45), .Z(n293) );
  XOR2_X1 U288 ( .A(n210), .B(n293), .Z(product[7]) );
  NAND2_X1 U289 ( .A1(n258), .A2(n40), .ZN(n294) );
  NAND2_X1 U290 ( .A1(n9), .A2(n45), .ZN(n295) );
  NAND2_X1 U291 ( .A1(n40), .A2(n45), .ZN(n296) );
  NAND3_X1 U292 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n8) );
  NAND2_X1 U293 ( .A1(n324), .A2(n360), .ZN(n297) );
  NAND2_X1 U294 ( .A1(n221), .A2(n360), .ZN(n298) );
  XOR2_X1 U295 ( .A(n223), .B(n71), .Z(n299) );
  XOR2_X1 U296 ( .A(n285), .B(n299), .Z(product[3]) );
  NAND2_X1 U297 ( .A1(n56), .A2(n13), .ZN(n300) );
  NAND2_X1 U298 ( .A1(n56), .A2(n71), .ZN(n301) );
  NAND2_X1 U299 ( .A1(n222), .A2(n71), .ZN(n302) );
  NAND3_X1 U300 ( .A1(n300), .A2(n302), .A3(n301), .ZN(n12) );
  OR2_X1 U301 ( .A1(n221), .A2(n325), .ZN(n304) );
  NAND2_X1 U302 ( .A1(n303), .A2(n304), .ZN(n95) );
  INV_X1 U303 ( .A(a[3]), .ZN(n315) );
  INV_X1 U304 ( .A(a[1]), .ZN(n317) );
  INV_X1 U305 ( .A(n306), .ZN(n305) );
  NOR2_X1 U306 ( .A1(n318), .A2(n306), .ZN(product[0]) );
  OAI22_X1 U307 ( .A1(n319), .A2(n320), .B1(n321), .B2(n318), .ZN(n99) );
  OAI22_X1 U308 ( .A1(n321), .A2(n320), .B1(n322), .B2(n318), .ZN(n98) );
  XNOR2_X1 U309 ( .A(b[6]), .B(a[1]), .ZN(n321) );
  OAI22_X1 U310 ( .A1(n318), .A2(n322), .B1(n320), .B2(n322), .ZN(n323) );
  XNOR2_X1 U311 ( .A(b[7]), .B(a[1]), .ZN(n322) );
  NOR2_X1 U312 ( .A1(n221), .A2(n306), .ZN(n96) );
  OAI22_X1 U313 ( .A1(n325), .A2(n297), .B1(n221), .B2(n326), .ZN(n94) );
  XNOR2_X1 U314 ( .A(b[1]), .B(a[3]), .ZN(n325) );
  OAI22_X1 U315 ( .A1(n326), .A2(n297), .B1(n221), .B2(n327), .ZN(n93) );
  XNOR2_X1 U316 ( .A(b[2]), .B(a[3]), .ZN(n326) );
  OAI22_X1 U317 ( .A1(n327), .A2(n298), .B1(n221), .B2(n328), .ZN(n92) );
  XNOR2_X1 U318 ( .A(b[3]), .B(a[3]), .ZN(n327) );
  OAI22_X1 U319 ( .A1(n328), .A2(n297), .B1(n221), .B2(n329), .ZN(n91) );
  XNOR2_X1 U320 ( .A(b[4]), .B(a[3]), .ZN(n328) );
  OAI22_X1 U321 ( .A1(n331), .A2(n221), .B1(n297), .B2(n331), .ZN(n330) );
  NOR2_X1 U322 ( .A1(n286), .A2(n306), .ZN(n88) );
  OAI22_X1 U323 ( .A1(n333), .A2(n334), .B1(n286), .B2(n335), .ZN(n87) );
  XNOR2_X1 U324 ( .A(a[5]), .B(n284), .ZN(n333) );
  OAI22_X1 U325 ( .A1(n335), .A2(n334), .B1(n286), .B2(n336), .ZN(n86) );
  XNOR2_X1 U326 ( .A(n220), .B(a[5]), .ZN(n335) );
  OAI22_X1 U327 ( .A1(n336), .A2(n334), .B1(n286), .B2(n337), .ZN(n85) );
  XNOR2_X1 U328 ( .A(b[2]), .B(a[5]), .ZN(n336) );
  OAI22_X1 U329 ( .A1(n337), .A2(n334), .B1(n286), .B2(n338), .ZN(n84) );
  XNOR2_X1 U330 ( .A(b[3]), .B(a[5]), .ZN(n337) );
  OAI22_X1 U331 ( .A1(n338), .A2(n334), .B1(n286), .B2(n339), .ZN(n83) );
  XNOR2_X1 U332 ( .A(b[4]), .B(a[5]), .ZN(n338) );
  OAI22_X1 U333 ( .A1(n339), .A2(n334), .B1(n286), .B2(n340), .ZN(n82) );
  XNOR2_X1 U334 ( .A(b[5]), .B(a[5]), .ZN(n339) );
  OAI22_X1 U335 ( .A1(n342), .A2(n286), .B1(n334), .B2(n342), .ZN(n341) );
  NOR2_X1 U336 ( .A1(n343), .A2(n306), .ZN(n80) );
  OAI22_X1 U337 ( .A1(n344), .A2(n345), .B1(n343), .B2(n346), .ZN(n79) );
  XNOR2_X1 U338 ( .A(a[7]), .B(n284), .ZN(n344) );
  OAI22_X1 U339 ( .A1(n347), .A2(n345), .B1(n343), .B2(n348), .ZN(n77) );
  OAI22_X1 U340 ( .A1(n348), .A2(n345), .B1(n343), .B2(n349), .ZN(n76) );
  XNOR2_X1 U341 ( .A(b[3]), .B(a[7]), .ZN(n348) );
  OAI22_X1 U342 ( .A1(n349), .A2(n345), .B1(n343), .B2(n350), .ZN(n75) );
  XNOR2_X1 U343 ( .A(b[4]), .B(a[7]), .ZN(n349) );
  OAI22_X1 U344 ( .A1(n350), .A2(n345), .B1(n343), .B2(n351), .ZN(n74) );
  XNOR2_X1 U345 ( .A(b[5]), .B(a[7]), .ZN(n350) );
  OAI22_X1 U346 ( .A1(n353), .A2(n343), .B1(n345), .B2(n353), .ZN(n352) );
  OAI21_X1 U347 ( .B1(n305), .B2(n317), .A(n320), .ZN(n72) );
  OAI21_X1 U348 ( .B1(n315), .B2(n298), .A(n354), .ZN(n71) );
  OR3_X1 U349 ( .A1(n221), .A2(n284), .A3(n315), .ZN(n354) );
  OAI21_X1 U350 ( .B1(n334), .B2(n312), .A(n355), .ZN(n70) );
  OR3_X1 U351 ( .A1(n332), .A2(n284), .A3(n312), .ZN(n355) );
  OAI21_X1 U352 ( .B1(n309), .B2(n345), .A(n356), .ZN(n69) );
  OR3_X1 U353 ( .A1(n343), .A2(n284), .A3(n309), .ZN(n356) );
  XNOR2_X1 U354 ( .A(n357), .B(n358), .ZN(n38) );
  OR2_X1 U355 ( .A1(n357), .A2(n358), .ZN(n37) );
  OAI22_X1 U356 ( .A1(n329), .A2(n298), .B1(n221), .B2(n359), .ZN(n358) );
  XNOR2_X1 U357 ( .A(b[5]), .B(a[3]), .ZN(n329) );
  OAI22_X1 U358 ( .A1(n346), .A2(n345), .B1(n343), .B2(n347), .ZN(n357) );
  XNOR2_X1 U359 ( .A(b[2]), .B(a[7]), .ZN(n347) );
  XNOR2_X1 U360 ( .A(n220), .B(a[7]), .ZN(n346) );
  OAI22_X1 U361 ( .A1(n359), .A2(n298), .B1(n221), .B2(n331), .ZN(n31) );
  XNOR2_X1 U362 ( .A(b[7]), .B(a[3]), .ZN(n331) );
  XNOR2_X1 U363 ( .A(b[6]), .B(a[3]), .ZN(n359) );
  OAI22_X1 U364 ( .A1(n340), .A2(n334), .B1(n286), .B2(n342), .ZN(n21) );
  XNOR2_X1 U365 ( .A(b[7]), .B(a[5]), .ZN(n342) );
  XNOR2_X1 U366 ( .A(n312), .B(a[4]), .ZN(n361) );
  XNOR2_X1 U367 ( .A(b[6]), .B(a[5]), .ZN(n340) );
  OAI22_X1 U368 ( .A1(n351), .A2(n345), .B1(n343), .B2(n353), .ZN(n15) );
  XNOR2_X1 U369 ( .A(b[7]), .B(a[7]), .ZN(n353) );
  XNOR2_X1 U370 ( .A(n309), .B(a[6]), .ZN(n362) );
  XNOR2_X1 U371 ( .A(b[6]), .B(a[7]), .ZN(n351) );
  OAI22_X1 U372 ( .A1(n305), .A2(n320), .B1(n363), .B2(n318), .ZN(n104) );
  OAI22_X1 U373 ( .A1(n206), .A2(n320), .B1(n364), .B2(n318), .ZN(n103) );
  XNOR2_X1 U374 ( .A(b[1]), .B(a[1]), .ZN(n363) );
  OAI22_X1 U375 ( .A1(n364), .A2(n320), .B1(n365), .B2(n318), .ZN(n102) );
  XNOR2_X1 U376 ( .A(b[2]), .B(a[1]), .ZN(n364) );
  OAI22_X1 U377 ( .A1(n365), .A2(n320), .B1(n366), .B2(n318), .ZN(n101) );
  XNOR2_X1 U378 ( .A(b[3]), .B(a[1]), .ZN(n365) );
  OAI22_X1 U379 ( .A1(n366), .A2(n320), .B1(n319), .B2(n318), .ZN(n100) );
  XNOR2_X1 U380 ( .A(b[5]), .B(a[1]), .ZN(n319) );
  NAND2_X1 U381 ( .A1(a[1]), .A2(n318), .ZN(n320) );
  XNOR2_X1 U382 ( .A(b[4]), .B(a[1]), .ZN(n366) );
endmodule


module mac_11 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   n6, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, n2, n4;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(n6), .QN(n2) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_11_DW01_add_0 add_356 ( .A(pipeline), .B({mac_out[15:1], n6}), .CI(1'b0), 
        .SUM(sum) );
  mac_11_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X2 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n4), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n4), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n4), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n4), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n4), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n4), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n4), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n4), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n4), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n4), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n4), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n4), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n4), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n4), .ZN(N6) );
  INV_X1 U18 ( .A(n2), .ZN(mac_out[0]) );
  AND2_X1 U19 ( .A1(sum[0]), .A2(n4), .ZN(N3) );
  AND2_X1 U20 ( .A1(sum[15]), .A2(n4), .ZN(N18) );
  INV_X1 U21 ( .A(clear_acc), .ZN(n4) );
endmodule


module mac_10_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72;
  wire   [15:1] carry;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n72) );
  XOR2_X1 U2 ( .A(B[15]), .B(A[15]), .Z(n1) );
  XOR2_X1 U3 ( .A(carry[15]), .B(n1), .Z(SUM[15]) );
  NAND2_X1 U4 ( .A1(carry[9]), .A2(A[9]), .ZN(n2) );
  NAND3_X1 U5 ( .A1(n69), .A2(n70), .A3(n71), .ZN(n3) );
  NAND3_X1 U6 ( .A1(n69), .A2(n70), .A3(n71), .ZN(n4) );
  XOR2_X1 U7 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR2_X1 U8 ( .A(n4), .B(n5), .Z(SUM[3]) );
  NAND2_X1 U9 ( .A1(n3), .A2(B[3]), .ZN(n6) );
  NAND2_X1 U10 ( .A1(carry[3]), .A2(A[3]), .ZN(n7) );
  NAND2_X1 U11 ( .A1(B[3]), .A2(A[3]), .ZN(n8) );
  NAND3_X1 U12 ( .A1(n6), .A2(n7), .A3(n8), .ZN(carry[4]) );
  NAND3_X1 U13 ( .A1(n61), .A2(n2), .A3(n63), .ZN(n9) );
  NAND3_X1 U14 ( .A1(n57), .A2(n58), .A3(n59), .ZN(n10) );
  NAND3_X1 U15 ( .A1(n28), .A2(n27), .A3(n29), .ZN(n11) );
  NAND3_X1 U16 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n12) );
  NAND3_X1 U17 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n13) );
  NAND3_X1 U18 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n14) );
  NAND3_X1 U19 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n15) );
  XOR2_X1 U20 ( .A(B[5]), .B(A[5]), .Z(n16) );
  XOR2_X1 U21 ( .A(carry[5]), .B(n16), .Z(SUM[5]) );
  NAND2_X1 U22 ( .A1(carry[5]), .A2(B[5]), .ZN(n17) );
  NAND2_X1 U23 ( .A1(carry[5]), .A2(A[5]), .ZN(n18) );
  NAND2_X1 U24 ( .A1(B[5]), .A2(A[5]), .ZN(n19) );
  NAND3_X1 U25 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[6]) );
  NAND3_X1 U26 ( .A1(n23), .A2(n24), .A3(n25), .ZN(n20) );
  NAND3_X1 U27 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n21) );
  XOR2_X1 U28 ( .A(B[6]), .B(A[6]), .Z(n22) );
  XOR2_X1 U29 ( .A(n15), .B(n22), .Z(SUM[6]) );
  NAND2_X1 U30 ( .A1(n14), .A2(B[6]), .ZN(n23) );
  NAND2_X1 U31 ( .A1(carry[6]), .A2(A[6]), .ZN(n24) );
  NAND2_X1 U32 ( .A1(B[6]), .A2(A[6]), .ZN(n25) );
  NAND3_X1 U33 ( .A1(n24), .A2(n23), .A3(n25), .ZN(carry[7]) );
  XOR2_X1 U34 ( .A(B[13]), .B(A[13]), .Z(n26) );
  XOR2_X1 U35 ( .A(n13), .B(n26), .Z(SUM[13]) );
  NAND2_X1 U36 ( .A1(n12), .A2(B[13]), .ZN(n27) );
  NAND2_X1 U37 ( .A1(carry[13]), .A2(A[13]), .ZN(n28) );
  NAND2_X1 U38 ( .A1(B[13]), .A2(A[13]), .ZN(n29) );
  NAND3_X1 U39 ( .A1(n27), .A2(n28), .A3(n29), .ZN(carry[14]) );
  XOR2_X1 U40 ( .A(B[14]), .B(A[14]), .Z(n30) );
  XOR2_X1 U41 ( .A(n11), .B(n30), .Z(SUM[14]) );
  NAND2_X1 U42 ( .A1(n11), .A2(B[14]), .ZN(n31) );
  NAND2_X1 U43 ( .A1(carry[14]), .A2(A[14]), .ZN(n32) );
  NAND2_X1 U44 ( .A1(B[14]), .A2(A[14]), .ZN(n33) );
  NAND3_X1 U45 ( .A1(n31), .A2(n32), .A3(n33), .ZN(carry[15]) );
  NAND3_X1 U46 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n34) );
  NAND3_X1 U47 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n35) );
  XOR2_X1 U48 ( .A(B[12]), .B(A[12]), .Z(n36) );
  XOR2_X1 U49 ( .A(n34), .B(n36), .Z(SUM[12]) );
  NAND2_X1 U50 ( .A1(n34), .A2(B[12]), .ZN(n37) );
  NAND2_X1 U51 ( .A1(carry[12]), .A2(A[12]), .ZN(n38) );
  NAND2_X1 U52 ( .A1(B[12]), .A2(A[12]), .ZN(n39) );
  NAND3_X1 U53 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[13]) );
  XOR2_X1 U54 ( .A(B[7]), .B(A[7]), .Z(n40) );
  XOR2_X1 U55 ( .A(n20), .B(n40), .Z(SUM[7]) );
  NAND2_X1 U56 ( .A1(n20), .A2(B[7]), .ZN(n41) );
  NAND2_X1 U57 ( .A1(carry[7]), .A2(A[7]), .ZN(n42) );
  NAND2_X1 U58 ( .A1(B[7]), .A2(A[7]), .ZN(n43) );
  NAND3_X1 U59 ( .A1(n41), .A2(n42), .A3(n43), .ZN(carry[8]) );
  NAND3_X1 U60 ( .A1(n61), .A2(n2), .A3(n63), .ZN(n44) );
  XOR2_X1 U61 ( .A(B[10]), .B(A[10]), .Z(n45) );
  XOR2_X1 U62 ( .A(n44), .B(n45), .Z(SUM[10]) );
  NAND2_X1 U63 ( .A1(n9), .A2(B[10]), .ZN(n46) );
  NAND2_X1 U64 ( .A1(carry[10]), .A2(A[10]), .ZN(n47) );
  NAND2_X1 U65 ( .A1(B[10]), .A2(A[10]), .ZN(n48) );
  NAND3_X1 U66 ( .A1(n47), .A2(n46), .A3(n48), .ZN(carry[11]) );
  XOR2_X1 U67 ( .A(B[11]), .B(A[11]), .Z(n49) );
  XOR2_X1 U68 ( .A(n21), .B(n49), .Z(SUM[11]) );
  NAND2_X1 U69 ( .A1(n21), .A2(B[11]), .ZN(n50) );
  NAND2_X1 U70 ( .A1(carry[11]), .A2(A[11]), .ZN(n51) );
  NAND2_X1 U71 ( .A1(B[11]), .A2(A[11]), .ZN(n52) );
  NAND3_X1 U72 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[12]) );
  NAND3_X1 U73 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n53) );
  NAND3_X1 U74 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n54) );
  NAND3_X1 U75 ( .A1(n57), .A2(n58), .A3(n59), .ZN(n55) );
  XOR2_X1 U76 ( .A(B[8]), .B(A[8]), .Z(n56) );
  XOR2_X1 U77 ( .A(n35), .B(n56), .Z(SUM[8]) );
  NAND2_X1 U78 ( .A1(n35), .A2(B[8]), .ZN(n57) );
  NAND2_X1 U79 ( .A1(carry[8]), .A2(A[8]), .ZN(n58) );
  NAND2_X1 U80 ( .A1(B[8]), .A2(A[8]), .ZN(n59) );
  NAND3_X1 U81 ( .A1(n57), .A2(n58), .A3(n59), .ZN(carry[9]) );
  XOR2_X1 U82 ( .A(B[9]), .B(A[9]), .Z(n60) );
  XOR2_X1 U83 ( .A(n55), .B(n60), .Z(SUM[9]) );
  NAND2_X1 U84 ( .A1(n10), .A2(B[9]), .ZN(n61) );
  NAND2_X1 U85 ( .A1(carry[9]), .A2(A[9]), .ZN(n62) );
  NAND2_X1 U86 ( .A1(B[9]), .A2(A[9]), .ZN(n63) );
  NAND3_X1 U87 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[10]) );
  XOR2_X1 U88 ( .A(B[1]), .B(A[1]), .Z(n64) );
  XOR2_X1 U89 ( .A(n72), .B(n64), .Z(SUM[1]) );
  NAND2_X1 U90 ( .A1(n72), .A2(B[1]), .ZN(n65) );
  NAND2_X1 U91 ( .A1(n72), .A2(A[1]), .ZN(n66) );
  NAND2_X1 U92 ( .A1(B[1]), .A2(A[1]), .ZN(n67) );
  NAND3_X1 U93 ( .A1(n65), .A2(n66), .A3(n67), .ZN(carry[2]) );
  XOR2_X1 U94 ( .A(B[2]), .B(A[2]), .Z(n68) );
  XOR2_X1 U95 ( .A(n54), .B(n68), .Z(SUM[2]) );
  NAND2_X1 U96 ( .A1(n53), .A2(B[2]), .ZN(n69) );
  NAND2_X1 U97 ( .A1(carry[2]), .A2(A[2]), .ZN(n70) );
  NAND2_X1 U98 ( .A1(B[2]), .A2(A[2]), .ZN(n71) );
  NAND3_X1 U99 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[3]) );
  XOR2_X1 U100 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_10_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n314), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n313), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n317), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n316), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n319), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  NAND3_X1 U157 ( .A1(n209), .A2(n210), .A3(n211), .ZN(n206) );
  NOR2_X1 U158 ( .A1(n291), .A2(n309), .ZN(n96) );
  CLKBUF_X1 U159 ( .A(n264), .Z(n207) );
  XOR2_X1 U160 ( .A(n103), .B(n96), .Z(n208) );
  XOR2_X1 U161 ( .A(n14), .B(n208), .Z(product[2]) );
  NAND2_X1 U162 ( .A1(n14), .A2(n103), .ZN(n209) );
  NAND2_X1 U163 ( .A1(n14), .A2(n96), .ZN(n210) );
  NAND2_X1 U164 ( .A1(n103), .A2(n96), .ZN(n211) );
  NAND3_X1 U165 ( .A1(n209), .A2(n210), .A3(n211), .ZN(n13) );
  AND2_X1 U166 ( .A1(n279), .A2(n102), .ZN(n212) );
  CLKBUF_X1 U167 ( .A(n273), .Z(n213) );
  CLKBUF_X1 U168 ( .A(n56), .Z(n214) );
  NAND3_X1 U169 ( .A1(n213), .A2(n274), .A3(n275), .ZN(n215) );
  CLKBUF_X1 U170 ( .A(n220), .Z(n216) );
  CLKBUF_X1 U171 ( .A(n206), .Z(n217) );
  NAND2_X1 U172 ( .A1(n6), .A2(n27), .ZN(n218) );
  CLKBUF_X1 U173 ( .A(n241), .Z(n219) );
  NAND3_X1 U174 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n220) );
  NAND2_X2 U175 ( .A1(n348), .A2(n367), .ZN(n350) );
  XOR2_X2 U176 ( .A(a[6]), .B(n315), .Z(n348) );
  CLKBUF_X1 U177 ( .A(n231), .Z(n221) );
  NAND3_X1 U178 ( .A1(n269), .A2(n268), .A3(n270), .ZN(n222) );
  XOR2_X1 U179 ( .A(n100), .B(n93), .Z(n223) );
  XOR2_X1 U180 ( .A(n52), .B(n223), .Z(n50) );
  NAND2_X1 U181 ( .A1(n227), .A2(n100), .ZN(n224) );
  NAND2_X1 U182 ( .A1(n227), .A2(n93), .ZN(n225) );
  NAND2_X1 U183 ( .A1(n100), .A2(n93), .ZN(n226) );
  NAND3_X1 U184 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n49) );
  XOR2_X1 U185 ( .A(n70), .B(n87), .Z(n227) );
  CLKBUF_X1 U186 ( .A(n301), .Z(n228) );
  CLKBUF_X1 U187 ( .A(n253), .Z(n229) );
  CLKBUF_X1 U188 ( .A(n218), .Z(n230) );
  NAND3_X1 U189 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n231) );
  CLKBUF_X1 U190 ( .A(n288), .Z(n232) );
  NAND3_X1 U191 ( .A1(n229), .A2(n254), .A3(n255), .ZN(n233) );
  XOR2_X1 U192 ( .A(n54), .B(n212), .Z(n234) );
  XOR2_X1 U193 ( .A(n216), .B(n234), .Z(product[4]) );
  NAND2_X1 U194 ( .A1(n220), .A2(n54), .ZN(n235) );
  NAND2_X1 U195 ( .A1(n12), .A2(n212), .ZN(n236) );
  NAND2_X1 U196 ( .A1(n54), .A2(n212), .ZN(n237) );
  NAND3_X1 U197 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n11) );
  NAND2_X2 U198 ( .A1(n337), .A2(n366), .ZN(n339) );
  CLKBUF_X1 U199 ( .A(n269), .Z(n238) );
  NAND3_X1 U200 ( .A1(n264), .A2(n218), .A3(n265), .ZN(n239) );
  NAND3_X1 U201 ( .A1(n207), .A2(n230), .A3(n265), .ZN(n240) );
  NAND3_X1 U202 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n241) );
  XOR2_X1 U203 ( .A(n20), .B(n23), .Z(n242) );
  XOR2_X1 U204 ( .A(n240), .B(n242), .Z(product[11]) );
  NAND2_X1 U205 ( .A1(n239), .A2(n20), .ZN(n243) );
  NAND2_X1 U206 ( .A1(n5), .A2(n23), .ZN(n244) );
  NAND2_X1 U207 ( .A1(n20), .A2(n23), .ZN(n245) );
  NAND3_X1 U208 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n4) );
  NAND3_X1 U209 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n246) );
  XOR2_X1 U210 ( .A(n214), .B(n71), .Z(n247) );
  XOR2_X1 U211 ( .A(n217), .B(n247), .Z(product[3]) );
  NAND2_X1 U212 ( .A1(n206), .A2(n56), .ZN(n248) );
  NAND2_X1 U213 ( .A1(n13), .A2(n71), .ZN(n249) );
  NAND2_X1 U214 ( .A1(n56), .A2(n71), .ZN(n250) );
  NAND3_X1 U215 ( .A1(n249), .A2(n248), .A3(n250), .ZN(n12) );
  CLKBUF_X1 U216 ( .A(n7), .Z(n251) );
  XOR2_X1 U217 ( .A(n18), .B(n19), .Z(n252) );
  XOR2_X1 U218 ( .A(n219), .B(n252), .Z(product[12]) );
  NAND2_X1 U219 ( .A1(n241), .A2(n18), .ZN(n253) );
  NAND2_X1 U220 ( .A1(n4), .A2(n19), .ZN(n254) );
  NAND2_X1 U221 ( .A1(n18), .A2(n19), .ZN(n255) );
  NAND3_X1 U222 ( .A1(n238), .A2(n268), .A3(n270), .ZN(n256) );
  NAND3_X1 U223 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n257) );
  AND3_X1 U224 ( .A1(n287), .A2(n286), .A3(n285), .ZN(product[15]) );
  NAND2_X1 U225 ( .A1(b[3]), .A2(a[1]), .ZN(n260) );
  NAND2_X1 U226 ( .A1(n259), .A2(n320), .ZN(n261) );
  NAND2_X1 U227 ( .A1(n260), .A2(n261), .ZN(n370) );
  INV_X1 U228 ( .A(b[3]), .ZN(n259) );
  XOR2_X1 U229 ( .A(n27), .B(n24), .Z(n262) );
  XOR2_X1 U230 ( .A(n256), .B(n262), .Z(product[10]) );
  NAND2_X1 U231 ( .A1(n6), .A2(n27), .ZN(n263) );
  NAND2_X1 U232 ( .A1(n222), .A2(n24), .ZN(n264) );
  NAND2_X1 U233 ( .A1(n27), .A2(n24), .ZN(n265) );
  NAND3_X1 U234 ( .A1(n264), .A2(n263), .A3(n265), .ZN(n5) );
  NAND3_X1 U235 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n266) );
  XOR2_X1 U236 ( .A(n33), .B(n28), .Z(n267) );
  XOR2_X1 U237 ( .A(n251), .B(n267), .Z(product[9]) );
  NAND2_X1 U238 ( .A1(n266), .A2(n33), .ZN(n268) );
  NAND2_X1 U239 ( .A1(n7), .A2(n28), .ZN(n269) );
  NAND2_X1 U240 ( .A1(n33), .A2(n28), .ZN(n270) );
  NAND3_X1 U241 ( .A1(n269), .A2(n268), .A3(n270), .ZN(n6) );
  INV_X1 U242 ( .A(n309), .ZN(n271) );
  INV_X1 U243 ( .A(n309), .ZN(n308) );
  XOR2_X1 U244 ( .A(n276), .B(a[3]), .Z(n330) );
  CLKBUF_X1 U245 ( .A(n95), .Z(n279) );
  XOR2_X1 U246 ( .A(n50), .B(n53), .Z(n272) );
  XOR2_X1 U247 ( .A(n221), .B(n272), .Z(product[5]) );
  NAND2_X1 U248 ( .A1(n231), .A2(n50), .ZN(n273) );
  NAND2_X1 U249 ( .A1(n11), .A2(n53), .ZN(n274) );
  NAND2_X1 U250 ( .A1(n50), .A2(n53), .ZN(n275) );
  NAND3_X1 U251 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n10) );
  INV_X1 U252 ( .A(b[1]), .ZN(n276) );
  INV_X1 U253 ( .A(n276), .ZN(n277) );
  XNOR2_X1 U254 ( .A(a[2]), .B(a[1]), .ZN(n327) );
  NAND3_X1 U255 ( .A1(n282), .A2(n281), .A3(n283), .ZN(n278) );
  XOR2_X1 U256 ( .A(n95), .B(n102), .Z(n56) );
  XOR2_X1 U257 ( .A(n17), .B(n310), .Z(n280) );
  XOR2_X1 U258 ( .A(n280), .B(n233), .Z(product[13]) );
  NAND2_X1 U259 ( .A1(n17), .A2(n310), .ZN(n281) );
  NAND2_X1 U260 ( .A1(n246), .A2(n17), .ZN(n282) );
  NAND2_X1 U261 ( .A1(n310), .A2(n246), .ZN(n283) );
  NAND3_X1 U262 ( .A1(n283), .A2(n282), .A3(n281), .ZN(n2) );
  XOR2_X1 U263 ( .A(n311), .B(n15), .Z(n284) );
  XOR2_X1 U264 ( .A(n278), .B(n284), .Z(product[14]) );
  NAND2_X1 U265 ( .A1(n311), .A2(n15), .ZN(n285) );
  NAND2_X1 U266 ( .A1(n2), .A2(n311), .ZN(n286) );
  NAND2_X1 U267 ( .A1(n2), .A2(n15), .ZN(n287) );
  NAND3_X1 U268 ( .A1(n305), .A2(n306), .A3(n307), .ZN(n288) );
  NAND3_X1 U269 ( .A1(n301), .A2(n302), .A3(n303), .ZN(n289) );
  NAND3_X1 U270 ( .A1(n228), .A2(n302), .A3(n303), .ZN(n290) );
  NAND2_X2 U271 ( .A1(n327), .A2(n365), .ZN(n329) );
  XNOR2_X2 U272 ( .A(a[4]), .B(a[3]), .ZN(n337) );
  XOR2_X1 U273 ( .A(n290), .B(n304), .Z(product[7]) );
  XOR2_X1 U274 ( .A(a[2]), .B(n320), .Z(n291) );
  XOR2_X1 U275 ( .A(a[2]), .B(n320), .Z(n292) );
  INV_X1 U276 ( .A(n15), .ZN(n310) );
  INV_X1 U277 ( .A(n335), .ZN(n317) );
  INV_X1 U278 ( .A(n21), .ZN(n313) );
  INV_X1 U279 ( .A(n346), .ZN(n314) );
  INV_X1 U280 ( .A(n326), .ZN(n319) );
  INV_X1 U281 ( .A(b[0]), .ZN(n309) );
  INV_X1 U282 ( .A(n357), .ZN(n311) );
  INV_X1 U283 ( .A(n31), .ZN(n316) );
  INV_X1 U284 ( .A(a[0]), .ZN(n321) );
  INV_X1 U285 ( .A(a[5]), .ZN(n315) );
  INV_X1 U286 ( .A(a[7]), .ZN(n312) );
  XOR2_X1 U287 ( .A(n34), .B(n39), .Z(n293) );
  XOR2_X1 U288 ( .A(n232), .B(n293), .Z(product[8]) );
  NAND2_X1 U289 ( .A1(n288), .A2(n34), .ZN(n294) );
  NAND2_X1 U290 ( .A1(n8), .A2(n39), .ZN(n295) );
  NAND2_X1 U291 ( .A1(n34), .A2(n39), .ZN(n296) );
  NAND3_X1 U292 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n7) );
  NAND2_X1 U293 ( .A1(b[1]), .A2(a[1]), .ZN(n298) );
  NAND2_X1 U294 ( .A1(n297), .A2(n320), .ZN(n299) );
  NAND2_X1 U295 ( .A1(n299), .A2(n298), .ZN(n368) );
  INV_X1 U296 ( .A(b[1]), .ZN(n297) );
  INV_X1 U297 ( .A(a[3]), .ZN(n318) );
  XOR2_X1 U298 ( .A(n46), .B(n49), .Z(n300) );
  XOR2_X1 U299 ( .A(n215), .B(n300), .Z(product[6]) );
  NAND2_X1 U300 ( .A1(n257), .A2(n46), .ZN(n301) );
  NAND2_X1 U301 ( .A1(n10), .A2(n49), .ZN(n302) );
  NAND2_X1 U302 ( .A1(n46), .A2(n49), .ZN(n303) );
  NAND3_X1 U303 ( .A1(n302), .A2(n301), .A3(n303), .ZN(n9) );
  XOR2_X1 U304 ( .A(n40), .B(n45), .Z(n304) );
  NAND2_X1 U305 ( .A1(n289), .A2(n40), .ZN(n305) );
  NAND2_X1 U306 ( .A1(n9), .A2(n45), .ZN(n306) );
  NAND2_X1 U307 ( .A1(n40), .A2(n45), .ZN(n307) );
  NAND3_X1 U308 ( .A1(n306), .A2(n305), .A3(n307), .ZN(n8) );
  INV_X1 U309 ( .A(a[1]), .ZN(n320) );
  NOR2_X1 U310 ( .A1(n321), .A2(n309), .ZN(product[0]) );
  OAI22_X1 U311 ( .A1(n322), .A2(n323), .B1(n324), .B2(n321), .ZN(n99) );
  OAI22_X1 U312 ( .A1(n324), .A2(n323), .B1(n325), .B2(n321), .ZN(n98) );
  XNOR2_X1 U313 ( .A(b[6]), .B(a[1]), .ZN(n324) );
  OAI22_X1 U314 ( .A1(n321), .A2(n325), .B1(n323), .B2(n325), .ZN(n326) );
  XNOR2_X1 U315 ( .A(b[7]), .B(a[1]), .ZN(n325) );
  OAI22_X1 U316 ( .A1(n328), .A2(n329), .B1(n292), .B2(n330), .ZN(n95) );
  XNOR2_X1 U317 ( .A(a[3]), .B(n308), .ZN(n328) );
  OAI22_X1 U318 ( .A1(n330), .A2(n329), .B1(n331), .B2(n292), .ZN(n94) );
  OAI22_X1 U319 ( .A1(n331), .A2(n329), .B1(n292), .B2(n332), .ZN(n93) );
  XNOR2_X1 U320 ( .A(b[2]), .B(a[3]), .ZN(n331) );
  OAI22_X1 U321 ( .A1(n332), .A2(n329), .B1(n291), .B2(n333), .ZN(n92) );
  XNOR2_X1 U322 ( .A(b[3]), .B(a[3]), .ZN(n332) );
  OAI22_X1 U323 ( .A1(n333), .A2(n329), .B1(n292), .B2(n334), .ZN(n91) );
  XNOR2_X1 U324 ( .A(b[4]), .B(a[3]), .ZN(n333) );
  OAI22_X1 U325 ( .A1(n336), .A2(n291), .B1(n329), .B2(n336), .ZN(n335) );
  NOR2_X1 U326 ( .A1(n337), .A2(n309), .ZN(n88) );
  OAI22_X1 U327 ( .A1(n338), .A2(n339), .B1(n337), .B2(n340), .ZN(n87) );
  XNOR2_X1 U328 ( .A(a[5]), .B(n271), .ZN(n338) );
  OAI22_X1 U329 ( .A1(n340), .A2(n339), .B1(n337), .B2(n341), .ZN(n86) );
  XNOR2_X1 U330 ( .A(n277), .B(a[5]), .ZN(n340) );
  OAI22_X1 U331 ( .A1(n341), .A2(n339), .B1(n337), .B2(n342), .ZN(n85) );
  XNOR2_X1 U332 ( .A(b[2]), .B(a[5]), .ZN(n341) );
  OAI22_X1 U333 ( .A1(n342), .A2(n339), .B1(n337), .B2(n343), .ZN(n84) );
  XNOR2_X1 U334 ( .A(b[3]), .B(a[5]), .ZN(n342) );
  OAI22_X1 U335 ( .A1(n343), .A2(n339), .B1(n337), .B2(n344), .ZN(n83) );
  XNOR2_X1 U336 ( .A(b[4]), .B(a[5]), .ZN(n343) );
  OAI22_X1 U337 ( .A1(n344), .A2(n339), .B1(n337), .B2(n345), .ZN(n82) );
  XNOR2_X1 U338 ( .A(b[5]), .B(a[5]), .ZN(n344) );
  OAI22_X1 U339 ( .A1(n347), .A2(n337), .B1(n339), .B2(n347), .ZN(n346) );
  NOR2_X1 U340 ( .A1(n348), .A2(n309), .ZN(n80) );
  OAI22_X1 U341 ( .A1(n349), .A2(n350), .B1(n348), .B2(n351), .ZN(n79) );
  XNOR2_X1 U342 ( .A(a[7]), .B(n271), .ZN(n349) );
  OAI22_X1 U343 ( .A1(n352), .A2(n350), .B1(n348), .B2(n353), .ZN(n77) );
  OAI22_X1 U344 ( .A1(n353), .A2(n350), .B1(n348), .B2(n354), .ZN(n76) );
  XNOR2_X1 U345 ( .A(b[3]), .B(a[7]), .ZN(n353) );
  OAI22_X1 U346 ( .A1(n354), .A2(n350), .B1(n348), .B2(n355), .ZN(n75) );
  XNOR2_X1 U347 ( .A(b[4]), .B(a[7]), .ZN(n354) );
  OAI22_X1 U348 ( .A1(n355), .A2(n350), .B1(n348), .B2(n356), .ZN(n74) );
  XNOR2_X1 U349 ( .A(b[5]), .B(a[7]), .ZN(n355) );
  OAI22_X1 U350 ( .A1(n358), .A2(n348), .B1(n350), .B2(n358), .ZN(n357) );
  OAI21_X1 U351 ( .B1(n308), .B2(n320), .A(n323), .ZN(n72) );
  OAI21_X1 U352 ( .B1(n318), .B2(n329), .A(n359), .ZN(n71) );
  OR3_X1 U353 ( .A1(n291), .A2(n271), .A3(n318), .ZN(n359) );
  OAI21_X1 U354 ( .B1(n315), .B2(n339), .A(n360), .ZN(n70) );
  OR3_X1 U355 ( .A1(n337), .A2(n271), .A3(n315), .ZN(n360) );
  OAI21_X1 U356 ( .B1(n312), .B2(n350), .A(n361), .ZN(n69) );
  OR3_X1 U357 ( .A1(n348), .A2(n271), .A3(n312), .ZN(n361) );
  XNOR2_X1 U358 ( .A(n362), .B(n363), .ZN(n38) );
  OR2_X1 U359 ( .A1(n362), .A2(n363), .ZN(n37) );
  OAI22_X1 U360 ( .A1(n334), .A2(n329), .B1(n292), .B2(n364), .ZN(n363) );
  XNOR2_X1 U361 ( .A(b[5]), .B(a[3]), .ZN(n334) );
  OAI22_X1 U362 ( .A1(n351), .A2(n350), .B1(n348), .B2(n352), .ZN(n362) );
  XNOR2_X1 U363 ( .A(b[2]), .B(a[7]), .ZN(n352) );
  XNOR2_X1 U364 ( .A(n277), .B(a[7]), .ZN(n351) );
  OAI22_X1 U365 ( .A1(n364), .A2(n329), .B1(n291), .B2(n336), .ZN(n31) );
  XNOR2_X1 U366 ( .A(b[7]), .B(a[3]), .ZN(n336) );
  XNOR2_X1 U367 ( .A(n318), .B(a[2]), .ZN(n365) );
  XNOR2_X1 U368 ( .A(b[6]), .B(a[3]), .ZN(n364) );
  OAI22_X1 U369 ( .A1(n345), .A2(n339), .B1(n337), .B2(n347), .ZN(n21) );
  XNOR2_X1 U370 ( .A(b[7]), .B(a[5]), .ZN(n347) );
  XNOR2_X1 U371 ( .A(n315), .B(a[4]), .ZN(n366) );
  XNOR2_X1 U372 ( .A(b[6]), .B(a[5]), .ZN(n345) );
  OAI22_X1 U373 ( .A1(n356), .A2(n350), .B1(n348), .B2(n358), .ZN(n15) );
  XNOR2_X1 U374 ( .A(b[7]), .B(a[7]), .ZN(n358) );
  XNOR2_X1 U375 ( .A(n312), .B(a[6]), .ZN(n367) );
  XNOR2_X1 U376 ( .A(b[6]), .B(a[7]), .ZN(n356) );
  OAI22_X1 U377 ( .A1(n308), .A2(n323), .B1(n368), .B2(n321), .ZN(n104) );
  OAI22_X1 U378 ( .A1(n368), .A2(n323), .B1(n369), .B2(n321), .ZN(n103) );
  OAI22_X1 U379 ( .A1(n369), .A2(n323), .B1(n370), .B2(n321), .ZN(n102) );
  XNOR2_X1 U380 ( .A(b[2]), .B(a[1]), .ZN(n369) );
  OAI22_X1 U381 ( .A1(n370), .A2(n323), .B1(n371), .B2(n321), .ZN(n101) );
  OAI22_X1 U382 ( .A1(n371), .A2(n323), .B1(n322), .B2(n321), .ZN(n100) );
  XNOR2_X1 U383 ( .A(b[5]), .B(a[1]), .ZN(n322) );
  NAND2_X1 U384 ( .A1(a[1]), .A2(n321), .ZN(n323) );
  XNOR2_X1 U385 ( .A(b[4]), .B(a[1]), .ZN(n371) );
endmodule


module mac_10 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_10_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_10_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_9_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;
  wire   [15:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .S(SUM[15]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n84) );
  CLKBUF_X1 U2 ( .A(n74), .Z(n1) );
  CLKBUF_X1 U3 ( .A(n61), .Z(n2) );
  NAND3_X1 U4 ( .A1(n23), .A2(n24), .A3(n25), .ZN(n3) );
  CLKBUF_X1 U5 ( .A(n48), .Z(n4) );
  NAND3_X1 U6 ( .A1(n13), .A2(n14), .A3(n15), .ZN(n5) );
  CLKBUF_X1 U7 ( .A(n3), .Z(n6) );
  NAND3_X1 U8 ( .A1(n73), .A2(n74), .A3(n75), .ZN(n7) );
  NAND3_X1 U9 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n8) );
  NAND3_X1 U10 ( .A1(n81), .A2(n82), .A3(n83), .ZN(n9) );
  CLKBUF_X1 U11 ( .A(n5), .Z(n10) );
  CLKBUF_X1 U12 ( .A(n33), .Z(n11) );
  XOR2_X1 U13 ( .A(B[5]), .B(A[5]), .Z(n12) );
  XOR2_X1 U14 ( .A(n6), .B(n12), .Z(SUM[5]) );
  NAND2_X1 U15 ( .A1(n3), .A2(B[5]), .ZN(n13) );
  NAND2_X1 U16 ( .A1(carry[5]), .A2(A[5]), .ZN(n14) );
  NAND2_X1 U17 ( .A1(B[5]), .A2(A[5]), .ZN(n15) );
  NAND3_X1 U18 ( .A1(n13), .A2(n14), .A3(n15), .ZN(carry[6]) );
  NAND3_X1 U19 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n16) );
  CLKBUF_X1 U20 ( .A(n8), .Z(n17) );
  XOR2_X1 U21 ( .A(B[3]), .B(A[3]), .Z(n18) );
  XOR2_X1 U22 ( .A(carry[3]), .B(n18), .Z(SUM[3]) );
  NAND2_X1 U23 ( .A1(n9), .A2(B[3]), .ZN(n19) );
  NAND2_X1 U24 ( .A1(n9), .A2(A[3]), .ZN(n20) );
  NAND2_X1 U25 ( .A1(B[3]), .A2(A[3]), .ZN(n21) );
  NAND3_X1 U26 ( .A1(n20), .A2(n19), .A3(n21), .ZN(carry[4]) );
  XOR2_X1 U27 ( .A(B[4]), .B(A[4]), .Z(n22) );
  XOR2_X1 U28 ( .A(n17), .B(n22), .Z(SUM[4]) );
  NAND2_X1 U29 ( .A1(n8), .A2(B[4]), .ZN(n23) );
  NAND2_X1 U30 ( .A1(carry[4]), .A2(A[4]), .ZN(n24) );
  NAND2_X1 U31 ( .A1(B[4]), .A2(A[4]), .ZN(n25) );
  NAND3_X1 U32 ( .A1(n23), .A2(n24), .A3(n25), .ZN(carry[5]) );
  CLKBUF_X1 U33 ( .A(n34), .Z(n26) );
  XOR2_X1 U34 ( .A(B[6]), .B(A[6]), .Z(n27) );
  XOR2_X1 U35 ( .A(n10), .B(n27), .Z(SUM[6]) );
  NAND2_X1 U36 ( .A1(n5), .A2(B[6]), .ZN(n28) );
  NAND2_X1 U37 ( .A1(carry[6]), .A2(A[6]), .ZN(n29) );
  NAND2_X1 U38 ( .A1(B[6]), .A2(A[6]), .ZN(n30) );
  NAND3_X1 U39 ( .A1(n28), .A2(n29), .A3(n30), .ZN(carry[7]) );
  NAND3_X1 U40 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n31) );
  NAND3_X1 U41 ( .A1(n47), .A2(n4), .A3(n49), .ZN(n32) );
  NAND3_X1 U42 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n33) );
  NAND3_X1 U43 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n34) );
  NAND3_X1 U44 ( .A1(n57), .A2(n58), .A3(n59), .ZN(n35) );
  XOR2_X1 U45 ( .A(B[7]), .B(A[7]), .Z(n36) );
  XOR2_X1 U46 ( .A(carry[7]), .B(n36), .Z(SUM[7]) );
  NAND2_X1 U47 ( .A1(n16), .A2(B[7]), .ZN(n37) );
  NAND2_X1 U48 ( .A1(n16), .A2(A[7]), .ZN(n38) );
  NAND2_X1 U49 ( .A1(B[7]), .A2(A[7]), .ZN(n39) );
  NAND3_X1 U50 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[8]) );
  XOR2_X1 U51 ( .A(B[13]), .B(A[13]), .Z(n40) );
  XOR2_X1 U52 ( .A(n32), .B(n40), .Z(SUM[13]) );
  NAND2_X1 U53 ( .A1(n31), .A2(B[13]), .ZN(n41) );
  NAND2_X1 U54 ( .A1(carry[13]), .A2(A[13]), .ZN(n42) );
  NAND2_X1 U55 ( .A1(B[13]), .A2(A[13]), .ZN(n43) );
  NAND3_X1 U56 ( .A1(n42), .A2(n41), .A3(n43), .ZN(carry[14]) );
  NAND3_X1 U57 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n44) );
  NAND3_X1 U58 ( .A1(n2), .A2(n62), .A3(n63), .ZN(n45) );
  XOR2_X1 U59 ( .A(B[12]), .B(A[12]), .Z(n46) );
  XOR2_X1 U60 ( .A(n45), .B(n46), .Z(SUM[12]) );
  NAND2_X1 U61 ( .A1(n44), .A2(B[12]), .ZN(n47) );
  NAND2_X1 U62 ( .A1(carry[12]), .A2(A[12]), .ZN(n48) );
  NAND2_X1 U63 ( .A1(B[12]), .A2(A[12]), .ZN(n49) );
  NAND3_X1 U64 ( .A1(n47), .A2(n48), .A3(n49), .ZN(carry[13]) );
  XOR2_X1 U65 ( .A(B[14]), .B(A[14]), .Z(n50) );
  XOR2_X1 U66 ( .A(n11), .B(n50), .Z(SUM[14]) );
  NAND2_X1 U67 ( .A1(n33), .A2(B[14]), .ZN(n51) );
  NAND2_X1 U68 ( .A1(carry[14]), .A2(A[14]), .ZN(n52) );
  NAND2_X1 U69 ( .A1(B[14]), .A2(A[14]), .ZN(n53) );
  NAND3_X1 U70 ( .A1(n51), .A2(n52), .A3(n53), .ZN(carry[15]) );
  CLKBUF_X1 U71 ( .A(n35), .Z(n54) );
  NAND3_X1 U72 ( .A1(n73), .A2(n1), .A3(n75), .ZN(n55) );
  XOR2_X1 U73 ( .A(B[10]), .B(A[10]), .Z(n56) );
  XOR2_X1 U74 ( .A(n55), .B(n56), .Z(SUM[10]) );
  NAND2_X1 U75 ( .A1(n7), .A2(B[10]), .ZN(n57) );
  NAND2_X1 U76 ( .A1(carry[10]), .A2(A[10]), .ZN(n58) );
  NAND2_X1 U77 ( .A1(B[10]), .A2(A[10]), .ZN(n59) );
  NAND3_X1 U78 ( .A1(n58), .A2(n57), .A3(n59), .ZN(carry[11]) );
  XOR2_X1 U79 ( .A(B[11]), .B(A[11]), .Z(n60) );
  XOR2_X1 U80 ( .A(n54), .B(n60), .Z(SUM[11]) );
  NAND2_X1 U81 ( .A1(n35), .A2(B[11]), .ZN(n61) );
  NAND2_X1 U82 ( .A1(carry[11]), .A2(A[11]), .ZN(n62) );
  NAND2_X1 U83 ( .A1(B[11]), .A2(A[11]), .ZN(n63) );
  NAND3_X1 U84 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[12]) );
  NAND3_X1 U85 ( .A1(n77), .A2(n78), .A3(n79), .ZN(n64) );
  NAND3_X1 U86 ( .A1(n77), .A2(n78), .A3(n79), .ZN(n65) );
  NAND3_X1 U87 ( .A1(n69), .A2(n70), .A3(n71), .ZN(n66) );
  NAND3_X1 U88 ( .A1(n69), .A2(n70), .A3(n71), .ZN(n67) );
  XOR2_X1 U89 ( .A(B[8]), .B(A[8]), .Z(n68) );
  XOR2_X1 U90 ( .A(n26), .B(n68), .Z(SUM[8]) );
  NAND2_X1 U91 ( .A1(n34), .A2(B[8]), .ZN(n69) );
  NAND2_X1 U92 ( .A1(carry[8]), .A2(A[8]), .ZN(n70) );
  NAND2_X1 U93 ( .A1(B[8]), .A2(A[8]), .ZN(n71) );
  NAND3_X1 U94 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[9]) );
  XOR2_X1 U95 ( .A(B[9]), .B(A[9]), .Z(n72) );
  XOR2_X1 U96 ( .A(n67), .B(n72), .Z(SUM[9]) );
  NAND2_X1 U97 ( .A1(n66), .A2(B[9]), .ZN(n73) );
  NAND2_X1 U98 ( .A1(carry[9]), .A2(A[9]), .ZN(n74) );
  NAND2_X1 U99 ( .A1(B[9]), .A2(A[9]), .ZN(n75) );
  NAND3_X1 U100 ( .A1(n73), .A2(n74), .A3(n75), .ZN(carry[10]) );
  XOR2_X1 U101 ( .A(B[1]), .B(A[1]), .Z(n76) );
  XOR2_X1 U102 ( .A(n84), .B(n76), .Z(SUM[1]) );
  NAND2_X1 U103 ( .A1(n84), .A2(B[1]), .ZN(n77) );
  NAND2_X1 U104 ( .A1(n84), .A2(A[1]), .ZN(n78) );
  NAND2_X1 U105 ( .A1(B[1]), .A2(A[1]), .ZN(n79) );
  NAND3_X1 U106 ( .A1(n77), .A2(n78), .A3(n79), .ZN(carry[2]) );
  XOR2_X1 U107 ( .A(B[2]), .B(A[2]), .Z(n80) );
  XOR2_X1 U108 ( .A(n65), .B(n80), .Z(SUM[2]) );
  NAND2_X1 U109 ( .A1(n64), .A2(B[2]), .ZN(n81) );
  NAND2_X1 U110 ( .A1(carry[2]), .A2(A[2]), .ZN(n82) );
  NAND2_X1 U111 ( .A1(B[2]), .A2(A[2]), .ZN(n83) );
  NAND3_X1 U112 ( .A1(n81), .A2(n82), .A3(n83), .ZN(carry[3]) );
  XOR2_X1 U113 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_9_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378;

  HA_X1 U15 ( .A(n208), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n321), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n320), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n324), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n323), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n326), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  NAND2_X1 U157 ( .A1(n334), .A2(n372), .ZN(n336) );
  INV_X1 U158 ( .A(n316), .ZN(n267) );
  NAND2_X1 U159 ( .A1(n50), .A2(n53), .ZN(n312) );
  INV_X1 U160 ( .A(n15), .ZN(n317) );
  CLKBUF_X1 U161 ( .A(n244), .Z(n206) );
  CLKBUF_X1 U162 ( .A(n314), .Z(n207) );
  OAI22_X1 U163 ( .A1(n267), .A2(n330), .B1(n375), .B2(n328), .ZN(n208) );
  AND2_X1 U164 ( .A1(n95), .A2(n102), .ZN(n209) );
  XNOR2_X1 U165 ( .A(n318), .B(n15), .ZN(n210) );
  XOR2_X1 U166 ( .A(n100), .B(n93), .Z(n211) );
  XOR2_X1 U167 ( .A(n52), .B(n211), .Z(n50) );
  NAND2_X1 U168 ( .A1(n52), .A2(n100), .ZN(n212) );
  NAND2_X1 U169 ( .A1(n52), .A2(n93), .ZN(n213) );
  NAND2_X1 U170 ( .A1(n100), .A2(n93), .ZN(n214) );
  NAND3_X1 U171 ( .A1(n212), .A2(n213), .A3(n214), .ZN(n49) );
  NAND3_X1 U172 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n215) );
  CLKBUF_X1 U173 ( .A(n8), .Z(n216) );
  XNOR2_X1 U174 ( .A(b[3]), .B(a[1]), .ZN(n217) );
  CLKBUF_X1 U175 ( .A(b[1]), .Z(n218) );
  AND2_X1 U176 ( .A1(n208), .A2(n72), .ZN(n219) );
  NAND3_X1 U177 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n220) );
  NAND3_X1 U178 ( .A1(n243), .A2(n206), .A3(n245), .ZN(n221) );
  NAND3_X1 U179 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n222) );
  NAND3_X1 U180 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n223) );
  NAND2_X1 U181 ( .A1(n219), .A2(n96), .ZN(n224) );
  NAND2_X1 U182 ( .A1(n219), .A2(n96), .ZN(n225) );
  INV_X1 U183 ( .A(n316), .ZN(n315) );
  CLKBUF_X1 U184 ( .A(n298), .Z(n226) );
  NAND3_X1 U185 ( .A1(n290), .A2(n289), .A3(n288), .ZN(n227) );
  NAND3_X1 U186 ( .A1(n302), .A2(n301), .A3(n303), .ZN(n228) );
  XOR2_X1 U187 ( .A(n95), .B(n102), .Z(n56) );
  XNOR2_X1 U188 ( .A(a[2]), .B(a[1]), .ZN(n334) );
  AND2_X1 U189 ( .A1(n104), .A2(n72), .ZN(n229) );
  NAND2_X1 U190 ( .A1(n269), .A2(n20), .ZN(n230) );
  CLKBUF_X1 U191 ( .A(n56), .Z(n231) );
  NAND2_X2 U192 ( .A1(n355), .A2(n374), .ZN(n357) );
  XOR2_X2 U193 ( .A(a[6]), .B(n322), .Z(n355) );
  CLKBUF_X1 U194 ( .A(n313), .Z(n232) );
  CLKBUF_X1 U195 ( .A(n310), .Z(n233) );
  BUF_X2 U196 ( .A(n344), .Z(n234) );
  XNOR2_X1 U197 ( .A(a[4]), .B(a[3]), .ZN(n344) );
  XNOR2_X1 U198 ( .A(n223), .B(n210), .ZN(product[14]) );
  AND3_X1 U199 ( .A1(n249), .A2(n248), .A3(n250), .ZN(product[15]) );
  CLKBUF_X1 U200 ( .A(n230), .Z(n236) );
  CLKBUF_X1 U201 ( .A(n261), .Z(n237) );
  XOR2_X1 U202 ( .A(n17), .B(n317), .Z(n238) );
  XOR2_X1 U203 ( .A(n3), .B(n238), .Z(product[13]) );
  NAND2_X1 U204 ( .A1(n227), .A2(n17), .ZN(n239) );
  NAND2_X1 U205 ( .A1(n227), .A2(n317), .ZN(n240) );
  NAND2_X1 U206 ( .A1(n17), .A2(n317), .ZN(n241) );
  NAND3_X1 U207 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n2) );
  XOR2_X1 U208 ( .A(n34), .B(n39), .Z(n242) );
  XOR2_X1 U209 ( .A(n216), .B(n242), .Z(product[8]) );
  NAND2_X1 U210 ( .A1(n228), .A2(n34), .ZN(n243) );
  NAND2_X1 U211 ( .A1(n8), .A2(n39), .ZN(n244) );
  NAND2_X1 U212 ( .A1(n34), .A2(n39), .ZN(n245) );
  NAND3_X1 U213 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n7) );
  NAND3_X1 U214 ( .A1(n254), .A2(n224), .A3(n256), .ZN(n246) );
  NAND3_X1 U215 ( .A1(n254), .A2(n225), .A3(n256), .ZN(n247) );
  NAND2_X1 U216 ( .A1(n2), .A2(n318), .ZN(n248) );
  NAND2_X1 U217 ( .A1(n222), .A2(n15), .ZN(n249) );
  NAND2_X1 U218 ( .A1(n318), .A2(n15), .ZN(n250) );
  CLKBUF_X1 U219 ( .A(n286), .Z(n251) );
  CLKBUF_X1 U220 ( .A(n280), .Z(n252) );
  XOR2_X1 U221 ( .A(n103), .B(n96), .Z(n253) );
  XOR2_X1 U222 ( .A(n229), .B(n253), .Z(product[2]) );
  NAND2_X1 U223 ( .A1(n229), .A2(n103), .ZN(n254) );
  NAND2_X1 U224 ( .A1(n14), .A2(n96), .ZN(n255) );
  NAND2_X1 U225 ( .A1(n103), .A2(n96), .ZN(n256) );
  NAND3_X1 U226 ( .A1(n255), .A2(n254), .A3(n256), .ZN(n13) );
  NAND3_X1 U227 ( .A1(n260), .A2(n237), .A3(n262), .ZN(n257) );
  CLKBUF_X1 U228 ( .A(n273), .Z(n258) );
  XOR2_X1 U229 ( .A(n33), .B(n28), .Z(n259) );
  XOR2_X1 U230 ( .A(n221), .B(n259), .Z(product[9]) );
  NAND2_X1 U231 ( .A1(n7), .A2(n33), .ZN(n260) );
  NAND2_X1 U232 ( .A1(n220), .A2(n28), .ZN(n261) );
  NAND2_X1 U233 ( .A1(n33), .A2(n28), .ZN(n262) );
  NAND3_X1 U234 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n6) );
  NAND3_X1 U235 ( .A1(n312), .A2(n313), .A3(n314), .ZN(n263) );
  NAND3_X1 U236 ( .A1(n312), .A2(n232), .A3(n207), .ZN(n264) );
  NAND3_X1 U237 ( .A1(n297), .A2(n298), .A3(n299), .ZN(n265) );
  NAND3_X1 U238 ( .A1(n297), .A2(n226), .A3(n299), .ZN(n266) );
  INV_X1 U239 ( .A(n267), .ZN(n268) );
  NAND3_X1 U240 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n269) );
  NAND3_X1 U241 ( .A1(n272), .A2(n258), .A3(n274), .ZN(n270) );
  XOR2_X1 U242 ( .A(n27), .B(n24), .Z(n271) );
  XOR2_X1 U243 ( .A(n257), .B(n271), .Z(product[10]) );
  NAND2_X1 U244 ( .A1(n215), .A2(n27), .ZN(n272) );
  NAND2_X1 U245 ( .A1(n6), .A2(n24), .ZN(n273) );
  NAND2_X1 U246 ( .A1(n27), .A2(n24), .ZN(n274) );
  NAND3_X1 U247 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n5) );
  NAND3_X1 U248 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n275) );
  NAND3_X1 U249 ( .A1(n278), .A2(n279), .A3(n252), .ZN(n276) );
  XOR2_X1 U250 ( .A(n247), .B(n71), .Z(n277) );
  XOR2_X1 U251 ( .A(n231), .B(n277), .Z(product[3]) );
  NAND2_X1 U252 ( .A1(n246), .A2(n56), .ZN(n278) );
  NAND2_X1 U253 ( .A1(n56), .A2(n71), .ZN(n279) );
  NAND2_X1 U254 ( .A1(n13), .A2(n71), .ZN(n280) );
  NAND3_X1 U255 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n12) );
  NAND3_X1 U256 ( .A1(n286), .A2(n285), .A3(n284), .ZN(n281) );
  NAND3_X1 U257 ( .A1(n284), .A2(n236), .A3(n251), .ZN(n282) );
  XOR2_X1 U258 ( .A(n20), .B(n23), .Z(n283) );
  XOR2_X1 U259 ( .A(n283), .B(n270), .Z(product[11]) );
  NAND2_X1 U260 ( .A1(n20), .A2(n23), .ZN(n284) );
  NAND2_X1 U261 ( .A1(n269), .A2(n20), .ZN(n285) );
  NAND2_X1 U262 ( .A1(n5), .A2(n23), .ZN(n286) );
  NAND3_X1 U263 ( .A1(n230), .A2(n286), .A3(n284), .ZN(n4) );
  XOR2_X1 U264 ( .A(n19), .B(n18), .Z(n287) );
  XOR2_X1 U265 ( .A(n287), .B(n282), .Z(product[12]) );
  NAND2_X1 U266 ( .A1(n19), .A2(n18), .ZN(n288) );
  NAND2_X1 U267 ( .A1(n281), .A2(n19), .ZN(n289) );
  NAND2_X1 U268 ( .A1(n4), .A2(n18), .ZN(n290) );
  NAND3_X1 U269 ( .A1(n288), .A2(n289), .A3(n290), .ZN(n3) );
  NAND3_X1 U270 ( .A1(n309), .A2(n308), .A3(n310), .ZN(n291) );
  NAND3_X1 U271 ( .A1(n308), .A2(n309), .A3(n233), .ZN(n292) );
  NAND2_X2 U272 ( .A1(n344), .A2(n373), .ZN(n346) );
  NAND2_X1 U273 ( .A1(n334), .A2(n372), .ZN(n293) );
  XOR2_X1 U274 ( .A(a[2]), .B(n327), .Z(n294) );
  XOR2_X1 U275 ( .A(a[2]), .B(n327), .Z(n295) );
  INV_X1 U276 ( .A(n342), .ZN(n324) );
  INV_X1 U277 ( .A(n21), .ZN(n320) );
  INV_X1 U278 ( .A(n353), .ZN(n321) );
  INV_X1 U279 ( .A(n333), .ZN(n326) );
  INV_X1 U280 ( .A(b[0]), .ZN(n316) );
  INV_X1 U281 ( .A(n364), .ZN(n318) );
  INV_X1 U282 ( .A(n31), .ZN(n323) );
  INV_X1 U283 ( .A(a[0]), .ZN(n328) );
  INV_X1 U284 ( .A(a[5]), .ZN(n322) );
  INV_X1 U285 ( .A(a[7]), .ZN(n319) );
  XOR2_X1 U286 ( .A(n46), .B(n49), .Z(n296) );
  XOR2_X1 U287 ( .A(n264), .B(n296), .Z(product[6]) );
  NAND2_X1 U288 ( .A1(n263), .A2(n46), .ZN(n297) );
  NAND2_X1 U289 ( .A1(n10), .A2(n49), .ZN(n298) );
  NAND2_X1 U290 ( .A1(n46), .A2(n49), .ZN(n299) );
  NAND3_X1 U291 ( .A1(n297), .A2(n298), .A3(n299), .ZN(n9) );
  XOR2_X1 U292 ( .A(n40), .B(n45), .Z(n300) );
  XOR2_X1 U293 ( .A(n266), .B(n300), .Z(product[7]) );
  NAND2_X1 U294 ( .A1(n265), .A2(n40), .ZN(n301) );
  NAND2_X1 U295 ( .A1(n9), .A2(n45), .ZN(n302) );
  NAND2_X1 U296 ( .A1(n40), .A2(n45), .ZN(n303) );
  NAND3_X1 U297 ( .A1(n301), .A2(n302), .A3(n303), .ZN(n8) );
  NAND2_X1 U298 ( .A1(b[1]), .A2(a[1]), .ZN(n305) );
  NAND2_X1 U299 ( .A1(n304), .A2(n327), .ZN(n306) );
  NAND2_X1 U300 ( .A1(n305), .A2(n306), .ZN(n375) );
  INV_X1 U301 ( .A(b[1]), .ZN(n304) );
  INV_X1 U302 ( .A(a[3]), .ZN(n325) );
  XOR2_X1 U303 ( .A(n54), .B(n209), .Z(n307) );
  XOR2_X1 U304 ( .A(n307), .B(n276), .Z(product[4]) );
  NAND2_X1 U305 ( .A1(n54), .A2(n209), .ZN(n308) );
  NAND2_X1 U306 ( .A1(n275), .A2(n54), .ZN(n309) );
  NAND2_X1 U307 ( .A1(n12), .A2(n209), .ZN(n310) );
  NAND3_X1 U308 ( .A1(n310), .A2(n309), .A3(n308), .ZN(n11) );
  XOR2_X1 U309 ( .A(n50), .B(n53), .Z(n311) );
  XOR2_X1 U310 ( .A(n311), .B(n292), .Z(product[5]) );
  NAND2_X1 U311 ( .A1(n50), .A2(n291), .ZN(n313) );
  NAND2_X1 U312 ( .A1(n11), .A2(n53), .ZN(n314) );
  NAND3_X1 U313 ( .A1(n312), .A2(n313), .A3(n314), .ZN(n10) );
  INV_X1 U314 ( .A(a[1]), .ZN(n327) );
  NOR2_X1 U315 ( .A1(n328), .A2(n268), .ZN(product[0]) );
  OAI22_X1 U316 ( .A1(n329), .A2(n330), .B1(n331), .B2(n328), .ZN(n99) );
  OAI22_X1 U317 ( .A1(n331), .A2(n330), .B1(n332), .B2(n328), .ZN(n98) );
  XNOR2_X1 U318 ( .A(b[6]), .B(a[1]), .ZN(n331) );
  OAI22_X1 U319 ( .A1(n328), .A2(n332), .B1(n330), .B2(n332), .ZN(n333) );
  XNOR2_X1 U320 ( .A(b[7]), .B(a[1]), .ZN(n332) );
  NOR2_X1 U321 ( .A1(n295), .A2(n268), .ZN(n96) );
  OAI22_X1 U322 ( .A1(n335), .A2(n336), .B1(n294), .B2(n337), .ZN(n95) );
  XNOR2_X1 U323 ( .A(a[3]), .B(n315), .ZN(n335) );
  OAI22_X1 U324 ( .A1(n337), .A2(n293), .B1(n294), .B2(n338), .ZN(n94) );
  XNOR2_X1 U325 ( .A(b[1]), .B(a[3]), .ZN(n337) );
  OAI22_X1 U326 ( .A1(n338), .A2(n336), .B1(n294), .B2(n339), .ZN(n93) );
  XNOR2_X1 U327 ( .A(b[2]), .B(a[3]), .ZN(n338) );
  OAI22_X1 U328 ( .A1(n339), .A2(n293), .B1(n295), .B2(n340), .ZN(n92) );
  XNOR2_X1 U329 ( .A(b[3]), .B(a[3]), .ZN(n339) );
  OAI22_X1 U330 ( .A1(n340), .A2(n293), .B1(n295), .B2(n341), .ZN(n91) );
  XNOR2_X1 U331 ( .A(b[4]), .B(a[3]), .ZN(n340) );
  OAI22_X1 U332 ( .A1(n343), .A2(n294), .B1(n336), .B2(n343), .ZN(n342) );
  NOR2_X1 U333 ( .A1(n234), .A2(n268), .ZN(n88) );
  OAI22_X1 U334 ( .A1(n345), .A2(n346), .B1(n234), .B2(n347), .ZN(n87) );
  XNOR2_X1 U335 ( .A(a[5]), .B(n267), .ZN(n345) );
  OAI22_X1 U336 ( .A1(n347), .A2(n346), .B1(n234), .B2(n348), .ZN(n86) );
  XNOR2_X1 U337 ( .A(n218), .B(a[5]), .ZN(n347) );
  OAI22_X1 U338 ( .A1(n348), .A2(n346), .B1(n234), .B2(n349), .ZN(n85) );
  XNOR2_X1 U339 ( .A(b[2]), .B(a[5]), .ZN(n348) );
  OAI22_X1 U340 ( .A1(n349), .A2(n346), .B1(n234), .B2(n350), .ZN(n84) );
  XNOR2_X1 U341 ( .A(b[3]), .B(a[5]), .ZN(n349) );
  OAI22_X1 U342 ( .A1(n350), .A2(n346), .B1(n234), .B2(n351), .ZN(n83) );
  XNOR2_X1 U343 ( .A(b[4]), .B(a[5]), .ZN(n350) );
  OAI22_X1 U344 ( .A1(n351), .A2(n346), .B1(n234), .B2(n352), .ZN(n82) );
  XNOR2_X1 U345 ( .A(b[5]), .B(a[5]), .ZN(n351) );
  OAI22_X1 U346 ( .A1(n354), .A2(n234), .B1(n346), .B2(n354), .ZN(n353) );
  NOR2_X1 U347 ( .A1(n355), .A2(n268), .ZN(n80) );
  OAI22_X1 U348 ( .A1(n356), .A2(n357), .B1(n355), .B2(n358), .ZN(n79) );
  XNOR2_X1 U349 ( .A(a[7]), .B(n267), .ZN(n356) );
  OAI22_X1 U350 ( .A1(n359), .A2(n357), .B1(n355), .B2(n360), .ZN(n77) );
  OAI22_X1 U351 ( .A1(n360), .A2(n357), .B1(n355), .B2(n361), .ZN(n76) );
  XNOR2_X1 U352 ( .A(b[3]), .B(a[7]), .ZN(n360) );
  OAI22_X1 U353 ( .A1(n361), .A2(n357), .B1(n355), .B2(n362), .ZN(n75) );
  XNOR2_X1 U354 ( .A(b[4]), .B(a[7]), .ZN(n361) );
  OAI22_X1 U355 ( .A1(n362), .A2(n357), .B1(n355), .B2(n363), .ZN(n74) );
  XNOR2_X1 U356 ( .A(b[5]), .B(a[7]), .ZN(n362) );
  OAI22_X1 U357 ( .A1(n365), .A2(n355), .B1(n357), .B2(n365), .ZN(n364) );
  OAI21_X1 U358 ( .B1(n315), .B2(n327), .A(n330), .ZN(n72) );
  OAI21_X1 U359 ( .B1(n325), .B2(n336), .A(n366), .ZN(n71) );
  OR3_X1 U360 ( .A1(n295), .A2(n267), .A3(n325), .ZN(n366) );
  OAI21_X1 U361 ( .B1(n322), .B2(n346), .A(n367), .ZN(n70) );
  OR3_X1 U362 ( .A1(n234), .A2(n315), .A3(n322), .ZN(n367) );
  OAI21_X1 U363 ( .B1(n319), .B2(n357), .A(n368), .ZN(n69) );
  OR3_X1 U364 ( .A1(n355), .A2(n267), .A3(n319), .ZN(n368) );
  XNOR2_X1 U365 ( .A(n369), .B(n370), .ZN(n38) );
  OR2_X1 U366 ( .A1(n369), .A2(n370), .ZN(n37) );
  OAI22_X1 U367 ( .A1(n341), .A2(n336), .B1(n294), .B2(n371), .ZN(n370) );
  XNOR2_X1 U368 ( .A(b[5]), .B(a[3]), .ZN(n341) );
  OAI22_X1 U369 ( .A1(n358), .A2(n357), .B1(n355), .B2(n359), .ZN(n369) );
  XNOR2_X1 U370 ( .A(b[2]), .B(a[7]), .ZN(n359) );
  XNOR2_X1 U371 ( .A(n218), .B(a[7]), .ZN(n358) );
  OAI22_X1 U372 ( .A1(n371), .A2(n293), .B1(n295), .B2(n343), .ZN(n31) );
  XNOR2_X1 U373 ( .A(b[7]), .B(a[3]), .ZN(n343) );
  XNOR2_X1 U374 ( .A(n325), .B(a[2]), .ZN(n372) );
  XNOR2_X1 U375 ( .A(b[6]), .B(a[3]), .ZN(n371) );
  OAI22_X1 U376 ( .A1(n352), .A2(n346), .B1(n234), .B2(n354), .ZN(n21) );
  XNOR2_X1 U377 ( .A(b[7]), .B(a[5]), .ZN(n354) );
  XNOR2_X1 U378 ( .A(n322), .B(a[4]), .ZN(n373) );
  XNOR2_X1 U379 ( .A(b[6]), .B(a[5]), .ZN(n352) );
  OAI22_X1 U380 ( .A1(n363), .A2(n357), .B1(n355), .B2(n365), .ZN(n15) );
  XNOR2_X1 U381 ( .A(b[7]), .B(a[7]), .ZN(n365) );
  XNOR2_X1 U382 ( .A(n319), .B(a[6]), .ZN(n374) );
  XNOR2_X1 U383 ( .A(b[6]), .B(a[7]), .ZN(n363) );
  OAI22_X1 U384 ( .A1(n267), .A2(n330), .B1(n375), .B2(n328), .ZN(n104) );
  OAI22_X1 U385 ( .A1(n375), .A2(n330), .B1(n376), .B2(n328), .ZN(n103) );
  OAI22_X1 U386 ( .A1(n376), .A2(n330), .B1(n377), .B2(n328), .ZN(n102) );
  XNOR2_X1 U387 ( .A(b[2]), .B(a[1]), .ZN(n376) );
  OAI22_X1 U388 ( .A1(n217), .A2(n330), .B1(n378), .B2(n328), .ZN(n101) );
  XNOR2_X1 U389 ( .A(b[3]), .B(a[1]), .ZN(n377) );
  OAI22_X1 U390 ( .A1(n378), .A2(n330), .B1(n329), .B2(n328), .ZN(n100) );
  XNOR2_X1 U391 ( .A(b[5]), .B(a[1]), .ZN(n329) );
  NAND2_X1 U392 ( .A1(a[1]), .A2(n328), .ZN(n330) );
  XNOR2_X1 U393 ( .A(b[4]), .B(a[1]), .ZN(n378) );
endmodule


module mac_9 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_9_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_9_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_8_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79;
  wire   [15:1] carry;

  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n79) );
  XOR2_X1 U2 ( .A(B[15]), .B(A[15]), .Z(n1) );
  XOR2_X1 U3 ( .A(carry[15]), .B(n1), .Z(SUM[15]) );
  NAND3_X1 U4 ( .A1(n9), .A2(n10), .A3(n11), .ZN(n2) );
  NAND3_X1 U5 ( .A1(n9), .A2(n10), .A3(n11), .ZN(n3) );
  NAND3_X1 U6 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n4) );
  NAND3_X1 U7 ( .A1(n68), .A2(n69), .A3(n70), .ZN(n5) );
  NAND3_X1 U8 ( .A1(n26), .A2(n25), .A3(n27), .ZN(n6) );
  NAND3_X1 U9 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n7) );
  XOR2_X1 U10 ( .A(B[3]), .B(A[3]), .Z(n8) );
  XOR2_X1 U11 ( .A(carry[3]), .B(n8), .Z(SUM[3]) );
  NAND2_X1 U12 ( .A1(carry[3]), .A2(B[3]), .ZN(n9) );
  NAND2_X1 U13 ( .A1(carry[3]), .A2(A[3]), .ZN(n10) );
  NAND2_X1 U14 ( .A1(B[3]), .A2(A[3]), .ZN(n11) );
  NAND3_X1 U15 ( .A1(n9), .A2(n10), .A3(n11), .ZN(carry[4]) );
  NAND3_X1 U16 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n12) );
  NAND3_X1 U17 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n13) );
  NAND3_X1 U18 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n14) );
  NAND3_X1 U19 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n15) );
  NAND3_X1 U20 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n16) );
  NAND3_X1 U21 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n17) );
  NAND3_X1 U22 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n18) );
  NAND3_X1 U23 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n19) );
  XOR2_X1 U24 ( .A(B[4]), .B(A[4]), .Z(n20) );
  XOR2_X1 U25 ( .A(n3), .B(n20), .Z(SUM[4]) );
  NAND2_X1 U26 ( .A1(n2), .A2(B[4]), .ZN(n21) );
  NAND2_X1 U27 ( .A1(carry[4]), .A2(A[4]), .ZN(n22) );
  NAND2_X1 U28 ( .A1(B[4]), .A2(A[4]), .ZN(n23) );
  NAND3_X1 U29 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[5]) );
  XOR2_X1 U30 ( .A(B[11]), .B(A[11]), .Z(n24) );
  XOR2_X1 U31 ( .A(n16), .B(n24), .Z(SUM[11]) );
  NAND2_X1 U32 ( .A1(n15), .A2(B[11]), .ZN(n25) );
  NAND2_X1 U33 ( .A1(carry[11]), .A2(A[11]), .ZN(n26) );
  NAND2_X1 U34 ( .A1(B[11]), .A2(A[11]), .ZN(n27) );
  NAND3_X1 U35 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[12]) );
  XOR2_X1 U36 ( .A(B[6]), .B(A[6]), .Z(n28) );
  XOR2_X1 U37 ( .A(n4), .B(n28), .Z(SUM[6]) );
  NAND2_X1 U38 ( .A1(carry[6]), .A2(B[6]), .ZN(n29) );
  NAND2_X1 U39 ( .A1(n19), .A2(A[6]), .ZN(n30) );
  NAND2_X1 U40 ( .A1(B[6]), .A2(A[6]), .ZN(n31) );
  NAND3_X1 U41 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[7]) );
  XOR2_X1 U42 ( .A(B[5]), .B(A[5]), .Z(n32) );
  XOR2_X1 U43 ( .A(n18), .B(n32), .Z(SUM[5]) );
  NAND2_X1 U44 ( .A1(n17), .A2(B[5]), .ZN(n33) );
  NAND2_X1 U45 ( .A1(carry[5]), .A2(A[5]), .ZN(n34) );
  NAND2_X1 U46 ( .A1(B[5]), .A2(A[5]), .ZN(n35) );
  NAND3_X1 U47 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[6]) );
  XOR2_X1 U48 ( .A(B[12]), .B(A[12]), .Z(n36) );
  XOR2_X1 U49 ( .A(n6), .B(n36), .Z(SUM[12]) );
  NAND2_X1 U50 ( .A1(n6), .A2(B[12]), .ZN(n37) );
  NAND2_X1 U51 ( .A1(carry[12]), .A2(A[12]), .ZN(n38) );
  NAND2_X1 U52 ( .A1(B[12]), .A2(A[12]), .ZN(n39) );
  NAND3_X1 U53 ( .A1(n38), .A2(n37), .A3(n39), .ZN(carry[13]) );
  NAND3_X1 U54 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n40) );
  NAND3_X1 U55 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n41) );
  NAND3_X1 U56 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n42) );
  NAND3_X1 U57 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n43) );
  NAND3_X1 U58 ( .A1(n68), .A2(n69), .A3(n70), .ZN(n44) );
  XOR2_X1 U59 ( .A(B[10]), .B(A[10]), .Z(n45) );
  XOR2_X1 U60 ( .A(n5), .B(n45), .Z(SUM[10]) );
  NAND2_X1 U61 ( .A1(carry[10]), .A2(B[10]), .ZN(n46) );
  NAND2_X1 U62 ( .A1(n44), .A2(A[10]), .ZN(n47) );
  NAND2_X1 U63 ( .A1(B[10]), .A2(A[10]), .ZN(n48) );
  NAND3_X1 U64 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[11]) );
  XOR2_X1 U65 ( .A(B[13]), .B(A[13]), .Z(n49) );
  XOR2_X1 U66 ( .A(n12), .B(n49), .Z(SUM[13]) );
  NAND2_X1 U67 ( .A1(n12), .A2(B[13]), .ZN(n50) );
  NAND2_X1 U68 ( .A1(carry[13]), .A2(A[13]), .ZN(n51) );
  NAND2_X1 U69 ( .A1(B[13]), .A2(A[13]), .ZN(n52) );
  XOR2_X1 U70 ( .A(B[7]), .B(A[7]), .Z(n53) );
  XOR2_X1 U71 ( .A(n14), .B(n53), .Z(SUM[7]) );
  NAND2_X1 U72 ( .A1(n13), .A2(B[7]), .ZN(n54) );
  NAND2_X1 U73 ( .A1(carry[7]), .A2(A[7]), .ZN(n55) );
  NAND2_X1 U74 ( .A1(B[7]), .A2(A[7]), .ZN(n56) );
  NAND3_X1 U75 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[8]) );
  NAND3_X1 U76 ( .A1(n72), .A2(n73), .A3(n74), .ZN(n57) );
  NAND3_X1 U77 ( .A1(n72), .A2(n73), .A3(n74), .ZN(n58) );
  XOR2_X1 U78 ( .A(B[14]), .B(A[14]), .Z(n59) );
  XOR2_X1 U79 ( .A(n43), .B(n59), .Z(SUM[14]) );
  NAND2_X1 U80 ( .A1(n43), .A2(B[14]), .ZN(n60) );
  NAND2_X1 U81 ( .A1(n42), .A2(A[14]), .ZN(n61) );
  NAND2_X1 U82 ( .A1(B[14]), .A2(A[14]), .ZN(n62) );
  NAND3_X1 U83 ( .A1(n60), .A2(n61), .A3(n62), .ZN(carry[15]) );
  XOR2_X1 U84 ( .A(B[8]), .B(A[8]), .Z(n63) );
  XOR2_X1 U85 ( .A(n41), .B(n63), .Z(SUM[8]) );
  NAND2_X1 U86 ( .A1(n40), .A2(B[8]), .ZN(n64) );
  NAND2_X1 U87 ( .A1(carry[8]), .A2(A[8]), .ZN(n65) );
  NAND2_X1 U88 ( .A1(B[8]), .A2(A[8]), .ZN(n66) );
  NAND3_X1 U89 ( .A1(n64), .A2(n65), .A3(n66), .ZN(carry[9]) );
  XOR2_X1 U90 ( .A(B[9]), .B(A[9]), .Z(n67) );
  XOR2_X1 U91 ( .A(n7), .B(n67), .Z(SUM[9]) );
  NAND2_X1 U92 ( .A1(n7), .A2(B[9]), .ZN(n68) );
  NAND2_X1 U93 ( .A1(carry[9]), .A2(A[9]), .ZN(n69) );
  NAND2_X1 U94 ( .A1(B[9]), .A2(A[9]), .ZN(n70) );
  NAND3_X1 U95 ( .A1(n68), .A2(n69), .A3(n70), .ZN(carry[10]) );
  XOR2_X1 U96 ( .A(B[1]), .B(A[1]), .Z(n71) );
  XOR2_X1 U97 ( .A(n79), .B(n71), .Z(SUM[1]) );
  NAND2_X1 U98 ( .A1(n79), .A2(B[1]), .ZN(n72) );
  NAND2_X1 U99 ( .A1(n79), .A2(A[1]), .ZN(n73) );
  NAND2_X1 U100 ( .A1(B[1]), .A2(A[1]), .ZN(n74) );
  NAND3_X1 U101 ( .A1(n72), .A2(n73), .A3(n74), .ZN(carry[2]) );
  XOR2_X1 U102 ( .A(B[2]), .B(A[2]), .Z(n75) );
  XOR2_X1 U103 ( .A(n58), .B(n75), .Z(SUM[2]) );
  NAND2_X1 U104 ( .A1(n57), .A2(B[2]), .ZN(n76) );
  NAND2_X1 U105 ( .A1(carry[2]), .A2(A[2]), .ZN(n77) );
  NAND2_X1 U106 ( .A1(B[2]), .A2(A[2]), .ZN(n78) );
  NAND3_X1 U107 ( .A1(n76), .A2(n77), .A3(n78), .ZN(carry[3]) );
  XOR2_X1 U108 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_8_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n17, n18, n19,
         n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76, n77,
         n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94, n96,
         n98, n99, n100, n101, n102, n103, n104, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370;

  FA_X1 U17 ( .A(n74), .B(n21), .CI(n314), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n313), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n317), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n316), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n319), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n92), .B(n80), .CI(n99), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  XNOR2_X1 U157 ( .A(n206), .B(n223), .ZN(product[14]) );
  AND3_X2 U158 ( .A1(n298), .A2(n299), .A3(n300), .ZN(n206) );
  BUF_X1 U159 ( .A(b[1]), .Z(n207) );
  BUF_X2 U160 ( .A(b[0]), .Z(n292) );
  NAND3_X1 U161 ( .A1(n303), .A2(n304), .A3(n305), .ZN(n49) );
  CLKBUF_X1 U162 ( .A(n242), .Z(n208) );
  CLKBUF_X1 U163 ( .A(n104), .Z(n209) );
  NAND3_X1 U164 ( .A1(n298), .A2(n299), .A3(n300), .ZN(n210) );
  NAND3_X1 U165 ( .A1(n298), .A2(n299), .A3(n300), .ZN(n211) );
  CLKBUF_X1 U166 ( .A(b[3]), .Z(n212) );
  CLKBUF_X1 U167 ( .A(n56), .Z(n213) );
  CLKBUF_X1 U168 ( .A(n233), .Z(n214) );
  NAND3_X1 U169 ( .A1(n283), .A2(n284), .A3(n285), .ZN(n215) );
  CLKBUF_X1 U170 ( .A(n239), .Z(n216) );
  NAND2_X1 U171 ( .A1(b[1]), .A2(a[1]), .ZN(n219) );
  NAND2_X1 U172 ( .A1(n217), .A2(n218), .ZN(n220) );
  NAND2_X1 U173 ( .A1(n219), .A2(n220), .ZN(n367) );
  INV_X1 U174 ( .A(b[1]), .ZN(n217) );
  INV_X1 U175 ( .A(a[1]), .ZN(n218) );
  AND2_X1 U176 ( .A1(n231), .A2(n234), .ZN(n221) );
  AND3_X1 U177 ( .A1(n224), .A2(n225), .A3(n226), .ZN(product[15]) );
  XOR2_X1 U178 ( .A(n311), .B(n15), .Z(n223) );
  NAND2_X1 U179 ( .A1(n211), .A2(n311), .ZN(n224) );
  NAND2_X1 U180 ( .A1(n210), .A2(n15), .ZN(n225) );
  NAND2_X1 U181 ( .A1(n311), .A2(n15), .ZN(n226) );
  CLKBUF_X1 U182 ( .A(n266), .Z(n227) );
  CLKBUF_X1 U183 ( .A(n347), .Z(n228) );
  XOR2_X1 U184 ( .A(a[6]), .B(n315), .Z(n347) );
  CLKBUF_X3 U185 ( .A(a[3]), .Z(n229) );
  XNOR2_X1 U186 ( .A(a[2]), .B(a[1]), .ZN(n230) );
  OAI22_X1 U187 ( .A1(n327), .A2(n328), .B1(n248), .B2(n329), .ZN(n231) );
  XOR2_X1 U188 ( .A(n209), .B(n72), .Z(product[1]) );
  NAND3_X1 U189 ( .A1(n264), .A2(n265), .A3(n227), .ZN(n232) );
  NAND2_X1 U190 ( .A1(n242), .A2(n40), .ZN(n233) );
  CLKBUF_X1 U191 ( .A(n102), .Z(n234) );
  XOR2_X1 U192 ( .A(n102), .B(n231), .Z(n56) );
  CLKBUF_X1 U193 ( .A(n212), .Z(n235) );
  NAND2_X1 U194 ( .A1(n18), .A2(n4), .ZN(n236) );
  AND2_X1 U195 ( .A1(n104), .A2(n72), .ZN(n237) );
  NAND3_X1 U196 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n238) );
  NAND3_X1 U197 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n239) );
  NAND3_X1 U198 ( .A1(n283), .A2(n284), .A3(n285), .ZN(n240) );
  NAND3_X1 U199 ( .A1(n287), .A2(n288), .A3(n289), .ZN(n241) );
  NAND3_X1 U200 ( .A1(n275), .A2(n276), .A3(n277), .ZN(n242) );
  NAND3_X1 U201 ( .A1(n255), .A2(n254), .A3(n256), .ZN(n243) );
  NAND3_X1 U202 ( .A1(n306), .A2(n307), .A3(n308), .ZN(n244) );
  NAND3_X1 U203 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n245) );
  CLKBUF_X1 U204 ( .A(n236), .Z(n246) );
  BUF_X2 U205 ( .A(n326), .Z(n247) );
  BUF_X2 U206 ( .A(n326), .Z(n248) );
  XNOR2_X1 U207 ( .A(a[2]), .B(a[1]), .ZN(n326) );
  XOR2_X1 U208 ( .A(n33), .B(n28), .Z(n249) );
  XOR2_X1 U209 ( .A(n245), .B(n249), .Z(product[9]) );
  NAND2_X1 U210 ( .A1(n245), .A2(n33), .ZN(n250) );
  NAND2_X1 U211 ( .A1(n7), .A2(n28), .ZN(n251) );
  NAND2_X1 U212 ( .A1(n33), .A2(n28), .ZN(n252) );
  NAND3_X1 U213 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n6) );
  XOR2_X1 U214 ( .A(n103), .B(n96), .Z(n253) );
  XOR2_X1 U215 ( .A(n237), .B(n253), .Z(product[2]) );
  NAND2_X1 U216 ( .A1(n103), .A2(n237), .ZN(n254) );
  NAND2_X1 U217 ( .A1(n237), .A2(n96), .ZN(n255) );
  NAND2_X1 U218 ( .A1(n103), .A2(n96), .ZN(n256) );
  NAND3_X1 U219 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n13) );
  XNOR2_X2 U220 ( .A(a[4]), .B(a[3]), .ZN(n336) );
  XOR2_X1 U221 ( .A(n27), .B(n24), .Z(n257) );
  XOR2_X1 U222 ( .A(n216), .B(n257), .Z(product[10]) );
  NAND2_X1 U223 ( .A1(n239), .A2(n27), .ZN(n258) );
  NAND2_X1 U224 ( .A1(n6), .A2(n24), .ZN(n259) );
  NAND2_X1 U225 ( .A1(n27), .A2(n24), .ZN(n260) );
  NAND3_X1 U226 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n5) );
  NAND3_X1 U227 ( .A1(n264), .A2(n266), .A3(n265), .ZN(n261) );
  XNOR2_X1 U228 ( .A(n207), .B(a[1]), .ZN(n262) );
  XOR2_X1 U229 ( .A(n213), .B(n71), .Z(n263) );
  XOR2_X1 U230 ( .A(n243), .B(n263), .Z(product[3]) );
  NAND2_X1 U231 ( .A1(n56), .A2(n243), .ZN(n264) );
  NAND2_X1 U232 ( .A1(n13), .A2(n71), .ZN(n265) );
  NAND2_X1 U233 ( .A1(n56), .A2(n71), .ZN(n266) );
  NAND3_X1 U234 ( .A1(n266), .A2(n265), .A3(n264), .ZN(n12) );
  NAND3_X1 U235 ( .A1(n233), .A2(n280), .A3(n281), .ZN(n267) );
  NAND3_X1 U236 ( .A1(n214), .A2(n280), .A3(n281), .ZN(n268) );
  NAND3_X1 U237 ( .A1(n287), .A2(n288), .A3(n289), .ZN(n269) );
  NAND2_X2 U238 ( .A1(n336), .A2(n365), .ZN(n338) );
  XOR2_X1 U239 ( .A(n34), .B(n39), .Z(n270) );
  XOR2_X1 U240 ( .A(n268), .B(n270), .Z(product[8]) );
  NAND2_X1 U241 ( .A1(n267), .A2(n34), .ZN(n271) );
  NAND2_X1 U242 ( .A1(n8), .A2(n39), .ZN(n272) );
  NAND2_X1 U243 ( .A1(n34), .A2(n39), .ZN(n273) );
  NAND3_X1 U244 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n7) );
  XOR2_X1 U245 ( .A(n46), .B(n49), .Z(n274) );
  XOR2_X1 U246 ( .A(n244), .B(n274), .Z(product[6]) );
  NAND2_X1 U247 ( .A1(n244), .A2(n46), .ZN(n275) );
  NAND2_X1 U248 ( .A1(n10), .A2(n49), .ZN(n276) );
  NAND2_X1 U249 ( .A1(n46), .A2(n49), .ZN(n277) );
  NAND3_X1 U250 ( .A1(n275), .A2(n276), .A3(n277), .ZN(n9) );
  XOR2_X1 U251 ( .A(n40), .B(n45), .Z(n278) );
  XOR2_X1 U252 ( .A(n208), .B(n278), .Z(product[7]) );
  NAND2_X1 U253 ( .A1(n242), .A2(n40), .ZN(n279) );
  NAND2_X1 U254 ( .A1(n9), .A2(n45), .ZN(n280) );
  NAND2_X1 U255 ( .A1(n40), .A2(n45), .ZN(n281) );
  NAND3_X1 U256 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n8) );
  XOR2_X1 U257 ( .A(n54), .B(n221), .Z(n282) );
  XOR2_X1 U258 ( .A(n232), .B(n282), .Z(product[4]) );
  NAND2_X1 U259 ( .A1(n12), .A2(n54), .ZN(n283) );
  NAND2_X1 U260 ( .A1(n261), .A2(n221), .ZN(n284) );
  NAND2_X1 U261 ( .A1(n54), .A2(n221), .ZN(n285) );
  NAND3_X1 U262 ( .A1(n283), .A2(n284), .A3(n285), .ZN(n11) );
  XOR2_X1 U263 ( .A(n23), .B(n20), .Z(n286) );
  XOR2_X1 U264 ( .A(n238), .B(n286), .Z(product[11]) );
  NAND2_X1 U265 ( .A1(n238), .A2(n23), .ZN(n287) );
  NAND2_X1 U266 ( .A1(n5), .A2(n20), .ZN(n288) );
  NAND2_X1 U267 ( .A1(n23), .A2(n20), .ZN(n289) );
  NAND3_X1 U268 ( .A1(n287), .A2(n288), .A3(n289), .ZN(n4) );
  NAND3_X1 U269 ( .A1(n236), .A2(n295), .A3(n294), .ZN(n290) );
  NAND3_X1 U270 ( .A1(n294), .A2(n295), .A3(n246), .ZN(n291) );
  XOR2_X1 U271 ( .A(n301), .B(n52), .Z(n50) );
  INV_X1 U272 ( .A(n15), .ZN(n310) );
  INV_X1 U273 ( .A(n345), .ZN(n314) );
  INV_X1 U274 ( .A(n21), .ZN(n313) );
  INV_X1 U275 ( .A(n325), .ZN(n319) );
  INV_X1 U276 ( .A(n334), .ZN(n317) );
  INV_X1 U277 ( .A(b[0]), .ZN(n309) );
  INV_X1 U278 ( .A(n356), .ZN(n311) );
  INV_X1 U279 ( .A(n31), .ZN(n316) );
  INV_X1 U280 ( .A(a[0]), .ZN(n320) );
  INV_X1 U281 ( .A(a[5]), .ZN(n315) );
  INV_X1 U282 ( .A(a[7]), .ZN(n312) );
  XOR2_X1 U283 ( .A(n19), .B(n18), .Z(n293) );
  XOR2_X1 U284 ( .A(n293), .B(n269), .Z(product[12]) );
  NAND2_X1 U285 ( .A1(n19), .A2(n18), .ZN(n294) );
  NAND2_X1 U286 ( .A1(n241), .A2(n19), .ZN(n295) );
  NAND2_X1 U287 ( .A1(n18), .A2(n4), .ZN(n296) );
  NAND3_X1 U288 ( .A1(n295), .A2(n296), .A3(n294), .ZN(n3) );
  XOR2_X1 U289 ( .A(n17), .B(n310), .Z(n297) );
  XOR2_X1 U290 ( .A(n297), .B(n291), .Z(product[13]) );
  NAND2_X1 U291 ( .A1(n17), .A2(n310), .ZN(n298) );
  NAND2_X1 U292 ( .A1(n17), .A2(n290), .ZN(n299) );
  NAND2_X1 U293 ( .A1(n310), .A2(n3), .ZN(n300) );
  XOR2_X1 U294 ( .A(n93), .B(n100), .Z(n301) );
  XOR2_X1 U295 ( .A(n53), .B(n240), .Z(n302) );
  XOR2_X1 U296 ( .A(n302), .B(n50), .Z(product[5]) );
  NAND2_X1 U297 ( .A1(n93), .A2(n100), .ZN(n303) );
  NAND2_X1 U298 ( .A1(n93), .A2(n52), .ZN(n304) );
  NAND2_X1 U299 ( .A1(n100), .A2(n52), .ZN(n305) );
  NAND2_X1 U300 ( .A1(n215), .A2(n53), .ZN(n306) );
  NAND2_X1 U301 ( .A1(n53), .A2(n50), .ZN(n307) );
  NAND2_X1 U302 ( .A1(n11), .A2(n50), .ZN(n308) );
  NAND3_X1 U303 ( .A1(n306), .A2(n307), .A3(n308), .ZN(n10) );
  INV_X1 U304 ( .A(a[3]), .ZN(n318) );
  NAND2_X2 U305 ( .A1(n230), .A2(n364), .ZN(n328) );
  NOR2_X1 U306 ( .A1(n320), .A2(n309), .ZN(product[0]) );
  OAI22_X1 U307 ( .A1(n321), .A2(n322), .B1(n323), .B2(n320), .ZN(n99) );
  OAI22_X1 U308 ( .A1(n323), .A2(n322), .B1(n324), .B2(n320), .ZN(n98) );
  XNOR2_X1 U309 ( .A(b[6]), .B(a[1]), .ZN(n323) );
  OAI22_X1 U310 ( .A1(n320), .A2(n324), .B1(n322), .B2(n324), .ZN(n325) );
  XNOR2_X1 U311 ( .A(b[7]), .B(a[1]), .ZN(n324) );
  NOR2_X1 U312 ( .A1(n247), .A2(n309), .ZN(n96) );
  XNOR2_X1 U313 ( .A(n229), .B(n292), .ZN(n327) );
  OAI22_X1 U314 ( .A1(n329), .A2(n328), .B1(n248), .B2(n330), .ZN(n94) );
  XNOR2_X1 U315 ( .A(b[1]), .B(n229), .ZN(n329) );
  OAI22_X1 U316 ( .A1(n330), .A2(n328), .B1(n247), .B2(n331), .ZN(n93) );
  XNOR2_X1 U317 ( .A(b[2]), .B(n229), .ZN(n330) );
  OAI22_X1 U318 ( .A1(n331), .A2(n328), .B1(n248), .B2(n332), .ZN(n92) );
  XNOR2_X1 U319 ( .A(n212), .B(n229), .ZN(n331) );
  OAI22_X1 U320 ( .A1(n332), .A2(n328), .B1(n248), .B2(n333), .ZN(n91) );
  XNOR2_X1 U321 ( .A(b[4]), .B(n229), .ZN(n332) );
  OAI22_X1 U322 ( .A1(n335), .A2(n247), .B1(n328), .B2(n335), .ZN(n334) );
  NOR2_X1 U323 ( .A1(n336), .A2(n309), .ZN(n88) );
  OAI22_X1 U324 ( .A1(n337), .A2(n338), .B1(n336), .B2(n339), .ZN(n87) );
  XNOR2_X1 U325 ( .A(a[5]), .B(n292), .ZN(n337) );
  OAI22_X1 U326 ( .A1(n339), .A2(n338), .B1(n336), .B2(n340), .ZN(n86) );
  XNOR2_X1 U327 ( .A(n207), .B(a[5]), .ZN(n339) );
  OAI22_X1 U328 ( .A1(n340), .A2(n338), .B1(n336), .B2(n341), .ZN(n85) );
  XNOR2_X1 U329 ( .A(b[2]), .B(a[5]), .ZN(n340) );
  OAI22_X1 U330 ( .A1(n341), .A2(n338), .B1(n336), .B2(n342), .ZN(n84) );
  XNOR2_X1 U331 ( .A(n235), .B(a[5]), .ZN(n341) );
  OAI22_X1 U332 ( .A1(n342), .A2(n338), .B1(n336), .B2(n343), .ZN(n83) );
  XNOR2_X1 U333 ( .A(b[4]), .B(a[5]), .ZN(n342) );
  OAI22_X1 U334 ( .A1(n343), .A2(n338), .B1(n336), .B2(n344), .ZN(n82) );
  XNOR2_X1 U335 ( .A(b[5]), .B(a[5]), .ZN(n343) );
  OAI22_X1 U336 ( .A1(n346), .A2(n336), .B1(n338), .B2(n346), .ZN(n345) );
  NOR2_X1 U337 ( .A1(n347), .A2(n309), .ZN(n80) );
  OAI22_X1 U338 ( .A1(n348), .A2(n349), .B1(n347), .B2(n350), .ZN(n79) );
  XNOR2_X1 U339 ( .A(a[7]), .B(n292), .ZN(n348) );
  OAI22_X1 U340 ( .A1(n351), .A2(n349), .B1(n228), .B2(n352), .ZN(n77) );
  OAI22_X1 U341 ( .A1(n352), .A2(n349), .B1(n228), .B2(n353), .ZN(n76) );
  XNOR2_X1 U342 ( .A(n235), .B(a[7]), .ZN(n352) );
  OAI22_X1 U343 ( .A1(n353), .A2(n349), .B1(n228), .B2(n354), .ZN(n75) );
  XNOR2_X1 U344 ( .A(b[4]), .B(a[7]), .ZN(n353) );
  OAI22_X1 U345 ( .A1(n354), .A2(n349), .B1(n228), .B2(n355), .ZN(n74) );
  XNOR2_X1 U346 ( .A(b[5]), .B(a[7]), .ZN(n354) );
  OAI22_X1 U347 ( .A1(n357), .A2(n228), .B1(n349), .B2(n357), .ZN(n356) );
  OAI21_X1 U348 ( .B1(n292), .B2(n218), .A(n322), .ZN(n72) );
  OAI21_X1 U349 ( .B1(n318), .B2(n328), .A(n358), .ZN(n71) );
  OR3_X1 U350 ( .A1(n247), .A2(n292), .A3(n318), .ZN(n358) );
  OAI21_X1 U351 ( .B1(n315), .B2(n338), .A(n359), .ZN(n70) );
  OR3_X1 U352 ( .A1(n336), .A2(n292), .A3(n315), .ZN(n359) );
  OAI21_X1 U353 ( .B1(n312), .B2(n349), .A(n360), .ZN(n69) );
  OR3_X1 U354 ( .A1(n347), .A2(n292), .A3(n312), .ZN(n360) );
  XNOR2_X1 U355 ( .A(n361), .B(n362), .ZN(n38) );
  OR2_X1 U356 ( .A1(n361), .A2(n362), .ZN(n37) );
  OAI22_X1 U357 ( .A1(n333), .A2(n328), .B1(n248), .B2(n363), .ZN(n362) );
  XNOR2_X1 U358 ( .A(b[5]), .B(n229), .ZN(n333) );
  OAI22_X1 U359 ( .A1(n350), .A2(n349), .B1(n228), .B2(n351), .ZN(n361) );
  XNOR2_X1 U360 ( .A(b[2]), .B(a[7]), .ZN(n351) );
  XNOR2_X1 U361 ( .A(n207), .B(a[7]), .ZN(n350) );
  OAI22_X1 U362 ( .A1(n363), .A2(n328), .B1(n247), .B2(n335), .ZN(n31) );
  XNOR2_X1 U363 ( .A(b[7]), .B(n229), .ZN(n335) );
  XNOR2_X1 U364 ( .A(n318), .B(a[2]), .ZN(n364) );
  XNOR2_X1 U365 ( .A(b[6]), .B(n229), .ZN(n363) );
  OAI22_X1 U366 ( .A1(n344), .A2(n338), .B1(n336), .B2(n346), .ZN(n21) );
  XNOR2_X1 U367 ( .A(b[7]), .B(a[5]), .ZN(n346) );
  XNOR2_X1 U368 ( .A(n315), .B(a[4]), .ZN(n365) );
  XNOR2_X1 U369 ( .A(b[6]), .B(a[5]), .ZN(n344) );
  OAI22_X1 U370 ( .A1(n355), .A2(n349), .B1(n228), .B2(n357), .ZN(n15) );
  XNOR2_X1 U371 ( .A(b[7]), .B(a[7]), .ZN(n357) );
  NAND2_X1 U372 ( .A1(n347), .A2(n366), .ZN(n349) );
  XNOR2_X1 U373 ( .A(n312), .B(a[6]), .ZN(n366) );
  XNOR2_X1 U374 ( .A(b[6]), .B(a[7]), .ZN(n355) );
  OAI22_X1 U375 ( .A1(n292), .A2(n322), .B1(n367), .B2(n320), .ZN(n104) );
  OAI22_X1 U376 ( .A1(n262), .A2(n322), .B1(n368), .B2(n320), .ZN(n103) );
  OAI22_X1 U377 ( .A1(n368), .A2(n322), .B1(n369), .B2(n320), .ZN(n102) );
  XNOR2_X1 U378 ( .A(b[2]), .B(a[1]), .ZN(n368) );
  OAI22_X1 U379 ( .A1(n322), .A2(n369), .B1(n370), .B2(n320), .ZN(n101) );
  XNOR2_X1 U380 ( .A(b[3]), .B(a[1]), .ZN(n369) );
  OAI22_X1 U381 ( .A1(n370), .A2(n322), .B1(n321), .B2(n320), .ZN(n100) );
  XNOR2_X1 U382 ( .A(b[5]), .B(a[1]), .ZN(n321) );
  NAND2_X1 U383 ( .A1(a[1]), .A2(n320), .ZN(n322) );
  XNOR2_X1 U384 ( .A(b[4]), .B(a[1]), .ZN(n370) );
endmodule


module mac_8 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  mac_8_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_8_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_7_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63;
  wire   [15:1] carry;

  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n63), .CO(carry[2]), .S(SUM[1]) );
  XNOR2_X1 U1 ( .A(B[15]), .B(A[15]), .ZN(n1) );
  CLKBUF_X1 U2 ( .A(carry[8]), .Z(n2) );
  XOR2_X1 U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR2_X1 U4 ( .A(n2), .B(n3), .Z(SUM[8]) );
  NAND2_X1 U5 ( .A1(carry[8]), .A2(B[8]), .ZN(n4) );
  NAND2_X1 U6 ( .A1(carry[8]), .A2(A[8]), .ZN(n5) );
  NAND2_X1 U7 ( .A1(B[8]), .A2(A[8]), .ZN(n6) );
  NAND3_X1 U8 ( .A1(n4), .A2(n5), .A3(n6), .ZN(carry[9]) );
  CLKBUF_X1 U9 ( .A(n46), .Z(n7) );
  FA_X1 U10 ( .A(A[1]), .B(B[1]), .CI(n63), .CO(n8) );
  FA_X1 U11 ( .A(A[1]), .B(B[1]), .CI(n63), .CO(n9) );
  AND2_X2 U12 ( .A1(B[0]), .A2(A[0]), .ZN(n63) );
  CLKBUF_X1 U13 ( .A(carry[11]), .Z(n10) );
  NAND3_X1 U14 ( .A1(n15), .A2(n16), .A3(n17), .ZN(n11) );
  NAND3_X1 U15 ( .A1(n15), .A2(n16), .A3(n17), .ZN(n12) );
  CLKBUF_X1 U16 ( .A(n34), .Z(n13) );
  XOR2_X1 U17 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR2_X1 U18 ( .A(n9), .B(n14), .Z(SUM[2]) );
  NAND2_X1 U19 ( .A1(n8), .A2(B[2]), .ZN(n15) );
  NAND2_X1 U20 ( .A1(carry[2]), .A2(A[2]), .ZN(n16) );
  NAND2_X1 U21 ( .A1(B[2]), .A2(A[2]), .ZN(n17) );
  NAND3_X1 U22 ( .A1(n15), .A2(n16), .A3(n17), .ZN(carry[3]) );
  NAND3_X1 U23 ( .A1(n20), .A2(n21), .A3(n22), .ZN(n18) );
  XOR2_X1 U24 ( .A(B[3]), .B(A[3]), .Z(n19) );
  XOR2_X1 U25 ( .A(n12), .B(n19), .Z(SUM[3]) );
  NAND2_X1 U26 ( .A1(n11), .A2(B[3]), .ZN(n20) );
  NAND2_X1 U27 ( .A1(carry[3]), .A2(A[3]), .ZN(n21) );
  NAND2_X1 U28 ( .A1(B[3]), .A2(A[3]), .ZN(n22) );
  NAND3_X1 U29 ( .A1(n20), .A2(n21), .A3(n22), .ZN(carry[4]) );
  NAND3_X1 U30 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n23) );
  NAND3_X1 U31 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n24) );
  NAND3_X1 U32 ( .A1(n31), .A2(n32), .A3(n33), .ZN(n25) );
  XNOR2_X1 U33 ( .A(carry[15]), .B(n1), .ZN(SUM[15]) );
  XOR2_X1 U34 ( .A(B[11]), .B(A[11]), .Z(n26) );
  XOR2_X1 U35 ( .A(n10), .B(n26), .Z(SUM[11]) );
  NAND2_X1 U36 ( .A1(carry[11]), .A2(B[11]), .ZN(n27) );
  NAND2_X1 U37 ( .A1(carry[11]), .A2(A[11]), .ZN(n28) );
  NAND2_X1 U38 ( .A1(B[11]), .A2(A[11]), .ZN(n29) );
  NAND3_X1 U39 ( .A1(n27), .A2(n28), .A3(n29), .ZN(carry[12]) );
  XOR2_X1 U40 ( .A(B[4]), .B(A[4]), .Z(n30) );
  XOR2_X1 U41 ( .A(n18), .B(n30), .Z(SUM[4]) );
  NAND2_X1 U42 ( .A1(n18), .A2(B[4]), .ZN(n31) );
  NAND2_X1 U43 ( .A1(carry[4]), .A2(A[4]), .ZN(n32) );
  NAND2_X1 U44 ( .A1(B[4]), .A2(A[4]), .ZN(n33) );
  NAND3_X1 U45 ( .A1(n31), .A2(n32), .A3(n33), .ZN(carry[5]) );
  NAND3_X1 U46 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n34) );
  NAND3_X1 U47 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n35) );
  XOR2_X1 U48 ( .A(B[12]), .B(A[12]), .Z(n36) );
  XOR2_X1 U49 ( .A(n24), .B(n36), .Z(SUM[12]) );
  NAND2_X1 U50 ( .A1(n23), .A2(B[12]), .ZN(n37) );
  NAND2_X1 U51 ( .A1(carry[12]), .A2(A[12]), .ZN(n38) );
  NAND2_X1 U52 ( .A1(B[12]), .A2(A[12]), .ZN(n39) );
  NAND3_X1 U53 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[13]) );
  XOR2_X1 U54 ( .A(B[5]), .B(A[5]), .Z(n40) );
  XOR2_X1 U55 ( .A(carry[5]), .B(n40), .Z(SUM[5]) );
  NAND2_X1 U56 ( .A1(n25), .A2(B[5]), .ZN(n41) );
  NAND2_X1 U57 ( .A1(n25), .A2(A[5]), .ZN(n42) );
  NAND2_X1 U58 ( .A1(B[5]), .A2(A[5]), .ZN(n43) );
  NAND3_X1 U59 ( .A1(n41), .A2(n42), .A3(n43), .ZN(carry[6]) );
  NAND3_X1 U60 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n44) );
  NAND3_X1 U61 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n45) );
  NAND3_X1 U62 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n46) );
  XOR2_X1 U63 ( .A(B[13]), .B(A[13]), .Z(n47) );
  XOR2_X1 U64 ( .A(n13), .B(n47), .Z(SUM[13]) );
  NAND2_X1 U65 ( .A1(n34), .A2(B[13]), .ZN(n48) );
  NAND2_X1 U66 ( .A1(carry[13]), .A2(A[13]), .ZN(n49) );
  NAND2_X1 U67 ( .A1(B[13]), .A2(A[13]), .ZN(n50) );
  XOR2_X1 U68 ( .A(B[6]), .B(A[6]), .Z(n51) );
  XOR2_X1 U69 ( .A(carry[6]), .B(n51), .Z(SUM[6]) );
  NAND2_X1 U70 ( .A1(n35), .A2(B[6]), .ZN(n52) );
  NAND2_X1 U71 ( .A1(n35), .A2(A[6]), .ZN(n53) );
  NAND2_X1 U72 ( .A1(B[6]), .A2(A[6]), .ZN(n54) );
  NAND3_X1 U73 ( .A1(n52), .A2(n53), .A3(n54), .ZN(carry[7]) );
  XOR2_X1 U74 ( .A(B[14]), .B(A[14]), .Z(n55) );
  XOR2_X1 U75 ( .A(n45), .B(n55), .Z(SUM[14]) );
  NAND2_X1 U76 ( .A1(n44), .A2(B[14]), .ZN(n56) );
  NAND2_X1 U77 ( .A1(n44), .A2(A[14]), .ZN(n57) );
  NAND2_X1 U78 ( .A1(B[14]), .A2(A[14]), .ZN(n58) );
  NAND3_X1 U79 ( .A1(n56), .A2(n57), .A3(n58), .ZN(carry[15]) );
  XOR2_X1 U80 ( .A(B[7]), .B(A[7]), .Z(n59) );
  XOR2_X1 U81 ( .A(n7), .B(n59), .Z(SUM[7]) );
  NAND2_X1 U82 ( .A1(n46), .A2(B[7]), .ZN(n60) );
  NAND2_X1 U83 ( .A1(carry[7]), .A2(A[7]), .ZN(n61) );
  NAND2_X1 U84 ( .A1(B[7]), .A2(A[7]), .ZN(n62) );
  NAND3_X1 U85 ( .A1(n60), .A2(n61), .A3(n62), .ZN(carry[8]) );
  XOR2_X1 U86 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_7_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n310), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n309), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n313), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n312), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n314), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  XOR2_X2 U157 ( .A(a[2]), .B(n315), .Z(n294) );
  CLKBUF_X1 U158 ( .A(b[1]), .Z(n206) );
  INV_X1 U159 ( .A(n15), .ZN(n306) );
  NAND3_X1 U160 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n207) );
  CLKBUF_X1 U161 ( .A(n363), .Z(n208) );
  CLKBUF_X1 U162 ( .A(n251), .Z(n209) );
  AND2_X1 U163 ( .A1(n227), .A2(n102), .ZN(n210) );
  CLKBUF_X1 U164 ( .A(n56), .Z(n211) );
  XNOR2_X1 U165 ( .A(a[2]), .B(a[1]), .ZN(n322) );
  CLKBUF_X1 U166 ( .A(n246), .Z(n212) );
  CLKBUF_X1 U167 ( .A(n301), .Z(n213) );
  CLKBUF_X1 U168 ( .A(n271), .Z(n214) );
  CLKBUF_X1 U169 ( .A(n14), .Z(n215) );
  NAND3_X1 U170 ( .A1(n301), .A2(n302), .A3(n303), .ZN(n216) );
  NAND3_X1 U171 ( .A1(n213), .A2(n302), .A3(n303), .ZN(n217) );
  BUF_X1 U172 ( .A(n305), .Z(n218) );
  XOR2_X1 U173 ( .A(n100), .B(n93), .Z(n219) );
  XOR2_X1 U174 ( .A(n52), .B(n219), .Z(n50) );
  NAND2_X1 U175 ( .A1(n52), .A2(n100), .ZN(n220) );
  NAND2_X1 U176 ( .A1(n52), .A2(n93), .ZN(n221) );
  NAND2_X1 U177 ( .A1(n100), .A2(n93), .ZN(n222) );
  NAND3_X1 U178 ( .A1(n220), .A2(n221), .A3(n222), .ZN(n49) );
  CLKBUF_X1 U179 ( .A(n262), .Z(n223) );
  NAND3_X1 U180 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n224) );
  NAND3_X1 U181 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n225) );
  NAND3_X1 U182 ( .A1(n214), .A2(n272), .A3(n273), .ZN(n226) );
  OAI22_X1 U183 ( .A1(n323), .A2(n324), .B1(n294), .B2(n325), .ZN(n227) );
  CLKBUF_X1 U184 ( .A(n277), .Z(n228) );
  NAND3_X1 U185 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n229) );
  CLKBUF_X1 U186 ( .A(n224), .Z(n230) );
  NAND3_X1 U187 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n231) );
  XOR2_X1 U188 ( .A(n23), .B(n20), .Z(n232) );
  XOR2_X1 U189 ( .A(n226), .B(n232), .Z(product[11]) );
  NAND2_X1 U190 ( .A1(n225), .A2(n23), .ZN(n233) );
  NAND2_X1 U191 ( .A1(n5), .A2(n20), .ZN(n234) );
  NAND2_X1 U192 ( .A1(n23), .A2(n20), .ZN(n235) );
  NAND3_X1 U193 ( .A1(n234), .A2(n233), .A3(n235), .ZN(n4) );
  XOR2_X1 U194 ( .A(n17), .B(n306), .Z(n236) );
  XOR2_X1 U195 ( .A(n217), .B(n236), .Z(product[13]) );
  NAND2_X1 U196 ( .A1(n216), .A2(n17), .ZN(n237) );
  NAND2_X1 U197 ( .A1(n3), .A2(n306), .ZN(n238) );
  NAND2_X1 U198 ( .A1(n17), .A2(n306), .ZN(n239) );
  NAND3_X1 U199 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n2) );
  NAND2_X1 U200 ( .A1(a[4]), .A2(a[3]), .ZN(n242) );
  NAND2_X1 U201 ( .A1(n240), .A2(n241), .ZN(n243) );
  NAND2_X2 U202 ( .A1(n242), .A2(n243), .ZN(n332) );
  INV_X1 U203 ( .A(a[4]), .ZN(n240) );
  INV_X1 U204 ( .A(a[3]), .ZN(n241) );
  NAND3_X1 U205 ( .A1(n281), .A2(n282), .A3(n283), .ZN(n244) );
  CLKBUF_X1 U206 ( .A(n260), .Z(n245) );
  NAND3_X1 U207 ( .A1(n255), .A2(n256), .A3(n254), .ZN(n246) );
  NAND3_X1 U208 ( .A1(n252), .A2(n251), .A3(n250), .ZN(n247) );
  NAND3_X1 U209 ( .A1(n250), .A2(n209), .A3(n252), .ZN(n248) );
  XOR2_X1 U210 ( .A(n103), .B(n96), .Z(n249) );
  XOR2_X1 U211 ( .A(n249), .B(n215), .Z(product[2]) );
  NAND2_X1 U212 ( .A1(n103), .A2(n96), .ZN(n250) );
  NAND2_X1 U213 ( .A1(n103), .A2(n14), .ZN(n251) );
  NAND2_X1 U214 ( .A1(n96), .A2(n14), .ZN(n252) );
  NAND3_X1 U215 ( .A1(n252), .A2(n251), .A3(n250), .ZN(n13) );
  XOR2_X1 U216 ( .A(n211), .B(n71), .Z(n253) );
  XOR2_X1 U217 ( .A(n253), .B(n248), .Z(product[3]) );
  NAND2_X1 U218 ( .A1(n56), .A2(n71), .ZN(n254) );
  NAND2_X1 U219 ( .A1(n56), .A2(n247), .ZN(n255) );
  NAND2_X1 U220 ( .A1(n13), .A2(n71), .ZN(n256) );
  NAND3_X1 U221 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n12) );
  INV_X2 U222 ( .A(n305), .ZN(n304) );
  XOR2_X1 U223 ( .A(a[3]), .B(n305), .Z(n323) );
  NAND3_X1 U224 ( .A1(n286), .A2(n287), .A3(n288), .ZN(n257) );
  NAND3_X1 U225 ( .A1(n277), .A2(n278), .A3(n279), .ZN(n258) );
  NAND3_X1 U226 ( .A1(n228), .A2(n278), .A3(n279), .ZN(n259) );
  NAND3_X1 U227 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n260) );
  XOR2_X1 U228 ( .A(n95), .B(n102), .Z(n56) );
  XOR2_X1 U229 ( .A(n54), .B(n210), .Z(n261) );
  XOR2_X1 U230 ( .A(n212), .B(n261), .Z(product[4]) );
  NAND2_X1 U231 ( .A1(n246), .A2(n54), .ZN(n262) );
  NAND2_X1 U232 ( .A1(n12), .A2(n210), .ZN(n263) );
  NAND2_X1 U233 ( .A1(n54), .A2(n210), .ZN(n264) );
  NAND3_X1 U234 ( .A1(n223), .A2(n263), .A3(n264), .ZN(n11) );
  XOR2_X1 U235 ( .A(n33), .B(n28), .Z(n265) );
  XOR2_X1 U236 ( .A(n259), .B(n265), .Z(product[9]) );
  NAND2_X1 U237 ( .A1(n258), .A2(n33), .ZN(n266) );
  NAND2_X1 U238 ( .A1(n7), .A2(n28), .ZN(n267) );
  NAND2_X1 U239 ( .A1(n33), .A2(n28), .ZN(n268) );
  NAND3_X1 U240 ( .A1(n267), .A2(n266), .A3(n268), .ZN(n6) );
  CLKBUF_X1 U241 ( .A(b[1]), .Z(n269) );
  XOR2_X1 U242 ( .A(n27), .B(n24), .Z(n270) );
  XOR2_X1 U243 ( .A(n245), .B(n270), .Z(product[10]) );
  NAND2_X1 U244 ( .A1(n260), .A2(n27), .ZN(n271) );
  NAND2_X1 U245 ( .A1(n6), .A2(n24), .ZN(n272) );
  NAND2_X1 U246 ( .A1(n27), .A2(n24), .ZN(n273) );
  NAND3_X1 U247 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n5) );
  NAND3_X1 U248 ( .A1(n290), .A2(n291), .A3(n292), .ZN(n274) );
  CLKBUF_X1 U249 ( .A(n244), .Z(n275) );
  XOR2_X1 U250 ( .A(n34), .B(n39), .Z(n276) );
  XOR2_X1 U251 ( .A(n274), .B(n276), .Z(product[8]) );
  NAND2_X1 U252 ( .A1(n274), .A2(n34), .ZN(n277) );
  NAND2_X1 U253 ( .A1(n8), .A2(n39), .ZN(n278) );
  NAND2_X1 U254 ( .A1(n34), .A2(n39), .ZN(n279) );
  NAND3_X1 U255 ( .A1(n277), .A2(n278), .A3(n279), .ZN(n7) );
  XOR2_X1 U256 ( .A(n50), .B(n53), .Z(n280) );
  XOR2_X1 U257 ( .A(n11), .B(n280), .Z(product[5]) );
  NAND2_X1 U258 ( .A1(n207), .A2(n50), .ZN(n281) );
  NAND2_X1 U259 ( .A1(n229), .A2(n53), .ZN(n282) );
  NAND2_X1 U260 ( .A1(n50), .A2(n53), .ZN(n283) );
  NAND3_X1 U261 ( .A1(n281), .A2(n282), .A3(n283), .ZN(n10) );
  CLKBUF_X1 U262 ( .A(n257), .Z(n284) );
  XOR2_X1 U263 ( .A(n46), .B(n49), .Z(n285) );
  XOR2_X1 U264 ( .A(n275), .B(n285), .Z(product[6]) );
  NAND2_X1 U265 ( .A1(n244), .A2(n46), .ZN(n286) );
  NAND2_X1 U266 ( .A1(n10), .A2(n49), .ZN(n287) );
  NAND2_X1 U267 ( .A1(n46), .A2(n49), .ZN(n288) );
  NAND3_X1 U268 ( .A1(n286), .A2(n287), .A3(n288), .ZN(n9) );
  XOR2_X1 U269 ( .A(n40), .B(n45), .Z(n289) );
  XOR2_X1 U270 ( .A(n284), .B(n289), .Z(product[7]) );
  NAND2_X1 U271 ( .A1(n257), .A2(n40), .ZN(n290) );
  NAND2_X1 U272 ( .A1(n9), .A2(n45), .ZN(n291) );
  NAND2_X1 U273 ( .A1(n40), .A2(n45), .ZN(n292) );
  NAND3_X1 U274 ( .A1(n290), .A2(n291), .A3(n292), .ZN(n8) );
  NAND2_X2 U275 ( .A1(n322), .A2(n360), .ZN(n324) );
  NAND2_X2 U276 ( .A1(n332), .A2(n361), .ZN(n334) );
  XOR2_X1 U277 ( .A(a[2]), .B(n315), .Z(n293) );
  XNOR2_X1 U278 ( .A(n231), .B(n295), .ZN(product[14]) );
  XNOR2_X1 U279 ( .A(n307), .B(n15), .ZN(n295) );
  XNOR2_X1 U280 ( .A(n230), .B(n296), .ZN(product[12]) );
  XNOR2_X1 U281 ( .A(n19), .B(n18), .ZN(n296) );
  AND3_X1 U282 ( .A1(n298), .A2(n299), .A3(n300), .ZN(product[15]) );
  INV_X1 U283 ( .A(n330), .ZN(n313) );
  OAI22_X1 U284 ( .A1(n351), .A2(n345), .B1(n343), .B2(n353), .ZN(n15) );
  INV_X1 U285 ( .A(n341), .ZN(n310) );
  INV_X1 U286 ( .A(n21), .ZN(n309) );
  INV_X1 U287 ( .A(n321), .ZN(n314) );
  INV_X1 U288 ( .A(n31), .ZN(n312) );
  INV_X1 U289 ( .A(b[0]), .ZN(n305) );
  INV_X1 U290 ( .A(a[0]), .ZN(n316) );
  INV_X1 U291 ( .A(a[5]), .ZN(n311) );
  INV_X1 U292 ( .A(a[7]), .ZN(n308) );
  NAND2_X1 U293 ( .A1(n231), .A2(n307), .ZN(n298) );
  NAND2_X1 U294 ( .A1(n2), .A2(n15), .ZN(n299) );
  NAND2_X1 U295 ( .A1(n307), .A2(n15), .ZN(n300) );
  NAND2_X1 U296 ( .A1(n224), .A2(n19), .ZN(n301) );
  NAND2_X1 U297 ( .A1(n4), .A2(n18), .ZN(n302) );
  NAND2_X1 U298 ( .A1(n19), .A2(n18), .ZN(n303) );
  NAND3_X1 U299 ( .A1(n301), .A2(n302), .A3(n303), .ZN(n3) );
  INV_X1 U300 ( .A(n352), .ZN(n307) );
  INV_X1 U301 ( .A(a[1]), .ZN(n315) );
  XOR2_X2 U302 ( .A(a[6]), .B(n311), .Z(n343) );
  NOR2_X1 U303 ( .A1(n316), .A2(n218), .ZN(product[0]) );
  OAI22_X1 U304 ( .A1(n317), .A2(n318), .B1(n319), .B2(n316), .ZN(n99) );
  OAI22_X1 U305 ( .A1(n319), .A2(n318), .B1(n320), .B2(n316), .ZN(n98) );
  XNOR2_X1 U306 ( .A(b[6]), .B(a[1]), .ZN(n319) );
  OAI22_X1 U307 ( .A1(n316), .A2(n320), .B1(n318), .B2(n320), .ZN(n321) );
  XNOR2_X1 U308 ( .A(b[7]), .B(a[1]), .ZN(n320) );
  NOR2_X1 U309 ( .A1(n293), .A2(n218), .ZN(n96) );
  OAI22_X1 U310 ( .A1(n323), .A2(n324), .B1(n294), .B2(n325), .ZN(n95) );
  OAI22_X1 U311 ( .A1(n325), .A2(n324), .B1(n294), .B2(n326), .ZN(n94) );
  XNOR2_X1 U312 ( .A(n206), .B(a[3]), .ZN(n325) );
  OAI22_X1 U313 ( .A1(n326), .A2(n324), .B1(n293), .B2(n327), .ZN(n93) );
  XNOR2_X1 U314 ( .A(b[2]), .B(a[3]), .ZN(n326) );
  OAI22_X1 U315 ( .A1(n327), .A2(n324), .B1(n294), .B2(n328), .ZN(n92) );
  XNOR2_X1 U316 ( .A(b[3]), .B(a[3]), .ZN(n327) );
  OAI22_X1 U317 ( .A1(n328), .A2(n324), .B1(n294), .B2(n329), .ZN(n91) );
  XNOR2_X1 U318 ( .A(b[4]), .B(a[3]), .ZN(n328) );
  OAI22_X1 U319 ( .A1(n331), .A2(n293), .B1(n324), .B2(n331), .ZN(n330) );
  NOR2_X1 U320 ( .A1(n332), .A2(n218), .ZN(n88) );
  OAI22_X1 U321 ( .A1(n333), .A2(n334), .B1(n332), .B2(n335), .ZN(n87) );
  XNOR2_X1 U322 ( .A(a[5]), .B(n304), .ZN(n333) );
  OAI22_X1 U323 ( .A1(n335), .A2(n334), .B1(n332), .B2(n336), .ZN(n86) );
  XNOR2_X1 U324 ( .A(n269), .B(a[5]), .ZN(n335) );
  OAI22_X1 U325 ( .A1(n336), .A2(n334), .B1(n332), .B2(n337), .ZN(n85) );
  XNOR2_X1 U326 ( .A(b[2]), .B(a[5]), .ZN(n336) );
  OAI22_X1 U327 ( .A1(n337), .A2(n334), .B1(n332), .B2(n338), .ZN(n84) );
  XNOR2_X1 U328 ( .A(b[3]), .B(a[5]), .ZN(n337) );
  OAI22_X1 U329 ( .A1(n338), .A2(n334), .B1(n332), .B2(n339), .ZN(n83) );
  XNOR2_X1 U330 ( .A(b[4]), .B(a[5]), .ZN(n338) );
  OAI22_X1 U331 ( .A1(n339), .A2(n334), .B1(n332), .B2(n340), .ZN(n82) );
  XNOR2_X1 U332 ( .A(b[5]), .B(a[5]), .ZN(n339) );
  OAI22_X1 U333 ( .A1(n342), .A2(n332), .B1(n334), .B2(n342), .ZN(n341) );
  NOR2_X1 U334 ( .A1(n343), .A2(n218), .ZN(n80) );
  OAI22_X1 U335 ( .A1(n344), .A2(n345), .B1(n343), .B2(n346), .ZN(n79) );
  XNOR2_X1 U336 ( .A(a[7]), .B(n304), .ZN(n344) );
  OAI22_X1 U337 ( .A1(n347), .A2(n345), .B1(n343), .B2(n348), .ZN(n77) );
  OAI22_X1 U338 ( .A1(n348), .A2(n345), .B1(n343), .B2(n349), .ZN(n76) );
  XNOR2_X1 U339 ( .A(b[3]), .B(a[7]), .ZN(n348) );
  OAI22_X1 U340 ( .A1(n349), .A2(n345), .B1(n343), .B2(n350), .ZN(n75) );
  XNOR2_X1 U341 ( .A(b[4]), .B(a[7]), .ZN(n349) );
  OAI22_X1 U342 ( .A1(n350), .A2(n345), .B1(n343), .B2(n351), .ZN(n74) );
  XNOR2_X1 U343 ( .A(b[5]), .B(a[7]), .ZN(n350) );
  OAI22_X1 U344 ( .A1(n353), .A2(n343), .B1(n345), .B2(n353), .ZN(n352) );
  OAI21_X1 U345 ( .B1(n304), .B2(n315), .A(n318), .ZN(n72) );
  OAI21_X1 U346 ( .B1(n241), .B2(n324), .A(n354), .ZN(n71) );
  OR3_X1 U347 ( .A1(n293), .A2(n304), .A3(n241), .ZN(n354) );
  OAI21_X1 U348 ( .B1(n311), .B2(n334), .A(n355), .ZN(n70) );
  OR3_X1 U349 ( .A1(n332), .A2(n304), .A3(n311), .ZN(n355) );
  OAI21_X1 U350 ( .B1(n308), .B2(n345), .A(n356), .ZN(n69) );
  OR3_X1 U351 ( .A1(n343), .A2(n304), .A3(n308), .ZN(n356) );
  XNOR2_X1 U352 ( .A(n357), .B(n358), .ZN(n38) );
  OR2_X1 U353 ( .A1(n357), .A2(n358), .ZN(n37) );
  OAI22_X1 U354 ( .A1(n329), .A2(n324), .B1(n293), .B2(n359), .ZN(n358) );
  XNOR2_X1 U355 ( .A(b[5]), .B(a[3]), .ZN(n329) );
  OAI22_X1 U356 ( .A1(n346), .A2(n345), .B1(n343), .B2(n347), .ZN(n357) );
  XNOR2_X1 U357 ( .A(b[2]), .B(a[7]), .ZN(n347) );
  XNOR2_X1 U358 ( .A(n269), .B(a[7]), .ZN(n346) );
  OAI22_X1 U359 ( .A1(n359), .A2(n324), .B1(n294), .B2(n331), .ZN(n31) );
  XNOR2_X1 U360 ( .A(b[7]), .B(a[3]), .ZN(n331) );
  XNOR2_X1 U361 ( .A(n241), .B(a[2]), .ZN(n360) );
  XNOR2_X1 U362 ( .A(b[6]), .B(a[3]), .ZN(n359) );
  OAI22_X1 U363 ( .A1(n340), .A2(n334), .B1(n332), .B2(n342), .ZN(n21) );
  XNOR2_X1 U364 ( .A(b[7]), .B(a[5]), .ZN(n342) );
  XNOR2_X1 U365 ( .A(n311), .B(a[4]), .ZN(n361) );
  XNOR2_X1 U366 ( .A(b[6]), .B(a[5]), .ZN(n340) );
  XNOR2_X1 U367 ( .A(b[7]), .B(a[7]), .ZN(n353) );
  NAND2_X1 U368 ( .A1(n343), .A2(n362), .ZN(n345) );
  XNOR2_X1 U369 ( .A(n308), .B(a[6]), .ZN(n362) );
  XNOR2_X1 U370 ( .A(b[6]), .B(a[7]), .ZN(n351) );
  OAI22_X1 U371 ( .A1(n304), .A2(n318), .B1(n363), .B2(n316), .ZN(n104) );
  OAI22_X1 U372 ( .A1(n208), .A2(n318), .B1(n364), .B2(n316), .ZN(n103) );
  XNOR2_X1 U373 ( .A(b[1]), .B(a[1]), .ZN(n363) );
  OAI22_X1 U374 ( .A1(n364), .A2(n318), .B1(n365), .B2(n316), .ZN(n102) );
  XNOR2_X1 U375 ( .A(b[2]), .B(a[1]), .ZN(n364) );
  OAI22_X1 U376 ( .A1(n365), .A2(n318), .B1(n366), .B2(n316), .ZN(n101) );
  XNOR2_X1 U377 ( .A(b[3]), .B(a[1]), .ZN(n365) );
  OAI22_X1 U378 ( .A1(n366), .A2(n318), .B1(n317), .B2(n316), .ZN(n100) );
  XNOR2_X1 U379 ( .A(b[5]), .B(a[1]), .ZN(n317) );
  NAND2_X1 U380 ( .A1(a[1]), .A2(n316), .ZN(n318) );
  XNOR2_X1 U381 ( .A(b[4]), .B(a[1]), .ZN(n366) );
endmodule


module mac_7 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_7_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_7_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_6_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;
  wire   [15:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .S(SUM[15]) );
  NAND3_X1 U1 ( .A1(n81), .A2(n82), .A3(n83), .ZN(n1) );
  NAND2_X1 U2 ( .A1(n7), .A2(B[11]), .ZN(n2) );
  AND2_X1 U3 ( .A1(B[0]), .A2(A[0]), .ZN(n84) );
  NAND3_X1 U4 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n3) );
  NAND3_X1 U5 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n4) );
  NAND3_X1 U6 ( .A1(n2), .A2(n51), .A3(n52), .ZN(n5) );
  CLKBUF_X1 U7 ( .A(n15), .Z(n6) );
  NAND3_X1 U8 ( .A1(n20), .A2(n21), .A3(n22), .ZN(n7) );
  NAND3_X1 U9 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n8) );
  NAND3_X1 U10 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n9) );
  NAND3_X1 U11 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n10) );
  CLKBUF_X1 U12 ( .A(n1), .Z(n11) );
  CLKBUF_X1 U13 ( .A(n3), .Z(n12) );
  NAND3_X1 U14 ( .A1(n32), .A2(n33), .A3(n34), .ZN(n13) );
  NAND3_X1 U15 ( .A1(n32), .A2(n33), .A3(n34), .ZN(n14) );
  NAND3_X1 U16 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n15) );
  CLKBUF_X1 U17 ( .A(n7), .Z(n16) );
  CLKBUF_X1 U18 ( .A(n8), .Z(n17) );
  CLKBUF_X1 U19 ( .A(n55), .Z(n18) );
  XOR2_X1 U20 ( .A(B[10]), .B(A[10]), .Z(n19) );
  XOR2_X1 U21 ( .A(n17), .B(n19), .Z(SUM[10]) );
  NAND2_X1 U22 ( .A1(n8), .A2(B[10]), .ZN(n20) );
  NAND2_X1 U23 ( .A1(carry[10]), .A2(A[10]), .ZN(n21) );
  NAND2_X1 U24 ( .A1(B[10]), .A2(A[10]), .ZN(n22) );
  NAND3_X1 U25 ( .A1(n20), .A2(n21), .A3(n22), .ZN(carry[11]) );
  XOR2_X1 U26 ( .A(B[8]), .B(A[8]), .Z(n23) );
  XOR2_X1 U27 ( .A(n11), .B(n23), .Z(SUM[8]) );
  NAND2_X1 U28 ( .A1(n1), .A2(B[8]), .ZN(n24) );
  NAND2_X1 U29 ( .A1(carry[8]), .A2(A[8]), .ZN(n25) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n26) );
  NAND3_X1 U31 ( .A1(n24), .A2(n25), .A3(n26), .ZN(carry[9]) );
  XOR2_X1 U32 ( .A(B[9]), .B(A[9]), .Z(n27) );
  XOR2_X1 U33 ( .A(n12), .B(n27), .Z(SUM[9]) );
  NAND2_X1 U34 ( .A1(n3), .A2(B[9]), .ZN(n28) );
  NAND2_X1 U35 ( .A1(carry[9]), .A2(A[9]), .ZN(n29) );
  NAND2_X1 U36 ( .A1(B[9]), .A2(A[9]), .ZN(n30) );
  NAND3_X1 U37 ( .A1(n28), .A2(n29), .A3(n30), .ZN(carry[10]) );
  XOR2_X1 U38 ( .A(B[1]), .B(A[1]), .Z(n31) );
  XOR2_X1 U39 ( .A(n84), .B(n31), .Z(SUM[1]) );
  NAND2_X1 U40 ( .A1(n84), .A2(B[1]), .ZN(n32) );
  NAND2_X1 U41 ( .A1(n84), .A2(A[1]), .ZN(n33) );
  NAND2_X1 U42 ( .A1(B[1]), .A2(A[1]), .ZN(n34) );
  NAND3_X1 U43 ( .A1(n32), .A2(n33), .A3(n34), .ZN(carry[2]) );
  XOR2_X1 U44 ( .A(B[3]), .B(A[3]), .Z(n35) );
  XOR2_X1 U45 ( .A(n6), .B(n35), .Z(SUM[3]) );
  NAND2_X1 U46 ( .A1(n15), .A2(B[3]), .ZN(n36) );
  NAND2_X1 U47 ( .A1(carry[3]), .A2(A[3]), .ZN(n37) );
  NAND2_X1 U48 ( .A1(B[3]), .A2(A[3]), .ZN(n38) );
  NAND3_X1 U49 ( .A1(n36), .A2(n37), .A3(n38), .ZN(carry[4]) );
  CLKBUF_X1 U50 ( .A(n67), .Z(n39) );
  CLKBUF_X1 U51 ( .A(n64), .Z(n40) );
  CLKBUF_X1 U52 ( .A(carry[13]), .Z(n41) );
  NAND3_X1 U53 ( .A1(n2), .A2(n51), .A3(n52), .ZN(n42) );
  NAND3_X1 U54 ( .A1(n54), .A2(n18), .A3(n56), .ZN(n43) );
  NAND3_X1 U55 ( .A1(n63), .A2(n40), .A3(n65), .ZN(n44) );
  XOR2_X1 U56 ( .A(B[2]), .B(A[2]), .Z(n45) );
  XOR2_X1 U57 ( .A(n14), .B(n45), .Z(SUM[2]) );
  NAND2_X1 U58 ( .A1(n13), .A2(B[2]), .ZN(n46) );
  NAND2_X1 U59 ( .A1(carry[2]), .A2(A[2]), .ZN(n47) );
  NAND2_X1 U60 ( .A1(B[2]), .A2(A[2]), .ZN(n48) );
  NAND3_X1 U61 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[3]) );
  XOR2_X1 U62 ( .A(B[11]), .B(A[11]), .Z(n49) );
  XOR2_X1 U63 ( .A(n16), .B(n49), .Z(SUM[11]) );
  NAND2_X1 U64 ( .A1(n7), .A2(B[11]), .ZN(n50) );
  NAND2_X1 U65 ( .A1(carry[11]), .A2(A[11]), .ZN(n51) );
  NAND2_X1 U66 ( .A1(B[11]), .A2(A[11]), .ZN(n52) );
  NAND3_X1 U67 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[12]) );
  XOR2_X1 U68 ( .A(B[4]), .B(A[4]), .Z(n53) );
  XOR2_X1 U69 ( .A(n10), .B(n53), .Z(SUM[4]) );
  NAND2_X1 U70 ( .A1(n9), .A2(B[4]), .ZN(n54) );
  NAND2_X1 U71 ( .A1(carry[4]), .A2(A[4]), .ZN(n55) );
  NAND2_X1 U72 ( .A1(B[4]), .A2(A[4]), .ZN(n56) );
  NAND3_X1 U73 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[5]) );
  NAND3_X1 U74 ( .A1(n60), .A2(n59), .A3(n61), .ZN(n57) );
  XOR2_X1 U75 ( .A(B[12]), .B(A[12]), .Z(n58) );
  XOR2_X1 U76 ( .A(n42), .B(n58), .Z(SUM[12]) );
  NAND2_X1 U77 ( .A1(n5), .A2(B[12]), .ZN(n59) );
  NAND2_X1 U78 ( .A1(carry[12]), .A2(A[12]), .ZN(n60) );
  NAND2_X1 U79 ( .A1(B[12]), .A2(A[12]), .ZN(n61) );
  NAND3_X1 U80 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[13]) );
  XOR2_X1 U81 ( .A(B[5]), .B(A[5]), .Z(n62) );
  XOR2_X1 U82 ( .A(n43), .B(n62), .Z(SUM[5]) );
  NAND2_X1 U83 ( .A1(carry[5]), .A2(B[5]), .ZN(n63) );
  NAND2_X1 U84 ( .A1(carry[5]), .A2(A[5]), .ZN(n64) );
  NAND2_X1 U85 ( .A1(B[5]), .A2(A[5]), .ZN(n65) );
  NAND3_X1 U86 ( .A1(n63), .A2(n64), .A3(n65), .ZN(carry[6]) );
  NAND3_X1 U87 ( .A1(n69), .A2(n70), .A3(n71), .ZN(n66) );
  NAND3_X1 U88 ( .A1(n73), .A2(n74), .A3(n75), .ZN(n67) );
  XOR2_X1 U89 ( .A(B[13]), .B(A[13]), .Z(n68) );
  XOR2_X1 U90 ( .A(n41), .B(n68), .Z(SUM[13]) );
  NAND2_X1 U91 ( .A1(n57), .A2(B[13]), .ZN(n69) );
  NAND2_X1 U92 ( .A1(carry[13]), .A2(A[13]), .ZN(n70) );
  NAND2_X1 U93 ( .A1(B[13]), .A2(A[13]), .ZN(n71) );
  NAND3_X1 U94 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[14]) );
  XOR2_X1 U95 ( .A(B[6]), .B(A[6]), .Z(n72) );
  XOR2_X1 U96 ( .A(n44), .B(n72), .Z(SUM[6]) );
  NAND2_X1 U97 ( .A1(n4), .A2(B[6]), .ZN(n73) );
  NAND2_X1 U98 ( .A1(carry[6]), .A2(A[6]), .ZN(n74) );
  NAND2_X1 U99 ( .A1(B[6]), .A2(A[6]), .ZN(n75) );
  NAND3_X1 U100 ( .A1(n73), .A2(n74), .A3(n75), .ZN(carry[7]) );
  XOR2_X1 U101 ( .A(B[14]), .B(A[14]), .Z(n76) );
  XOR2_X1 U102 ( .A(carry[14]), .B(n76), .Z(SUM[14]) );
  NAND2_X1 U103 ( .A1(n66), .A2(B[14]), .ZN(n77) );
  NAND2_X1 U104 ( .A1(n66), .A2(A[14]), .ZN(n78) );
  NAND2_X1 U105 ( .A1(B[14]), .A2(A[14]), .ZN(n79) );
  NAND3_X1 U106 ( .A1(n77), .A2(n78), .A3(n79), .ZN(carry[15]) );
  XOR2_X1 U107 ( .A(B[7]), .B(A[7]), .Z(n80) );
  XOR2_X1 U108 ( .A(n39), .B(n80), .Z(SUM[7]) );
  NAND2_X1 U109 ( .A1(n67), .A2(B[7]), .ZN(n81) );
  NAND2_X1 U110 ( .A1(carry[7]), .A2(A[7]), .ZN(n82) );
  NAND2_X1 U111 ( .A1(B[7]), .A2(A[7]), .ZN(n83) );
  NAND3_X1 U112 ( .A1(n81), .A2(n82), .A3(n83), .ZN(carry[8]) );
  XOR2_X1 U113 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_6_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18, n19,
         n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76, n77,
         n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94, n95,
         n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n312), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n311), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n315), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n314), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n317), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n94), .B(n88), .CI(n101), .CO(n53), .S(n54) );
  NAND2_X1 U157 ( .A1(n335), .A2(n364), .ZN(n337) );
  AND2_X1 U158 ( .A1(n207), .A2(n102), .ZN(n206) );
  OAI22_X1 U159 ( .A1(n326), .A2(n327), .B1(n297), .B2(n328), .ZN(n207) );
  CLKBUF_X1 U160 ( .A(a[5]), .Z(n208) );
  INV_X1 U161 ( .A(n306), .ZN(n209) );
  XOR2_X1 U162 ( .A(n95), .B(n102), .Z(n56) );
  CLKBUF_X1 U163 ( .A(b[3]), .Z(n210) );
  NAND2_X2 U164 ( .A1(n230), .A2(n231), .ZN(n211) );
  NAND2_X1 U165 ( .A1(n230), .A2(n231), .ZN(n335) );
  NAND3_X1 U166 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n212) );
  CLKBUF_X1 U167 ( .A(n270), .Z(n213) );
  CLKBUF_X1 U168 ( .A(n56), .Z(n214) );
  XNOR2_X1 U169 ( .A(b[1]), .B(a[1]), .ZN(n215) );
  AND2_X1 U170 ( .A1(n104), .A2(n72), .ZN(n216) );
  CLKBUF_X1 U171 ( .A(n301), .Z(n217) );
  CLKBUF_X1 U172 ( .A(n268), .Z(n218) );
  CLKBUF_X1 U173 ( .A(b[1]), .Z(n219) );
  CLKBUF_X1 U174 ( .A(b[1]), .Z(n220) );
  NAND3_X1 U175 ( .A1(n282), .A2(n281), .A3(n283), .ZN(n221) );
  CLKBUF_X1 U176 ( .A(n305), .Z(n222) );
  CLKBUF_X1 U177 ( .A(n4), .Z(n223) );
  CLKBUF_X1 U178 ( .A(n295), .Z(n224) );
  NAND3_X1 U179 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n225) );
  NAND3_X1 U180 ( .A1(n237), .A2(n236), .A3(n238), .ZN(n226) );
  NAND3_X1 U181 ( .A1(n294), .A2(n224), .A3(n296), .ZN(n227) );
  NAND2_X1 U182 ( .A1(a[4]), .A2(a[3]), .ZN(n230) );
  NAND2_X1 U183 ( .A1(n228), .A2(n229), .ZN(n231) );
  INV_X1 U184 ( .A(a[4]), .ZN(n228) );
  INV_X1 U185 ( .A(a[3]), .ZN(n229) );
  CLKBUF_X1 U186 ( .A(n7), .Z(n232) );
  NAND3_X1 U187 ( .A1(n259), .A2(n258), .A3(n260), .ZN(n233) );
  NAND3_X1 U188 ( .A1(n244), .A2(n243), .A3(n245), .ZN(n234) );
  XOR2_X1 U189 ( .A(n34), .B(n39), .Z(n235) );
  XOR2_X1 U190 ( .A(n227), .B(n235), .Z(product[8]) );
  NAND2_X1 U191 ( .A1(n212), .A2(n34), .ZN(n236) );
  NAND2_X1 U192 ( .A1(n8), .A2(n39), .ZN(n237) );
  NAND2_X1 U193 ( .A1(n34), .A2(n39), .ZN(n238) );
  NAND3_X1 U194 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n7) );
  CLKBUF_X1 U195 ( .A(n273), .Z(n239) );
  CLKBUF_X1 U196 ( .A(n5), .Z(n240) );
  CLKBUF_X1 U197 ( .A(n234), .Z(n241) );
  XOR2_X1 U198 ( .A(n33), .B(n28), .Z(n242) );
  XOR2_X1 U199 ( .A(n232), .B(n242), .Z(product[9]) );
  NAND2_X1 U200 ( .A1(n7), .A2(n33), .ZN(n243) );
  NAND2_X1 U201 ( .A1(n226), .A2(n28), .ZN(n244) );
  NAND2_X1 U202 ( .A1(n33), .A2(n28), .ZN(n245) );
  NAND3_X1 U203 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n6) );
  XOR2_X1 U204 ( .A(n103), .B(n96), .Z(n246) );
  XOR2_X1 U205 ( .A(n216), .B(n246), .Z(product[2]) );
  NAND2_X1 U206 ( .A1(n216), .A2(n103), .ZN(n247) );
  NAND2_X1 U207 ( .A1(n14), .A2(n96), .ZN(n248) );
  NAND2_X1 U208 ( .A1(n103), .A2(n96), .ZN(n249) );
  NAND3_X1 U209 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n13) );
  NAND3_X1 U210 ( .A1(n273), .A2(n272), .A3(n274), .ZN(n250) );
  NAND3_X1 U211 ( .A1(n239), .A2(n272), .A3(n274), .ZN(n251) );
  CLKBUF_X1 U212 ( .A(n304), .Z(n252) );
  CLKBUF_X1 U213 ( .A(n300), .Z(n253) );
  XNOR2_X1 U214 ( .A(n221), .B(n254), .ZN(product[14]) );
  XNOR2_X1 U215 ( .A(n309), .B(n15), .ZN(n254) );
  NAND3_X1 U216 ( .A1(n265), .A2(n264), .A3(n266), .ZN(n255) );
  AND3_X1 U217 ( .A1(n286), .A2(n285), .A3(n284), .ZN(product[15]) );
  XOR2_X1 U218 ( .A(n27), .B(n24), .Z(n257) );
  XOR2_X1 U219 ( .A(n241), .B(n257), .Z(product[10]) );
  NAND2_X1 U220 ( .A1(n6), .A2(n27), .ZN(n258) );
  NAND2_X1 U221 ( .A1(n234), .A2(n24), .ZN(n259) );
  NAND2_X1 U222 ( .A1(n27), .A2(n24), .ZN(n260) );
  NAND3_X1 U223 ( .A1(n259), .A2(n258), .A3(n260), .ZN(n5) );
  NAND3_X1 U224 ( .A1(n268), .A2(n269), .A3(n270), .ZN(n261) );
  NAND3_X1 U225 ( .A1(n218), .A2(n269), .A3(n213), .ZN(n262) );
  XOR2_X1 U226 ( .A(n23), .B(n20), .Z(n263) );
  XOR2_X1 U227 ( .A(n240), .B(n263), .Z(product[11]) );
  NAND2_X1 U228 ( .A1(n233), .A2(n23), .ZN(n264) );
  NAND2_X1 U229 ( .A1(n5), .A2(n20), .ZN(n265) );
  NAND2_X1 U230 ( .A1(n23), .A2(n20), .ZN(n266) );
  NAND3_X1 U231 ( .A1(n265), .A2(n264), .A3(n266), .ZN(n4) );
  XOR2_X1 U232 ( .A(n214), .B(n71), .Z(n267) );
  XOR2_X1 U233 ( .A(n13), .B(n267), .Z(product[3]) );
  NAND2_X1 U234 ( .A1(n13), .A2(n56), .ZN(n268) );
  NAND2_X1 U235 ( .A1(n225), .A2(n71), .ZN(n269) );
  NAND2_X1 U236 ( .A1(n56), .A2(n71), .ZN(n270) );
  NAND3_X1 U237 ( .A1(n268), .A2(n269), .A3(n270), .ZN(n12) );
  XOR2_X1 U238 ( .A(n18), .B(n19), .Z(n271) );
  XOR2_X1 U239 ( .A(n223), .B(n271), .Z(product[12]) );
  NAND2_X1 U240 ( .A1(n255), .A2(n18), .ZN(n272) );
  NAND2_X1 U241 ( .A1(n4), .A2(n19), .ZN(n273) );
  NAND2_X1 U242 ( .A1(n18), .A2(n19), .ZN(n274) );
  NAND3_X1 U243 ( .A1(n305), .A2(n304), .A3(n303), .ZN(n275) );
  NAND3_X1 U244 ( .A1(n303), .A2(n252), .A3(n222), .ZN(n276) );
  NAND3_X1 U245 ( .A1(n290), .A2(n291), .A3(n292), .ZN(n277) );
  NAND3_X1 U246 ( .A1(n282), .A2(n283), .A3(n281), .ZN(n278) );
  NAND3_X1 U247 ( .A1(n283), .A2(n281), .A3(n282), .ZN(n279) );
  XOR2_X1 U248 ( .A(n17), .B(n308), .Z(n280) );
  XOR2_X1 U249 ( .A(n280), .B(n251), .Z(product[13]) );
  NAND2_X1 U250 ( .A1(n17), .A2(n308), .ZN(n281) );
  NAND2_X1 U251 ( .A1(n17), .A2(n250), .ZN(n282) );
  NAND2_X1 U252 ( .A1(n308), .A2(n250), .ZN(n283) );
  NAND2_X1 U253 ( .A1(n309), .A2(n15), .ZN(n284) );
  NAND2_X1 U254 ( .A1(n279), .A2(n309), .ZN(n285) );
  NAND2_X1 U255 ( .A1(n278), .A2(n15), .ZN(n286) );
  NAND3_X1 U256 ( .A1(n300), .A2(n301), .A3(n299), .ZN(n287) );
  NAND3_X1 U257 ( .A1(n299), .A2(n253), .A3(n217), .ZN(n288) );
  XOR2_X1 U258 ( .A(n46), .B(n49), .Z(n289) );
  XOR2_X1 U259 ( .A(n276), .B(n289), .Z(product[6]) );
  NAND2_X1 U260 ( .A1(n275), .A2(n46), .ZN(n290) );
  NAND2_X1 U261 ( .A1(n10), .A2(n49), .ZN(n291) );
  NAND2_X1 U262 ( .A1(n46), .A2(n49), .ZN(n292) );
  NAND3_X1 U263 ( .A1(n290), .A2(n291), .A3(n292), .ZN(n9) );
  XOR2_X1 U264 ( .A(n40), .B(n45), .Z(n293) );
  XOR2_X1 U265 ( .A(n9), .B(n293), .Z(product[7]) );
  NAND2_X1 U266 ( .A1(n277), .A2(n40), .ZN(n294) );
  NAND2_X1 U267 ( .A1(n277), .A2(n45), .ZN(n295) );
  NAND2_X1 U268 ( .A1(n40), .A2(n45), .ZN(n296) );
  NAND3_X1 U269 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n8) );
  XNOR2_X2 U270 ( .A(a[2]), .B(a[1]), .ZN(n297) );
  XNOR2_X1 U271 ( .A(a[2]), .B(a[1]), .ZN(n325) );
  INV_X1 U272 ( .A(n15), .ZN(n308) );
  INV_X1 U273 ( .A(n21), .ZN(n311) );
  INV_X1 U274 ( .A(n344), .ZN(n312) );
  INV_X1 U275 ( .A(n324), .ZN(n317) );
  INV_X1 U276 ( .A(n333), .ZN(n315) );
  INV_X1 U277 ( .A(n31), .ZN(n314) );
  INV_X1 U278 ( .A(n355), .ZN(n309) );
  INV_X1 U279 ( .A(a[0]), .ZN(n319) );
  INV_X1 U280 ( .A(a[5]), .ZN(n313) );
  INV_X1 U281 ( .A(a[7]), .ZN(n310) );
  INV_X1 U282 ( .A(a[3]), .ZN(n316) );
  INV_X1 U283 ( .A(b[0]), .ZN(n307) );
  XOR2_X1 U284 ( .A(n54), .B(n206), .Z(n298) );
  XOR2_X1 U285 ( .A(n298), .B(n262), .Z(product[4]) );
  NAND2_X1 U286 ( .A1(n54), .A2(n206), .ZN(n299) );
  NAND2_X1 U287 ( .A1(n261), .A2(n54), .ZN(n300) );
  NAND2_X1 U288 ( .A1(n12), .A2(n206), .ZN(n301) );
  NAND3_X1 U289 ( .A1(n299), .A2(n300), .A3(n301), .ZN(n11) );
  XOR2_X1 U290 ( .A(n50), .B(n53), .Z(n302) );
  XOR2_X1 U291 ( .A(n302), .B(n288), .Z(product[5]) );
  NAND2_X1 U292 ( .A1(n50), .A2(n53), .ZN(n303) );
  NAND2_X1 U293 ( .A1(n50), .A2(n287), .ZN(n304) );
  NAND2_X1 U294 ( .A1(n11), .A2(n53), .ZN(n305) );
  NAND3_X1 U295 ( .A1(n304), .A2(n303), .A3(n305), .ZN(n10) );
  INV_X1 U296 ( .A(a[1]), .ZN(n318) );
  NAND2_X2 U297 ( .A1(n325), .A2(n363), .ZN(n327) );
  XOR2_X2 U298 ( .A(a[6]), .B(n313), .Z(n346) );
  INV_X1 U299 ( .A(n307), .ZN(n306) );
  NOR2_X1 U300 ( .A1(n319), .A2(n209), .ZN(product[0]) );
  OAI22_X1 U301 ( .A1(n320), .A2(n321), .B1(n322), .B2(n319), .ZN(n99) );
  OAI22_X1 U302 ( .A1(n322), .A2(n321), .B1(n323), .B2(n319), .ZN(n98) );
  XNOR2_X1 U303 ( .A(b[6]), .B(a[1]), .ZN(n322) );
  OAI22_X1 U304 ( .A1(n319), .A2(n323), .B1(n321), .B2(n323), .ZN(n324) );
  XNOR2_X1 U305 ( .A(b[7]), .B(a[1]), .ZN(n323) );
  NOR2_X1 U306 ( .A1(n297), .A2(n307), .ZN(n96) );
  OAI22_X1 U307 ( .A1(n326), .A2(n327), .B1(n297), .B2(n328), .ZN(n95) );
  XNOR2_X1 U308 ( .A(a[3]), .B(b[0]), .ZN(n326) );
  OAI22_X1 U309 ( .A1(n328), .A2(n327), .B1(n297), .B2(n329), .ZN(n94) );
  XNOR2_X1 U310 ( .A(n219), .B(a[3]), .ZN(n328) );
  OAI22_X1 U311 ( .A1(n329), .A2(n327), .B1(n297), .B2(n330), .ZN(n93) );
  XNOR2_X1 U312 ( .A(b[2]), .B(a[3]), .ZN(n329) );
  OAI22_X1 U313 ( .A1(n330), .A2(n327), .B1(n297), .B2(n331), .ZN(n92) );
  XNOR2_X1 U314 ( .A(n210), .B(a[3]), .ZN(n330) );
  OAI22_X1 U315 ( .A1(n331), .A2(n327), .B1(n297), .B2(n332), .ZN(n91) );
  XNOR2_X1 U316 ( .A(b[4]), .B(a[3]), .ZN(n331) );
  OAI22_X1 U317 ( .A1(n334), .A2(n297), .B1(n327), .B2(n334), .ZN(n333) );
  NOR2_X1 U318 ( .A1(n211), .A2(n209), .ZN(n88) );
  OAI22_X1 U319 ( .A1(n336), .A2(n337), .B1(n211), .B2(n338), .ZN(n87) );
  XNOR2_X1 U320 ( .A(a[5]), .B(n306), .ZN(n336) );
  OAI22_X1 U321 ( .A1(n338), .A2(n337), .B1(n211), .B2(n339), .ZN(n86) );
  XNOR2_X1 U322 ( .A(n220), .B(a[5]), .ZN(n338) );
  OAI22_X1 U323 ( .A1(n339), .A2(n337), .B1(n211), .B2(n340), .ZN(n85) );
  XNOR2_X1 U324 ( .A(b[2]), .B(a[5]), .ZN(n339) );
  OAI22_X1 U325 ( .A1(n340), .A2(n337), .B1(n211), .B2(n341), .ZN(n84) );
  XNOR2_X1 U326 ( .A(n210), .B(a[5]), .ZN(n340) );
  OAI22_X1 U327 ( .A1(n341), .A2(n337), .B1(n211), .B2(n342), .ZN(n83) );
  XNOR2_X1 U328 ( .A(b[4]), .B(n208), .ZN(n341) );
  OAI22_X1 U329 ( .A1(n342), .A2(n337), .B1(n211), .B2(n343), .ZN(n82) );
  XNOR2_X1 U330 ( .A(b[5]), .B(n208), .ZN(n342) );
  OAI22_X1 U331 ( .A1(n345), .A2(n211), .B1(n337), .B2(n345), .ZN(n344) );
  NOR2_X1 U332 ( .A1(n346), .A2(n209), .ZN(n80) );
  OAI22_X1 U333 ( .A1(n347), .A2(n348), .B1(n346), .B2(n349), .ZN(n79) );
  XNOR2_X1 U334 ( .A(a[7]), .B(n306), .ZN(n347) );
  OAI22_X1 U335 ( .A1(n350), .A2(n348), .B1(n346), .B2(n351), .ZN(n77) );
  OAI22_X1 U336 ( .A1(n351), .A2(n348), .B1(n346), .B2(n352), .ZN(n76) );
  XNOR2_X1 U337 ( .A(n210), .B(a[7]), .ZN(n351) );
  OAI22_X1 U338 ( .A1(n352), .A2(n348), .B1(n346), .B2(n353), .ZN(n75) );
  XNOR2_X1 U339 ( .A(b[4]), .B(a[7]), .ZN(n352) );
  OAI22_X1 U340 ( .A1(n353), .A2(n348), .B1(n346), .B2(n354), .ZN(n74) );
  XNOR2_X1 U341 ( .A(b[5]), .B(a[7]), .ZN(n353) );
  OAI22_X1 U342 ( .A1(n356), .A2(n346), .B1(n348), .B2(n356), .ZN(n355) );
  OAI21_X1 U343 ( .B1(b[0]), .B2(n318), .A(n321), .ZN(n72) );
  OAI21_X1 U344 ( .B1(n316), .B2(n327), .A(n357), .ZN(n71) );
  OR3_X1 U345 ( .A1(n297), .A2(n306), .A3(n316), .ZN(n357) );
  OAI21_X1 U346 ( .B1(n313), .B2(n337), .A(n358), .ZN(n70) );
  OR3_X1 U347 ( .A1(n335), .A2(n306), .A3(n313), .ZN(n358) );
  OAI21_X1 U348 ( .B1(n310), .B2(n348), .A(n359), .ZN(n69) );
  OR3_X1 U349 ( .A1(n346), .A2(n306), .A3(n310), .ZN(n359) );
  XNOR2_X1 U350 ( .A(n360), .B(n361), .ZN(n38) );
  OR2_X1 U351 ( .A1(n360), .A2(n361), .ZN(n37) );
  OAI22_X1 U352 ( .A1(n332), .A2(n327), .B1(n297), .B2(n362), .ZN(n361) );
  XNOR2_X1 U353 ( .A(b[5]), .B(a[3]), .ZN(n332) );
  OAI22_X1 U354 ( .A1(n349), .A2(n348), .B1(n346), .B2(n350), .ZN(n360) );
  XNOR2_X1 U355 ( .A(b[2]), .B(a[7]), .ZN(n350) );
  XNOR2_X1 U356 ( .A(b[1]), .B(a[7]), .ZN(n349) );
  OAI22_X1 U357 ( .A1(n362), .A2(n327), .B1(n297), .B2(n334), .ZN(n31) );
  XNOR2_X1 U358 ( .A(b[7]), .B(a[3]), .ZN(n334) );
  XNOR2_X1 U359 ( .A(n316), .B(a[2]), .ZN(n363) );
  XNOR2_X1 U360 ( .A(b[6]), .B(a[3]), .ZN(n362) );
  OAI22_X1 U361 ( .A1(n343), .A2(n337), .B1(n211), .B2(n345), .ZN(n21) );
  XNOR2_X1 U362 ( .A(b[7]), .B(n208), .ZN(n345) );
  XNOR2_X1 U363 ( .A(n313), .B(a[4]), .ZN(n364) );
  XNOR2_X1 U364 ( .A(b[6]), .B(n208), .ZN(n343) );
  OAI22_X1 U365 ( .A1(n354), .A2(n348), .B1(n346), .B2(n356), .ZN(n15) );
  XNOR2_X1 U366 ( .A(b[7]), .B(a[7]), .ZN(n356) );
  NAND2_X1 U367 ( .A1(n346), .A2(n365), .ZN(n348) );
  XNOR2_X1 U368 ( .A(n310), .B(a[6]), .ZN(n365) );
  XNOR2_X1 U369 ( .A(b[6]), .B(a[7]), .ZN(n354) );
  OAI22_X1 U370 ( .A1(b[0]), .A2(n321), .B1(n366), .B2(n319), .ZN(n104) );
  OAI22_X1 U371 ( .A1(n215), .A2(n321), .B1(n367), .B2(n319), .ZN(n103) );
  XNOR2_X1 U372 ( .A(b[1]), .B(a[1]), .ZN(n366) );
  OAI22_X1 U373 ( .A1(n367), .A2(n321), .B1(n368), .B2(n319), .ZN(n102) );
  XNOR2_X1 U374 ( .A(b[2]), .B(a[1]), .ZN(n367) );
  OAI22_X1 U375 ( .A1(n368), .A2(n321), .B1(n369), .B2(n319), .ZN(n101) );
  XNOR2_X1 U376 ( .A(b[3]), .B(a[1]), .ZN(n368) );
  OAI22_X1 U377 ( .A1(n369), .A2(n321), .B1(n320), .B2(n319), .ZN(n100) );
  XNOR2_X1 U378 ( .A(b[5]), .B(a[1]), .ZN(n320) );
  NAND2_X1 U379 ( .A1(a[1]), .A2(n319), .ZN(n321) );
  XNOR2_X1 U380 ( .A(b[4]), .B(a[1]), .ZN(n369) );
endmodule


module mac_6 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   n6, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, n2, n4;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(n6), .QN(n2) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_6_DW01_add_0 add_356 ( .A(pipeline), .B({mac_out[15:1], n6}), .CI(1'b0), 
        .SUM(sum) );
  mac_6_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n4), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n4), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n4), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n4), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n4), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n4), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n4), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n4), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n4), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n4), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n4), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n4), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n4), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n4), .ZN(N6) );
  INV_X1 U18 ( .A(n2), .ZN(mac_out[0]) );
  AND2_X1 U19 ( .A1(sum[0]), .A2(n4), .ZN(N3) );
  AND2_X1 U20 ( .A1(sum[15]), .A2(n4), .ZN(N18) );
  INV_X1 U21 ( .A(clear_acc), .ZN(n4) );
endmodule


module mac_5_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73;
  wire   [15:1] carry;

  CLKBUF_X1 U1 ( .A(carry[6]), .Z(n1) );
  NAND2_X1 U2 ( .A1(A[13]), .A2(B[13]), .ZN(n14) );
  AND2_X1 U3 ( .A1(B[0]), .A2(A[0]), .ZN(n73) );
  XOR2_X1 U4 ( .A(B[15]), .B(A[15]), .Z(n2) );
  XOR2_X1 U5 ( .A(carry[15]), .B(n2), .Z(SUM[15]) );
  NAND3_X1 U6 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n3) );
  XOR2_X1 U7 ( .A(B[4]), .B(A[4]), .Z(n4) );
  XOR2_X1 U8 ( .A(carry[4]), .B(n4), .Z(SUM[4]) );
  NAND2_X1 U9 ( .A1(carry[4]), .A2(B[4]), .ZN(n5) );
  NAND2_X1 U10 ( .A1(carry[4]), .A2(A[4]), .ZN(n6) );
  NAND2_X1 U11 ( .A1(B[4]), .A2(A[4]), .ZN(n7) );
  NAND3_X1 U12 ( .A1(n5), .A2(n6), .A3(n7), .ZN(carry[5]) );
  CLKBUF_X1 U13 ( .A(n40), .Z(n8) );
  XOR2_X1 U14 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U15 ( .A(carry[3]), .B(n9), .Z(SUM[3]) );
  NAND2_X1 U16 ( .A1(carry[3]), .A2(B[3]), .ZN(n10) );
  NAND2_X1 U17 ( .A1(carry[3]), .A2(A[3]), .ZN(n11) );
  NAND2_X1 U18 ( .A1(B[3]), .A2(A[3]), .ZN(n12) );
  NAND3_X1 U19 ( .A1(n10), .A2(n11), .A3(n12), .ZN(carry[4]) );
  XOR2_X1 U20 ( .A(A[13]), .B(B[13]), .Z(n13) );
  XOR2_X1 U21 ( .A(n13), .B(carry[13]), .Z(SUM[13]) );
  NAND2_X1 U22 ( .A1(A[13]), .A2(carry[13]), .ZN(n15) );
  NAND2_X1 U23 ( .A1(B[13]), .A2(carry[13]), .ZN(n16) );
  NAND3_X1 U24 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[14]) );
  XOR2_X1 U25 ( .A(A[14]), .B(B[14]), .Z(n17) );
  XOR2_X1 U26 ( .A(n17), .B(carry[14]), .Z(SUM[14]) );
  NAND2_X1 U27 ( .A1(A[14]), .A2(B[14]), .ZN(n18) );
  NAND2_X1 U28 ( .A1(A[14]), .A2(carry[14]), .ZN(n19) );
  NAND2_X1 U29 ( .A1(B[14]), .A2(carry[14]), .ZN(n20) );
  NAND3_X1 U30 ( .A1(n18), .A2(n19), .A3(n20), .ZN(carry[15]) );
  CLKBUF_X1 U31 ( .A(n32), .Z(n21) );
  XOR2_X1 U32 ( .A(B[5]), .B(A[5]), .Z(n22) );
  XOR2_X1 U33 ( .A(carry[5]), .B(n22), .Z(SUM[5]) );
  NAND2_X1 U34 ( .A1(carry[5]), .A2(B[5]), .ZN(n23) );
  NAND2_X1 U35 ( .A1(carry[5]), .A2(A[5]), .ZN(n24) );
  NAND2_X1 U36 ( .A1(B[5]), .A2(A[5]), .ZN(n25) );
  NAND3_X1 U37 ( .A1(n23), .A2(n24), .A3(n25), .ZN(carry[6]) );
  NAND3_X1 U38 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n26) );
  NAND3_X1 U39 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n27) );
  XOR2_X1 U40 ( .A(B[6]), .B(A[6]), .Z(n28) );
  XOR2_X1 U41 ( .A(n1), .B(n28), .Z(SUM[6]) );
  NAND2_X1 U42 ( .A1(carry[6]), .A2(B[6]), .ZN(n29) );
  NAND2_X1 U43 ( .A1(carry[6]), .A2(A[6]), .ZN(n30) );
  NAND2_X1 U44 ( .A1(B[6]), .A2(A[6]), .ZN(n31) );
  NAND3_X1 U45 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[7]) );
  NAND3_X1 U46 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n32) );
  NAND3_X1 U47 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n33) );
  XOR2_X1 U48 ( .A(B[12]), .B(A[12]), .Z(n34) );
  XOR2_X1 U49 ( .A(n21), .B(n34), .Z(SUM[12]) );
  NAND2_X1 U50 ( .A1(n32), .A2(B[12]), .ZN(n35) );
  NAND2_X1 U51 ( .A1(carry[12]), .A2(A[12]), .ZN(n36) );
  NAND2_X1 U52 ( .A1(B[12]), .A2(A[12]), .ZN(n37) );
  NAND3_X1 U53 ( .A1(n35), .A2(n36), .A3(n37), .ZN(carry[13]) );
  XOR2_X1 U54 ( .A(B[7]), .B(A[7]), .Z(n38) );
  XOR2_X1 U55 ( .A(carry[7]), .B(n38), .Z(SUM[7]) );
  NAND2_X1 U56 ( .A1(n26), .A2(B[7]), .ZN(n39) );
  NAND2_X1 U57 ( .A1(n26), .A2(A[7]), .ZN(n40) );
  NAND2_X1 U58 ( .A1(B[7]), .A2(A[7]), .ZN(n41) );
  NAND3_X1 U59 ( .A1(n39), .A2(n8), .A3(n41), .ZN(carry[8]) );
  CLKBUF_X1 U60 ( .A(n27), .Z(n42) );
  NAND3_X1 U61 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n43) );
  NAND3_X1 U62 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n44) );
  XOR2_X1 U63 ( .A(B[10]), .B(A[10]), .Z(n45) );
  XOR2_X1 U64 ( .A(n44), .B(n45), .Z(SUM[10]) );
  NAND2_X1 U65 ( .A1(n43), .A2(B[10]), .ZN(n46) );
  NAND2_X1 U66 ( .A1(carry[10]), .A2(A[10]), .ZN(n47) );
  NAND2_X1 U67 ( .A1(B[10]), .A2(A[10]), .ZN(n48) );
  NAND3_X1 U68 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[11]) );
  XOR2_X1 U69 ( .A(B[11]), .B(A[11]), .Z(n49) );
  XOR2_X1 U70 ( .A(n42), .B(n49), .Z(SUM[11]) );
  NAND2_X1 U71 ( .A1(n27), .A2(B[11]), .ZN(n50) );
  NAND2_X1 U72 ( .A1(carry[11]), .A2(A[11]), .ZN(n51) );
  NAND2_X1 U73 ( .A1(B[11]), .A2(A[11]), .ZN(n52) );
  NAND3_X1 U74 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[12]) );
  NAND3_X1 U75 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n53) );
  NAND3_X1 U76 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n54) );
  NAND3_X1 U77 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n55) );
  NAND3_X1 U78 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n56) );
  XOR2_X1 U79 ( .A(B[8]), .B(A[8]), .Z(n57) );
  XOR2_X1 U80 ( .A(carry[8]), .B(n57), .Z(SUM[8]) );
  NAND2_X1 U81 ( .A1(n3), .A2(B[8]), .ZN(n58) );
  NAND2_X1 U82 ( .A1(n33), .A2(A[8]), .ZN(n59) );
  NAND2_X1 U83 ( .A1(B[8]), .A2(A[8]), .ZN(n60) );
  NAND3_X1 U84 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[9]) );
  XOR2_X1 U85 ( .A(B[9]), .B(A[9]), .Z(n61) );
  XOR2_X1 U86 ( .A(n56), .B(n61), .Z(SUM[9]) );
  NAND2_X1 U87 ( .A1(n55), .A2(B[9]), .ZN(n62) );
  NAND2_X1 U88 ( .A1(carry[9]), .A2(A[9]), .ZN(n63) );
  NAND2_X1 U89 ( .A1(B[9]), .A2(A[9]), .ZN(n64) );
  NAND3_X1 U90 ( .A1(n62), .A2(n63), .A3(n64), .ZN(carry[10]) );
  XOR2_X1 U91 ( .A(B[1]), .B(A[1]), .Z(n65) );
  XOR2_X1 U92 ( .A(n73), .B(n65), .Z(SUM[1]) );
  NAND2_X1 U93 ( .A1(n73), .A2(B[1]), .ZN(n66) );
  NAND2_X1 U94 ( .A1(n73), .A2(A[1]), .ZN(n67) );
  NAND2_X1 U95 ( .A1(B[1]), .A2(A[1]), .ZN(n68) );
  NAND3_X1 U96 ( .A1(n66), .A2(n67), .A3(n68), .ZN(carry[2]) );
  XOR2_X1 U97 ( .A(B[2]), .B(A[2]), .Z(n69) );
  XOR2_X1 U98 ( .A(n54), .B(n69), .Z(SUM[2]) );
  NAND2_X1 U99 ( .A1(n53), .A2(B[2]), .ZN(n70) );
  NAND2_X1 U100 ( .A1(carry[2]), .A2(A[2]), .ZN(n71) );
  NAND2_X1 U101 ( .A1(B[2]), .A2(A[2]), .ZN(n72) );
  NAND3_X1 U102 ( .A1(n70), .A2(n71), .A3(n72), .ZN(carry[3]) );
  XOR2_X1 U103 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_5_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n317), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n316), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n320), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n319), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n322), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  NAND2_X1 U157 ( .A1(n339), .A2(n368), .ZN(n341) );
  CLKBUF_X1 U158 ( .A(n265), .Z(n206) );
  NAND2_X1 U159 ( .A1(n8), .A2(n39), .ZN(n207) );
  CLKBUF_X1 U160 ( .A(n230), .Z(n208) );
  CLKBUF_X1 U161 ( .A(b[1]), .Z(n209) );
  CLKBUF_X1 U162 ( .A(n252), .Z(n210) );
  XNOR2_X1 U163 ( .A(n209), .B(n222), .ZN(n211) );
  AND2_X1 U164 ( .A1(n262), .A2(n102), .ZN(n212) );
  INV_X1 U165 ( .A(n311), .ZN(n213) );
  CLKBUF_X1 U166 ( .A(n284), .Z(n214) );
  NAND2_X2 U167 ( .A1(n246), .A2(n247), .ZN(n215) );
  NAND2_X1 U168 ( .A1(n246), .A2(n247), .ZN(n339) );
  NAND3_X1 U169 ( .A1(n284), .A2(n285), .A3(n286), .ZN(n216) );
  NAND3_X1 U170 ( .A1(n257), .A2(n207), .A3(n259), .ZN(n217) );
  NAND2_X1 U171 ( .A1(n253), .A2(n20), .ZN(n218) );
  NAND3_X1 U172 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n219) );
  CLKBUF_X1 U173 ( .A(n309), .Z(n220) );
  CLKBUF_X1 U174 ( .A(b[1]), .Z(n221) );
  BUF_X2 U175 ( .A(a[1]), .Z(n222) );
  NAND3_X1 U176 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n223) );
  NAND3_X1 U177 ( .A1(n229), .A2(n208), .A3(n231), .ZN(n224) );
  CLKBUF_X1 U178 ( .A(b[1]), .Z(n289) );
  CLKBUF_X1 U179 ( .A(n56), .Z(n225) );
  XNOR2_X1 U180 ( .A(a[6]), .B(a[5]), .ZN(n350) );
  XNOR2_X1 U181 ( .A(a[6]), .B(a[5]), .ZN(n226) );
  NAND3_X1 U182 ( .A1(n268), .A2(n269), .A3(n270), .ZN(n227) );
  XOR2_X1 U183 ( .A(n103), .B(n96), .Z(n228) );
  XOR2_X1 U184 ( .A(n14), .B(n228), .Z(product[2]) );
  NAND2_X1 U185 ( .A1(n14), .A2(n103), .ZN(n229) );
  NAND2_X1 U186 ( .A1(n14), .A2(n96), .ZN(n230) );
  NAND2_X1 U187 ( .A1(n103), .A2(n96), .ZN(n231) );
  NAND3_X1 U188 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n13) );
  CLKBUF_X1 U189 ( .A(n207), .Z(n232) );
  NAND3_X1 U190 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n233) );
  NAND3_X1 U191 ( .A1(n264), .A2(n206), .A3(n266), .ZN(n234) );
  NAND2_X1 U192 ( .A1(n280), .A2(n19), .ZN(n235) );
  XOR2_X1 U193 ( .A(n50), .B(n53), .Z(n236) );
  XOR2_X1 U194 ( .A(n234), .B(n236), .Z(product[5]) );
  NAND2_X1 U195 ( .A1(n233), .A2(n50), .ZN(n237) );
  NAND2_X1 U196 ( .A1(n11), .A2(n53), .ZN(n238) );
  NAND2_X1 U197 ( .A1(n50), .A2(n53), .ZN(n239) );
  NAND3_X1 U198 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n10) );
  NAND3_X1 U199 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n240) );
  NAND3_X1 U200 ( .A1(n250), .A2(n251), .A3(n210), .ZN(n241) );
  NAND3_X1 U201 ( .A1(n220), .A2(n235), .A3(n310), .ZN(n242) );
  CLKBUF_X1 U202 ( .A(n218), .Z(n243) );
  NAND2_X1 U203 ( .A1(a[4]), .A2(a[3]), .ZN(n246) );
  NAND2_X1 U204 ( .A1(n244), .A2(n245), .ZN(n247) );
  INV_X1 U205 ( .A(a[4]), .ZN(n244) );
  INV_X1 U206 ( .A(a[3]), .ZN(n245) );
  NAND3_X1 U207 ( .A1(n273), .A2(n272), .A3(n274), .ZN(n248) );
  XOR2_X1 U208 ( .A(n224), .B(n71), .Z(n249) );
  XOR2_X1 U209 ( .A(n225), .B(n249), .Z(product[3]) );
  NAND2_X1 U210 ( .A1(n56), .A2(n223), .ZN(n250) );
  NAND2_X1 U211 ( .A1(n56), .A2(n71), .ZN(n251) );
  NAND2_X1 U212 ( .A1(n13), .A2(n71), .ZN(n252) );
  NAND3_X1 U213 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n12) );
  CLKBUF_X1 U214 ( .A(n95), .Z(n262) );
  NAND3_X1 U215 ( .A1(n277), .A2(n278), .A3(n279), .ZN(n253) );
  NAND3_X1 U216 ( .A1(n214), .A2(n285), .A3(n286), .ZN(n254) );
  NAND3_X1 U217 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n255) );
  XOR2_X1 U218 ( .A(n34), .B(n39), .Z(n256) );
  XOR2_X1 U219 ( .A(n254), .B(n256), .Z(product[8]) );
  NAND2_X1 U220 ( .A1(n216), .A2(n34), .ZN(n257) );
  NAND2_X1 U221 ( .A1(n8), .A2(n39), .ZN(n258) );
  NAND2_X1 U222 ( .A1(n34), .A2(n39), .ZN(n259) );
  NAND3_X1 U223 ( .A1(n257), .A2(n232), .A3(n259), .ZN(n7) );
  CLKBUF_X1 U224 ( .A(n227), .Z(n260) );
  CLKBUF_X1 U225 ( .A(n6), .Z(n261) );
  XOR2_X1 U226 ( .A(n102), .B(n95), .Z(n56) );
  XOR2_X1 U227 ( .A(n54), .B(n212), .Z(n263) );
  XOR2_X1 U228 ( .A(n241), .B(n263), .Z(product[4]) );
  NAND2_X1 U229 ( .A1(n240), .A2(n54), .ZN(n264) );
  NAND2_X1 U230 ( .A1(n12), .A2(n212), .ZN(n265) );
  NAND2_X1 U231 ( .A1(n54), .A2(n212), .ZN(n266) );
  NAND3_X1 U232 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n11) );
  XOR2_X1 U233 ( .A(n46), .B(n49), .Z(n267) );
  XOR2_X1 U234 ( .A(n10), .B(n267), .Z(product[6]) );
  NAND2_X1 U235 ( .A1(n219), .A2(n46), .ZN(n268) );
  NAND2_X1 U236 ( .A1(n219), .A2(n49), .ZN(n269) );
  NAND2_X1 U237 ( .A1(n46), .A2(n49), .ZN(n270) );
  NAND3_X1 U238 ( .A1(n268), .A2(n269), .A3(n270), .ZN(n9) );
  XOR2_X1 U239 ( .A(n33), .B(n28), .Z(n271) );
  XOR2_X1 U240 ( .A(n7), .B(n271), .Z(product[9]) );
  NAND2_X1 U241 ( .A1(n217), .A2(n33), .ZN(n272) );
  NAND2_X1 U242 ( .A1(n255), .A2(n28), .ZN(n273) );
  NAND2_X1 U243 ( .A1(n33), .A2(n28), .ZN(n274) );
  NAND3_X1 U244 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n6) );
  CLKBUF_X1 U245 ( .A(n253), .Z(n275) );
  XOR2_X1 U246 ( .A(n27), .B(n24), .Z(n276) );
  XOR2_X1 U247 ( .A(n261), .B(n276), .Z(product[10]) );
  NAND2_X1 U248 ( .A1(n6), .A2(n27), .ZN(n277) );
  NAND2_X1 U249 ( .A1(n248), .A2(n24), .ZN(n278) );
  NAND2_X1 U250 ( .A1(n27), .A2(n24), .ZN(n279) );
  NAND3_X1 U251 ( .A1(n277), .A2(n278), .A3(n279), .ZN(n5) );
  NAND3_X1 U252 ( .A1(n291), .A2(n292), .A3(n293), .ZN(n280) );
  NAND3_X1 U253 ( .A1(n243), .A2(n292), .A3(n293), .ZN(n281) );
  NAND3_X1 U254 ( .A1(n296), .A2(n295), .A3(n297), .ZN(n282) );
  INV_X2 U255 ( .A(n312), .ZN(n311) );
  XOR2_X1 U256 ( .A(n40), .B(n45), .Z(n283) );
  XOR2_X1 U257 ( .A(n260), .B(n283), .Z(product[7]) );
  NAND2_X1 U258 ( .A1(n227), .A2(n40), .ZN(n284) );
  NAND2_X1 U259 ( .A1(n9), .A2(n45), .ZN(n285) );
  NAND2_X1 U260 ( .A1(n40), .A2(n45), .ZN(n286) );
  NAND3_X1 U261 ( .A1(n284), .A2(n285), .A3(n286), .ZN(n8) );
  NAND3_X1 U262 ( .A1(n309), .A2(n308), .A3(n310), .ZN(n287) );
  NAND3_X1 U263 ( .A1(n235), .A2(n309), .A3(n310), .ZN(n288) );
  XOR2_X1 U264 ( .A(n20), .B(n23), .Z(n290) );
  XOR2_X1 U265 ( .A(n275), .B(n290), .Z(product[11]) );
  NAND2_X1 U266 ( .A1(n253), .A2(n20), .ZN(n291) );
  NAND2_X1 U267 ( .A1(n5), .A2(n23), .ZN(n292) );
  NAND2_X1 U268 ( .A1(n20), .A2(n23), .ZN(n293) );
  NAND3_X1 U269 ( .A1(n218), .A2(n292), .A3(n293), .ZN(n4) );
  XOR2_X1 U270 ( .A(n313), .B(n17), .Z(n294) );
  XOR2_X1 U271 ( .A(n242), .B(n294), .Z(product[13]) );
  NAND2_X1 U272 ( .A1(n287), .A2(n313), .ZN(n295) );
  NAND2_X1 U273 ( .A1(n288), .A2(n17), .ZN(n296) );
  NAND2_X1 U274 ( .A1(n313), .A2(n17), .ZN(n297) );
  NAND3_X1 U275 ( .A1(n295), .A2(n296), .A3(n297), .ZN(n2) );
  NAND2_X1 U276 ( .A1(a[2]), .A2(a[1]), .ZN(n300) );
  NAND2_X1 U277 ( .A1(n298), .A2(n299), .ZN(n301) );
  NAND2_X2 U278 ( .A1(n300), .A2(n301), .ZN(n329) );
  INV_X1 U279 ( .A(a[2]), .ZN(n298) );
  INV_X1 U280 ( .A(a[1]), .ZN(n299) );
  NAND2_X2 U281 ( .A1(n367), .A2(n329), .ZN(n331) );
  INV_X1 U282 ( .A(n15), .ZN(n313) );
  XNOR2_X1 U283 ( .A(n281), .B(n302), .ZN(product[12]) );
  XNOR2_X1 U284 ( .A(n19), .B(n18), .ZN(n302) );
  XNOR2_X1 U285 ( .A(n2), .B(n303), .ZN(product[14]) );
  XNOR2_X1 U286 ( .A(n314), .B(n15), .ZN(n303) );
  AND3_X1 U287 ( .A1(n306), .A2(n305), .A3(n307), .ZN(product[15]) );
  OAI22_X1 U288 ( .A1(n358), .A2(n352), .B1(n226), .B2(n360), .ZN(n15) );
  INV_X1 U289 ( .A(n337), .ZN(n320) );
  INV_X1 U290 ( .A(n348), .ZN(n317) );
  INV_X1 U291 ( .A(n21), .ZN(n316) );
  INV_X1 U292 ( .A(n328), .ZN(n322) );
  INV_X1 U293 ( .A(n31), .ZN(n319) );
  INV_X1 U294 ( .A(a[0]), .ZN(n323) );
  INV_X1 U295 ( .A(a[5]), .ZN(n318) );
  INV_X1 U296 ( .A(a[7]), .ZN(n315) );
  INV_X1 U297 ( .A(b[0]), .ZN(n312) );
  NAND2_X1 U298 ( .A1(n282), .A2(n314), .ZN(n305) );
  NAND2_X1 U299 ( .A1(n282), .A2(n15), .ZN(n306) );
  NAND2_X1 U300 ( .A1(n314), .A2(n15), .ZN(n307) );
  NAND2_X1 U301 ( .A1(n280), .A2(n19), .ZN(n308) );
  NAND2_X1 U302 ( .A1(n4), .A2(n18), .ZN(n309) );
  NAND2_X1 U303 ( .A1(n19), .A2(n18), .ZN(n310) );
  INV_X1 U304 ( .A(n359), .ZN(n314) );
  INV_X1 U305 ( .A(a[3]), .ZN(n321) );
  NOR2_X1 U306 ( .A1(n323), .A2(n213), .ZN(product[0]) );
  OAI22_X1 U307 ( .A1(n324), .A2(n325), .B1(n326), .B2(n323), .ZN(n99) );
  OAI22_X1 U308 ( .A1(n326), .A2(n325), .B1(n327), .B2(n323), .ZN(n98) );
  XNOR2_X1 U309 ( .A(b[6]), .B(n222), .ZN(n326) );
  OAI22_X1 U310 ( .A1(n323), .A2(n327), .B1(n325), .B2(n327), .ZN(n328) );
  XNOR2_X1 U311 ( .A(b[7]), .B(n222), .ZN(n327) );
  NOR2_X1 U312 ( .A1(n329), .A2(n312), .ZN(n96) );
  OAI22_X1 U313 ( .A1(n330), .A2(n331), .B1(n329), .B2(n332), .ZN(n95) );
  XNOR2_X1 U314 ( .A(a[3]), .B(n311), .ZN(n330) );
  OAI22_X1 U315 ( .A1(n331), .A2(n332), .B1(n329), .B2(n333), .ZN(n94) );
  XNOR2_X1 U316 ( .A(n221), .B(a[3]), .ZN(n332) );
  OAI22_X1 U317 ( .A1(n333), .A2(n331), .B1(n329), .B2(n334), .ZN(n93) );
  XNOR2_X1 U318 ( .A(b[2]), .B(a[3]), .ZN(n333) );
  OAI22_X1 U319 ( .A1(n334), .A2(n331), .B1(n329), .B2(n335), .ZN(n92) );
  XNOR2_X1 U320 ( .A(b[3]), .B(a[3]), .ZN(n334) );
  OAI22_X1 U321 ( .A1(n335), .A2(n331), .B1(n329), .B2(n336), .ZN(n91) );
  XNOR2_X1 U322 ( .A(b[4]), .B(a[3]), .ZN(n335) );
  OAI22_X1 U323 ( .A1(n338), .A2(n329), .B1(n331), .B2(n338), .ZN(n337) );
  NOR2_X1 U324 ( .A1(n215), .A2(n213), .ZN(n88) );
  OAI22_X1 U325 ( .A1(n340), .A2(n341), .B1(n215), .B2(n342), .ZN(n87) );
  XNOR2_X1 U326 ( .A(a[5]), .B(n311), .ZN(n340) );
  OAI22_X1 U327 ( .A1(n342), .A2(n341), .B1(n215), .B2(n343), .ZN(n86) );
  XNOR2_X1 U328 ( .A(n289), .B(a[5]), .ZN(n342) );
  OAI22_X1 U329 ( .A1(n343), .A2(n341), .B1(n215), .B2(n344), .ZN(n85) );
  XNOR2_X1 U330 ( .A(b[2]), .B(a[5]), .ZN(n343) );
  OAI22_X1 U331 ( .A1(n344), .A2(n341), .B1(n215), .B2(n345), .ZN(n84) );
  XNOR2_X1 U332 ( .A(b[3]), .B(a[5]), .ZN(n344) );
  OAI22_X1 U333 ( .A1(n345), .A2(n341), .B1(n215), .B2(n346), .ZN(n83) );
  XNOR2_X1 U334 ( .A(b[4]), .B(a[5]), .ZN(n345) );
  OAI22_X1 U335 ( .A1(n346), .A2(n341), .B1(n215), .B2(n347), .ZN(n82) );
  XNOR2_X1 U336 ( .A(b[5]), .B(a[5]), .ZN(n346) );
  OAI22_X1 U337 ( .A1(n349), .A2(n215), .B1(n341), .B2(n349), .ZN(n348) );
  NOR2_X1 U338 ( .A1(n350), .A2(n213), .ZN(n80) );
  OAI22_X1 U339 ( .A1(n351), .A2(n352), .B1(n226), .B2(n353), .ZN(n79) );
  XNOR2_X1 U340 ( .A(a[7]), .B(n311), .ZN(n351) );
  OAI22_X1 U341 ( .A1(n354), .A2(n352), .B1(n226), .B2(n355), .ZN(n77) );
  OAI22_X1 U342 ( .A1(n355), .A2(n352), .B1(n226), .B2(n356), .ZN(n76) );
  XNOR2_X1 U343 ( .A(b[3]), .B(a[7]), .ZN(n355) );
  OAI22_X1 U344 ( .A1(n356), .A2(n352), .B1(n226), .B2(n357), .ZN(n75) );
  XNOR2_X1 U345 ( .A(b[4]), .B(a[7]), .ZN(n356) );
  OAI22_X1 U346 ( .A1(n357), .A2(n352), .B1(n226), .B2(n358), .ZN(n74) );
  XNOR2_X1 U347 ( .A(b[5]), .B(a[7]), .ZN(n357) );
  OAI22_X1 U348 ( .A1(n360), .A2(n226), .B1(n352), .B2(n360), .ZN(n359) );
  OAI21_X1 U349 ( .B1(n311), .B2(n299), .A(n325), .ZN(n72) );
  OAI21_X1 U350 ( .B1(n321), .B2(n331), .A(n361), .ZN(n71) );
  OR3_X1 U351 ( .A1(n329), .A2(n311), .A3(n321), .ZN(n361) );
  OAI21_X1 U352 ( .B1(n318), .B2(n341), .A(n362), .ZN(n70) );
  OR3_X1 U353 ( .A1(n339), .A2(n311), .A3(n318), .ZN(n362) );
  OAI21_X1 U354 ( .B1(n315), .B2(n352), .A(n363), .ZN(n69) );
  OR3_X1 U355 ( .A1(n226), .A2(n311), .A3(n315), .ZN(n363) );
  XNOR2_X1 U356 ( .A(n364), .B(n365), .ZN(n38) );
  OR2_X1 U357 ( .A1(n364), .A2(n365), .ZN(n37) );
  OAI22_X1 U358 ( .A1(n336), .A2(n331), .B1(n329), .B2(n366), .ZN(n365) );
  XNOR2_X1 U359 ( .A(b[5]), .B(a[3]), .ZN(n336) );
  OAI22_X1 U360 ( .A1(n353), .A2(n352), .B1(n226), .B2(n354), .ZN(n364) );
  XNOR2_X1 U361 ( .A(b[2]), .B(a[7]), .ZN(n354) );
  XNOR2_X1 U362 ( .A(n289), .B(a[7]), .ZN(n353) );
  OAI22_X1 U363 ( .A1(n366), .A2(n331), .B1(n329), .B2(n338), .ZN(n31) );
  XNOR2_X1 U364 ( .A(b[7]), .B(a[3]), .ZN(n338) );
  XNOR2_X1 U365 ( .A(n321), .B(a[2]), .ZN(n367) );
  XNOR2_X1 U366 ( .A(b[6]), .B(a[3]), .ZN(n366) );
  OAI22_X1 U367 ( .A1(n347), .A2(n341), .B1(n215), .B2(n349), .ZN(n21) );
  XNOR2_X1 U368 ( .A(b[7]), .B(a[5]), .ZN(n349) );
  XNOR2_X1 U369 ( .A(n318), .B(a[4]), .ZN(n368) );
  XNOR2_X1 U370 ( .A(b[6]), .B(a[5]), .ZN(n347) );
  XNOR2_X1 U371 ( .A(b[7]), .B(a[7]), .ZN(n360) );
  NAND2_X1 U372 ( .A1(n350), .A2(n369), .ZN(n352) );
  XNOR2_X1 U373 ( .A(n315), .B(a[6]), .ZN(n369) );
  XNOR2_X1 U374 ( .A(b[6]), .B(a[7]), .ZN(n358) );
  OAI22_X1 U375 ( .A1(n311), .A2(n325), .B1(n370), .B2(n323), .ZN(n104) );
  OAI22_X1 U376 ( .A1(n211), .A2(n325), .B1(n371), .B2(n323), .ZN(n103) );
  XNOR2_X1 U377 ( .A(b[1]), .B(n222), .ZN(n370) );
  OAI22_X1 U378 ( .A1(n371), .A2(n325), .B1(n372), .B2(n323), .ZN(n102) );
  XNOR2_X1 U379 ( .A(b[2]), .B(n222), .ZN(n371) );
  OAI22_X1 U380 ( .A1(n372), .A2(n325), .B1(n373), .B2(n323), .ZN(n101) );
  XNOR2_X1 U381 ( .A(b[3]), .B(n222), .ZN(n372) );
  OAI22_X1 U382 ( .A1(n373), .A2(n325), .B1(n324), .B2(n323), .ZN(n100) );
  XNOR2_X1 U383 ( .A(b[5]), .B(n222), .ZN(n324) );
  NAND2_X1 U384 ( .A1(n222), .A2(n323), .ZN(n325) );
  XNOR2_X1 U385 ( .A(b[4]), .B(n222), .ZN(n373) );
endmodule


module mac_5 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_5_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_5_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_4_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83;
  wire   [15:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .S(SUM[15]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n83) );
  NAND3_X1 U2 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n1) );
  NAND3_X1 U3 ( .A1(n10), .A2(n11), .A3(n12), .ZN(n2) );
  NAND3_X1 U4 ( .A1(n72), .A2(n73), .A3(n74), .ZN(n3) );
  NAND3_X1 U5 ( .A1(n72), .A2(n73), .A3(n74), .ZN(n4) );
  NAND3_X1 U6 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n5) );
  NAND3_X1 U7 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n6) );
  CLKBUF_X1 U8 ( .A(n2), .Z(n7) );
  CLKBUF_X1 U9 ( .A(carry[14]), .Z(n8) );
  XOR2_X1 U10 ( .A(B[10]), .B(A[10]), .Z(n9) );
  XOR2_X1 U11 ( .A(n4), .B(n9), .Z(SUM[10]) );
  NAND2_X1 U12 ( .A1(n3), .A2(B[10]), .ZN(n10) );
  NAND2_X1 U13 ( .A1(carry[10]), .A2(A[10]), .ZN(n11) );
  NAND2_X1 U14 ( .A1(B[10]), .A2(A[10]), .ZN(n12) );
  NAND3_X1 U15 ( .A1(n10), .A2(n11), .A3(n12), .ZN(carry[11]) );
  CLKBUF_X1 U16 ( .A(n1), .Z(n13) );
  NAND3_X1 U17 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n14) );
  NAND3_X1 U18 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n15) );
  NAND3_X1 U19 ( .A1(n20), .A2(n21), .A3(n22), .ZN(n16) );
  NAND3_X1 U20 ( .A1(n20), .A2(n21), .A3(n22), .ZN(n17) );
  NAND3_X1 U21 ( .A1(n68), .A2(n69), .A3(n70), .ZN(n18) );
  XOR2_X1 U22 ( .A(B[4]), .B(A[4]), .Z(n19) );
  XOR2_X1 U23 ( .A(n15), .B(n19), .Z(SUM[4]) );
  NAND2_X1 U24 ( .A1(n14), .A2(B[4]), .ZN(n20) );
  NAND2_X1 U25 ( .A1(carry[4]), .A2(A[4]), .ZN(n21) );
  NAND2_X1 U26 ( .A1(B[4]), .A2(A[4]), .ZN(n22) );
  NAND3_X1 U27 ( .A1(n20), .A2(n21), .A3(n22), .ZN(carry[5]) );
  CLKBUF_X1 U28 ( .A(carry[7]), .Z(n23) );
  NAND3_X1 U29 ( .A1(n80), .A2(n81), .A3(n82), .ZN(n24) );
  XOR2_X1 U30 ( .A(B[3]), .B(A[3]), .Z(n25) );
  XOR2_X1 U31 ( .A(n24), .B(n25), .Z(SUM[3]) );
  NAND2_X1 U32 ( .A1(n24), .A2(B[3]), .ZN(n26) );
  NAND2_X1 U33 ( .A1(carry[3]), .A2(A[3]), .ZN(n27) );
  NAND2_X1 U34 ( .A1(B[3]), .A2(A[3]), .ZN(n28) );
  NAND3_X1 U35 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[4]) );
  CLKBUF_X1 U36 ( .A(n40), .Z(n29) );
  CLKBUF_X1 U37 ( .A(n51), .Z(n30) );
  CLKBUF_X1 U38 ( .A(n77), .Z(n31) );
  XOR2_X1 U39 ( .A(B[11]), .B(A[11]), .Z(n32) );
  XOR2_X1 U40 ( .A(n7), .B(n32), .Z(SUM[11]) );
  NAND2_X1 U41 ( .A1(n2), .A2(B[11]), .ZN(n33) );
  NAND2_X1 U42 ( .A1(carry[11]), .A2(A[11]), .ZN(n34) );
  NAND2_X1 U43 ( .A1(B[11]), .A2(A[11]), .ZN(n35) );
  NAND3_X1 U44 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[12]) );
  XOR2_X1 U45 ( .A(B[5]), .B(A[5]), .Z(n36) );
  XOR2_X1 U46 ( .A(n17), .B(n36), .Z(SUM[5]) );
  NAND2_X1 U47 ( .A1(n16), .A2(B[5]), .ZN(n37) );
  NAND2_X1 U48 ( .A1(carry[5]), .A2(A[5]), .ZN(n38) );
  NAND2_X1 U49 ( .A1(B[5]), .A2(A[5]), .ZN(n39) );
  NAND3_X1 U50 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[6]) );
  NAND3_X1 U51 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n40) );
  NAND3_X1 U52 ( .A1(n48), .A2(n47), .A3(n49), .ZN(n41) );
  XOR2_X1 U53 ( .A(B[12]), .B(A[12]), .Z(n42) );
  XOR2_X1 U54 ( .A(n13), .B(n42), .Z(SUM[12]) );
  NAND2_X1 U55 ( .A1(n1), .A2(B[12]), .ZN(n43) );
  NAND2_X1 U56 ( .A1(carry[12]), .A2(A[12]), .ZN(n44) );
  NAND2_X1 U57 ( .A1(B[12]), .A2(A[12]), .ZN(n45) );
  NAND3_X1 U58 ( .A1(n44), .A2(n43), .A3(n45), .ZN(carry[13]) );
  XOR2_X1 U59 ( .A(B[6]), .B(A[6]), .Z(n46) );
  XOR2_X1 U60 ( .A(n6), .B(n46), .Z(SUM[6]) );
  NAND2_X1 U61 ( .A1(n5), .A2(B[6]), .ZN(n47) );
  NAND2_X1 U62 ( .A1(carry[6]), .A2(A[6]), .ZN(n48) );
  NAND2_X1 U63 ( .A1(B[6]), .A2(A[6]), .ZN(n49) );
  NAND3_X1 U64 ( .A1(n47), .A2(n48), .A3(n49), .ZN(carry[7]) );
  NAND3_X1 U65 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n50) );
  NAND3_X1 U66 ( .A1(n57), .A2(n58), .A3(n59), .ZN(n51) );
  XOR2_X1 U67 ( .A(B[13]), .B(A[13]), .Z(n52) );
  XOR2_X1 U68 ( .A(n29), .B(n52), .Z(SUM[13]) );
  NAND2_X1 U69 ( .A1(n40), .A2(B[13]), .ZN(n53) );
  NAND2_X1 U70 ( .A1(carry[13]), .A2(A[13]), .ZN(n54) );
  NAND2_X1 U71 ( .A1(B[13]), .A2(A[13]), .ZN(n55) );
  NAND3_X1 U72 ( .A1(n53), .A2(n54), .A3(n55), .ZN(carry[14]) );
  XOR2_X1 U73 ( .A(B[7]), .B(A[7]), .Z(n56) );
  XOR2_X1 U74 ( .A(n23), .B(n56), .Z(SUM[7]) );
  NAND2_X1 U75 ( .A1(n41), .A2(B[7]), .ZN(n57) );
  NAND2_X1 U76 ( .A1(carry[7]), .A2(A[7]), .ZN(n58) );
  NAND2_X1 U77 ( .A1(B[7]), .A2(A[7]), .ZN(n59) );
  NAND3_X1 U78 ( .A1(n57), .A2(n58), .A3(n59), .ZN(carry[8]) );
  NAND3_X1 U79 ( .A1(n77), .A2(n76), .A3(n78), .ZN(n60) );
  NAND3_X1 U80 ( .A1(n76), .A2(n31), .A3(n78), .ZN(n61) );
  XOR2_X1 U81 ( .A(B[14]), .B(A[14]), .Z(n62) );
  XOR2_X1 U82 ( .A(n8), .B(n62), .Z(SUM[14]) );
  NAND2_X1 U83 ( .A1(carry[14]), .A2(B[14]), .ZN(n63) );
  NAND2_X1 U84 ( .A1(n50), .A2(A[14]), .ZN(n64) );
  NAND2_X1 U85 ( .A1(B[14]), .A2(A[14]), .ZN(n65) );
  NAND3_X1 U86 ( .A1(n63), .A2(n64), .A3(n65), .ZN(carry[15]) );
  CLKBUF_X1 U87 ( .A(n18), .Z(n66) );
  XOR2_X1 U88 ( .A(B[8]), .B(A[8]), .Z(n67) );
  XOR2_X1 U89 ( .A(n30), .B(n67), .Z(SUM[8]) );
  NAND2_X1 U90 ( .A1(n51), .A2(B[8]), .ZN(n68) );
  NAND2_X1 U91 ( .A1(carry[8]), .A2(A[8]), .ZN(n69) );
  NAND2_X1 U92 ( .A1(B[8]), .A2(A[8]), .ZN(n70) );
  NAND3_X1 U93 ( .A1(n68), .A2(n69), .A3(n70), .ZN(carry[9]) );
  XOR2_X1 U94 ( .A(B[9]), .B(A[9]), .Z(n71) );
  XOR2_X1 U95 ( .A(n66), .B(n71), .Z(SUM[9]) );
  NAND2_X1 U96 ( .A1(n18), .A2(B[9]), .ZN(n72) );
  NAND2_X1 U97 ( .A1(carry[9]), .A2(A[9]), .ZN(n73) );
  NAND2_X1 U98 ( .A1(B[9]), .A2(A[9]), .ZN(n74) );
  NAND3_X1 U99 ( .A1(n72), .A2(n73), .A3(n74), .ZN(carry[10]) );
  XOR2_X1 U100 ( .A(B[1]), .B(A[1]), .Z(n75) );
  XOR2_X1 U101 ( .A(n83), .B(n75), .Z(SUM[1]) );
  NAND2_X1 U102 ( .A1(n83), .A2(B[1]), .ZN(n76) );
  NAND2_X1 U103 ( .A1(n83), .A2(A[1]), .ZN(n77) );
  NAND2_X1 U104 ( .A1(B[1]), .A2(A[1]), .ZN(n78) );
  NAND3_X1 U105 ( .A1(n76), .A2(n77), .A3(n78), .ZN(carry[2]) );
  XOR2_X1 U106 ( .A(B[2]), .B(A[2]), .Z(n79) );
  XOR2_X1 U107 ( .A(n61), .B(n79), .Z(SUM[2]) );
  NAND2_X1 U108 ( .A1(n60), .A2(B[2]), .ZN(n80) );
  NAND2_X1 U109 ( .A1(carry[2]), .A2(A[2]), .ZN(n81) );
  NAND2_X1 U110 ( .A1(B[2]), .A2(A[2]), .ZN(n82) );
  NAND3_X1 U111 ( .A1(n80), .A2(n81), .A3(n82), .ZN(carry[3]) );
  XOR2_X1 U112 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_4_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74,
         n75, n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92,
         n93, n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n311), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n310), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n314), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n313), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n316), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  CLKBUF_X1 U157 ( .A(n336), .Z(n206) );
  NAND2_X1 U158 ( .A1(n334), .A2(n363), .ZN(n336) );
  BUF_X1 U159 ( .A(n306), .Z(n268) );
  CLKBUF_X1 U160 ( .A(n365), .Z(n207) );
  CLKBUF_X1 U161 ( .A(a[1]), .Z(n208) );
  NAND3_X1 U162 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n209) );
  NAND2_X2 U163 ( .A1(n285), .A2(n286), .ZN(n210) );
  NAND2_X1 U164 ( .A1(n285), .A2(n286), .ZN(n334) );
  NAND3_X1 U165 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n211) );
  NAND3_X1 U166 ( .A1(n222), .A2(n221), .A3(n223), .ZN(n212) );
  CLKBUF_X1 U167 ( .A(n256), .Z(n213) );
  CLKBUF_X1 U168 ( .A(n56), .Z(n214) );
  NAND3_X1 U169 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n215) );
  NAND3_X1 U170 ( .A1(n213), .A2(n257), .A3(n258), .ZN(n216) );
  CLKBUF_X1 U171 ( .A(n212), .Z(n217) );
  CLKBUF_X1 U172 ( .A(n302), .Z(n218) );
  NAND2_X1 U173 ( .A1(n230), .A2(n19), .ZN(n219) );
  XOR2_X1 U174 ( .A(n46), .B(n49), .Z(n220) );
  XOR2_X1 U175 ( .A(n216), .B(n220), .Z(product[6]) );
  NAND2_X1 U176 ( .A1(n215), .A2(n46), .ZN(n221) );
  NAND2_X1 U177 ( .A1(n10), .A2(n49), .ZN(n222) );
  NAND2_X1 U178 ( .A1(n46), .A2(n49), .ZN(n223) );
  NAND3_X1 U179 ( .A1(n221), .A2(n222), .A3(n223), .ZN(n9) );
  CLKBUF_X1 U180 ( .A(n240), .Z(n224) );
  CLKBUF_X1 U181 ( .A(b[1]), .Z(n225) );
  XOR2_X2 U182 ( .A(a[6]), .B(n312), .Z(n345) );
  CLKBUF_X1 U183 ( .A(n272), .Z(n226) );
  NAND3_X1 U184 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n227) );
  NAND3_X1 U185 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n228) );
  CLKBUF_X1 U186 ( .A(n245), .Z(n229) );
  NAND3_X1 U187 ( .A1(n302), .A2(n303), .A3(n304), .ZN(n230) );
  NAND3_X1 U188 ( .A1(n278), .A2(n277), .A3(n276), .ZN(n231) );
  NAND3_X1 U189 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n232) );
  XNOR2_X1 U190 ( .A(n233), .B(n231), .ZN(product[14]) );
  XNOR2_X1 U191 ( .A(n308), .B(n15), .ZN(n233) );
  NAND3_X1 U192 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n234) );
  XOR2_X1 U193 ( .A(n40), .B(n45), .Z(n235) );
  XOR2_X1 U194 ( .A(n217), .B(n235), .Z(product[7]) );
  NAND2_X1 U195 ( .A1(n212), .A2(n40), .ZN(n236) );
  NAND2_X1 U196 ( .A1(n9), .A2(n45), .ZN(n237) );
  NAND2_X1 U197 ( .A1(n40), .A2(n45), .ZN(n238) );
  NAND3_X1 U198 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n8) );
  XOR2_X1 U199 ( .A(n214), .B(n71), .Z(n239) );
  XOR2_X1 U200 ( .A(n232), .B(n239), .Z(product[3]) );
  NAND2_X1 U201 ( .A1(n232), .A2(n56), .ZN(n240) );
  NAND2_X1 U202 ( .A1(n13), .A2(n71), .ZN(n241) );
  NAND2_X1 U203 ( .A1(n56), .A2(n71), .ZN(n242) );
  NAND3_X1 U204 ( .A1(n224), .A2(n241), .A3(n242), .ZN(n12) );
  NAND3_X1 U205 ( .A1(n226), .A2(n219), .A3(n274), .ZN(n243) );
  NAND3_X1 U206 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n244) );
  NAND3_X1 U207 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n245) );
  NAND3_X1 U208 ( .A1(n299), .A2(n298), .A3(n300), .ZN(n246) );
  XOR2_X1 U209 ( .A(n54), .B(n55), .Z(n247) );
  XOR2_X1 U210 ( .A(n12), .B(n247), .Z(product[4]) );
  NAND2_X1 U211 ( .A1(n209), .A2(n54), .ZN(n248) );
  NAND2_X1 U212 ( .A1(n227), .A2(n55), .ZN(n249) );
  NAND2_X1 U213 ( .A1(n54), .A2(n55), .ZN(n250) );
  NAND3_X1 U214 ( .A1(n249), .A2(n248), .A3(n250), .ZN(n11) );
  XOR2_X1 U215 ( .A(n34), .B(n39), .Z(n251) );
  XOR2_X1 U216 ( .A(n8), .B(n251), .Z(product[8]) );
  NAND2_X1 U217 ( .A1(n211), .A2(n34), .ZN(n252) );
  NAND2_X1 U218 ( .A1(n228), .A2(n39), .ZN(n253) );
  NAND2_X1 U219 ( .A1(n34), .A2(n39), .ZN(n254) );
  NAND3_X1 U220 ( .A1(n253), .A2(n252), .A3(n254), .ZN(n7) );
  XOR2_X1 U221 ( .A(n50), .B(n53), .Z(n255) );
  XOR2_X1 U222 ( .A(n244), .B(n255), .Z(product[5]) );
  NAND2_X1 U223 ( .A1(n244), .A2(n50), .ZN(n256) );
  NAND2_X1 U224 ( .A1(n11), .A2(n53), .ZN(n257) );
  NAND2_X1 U225 ( .A1(n50), .A2(n53), .ZN(n258) );
  NAND3_X1 U226 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n10) );
  CLKBUF_X1 U227 ( .A(n246), .Z(n259) );
  CLKBUF_X1 U228 ( .A(n6), .Z(n260) );
  XOR2_X1 U229 ( .A(n33), .B(n28), .Z(n261) );
  XOR2_X1 U230 ( .A(n229), .B(n261), .Z(product[9]) );
  NAND2_X1 U231 ( .A1(n245), .A2(n33), .ZN(n262) );
  NAND2_X1 U232 ( .A1(n7), .A2(n28), .ZN(n263) );
  NAND2_X1 U233 ( .A1(n33), .A2(n28), .ZN(n264) );
  NAND3_X1 U234 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n6) );
  NAND3_X1 U235 ( .A1(n278), .A2(n277), .A3(n276), .ZN(n265) );
  NAND3_X1 U236 ( .A1(n218), .A2(n303), .A3(n304), .ZN(n266) );
  NAND3_X1 U237 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n267) );
  AND3_X1 U238 ( .A1(n281), .A2(n280), .A3(n279), .ZN(product[15]) );
  AND2_X1 U239 ( .A1(n104), .A2(n72), .ZN(n270) );
  XOR2_X1 U240 ( .A(n18), .B(n19), .Z(n271) );
  XOR2_X1 U241 ( .A(n266), .B(n271), .Z(product[12]) );
  NAND2_X1 U242 ( .A1(n4), .A2(n18), .ZN(n272) );
  NAND2_X1 U243 ( .A1(n230), .A2(n19), .ZN(n273) );
  NAND2_X1 U244 ( .A1(n18), .A2(n19), .ZN(n274) );
  NAND3_X1 U245 ( .A1(n219), .A2(n272), .A3(n274), .ZN(n3) );
  NAND2_X2 U246 ( .A1(n324), .A2(n362), .ZN(n326) );
  XOR2_X1 U247 ( .A(n17), .B(n307), .Z(n275) );
  XOR2_X1 U248 ( .A(n275), .B(n243), .Z(product[13]) );
  NAND2_X1 U249 ( .A1(n17), .A2(n307), .ZN(n276) );
  NAND2_X1 U250 ( .A1(n17), .A2(n267), .ZN(n277) );
  NAND2_X1 U251 ( .A1(n307), .A2(n3), .ZN(n278) );
  NAND3_X1 U252 ( .A1(n278), .A2(n277), .A3(n276), .ZN(n2) );
  NAND2_X1 U253 ( .A1(n308), .A2(n15), .ZN(n279) );
  NAND2_X1 U254 ( .A1(n2), .A2(n308), .ZN(n280) );
  NAND2_X1 U255 ( .A1(n265), .A2(n15), .ZN(n281) );
  INV_X1 U256 ( .A(n306), .ZN(n282) );
  NAND2_X1 U257 ( .A1(a[4]), .A2(a[3]), .ZN(n285) );
  NAND2_X1 U258 ( .A1(n283), .A2(n284), .ZN(n286) );
  INV_X1 U259 ( .A(a[4]), .ZN(n283) );
  INV_X1 U260 ( .A(a[3]), .ZN(n284) );
  NAND2_X1 U261 ( .A1(n291), .A2(n292), .ZN(n287) );
  NAND2_X1 U262 ( .A1(n291), .A2(n292), .ZN(n288) );
  NAND2_X1 U263 ( .A1(n291), .A2(n292), .ZN(n324) );
  NAND2_X1 U264 ( .A1(a[2]), .A2(a[1]), .ZN(n291) );
  NAND2_X1 U265 ( .A1(n289), .A2(n290), .ZN(n292) );
  INV_X1 U266 ( .A(a[2]), .ZN(n289) );
  INV_X1 U267 ( .A(a[1]), .ZN(n290) );
  INV_X1 U268 ( .A(n15), .ZN(n307) );
  INV_X1 U269 ( .A(n21), .ZN(n310) );
  INV_X1 U270 ( .A(n343), .ZN(n311) );
  INV_X1 U271 ( .A(n323), .ZN(n316) );
  INV_X1 U272 ( .A(n332), .ZN(n314) );
  INV_X1 U273 ( .A(n31), .ZN(n313) );
  INV_X1 U274 ( .A(n354), .ZN(n308) );
  INV_X1 U275 ( .A(a[0]), .ZN(n318) );
  INV_X1 U276 ( .A(a[5]), .ZN(n312) );
  INV_X1 U277 ( .A(a[7]), .ZN(n309) );
  XOR2_X1 U278 ( .A(n103), .B(n96), .Z(n293) );
  XOR2_X1 U279 ( .A(n270), .B(n293), .Z(product[2]) );
  NAND2_X1 U280 ( .A1(n270), .A2(n103), .ZN(n294) );
  NAND2_X1 U281 ( .A1(n14), .A2(n96), .ZN(n295) );
  NAND2_X1 U282 ( .A1(n103), .A2(n96), .ZN(n296) );
  NAND3_X1 U283 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n13) );
  XOR2_X1 U284 ( .A(n27), .B(n24), .Z(n297) );
  XOR2_X1 U285 ( .A(n260), .B(n297), .Z(product[10]) );
  NAND2_X1 U286 ( .A1(n234), .A2(n27), .ZN(n298) );
  NAND2_X1 U287 ( .A1(n6), .A2(n24), .ZN(n299) );
  NAND2_X1 U288 ( .A1(n27), .A2(n24), .ZN(n300) );
  NAND3_X1 U289 ( .A1(n299), .A2(n298), .A3(n300), .ZN(n5) );
  XOR2_X1 U290 ( .A(n23), .B(n20), .Z(n301) );
  XOR2_X1 U291 ( .A(n259), .B(n301), .Z(product[11]) );
  NAND2_X1 U292 ( .A1(n246), .A2(n23), .ZN(n302) );
  NAND2_X1 U293 ( .A1(n5), .A2(n20), .ZN(n303) );
  NAND2_X1 U294 ( .A1(n23), .A2(n20), .ZN(n304) );
  NAND3_X1 U295 ( .A1(n302), .A2(n303), .A3(n304), .ZN(n4) );
  INV_X1 U296 ( .A(b[0]), .ZN(n306) );
  INV_X1 U297 ( .A(a[3]), .ZN(n315) );
  INV_X1 U298 ( .A(a[1]), .ZN(n317) );
  INV_X1 U299 ( .A(n306), .ZN(n305) );
  NOR2_X1 U300 ( .A1(n318), .A2(n268), .ZN(product[0]) );
  OAI22_X1 U301 ( .A1(n319), .A2(n320), .B1(n321), .B2(n318), .ZN(n99) );
  OAI22_X1 U302 ( .A1(n321), .A2(n320), .B1(n322), .B2(n318), .ZN(n98) );
  XNOR2_X1 U303 ( .A(b[6]), .B(n208), .ZN(n321) );
  OAI22_X1 U304 ( .A1(n318), .A2(n322), .B1(n320), .B2(n322), .ZN(n323) );
  XNOR2_X1 U305 ( .A(b[7]), .B(n208), .ZN(n322) );
  NOR2_X1 U306 ( .A1(n287), .A2(n268), .ZN(n96) );
  OAI22_X1 U307 ( .A1(n325), .A2(n326), .B1(n287), .B2(n327), .ZN(n95) );
  XNOR2_X1 U308 ( .A(a[3]), .B(n305), .ZN(n325) );
  OAI22_X1 U309 ( .A1(n327), .A2(n326), .B1(n288), .B2(n328), .ZN(n94) );
  XNOR2_X1 U310 ( .A(b[1]), .B(a[3]), .ZN(n327) );
  OAI22_X1 U311 ( .A1(n328), .A2(n326), .B1(n288), .B2(n329), .ZN(n93) );
  XNOR2_X1 U312 ( .A(b[2]), .B(a[3]), .ZN(n328) );
  OAI22_X1 U313 ( .A1(n329), .A2(n326), .B1(n287), .B2(n330), .ZN(n92) );
  XNOR2_X1 U314 ( .A(b[3]), .B(a[3]), .ZN(n329) );
  OAI22_X1 U315 ( .A1(n330), .A2(n326), .B1(n287), .B2(n331), .ZN(n91) );
  XNOR2_X1 U316 ( .A(b[4]), .B(a[3]), .ZN(n330) );
  OAI22_X1 U317 ( .A1(n333), .A2(n288), .B1(n326), .B2(n333), .ZN(n332) );
  NOR2_X1 U318 ( .A1(n210), .A2(n268), .ZN(n88) );
  OAI22_X1 U319 ( .A1(n335), .A2(n336), .B1(n210), .B2(n337), .ZN(n87) );
  XNOR2_X1 U320 ( .A(a[5]), .B(n282), .ZN(n335) );
  OAI22_X1 U321 ( .A1(n337), .A2(n336), .B1(n210), .B2(n338), .ZN(n86) );
  XNOR2_X1 U322 ( .A(b[1]), .B(a[5]), .ZN(n337) );
  OAI22_X1 U323 ( .A1(n338), .A2(n336), .B1(n210), .B2(n339), .ZN(n85) );
  XNOR2_X1 U324 ( .A(b[2]), .B(a[5]), .ZN(n338) );
  OAI22_X1 U325 ( .A1(n339), .A2(n336), .B1(n210), .B2(n340), .ZN(n84) );
  XNOR2_X1 U326 ( .A(b[3]), .B(a[5]), .ZN(n339) );
  OAI22_X1 U327 ( .A1(n340), .A2(n336), .B1(n210), .B2(n341), .ZN(n83) );
  XNOR2_X1 U328 ( .A(b[4]), .B(a[5]), .ZN(n340) );
  OAI22_X1 U329 ( .A1(n341), .A2(n336), .B1(n210), .B2(n342), .ZN(n82) );
  XNOR2_X1 U330 ( .A(b[5]), .B(a[5]), .ZN(n341) );
  OAI22_X1 U331 ( .A1(n344), .A2(n210), .B1(n206), .B2(n344), .ZN(n343) );
  NOR2_X1 U332 ( .A1(n345), .A2(n268), .ZN(n80) );
  OAI22_X1 U333 ( .A1(n346), .A2(n347), .B1(n345), .B2(n348), .ZN(n79) );
  XNOR2_X1 U334 ( .A(a[7]), .B(n282), .ZN(n346) );
  OAI22_X1 U335 ( .A1(n349), .A2(n347), .B1(n345), .B2(n350), .ZN(n77) );
  OAI22_X1 U336 ( .A1(n350), .A2(n347), .B1(n345), .B2(n351), .ZN(n76) );
  XNOR2_X1 U337 ( .A(b[3]), .B(a[7]), .ZN(n350) );
  OAI22_X1 U338 ( .A1(n351), .A2(n347), .B1(n345), .B2(n352), .ZN(n75) );
  XNOR2_X1 U339 ( .A(b[4]), .B(a[7]), .ZN(n351) );
  OAI22_X1 U340 ( .A1(n352), .A2(n347), .B1(n345), .B2(n353), .ZN(n74) );
  XNOR2_X1 U341 ( .A(b[5]), .B(a[7]), .ZN(n352) );
  OAI22_X1 U342 ( .A1(n355), .A2(n345), .B1(n347), .B2(n355), .ZN(n354) );
  OAI21_X1 U343 ( .B1(n305), .B2(n317), .A(n320), .ZN(n72) );
  OAI21_X1 U344 ( .B1(n315), .B2(n326), .A(n356), .ZN(n71) );
  OR3_X1 U345 ( .A1(n288), .A2(n282), .A3(n315), .ZN(n356) );
  OAI21_X1 U346 ( .B1(n312), .B2(n336), .A(n357), .ZN(n70) );
  OR3_X1 U347 ( .A1(n334), .A2(n305), .A3(n312), .ZN(n357) );
  OAI21_X1 U348 ( .B1(n309), .B2(n347), .A(n358), .ZN(n69) );
  OR3_X1 U349 ( .A1(n345), .A2(n282), .A3(n309), .ZN(n358) );
  XNOR2_X1 U350 ( .A(n359), .B(n360), .ZN(n38) );
  OR2_X1 U351 ( .A1(n359), .A2(n360), .ZN(n37) );
  OAI22_X1 U352 ( .A1(n331), .A2(n326), .B1(n288), .B2(n361), .ZN(n360) );
  XNOR2_X1 U353 ( .A(b[5]), .B(a[3]), .ZN(n331) );
  OAI22_X1 U354 ( .A1(n348), .A2(n347), .B1(n345), .B2(n349), .ZN(n359) );
  XNOR2_X1 U355 ( .A(b[2]), .B(a[7]), .ZN(n349) );
  XNOR2_X1 U356 ( .A(n225), .B(a[7]), .ZN(n348) );
  OAI22_X1 U357 ( .A1(n361), .A2(n326), .B1(n287), .B2(n333), .ZN(n31) );
  XNOR2_X1 U358 ( .A(b[7]), .B(a[3]), .ZN(n333) );
  XNOR2_X1 U359 ( .A(n315), .B(a[2]), .ZN(n362) );
  XNOR2_X1 U360 ( .A(b[6]), .B(a[3]), .ZN(n361) );
  OAI22_X1 U361 ( .A1(n342), .A2(n206), .B1(n210), .B2(n344), .ZN(n21) );
  XNOR2_X1 U362 ( .A(b[7]), .B(a[5]), .ZN(n344) );
  XNOR2_X1 U363 ( .A(n312), .B(a[4]), .ZN(n363) );
  XNOR2_X1 U364 ( .A(b[6]), .B(a[5]), .ZN(n342) );
  OAI22_X1 U365 ( .A1(n353), .A2(n347), .B1(n345), .B2(n355), .ZN(n15) );
  XNOR2_X1 U366 ( .A(b[7]), .B(a[7]), .ZN(n355) );
  NAND2_X1 U367 ( .A1(n345), .A2(n364), .ZN(n347) );
  XNOR2_X1 U368 ( .A(n309), .B(a[6]), .ZN(n364) );
  XNOR2_X1 U369 ( .A(b[6]), .B(a[7]), .ZN(n353) );
  OAI22_X1 U370 ( .A1(n305), .A2(n320), .B1(n365), .B2(n318), .ZN(n104) );
  OAI22_X1 U371 ( .A1(n207), .A2(n320), .B1(n366), .B2(n318), .ZN(n103) );
  XNOR2_X1 U372 ( .A(b[1]), .B(a[1]), .ZN(n365) );
  OAI22_X1 U373 ( .A1(n366), .A2(n320), .B1(n367), .B2(n318), .ZN(n102) );
  XNOR2_X1 U374 ( .A(b[2]), .B(a[1]), .ZN(n366) );
  OAI22_X1 U375 ( .A1(n320), .A2(n367), .B1(n368), .B2(n318), .ZN(n101) );
  XNOR2_X1 U376 ( .A(b[3]), .B(a[1]), .ZN(n367) );
  OAI22_X1 U377 ( .A1(n368), .A2(n320), .B1(n319), .B2(n318), .ZN(n100) );
  XNOR2_X1 U378 ( .A(b[5]), .B(n208), .ZN(n319) );
  NAND2_X1 U379 ( .A1(a[1]), .A2(n318), .ZN(n320) );
  XNOR2_X1 U380 ( .A(b[4]), .B(a[1]), .ZN(n368) );
endmodule


module mac_4 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   n6, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, n2, n4;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(n6), .QN(n2) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  mac_4_DW01_add_0 add_356 ( .A(pipeline), .B({mac_out[15:1], n6}), .CI(1'b0), 
        .SUM(sum) );
  mac_4_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n4), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n4), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n4), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n4), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n4), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n4), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n4), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n4), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n4), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n4), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n4), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n4), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n4), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n4), .ZN(N6) );
  INV_X1 U18 ( .A(n2), .ZN(mac_out[0]) );
  AND2_X1 U19 ( .A1(sum[0]), .A2(n4), .ZN(N3) );
  AND2_X1 U20 ( .A1(sum[15]), .A2(n4), .ZN(N18) );
  INV_X1 U21 ( .A(clear_acc), .ZN(n4) );
endmodule


module mac_3_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88;
  wire   [15:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .S(SUM[15]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  NAND2_X1 U1 ( .A1(n88), .A2(A[1]), .ZN(n1) );
  CLKBUF_X1 U2 ( .A(n11), .Z(n2) );
  CLKBUF_X1 U3 ( .A(n14), .Z(n3) );
  CLKBUF_X1 U4 ( .A(n42), .Z(n4) );
  CLKBUF_X1 U5 ( .A(n47), .Z(n5) );
  CLKBUF_X1 U6 ( .A(n59), .Z(n6) );
  CLKBUF_X1 U7 ( .A(carry[5]), .Z(n7) );
  NAND3_X1 U8 ( .A1(n73), .A2(n74), .A3(n75), .ZN(n8) );
  NAND3_X1 U9 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n9) );
  NAND3_X1 U10 ( .A1(n58), .A2(n6), .A3(n60), .ZN(n10) );
  NAND3_X1 U11 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n11) );
  NAND3_X1 U12 ( .A1(n69), .A2(n1), .A3(n71), .ZN(n12) );
  NAND3_X1 U13 ( .A1(n69), .A2(n1), .A3(n71), .ZN(n13) );
  NAND3_X1 U14 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n14) );
  NAND3_X1 U15 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n15) );
  CLKBUF_X1 U16 ( .A(n78), .Z(n16) );
  XOR2_X1 U17 ( .A(B[10]), .B(A[10]), .Z(n17) );
  XOR2_X1 U18 ( .A(n10), .B(n17), .Z(SUM[10]) );
  NAND2_X1 U19 ( .A1(n9), .A2(B[10]), .ZN(n18) );
  NAND2_X1 U20 ( .A1(carry[10]), .A2(A[10]), .ZN(n19) );
  NAND2_X1 U21 ( .A1(B[10]), .A2(A[10]), .ZN(n20) );
  NAND3_X1 U22 ( .A1(n18), .A2(n19), .A3(n20), .ZN(carry[11]) );
  XOR2_X1 U23 ( .A(B[2]), .B(A[2]), .Z(n21) );
  XOR2_X1 U24 ( .A(n13), .B(n21), .Z(SUM[2]) );
  NAND2_X1 U25 ( .A1(n12), .A2(B[2]), .ZN(n22) );
  NAND2_X1 U26 ( .A1(carry[2]), .A2(A[2]), .ZN(n23) );
  NAND2_X1 U27 ( .A1(B[2]), .A2(A[2]), .ZN(n24) );
  NAND3_X1 U28 ( .A1(n22), .A2(n23), .A3(n24), .ZN(carry[3]) );
  NAND3_X1 U29 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n25) );
  NAND3_X1 U30 ( .A1(n4), .A2(n43), .A3(n44), .ZN(n26) );
  NAND3_X1 U31 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n27) );
  NAND3_X1 U32 ( .A1(n46), .A2(n5), .A3(n48), .ZN(n28) );
  CLKBUF_X1 U33 ( .A(n74), .Z(n29) );
  CLKBUF_X1 U34 ( .A(n52), .Z(n30) );
  XOR2_X1 U35 ( .A(B[3]), .B(A[3]), .Z(n31) );
  XOR2_X1 U36 ( .A(n3), .B(n31), .Z(SUM[3]) );
  NAND2_X1 U37 ( .A1(n14), .A2(B[3]), .ZN(n32) );
  NAND2_X1 U38 ( .A1(carry[3]), .A2(A[3]), .ZN(n33) );
  NAND2_X1 U39 ( .A1(B[3]), .A2(A[3]), .ZN(n34) );
  NAND3_X1 U40 ( .A1(n32), .A2(n33), .A3(n34), .ZN(carry[4]) );
  NAND3_X1 U41 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n35) );
  AND2_X1 U42 ( .A1(B[0]), .A2(A[0]), .ZN(n36) );
  AND2_X1 U43 ( .A1(A[0]), .A2(B[0]), .ZN(n37) );
  AND2_X1 U44 ( .A1(B[0]), .A2(A[0]), .ZN(n88) );
  CLKBUF_X1 U45 ( .A(n65), .Z(n38) );
  CLKBUF_X1 U46 ( .A(A[0]), .Z(n39) );
  NAND3_X1 U47 ( .A1(n86), .A2(n85), .A3(n87), .ZN(n40) );
  XOR2_X1 U48 ( .A(B[11]), .B(A[11]), .Z(n41) );
  XOR2_X1 U49 ( .A(n2), .B(n41), .Z(SUM[11]) );
  NAND2_X1 U50 ( .A1(n11), .A2(B[11]), .ZN(n42) );
  NAND2_X1 U51 ( .A1(carry[11]), .A2(A[11]), .ZN(n43) );
  NAND2_X1 U52 ( .A1(B[11]), .A2(A[11]), .ZN(n44) );
  NAND3_X1 U53 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[12]) );
  XOR2_X1 U54 ( .A(B[5]), .B(A[5]), .Z(n45) );
  XOR2_X1 U55 ( .A(n7), .B(n45), .Z(SUM[5]) );
  NAND2_X1 U56 ( .A1(carry[5]), .A2(B[5]), .ZN(n46) );
  NAND2_X1 U57 ( .A1(carry[5]), .A2(A[5]), .ZN(n47) );
  NAND2_X1 U58 ( .A1(B[5]), .A2(A[5]), .ZN(n48) );
  NAND3_X1 U59 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[6]) );
  NAND3_X1 U60 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n49) );
  XOR2_X1 U61 ( .A(B[12]), .B(A[12]), .Z(n50) );
  XOR2_X1 U62 ( .A(n26), .B(n50), .Z(SUM[12]) );
  NAND2_X1 U63 ( .A1(n25), .A2(B[12]), .ZN(n51) );
  NAND2_X1 U64 ( .A1(carry[12]), .A2(A[12]), .ZN(n52) );
  NAND2_X1 U65 ( .A1(B[12]), .A2(A[12]), .ZN(n53) );
  NAND3_X1 U66 ( .A1(n51), .A2(n30), .A3(n53), .ZN(carry[13]) );
  NAND3_X1 U67 ( .A1(n77), .A2(n78), .A3(n79), .ZN(n54) );
  NAND3_X1 U68 ( .A1(n77), .A2(n16), .A3(n79), .ZN(n55) );
  NAND3_X1 U69 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n56) );
  XOR2_X1 U70 ( .A(B[9]), .B(A[9]), .Z(n57) );
  XOR2_X1 U71 ( .A(carry[9]), .B(n57), .Z(SUM[9]) );
  NAND2_X1 U72 ( .A1(n35), .A2(B[9]), .ZN(n58) );
  NAND2_X1 U73 ( .A1(n56), .A2(A[9]), .ZN(n59) );
  NAND2_X1 U74 ( .A1(B[9]), .A2(A[9]), .ZN(n60) );
  NAND3_X1 U75 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[10]) );
  NAND3_X1 U76 ( .A1(n73), .A2(n29), .A3(n75), .ZN(n61) );
  NAND3_X1 U77 ( .A1(n73), .A2(n74), .A3(n75), .ZN(n62) );
  CLKBUF_X1 U78 ( .A(n40), .Z(n63) );
  XOR2_X1 U79 ( .A(B[8]), .B(A[8]), .Z(n64) );
  XOR2_X1 U80 ( .A(n63), .B(n64), .Z(SUM[8]) );
  NAND2_X1 U81 ( .A1(n40), .A2(B[8]), .ZN(n65) );
  NAND2_X1 U82 ( .A1(carry[8]), .A2(A[8]), .ZN(n66) );
  NAND2_X1 U83 ( .A1(B[8]), .A2(A[8]), .ZN(n67) );
  NAND3_X1 U84 ( .A1(n38), .A2(n66), .A3(n67), .ZN(carry[9]) );
  XOR2_X1 U85 ( .A(B[1]), .B(A[1]), .Z(n68) );
  XOR2_X1 U86 ( .A(n37), .B(n68), .Z(SUM[1]) );
  NAND2_X1 U87 ( .A1(n36), .A2(B[1]), .ZN(n69) );
  NAND2_X1 U88 ( .A1(n88), .A2(A[1]), .ZN(n70) );
  NAND2_X1 U89 ( .A1(B[1]), .A2(A[1]), .ZN(n71) );
  NAND3_X1 U90 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[2]) );
  XOR2_X1 U91 ( .A(B[13]), .B(A[13]), .Z(n72) );
  XOR2_X1 U92 ( .A(carry[13]), .B(n72), .Z(SUM[13]) );
  NAND2_X1 U93 ( .A1(n15), .A2(B[13]), .ZN(n73) );
  NAND2_X1 U94 ( .A1(n49), .A2(A[13]), .ZN(n74) );
  NAND2_X1 U95 ( .A1(B[13]), .A2(A[13]), .ZN(n75) );
  XOR2_X1 U96 ( .A(B[6]), .B(A[6]), .Z(n76) );
  XOR2_X1 U97 ( .A(n28), .B(n76), .Z(SUM[6]) );
  NAND2_X1 U98 ( .A1(n27), .A2(B[6]), .ZN(n77) );
  NAND2_X1 U99 ( .A1(carry[6]), .A2(A[6]), .ZN(n78) );
  NAND2_X1 U100 ( .A1(B[6]), .A2(A[6]), .ZN(n79) );
  NAND3_X1 U101 ( .A1(n77), .A2(n78), .A3(n79), .ZN(carry[7]) );
  XOR2_X1 U102 ( .A(B[14]), .B(A[14]), .Z(n80) );
  XOR2_X1 U103 ( .A(n61), .B(n80), .Z(SUM[14]) );
  NAND2_X1 U104 ( .A1(n8), .A2(B[14]), .ZN(n81) );
  NAND2_X1 U105 ( .A1(n62), .A2(A[14]), .ZN(n82) );
  NAND2_X1 U106 ( .A1(B[14]), .A2(A[14]), .ZN(n83) );
  NAND3_X1 U107 ( .A1(n81), .A2(n82), .A3(n83), .ZN(carry[15]) );
  XOR2_X1 U108 ( .A(B[7]), .B(A[7]), .Z(n84) );
  XOR2_X1 U109 ( .A(n55), .B(n84), .Z(SUM[7]) );
  NAND2_X1 U110 ( .A1(n54), .A2(B[7]), .ZN(n85) );
  NAND2_X1 U111 ( .A1(carry[7]), .A2(A[7]), .ZN(n86) );
  NAND2_X1 U112 ( .A1(B[7]), .A2(A[7]), .ZN(n87) );
  NAND3_X1 U113 ( .A1(n85), .A2(n86), .A3(n87), .ZN(carry[8]) );
  XOR2_X1 U114 ( .A(B[0]), .B(n39), .Z(SUM[0]) );
endmodule


module mac_3_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74,
         n75, n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92,
         n93, n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206,
         n207, n208, n209, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n303), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n302), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n306), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n305), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n308), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  CLKBUF_X1 U157 ( .A(n103), .Z(n206) );
  NAND2_X1 U158 ( .A1(n3), .A2(n17), .ZN(n207) );
  CLKBUF_X1 U159 ( .A(b[1]), .Z(n219) );
  NAND2_X1 U160 ( .A1(n227), .A2(n33), .ZN(n208) );
  CLKBUF_X1 U161 ( .A(n226), .Z(n209) );
  AND3_X1 U162 ( .A1(n250), .A2(n249), .A3(n248), .ZN(product[15]) );
  CLKBUF_X1 U163 ( .A(n208), .Z(n211) );
  NAND3_X1 U164 ( .A1(n290), .A2(n291), .A3(n292), .ZN(n212) );
  CLKBUF_X1 U165 ( .A(n281), .Z(n213) );
  NAND3_X1 U166 ( .A1(n208), .A2(n259), .A3(n260), .ZN(n214) );
  NAND3_X1 U167 ( .A1(n211), .A2(n259), .A3(n260), .ZN(n215) );
  XOR2_X1 U168 ( .A(a[3]), .B(n298), .Z(n317) );
  CLKBUF_X1 U169 ( .A(n269), .Z(n216) );
  AND2_X1 U170 ( .A1(n104), .A2(n72), .ZN(n217) );
  CLKBUF_X1 U171 ( .A(n227), .Z(n218) );
  XNOR2_X1 U172 ( .A(n220), .B(n243), .ZN(product[14]) );
  XNOR2_X1 U173 ( .A(n300), .B(n15), .ZN(n220) );
  CLKBUF_X1 U174 ( .A(n241), .Z(n221) );
  CLKBUF_X1 U175 ( .A(n270), .Z(n222) );
  NAND3_X1 U176 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n223) );
  CLKBUF_X1 U177 ( .A(n219), .Z(n224) );
  NAND3_X1 U178 ( .A1(n280), .A2(n213), .A3(n282), .ZN(n225) );
  NAND3_X1 U179 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n226) );
  NAND3_X1 U180 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n227) );
  NAND3_X1 U181 ( .A1(n281), .A2(n280), .A3(n282), .ZN(n228) );
  CLKBUF_X1 U182 ( .A(n56), .Z(n229) );
  BUF_X2 U183 ( .A(n316), .Z(n230) );
  XNOR2_X1 U184 ( .A(a[1]), .B(a[2]), .ZN(n316) );
  NAND3_X1 U185 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n231) );
  XOR2_X1 U186 ( .A(n34), .B(n39), .Z(n232) );
  XOR2_X1 U187 ( .A(n209), .B(n232), .Z(product[8]) );
  NAND2_X1 U188 ( .A1(n226), .A2(n34), .ZN(n233) );
  NAND2_X1 U189 ( .A1(n8), .A2(n39), .ZN(n234) );
  NAND2_X1 U190 ( .A1(n34), .A2(n39), .ZN(n235) );
  NAND3_X1 U191 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n7) );
  XOR2_X1 U192 ( .A(n206), .B(n96), .Z(n236) );
  XOR2_X1 U193 ( .A(n217), .B(n236), .Z(product[2]) );
  NAND2_X1 U194 ( .A1(n217), .A2(n103), .ZN(n237) );
  NAND2_X1 U195 ( .A1(n14), .A2(n96), .ZN(n238) );
  NAND2_X1 U196 ( .A1(n103), .A2(n96), .ZN(n239) );
  NAND3_X1 U197 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n13) );
  NAND3_X1 U198 ( .A1(n284), .A2(n285), .A3(n286), .ZN(n240) );
  NAND3_X1 U199 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n241) );
  NAND3_X1 U200 ( .A1(n207), .A2(n247), .A3(n245), .ZN(n242) );
  NAND3_X1 U201 ( .A1(n207), .A2(n245), .A3(n247), .ZN(n243) );
  XOR2_X1 U202 ( .A(n17), .B(n299), .Z(n244) );
  XOR2_X1 U203 ( .A(n244), .B(n225), .Z(product[13]) );
  NAND2_X1 U204 ( .A1(n17), .A2(n299), .ZN(n245) );
  NAND2_X1 U205 ( .A1(n3), .A2(n17), .ZN(n246) );
  NAND2_X1 U206 ( .A1(n299), .A2(n228), .ZN(n247) );
  NAND3_X1 U207 ( .A1(n247), .A2(n246), .A3(n245), .ZN(n2) );
  NAND2_X1 U208 ( .A1(n300), .A2(n15), .ZN(n248) );
  NAND2_X1 U209 ( .A1(n300), .A2(n2), .ZN(n249) );
  NAND2_X1 U210 ( .A1(n15), .A2(n242), .ZN(n250) );
  XOR2_X1 U211 ( .A(n93), .B(n100), .Z(n251) );
  XOR2_X1 U212 ( .A(n52), .B(n251), .Z(n50) );
  NAND2_X1 U213 ( .A1(n256), .A2(n93), .ZN(n252) );
  NAND2_X1 U214 ( .A1(n256), .A2(n100), .ZN(n253) );
  NAND2_X1 U215 ( .A1(n93), .A2(n100), .ZN(n254) );
  NAND3_X1 U216 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n49) );
  CLKBUF_X1 U217 ( .A(n4), .Z(n255) );
  XOR2_X1 U218 ( .A(n70), .B(n87), .Z(n256) );
  XOR2_X1 U219 ( .A(n33), .B(n28), .Z(n257) );
  XOR2_X1 U220 ( .A(n218), .B(n257), .Z(product[9]) );
  NAND2_X1 U221 ( .A1(n227), .A2(n33), .ZN(n258) );
  NAND2_X1 U222 ( .A1(n7), .A2(n28), .ZN(n259) );
  NAND2_X1 U223 ( .A1(n33), .A2(n28), .ZN(n260) );
  NAND3_X1 U224 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n6) );
  XOR2_X1 U225 ( .A(n23), .B(n20), .Z(n261) );
  XOR2_X1 U226 ( .A(n221), .B(n261), .Z(product[11]) );
  NAND2_X1 U227 ( .A1(n241), .A2(n23), .ZN(n262) );
  NAND2_X1 U228 ( .A1(n5), .A2(n20), .ZN(n263) );
  NAND2_X1 U229 ( .A1(n23), .A2(n20), .ZN(n264) );
  NAND3_X1 U230 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n4) );
  XOR2_X1 U231 ( .A(n27), .B(n24), .Z(n265) );
  XOR2_X1 U232 ( .A(n215), .B(n265), .Z(product[10]) );
  NAND2_X1 U233 ( .A1(n214), .A2(n27), .ZN(n266) );
  NAND2_X1 U234 ( .A1(n6), .A2(n24), .ZN(n267) );
  NAND2_X1 U235 ( .A1(n27), .A2(n24), .ZN(n268) );
  NAND3_X1 U236 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n5) );
  NAND3_X1 U237 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n269) );
  NAND3_X1 U238 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n270) );
  XOR2_X1 U239 ( .A(n46), .B(n49), .Z(n271) );
  XOR2_X1 U240 ( .A(n222), .B(n271), .Z(product[6]) );
  NAND2_X1 U241 ( .A1(n270), .A2(n46), .ZN(n272) );
  NAND2_X1 U242 ( .A1(n10), .A2(n49), .ZN(n273) );
  NAND2_X1 U243 ( .A1(n46), .A2(n49), .ZN(n274) );
  NAND3_X1 U244 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n9) );
  XOR2_X1 U245 ( .A(n40), .B(n45), .Z(n275) );
  XOR2_X1 U246 ( .A(n216), .B(n275), .Z(product[7]) );
  NAND2_X1 U247 ( .A1(n269), .A2(n40), .ZN(n276) );
  NAND2_X1 U248 ( .A1(n9), .A2(n45), .ZN(n277) );
  NAND2_X1 U249 ( .A1(n40), .A2(n45), .ZN(n278) );
  NAND3_X1 U250 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n8) );
  INV_X2 U251 ( .A(n298), .ZN(n297) );
  XOR2_X1 U252 ( .A(n18), .B(n19), .Z(n279) );
  XOR2_X1 U253 ( .A(n255), .B(n279), .Z(product[12]) );
  NAND2_X1 U254 ( .A1(n231), .A2(n18), .ZN(n280) );
  NAND2_X1 U255 ( .A1(n4), .A2(n19), .ZN(n281) );
  NAND2_X1 U256 ( .A1(n18), .A2(n19), .ZN(n282) );
  NAND3_X1 U257 ( .A1(n281), .A2(n280), .A3(n282), .ZN(n3) );
  XOR2_X1 U258 ( .A(n229), .B(n71), .Z(n283) );
  XOR2_X1 U259 ( .A(n223), .B(n283), .Z(product[3]) );
  NAND2_X1 U260 ( .A1(n223), .A2(n56), .ZN(n284) );
  NAND2_X1 U261 ( .A1(n13), .A2(n71), .ZN(n285) );
  NAND2_X1 U262 ( .A1(n56), .A2(n71), .ZN(n286) );
  NAND3_X1 U263 ( .A1(n284), .A2(n286), .A3(n285), .ZN(n12) );
  XNOR2_X2 U264 ( .A(a[4]), .B(a[3]), .ZN(n326) );
  CLKBUF_X1 U265 ( .A(n212), .Z(n287) );
  XNOR2_X1 U266 ( .A(n219), .B(a[1]), .ZN(n288) );
  INV_X1 U267 ( .A(n15), .ZN(n299) );
  INV_X1 U268 ( .A(n21), .ZN(n302) );
  INV_X1 U269 ( .A(n335), .ZN(n303) );
  INV_X1 U270 ( .A(n315), .ZN(n308) );
  INV_X1 U271 ( .A(n324), .ZN(n306) );
  INV_X1 U272 ( .A(n346), .ZN(n300) );
  INV_X1 U273 ( .A(n31), .ZN(n305) );
  NAND2_X1 U274 ( .A1(n326), .A2(n355), .ZN(n328) );
  INV_X1 U275 ( .A(a[0]), .ZN(n310) );
  INV_X1 U276 ( .A(a[5]), .ZN(n304) );
  INV_X1 U277 ( .A(a[7]), .ZN(n301) );
  INV_X1 U278 ( .A(b[0]), .ZN(n298) );
  XOR2_X1 U279 ( .A(n54), .B(n55), .Z(n289) );
  XOR2_X1 U280 ( .A(n12), .B(n289), .Z(product[4]) );
  NAND2_X1 U281 ( .A1(n240), .A2(n54), .ZN(n290) );
  NAND2_X1 U282 ( .A1(n12), .A2(n55), .ZN(n291) );
  NAND2_X1 U283 ( .A1(n54), .A2(n55), .ZN(n292) );
  NAND3_X1 U284 ( .A1(n290), .A2(n291), .A3(n292), .ZN(n11) );
  XOR2_X1 U285 ( .A(n50), .B(n53), .Z(n293) );
  XOR2_X1 U286 ( .A(n287), .B(n293), .Z(product[5]) );
  NAND2_X1 U287 ( .A1(n212), .A2(n50), .ZN(n294) );
  NAND2_X1 U288 ( .A1(n11), .A2(n53), .ZN(n295) );
  NAND2_X1 U289 ( .A1(n50), .A2(n53), .ZN(n296) );
  NAND3_X1 U290 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n10) );
  INV_X1 U291 ( .A(a[3]), .ZN(n307) );
  INV_X1 U292 ( .A(a[1]), .ZN(n309) );
  NAND2_X2 U293 ( .A1(n316), .A2(n354), .ZN(n318) );
  XOR2_X2 U294 ( .A(a[6]), .B(n304), .Z(n337) );
  NOR2_X1 U295 ( .A1(n310), .A2(n298), .ZN(product[0]) );
  OAI22_X1 U296 ( .A1(n311), .A2(n312), .B1(n313), .B2(n310), .ZN(n99) );
  OAI22_X1 U297 ( .A1(n313), .A2(n312), .B1(n314), .B2(n310), .ZN(n98) );
  XNOR2_X1 U298 ( .A(b[6]), .B(a[1]), .ZN(n313) );
  OAI22_X1 U299 ( .A1(n310), .A2(n314), .B1(n312), .B2(n314), .ZN(n315) );
  XNOR2_X1 U300 ( .A(b[7]), .B(a[1]), .ZN(n314) );
  NOR2_X1 U301 ( .A1(n230), .A2(n298), .ZN(n96) );
  OAI22_X1 U302 ( .A1(n317), .A2(n318), .B1(n230), .B2(n319), .ZN(n95) );
  OAI22_X1 U303 ( .A1(n319), .A2(n318), .B1(n230), .B2(n320), .ZN(n94) );
  XNOR2_X1 U304 ( .A(b[1]), .B(a[3]), .ZN(n319) );
  OAI22_X1 U305 ( .A1(n320), .A2(n318), .B1(n230), .B2(n321), .ZN(n93) );
  XNOR2_X1 U306 ( .A(b[2]), .B(a[3]), .ZN(n320) );
  OAI22_X1 U307 ( .A1(n321), .A2(n318), .B1(n230), .B2(n322), .ZN(n92) );
  XNOR2_X1 U308 ( .A(b[3]), .B(a[3]), .ZN(n321) );
  OAI22_X1 U309 ( .A1(n322), .A2(n318), .B1(n230), .B2(n323), .ZN(n91) );
  XNOR2_X1 U310 ( .A(b[4]), .B(a[3]), .ZN(n322) );
  OAI22_X1 U311 ( .A1(n325), .A2(n230), .B1(n318), .B2(n325), .ZN(n324) );
  NOR2_X1 U312 ( .A1(n326), .A2(n298), .ZN(n88) );
  OAI22_X1 U313 ( .A1(n327), .A2(n328), .B1(n326), .B2(n329), .ZN(n87) );
  XNOR2_X1 U314 ( .A(a[5]), .B(n297), .ZN(n327) );
  OAI22_X1 U315 ( .A1(n329), .A2(n328), .B1(n326), .B2(n330), .ZN(n86) );
  XNOR2_X1 U316 ( .A(n219), .B(a[5]), .ZN(n329) );
  OAI22_X1 U317 ( .A1(n330), .A2(n328), .B1(n326), .B2(n331), .ZN(n85) );
  XNOR2_X1 U318 ( .A(b[2]), .B(a[5]), .ZN(n330) );
  OAI22_X1 U319 ( .A1(n331), .A2(n328), .B1(n326), .B2(n332), .ZN(n84) );
  XNOR2_X1 U320 ( .A(b[3]), .B(a[5]), .ZN(n331) );
  OAI22_X1 U321 ( .A1(n332), .A2(n328), .B1(n326), .B2(n333), .ZN(n83) );
  XNOR2_X1 U322 ( .A(b[4]), .B(a[5]), .ZN(n332) );
  OAI22_X1 U323 ( .A1(n333), .A2(n328), .B1(n326), .B2(n334), .ZN(n82) );
  XNOR2_X1 U324 ( .A(b[5]), .B(a[5]), .ZN(n333) );
  OAI22_X1 U325 ( .A1(n336), .A2(n326), .B1(n328), .B2(n336), .ZN(n335) );
  NOR2_X1 U326 ( .A1(n337), .A2(n298), .ZN(n80) );
  OAI22_X1 U327 ( .A1(n338), .A2(n339), .B1(n337), .B2(n340), .ZN(n79) );
  XNOR2_X1 U328 ( .A(a[7]), .B(n297), .ZN(n338) );
  OAI22_X1 U329 ( .A1(n341), .A2(n339), .B1(n337), .B2(n342), .ZN(n77) );
  OAI22_X1 U330 ( .A1(n342), .A2(n339), .B1(n337), .B2(n343), .ZN(n76) );
  XNOR2_X1 U331 ( .A(b[3]), .B(a[7]), .ZN(n342) );
  OAI22_X1 U332 ( .A1(n343), .A2(n339), .B1(n337), .B2(n344), .ZN(n75) );
  XNOR2_X1 U333 ( .A(b[4]), .B(a[7]), .ZN(n343) );
  OAI22_X1 U334 ( .A1(n344), .A2(n339), .B1(n337), .B2(n345), .ZN(n74) );
  XNOR2_X1 U335 ( .A(b[5]), .B(a[7]), .ZN(n344) );
  OAI22_X1 U336 ( .A1(n347), .A2(n337), .B1(n339), .B2(n347), .ZN(n346) );
  OAI21_X1 U337 ( .B1(n297), .B2(n309), .A(n312), .ZN(n72) );
  OAI21_X1 U338 ( .B1(n307), .B2(n318), .A(n348), .ZN(n71) );
  OR3_X1 U339 ( .A1(n230), .A2(n297), .A3(n307), .ZN(n348) );
  OAI21_X1 U340 ( .B1(n304), .B2(n328), .A(n349), .ZN(n70) );
  OR3_X1 U341 ( .A1(n326), .A2(n297), .A3(n304), .ZN(n349) );
  OAI21_X1 U342 ( .B1(n301), .B2(n339), .A(n350), .ZN(n69) );
  OR3_X1 U343 ( .A1(n337), .A2(n297), .A3(n301), .ZN(n350) );
  XNOR2_X1 U344 ( .A(n351), .B(n352), .ZN(n38) );
  OR2_X1 U345 ( .A1(n351), .A2(n352), .ZN(n37) );
  OAI22_X1 U346 ( .A1(n323), .A2(n318), .B1(n230), .B2(n353), .ZN(n352) );
  XNOR2_X1 U347 ( .A(b[5]), .B(a[3]), .ZN(n323) );
  OAI22_X1 U348 ( .A1(n340), .A2(n339), .B1(n337), .B2(n341), .ZN(n351) );
  XNOR2_X1 U349 ( .A(b[2]), .B(a[7]), .ZN(n341) );
  XNOR2_X1 U350 ( .A(n224), .B(a[7]), .ZN(n340) );
  OAI22_X1 U351 ( .A1(n353), .A2(n318), .B1(n230), .B2(n325), .ZN(n31) );
  XNOR2_X1 U352 ( .A(b[7]), .B(a[3]), .ZN(n325) );
  XNOR2_X1 U353 ( .A(n307), .B(a[2]), .ZN(n354) );
  XNOR2_X1 U354 ( .A(b[6]), .B(a[3]), .ZN(n353) );
  OAI22_X1 U355 ( .A1(n334), .A2(n328), .B1(n326), .B2(n336), .ZN(n21) );
  XNOR2_X1 U356 ( .A(b[7]), .B(a[5]), .ZN(n336) );
  XNOR2_X1 U357 ( .A(n304), .B(a[4]), .ZN(n355) );
  XNOR2_X1 U358 ( .A(b[6]), .B(a[5]), .ZN(n334) );
  OAI22_X1 U359 ( .A1(n345), .A2(n339), .B1(n337), .B2(n347), .ZN(n15) );
  XNOR2_X1 U360 ( .A(b[7]), .B(a[7]), .ZN(n347) );
  NAND2_X1 U361 ( .A1(n337), .A2(n356), .ZN(n339) );
  XNOR2_X1 U362 ( .A(n301), .B(a[6]), .ZN(n356) );
  XNOR2_X1 U363 ( .A(b[6]), .B(a[7]), .ZN(n345) );
  OAI22_X1 U364 ( .A1(n297), .A2(n312), .B1(n357), .B2(n310), .ZN(n104) );
  OAI22_X1 U365 ( .A1(n288), .A2(n312), .B1(n358), .B2(n310), .ZN(n103) );
  XNOR2_X1 U366 ( .A(b[1]), .B(a[1]), .ZN(n357) );
  OAI22_X1 U367 ( .A1(n358), .A2(n312), .B1(n359), .B2(n310), .ZN(n102) );
  XNOR2_X1 U368 ( .A(b[2]), .B(a[1]), .ZN(n358) );
  OAI22_X1 U369 ( .A1(n359), .A2(n312), .B1(n360), .B2(n310), .ZN(n101) );
  XNOR2_X1 U370 ( .A(b[3]), .B(a[1]), .ZN(n359) );
  OAI22_X1 U371 ( .A1(n360), .A2(n312), .B1(n311), .B2(n310), .ZN(n100) );
  XNOR2_X1 U372 ( .A(b[5]), .B(a[1]), .ZN(n311) );
  NAND2_X1 U373 ( .A1(a[1]), .A2(n310), .ZN(n312) );
  XNOR2_X1 U374 ( .A(b[4]), .B(a[1]), .ZN(n360) );
endmodule


module mac_3 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   n6, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, n2, n4;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(n6), .QN(n2) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_3_DW01_add_0 add_356 ( .A(pipeline), .B({mac_out[15:1], n6}), .CI(1'b0), 
        .SUM(sum) );
  mac_3_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n4), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n4), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n4), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n4), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n4), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n4), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n4), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n4), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n4), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n4), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n4), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n4), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n4), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n4), .ZN(N6) );
  INV_X1 U18 ( .A(n2), .ZN(mac_out[0]) );
  AND2_X1 U19 ( .A1(sum[0]), .A2(n4), .ZN(N3) );
  AND2_X1 U20 ( .A1(sum[15]), .A2(n4), .ZN(N18) );
  INV_X1 U21 ( .A(clear_acc), .ZN(n4) );
endmodule


module mac_2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75;
  wire   [15:1] carry;

  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n75) );
  XOR2_X1 U2 ( .A(B[15]), .B(A[15]), .Z(n1) );
  XOR2_X1 U3 ( .A(carry[15]), .B(n1), .Z(SUM[15]) );
  NAND3_X1 U4 ( .A1(n8), .A2(n9), .A3(n10), .ZN(n2) );
  NAND3_X1 U5 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n3) );
  NAND3_X1 U6 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n4) );
  NAND3_X1 U7 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n5) );
  NAND3_X1 U8 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n6) );
  XOR2_X1 U9 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR2_X1 U10 ( .A(n3), .B(n7), .Z(SUM[6]) );
  NAND2_X1 U11 ( .A1(n3), .A2(B[6]), .ZN(n8) );
  NAND2_X1 U12 ( .A1(carry[6]), .A2(A[6]), .ZN(n9) );
  NAND2_X1 U13 ( .A1(B[6]), .A2(A[6]), .ZN(n10) );
  NAND3_X1 U14 ( .A1(n8), .A2(n9), .A3(n10), .ZN(carry[7]) );
  XOR2_X1 U15 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR2_X1 U16 ( .A(n5), .B(n11), .Z(SUM[4]) );
  NAND2_X1 U17 ( .A1(n4), .A2(B[4]), .ZN(n12) );
  NAND2_X1 U18 ( .A1(carry[4]), .A2(A[4]), .ZN(n13) );
  NAND2_X1 U19 ( .A1(B[4]), .A2(A[4]), .ZN(n14) );
  NAND3_X1 U20 ( .A1(n12), .A2(n13), .A3(n14), .ZN(carry[5]) );
  NAND3_X1 U21 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n15) );
  NAND3_X1 U22 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n16) );
  XOR2_X1 U23 ( .A(B[5]), .B(A[5]), .Z(n17) );
  XOR2_X1 U24 ( .A(carry[5]), .B(n17), .Z(SUM[5]) );
  NAND2_X1 U25 ( .A1(carry[5]), .A2(B[5]), .ZN(n18) );
  NAND2_X1 U26 ( .A1(carry[5]), .A2(A[5]), .ZN(n19) );
  NAND2_X1 U27 ( .A1(B[5]), .A2(A[5]), .ZN(n20) );
  NAND3_X1 U28 ( .A1(n18), .A2(n19), .A3(n20), .ZN(carry[6]) );
  NAND3_X1 U29 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n21) );
  NAND3_X1 U30 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n22) );
  XOR2_X1 U31 ( .A(B[7]), .B(A[7]), .Z(n23) );
  XOR2_X1 U32 ( .A(n2), .B(n23), .Z(SUM[7]) );
  NAND2_X1 U33 ( .A1(n2), .A2(B[7]), .ZN(n24) );
  NAND2_X1 U34 ( .A1(carry[7]), .A2(A[7]), .ZN(n25) );
  NAND2_X1 U35 ( .A1(B[7]), .A2(A[7]), .ZN(n26) );
  NAND3_X1 U36 ( .A1(n24), .A2(n25), .A3(n26), .ZN(carry[8]) );
  XOR2_X1 U37 ( .A(B[13]), .B(A[13]), .Z(n27) );
  XOR2_X1 U38 ( .A(n16), .B(n27), .Z(SUM[13]) );
  NAND2_X1 U39 ( .A1(n15), .A2(B[13]), .ZN(n28) );
  NAND2_X1 U40 ( .A1(carry[13]), .A2(A[13]), .ZN(n29) );
  NAND2_X1 U41 ( .A1(B[13]), .A2(A[13]), .ZN(n30) );
  NAND3_X1 U42 ( .A1(n29), .A2(n28), .A3(n30), .ZN(carry[14]) );
  NAND3_X1 U43 ( .A1(n72), .A2(n73), .A3(n74), .ZN(n31) );
  XOR2_X1 U44 ( .A(B[3]), .B(A[3]), .Z(n32) );
  XOR2_X1 U45 ( .A(n31), .B(n32), .Z(SUM[3]) );
  NAND2_X1 U46 ( .A1(n31), .A2(B[3]), .ZN(n33) );
  NAND2_X1 U47 ( .A1(carry[3]), .A2(A[3]), .ZN(n34) );
  NAND2_X1 U48 ( .A1(B[3]), .A2(A[3]), .ZN(n35) );
  NAND3_X1 U49 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[4]) );
  NAND3_X1 U50 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n36) );
  NAND3_X1 U51 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n37) );
  XOR2_X1 U52 ( .A(B[12]), .B(A[12]), .Z(n38) );
  XOR2_X1 U53 ( .A(n37), .B(n38), .Z(SUM[12]) );
  NAND2_X1 U54 ( .A1(n36), .A2(B[12]), .ZN(n39) );
  NAND2_X1 U55 ( .A1(carry[12]), .A2(A[12]), .ZN(n40) );
  NAND2_X1 U56 ( .A1(B[12]), .A2(A[12]), .ZN(n41) );
  NAND3_X1 U57 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[13]) );
  XOR2_X1 U58 ( .A(B[14]), .B(A[14]), .Z(n42) );
  XOR2_X1 U59 ( .A(n6), .B(n42), .Z(SUM[14]) );
  NAND2_X1 U60 ( .A1(n6), .A2(B[14]), .ZN(n43) );
  NAND2_X1 U61 ( .A1(carry[14]), .A2(A[14]), .ZN(n44) );
  NAND2_X1 U62 ( .A1(B[14]), .A2(A[14]), .ZN(n45) );
  NAND3_X1 U63 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[15]) );
  NAND3_X1 U64 ( .A1(n65), .A2(n64), .A3(n66), .ZN(n46) );
  NAND3_X1 U65 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n47) );
  XOR2_X1 U66 ( .A(B[10]), .B(A[10]), .Z(n48) );
  XOR2_X1 U67 ( .A(n47), .B(n48), .Z(SUM[10]) );
  NAND2_X1 U68 ( .A1(n46), .A2(B[10]), .ZN(n49) );
  NAND2_X1 U69 ( .A1(carry[10]), .A2(A[10]), .ZN(n50) );
  NAND2_X1 U70 ( .A1(B[10]), .A2(A[10]), .ZN(n51) );
  NAND3_X1 U71 ( .A1(n49), .A2(n50), .A3(n51), .ZN(carry[11]) );
  XOR2_X1 U72 ( .A(B[11]), .B(A[11]), .Z(n52) );
  XOR2_X1 U73 ( .A(n21), .B(n52), .Z(SUM[11]) );
  NAND2_X1 U74 ( .A1(n21), .A2(B[11]), .ZN(n53) );
  NAND2_X1 U75 ( .A1(carry[11]), .A2(A[11]), .ZN(n54) );
  NAND2_X1 U76 ( .A1(B[11]), .A2(A[11]), .ZN(n55) );
  NAND3_X1 U77 ( .A1(n53), .A2(n54), .A3(n55), .ZN(carry[12]) );
  NAND3_X1 U78 ( .A1(n68), .A2(n69), .A3(n70), .ZN(n56) );
  NAND3_X1 U79 ( .A1(n68), .A2(n69), .A3(n70), .ZN(n57) );
  NAND3_X1 U80 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n58) );
  XOR2_X1 U81 ( .A(B[8]), .B(A[8]), .Z(n59) );
  XOR2_X1 U82 ( .A(n22), .B(n59), .Z(SUM[8]) );
  NAND2_X1 U83 ( .A1(n22), .A2(B[8]), .ZN(n60) );
  NAND2_X1 U84 ( .A1(carry[8]), .A2(A[8]), .ZN(n61) );
  NAND2_X1 U85 ( .A1(B[8]), .A2(A[8]), .ZN(n62) );
  NAND3_X1 U86 ( .A1(n60), .A2(n61), .A3(n62), .ZN(carry[9]) );
  XOR2_X1 U87 ( .A(B[9]), .B(A[9]), .Z(n63) );
  XOR2_X1 U88 ( .A(carry[9]), .B(n63), .Z(SUM[9]) );
  NAND2_X1 U89 ( .A1(n58), .A2(B[9]), .ZN(n64) );
  NAND2_X1 U90 ( .A1(carry[9]), .A2(A[9]), .ZN(n65) );
  NAND2_X1 U91 ( .A1(B[9]), .A2(A[9]), .ZN(n66) );
  NAND3_X1 U92 ( .A1(n65), .A2(n64), .A3(n66), .ZN(carry[10]) );
  XOR2_X1 U93 ( .A(B[1]), .B(A[1]), .Z(n67) );
  XOR2_X1 U94 ( .A(n75), .B(n67), .Z(SUM[1]) );
  NAND2_X1 U95 ( .A1(n75), .A2(B[1]), .ZN(n68) );
  NAND2_X1 U96 ( .A1(n75), .A2(A[1]), .ZN(n69) );
  NAND2_X1 U97 ( .A1(B[1]), .A2(A[1]), .ZN(n70) );
  NAND3_X1 U98 ( .A1(n68), .A2(n69), .A3(n70), .ZN(carry[2]) );
  XOR2_X1 U99 ( .A(B[2]), .B(A[2]), .Z(n71) );
  XOR2_X1 U100 ( .A(n57), .B(n71), .Z(SUM[2]) );
  NAND2_X1 U101 ( .A1(n56), .A2(B[2]), .ZN(n72) );
  NAND2_X1 U102 ( .A1(carry[2]), .A2(A[2]), .ZN(n73) );
  NAND2_X1 U103 ( .A1(B[2]), .A2(A[2]), .ZN(n74) );
  NAND3_X1 U104 ( .A1(n72), .A2(n73), .A3(n74), .ZN(carry[3]) );
  XOR2_X1 U105 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_2_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n209, n210, n211, n212, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n309), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n308), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n312), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n311), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n314), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  CLKBUF_X1 U157 ( .A(n277), .Z(n206) );
  NAND3_X1 U158 ( .A1(n297), .A2(n298), .A3(n299), .ZN(n49) );
  NAND2_X2 U159 ( .A1(n331), .A2(n360), .ZN(n333) );
  INV_X1 U160 ( .A(n284), .ZN(n207) );
  AND2_X1 U161 ( .A1(n212), .A2(n102), .ZN(n208) );
  XNOR2_X1 U162 ( .A(n306), .B(n15), .ZN(n209) );
  NAND2_X1 U163 ( .A1(n251), .A2(n33), .ZN(n210) );
  NAND3_X1 U164 ( .A1(n292), .A2(n293), .A3(n294), .ZN(n211) );
  XOR2_X1 U165 ( .A(n95), .B(n102), .Z(n56) );
  OAI22_X1 U166 ( .A1(n322), .A2(n323), .B1(n282), .B2(n324), .ZN(n212) );
  XNOR2_X1 U167 ( .A(n211), .B(n209), .ZN(product[14]) );
  AND3_X1 U168 ( .A1(n216), .A2(n217), .A3(n218), .ZN(product[15]) );
  NAND3_X1 U169 ( .A1(n292), .A2(n293), .A3(n294), .ZN(n214) );
  CLKBUF_X1 U170 ( .A(n56), .Z(n215) );
  NAND2_X1 U171 ( .A1(n214), .A2(n306), .ZN(n216) );
  NAND2_X1 U172 ( .A1(n2), .A2(n15), .ZN(n217) );
  NAND2_X1 U173 ( .A1(n306), .A2(n15), .ZN(n218) );
  NAND2_X1 U174 ( .A1(n251), .A2(n33), .ZN(n219) );
  NAND3_X1 U175 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n220) );
  NAND3_X1 U176 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n221) );
  NAND3_X1 U177 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n222) );
  NAND3_X1 U178 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n223) );
  XOR2_X1 U179 ( .A(n54), .B(n208), .Z(n224) );
  XOR2_X1 U180 ( .A(n12), .B(n224), .Z(product[4]) );
  NAND2_X1 U181 ( .A1(n220), .A2(n54), .ZN(n225) );
  NAND2_X1 U182 ( .A1(n220), .A2(n208), .ZN(n226) );
  NAND2_X1 U183 ( .A1(n54), .A2(n208), .ZN(n227) );
  NAND3_X1 U184 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n11) );
  CLKBUF_X1 U185 ( .A(n236), .Z(n228) );
  NAND2_X2 U186 ( .A1(n342), .A2(n361), .ZN(n344) );
  XOR2_X2 U187 ( .A(a[6]), .B(n310), .Z(n342) );
  CLKBUF_X1 U188 ( .A(n261), .Z(n229) );
  CLKBUF_X1 U189 ( .A(n290), .Z(n230) );
  NAND3_X1 U190 ( .A1(n288), .A2(n289), .A3(n230), .ZN(n231) );
  AND2_X1 U191 ( .A1(n104), .A2(n72), .ZN(n232) );
  CLKBUF_X1 U192 ( .A(n210), .Z(n233) );
  NAND3_X1 U193 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n234) );
  CLKBUF_X1 U194 ( .A(n222), .Z(n235) );
  NAND3_X1 U195 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n236) );
  XOR2_X1 U196 ( .A(n20), .B(n23), .Z(n237) );
  XOR2_X1 U197 ( .A(n228), .B(n237), .Z(product[11]) );
  NAND2_X1 U198 ( .A1(n236), .A2(n20), .ZN(n238) );
  NAND2_X1 U199 ( .A1(n5), .A2(n23), .ZN(n239) );
  NAND2_X1 U200 ( .A1(n20), .A2(n23), .ZN(n240) );
  NAND3_X1 U201 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n4) );
  NAND3_X1 U202 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n241) );
  XOR2_X1 U203 ( .A(n103), .B(n96), .Z(n242) );
  XOR2_X1 U204 ( .A(n232), .B(n242), .Z(product[2]) );
  NAND2_X1 U205 ( .A1(n232), .A2(n103), .ZN(n243) );
  NAND2_X1 U206 ( .A1(n14), .A2(n96), .ZN(n244) );
  NAND2_X1 U207 ( .A1(n103), .A2(n96), .ZN(n245) );
  NAND3_X1 U208 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n13) );
  CLKBUF_X1 U209 ( .A(b[1]), .Z(n246) );
  XOR2_X1 U210 ( .A(n215), .B(n71), .Z(n247) );
  XOR2_X1 U211 ( .A(n241), .B(n247), .Z(product[3]) );
  NAND2_X1 U212 ( .A1(n241), .A2(n56), .ZN(n248) );
  NAND2_X1 U213 ( .A1(n13), .A2(n71), .ZN(n249) );
  NAND2_X1 U214 ( .A1(n56), .A2(n71), .ZN(n250) );
  NAND3_X1 U215 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n12) );
  NAND3_X1 U216 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n251) );
  CLKBUF_X1 U217 ( .A(n4), .Z(n252) );
  NAND3_X1 U218 ( .A1(n210), .A2(n268), .A3(n269), .ZN(n253) );
  NAND3_X1 U219 ( .A1(n233), .A2(n268), .A3(n269), .ZN(n254) );
  NAND3_X1 U220 ( .A1(n276), .A2(n206), .A3(n278), .ZN(n255) );
  XOR2_X1 U221 ( .A(n27), .B(n24), .Z(n256) );
  XOR2_X1 U222 ( .A(n254), .B(n256), .Z(product[10]) );
  NAND2_X1 U223 ( .A1(n253), .A2(n27), .ZN(n257) );
  NAND2_X1 U224 ( .A1(n6), .A2(n24), .ZN(n258) );
  NAND2_X1 U225 ( .A1(n27), .A2(n24), .ZN(n259) );
  NAND3_X1 U226 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n5) );
  CLKBUF_X1 U227 ( .A(n251), .Z(n260) );
  NAND3_X1 U228 ( .A1(n300), .A2(n301), .A3(n302), .ZN(n261) );
  NAND3_X1 U229 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n262) );
  XOR2_X1 U230 ( .A(n34), .B(n39), .Z(n263) );
  XOR2_X1 U231 ( .A(n255), .B(n263), .Z(product[8]) );
  NAND2_X1 U232 ( .A1(n221), .A2(n34), .ZN(n264) );
  NAND2_X1 U233 ( .A1(n8), .A2(n39), .ZN(n265) );
  NAND2_X1 U234 ( .A1(n34), .A2(n39), .ZN(n266) );
  NAND3_X1 U235 ( .A1(n265), .A2(n264), .A3(n266), .ZN(n7) );
  XOR2_X1 U236 ( .A(n33), .B(n28), .Z(n267) );
  XOR2_X1 U237 ( .A(n260), .B(n267), .Z(product[9]) );
  NAND2_X1 U238 ( .A1(n7), .A2(n28), .ZN(n268) );
  NAND2_X1 U239 ( .A1(n33), .A2(n28), .ZN(n269) );
  NAND3_X1 U240 ( .A1(n219), .A2(n268), .A3(n269), .ZN(n6) );
  INV_X1 U241 ( .A(b[0]), .ZN(n270) );
  XOR2_X1 U242 ( .A(n46), .B(n49), .Z(n271) );
  XOR2_X1 U243 ( .A(n229), .B(n271), .Z(product[6]) );
  NAND2_X1 U244 ( .A1(n261), .A2(n46), .ZN(n272) );
  NAND2_X1 U245 ( .A1(n10), .A2(n49), .ZN(n273) );
  NAND2_X1 U246 ( .A1(n46), .A2(n49), .ZN(n274) );
  NAND3_X1 U247 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n9) );
  XOR2_X1 U248 ( .A(n40), .B(n45), .Z(n275) );
  XOR2_X1 U249 ( .A(n262), .B(n275), .Z(product[7]) );
  NAND2_X1 U250 ( .A1(n223), .A2(n40), .ZN(n276) );
  NAND2_X1 U251 ( .A1(n9), .A2(n45), .ZN(n277) );
  NAND2_X1 U252 ( .A1(n40), .A2(n45), .ZN(n278) );
  NAND3_X1 U253 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n8) );
  XNOR2_X1 U254 ( .A(b[1]), .B(n207), .ZN(n279) );
  NAND2_X2 U255 ( .A1(n321), .A2(n359), .ZN(n323) );
  INV_X2 U256 ( .A(n270), .ZN(n303) );
  NAND3_X1 U257 ( .A1(n290), .A2(n289), .A3(n288), .ZN(n280) );
  XNOR2_X2 U258 ( .A(a[4]), .B(a[3]), .ZN(n331) );
  NAND2_X1 U259 ( .A1(n285), .A2(n286), .ZN(n281) );
  NAND2_X1 U260 ( .A1(n285), .A2(n286), .ZN(n282) );
  NAND2_X1 U261 ( .A1(n285), .A2(n286), .ZN(n321) );
  NAND2_X1 U262 ( .A1(a[2]), .A2(a[1]), .ZN(n285) );
  NAND2_X1 U263 ( .A1(n283), .A2(n284), .ZN(n286) );
  INV_X1 U264 ( .A(a[2]), .ZN(n283) );
  INV_X1 U265 ( .A(a[1]), .ZN(n284) );
  XOR2_X1 U266 ( .A(n295), .B(n52), .Z(n50) );
  INV_X1 U267 ( .A(n15), .ZN(n305) );
  INV_X1 U268 ( .A(n340), .ZN(n309) );
  INV_X1 U269 ( .A(n21), .ZN(n308) );
  INV_X1 U270 ( .A(n320), .ZN(n314) );
  INV_X1 U271 ( .A(n329), .ZN(n312) );
  INV_X1 U272 ( .A(n351), .ZN(n306) );
  INV_X1 U273 ( .A(n31), .ZN(n311) );
  INV_X1 U274 ( .A(a[0]), .ZN(n315) );
  INV_X1 U275 ( .A(a[5]), .ZN(n310) );
  INV_X1 U276 ( .A(a[7]), .ZN(n307) );
  INV_X1 U277 ( .A(b[0]), .ZN(n304) );
  XOR2_X1 U278 ( .A(n19), .B(n18), .Z(n287) );
  XOR2_X1 U279 ( .A(n287), .B(n252), .Z(product[12]) );
  NAND2_X1 U280 ( .A1(n19), .A2(n18), .ZN(n288) );
  NAND2_X1 U281 ( .A1(n19), .A2(n234), .ZN(n289) );
  NAND2_X1 U282 ( .A1(n18), .A2(n4), .ZN(n290) );
  NAND3_X1 U283 ( .A1(n290), .A2(n289), .A3(n288), .ZN(n3) );
  XOR2_X1 U284 ( .A(n17), .B(n305), .Z(n291) );
  XOR2_X1 U285 ( .A(n291), .B(n231), .Z(product[13]) );
  NAND2_X1 U286 ( .A1(n17), .A2(n305), .ZN(n292) );
  NAND2_X1 U287 ( .A1(n17), .A2(n280), .ZN(n293) );
  NAND2_X1 U288 ( .A1(n305), .A2(n3), .ZN(n294) );
  NAND3_X1 U289 ( .A1(n292), .A2(n293), .A3(n294), .ZN(n2) );
  XOR2_X1 U290 ( .A(n93), .B(n100), .Z(n295) );
  XOR2_X1 U291 ( .A(n53), .B(n235), .Z(n296) );
  XOR2_X1 U292 ( .A(n296), .B(n50), .Z(product[5]) );
  NAND2_X1 U293 ( .A1(n93), .A2(n100), .ZN(n297) );
  NAND2_X1 U294 ( .A1(n93), .A2(n52), .ZN(n298) );
  NAND2_X1 U295 ( .A1(n100), .A2(n52), .ZN(n299) );
  NAND2_X1 U296 ( .A1(n53), .A2(n222), .ZN(n300) );
  NAND2_X1 U297 ( .A1(n53), .A2(n50), .ZN(n301) );
  NAND2_X1 U298 ( .A1(n11), .A2(n50), .ZN(n302) );
  NAND3_X1 U299 ( .A1(n300), .A2(n301), .A3(n302), .ZN(n10) );
  INV_X1 U300 ( .A(a[3]), .ZN(n313) );
  NOR2_X1 U301 ( .A1(n315), .A2(n304), .ZN(product[0]) );
  OAI22_X1 U302 ( .A1(n316), .A2(n317), .B1(n318), .B2(n315), .ZN(n99) );
  OAI22_X1 U303 ( .A1(n318), .A2(n317), .B1(n319), .B2(n315), .ZN(n98) );
  XNOR2_X1 U304 ( .A(b[6]), .B(n207), .ZN(n318) );
  OAI22_X1 U305 ( .A1(n315), .A2(n319), .B1(n317), .B2(n319), .ZN(n320) );
  XNOR2_X1 U306 ( .A(b[7]), .B(n207), .ZN(n319) );
  NOR2_X1 U307 ( .A1(n281), .A2(n304), .ZN(n96) );
  OAI22_X1 U308 ( .A1(n322), .A2(n323), .B1(n282), .B2(n324), .ZN(n95) );
  XNOR2_X1 U309 ( .A(a[3]), .B(n303), .ZN(n322) );
  OAI22_X1 U310 ( .A1(n324), .A2(n323), .B1(n282), .B2(n325), .ZN(n94) );
  XNOR2_X1 U311 ( .A(b[1]), .B(a[3]), .ZN(n324) );
  OAI22_X1 U312 ( .A1(n325), .A2(n323), .B1(n281), .B2(n326), .ZN(n93) );
  XNOR2_X1 U313 ( .A(b[2]), .B(a[3]), .ZN(n325) );
  OAI22_X1 U314 ( .A1(n326), .A2(n323), .B1(n282), .B2(n327), .ZN(n92) );
  XNOR2_X1 U315 ( .A(b[3]), .B(a[3]), .ZN(n326) );
  OAI22_X1 U316 ( .A1(n327), .A2(n323), .B1(n282), .B2(n328), .ZN(n91) );
  XNOR2_X1 U317 ( .A(b[4]), .B(a[3]), .ZN(n327) );
  OAI22_X1 U318 ( .A1(n330), .A2(n281), .B1(n323), .B2(n330), .ZN(n329) );
  NOR2_X1 U319 ( .A1(n331), .A2(n304), .ZN(n88) );
  OAI22_X1 U320 ( .A1(n332), .A2(n333), .B1(n331), .B2(n334), .ZN(n87) );
  XNOR2_X1 U321 ( .A(a[5]), .B(n303), .ZN(n332) );
  OAI22_X1 U322 ( .A1(n334), .A2(n333), .B1(n331), .B2(n335), .ZN(n86) );
  XNOR2_X1 U323 ( .A(b[1]), .B(a[5]), .ZN(n334) );
  OAI22_X1 U324 ( .A1(n335), .A2(n333), .B1(n331), .B2(n336), .ZN(n85) );
  XNOR2_X1 U325 ( .A(b[2]), .B(a[5]), .ZN(n335) );
  OAI22_X1 U326 ( .A1(n336), .A2(n333), .B1(n331), .B2(n337), .ZN(n84) );
  XNOR2_X1 U327 ( .A(b[3]), .B(a[5]), .ZN(n336) );
  OAI22_X1 U328 ( .A1(n337), .A2(n333), .B1(n331), .B2(n338), .ZN(n83) );
  XNOR2_X1 U329 ( .A(b[4]), .B(a[5]), .ZN(n337) );
  OAI22_X1 U330 ( .A1(n338), .A2(n333), .B1(n331), .B2(n339), .ZN(n82) );
  XNOR2_X1 U331 ( .A(b[5]), .B(a[5]), .ZN(n338) );
  OAI22_X1 U332 ( .A1(n341), .A2(n331), .B1(n333), .B2(n341), .ZN(n340) );
  NOR2_X1 U333 ( .A1(n342), .A2(n304), .ZN(n80) );
  OAI22_X1 U334 ( .A1(n343), .A2(n344), .B1(n342), .B2(n345), .ZN(n79) );
  XNOR2_X1 U335 ( .A(a[7]), .B(n303), .ZN(n343) );
  OAI22_X1 U336 ( .A1(n346), .A2(n344), .B1(n342), .B2(n347), .ZN(n77) );
  OAI22_X1 U337 ( .A1(n347), .A2(n344), .B1(n342), .B2(n348), .ZN(n76) );
  XNOR2_X1 U338 ( .A(b[3]), .B(a[7]), .ZN(n347) );
  OAI22_X1 U339 ( .A1(n348), .A2(n344), .B1(n342), .B2(n349), .ZN(n75) );
  XNOR2_X1 U340 ( .A(b[4]), .B(a[7]), .ZN(n348) );
  OAI22_X1 U341 ( .A1(n349), .A2(n344), .B1(n342), .B2(n350), .ZN(n74) );
  XNOR2_X1 U342 ( .A(b[5]), .B(a[7]), .ZN(n349) );
  OAI22_X1 U343 ( .A1(n352), .A2(n342), .B1(n344), .B2(n352), .ZN(n351) );
  OAI21_X1 U344 ( .B1(n303), .B2(n284), .A(n317), .ZN(n72) );
  OAI21_X1 U345 ( .B1(n313), .B2(n323), .A(n353), .ZN(n71) );
  OR3_X1 U346 ( .A1(n281), .A2(n303), .A3(n313), .ZN(n353) );
  OAI21_X1 U347 ( .B1(n310), .B2(n333), .A(n354), .ZN(n70) );
  OR3_X1 U348 ( .A1(n331), .A2(n303), .A3(n310), .ZN(n354) );
  OAI21_X1 U349 ( .B1(n307), .B2(n344), .A(n355), .ZN(n69) );
  OR3_X1 U350 ( .A1(n342), .A2(n303), .A3(n307), .ZN(n355) );
  XNOR2_X1 U351 ( .A(n356), .B(n357), .ZN(n38) );
  OR2_X1 U352 ( .A1(n356), .A2(n357), .ZN(n37) );
  OAI22_X1 U353 ( .A1(n328), .A2(n323), .B1(n281), .B2(n358), .ZN(n357) );
  XNOR2_X1 U354 ( .A(b[5]), .B(a[3]), .ZN(n328) );
  OAI22_X1 U355 ( .A1(n345), .A2(n344), .B1(n342), .B2(n346), .ZN(n356) );
  XNOR2_X1 U356 ( .A(b[2]), .B(a[7]), .ZN(n346) );
  XNOR2_X1 U357 ( .A(n246), .B(a[7]), .ZN(n345) );
  OAI22_X1 U358 ( .A1(n358), .A2(n323), .B1(n282), .B2(n330), .ZN(n31) );
  XNOR2_X1 U359 ( .A(b[7]), .B(a[3]), .ZN(n330) );
  XNOR2_X1 U360 ( .A(n313), .B(a[2]), .ZN(n359) );
  XNOR2_X1 U361 ( .A(b[6]), .B(a[3]), .ZN(n358) );
  OAI22_X1 U362 ( .A1(n339), .A2(n333), .B1(n331), .B2(n341), .ZN(n21) );
  XNOR2_X1 U363 ( .A(b[7]), .B(a[5]), .ZN(n341) );
  XNOR2_X1 U364 ( .A(n310), .B(a[4]), .ZN(n360) );
  XNOR2_X1 U365 ( .A(b[6]), .B(a[5]), .ZN(n339) );
  OAI22_X1 U366 ( .A1(n350), .A2(n344), .B1(n342), .B2(n352), .ZN(n15) );
  XNOR2_X1 U367 ( .A(b[7]), .B(a[7]), .ZN(n352) );
  XNOR2_X1 U368 ( .A(n307), .B(a[6]), .ZN(n361) );
  XNOR2_X1 U369 ( .A(b[6]), .B(a[7]), .ZN(n350) );
  OAI22_X1 U370 ( .A1(n303), .A2(n317), .B1(n362), .B2(n315), .ZN(n104) );
  OAI22_X1 U371 ( .A1(n279), .A2(n317), .B1(n363), .B2(n315), .ZN(n103) );
  XNOR2_X1 U372 ( .A(b[1]), .B(a[1]), .ZN(n362) );
  OAI22_X1 U373 ( .A1(n363), .A2(n317), .B1(n364), .B2(n315), .ZN(n102) );
  XNOR2_X1 U374 ( .A(b[2]), .B(a[1]), .ZN(n363) );
  OAI22_X1 U375 ( .A1(n364), .A2(n317), .B1(n365), .B2(n315), .ZN(n101) );
  XNOR2_X1 U376 ( .A(b[3]), .B(a[1]), .ZN(n364) );
  OAI22_X1 U377 ( .A1(n365), .A2(n317), .B1(n316), .B2(n315), .ZN(n100) );
  XNOR2_X1 U378 ( .A(b[5]), .B(n207), .ZN(n316) );
  NAND2_X1 U379 ( .A1(a[1]), .A2(n315), .ZN(n317) );
  XNOR2_X1 U380 ( .A(b[4]), .B(a[1]), .ZN(n365) );
endmodule


module mac_2 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_2_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_2_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72;
  wire   [15:1] carry;

  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n72) );
  XOR2_X1 U2 ( .A(B[15]), .B(A[15]), .Z(n1) );
  XOR2_X1 U3 ( .A(carry[15]), .B(n1), .Z(SUM[15]) );
  NAND3_X1 U4 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n2) );
  XOR2_X1 U5 ( .A(B[2]), .B(A[2]), .Z(n3) );
  XOR2_X1 U6 ( .A(carry[2]), .B(n3), .Z(SUM[2]) );
  NAND2_X1 U7 ( .A1(carry[2]), .A2(B[2]), .ZN(n4) );
  NAND2_X1 U8 ( .A1(carry[2]), .A2(A[2]), .ZN(n5) );
  NAND2_X1 U9 ( .A1(B[2]), .A2(A[2]), .ZN(n6) );
  NAND3_X1 U10 ( .A1(n4), .A2(n5), .A3(n6), .ZN(carry[3]) );
  NAND3_X1 U11 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n7) );
  NAND3_X1 U12 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n8) );
  NAND3_X1 U13 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n9) );
  NAND2_X1 U14 ( .A1(n40), .A2(B[13]), .ZN(n10) );
  NAND3_X1 U15 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n11) );
  NAND3_X1 U16 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n12) );
  XOR2_X1 U17 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR2_X1 U18 ( .A(carry[3]), .B(n13), .Z(SUM[3]) );
  NAND2_X1 U19 ( .A1(carry[3]), .A2(B[3]), .ZN(n14) );
  NAND2_X1 U20 ( .A1(carry[3]), .A2(A[3]), .ZN(n15) );
  NAND2_X1 U21 ( .A1(B[3]), .A2(A[3]), .ZN(n16) );
  NAND3_X1 U22 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[4]) );
  XOR2_X1 U23 ( .A(B[9]), .B(A[9]), .Z(n17) );
  XOR2_X1 U24 ( .A(n2), .B(n17), .Z(SUM[9]) );
  NAND2_X1 U25 ( .A1(n2), .A2(B[9]), .ZN(n18) );
  NAND2_X1 U26 ( .A1(carry[9]), .A2(A[9]), .ZN(n19) );
  NAND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .ZN(n20) );
  NAND3_X1 U28 ( .A1(n18), .A2(n19), .A3(n20), .ZN(carry[10]) );
  XOR2_X1 U29 ( .A(B[10]), .B(A[10]), .Z(n21) );
  XOR2_X1 U30 ( .A(n7), .B(n21), .Z(SUM[10]) );
  NAND2_X1 U31 ( .A1(n7), .A2(B[10]), .ZN(n22) );
  NAND2_X1 U32 ( .A1(carry[10]), .A2(A[10]), .ZN(n23) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n24) );
  NAND3_X1 U34 ( .A1(n22), .A2(n23), .A3(n24), .ZN(carry[11]) );
  NAND3_X1 U35 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n25) );
  NAND3_X1 U36 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n26) );
  NAND3_X1 U37 ( .A1(n10), .A2(n58), .A3(n59), .ZN(n27) );
  XOR2_X1 U38 ( .A(B[4]), .B(A[4]), .Z(n28) );
  XOR2_X1 U39 ( .A(n9), .B(n28), .Z(SUM[4]) );
  NAND2_X1 U40 ( .A1(carry[4]), .A2(B[4]), .ZN(n29) );
  NAND2_X1 U41 ( .A1(n8), .A2(A[4]), .ZN(n30) );
  NAND2_X1 U42 ( .A1(B[4]), .A2(A[4]), .ZN(n31) );
  NAND3_X1 U43 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[5]) );
  XOR2_X1 U44 ( .A(B[11]), .B(A[11]), .Z(n32) );
  XOR2_X1 U45 ( .A(n11), .B(n32), .Z(SUM[11]) );
  NAND2_X1 U46 ( .A1(n11), .A2(B[11]), .ZN(n33) );
  NAND2_X1 U47 ( .A1(carry[11]), .A2(A[11]), .ZN(n34) );
  NAND2_X1 U48 ( .A1(B[11]), .A2(A[11]), .ZN(n35) );
  NAND3_X1 U49 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[12]) );
  XOR2_X1 U50 ( .A(B[5]), .B(A[5]), .Z(n36) );
  XOR2_X1 U51 ( .A(n26), .B(n36), .Z(SUM[5]) );
  NAND2_X1 U52 ( .A1(carry[5]), .A2(B[5]), .ZN(n37) );
  NAND2_X1 U53 ( .A1(carry[5]), .A2(A[5]), .ZN(n38) );
  NAND2_X1 U54 ( .A1(B[5]), .A2(A[5]), .ZN(n39) );
  NAND3_X1 U55 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[6]) );
  NAND3_X1 U56 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n40) );
  XOR2_X1 U57 ( .A(B[12]), .B(A[12]), .Z(n41) );
  XOR2_X1 U58 ( .A(n25), .B(n41), .Z(SUM[12]) );
  NAND2_X1 U59 ( .A1(n25), .A2(B[12]), .ZN(n42) );
  NAND2_X1 U60 ( .A1(carry[12]), .A2(A[12]), .ZN(n43) );
  NAND2_X1 U61 ( .A1(B[12]), .A2(A[12]), .ZN(n44) );
  NAND3_X1 U62 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[13]) );
  NAND3_X1 U63 ( .A1(n10), .A2(n58), .A3(n59), .ZN(n45) );
  NAND3_X1 U64 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n46) );
  NAND3_X1 U65 ( .A1(n69), .A2(n70), .A3(n71), .ZN(n47) );
  XOR2_X1 U66 ( .A(B[8]), .B(A[8]), .Z(n48) );
  XOR2_X1 U67 ( .A(n47), .B(n48), .Z(SUM[8]) );
  NAND2_X1 U68 ( .A1(n47), .A2(B[8]), .ZN(n49) );
  NAND2_X1 U69 ( .A1(carry[8]), .A2(A[8]), .ZN(n50) );
  NAND2_X1 U70 ( .A1(B[8]), .A2(A[8]), .ZN(n51) );
  NAND3_X1 U71 ( .A1(n49), .A2(n50), .A3(n51), .ZN(carry[9]) );
  XOR2_X1 U72 ( .A(B[1]), .B(A[1]), .Z(n52) );
  XOR2_X1 U73 ( .A(n72), .B(n52), .Z(SUM[1]) );
  NAND2_X1 U74 ( .A1(n72), .A2(B[1]), .ZN(n53) );
  NAND2_X1 U75 ( .A1(n72), .A2(A[1]), .ZN(n54) );
  NAND2_X1 U76 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  NAND3_X1 U77 ( .A1(n53), .A2(n54), .A3(n55), .ZN(carry[2]) );
  XOR2_X1 U78 ( .A(B[13]), .B(A[13]), .Z(n56) );
  XOR2_X1 U79 ( .A(n40), .B(n56), .Z(SUM[13]) );
  NAND2_X1 U80 ( .A1(n40), .A2(B[13]), .ZN(n57) );
  NAND2_X1 U81 ( .A1(carry[13]), .A2(A[13]), .ZN(n58) );
  NAND2_X1 U82 ( .A1(B[13]), .A2(A[13]), .ZN(n59) );
  NAND3_X1 U83 ( .A1(n57), .A2(n58), .A3(n59), .ZN(carry[14]) );
  XOR2_X1 U84 ( .A(B[6]), .B(A[6]), .Z(n60) );
  XOR2_X1 U85 ( .A(n12), .B(n60), .Z(SUM[6]) );
  NAND2_X1 U86 ( .A1(n12), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U87 ( .A1(carry[6]), .A2(A[6]), .ZN(n62) );
  NAND2_X1 U88 ( .A1(B[6]), .A2(A[6]), .ZN(n63) );
  NAND3_X1 U89 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[7]) );
  XOR2_X1 U90 ( .A(B[14]), .B(A[14]), .Z(n64) );
  XOR2_X1 U91 ( .A(n27), .B(n64), .Z(SUM[14]) );
  NAND2_X1 U92 ( .A1(n45), .A2(B[14]), .ZN(n65) );
  NAND2_X1 U93 ( .A1(carry[14]), .A2(A[14]), .ZN(n66) );
  NAND2_X1 U94 ( .A1(B[14]), .A2(A[14]), .ZN(n67) );
  NAND3_X1 U95 ( .A1(n65), .A2(n66), .A3(n67), .ZN(carry[15]) );
  XOR2_X1 U96 ( .A(B[7]), .B(A[7]), .Z(n68) );
  XOR2_X1 U97 ( .A(n46), .B(n68), .Z(SUM[7]) );
  NAND2_X1 U98 ( .A1(n46), .A2(B[7]), .ZN(n69) );
  NAND2_X1 U99 ( .A1(carry[7]), .A2(A[7]), .ZN(n70) );
  NAND2_X1 U100 ( .A1(B[7]), .A2(A[7]), .ZN(n71) );
  NAND3_X1 U101 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[8]) );
  XOR2_X1 U102 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_1_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n306), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n305), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n309), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n308), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n311), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  NAND3_X1 U157 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n49) );
  AND2_X1 U158 ( .A1(n95), .A2(n214), .ZN(n206) );
  NAND2_X1 U159 ( .A1(n3), .A2(n302), .ZN(n207) );
  NAND3_X1 U160 ( .A1(n207), .A2(n264), .A3(n265), .ZN(n208) );
  CLKBUF_X1 U161 ( .A(n243), .Z(n209) );
  CLKBUF_X1 U162 ( .A(n280), .Z(n210) );
  NAND3_X1 U163 ( .A1(n217), .A2(n218), .A3(n219), .ZN(n211) );
  NAND3_X1 U164 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n212) );
  NAND3_X1 U165 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n213) );
  XOR2_X1 U166 ( .A(n95), .B(n102), .Z(n56) );
  CLKBUF_X1 U167 ( .A(n102), .Z(n214) );
  XNOR2_X1 U168 ( .A(a[4]), .B(a[3]), .ZN(n328) );
  CLKBUF_X1 U169 ( .A(n211), .Z(n215) );
  XOR2_X1 U170 ( .A(n46), .B(n49), .Z(n216) );
  XOR2_X1 U171 ( .A(n213), .B(n216), .Z(product[6]) );
  NAND2_X1 U172 ( .A1(n212), .A2(n46), .ZN(n217) );
  NAND2_X1 U173 ( .A1(n10), .A2(n49), .ZN(n218) );
  NAND2_X1 U174 ( .A1(n46), .A2(n49), .ZN(n219) );
  NAND3_X1 U175 ( .A1(n217), .A2(n218), .A3(n219), .ZN(n9) );
  NAND3_X1 U176 ( .A1(n280), .A2(n281), .A3(n282), .ZN(n220) );
  NAND3_X1 U177 ( .A1(n210), .A2(n281), .A3(n282), .ZN(n221) );
  XOR2_X1 U178 ( .A(a[3]), .B(n301), .Z(n319) );
  NAND2_X2 U179 ( .A1(n339), .A2(n358), .ZN(n341) );
  XOR2_X2 U180 ( .A(a[6]), .B(n307), .Z(n339) );
  CLKBUF_X1 U181 ( .A(n256), .Z(n222) );
  CLKBUF_X1 U182 ( .A(n286), .Z(n223) );
  CLKBUF_X1 U183 ( .A(n56), .Z(n224) );
  AND2_X1 U184 ( .A1(n104), .A2(n72), .ZN(n225) );
  NAND3_X1 U185 ( .A1(n268), .A2(n267), .A3(n269), .ZN(n226) );
  CLKBUF_X1 U186 ( .A(n251), .Z(n227) );
  CLKBUF_X1 U187 ( .A(n298), .Z(n228) );
  CLKBUF_X1 U188 ( .A(n284), .Z(n229) );
  NAND3_X1 U189 ( .A1(n228), .A2(n297), .A3(n299), .ZN(n230) );
  NAND3_X1 U190 ( .A1(n248), .A2(n247), .A3(n249), .ZN(n231) );
  XOR2_X1 U191 ( .A(n93), .B(n100), .Z(n232) );
  XOR2_X1 U192 ( .A(n52), .B(n232), .Z(n50) );
  NAND2_X1 U193 ( .A1(n236), .A2(n93), .ZN(n233) );
  NAND2_X1 U194 ( .A1(n236), .A2(n100), .ZN(n234) );
  NAND2_X1 U195 ( .A1(n93), .A2(n100), .ZN(n235) );
  CLKBUF_X1 U196 ( .A(n52), .Z(n236) );
  NAND2_X2 U197 ( .A1(n289), .A2(n290), .ZN(n237) );
  NAND2_X1 U198 ( .A1(n289), .A2(n290), .ZN(n318) );
  NAND2_X2 U199 ( .A1(a[1]), .A2(n312), .ZN(n314) );
  NAND3_X1 U200 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n238) );
  NAND3_X1 U201 ( .A1(n284), .A2(n285), .A3(n286), .ZN(n239) );
  NAND3_X1 U202 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n240) );
  CLKBUF_X1 U203 ( .A(n231), .Z(n241) );
  XOR2_X1 U204 ( .A(n40), .B(n45), .Z(n242) );
  XOR2_X1 U205 ( .A(n215), .B(n242), .Z(product[7]) );
  NAND2_X1 U206 ( .A1(n211), .A2(n40), .ZN(n243) );
  NAND2_X1 U207 ( .A1(n9), .A2(n45), .ZN(n244) );
  NAND2_X1 U208 ( .A1(n40), .A2(n45), .ZN(n245) );
  NAND3_X1 U209 ( .A1(n209), .A2(n244), .A3(n245), .ZN(n8) );
  XOR2_X1 U210 ( .A(n20), .B(n23), .Z(n246) );
  XOR2_X1 U211 ( .A(n221), .B(n246), .Z(product[11]) );
  NAND2_X1 U212 ( .A1(n5), .A2(n20), .ZN(n247) );
  NAND2_X1 U213 ( .A1(n220), .A2(n23), .ZN(n248) );
  NAND2_X1 U214 ( .A1(n20), .A2(n23), .ZN(n249) );
  NAND3_X1 U215 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n4) );
  NAND3_X1 U216 ( .A1(n298), .A2(n297), .A3(n299), .ZN(n250) );
  NAND3_X1 U217 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n251) );
  XOR2_X1 U218 ( .A(n34), .B(n39), .Z(n252) );
  XOR2_X1 U219 ( .A(n8), .B(n252), .Z(product[8]) );
  NAND2_X1 U220 ( .A1(n240), .A2(n34), .ZN(n253) );
  NAND2_X1 U221 ( .A1(n240), .A2(n39), .ZN(n254) );
  NAND2_X1 U222 ( .A1(n34), .A2(n39), .ZN(n255) );
  NAND3_X1 U223 ( .A1(n254), .A2(n253), .A3(n255), .ZN(n7) );
  NAND3_X1 U224 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n256) );
  NAND3_X1 U225 ( .A1(n207), .A2(n264), .A3(n265), .ZN(n257) );
  XOR2_X1 U226 ( .A(n54), .B(n206), .Z(n258) );
  XOR2_X1 U227 ( .A(n12), .B(n258), .Z(product[4]) );
  NAND2_X1 U228 ( .A1(n239), .A2(n54), .ZN(n259) );
  NAND2_X1 U229 ( .A1(n239), .A2(n206), .ZN(n260) );
  NAND2_X1 U230 ( .A1(n54), .A2(n206), .ZN(n261) );
  NAND3_X1 U231 ( .A1(n260), .A2(n259), .A3(n261), .ZN(n11) );
  XOR2_X1 U232 ( .A(n302), .B(n17), .Z(n262) );
  XOR2_X1 U233 ( .A(n230), .B(n262), .Z(product[13]) );
  NAND2_X1 U234 ( .A1(n3), .A2(n302), .ZN(n263) );
  NAND2_X1 U235 ( .A1(n250), .A2(n17), .ZN(n264) );
  NAND2_X1 U236 ( .A1(n302), .A2(n17), .ZN(n265) );
  NAND3_X1 U237 ( .A1(n264), .A2(n263), .A3(n265), .ZN(n2) );
  XOR2_X1 U238 ( .A(n103), .B(n96), .Z(n266) );
  XOR2_X1 U239 ( .A(n225), .B(n266), .Z(product[2]) );
  NAND2_X1 U240 ( .A1(n225), .A2(n103), .ZN(n267) );
  NAND2_X1 U241 ( .A1(n14), .A2(n96), .ZN(n268) );
  NAND2_X1 U242 ( .A1(n103), .A2(n96), .ZN(n269) );
  NAND3_X1 U243 ( .A1(n267), .A2(n268), .A3(n269), .ZN(n13) );
  CLKBUF_X1 U244 ( .A(n238), .Z(n270) );
  XOR2_X1 U245 ( .A(n50), .B(n53), .Z(n271) );
  XOR2_X1 U246 ( .A(n222), .B(n271), .Z(product[5]) );
  NAND2_X1 U247 ( .A1(n256), .A2(n50), .ZN(n272) );
  NAND2_X1 U248 ( .A1(n11), .A2(n53), .ZN(n273) );
  NAND2_X1 U249 ( .A1(n50), .A2(n53), .ZN(n274) );
  NAND3_X1 U250 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n10) );
  XOR2_X1 U251 ( .A(n33), .B(n28), .Z(n275) );
  XOR2_X1 U252 ( .A(n227), .B(n275), .Z(product[9]) );
  NAND2_X1 U253 ( .A1(n251), .A2(n33), .ZN(n276) );
  NAND2_X1 U254 ( .A1(n7), .A2(n28), .ZN(n277) );
  NAND2_X1 U255 ( .A1(n33), .A2(n28), .ZN(n278) );
  NAND3_X1 U256 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n6) );
  XOR2_X1 U257 ( .A(n27), .B(n24), .Z(n279) );
  XOR2_X1 U258 ( .A(n270), .B(n279), .Z(product[10]) );
  NAND2_X1 U259 ( .A1(n238), .A2(n27), .ZN(n280) );
  NAND2_X1 U260 ( .A1(n6), .A2(n24), .ZN(n281) );
  NAND2_X1 U261 ( .A1(n27), .A2(n24), .ZN(n282) );
  NAND3_X1 U262 ( .A1(n280), .A2(n281), .A3(n282), .ZN(n5) );
  XOR2_X1 U263 ( .A(n224), .B(n71), .Z(n283) );
  XOR2_X1 U264 ( .A(n226), .B(n283), .Z(product[3]) );
  NAND2_X1 U265 ( .A1(n226), .A2(n56), .ZN(n284) );
  NAND2_X1 U266 ( .A1(n13), .A2(n71), .ZN(n285) );
  NAND2_X1 U267 ( .A1(n56), .A2(n71), .ZN(n286) );
  NAND3_X1 U268 ( .A1(n229), .A2(n285), .A3(n223), .ZN(n12) );
  INV_X2 U269 ( .A(n301), .ZN(n300) );
  NAND2_X2 U270 ( .A1(n328), .A2(n357), .ZN(n330) );
  NAND2_X1 U271 ( .A1(a[2]), .A2(a[1]), .ZN(n289) );
  NAND2_X1 U272 ( .A1(n287), .A2(n288), .ZN(n290) );
  INV_X1 U273 ( .A(a[2]), .ZN(n287) );
  INV_X1 U274 ( .A(a[1]), .ZN(n288) );
  NAND2_X2 U275 ( .A1(n318), .A2(n356), .ZN(n320) );
  INV_X1 U276 ( .A(n15), .ZN(n302) );
  XNOR2_X1 U277 ( .A(n241), .B(n291), .ZN(product[12]) );
  XNOR2_X1 U278 ( .A(n19), .B(n18), .ZN(n291) );
  XNOR2_X1 U279 ( .A(n208), .B(n292), .ZN(product[14]) );
  XNOR2_X1 U280 ( .A(n303), .B(n15), .ZN(n292) );
  AND3_X1 U281 ( .A1(n295), .A2(n294), .A3(n296), .ZN(product[15]) );
  OAI22_X1 U282 ( .A1(n347), .A2(n341), .B1(n339), .B2(n349), .ZN(n15) );
  INV_X1 U283 ( .A(n326), .ZN(n309) );
  INV_X1 U284 ( .A(n337), .ZN(n306) );
  INV_X1 U285 ( .A(n21), .ZN(n305) );
  INV_X1 U286 ( .A(n317), .ZN(n311) );
  INV_X1 U287 ( .A(n31), .ZN(n308) );
  INV_X1 U288 ( .A(a[0]), .ZN(n312) );
  INV_X1 U289 ( .A(a[5]), .ZN(n307) );
  INV_X1 U290 ( .A(a[7]), .ZN(n304) );
  INV_X1 U291 ( .A(b[0]), .ZN(n301) );
  NAND2_X1 U292 ( .A1(n2), .A2(n303), .ZN(n294) );
  NAND2_X1 U293 ( .A1(n257), .A2(n15), .ZN(n295) );
  NAND2_X1 U294 ( .A1(n303), .A2(n15), .ZN(n296) );
  NAND2_X1 U295 ( .A1(n4), .A2(n19), .ZN(n297) );
  NAND2_X1 U296 ( .A1(n231), .A2(n18), .ZN(n298) );
  NAND2_X1 U297 ( .A1(n19), .A2(n18), .ZN(n299) );
  NAND3_X1 U298 ( .A1(n298), .A2(n297), .A3(n299), .ZN(n3) );
  INV_X1 U299 ( .A(n348), .ZN(n303) );
  INV_X1 U300 ( .A(a[3]), .ZN(n310) );
  NOR2_X1 U301 ( .A1(n312), .A2(n301), .ZN(product[0]) );
  OAI22_X1 U302 ( .A1(n313), .A2(n314), .B1(n315), .B2(n312), .ZN(n99) );
  OAI22_X1 U303 ( .A1(n315), .A2(n314), .B1(n316), .B2(n312), .ZN(n98) );
  XNOR2_X1 U304 ( .A(b[6]), .B(a[1]), .ZN(n315) );
  OAI22_X1 U305 ( .A1(n312), .A2(n316), .B1(n314), .B2(n316), .ZN(n317) );
  XNOR2_X1 U306 ( .A(b[7]), .B(a[1]), .ZN(n316) );
  NOR2_X1 U307 ( .A1(n237), .A2(n301), .ZN(n96) );
  OAI22_X1 U308 ( .A1(n319), .A2(n320), .B1(n237), .B2(n321), .ZN(n95) );
  OAI22_X1 U309 ( .A1(n321), .A2(n320), .B1(n237), .B2(n322), .ZN(n94) );
  XNOR2_X1 U310 ( .A(b[1]), .B(a[3]), .ZN(n321) );
  OAI22_X1 U311 ( .A1(n322), .A2(n320), .B1(n237), .B2(n323), .ZN(n93) );
  XNOR2_X1 U312 ( .A(b[2]), .B(a[3]), .ZN(n322) );
  OAI22_X1 U313 ( .A1(n323), .A2(n320), .B1(n237), .B2(n324), .ZN(n92) );
  XNOR2_X1 U314 ( .A(b[3]), .B(a[3]), .ZN(n323) );
  OAI22_X1 U315 ( .A1(n324), .A2(n320), .B1(n237), .B2(n325), .ZN(n91) );
  XNOR2_X1 U316 ( .A(b[4]), .B(a[3]), .ZN(n324) );
  OAI22_X1 U317 ( .A1(n327), .A2(n237), .B1(n320), .B2(n327), .ZN(n326) );
  NOR2_X1 U318 ( .A1(n328), .A2(n301), .ZN(n88) );
  OAI22_X1 U319 ( .A1(n329), .A2(n330), .B1(n328), .B2(n331), .ZN(n87) );
  XNOR2_X1 U320 ( .A(a[5]), .B(n300), .ZN(n329) );
  OAI22_X1 U321 ( .A1(n331), .A2(n330), .B1(n328), .B2(n332), .ZN(n86) );
  XNOR2_X1 U322 ( .A(b[1]), .B(a[5]), .ZN(n331) );
  OAI22_X1 U323 ( .A1(n332), .A2(n330), .B1(n328), .B2(n333), .ZN(n85) );
  XNOR2_X1 U324 ( .A(b[2]), .B(a[5]), .ZN(n332) );
  OAI22_X1 U325 ( .A1(n333), .A2(n330), .B1(n328), .B2(n334), .ZN(n84) );
  XNOR2_X1 U326 ( .A(b[3]), .B(a[5]), .ZN(n333) );
  OAI22_X1 U327 ( .A1(n334), .A2(n330), .B1(n328), .B2(n335), .ZN(n83) );
  XNOR2_X1 U328 ( .A(b[4]), .B(a[5]), .ZN(n334) );
  OAI22_X1 U329 ( .A1(n335), .A2(n330), .B1(n328), .B2(n336), .ZN(n82) );
  XNOR2_X1 U330 ( .A(b[5]), .B(a[5]), .ZN(n335) );
  OAI22_X1 U331 ( .A1(n338), .A2(n328), .B1(n330), .B2(n338), .ZN(n337) );
  NOR2_X1 U332 ( .A1(n339), .A2(n301), .ZN(n80) );
  OAI22_X1 U333 ( .A1(n340), .A2(n341), .B1(n339), .B2(n342), .ZN(n79) );
  XNOR2_X1 U334 ( .A(a[7]), .B(n300), .ZN(n340) );
  OAI22_X1 U335 ( .A1(n343), .A2(n341), .B1(n339), .B2(n344), .ZN(n77) );
  OAI22_X1 U336 ( .A1(n344), .A2(n341), .B1(n339), .B2(n345), .ZN(n76) );
  XNOR2_X1 U337 ( .A(b[3]), .B(a[7]), .ZN(n344) );
  OAI22_X1 U338 ( .A1(n345), .A2(n341), .B1(n339), .B2(n346), .ZN(n75) );
  XNOR2_X1 U339 ( .A(b[4]), .B(a[7]), .ZN(n345) );
  OAI22_X1 U340 ( .A1(n346), .A2(n341), .B1(n339), .B2(n347), .ZN(n74) );
  XNOR2_X1 U341 ( .A(b[5]), .B(a[7]), .ZN(n346) );
  OAI22_X1 U342 ( .A1(n349), .A2(n339), .B1(n341), .B2(n349), .ZN(n348) );
  OAI21_X1 U343 ( .B1(n300), .B2(n288), .A(n314), .ZN(n72) );
  OAI21_X1 U344 ( .B1(n310), .B2(n320), .A(n350), .ZN(n71) );
  OR3_X1 U345 ( .A1(n237), .A2(n300), .A3(n310), .ZN(n350) );
  OAI21_X1 U346 ( .B1(n307), .B2(n330), .A(n351), .ZN(n70) );
  OR3_X1 U347 ( .A1(n328), .A2(n300), .A3(n307), .ZN(n351) );
  OAI21_X1 U348 ( .B1(n304), .B2(n341), .A(n352), .ZN(n69) );
  OR3_X1 U349 ( .A1(n339), .A2(n300), .A3(n304), .ZN(n352) );
  XNOR2_X1 U350 ( .A(n353), .B(n354), .ZN(n38) );
  OR2_X1 U351 ( .A1(n353), .A2(n354), .ZN(n37) );
  OAI22_X1 U352 ( .A1(n325), .A2(n320), .B1(n237), .B2(n355), .ZN(n354) );
  XNOR2_X1 U353 ( .A(b[5]), .B(a[3]), .ZN(n325) );
  OAI22_X1 U354 ( .A1(n342), .A2(n341), .B1(n339), .B2(n343), .ZN(n353) );
  XNOR2_X1 U355 ( .A(b[2]), .B(a[7]), .ZN(n343) );
  XNOR2_X1 U356 ( .A(b[1]), .B(a[7]), .ZN(n342) );
  OAI22_X1 U357 ( .A1(n355), .A2(n320), .B1(n237), .B2(n327), .ZN(n31) );
  XNOR2_X1 U358 ( .A(b[7]), .B(a[3]), .ZN(n327) );
  XNOR2_X1 U359 ( .A(n310), .B(a[2]), .ZN(n356) );
  XNOR2_X1 U360 ( .A(b[6]), .B(a[3]), .ZN(n355) );
  OAI22_X1 U361 ( .A1(n336), .A2(n330), .B1(n328), .B2(n338), .ZN(n21) );
  XNOR2_X1 U362 ( .A(b[7]), .B(a[5]), .ZN(n338) );
  XNOR2_X1 U363 ( .A(n307), .B(a[4]), .ZN(n357) );
  XNOR2_X1 U364 ( .A(b[6]), .B(a[5]), .ZN(n336) );
  XNOR2_X1 U365 ( .A(b[7]), .B(a[7]), .ZN(n349) );
  XNOR2_X1 U366 ( .A(n304), .B(a[6]), .ZN(n358) );
  XNOR2_X1 U367 ( .A(b[6]), .B(a[7]), .ZN(n347) );
  OAI22_X1 U368 ( .A1(n300), .A2(n314), .B1(n359), .B2(n312), .ZN(n104) );
  OAI22_X1 U369 ( .A1(n359), .A2(n314), .B1(n360), .B2(n312), .ZN(n103) );
  XNOR2_X1 U370 ( .A(b[1]), .B(a[1]), .ZN(n359) );
  OAI22_X1 U371 ( .A1(n360), .A2(n314), .B1(n361), .B2(n312), .ZN(n102) );
  XNOR2_X1 U372 ( .A(b[2]), .B(a[1]), .ZN(n360) );
  OAI22_X1 U373 ( .A1(n314), .A2(n361), .B1(n362), .B2(n312), .ZN(n101) );
  XNOR2_X1 U374 ( .A(b[3]), .B(a[1]), .ZN(n361) );
  OAI22_X1 U375 ( .A1(n362), .A2(n314), .B1(n313), .B2(n312), .ZN(n100) );
  XNOR2_X1 U376 ( .A(b[5]), .B(a[1]), .ZN(n313) );
  XNOR2_X1 U377 ( .A(b[4]), .B(a[1]), .ZN(n362) );
endmodule


module mac_1 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n2;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  mac_1_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_1_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  AND2_X1 U3 ( .A1(sum[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U4 ( .A1(sum[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U6 ( .A1(sum[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U10 ( .A1(sum[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U11 ( .A1(sum[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U12 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U13 ( .A1(sum[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U14 ( .A1(sum[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U15 ( .A1(sum[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U16 ( .A1(sum[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U17 ( .A1(sum[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U18 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n2), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n2) );
endmodule


module mac_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65;
  wire   [15:1] carry;

  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n65), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(carry[9]), .Z(n1) );
  XNOR2_X1 U2 ( .A(B[15]), .B(A[15]), .ZN(n2) );
  NAND3_X1 U3 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n3) );
  NAND3_X1 U4 ( .A1(n20), .A2(n21), .A3(n22), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(carry[10]), .Z(n5) );
  NAND3_X1 U6 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n6) );
  NAND3_X1 U7 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n7) );
  CLKBUF_X1 U8 ( .A(n4), .Z(n8) );
  CLKBUF_X1 U9 ( .A(n3), .Z(n9) );
  XOR2_X1 U10 ( .A(B[8]), .B(A[8]), .Z(n10) );
  XOR2_X1 U11 ( .A(carry[8]), .B(n10), .Z(SUM[8]) );
  NAND2_X1 U12 ( .A1(carry[8]), .A2(B[8]), .ZN(n11) );
  NAND2_X1 U13 ( .A1(carry[8]), .A2(A[8]), .ZN(n12) );
  NAND2_X1 U14 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND3_X1 U15 ( .A1(n11), .A2(n12), .A3(n13), .ZN(carry[9]) );
  CLKBUF_X1 U16 ( .A(n48), .Z(n14) );
  XOR2_X1 U17 ( .A(B[9]), .B(A[9]), .Z(n15) );
  XOR2_X1 U18 ( .A(n1), .B(n15), .Z(SUM[9]) );
  NAND2_X1 U19 ( .A1(carry[9]), .A2(B[9]), .ZN(n16) );
  NAND2_X1 U20 ( .A1(carry[9]), .A2(A[9]), .ZN(n17) );
  NAND2_X1 U21 ( .A1(B[9]), .A2(A[9]), .ZN(n18) );
  NAND3_X1 U22 ( .A1(n16), .A2(n17), .A3(n18), .ZN(carry[10]) );
  XOR2_X1 U23 ( .A(B[10]), .B(A[10]), .Z(n19) );
  XOR2_X1 U24 ( .A(n5), .B(n19), .Z(SUM[10]) );
  NAND2_X1 U25 ( .A1(carry[10]), .A2(B[10]), .ZN(n20) );
  NAND2_X1 U26 ( .A1(carry[10]), .A2(A[10]), .ZN(n21) );
  NAND2_X1 U27 ( .A1(B[10]), .A2(A[10]), .ZN(n22) );
  NAND3_X1 U28 ( .A1(n20), .A2(n21), .A3(n22), .ZN(carry[11]) );
  XOR2_X1 U29 ( .A(B[3]), .B(A[3]), .Z(n23) );
  XOR2_X1 U30 ( .A(carry[3]), .B(n23), .Z(SUM[3]) );
  NAND2_X1 U31 ( .A1(carry[3]), .A2(B[3]), .ZN(n24) );
  NAND2_X1 U32 ( .A1(carry[3]), .A2(A[3]), .ZN(n25) );
  NAND2_X1 U33 ( .A1(B[3]), .A2(A[3]), .ZN(n26) );
  NAND3_X1 U34 ( .A1(n24), .A2(n25), .A3(n26), .ZN(carry[4]) );
  NAND3_X1 U35 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n27) );
  XOR2_X1 U36 ( .A(B[11]), .B(A[11]), .Z(n28) );
  XOR2_X1 U37 ( .A(n8), .B(n28), .Z(SUM[11]) );
  NAND2_X1 U38 ( .A1(n4), .A2(B[11]), .ZN(n29) );
  NAND2_X1 U39 ( .A1(carry[11]), .A2(A[11]), .ZN(n30) );
  NAND2_X1 U40 ( .A1(B[11]), .A2(A[11]), .ZN(n31) );
  NAND3_X1 U41 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[12]) );
  XOR2_X1 U42 ( .A(B[4]), .B(A[4]), .Z(n32) );
  XOR2_X1 U43 ( .A(n7), .B(n32), .Z(SUM[4]) );
  NAND2_X1 U44 ( .A1(n6), .A2(B[4]), .ZN(n33) );
  NAND2_X1 U45 ( .A1(carry[4]), .A2(A[4]), .ZN(n34) );
  NAND2_X1 U46 ( .A1(B[4]), .A2(A[4]), .ZN(n35) );
  NAND3_X1 U47 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[5]) );
  NAND3_X1 U48 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n36) );
  NAND3_X1 U49 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n37) );
  XOR2_X1 U50 ( .A(B[12]), .B(A[12]), .Z(n38) );
  XOR2_X1 U51 ( .A(n9), .B(n38), .Z(SUM[12]) );
  NAND2_X1 U52 ( .A1(n3), .A2(B[12]), .ZN(n39) );
  NAND2_X1 U53 ( .A1(carry[12]), .A2(A[12]), .ZN(n40) );
  NAND2_X1 U54 ( .A1(B[12]), .A2(A[12]), .ZN(n41) );
  NAND3_X1 U55 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[13]) );
  XOR2_X1 U56 ( .A(B[5]), .B(A[5]), .Z(n42) );
  XOR2_X1 U57 ( .A(n27), .B(n42), .Z(SUM[5]) );
  NAND2_X1 U58 ( .A1(n27), .A2(B[5]), .ZN(n43) );
  NAND2_X1 U59 ( .A1(carry[5]), .A2(A[5]), .ZN(n44) );
  NAND2_X1 U60 ( .A1(B[5]), .A2(A[5]), .ZN(n45) );
  NAND3_X1 U61 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[6]) );
  XNOR2_X1 U62 ( .A(carry[15]), .B(n2), .ZN(SUM[15]) );
  NAND3_X1 U63 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n46) );
  NAND3_X1 U64 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n47) );
  NAND3_X1 U65 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n48) );
  XOR2_X1 U66 ( .A(B[13]), .B(A[13]), .Z(n49) );
  XOR2_X1 U67 ( .A(carry[13]), .B(n49), .Z(SUM[13]) );
  NAND2_X1 U68 ( .A1(n36), .A2(B[13]), .ZN(n50) );
  NAND2_X1 U69 ( .A1(carry[13]), .A2(A[13]), .ZN(n51) );
  NAND2_X1 U70 ( .A1(B[13]), .A2(A[13]), .ZN(n52) );
  XOR2_X1 U71 ( .A(B[6]), .B(A[6]), .Z(n53) );
  XOR2_X1 U72 ( .A(carry[6]), .B(n53), .Z(SUM[6]) );
  NAND2_X1 U73 ( .A1(n37), .A2(B[6]), .ZN(n54) );
  NAND2_X1 U74 ( .A1(carry[6]), .A2(A[6]), .ZN(n55) );
  NAND2_X1 U75 ( .A1(B[6]), .A2(A[6]), .ZN(n56) );
  NAND3_X1 U76 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[7]) );
  XOR2_X1 U77 ( .A(B[14]), .B(A[14]), .Z(n57) );
  XOR2_X1 U78 ( .A(n47), .B(n57), .Z(SUM[14]) );
  NAND2_X1 U79 ( .A1(n46), .A2(B[14]), .ZN(n58) );
  NAND2_X1 U80 ( .A1(n46), .A2(A[14]), .ZN(n59) );
  NAND2_X1 U81 ( .A1(B[14]), .A2(A[14]), .ZN(n60) );
  NAND3_X1 U82 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[15]) );
  XOR2_X1 U83 ( .A(B[7]), .B(A[7]), .Z(n61) );
  XOR2_X1 U84 ( .A(n14), .B(n61), .Z(SUM[7]) );
  NAND2_X1 U85 ( .A1(n48), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U86 ( .A1(carry[7]), .A2(A[7]), .ZN(n63) );
  NAND2_X1 U87 ( .A1(B[7]), .A2(A[7]), .ZN(n64) );
  NAND3_X1 U88 ( .A1(n62), .A2(n63), .A3(n64), .ZN(carry[8]) );
  AND2_X1 U89 ( .A1(B[0]), .A2(A[0]), .ZN(n65) );
  XOR2_X1 U90 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module mac_0_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n312), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n311), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n315), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n314), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n317), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n88), .B(n101), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n102), .B(n95), .CO(n55), .S(n56) );
  NAND2_X1 U157 ( .A1(n335), .A2(n364), .ZN(n337) );
  INV_X1 U158 ( .A(n20), .ZN(n287) );
  CLKBUF_X1 U159 ( .A(b[1]), .Z(n268) );
  CLKBUF_X1 U160 ( .A(a[5]), .Z(n206) );
  NAND3_X1 U161 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n207) );
  NAND3_X1 U162 ( .A1(n283), .A2(n282), .A3(n281), .ZN(n208) );
  NAND2_X1 U163 ( .A1(n8), .A2(n39), .ZN(n209) );
  NAND2_X2 U164 ( .A1(n236), .A2(n237), .ZN(n210) );
  INV_X2 U165 ( .A(n316), .ZN(n211) );
  NAND2_X1 U166 ( .A1(n236), .A2(n237), .ZN(n335) );
  AND2_X1 U167 ( .A1(n104), .A2(n72), .ZN(n212) );
  CLKBUF_X1 U168 ( .A(n257), .Z(n213) );
  CLKBUF_X1 U169 ( .A(n262), .Z(n214) );
  INV_X1 U170 ( .A(n307), .ZN(n306) );
  CLKBUF_X1 U171 ( .A(n209), .Z(n215) );
  NAND3_X1 U172 ( .A1(n262), .A2(n261), .A3(n263), .ZN(n216) );
  NAND3_X1 U173 ( .A1(n214), .A2(n261), .A3(n263), .ZN(n217) );
  NAND3_X1 U174 ( .A1(n272), .A2(n209), .A3(n274), .ZN(n218) );
  NAND3_X1 U175 ( .A1(n272), .A2(n215), .A3(n274), .ZN(n219) );
  NAND3_X1 U176 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n220) );
  NAND3_X1 U177 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n221) );
  OR2_X1 U178 ( .A1(n288), .A2(n287), .ZN(n222) );
  CLKBUF_X1 U179 ( .A(n9), .Z(n223) );
  CLKBUF_X1 U180 ( .A(n248), .Z(n224) );
  CLKBUF_X1 U181 ( .A(n299), .Z(n225) );
  OR2_X1 U182 ( .A1(n288), .A2(n287), .ZN(n299) );
  NAND3_X1 U183 ( .A1(n247), .A2(n224), .A3(n249), .ZN(n226) );
  NAND3_X1 U184 ( .A1(n231), .A2(n230), .A3(n232), .ZN(n227) );
  NAND3_X1 U185 ( .A1(n265), .A2(n266), .A3(n267), .ZN(n228) );
  XOR2_X1 U186 ( .A(n46), .B(n49), .Z(n229) );
  XOR2_X1 U187 ( .A(n226), .B(n229), .Z(product[6]) );
  NAND2_X1 U188 ( .A1(n207), .A2(n46), .ZN(n230) );
  NAND2_X1 U189 ( .A1(n10), .A2(n49), .ZN(n231) );
  NAND2_X1 U190 ( .A1(n46), .A2(n49), .ZN(n232) );
  NAND3_X1 U191 ( .A1(n230), .A2(n231), .A3(n232), .ZN(n9) );
  NAND3_X1 U192 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n233) );
  NAND3_X1 U193 ( .A1(n255), .A2(n256), .A3(n213), .ZN(n234) );
  NAND2_X1 U194 ( .A1(a[4]), .A2(a[3]), .ZN(n236) );
  NAND2_X1 U195 ( .A1(n235), .A2(n316), .ZN(n237) );
  INV_X1 U196 ( .A(a[4]), .ZN(n235) );
  XOR2_X1 U197 ( .A(n103), .B(n96), .Z(n238) );
  XOR2_X1 U198 ( .A(n212), .B(n238), .Z(product[2]) );
  NAND2_X1 U199 ( .A1(n212), .A2(n103), .ZN(n239) );
  NAND2_X1 U200 ( .A1(n14), .A2(n96), .ZN(n240) );
  NAND2_X1 U201 ( .A1(n103), .A2(n96), .ZN(n241) );
  NAND3_X1 U202 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n13) );
  CLKBUF_X1 U203 ( .A(b[1]), .Z(n242) );
  CLKBUF_X1 U204 ( .A(n228), .Z(n243) );
  NAND3_X1 U205 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n244) );
  NAND3_X1 U206 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n245) );
  XOR2_X1 U207 ( .A(n50), .B(n53), .Z(n246) );
  XOR2_X1 U208 ( .A(n234), .B(n246), .Z(product[5]) );
  NAND2_X1 U209 ( .A1(n233), .A2(n50), .ZN(n247) );
  NAND2_X1 U210 ( .A1(n11), .A2(n53), .ZN(n248) );
  NAND2_X1 U211 ( .A1(n50), .A2(n53), .ZN(n249) );
  NAND3_X1 U212 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n10) );
  XOR2_X1 U213 ( .A(n221), .B(n71), .Z(n250) );
  XOR2_X1 U214 ( .A(n56), .B(n250), .Z(product[3]) );
  NAND2_X1 U215 ( .A1(n220), .A2(n56), .ZN(n251) );
  NAND2_X1 U216 ( .A1(n56), .A2(n71), .ZN(n252) );
  NAND2_X1 U217 ( .A1(n13), .A2(n71), .ZN(n253) );
  NAND3_X1 U218 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n12) );
  XOR2_X1 U219 ( .A(n245), .B(n55), .Z(n254) );
  XOR2_X1 U220 ( .A(n54), .B(n254), .Z(product[4]) );
  NAND2_X1 U221 ( .A1(n244), .A2(n54), .ZN(n255) );
  NAND2_X1 U222 ( .A1(n54), .A2(n55), .ZN(n256) );
  NAND2_X1 U223 ( .A1(n12), .A2(n55), .ZN(n257) );
  NAND3_X1 U224 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n11) );
  XNOR2_X1 U225 ( .A(n258), .B(n277), .ZN(product[14]) );
  XNOR2_X1 U226 ( .A(n309), .B(n15), .ZN(n258) );
  AND3_X1 U227 ( .A1(n286), .A2(n285), .A3(n284), .ZN(product[15]) );
  XOR2_X1 U228 ( .A(n40), .B(n45), .Z(n260) );
  XOR2_X1 U229 ( .A(n223), .B(n260), .Z(product[7]) );
  NAND2_X1 U230 ( .A1(n227), .A2(n40), .ZN(n261) );
  NAND2_X1 U231 ( .A1(n9), .A2(n45), .ZN(n262) );
  NAND2_X1 U232 ( .A1(n40), .A2(n45), .ZN(n263) );
  NAND3_X1 U233 ( .A1(n262), .A2(n261), .A3(n263), .ZN(n8) );
  XOR2_X1 U234 ( .A(n33), .B(n28), .Z(n264) );
  XOR2_X1 U235 ( .A(n219), .B(n264), .Z(product[9]) );
  NAND2_X1 U236 ( .A1(n218), .A2(n33), .ZN(n265) );
  NAND2_X1 U237 ( .A1(n7), .A2(n28), .ZN(n266) );
  NAND2_X1 U238 ( .A1(n33), .A2(n28), .ZN(n267) );
  NAND3_X1 U239 ( .A1(n266), .A2(n265), .A3(n267), .ZN(n6) );
  INV_X1 U240 ( .A(n307), .ZN(n269) );
  INV_X1 U241 ( .A(n269), .ZN(n270) );
  XOR2_X1 U242 ( .A(n34), .B(n39), .Z(n271) );
  XOR2_X1 U243 ( .A(n217), .B(n271), .Z(product[8]) );
  NAND2_X1 U244 ( .A1(n216), .A2(n34), .ZN(n272) );
  NAND2_X1 U245 ( .A1(n8), .A2(n39), .ZN(n273) );
  NAND2_X1 U246 ( .A1(n34), .A2(n39), .ZN(n274) );
  NAND3_X1 U247 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n7) );
  NAND3_X1 U248 ( .A1(n304), .A2(n302), .A3(n303), .ZN(n275) );
  NAND3_X1 U249 ( .A1(n302), .A2(n303), .A3(n304), .ZN(n276) );
  NAND3_X1 U250 ( .A1(n281), .A2(n282), .A3(n283), .ZN(n277) );
  XNOR2_X1 U251 ( .A(a[2]), .B(a[1]), .ZN(n278) );
  XNOR2_X1 U252 ( .A(a[2]), .B(a[1]), .ZN(n279) );
  XNOR2_X1 U253 ( .A(a[2]), .B(a[1]), .ZN(n325) );
  XOR2_X1 U254 ( .A(n17), .B(n308), .Z(n280) );
  XOR2_X1 U255 ( .A(n280), .B(n276), .Z(product[13]) );
  NAND2_X1 U256 ( .A1(n17), .A2(n308), .ZN(n281) );
  NAND2_X1 U257 ( .A1(n275), .A2(n17), .ZN(n282) );
  NAND2_X1 U258 ( .A1(n308), .A2(n3), .ZN(n283) );
  NAND3_X1 U259 ( .A1(n283), .A2(n282), .A3(n281), .ZN(n2) );
  NAND2_X1 U260 ( .A1(n309), .A2(n15), .ZN(n284) );
  NAND2_X1 U261 ( .A1(n2), .A2(n309), .ZN(n285) );
  NAND2_X1 U262 ( .A1(n208), .A2(n15), .ZN(n286) );
  AND3_X1 U263 ( .A1(n293), .A2(n292), .A3(n294), .ZN(n288) );
  NAND3_X1 U264 ( .A1(n293), .A2(n292), .A3(n294), .ZN(n289) );
  CLKBUF_X1 U265 ( .A(b[3]), .Z(n290) );
  XOR2_X1 U266 ( .A(n27), .B(n24), .Z(n291) );
  XOR2_X1 U267 ( .A(n243), .B(n291), .Z(product[10]) );
  NAND2_X1 U268 ( .A1(n6), .A2(n27), .ZN(n292) );
  NAND2_X1 U269 ( .A1(n228), .A2(n24), .ZN(n293) );
  NAND2_X1 U270 ( .A1(n27), .A2(n24), .ZN(n294) );
  NAND3_X1 U271 ( .A1(n300), .A2(n222), .A3(n298), .ZN(n295) );
  NAND3_X1 U272 ( .A1(n298), .A2(n225), .A3(n300), .ZN(n296) );
  INV_X1 U273 ( .A(n15), .ZN(n308) );
  INV_X1 U274 ( .A(n344), .ZN(n312) );
  INV_X1 U275 ( .A(n21), .ZN(n311) );
  INV_X1 U276 ( .A(n324), .ZN(n317) );
  INV_X1 U277 ( .A(n333), .ZN(n315) );
  INV_X1 U278 ( .A(n31), .ZN(n314) );
  INV_X1 U279 ( .A(n355), .ZN(n309) );
  INV_X1 U280 ( .A(a[0]), .ZN(n319) );
  INV_X1 U281 ( .A(a[5]), .ZN(n313) );
  INV_X1 U282 ( .A(a[7]), .ZN(n310) );
  XOR2_X1 U283 ( .A(n20), .B(n23), .Z(n297) );
  XOR2_X1 U284 ( .A(n297), .B(n289), .Z(product[11]) );
  NAND2_X1 U285 ( .A1(n20), .A2(n23), .ZN(n298) );
  NAND2_X1 U286 ( .A1(n23), .A2(n289), .ZN(n300) );
  NAND3_X1 U287 ( .A1(n298), .A2(n299), .A3(n300), .ZN(n4) );
  XOR2_X1 U288 ( .A(n19), .B(n18), .Z(n301) );
  XOR2_X1 U289 ( .A(n301), .B(n296), .Z(product[12]) );
  NAND2_X1 U290 ( .A1(n19), .A2(n18), .ZN(n302) );
  NAND2_X1 U291 ( .A1(n295), .A2(n19), .ZN(n303) );
  NAND2_X1 U292 ( .A1(n4), .A2(n18), .ZN(n304) );
  NAND3_X1 U293 ( .A1(n304), .A2(n302), .A3(n303), .ZN(n3) );
  XNOR2_X1 U294 ( .A(n242), .B(a[1]), .ZN(n305) );
  INV_X1 U295 ( .A(b[0]), .ZN(n307) );
  INV_X1 U296 ( .A(a[3]), .ZN(n316) );
  INV_X1 U297 ( .A(a[1]), .ZN(n318) );
  NAND2_X2 U298 ( .A1(n325), .A2(n363), .ZN(n327) );
  XOR2_X2 U299 ( .A(a[6]), .B(n313), .Z(n346) );
  NOR2_X1 U300 ( .A1(n319), .A2(n270), .ZN(product[0]) );
  OAI22_X1 U301 ( .A1(n320), .A2(n321), .B1(n322), .B2(n319), .ZN(n99) );
  OAI22_X1 U302 ( .A1(n322), .A2(n321), .B1(n323), .B2(n319), .ZN(n98) );
  XNOR2_X1 U303 ( .A(b[6]), .B(a[1]), .ZN(n322) );
  OAI22_X1 U304 ( .A1(n319), .A2(n323), .B1(n321), .B2(n323), .ZN(n324) );
  XNOR2_X1 U305 ( .A(b[7]), .B(a[1]), .ZN(n323) );
  NOR2_X1 U306 ( .A1(n279), .A2(n270), .ZN(n96) );
  OAI22_X1 U307 ( .A1(n326), .A2(n327), .B1(n328), .B2(n278), .ZN(n95) );
  XNOR2_X1 U308 ( .A(n211), .B(n306), .ZN(n326) );
  OAI22_X1 U309 ( .A1(n328), .A2(n327), .B1(n278), .B2(n329), .ZN(n94) );
  XNOR2_X1 U310 ( .A(b[1]), .B(a[3]), .ZN(n328) );
  OAI22_X1 U311 ( .A1(n329), .A2(n327), .B1(n278), .B2(n330), .ZN(n93) );
  XNOR2_X1 U312 ( .A(b[2]), .B(n211), .ZN(n329) );
  OAI22_X1 U313 ( .A1(n330), .A2(n327), .B1(n279), .B2(n331), .ZN(n92) );
  XNOR2_X1 U314 ( .A(n290), .B(n211), .ZN(n330) );
  OAI22_X1 U315 ( .A1(n331), .A2(n327), .B1(n279), .B2(n332), .ZN(n91) );
  XNOR2_X1 U316 ( .A(b[4]), .B(n211), .ZN(n331) );
  OAI22_X1 U317 ( .A1(n334), .A2(n279), .B1(n327), .B2(n334), .ZN(n333) );
  NOR2_X1 U318 ( .A1(n210), .A2(n270), .ZN(n88) );
  OAI22_X1 U319 ( .A1(n336), .A2(n337), .B1(n210), .B2(n338), .ZN(n87) );
  XNOR2_X1 U320 ( .A(a[5]), .B(n269), .ZN(n336) );
  OAI22_X1 U321 ( .A1(n338), .A2(n337), .B1(n210), .B2(n339), .ZN(n86) );
  XNOR2_X1 U322 ( .A(n268), .B(a[5]), .ZN(n338) );
  OAI22_X1 U323 ( .A1(n339), .A2(n337), .B1(n210), .B2(n340), .ZN(n85) );
  XNOR2_X1 U324 ( .A(b[2]), .B(a[5]), .ZN(n339) );
  OAI22_X1 U325 ( .A1(n340), .A2(n337), .B1(n210), .B2(n341), .ZN(n84) );
  XNOR2_X1 U326 ( .A(n290), .B(a[5]), .ZN(n340) );
  OAI22_X1 U327 ( .A1(n341), .A2(n337), .B1(n210), .B2(n342), .ZN(n83) );
  XNOR2_X1 U328 ( .A(b[4]), .B(n206), .ZN(n341) );
  OAI22_X1 U329 ( .A1(n342), .A2(n337), .B1(n210), .B2(n343), .ZN(n82) );
  XNOR2_X1 U330 ( .A(b[5]), .B(n206), .ZN(n342) );
  OAI22_X1 U331 ( .A1(n345), .A2(n210), .B1(n337), .B2(n345), .ZN(n344) );
  NOR2_X1 U332 ( .A1(n346), .A2(n270), .ZN(n80) );
  OAI22_X1 U333 ( .A1(n347), .A2(n348), .B1(n346), .B2(n349), .ZN(n79) );
  XNOR2_X1 U334 ( .A(a[7]), .B(n269), .ZN(n347) );
  OAI22_X1 U335 ( .A1(n350), .A2(n348), .B1(n346), .B2(n351), .ZN(n77) );
  OAI22_X1 U336 ( .A1(n351), .A2(n348), .B1(n346), .B2(n352), .ZN(n76) );
  XNOR2_X1 U337 ( .A(n290), .B(a[7]), .ZN(n351) );
  OAI22_X1 U338 ( .A1(n352), .A2(n348), .B1(n346), .B2(n353), .ZN(n75) );
  XNOR2_X1 U339 ( .A(b[4]), .B(a[7]), .ZN(n352) );
  OAI22_X1 U340 ( .A1(n353), .A2(n348), .B1(n346), .B2(n354), .ZN(n74) );
  XNOR2_X1 U341 ( .A(b[5]), .B(a[7]), .ZN(n353) );
  OAI22_X1 U342 ( .A1(n356), .A2(n346), .B1(n348), .B2(n356), .ZN(n355) );
  OAI21_X1 U343 ( .B1(n306), .B2(n318), .A(n321), .ZN(n72) );
  OAI21_X1 U344 ( .B1(n316), .B2(n327), .A(n357), .ZN(n71) );
  OR3_X1 U345 ( .A1(n279), .A2(n269), .A3(n316), .ZN(n357) );
  OAI21_X1 U346 ( .B1(n313), .B2(n337), .A(n358), .ZN(n70) );
  OR3_X1 U347 ( .A1(n335), .A2(n269), .A3(n313), .ZN(n358) );
  OAI21_X1 U348 ( .B1(n310), .B2(n348), .A(n359), .ZN(n69) );
  OR3_X1 U349 ( .A1(n346), .A2(n269), .A3(n310), .ZN(n359) );
  XNOR2_X1 U350 ( .A(n360), .B(n361), .ZN(n38) );
  OR2_X1 U351 ( .A1(n360), .A2(n361), .ZN(n37) );
  OAI22_X1 U352 ( .A1(n332), .A2(n327), .B1(n278), .B2(n362), .ZN(n361) );
  XNOR2_X1 U353 ( .A(b[5]), .B(n211), .ZN(n332) );
  OAI22_X1 U354 ( .A1(n349), .A2(n348), .B1(n346), .B2(n350), .ZN(n360) );
  XNOR2_X1 U355 ( .A(b[2]), .B(a[7]), .ZN(n350) );
  XNOR2_X1 U356 ( .A(n268), .B(a[7]), .ZN(n349) );
  OAI22_X1 U357 ( .A1(n362), .A2(n327), .B1(n278), .B2(n334), .ZN(n31) );
  XNOR2_X1 U358 ( .A(b[7]), .B(n211), .ZN(n334) );
  XNOR2_X1 U359 ( .A(n316), .B(a[2]), .ZN(n363) );
  XNOR2_X1 U360 ( .A(b[6]), .B(n211), .ZN(n362) );
  OAI22_X1 U361 ( .A1(n343), .A2(n337), .B1(n210), .B2(n345), .ZN(n21) );
  XNOR2_X1 U362 ( .A(b[7]), .B(n206), .ZN(n345) );
  XNOR2_X1 U363 ( .A(n313), .B(a[4]), .ZN(n364) );
  XNOR2_X1 U364 ( .A(b[6]), .B(n206), .ZN(n343) );
  OAI22_X1 U365 ( .A1(n354), .A2(n348), .B1(n346), .B2(n356), .ZN(n15) );
  XNOR2_X1 U366 ( .A(b[7]), .B(a[7]), .ZN(n356) );
  NAND2_X1 U367 ( .A1(n346), .A2(n365), .ZN(n348) );
  XNOR2_X1 U368 ( .A(n310), .B(a[6]), .ZN(n365) );
  XNOR2_X1 U369 ( .A(b[6]), .B(a[7]), .ZN(n354) );
  OAI22_X1 U370 ( .A1(n306), .A2(n321), .B1(n366), .B2(n319), .ZN(n104) );
  OAI22_X1 U371 ( .A1(n305), .A2(n321), .B1(n367), .B2(n319), .ZN(n103) );
  XNOR2_X1 U372 ( .A(b[1]), .B(a[1]), .ZN(n366) );
  OAI22_X1 U373 ( .A1(n367), .A2(n321), .B1(n368), .B2(n319), .ZN(n102) );
  XNOR2_X1 U374 ( .A(b[2]), .B(a[1]), .ZN(n367) );
  OAI22_X1 U375 ( .A1(n368), .A2(n321), .B1(n369), .B2(n319), .ZN(n101) );
  XNOR2_X1 U376 ( .A(b[3]), .B(a[1]), .ZN(n368) );
  OAI22_X1 U377 ( .A1(n369), .A2(n321), .B1(n320), .B2(n319), .ZN(n100) );
  XNOR2_X1 U378 ( .A(b[5]), .B(a[1]), .ZN(n320) );
  NAND2_X1 U379 ( .A1(a[1]), .A2(n319), .ZN(n321) );
  XNOR2_X1 U380 ( .A(b[4]), .B(a[1]), .ZN(n369) );
endmodule


module mac_0 ( clk, clear_acc, a, b, mac_out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] mac_out;
  input clk, clear_acc;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         n3;
  wire   [15:0] mul;
  wire   [15:0] pipeline;
  wire   [15:0] sum;

  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  mac_0_DW01_add_0 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  mac_0_DW_mult_tc_0 mult_355 ( .a(a), .b(b), .product(mul) );
  SDFF_X1 \mac_out_reg[0]  ( .D(1'b0), .SI(n3), .SE(sum[0]), .CK(clk), .Q(
        mac_out[0]) );
  AND2_X1 U4 ( .A1(sum[12]), .A2(n3), .ZN(N15) );
  AND2_X1 U6 ( .A1(sum[11]), .A2(n3), .ZN(N14) );
  AND2_X1 U7 ( .A1(sum[10]), .A2(n3), .ZN(N13) );
  AND2_X1 U8 ( .A1(sum[14]), .A2(n3), .ZN(N17) );
  AND2_X1 U9 ( .A1(sum[13]), .A2(n3), .ZN(N16) );
  AND2_X1 U10 ( .A1(sum[9]), .A2(n3), .ZN(N12) );
  AND2_X1 U11 ( .A1(sum[8]), .A2(n3), .ZN(N11) );
  AND2_X1 U12 ( .A1(sum[7]), .A2(n3), .ZN(N10) );
  AND2_X1 U13 ( .A1(sum[2]), .A2(n3), .ZN(N5) );
  AND2_X1 U14 ( .A1(sum[1]), .A2(n3), .ZN(N4) );
  AND2_X1 U15 ( .A1(sum[6]), .A2(n3), .ZN(N9) );
  AND2_X1 U16 ( .A1(sum[5]), .A2(n3), .ZN(N8) );
  AND2_X1 U17 ( .A1(sum[4]), .A2(n3), .ZN(N7) );
  AND2_X1 U18 ( .A1(sum[3]), .A2(n3), .ZN(N6) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n3), .ZN(N18) );
  INV_X1 U20 ( .A(clear_acc), .ZN(n3) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_31 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;

  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  INV_X1 U3 ( .A(n19), .ZN(n17) );
  NAND3_X1 U4 ( .A1(n35), .A2(wr_en), .A3(n36), .ZN(n19) );
  NOR2_X1 U5 ( .A1(addr[1]), .A2(addr[0]), .ZN(n35) );
  NOR4_X1 U6 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n36) );
  INV_X1 U7 ( .A(n18), .ZN(n16) );
  INV_X1 U8 ( .A(n20), .ZN(n15) );
  AOI22_X1 U9 ( .A1(\mem[0][1] ), .A2(n19), .B1(data_in[1]), .B2(n17), .ZN(n20) );
  INV_X1 U10 ( .A(n21), .ZN(n14) );
  AOI22_X1 U11 ( .A1(\mem[0][2] ), .A2(n19), .B1(data_in[2]), .B2(n17), .ZN(
        n21) );
  INV_X1 U12 ( .A(n22), .ZN(n13) );
  AOI22_X1 U13 ( .A1(\mem[0][3] ), .A2(n19), .B1(data_in[3]), .B2(n17), .ZN(
        n22) );
  INV_X1 U14 ( .A(n23), .ZN(n12) );
  AOI22_X1 U15 ( .A1(\mem[0][4] ), .A2(n19), .B1(data_in[4]), .B2(n17), .ZN(
        n23) );
  INV_X1 U16 ( .A(n24), .ZN(n11) );
  AOI22_X1 U17 ( .A1(\mem[0][5] ), .A2(n19), .B1(data_in[5]), .B2(n17), .ZN(
        n24) );
  INV_X1 U18 ( .A(n25), .ZN(n10) );
  AOI22_X1 U19 ( .A1(\mem[0][6] ), .A2(n19), .B1(data_in[6]), .B2(n17), .ZN(
        n25) );
  INV_X1 U20 ( .A(n26), .ZN(n9) );
  AOI22_X1 U21 ( .A1(\mem[0][7] ), .A2(n19), .B1(data_in[7]), .B2(n17), .ZN(
        n26) );
  INV_X1 U22 ( .A(n27), .ZN(n8) );
  AOI22_X1 U23 ( .A1(\mem[0][8] ), .A2(n19), .B1(data_in[8]), .B2(n17), .ZN(
        n27) );
  INV_X1 U24 ( .A(n28), .ZN(n7) );
  AOI22_X1 U25 ( .A1(\mem[0][9] ), .A2(n19), .B1(data_in[9]), .B2(n17), .ZN(
        n28) );
  INV_X1 U26 ( .A(n29), .ZN(n6) );
  AOI22_X1 U27 ( .A1(\mem[0][10] ), .A2(n19), .B1(data_in[10]), .B2(n17), .ZN(
        n29) );
  INV_X1 U28 ( .A(n30), .ZN(n5) );
  AOI22_X1 U29 ( .A1(\mem[0][11] ), .A2(n19), .B1(data_in[11]), .B2(n17), .ZN(
        n30) );
  INV_X1 U30 ( .A(n31), .ZN(n4) );
  AOI22_X1 U31 ( .A1(\mem[0][12] ), .A2(n19), .B1(data_in[12]), .B2(n17), .ZN(
        n31) );
  INV_X1 U32 ( .A(n32), .ZN(n3) );
  AOI22_X1 U33 ( .A1(\mem[0][13] ), .A2(n19), .B1(data_in[13]), .B2(n17), .ZN(
        n32) );
  INV_X1 U34 ( .A(n33), .ZN(n2) );
  AOI22_X1 U35 ( .A1(\mem[0][14] ), .A2(n19), .B1(data_in[14]), .B2(n17), .ZN(
        n33) );
  INV_X1 U36 ( .A(n34), .ZN(n1) );
  AOI22_X1 U37 ( .A1(\mem[0][15] ), .A2(n19), .B1(data_in[15]), .B2(n17), .ZN(
        n34) );
  AOI22_X1 U38 ( .A1(\mem[0][0] ), .A2(n19), .B1(data_in[0]), .B2(n17), .ZN(
        n18) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_30 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_29 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_28 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_27 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_26 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_25 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_24 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_23 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_22 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_21 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NAND3_X1 U4 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  NOR2_X1 U5 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U6 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U7 ( .A(n55), .ZN(n16) );
  INV_X1 U8 ( .A(n53), .ZN(n15) );
  AOI22_X1 U9 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U10 ( .A(n52), .ZN(n14) );
  AOI22_X1 U11 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U12 ( .A(n51), .ZN(n13) );
  AOI22_X1 U13 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U14 ( .A(n50), .ZN(n12) );
  AOI22_X1 U15 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U16 ( .A(n49), .ZN(n11) );
  AOI22_X1 U17 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U18 ( .A(n48), .ZN(n10) );
  AOI22_X1 U19 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U20 ( .A(n47), .ZN(n9) );
  AOI22_X1 U21 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U22 ( .A(n46), .ZN(n8) );
  AOI22_X1 U23 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U24 ( .A(n45), .ZN(n7) );
  AOI22_X1 U25 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U26 ( .A(n44), .ZN(n6) );
  AOI22_X1 U27 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U28 ( .A(n43), .ZN(n5) );
  AOI22_X1 U29 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U30 ( .A(n42), .ZN(n4) );
  AOI22_X1 U31 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U32 ( .A(n41), .ZN(n3) );
  AOI22_X1 U33 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U34 ( .A(n40), .ZN(n2) );
  AOI22_X1 U35 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U36 ( .A(n39), .ZN(n1) );
  AOI22_X1 U37 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U38 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_20 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NAND3_X1 U4 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  NOR2_X1 U5 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U6 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U7 ( .A(n55), .ZN(n16) );
  INV_X1 U8 ( .A(n53), .ZN(n15) );
  AOI22_X1 U9 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U10 ( .A(n52), .ZN(n14) );
  AOI22_X1 U11 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U12 ( .A(n51), .ZN(n13) );
  AOI22_X1 U13 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U14 ( .A(n50), .ZN(n12) );
  AOI22_X1 U15 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U16 ( .A(n49), .ZN(n11) );
  AOI22_X1 U17 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U18 ( .A(n48), .ZN(n10) );
  AOI22_X1 U19 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U20 ( .A(n47), .ZN(n9) );
  AOI22_X1 U21 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U22 ( .A(n46), .ZN(n8) );
  AOI22_X1 U23 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U24 ( .A(n45), .ZN(n7) );
  AOI22_X1 U25 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U26 ( .A(n44), .ZN(n6) );
  AOI22_X1 U27 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U28 ( .A(n43), .ZN(n5) );
  AOI22_X1 U29 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U30 ( .A(n42), .ZN(n4) );
  AOI22_X1 U31 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U32 ( .A(n41), .ZN(n3) );
  AOI22_X1 U33 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U34 ( .A(n40), .ZN(n2) );
  AOI22_X1 U35 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U36 ( .A(n39), .ZN(n1) );
  AOI22_X1 U37 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U38 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_19 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NAND3_X1 U4 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  NOR2_X1 U5 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U6 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U7 ( .A(n55), .ZN(n16) );
  INV_X1 U8 ( .A(n53), .ZN(n15) );
  AOI22_X1 U9 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U10 ( .A(n52), .ZN(n14) );
  AOI22_X1 U11 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U12 ( .A(n51), .ZN(n13) );
  AOI22_X1 U13 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U14 ( .A(n50), .ZN(n12) );
  AOI22_X1 U15 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U16 ( .A(n49), .ZN(n11) );
  AOI22_X1 U17 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U18 ( .A(n48), .ZN(n10) );
  AOI22_X1 U19 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U20 ( .A(n47), .ZN(n9) );
  AOI22_X1 U21 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U22 ( .A(n46), .ZN(n8) );
  AOI22_X1 U23 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U24 ( .A(n45), .ZN(n7) );
  AOI22_X1 U25 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U26 ( .A(n44), .ZN(n6) );
  AOI22_X1 U27 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U28 ( .A(n43), .ZN(n5) );
  AOI22_X1 U29 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U30 ( .A(n42), .ZN(n4) );
  AOI22_X1 U31 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U32 ( .A(n41), .ZN(n3) );
  AOI22_X1 U33 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U34 ( .A(n40), .ZN(n2) );
  AOI22_X1 U35 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U36 ( .A(n39), .ZN(n1) );
  AOI22_X1 U37 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U38 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_18 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_17 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_16 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_15 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_14 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_13 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_12 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_11 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_10 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_9 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NAND3_X1 U4 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  NOR2_X1 U5 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U6 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U7 ( .A(n55), .ZN(n16) );
  INV_X1 U8 ( .A(n53), .ZN(n15) );
  AOI22_X1 U9 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U10 ( .A(n52), .ZN(n14) );
  AOI22_X1 U11 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U12 ( .A(n51), .ZN(n13) );
  AOI22_X1 U13 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U14 ( .A(n50), .ZN(n12) );
  AOI22_X1 U15 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U16 ( .A(n49), .ZN(n11) );
  AOI22_X1 U17 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U18 ( .A(n48), .ZN(n10) );
  AOI22_X1 U19 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U20 ( .A(n47), .ZN(n9) );
  AOI22_X1 U21 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U22 ( .A(n46), .ZN(n8) );
  AOI22_X1 U23 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U24 ( .A(n45), .ZN(n7) );
  AOI22_X1 U25 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U26 ( .A(n44), .ZN(n6) );
  AOI22_X1 U27 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U28 ( .A(n43), .ZN(n5) );
  AOI22_X1 U29 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U30 ( .A(n42), .ZN(n4) );
  AOI22_X1 U31 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U32 ( .A(n41), .ZN(n3) );
  AOI22_X1 U33 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U34 ( .A(n40), .ZN(n2) );
  AOI22_X1 U35 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U36 ( .A(n39), .ZN(n1) );
  AOI22_X1 U37 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U38 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_8 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NAND3_X1 U4 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  NOR2_X1 U5 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U6 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U7 ( .A(n55), .ZN(n16) );
  INV_X1 U8 ( .A(n53), .ZN(n15) );
  AOI22_X1 U9 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U10 ( .A(n52), .ZN(n14) );
  AOI22_X1 U11 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U12 ( .A(n51), .ZN(n13) );
  AOI22_X1 U13 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U14 ( .A(n50), .ZN(n12) );
  AOI22_X1 U15 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U16 ( .A(n49), .ZN(n11) );
  AOI22_X1 U17 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U18 ( .A(n48), .ZN(n10) );
  AOI22_X1 U19 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U20 ( .A(n47), .ZN(n9) );
  AOI22_X1 U21 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U22 ( .A(n46), .ZN(n8) );
  AOI22_X1 U23 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U24 ( .A(n45), .ZN(n7) );
  AOI22_X1 U25 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U26 ( .A(n44), .ZN(n6) );
  AOI22_X1 U27 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U28 ( .A(n43), .ZN(n5) );
  AOI22_X1 U29 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U30 ( .A(n42), .ZN(n4) );
  AOI22_X1 U31 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U32 ( .A(n41), .ZN(n3) );
  AOI22_X1 U33 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U34 ( .A(n40), .ZN(n2) );
  AOI22_X1 U35 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U36 ( .A(n39), .ZN(n1) );
  AOI22_X1 U37 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U38 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_7 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NAND3_X1 U4 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  NOR2_X1 U5 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U6 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U7 ( .A(n55), .ZN(n16) );
  INV_X1 U8 ( .A(n53), .ZN(n15) );
  AOI22_X1 U9 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U10 ( .A(n52), .ZN(n14) );
  AOI22_X1 U11 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U12 ( .A(n51), .ZN(n13) );
  AOI22_X1 U13 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U14 ( .A(n50), .ZN(n12) );
  AOI22_X1 U15 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U16 ( .A(n49), .ZN(n11) );
  AOI22_X1 U17 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U18 ( .A(n48), .ZN(n10) );
  AOI22_X1 U19 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U20 ( .A(n47), .ZN(n9) );
  AOI22_X1 U21 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U22 ( .A(n46), .ZN(n8) );
  AOI22_X1 U23 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U24 ( .A(n45), .ZN(n7) );
  AOI22_X1 U25 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U26 ( .A(n44), .ZN(n6) );
  AOI22_X1 U27 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U28 ( .A(n43), .ZN(n5) );
  AOI22_X1 U29 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U30 ( .A(n42), .ZN(n4) );
  AOI22_X1 U31 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U32 ( .A(n41), .ZN(n3) );
  AOI22_X1 U33 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U34 ( .A(n40), .ZN(n2) );
  AOI22_X1 U35 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U36 ( .A(n39), .ZN(n1) );
  AOI22_X1 U37 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U38 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_6 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_5 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_4 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_3 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  NAND3_X1 U38 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NOR2_X1 U4 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U5 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U6 ( .A(n55), .ZN(n16) );
  INV_X1 U7 ( .A(n53), .ZN(n15) );
  AOI22_X1 U8 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U9 ( .A(n52), .ZN(n14) );
  AOI22_X1 U10 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U11 ( .A(n51), .ZN(n13) );
  AOI22_X1 U12 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U13 ( .A(n50), .ZN(n12) );
  AOI22_X1 U14 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U15 ( .A(n49), .ZN(n11) );
  AOI22_X1 U16 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U17 ( .A(n48), .ZN(n10) );
  AOI22_X1 U18 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U19 ( .A(n47), .ZN(n9) );
  AOI22_X1 U20 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U21 ( .A(n46), .ZN(n8) );
  AOI22_X1 U22 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U23 ( .A(n45), .ZN(n7) );
  AOI22_X1 U24 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U25 ( .A(n44), .ZN(n6) );
  AOI22_X1 U26 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U27 ( .A(n43), .ZN(n5) );
  AOI22_X1 U28 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U29 ( .A(n42), .ZN(n4) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U31 ( .A(n41), .ZN(n3) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U33 ( .A(n40), .ZN(n2) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U35 ( .A(n39), .ZN(n1) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U37 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_2 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NAND3_X1 U4 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  NOR2_X1 U5 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U6 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U7 ( .A(n55), .ZN(n16) );
  INV_X1 U8 ( .A(n53), .ZN(n15) );
  AOI22_X1 U9 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U10 ( .A(n52), .ZN(n14) );
  AOI22_X1 U11 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U12 ( .A(n51), .ZN(n13) );
  AOI22_X1 U13 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U14 ( .A(n50), .ZN(n12) );
  AOI22_X1 U15 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U16 ( .A(n49), .ZN(n11) );
  AOI22_X1 U17 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U18 ( .A(n48), .ZN(n10) );
  AOI22_X1 U19 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U20 ( .A(n47), .ZN(n9) );
  AOI22_X1 U21 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U22 ( .A(n46), .ZN(n8) );
  AOI22_X1 U23 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U24 ( .A(n45), .ZN(n7) );
  AOI22_X1 U25 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U26 ( .A(n44), .ZN(n6) );
  AOI22_X1 U27 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U28 ( .A(n43), .ZN(n5) );
  AOI22_X1 U29 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U30 ( .A(n42), .ZN(n4) );
  AOI22_X1 U31 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U32 ( .A(n41), .ZN(n3) );
  AOI22_X1 U33 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U34 ( .A(n40), .ZN(n2) );
  AOI22_X1 U35 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U36 ( .A(n39), .ZN(n1) );
  AOI22_X1 U37 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U38 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_1 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NAND3_X1 U4 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  NOR2_X1 U5 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U6 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U7 ( .A(n55), .ZN(n16) );
  INV_X1 U8 ( .A(n53), .ZN(n15) );
  AOI22_X1 U9 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U10 ( .A(n52), .ZN(n14) );
  AOI22_X1 U11 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U12 ( .A(n51), .ZN(n13) );
  AOI22_X1 U13 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U14 ( .A(n50), .ZN(n12) );
  AOI22_X1 U15 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U16 ( .A(n49), .ZN(n11) );
  AOI22_X1 U17 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U18 ( .A(n48), .ZN(n10) );
  AOI22_X1 U19 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U20 ( .A(n47), .ZN(n9) );
  AOI22_X1 U21 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U22 ( .A(n46), .ZN(n8) );
  AOI22_X1 U23 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U24 ( .A(n45), .ZN(n7) );
  AOI22_X1 U25 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U26 ( .A(n44), .ZN(n6) );
  AOI22_X1 U27 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U28 ( .A(n43), .ZN(n5) );
  AOI22_X1 U29 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U30 ( .A(n42), .ZN(n4) );
  AOI22_X1 U31 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U32 ( .A(n41), .ZN(n3) );
  AOI22_X1 U33 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U34 ( .A(n40), .ZN(n2) );
  AOI22_X1 U35 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U36 ( .A(n39), .ZN(n1) );
  AOI22_X1 U37 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U38 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module memory_WIDTH16_SIZE1_LOGSIZE6_0 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;

  DFF_X1 \mem_reg[0][15]  ( .D(n1), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n2), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n3), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n4), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n5), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n6), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n7), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n8), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n9), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n10), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n11), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n12), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n13), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n14), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n15), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n16), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  INV_X1 U3 ( .A(n54), .ZN(n17) );
  NAND3_X1 U4 ( .A1(n38), .A2(wr_en), .A3(n37), .ZN(n54) );
  NOR2_X1 U5 ( .A1(addr[1]), .A2(addr[0]), .ZN(n38) );
  NOR4_X1 U6 ( .A1(addr[5]), .A2(addr[4]), .A3(addr[3]), .A4(addr[2]), .ZN(n37) );
  INV_X1 U7 ( .A(n55), .ZN(n16) );
  INV_X1 U8 ( .A(n53), .ZN(n15) );
  AOI22_X1 U9 ( .A1(\mem[0][1] ), .A2(n54), .B1(data_in[1]), .B2(n17), .ZN(n53) );
  INV_X1 U10 ( .A(n52), .ZN(n14) );
  AOI22_X1 U11 ( .A1(\mem[0][2] ), .A2(n54), .B1(data_in[2]), .B2(n17), .ZN(
        n52) );
  INV_X1 U12 ( .A(n51), .ZN(n13) );
  AOI22_X1 U13 ( .A1(\mem[0][3] ), .A2(n54), .B1(data_in[3]), .B2(n17), .ZN(
        n51) );
  INV_X1 U14 ( .A(n50), .ZN(n12) );
  AOI22_X1 U15 ( .A1(\mem[0][4] ), .A2(n54), .B1(data_in[4]), .B2(n17), .ZN(
        n50) );
  INV_X1 U16 ( .A(n49), .ZN(n11) );
  AOI22_X1 U17 ( .A1(\mem[0][5] ), .A2(n54), .B1(data_in[5]), .B2(n17), .ZN(
        n49) );
  INV_X1 U18 ( .A(n48), .ZN(n10) );
  AOI22_X1 U19 ( .A1(\mem[0][6] ), .A2(n54), .B1(data_in[6]), .B2(n17), .ZN(
        n48) );
  INV_X1 U20 ( .A(n47), .ZN(n9) );
  AOI22_X1 U21 ( .A1(\mem[0][7] ), .A2(n54), .B1(data_in[7]), .B2(n17), .ZN(
        n47) );
  INV_X1 U22 ( .A(n46), .ZN(n8) );
  AOI22_X1 U23 ( .A1(\mem[0][8] ), .A2(n54), .B1(data_in[8]), .B2(n17), .ZN(
        n46) );
  INV_X1 U24 ( .A(n45), .ZN(n7) );
  AOI22_X1 U25 ( .A1(\mem[0][9] ), .A2(n54), .B1(data_in[9]), .B2(n17), .ZN(
        n45) );
  INV_X1 U26 ( .A(n44), .ZN(n6) );
  AOI22_X1 U27 ( .A1(\mem[0][10] ), .A2(n54), .B1(data_in[10]), .B2(n17), .ZN(
        n44) );
  INV_X1 U28 ( .A(n43), .ZN(n5) );
  AOI22_X1 U29 ( .A1(\mem[0][11] ), .A2(n54), .B1(data_in[11]), .B2(n17), .ZN(
        n43) );
  INV_X1 U30 ( .A(n42), .ZN(n4) );
  AOI22_X1 U31 ( .A1(\mem[0][12] ), .A2(n54), .B1(data_in[12]), .B2(n17), .ZN(
        n42) );
  INV_X1 U32 ( .A(n41), .ZN(n3) );
  AOI22_X1 U33 ( .A1(\mem[0][13] ), .A2(n54), .B1(data_in[13]), .B2(n17), .ZN(
        n41) );
  INV_X1 U34 ( .A(n40), .ZN(n2) );
  AOI22_X1 U35 ( .A1(\mem[0][14] ), .A2(n54), .B1(data_in[14]), .B2(n17), .ZN(
        n40) );
  INV_X1 U36 ( .A(n39), .ZN(n1) );
  AOI22_X1 U37 ( .A1(\mem[0][15] ), .A2(n54), .B1(data_in[15]), .B2(n17), .ZN(
        n39) );
  AOI22_X1 U38 ( .A1(\mem[0][0] ), .A2(n54), .B1(data_in[0]), .B2(n17), .ZN(
        n55) );
endmodule


module datapath ( clk, wr_en_x, clear_acc, wr_en_y, addr_x, addr_y, .addr_a({
        \addr_a[31][5] , \addr_a[31][4] , \addr_a[31][3] , \addr_a[31][2] , 
        \addr_a[31][1] , \addr_a[31][0] , \addr_a[30][5] , \addr_a[30][4] , 
        \addr_a[30][3] , \addr_a[30][2] , \addr_a[30][1] , \addr_a[30][0] , 
        \addr_a[29][5] , \addr_a[29][4] , \addr_a[29][3] , \addr_a[29][2] , 
        \addr_a[29][1] , \addr_a[29][0] , \addr_a[28][5] , \addr_a[28][4] , 
        \addr_a[28][3] , \addr_a[28][2] , \addr_a[28][1] , \addr_a[28][0] , 
        \addr_a[27][5] , \addr_a[27][4] , \addr_a[27][3] , \addr_a[27][2] , 
        \addr_a[27][1] , \addr_a[27][0] , \addr_a[26][5] , \addr_a[26][4] , 
        \addr_a[26][3] , \addr_a[26][2] , \addr_a[26][1] , \addr_a[26][0] , 
        \addr_a[25][5] , \addr_a[25][4] , \addr_a[25][3] , \addr_a[25][2] , 
        \addr_a[25][1] , \addr_a[25][0] , \addr_a[24][5] , \addr_a[24][4] , 
        \addr_a[24][3] , \addr_a[24][2] , \addr_a[24][1] , \addr_a[24][0] , 
        \addr_a[23][5] , \addr_a[23][4] , \addr_a[23][3] , \addr_a[23][2] , 
        \addr_a[23][1] , \addr_a[23][0] , \addr_a[22][5] , \addr_a[22][4] , 
        \addr_a[22][3] , \addr_a[22][2] , \addr_a[22][1] , \addr_a[22][0] , 
        \addr_a[21][5] , \addr_a[21][4] , \addr_a[21][3] , \addr_a[21][2] , 
        \addr_a[21][1] , \addr_a[21][0] , \addr_a[20][5] , \addr_a[20][4] , 
        \addr_a[20][3] , \addr_a[20][2] , \addr_a[20][1] , \addr_a[20][0] , 
        \addr_a[19][5] , \addr_a[19][4] , \addr_a[19][3] , \addr_a[19][2] , 
        \addr_a[19][1] , \addr_a[19][0] , \addr_a[18][5] , \addr_a[18][4] , 
        \addr_a[18][3] , \addr_a[18][2] , \addr_a[18][1] , \addr_a[18][0] , 
        \addr_a[17][5] , \addr_a[17][4] , \addr_a[17][3] , \addr_a[17][2] , 
        \addr_a[17][1] , \addr_a[17][0] , \addr_a[16][5] , \addr_a[16][4] , 
        \addr_a[16][3] , \addr_a[16][2] , \addr_a[16][1] , \addr_a[16][0] , 
        \addr_a[15][5] , \addr_a[15][4] , \addr_a[15][3] , \addr_a[15][2] , 
        \addr_a[15][1] , \addr_a[15][0] , \addr_a[14][5] , \addr_a[14][4] , 
        \addr_a[14][3] , \addr_a[14][2] , \addr_a[14][1] , \addr_a[14][0] , 
        \addr_a[13][5] , \addr_a[13][4] , \addr_a[13][3] , \addr_a[13][2] , 
        \addr_a[13][1] , \addr_a[13][0] , \addr_a[12][5] , \addr_a[12][4] , 
        \addr_a[12][3] , \addr_a[12][2] , \addr_a[12][1] , \addr_a[12][0] , 
        \addr_a[11][5] , \addr_a[11][4] , \addr_a[11][3] , \addr_a[11][2] , 
        \addr_a[11][1] , \addr_a[11][0] , \addr_a[10][5] , \addr_a[10][4] , 
        \addr_a[10][3] , \addr_a[10][2] , \addr_a[10][1] , \addr_a[10][0] , 
        \addr_a[9][5] , \addr_a[9][4] , \addr_a[9][3] , \addr_a[9][2] , 
        \addr_a[9][1] , \addr_a[9][0] , \addr_a[8][5] , \addr_a[8][4] , 
        \addr_a[8][3] , \addr_a[8][2] , \addr_a[8][1] , \addr_a[8][0] , 
        \addr_a[7][5] , \addr_a[7][4] , \addr_a[7][3] , \addr_a[7][2] , 
        \addr_a[7][1] , \addr_a[7][0] , \addr_a[6][5] , \addr_a[6][4] , 
        \addr_a[6][3] , \addr_a[6][2] , \addr_a[6][1] , \addr_a[6][0] , 
        \addr_a[5][5] , \addr_a[5][4] , \addr_a[5][3] , \addr_a[5][2] , 
        \addr_a[5][1] , \addr_a[5][0] , \addr_a[4][5] , \addr_a[4][4] , 
        \addr_a[4][3] , \addr_a[4][2] , \addr_a[4][1] , \addr_a[4][0] , 
        \addr_a[3][5] , \addr_a[3][4] , \addr_a[3][3] , \addr_a[3][2] , 
        \addr_a[3][1] , \addr_a[3][0] , \addr_a[2][5] , \addr_a[2][4] , 
        \addr_a[2][3] , \addr_a[2][2] , \addr_a[2][1] , \addr_a[2][0] , 
        \addr_a[1][5] , \addr_a[1][4] , \addr_a[1][3] , \addr_a[1][2] , 
        \addr_a[1][1] , \addr_a[1][0] , \addr_a[0][5] , \addr_a[0][4] , 
        \addr_a[0][3] , \addr_a[0][2] , \addr_a[0][1] , \addr_a[0][0] }), 
        data_in, wr_en_a, data_out );
  input [5:0] addr_x;
  input [5:0] addr_y;
  input [7:0] data_in;
  input [31:0] wr_en_a;
  output [15:0] data_out;
  input clk, wr_en_x, clear_acc, wr_en_y, \addr_a[31][5] , \addr_a[31][4] ,
         \addr_a[31][3] , \addr_a[31][2] , \addr_a[31][1] , \addr_a[31][0] ,
         \addr_a[30][5] , \addr_a[30][4] , \addr_a[30][3] , \addr_a[30][2] ,
         \addr_a[30][1] , \addr_a[30][0] , \addr_a[29][5] , \addr_a[29][4] ,
         \addr_a[29][3] , \addr_a[29][2] , \addr_a[29][1] , \addr_a[29][0] ,
         \addr_a[28][5] , \addr_a[28][4] , \addr_a[28][3] , \addr_a[28][2] ,
         \addr_a[28][1] , \addr_a[28][0] , \addr_a[27][5] , \addr_a[27][4] ,
         \addr_a[27][3] , \addr_a[27][2] , \addr_a[27][1] , \addr_a[27][0] ,
         \addr_a[26][5] , \addr_a[26][4] , \addr_a[26][3] , \addr_a[26][2] ,
         \addr_a[26][1] , \addr_a[26][0] , \addr_a[25][5] , \addr_a[25][4] ,
         \addr_a[25][3] , \addr_a[25][2] , \addr_a[25][1] , \addr_a[25][0] ,
         \addr_a[24][5] , \addr_a[24][4] , \addr_a[24][3] , \addr_a[24][2] ,
         \addr_a[24][1] , \addr_a[24][0] , \addr_a[23][5] , \addr_a[23][4] ,
         \addr_a[23][3] , \addr_a[23][2] , \addr_a[23][1] , \addr_a[23][0] ,
         \addr_a[22][5] , \addr_a[22][4] , \addr_a[22][3] , \addr_a[22][2] ,
         \addr_a[22][1] , \addr_a[22][0] , \addr_a[21][5] , \addr_a[21][4] ,
         \addr_a[21][3] , \addr_a[21][2] , \addr_a[21][1] , \addr_a[21][0] ,
         \addr_a[20][5] , \addr_a[20][4] , \addr_a[20][3] , \addr_a[20][2] ,
         \addr_a[20][1] , \addr_a[20][0] , \addr_a[19][5] , \addr_a[19][4] ,
         \addr_a[19][3] , \addr_a[19][2] , \addr_a[19][1] , \addr_a[19][0] ,
         \addr_a[18][5] , \addr_a[18][4] , \addr_a[18][3] , \addr_a[18][2] ,
         \addr_a[18][1] , \addr_a[18][0] , \addr_a[17][5] , \addr_a[17][4] ,
         \addr_a[17][3] , \addr_a[17][2] , \addr_a[17][1] , \addr_a[17][0] ,
         \addr_a[16][5] , \addr_a[16][4] , \addr_a[16][3] , \addr_a[16][2] ,
         \addr_a[16][1] , \addr_a[16][0] , \addr_a[15][5] , \addr_a[15][4] ,
         \addr_a[15][3] , \addr_a[15][2] , \addr_a[15][1] , \addr_a[15][0] ,
         \addr_a[14][5] , \addr_a[14][4] , \addr_a[14][3] , \addr_a[14][2] ,
         \addr_a[14][1] , \addr_a[14][0] , \addr_a[13][5] , \addr_a[13][4] ,
         \addr_a[13][3] , \addr_a[13][2] , \addr_a[13][1] , \addr_a[13][0] ,
         \addr_a[12][5] , \addr_a[12][4] , \addr_a[12][3] , \addr_a[12][2] ,
         \addr_a[12][1] , \addr_a[12][0] , \addr_a[11][5] , \addr_a[11][4] ,
         \addr_a[11][3] , \addr_a[11][2] , \addr_a[11][1] , \addr_a[11][0] ,
         \addr_a[10][5] , \addr_a[10][4] , \addr_a[10][3] , \addr_a[10][2] ,
         \addr_a[10][1] , \addr_a[10][0] , \addr_a[9][5] , \addr_a[9][4] ,
         \addr_a[9][3] , \addr_a[9][2] , \addr_a[9][1] , \addr_a[9][0] ,
         \addr_a[8][5] , \addr_a[8][4] , \addr_a[8][3] , \addr_a[8][2] ,
         \addr_a[8][1] , \addr_a[8][0] , \addr_a[7][5] , \addr_a[7][4] ,
         \addr_a[7][3] , \addr_a[7][2] , \addr_a[7][1] , \addr_a[7][0] ,
         \addr_a[6][5] , \addr_a[6][4] , \addr_a[6][3] , \addr_a[6][2] ,
         \addr_a[6][1] , \addr_a[6][0] , \addr_a[5][5] , \addr_a[5][4] ,
         \addr_a[5][3] , \addr_a[5][2] , \addr_a[5][1] , \addr_a[5][0] ,
         \addr_a[4][5] , \addr_a[4][4] , \addr_a[4][3] , \addr_a[4][2] ,
         \addr_a[4][1] , \addr_a[4][0] , \addr_a[3][5] , \addr_a[3][4] ,
         \addr_a[3][3] , \addr_a[3][2] , \addr_a[3][1] , \addr_a[3][0] ,
         \addr_a[2][5] , \addr_a[2][4] , \addr_a[2][3] , \addr_a[2][2] ,
         \addr_a[2][1] , \addr_a[2][0] , \addr_a[1][5] , \addr_a[1][4] ,
         \addr_a[1][3] , \addr_a[1][2] , \addr_a[1][1] , \addr_a[1][0] ,
         \addr_a[0][5] , \addr_a[0][4] , \addr_a[0][3] , \addr_a[0][2] ,
         \addr_a[0][1] , \addr_a[0][0] ;
  wire   \matrix_out[31][7] , \matrix_out[31][6] , \matrix_out[31][5] ,
         \matrix_out[31][4] , \matrix_out[31][3] , \matrix_out[31][2] ,
         \matrix_out[31][1] , \matrix_out[31][0] , \matrix_out[30][7] ,
         \matrix_out[30][6] , \matrix_out[30][5] , \matrix_out[30][4] ,
         \matrix_out[30][3] , \matrix_out[30][2] , \matrix_out[30][1] ,
         \matrix_out[30][0] , \matrix_out[29][7] , \matrix_out[29][6] ,
         \matrix_out[29][5] , \matrix_out[29][4] , \matrix_out[29][3] ,
         \matrix_out[29][2] , \matrix_out[29][1] , \matrix_out[29][0] ,
         \matrix_out[28][7] , \matrix_out[28][6] , \matrix_out[28][5] ,
         \matrix_out[28][4] , \matrix_out[28][3] , \matrix_out[28][2] ,
         \matrix_out[28][1] , \matrix_out[28][0] , \matrix_out[27][7] ,
         \matrix_out[27][6] , \matrix_out[27][5] , \matrix_out[27][4] ,
         \matrix_out[27][3] , \matrix_out[27][2] , \matrix_out[27][1] ,
         \matrix_out[27][0] , \matrix_out[26][7] , \matrix_out[26][6] ,
         \matrix_out[26][5] , \matrix_out[26][4] , \matrix_out[26][3] ,
         \matrix_out[26][2] , \matrix_out[26][1] , \matrix_out[26][0] ,
         \matrix_out[25][7] , \matrix_out[25][6] , \matrix_out[25][5] ,
         \matrix_out[25][4] , \matrix_out[25][3] , \matrix_out[25][2] ,
         \matrix_out[25][1] , \matrix_out[25][0] , \matrix_out[24][7] ,
         \matrix_out[24][6] , \matrix_out[24][5] , \matrix_out[24][4] ,
         \matrix_out[24][3] , \matrix_out[24][2] , \matrix_out[24][1] ,
         \matrix_out[24][0] , \matrix_out[23][7] , \matrix_out[23][6] ,
         \matrix_out[23][5] , \matrix_out[23][4] , \matrix_out[23][3] ,
         \matrix_out[23][2] , \matrix_out[23][1] , \matrix_out[23][0] ,
         \matrix_out[22][7] , \matrix_out[22][6] , \matrix_out[22][5] ,
         \matrix_out[22][4] , \matrix_out[22][3] , \matrix_out[22][2] ,
         \matrix_out[22][1] , \matrix_out[22][0] , \matrix_out[21][7] ,
         \matrix_out[21][6] , \matrix_out[21][5] , \matrix_out[21][4] ,
         \matrix_out[21][3] , \matrix_out[21][2] , \matrix_out[21][1] ,
         \matrix_out[21][0] , \matrix_out[20][7] , \matrix_out[20][6] ,
         \matrix_out[20][5] , \matrix_out[20][4] , \matrix_out[20][3] ,
         \matrix_out[20][2] , \matrix_out[20][1] , \matrix_out[20][0] ,
         \matrix_out[19][7] , \matrix_out[19][6] , \matrix_out[19][5] ,
         \matrix_out[19][4] , \matrix_out[19][3] , \matrix_out[19][2] ,
         \matrix_out[19][1] , \matrix_out[19][0] , \matrix_out[18][7] ,
         \matrix_out[18][6] , \matrix_out[18][5] , \matrix_out[18][4] ,
         \matrix_out[18][3] , \matrix_out[18][2] , \matrix_out[18][1] ,
         \matrix_out[18][0] , \matrix_out[17][7] , \matrix_out[17][6] ,
         \matrix_out[17][5] , \matrix_out[17][4] , \matrix_out[17][3] ,
         \matrix_out[17][2] , \matrix_out[17][1] , \matrix_out[17][0] ,
         \matrix_out[16][7] , \matrix_out[16][6] , \matrix_out[16][5] ,
         \matrix_out[16][4] , \matrix_out[16][3] , \matrix_out[16][2] ,
         \matrix_out[16][1] , \matrix_out[16][0] , \matrix_out[15][7] ,
         \matrix_out[15][6] , \matrix_out[15][5] , \matrix_out[15][4] ,
         \matrix_out[15][3] , \matrix_out[15][2] , \matrix_out[15][1] ,
         \matrix_out[15][0] , \matrix_out[14][7] , \matrix_out[14][6] ,
         \matrix_out[14][5] , \matrix_out[14][4] , \matrix_out[14][3] ,
         \matrix_out[14][2] , \matrix_out[14][1] , \matrix_out[14][0] ,
         \matrix_out[13][7] , \matrix_out[13][6] , \matrix_out[13][5] ,
         \matrix_out[13][4] , \matrix_out[13][3] , \matrix_out[13][2] ,
         \matrix_out[13][1] , \matrix_out[13][0] , \matrix_out[12][7] ,
         \matrix_out[12][6] , \matrix_out[12][5] , \matrix_out[12][4] ,
         \matrix_out[12][3] , \matrix_out[12][2] , \matrix_out[12][1] ,
         \matrix_out[12][0] , \matrix_out[11][7] , \matrix_out[11][6] ,
         \matrix_out[11][5] , \matrix_out[11][4] , \matrix_out[11][3] ,
         \matrix_out[11][2] , \matrix_out[11][1] , \matrix_out[11][0] ,
         \matrix_out[10][7] , \matrix_out[10][6] , \matrix_out[10][5] ,
         \matrix_out[10][4] , \matrix_out[10][3] , \matrix_out[10][2] ,
         \matrix_out[10][1] , \matrix_out[10][0] , \matrix_out[9][7] ,
         \matrix_out[9][6] , \matrix_out[9][5] , \matrix_out[9][4] ,
         \matrix_out[9][3] , \matrix_out[9][2] , \matrix_out[9][1] ,
         \matrix_out[9][0] , \matrix_out[8][7] , \matrix_out[8][6] ,
         \matrix_out[8][5] , \matrix_out[8][4] , \matrix_out[8][3] ,
         \matrix_out[8][2] , \matrix_out[8][1] , \matrix_out[8][0] ,
         \matrix_out[7][7] , \matrix_out[7][6] , \matrix_out[7][5] ,
         \matrix_out[7][4] , \matrix_out[7][3] , \matrix_out[7][2] ,
         \matrix_out[7][1] , \matrix_out[7][0] , \matrix_out[6][7] ,
         \matrix_out[6][6] , \matrix_out[6][5] , \matrix_out[6][4] ,
         \matrix_out[6][3] , \matrix_out[6][2] , \matrix_out[6][1] ,
         \matrix_out[6][0] , \matrix_out[5][7] , \matrix_out[5][6] ,
         \matrix_out[5][5] , \matrix_out[5][4] , \matrix_out[5][3] ,
         \matrix_out[5][2] , \matrix_out[5][1] , \matrix_out[5][0] ,
         \matrix_out[4][7] , \matrix_out[4][6] , \matrix_out[4][5] ,
         \matrix_out[4][4] , \matrix_out[4][3] , \matrix_out[4][2] ,
         \matrix_out[4][1] , \matrix_out[4][0] , \matrix_out[3][7] ,
         \matrix_out[3][6] , \matrix_out[3][5] , \matrix_out[3][4] ,
         \matrix_out[3][3] , \matrix_out[3][2] , \matrix_out[3][1] ,
         \matrix_out[3][0] , \matrix_out[2][7] , \matrix_out[2][6] ,
         \matrix_out[2][5] , \matrix_out[2][4] , \matrix_out[2][3] ,
         \matrix_out[2][2] , \matrix_out[2][1] , \matrix_out[2][0] ,
         \matrix_out[1][7] , \matrix_out[1][6] , \matrix_out[1][5] ,
         \matrix_out[1][4] , \matrix_out[1][3] , \matrix_out[1][2] ,
         \matrix_out[1][1] , \matrix_out[1][0] , \matrix_out[0][7] ,
         \matrix_out[0][6] , \matrix_out[0][5] , \matrix_out[0][4] ,
         \matrix_out[0][3] , \matrix_out[0][2] , \matrix_out[0][1] ,
         \matrix_out[0][0] , \mac_out[31][15] , \mac_out[31][14] ,
         \mac_out[31][13] , \mac_out[31][12] , \mac_out[31][11] ,
         \mac_out[31][10] , \mac_out[31][9] , \mac_out[31][8] ,
         \mac_out[31][7] , \mac_out[31][6] , \mac_out[31][5] ,
         \mac_out[31][4] , \mac_out[31][3] , \mac_out[31][2] ,
         \mac_out[31][1] , \mac_out[31][0] , \mac_out[30][15] ,
         \mac_out[30][14] , \mac_out[30][13] , \mac_out[30][12] ,
         \mac_out[30][11] , \mac_out[30][10] , \mac_out[30][9] ,
         \mac_out[30][8] , \mac_out[30][7] , \mac_out[30][6] ,
         \mac_out[30][5] , \mac_out[30][4] , \mac_out[30][3] ,
         \mac_out[30][2] , \mac_out[30][1] , \mac_out[30][0] ,
         \mac_out[29][15] , \mac_out[29][14] , \mac_out[29][13] ,
         \mac_out[29][12] , \mac_out[29][11] , \mac_out[29][10] ,
         \mac_out[29][9] , \mac_out[29][8] , \mac_out[29][7] ,
         \mac_out[29][6] , \mac_out[29][5] , \mac_out[29][4] ,
         \mac_out[29][3] , \mac_out[29][2] , \mac_out[29][1] ,
         \mac_out[29][0] , \mac_out[28][15] , \mac_out[28][14] ,
         \mac_out[28][13] , \mac_out[28][12] , \mac_out[28][11] ,
         \mac_out[28][10] , \mac_out[28][9] , \mac_out[28][8] ,
         \mac_out[28][7] , \mac_out[28][6] , \mac_out[28][5] ,
         \mac_out[28][4] , \mac_out[28][3] , \mac_out[28][2] ,
         \mac_out[28][1] , \mac_out[28][0] , \mac_out[27][15] ,
         \mac_out[27][14] , \mac_out[27][13] , \mac_out[27][12] ,
         \mac_out[27][11] , \mac_out[27][10] , \mac_out[27][9] ,
         \mac_out[27][8] , \mac_out[27][7] , \mac_out[27][6] ,
         \mac_out[27][5] , \mac_out[27][4] , \mac_out[27][3] ,
         \mac_out[27][2] , \mac_out[27][1] , \mac_out[27][0] ,
         \mac_out[26][15] , \mac_out[26][14] , \mac_out[26][13] ,
         \mac_out[26][12] , \mac_out[26][11] , \mac_out[26][10] ,
         \mac_out[26][9] , \mac_out[26][8] , \mac_out[26][7] ,
         \mac_out[26][6] , \mac_out[26][5] , \mac_out[26][4] ,
         \mac_out[26][3] , \mac_out[26][2] , \mac_out[26][1] ,
         \mac_out[26][0] , \mac_out[25][15] , \mac_out[25][14] ,
         \mac_out[25][13] , \mac_out[25][12] , \mac_out[25][11] ,
         \mac_out[25][10] , \mac_out[25][9] , \mac_out[25][8] ,
         \mac_out[25][7] , \mac_out[25][6] , \mac_out[25][5] ,
         \mac_out[25][4] , \mac_out[25][3] , \mac_out[25][2] ,
         \mac_out[25][1] , \mac_out[25][0] , \mac_out[24][15] ,
         \mac_out[24][14] , \mac_out[24][13] , \mac_out[24][12] ,
         \mac_out[24][11] , \mac_out[24][10] , \mac_out[24][9] ,
         \mac_out[24][8] , \mac_out[24][7] , \mac_out[24][6] ,
         \mac_out[24][5] , \mac_out[24][4] , \mac_out[24][3] ,
         \mac_out[24][2] , \mac_out[24][1] , \mac_out[24][0] ,
         \mac_out[23][15] , \mac_out[23][14] , \mac_out[23][13] ,
         \mac_out[23][12] , \mac_out[23][11] , \mac_out[23][10] ,
         \mac_out[23][9] , \mac_out[23][8] , \mac_out[23][7] ,
         \mac_out[23][6] , \mac_out[23][5] , \mac_out[23][4] ,
         \mac_out[23][3] , \mac_out[23][2] , \mac_out[23][1] ,
         \mac_out[23][0] , \mac_out[22][15] , \mac_out[22][14] ,
         \mac_out[22][13] , \mac_out[22][12] , \mac_out[22][11] ,
         \mac_out[22][10] , \mac_out[22][9] , \mac_out[22][8] ,
         \mac_out[22][7] , \mac_out[22][6] , \mac_out[22][5] ,
         \mac_out[22][4] , \mac_out[22][3] , \mac_out[22][2] ,
         \mac_out[22][1] , \mac_out[22][0] , \mac_out[21][15] ,
         \mac_out[21][14] , \mac_out[21][13] , \mac_out[21][12] ,
         \mac_out[21][11] , \mac_out[21][10] , \mac_out[21][9] ,
         \mac_out[21][8] , \mac_out[21][7] , \mac_out[21][6] ,
         \mac_out[21][5] , \mac_out[21][4] , \mac_out[21][3] ,
         \mac_out[21][2] , \mac_out[21][1] , \mac_out[21][0] ,
         \mac_out[20][15] , \mac_out[20][14] , \mac_out[20][13] ,
         \mac_out[20][12] , \mac_out[20][11] , \mac_out[20][10] ,
         \mac_out[20][9] , \mac_out[20][8] , \mac_out[20][7] ,
         \mac_out[20][6] , \mac_out[20][5] , \mac_out[20][4] ,
         \mac_out[20][3] , \mac_out[20][2] , \mac_out[20][1] ,
         \mac_out[20][0] , \mac_out[19][15] , \mac_out[19][14] ,
         \mac_out[19][13] , \mac_out[19][12] , \mac_out[19][11] ,
         \mac_out[19][10] , \mac_out[19][9] , \mac_out[19][8] ,
         \mac_out[19][7] , \mac_out[19][6] , \mac_out[19][5] ,
         \mac_out[19][4] , \mac_out[19][3] , \mac_out[19][2] ,
         \mac_out[19][1] , \mac_out[19][0] , \mac_out[18][15] ,
         \mac_out[18][14] , \mac_out[18][13] , \mac_out[18][12] ,
         \mac_out[18][11] , \mac_out[18][10] , \mac_out[18][9] ,
         \mac_out[18][8] , \mac_out[18][7] , \mac_out[18][6] ,
         \mac_out[18][5] , \mac_out[18][4] , \mac_out[18][3] ,
         \mac_out[18][2] , \mac_out[18][1] , \mac_out[18][0] ,
         \mac_out[17][15] , \mac_out[17][14] , \mac_out[17][13] ,
         \mac_out[17][12] , \mac_out[17][11] , \mac_out[17][10] ,
         \mac_out[17][9] , \mac_out[17][8] , \mac_out[17][7] ,
         \mac_out[17][6] , \mac_out[17][5] , \mac_out[17][4] ,
         \mac_out[17][3] , \mac_out[17][2] , \mac_out[17][1] ,
         \mac_out[17][0] , \mac_out[16][15] , \mac_out[16][14] ,
         \mac_out[16][13] , \mac_out[16][12] , \mac_out[16][11] ,
         \mac_out[16][10] , \mac_out[16][9] , \mac_out[16][8] ,
         \mac_out[16][7] , \mac_out[16][6] , \mac_out[16][5] ,
         \mac_out[16][4] , \mac_out[16][3] , \mac_out[16][2] ,
         \mac_out[16][1] , \mac_out[16][0] , \mac_out[15][15] ,
         \mac_out[15][14] , \mac_out[15][13] , \mac_out[15][12] ,
         \mac_out[15][11] , \mac_out[15][10] , \mac_out[15][9] ,
         \mac_out[15][8] , \mac_out[15][7] , \mac_out[15][6] ,
         \mac_out[15][5] , \mac_out[15][4] , \mac_out[15][3] ,
         \mac_out[15][2] , \mac_out[15][1] , \mac_out[15][0] ,
         \mac_out[14][15] , \mac_out[14][14] , \mac_out[14][13] ,
         \mac_out[14][12] , \mac_out[14][11] , \mac_out[14][10] ,
         \mac_out[14][9] , \mac_out[14][8] , \mac_out[14][7] ,
         \mac_out[14][6] , \mac_out[14][5] , \mac_out[14][4] ,
         \mac_out[14][3] , \mac_out[14][2] , \mac_out[14][1] ,
         \mac_out[14][0] , \mac_out[13][15] , \mac_out[13][14] ,
         \mac_out[13][13] , \mac_out[13][12] , \mac_out[13][11] ,
         \mac_out[13][10] , \mac_out[13][9] , \mac_out[13][8] ,
         \mac_out[13][7] , \mac_out[13][6] , \mac_out[13][5] ,
         \mac_out[13][4] , \mac_out[13][3] , \mac_out[13][2] ,
         \mac_out[13][1] , \mac_out[13][0] , \mac_out[12][15] ,
         \mac_out[12][14] , \mac_out[12][13] , \mac_out[12][12] ,
         \mac_out[12][11] , \mac_out[12][10] , \mac_out[12][9] ,
         \mac_out[12][8] , \mac_out[12][7] , \mac_out[12][6] ,
         \mac_out[12][5] , \mac_out[12][4] , \mac_out[12][3] ,
         \mac_out[12][2] , \mac_out[12][1] , \mac_out[12][0] ,
         \mac_out[11][15] , \mac_out[11][14] , \mac_out[11][13] ,
         \mac_out[11][12] , \mac_out[11][11] , \mac_out[11][10] ,
         \mac_out[11][9] , \mac_out[11][8] , \mac_out[11][7] ,
         \mac_out[11][6] , \mac_out[11][5] , \mac_out[11][4] ,
         \mac_out[11][3] , \mac_out[11][2] , \mac_out[11][1] ,
         \mac_out[11][0] , \mac_out[10][15] , \mac_out[10][14] ,
         \mac_out[10][13] , \mac_out[10][12] , \mac_out[10][11] ,
         \mac_out[10][10] , \mac_out[10][9] , \mac_out[10][8] ,
         \mac_out[10][7] , \mac_out[10][6] , \mac_out[10][5] ,
         \mac_out[10][4] , \mac_out[10][3] , \mac_out[10][2] ,
         \mac_out[10][1] , \mac_out[10][0] , \mac_out[9][15] ,
         \mac_out[9][14] , \mac_out[9][13] , \mac_out[9][12] ,
         \mac_out[9][11] , \mac_out[9][10] , \mac_out[9][9] , \mac_out[9][8] ,
         \mac_out[9][7] , \mac_out[9][6] , \mac_out[9][5] , \mac_out[9][4] ,
         \mac_out[9][3] , \mac_out[9][2] , \mac_out[9][1] , \mac_out[9][0] ,
         \mac_out[8][15] , \mac_out[8][14] , \mac_out[8][13] ,
         \mac_out[8][12] , \mac_out[8][11] , \mac_out[8][10] , \mac_out[8][9] ,
         \mac_out[8][8] , \mac_out[8][7] , \mac_out[8][6] , \mac_out[8][5] ,
         \mac_out[8][4] , \mac_out[8][3] , \mac_out[8][2] , \mac_out[8][1] ,
         \mac_out[8][0] , \mac_out[7][15] , \mac_out[7][14] , \mac_out[7][13] ,
         \mac_out[7][12] , \mac_out[7][11] , \mac_out[7][10] , \mac_out[7][9] ,
         \mac_out[7][8] , \mac_out[7][7] , \mac_out[7][6] , \mac_out[7][5] ,
         \mac_out[7][4] , \mac_out[7][3] , \mac_out[7][2] , \mac_out[7][1] ,
         \mac_out[7][0] , \mac_out[6][15] , \mac_out[6][14] , \mac_out[6][13] ,
         \mac_out[6][12] , \mac_out[6][11] , \mac_out[6][10] , \mac_out[6][9] ,
         \mac_out[6][8] , \mac_out[6][7] , \mac_out[6][6] , \mac_out[6][5] ,
         \mac_out[6][4] , \mac_out[6][3] , \mac_out[6][2] , \mac_out[6][1] ,
         \mac_out[6][0] , \mac_out[5][15] , \mac_out[5][14] , \mac_out[5][13] ,
         \mac_out[5][12] , \mac_out[5][11] , \mac_out[5][10] , \mac_out[5][9] ,
         \mac_out[5][8] , \mac_out[5][7] , \mac_out[5][6] , \mac_out[5][5] ,
         \mac_out[5][4] , \mac_out[5][3] , \mac_out[5][2] , \mac_out[5][1] ,
         \mac_out[5][0] , \mac_out[4][15] , \mac_out[4][14] , \mac_out[4][13] ,
         \mac_out[4][12] , \mac_out[4][11] , \mac_out[4][10] , \mac_out[4][9] ,
         \mac_out[4][8] , \mac_out[4][7] , \mac_out[4][6] , \mac_out[4][5] ,
         \mac_out[4][4] , \mac_out[4][3] , \mac_out[4][2] , \mac_out[4][1] ,
         \mac_out[4][0] , \mac_out[3][15] , \mac_out[3][14] , \mac_out[3][13] ,
         \mac_out[3][12] , \mac_out[3][11] , \mac_out[3][10] , \mac_out[3][9] ,
         \mac_out[3][8] , \mac_out[3][7] , \mac_out[3][6] , \mac_out[3][5] ,
         \mac_out[3][4] , \mac_out[3][3] , \mac_out[3][2] , \mac_out[3][1] ,
         \mac_out[3][0] , \mac_out[2][15] , \mac_out[2][14] , \mac_out[2][13] ,
         \mac_out[2][12] , \mac_out[2][11] , \mac_out[2][10] , \mac_out[2][9] ,
         \mac_out[2][8] , \mac_out[2][7] , \mac_out[2][6] , \mac_out[2][5] ,
         \mac_out[2][4] , \mac_out[2][3] , \mac_out[2][2] , \mac_out[2][1] ,
         \mac_out[2][0] , \mac_out[1][15] , \mac_out[1][14] , \mac_out[1][13] ,
         \mac_out[1][12] , \mac_out[1][11] , \mac_out[1][10] , \mac_out[1][9] ,
         \mac_out[1][8] , \mac_out[1][7] , \mac_out[1][6] , \mac_out[1][5] ,
         \mac_out[1][4] , \mac_out[1][3] , \mac_out[1][2] , \mac_out[1][1] ,
         \mac_out[1][0] , \mac_out[0][15] , \mac_out[0][14] , \mac_out[0][13] ,
         \mac_out[0][12] , \mac_out[0][11] , \mac_out[0][10] , \mac_out[0][9] ,
         \mac_out[0][8] , \mac_out[0][7] , \mac_out[0][6] , \mac_out[0][5] ,
         \mac_out[0][4] , \mac_out[0][3] , \mac_out[0][2] , \mac_out[0][1] ,
         \mac_out[0][0] , \mux[31][15] , \mux[31][14] , \mux[31][13] ,
         \mux[31][12] , \mux[31][11] , \mux[31][10] , \mux[31][9] ,
         \mux[31][8] , \mux[31][7] , \mux[31][6] , \mux[31][5] , \mux[31][4] ,
         \mux[31][3] , \mux[31][2] , \mux[31][1] , \mux[31][0] , \mux[30][15] ,
         \mux[30][14] , \mux[30][13] , \mux[30][12] , \mux[30][11] ,
         \mux[30][10] , \mux[30][9] , \mux[30][8] , \mux[30][7] , \mux[30][6] ,
         \mux[30][5] , \mux[30][4] , \mux[30][3] , \mux[30][2] , \mux[30][1] ,
         \mux[30][0] , \mux[29][15] , \mux[29][14] , \mux[29][13] ,
         \mux[29][12] , \mux[29][11] , \mux[29][10] , \mux[29][9] ,
         \mux[29][8] , \mux[29][7] , \mux[29][6] , \mux[29][5] , \mux[29][4] ,
         \mux[29][3] , \mux[29][2] , \mux[29][1] , \mux[29][0] , \mux[28][15] ,
         \mux[28][14] , \mux[28][13] , \mux[28][12] , \mux[28][11] ,
         \mux[28][10] , \mux[28][9] , \mux[28][8] , \mux[28][7] , \mux[28][6] ,
         \mux[28][5] , \mux[28][4] , \mux[28][3] , \mux[28][2] , \mux[28][1] ,
         \mux[28][0] , \mux[27][15] , \mux[27][14] , \mux[27][13] ,
         \mux[27][12] , \mux[27][11] , \mux[27][10] , \mux[27][9] ,
         \mux[27][8] , \mux[27][7] , \mux[27][6] , \mux[27][5] , \mux[27][4] ,
         \mux[27][3] , \mux[27][2] , \mux[27][1] , \mux[27][0] , \mux[26][15] ,
         \mux[26][14] , \mux[26][13] , \mux[26][12] , \mux[26][11] ,
         \mux[26][10] , \mux[26][9] , \mux[26][8] , \mux[26][7] , \mux[26][6] ,
         \mux[26][5] , \mux[26][4] , \mux[26][3] , \mux[26][2] , \mux[26][1] ,
         \mux[26][0] , \mux[25][15] , \mux[25][14] , \mux[25][13] ,
         \mux[25][12] , \mux[25][11] , \mux[25][10] , \mux[25][9] ,
         \mux[25][8] , \mux[25][7] , \mux[25][6] , \mux[25][5] , \mux[25][4] ,
         \mux[25][3] , \mux[25][2] , \mux[25][1] , \mux[25][0] , \mux[24][15] ,
         \mux[24][14] , \mux[24][13] , \mux[24][12] , \mux[24][11] ,
         \mux[24][10] , \mux[24][9] , \mux[24][8] , \mux[24][7] , \mux[24][6] ,
         \mux[24][5] , \mux[24][4] , \mux[24][3] , \mux[24][2] , \mux[24][1] ,
         \mux[24][0] , \mux[23][15] , \mux[23][14] , \mux[23][13] ,
         \mux[23][12] , \mux[23][11] , \mux[23][10] , \mux[23][9] ,
         \mux[23][8] , \mux[23][7] , \mux[23][6] , \mux[23][5] , \mux[23][4] ,
         \mux[23][3] , \mux[23][2] , \mux[23][1] , \mux[23][0] , \mux[22][15] ,
         \mux[22][14] , \mux[22][13] , \mux[22][12] , \mux[22][11] ,
         \mux[22][10] , \mux[22][9] , \mux[22][8] , \mux[22][7] , \mux[22][6] ,
         \mux[22][5] , \mux[22][4] , \mux[22][3] , \mux[22][2] , \mux[22][1] ,
         \mux[22][0] , \mux[21][15] , \mux[21][14] , \mux[21][13] ,
         \mux[21][12] , \mux[21][11] , \mux[21][10] , \mux[21][9] ,
         \mux[21][8] , \mux[21][7] , \mux[21][6] , \mux[21][5] , \mux[21][4] ,
         \mux[21][3] , \mux[21][2] , \mux[21][1] , \mux[21][0] , \mux[20][15] ,
         \mux[20][14] , \mux[20][13] , \mux[20][12] , \mux[20][11] ,
         \mux[20][10] , \mux[20][9] , \mux[20][8] , \mux[20][7] , \mux[20][6] ,
         \mux[20][5] , \mux[20][4] , \mux[20][3] , \mux[20][2] , \mux[20][1] ,
         \mux[20][0] , \mux[19][15] , \mux[19][14] , \mux[19][13] ,
         \mux[19][12] , \mux[19][11] , \mux[19][10] , \mux[19][9] ,
         \mux[19][8] , \mux[19][7] , \mux[19][6] , \mux[19][5] , \mux[19][4] ,
         \mux[19][3] , \mux[19][2] , \mux[19][1] , \mux[19][0] , \mux[18][15] ,
         \mux[18][14] , \mux[18][13] , \mux[18][12] , \mux[18][11] ,
         \mux[18][10] , \mux[18][9] , \mux[18][8] , \mux[18][7] , \mux[18][6] ,
         \mux[18][5] , \mux[18][4] , \mux[18][3] , \mux[18][2] , \mux[18][1] ,
         \mux[18][0] , \mux[17][15] , \mux[17][14] , \mux[17][13] ,
         \mux[17][12] , \mux[17][11] , \mux[17][10] , \mux[17][9] ,
         \mux[17][8] , \mux[17][7] , \mux[17][6] , \mux[17][5] , \mux[17][4] ,
         \mux[17][3] , \mux[17][2] , \mux[17][1] , \mux[17][0] , \mux[16][15] ,
         \mux[16][14] , \mux[16][13] , \mux[16][12] , \mux[16][11] ,
         \mux[16][10] , \mux[16][9] , \mux[16][8] , \mux[16][7] , \mux[16][6] ,
         \mux[16][5] , \mux[16][4] , \mux[16][3] , \mux[16][2] , \mux[16][1] ,
         \mux[16][0] , \mux[15][15] , \mux[15][14] , \mux[15][13] ,
         \mux[15][12] , \mux[15][11] , \mux[15][10] , \mux[15][9] ,
         \mux[15][8] , \mux[15][7] , \mux[15][6] , \mux[15][5] , \mux[15][4] ,
         \mux[15][3] , \mux[15][2] , \mux[15][1] , \mux[15][0] , \mux[14][15] ,
         \mux[14][14] , \mux[14][13] , \mux[14][12] , \mux[14][11] ,
         \mux[14][10] , \mux[14][9] , \mux[14][8] , \mux[14][7] , \mux[14][6] ,
         \mux[14][5] , \mux[14][4] , \mux[14][3] , \mux[14][2] , \mux[14][1] ,
         \mux[14][0] , \mux[13][15] , \mux[13][14] , \mux[13][13] ,
         \mux[13][12] , \mux[13][11] , \mux[13][10] , \mux[13][9] ,
         \mux[13][8] , \mux[13][7] , \mux[13][6] , \mux[13][5] , \mux[13][4] ,
         \mux[13][3] , \mux[13][2] , \mux[13][1] , \mux[13][0] , \mux[12][15] ,
         \mux[12][14] , \mux[12][13] , \mux[12][12] , \mux[12][11] ,
         \mux[12][10] , \mux[12][9] , \mux[12][8] , \mux[12][7] , \mux[12][6] ,
         \mux[12][5] , \mux[12][4] , \mux[12][3] , \mux[12][2] , \mux[12][1] ,
         \mux[12][0] , \mux[11][15] , \mux[11][14] , \mux[11][13] ,
         \mux[11][12] , \mux[11][11] , \mux[11][10] , \mux[11][9] ,
         \mux[11][8] , \mux[11][7] , \mux[11][6] , \mux[11][5] , \mux[11][4] ,
         \mux[11][3] , \mux[11][2] , \mux[11][1] , \mux[11][0] , \mux[10][15] ,
         \mux[10][14] , \mux[10][13] , \mux[10][12] , \mux[10][11] ,
         \mux[10][10] , \mux[10][9] , \mux[10][8] , \mux[10][7] , \mux[10][6] ,
         \mux[10][5] , \mux[10][4] , \mux[10][3] , \mux[10][2] , \mux[10][1] ,
         \mux[10][0] , \mux[9][15] , \mux[9][14] , \mux[9][13] , \mux[9][12] ,
         \mux[9][11] , \mux[9][10] , \mux[9][9] , \mux[9][8] , \mux[9][7] ,
         \mux[9][6] , \mux[9][5] , \mux[9][4] , \mux[9][3] , \mux[9][2] ,
         \mux[9][1] , \mux[9][0] , \mux[8][15] , \mux[8][14] , \mux[8][13] ,
         \mux[8][12] , \mux[8][11] , \mux[8][10] , \mux[8][9] , \mux[8][8] ,
         \mux[8][7] , \mux[8][6] , \mux[8][5] , \mux[8][4] , \mux[8][3] ,
         \mux[8][2] , \mux[8][1] , \mux[8][0] , \mux[7][15] , \mux[7][14] ,
         \mux[7][13] , \mux[7][12] , \mux[7][11] , \mux[7][10] , \mux[7][9] ,
         \mux[7][8] , \mux[7][7] , \mux[7][6] , \mux[7][5] , \mux[7][4] ,
         \mux[7][3] , \mux[7][2] , \mux[7][1] , \mux[7][0] , \mux[6][15] ,
         \mux[6][14] , \mux[6][13] , \mux[6][12] , \mux[6][11] , \mux[6][10] ,
         \mux[6][9] , \mux[6][8] , \mux[6][7] , \mux[6][6] , \mux[6][5] ,
         \mux[6][4] , \mux[6][3] , \mux[6][2] , \mux[6][1] , \mux[6][0] ,
         \mux[5][15] , \mux[5][14] , \mux[5][13] , \mux[5][12] , \mux[5][11] ,
         \mux[5][10] , \mux[5][9] , \mux[5][8] , \mux[5][7] , \mux[5][6] ,
         \mux[5][5] , \mux[5][4] , \mux[5][3] , \mux[5][2] , \mux[5][1] ,
         \mux[5][0] , \mux[4][15] , \mux[4][14] , \mux[4][13] , \mux[4][12] ,
         \mux[4][11] , \mux[4][10] , \mux[4][9] , \mux[4][8] , \mux[4][7] ,
         \mux[4][6] , \mux[4][5] , \mux[4][4] , \mux[4][3] , \mux[4][2] ,
         \mux[4][1] , \mux[4][0] , \mux[3][15] , \mux[3][14] , \mux[3][13] ,
         \mux[3][12] , \mux[3][11] , \mux[3][10] , \mux[3][9] , \mux[3][8] ,
         \mux[3][7] , \mux[3][6] , \mux[3][5] , \mux[3][4] , \mux[3][3] ,
         \mux[3][2] , \mux[3][1] , \mux[3][0] , \mux[2][15] , \mux[2][14] ,
         \mux[2][13] , \mux[2][12] , \mux[2][11] , \mux[2][10] , \mux[2][9] ,
         \mux[2][8] , \mux[2][7] , \mux[2][6] , \mux[2][5] , \mux[2][4] ,
         \mux[2][3] , \mux[2][2] , \mux[2][1] , \mux[2][0] , \mux[1][15] ,
         \mux[1][14] , \mux[1][13] , \mux[1][12] , \mux[1][11] , \mux[1][10] ,
         \mux[1][9] , \mux[1][8] , \mux[1][7] , \mux[1][6] , \mux[1][5] ,
         \mux[1][4] , \mux[1][3] , \mux[1][2] , \mux[1][1] , \mux[1][0] ,
         \mux[0][15] , \mux[0][14] , \mux[0][13] , \mux[0][12] , \mux[0][11] ,
         \mux[0][10] , \mux[0][9] , \mux[0][8] , \mux[0][7] , \mux[0][6] ,
         \mux[0][5] , \mux[0][4] , \mux[0][3] , \mux[0][2] , \mux[0][1] ,
         \mux[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560;
  wire   [7:0] vector_out;

  memory_WIDTH8_SIZE32_LOGSIZE6_32 \matrix[0]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[0][7] , \matrix_out[0][6] , \matrix_out[0][5] , 
        \matrix_out[0][4] , \matrix_out[0][3] , \matrix_out[0][2] , 
        \matrix_out[0][1] , \matrix_out[0][0] }), .addr({\addr_a[0][5] , 
        \addr_a[0][4] , \addr_a[0][3] , \addr_a[0][2] , \addr_a[0][1] , 
        \addr_a[0][0] }), .wr_en(wr_en_a[0]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_31 \matrix[1]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[1][7] , \matrix_out[1][6] , \matrix_out[1][5] , 
        \matrix_out[1][4] , \matrix_out[1][3] , \matrix_out[1][2] , 
        \matrix_out[1][1] , \matrix_out[1][0] }), .addr({\addr_a[1][5] , 
        \addr_a[1][4] , \addr_a[1][3] , \addr_a[1][2] , \addr_a[1][1] , 
        \addr_a[1][0] }), .wr_en(wr_en_a[1]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_30 \matrix[2]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[2][7] , \matrix_out[2][6] , \matrix_out[2][5] , 
        \matrix_out[2][4] , \matrix_out[2][3] , \matrix_out[2][2] , 
        \matrix_out[2][1] , \matrix_out[2][0] }), .addr({\addr_a[2][5] , 
        \addr_a[2][4] , \addr_a[2][3] , \addr_a[2][2] , \addr_a[2][1] , 
        \addr_a[2][0] }), .wr_en(wr_en_a[2]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_29 \matrix[3]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[3][7] , \matrix_out[3][6] , \matrix_out[3][5] , 
        \matrix_out[3][4] , \matrix_out[3][3] , \matrix_out[3][2] , 
        \matrix_out[3][1] , \matrix_out[3][0] }), .addr({\addr_a[3][5] , 
        \addr_a[3][4] , \addr_a[3][3] , \addr_a[3][2] , \addr_a[3][1] , 
        \addr_a[3][0] }), .wr_en(wr_en_a[3]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_28 \matrix[4]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[4][7] , \matrix_out[4][6] , \matrix_out[4][5] , 
        \matrix_out[4][4] , \matrix_out[4][3] , \matrix_out[4][2] , 
        \matrix_out[4][1] , \matrix_out[4][0] }), .addr({\addr_a[4][5] , 
        \addr_a[4][4] , \addr_a[4][3] , \addr_a[4][2] , \addr_a[4][1] , 
        \addr_a[4][0] }), .wr_en(wr_en_a[4]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_27 \matrix[5]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[5][7] , \matrix_out[5][6] , \matrix_out[5][5] , 
        \matrix_out[5][4] , \matrix_out[5][3] , \matrix_out[5][2] , 
        \matrix_out[5][1] , \matrix_out[5][0] }), .addr({\addr_a[5][5] , 
        \addr_a[5][4] , \addr_a[5][3] , \addr_a[5][2] , \addr_a[5][1] , 
        \addr_a[5][0] }), .wr_en(wr_en_a[5]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_26 \matrix[6]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[6][7] , \matrix_out[6][6] , \matrix_out[6][5] , 
        \matrix_out[6][4] , \matrix_out[6][3] , \matrix_out[6][2] , 
        \matrix_out[6][1] , \matrix_out[6][0] }), .addr({\addr_a[6][5] , 
        \addr_a[6][4] , \addr_a[6][3] , \addr_a[6][2] , \addr_a[6][1] , 
        \addr_a[6][0] }), .wr_en(wr_en_a[6]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_25 \matrix[7]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[7][7] , \matrix_out[7][6] , \matrix_out[7][5] , 
        \matrix_out[7][4] , \matrix_out[7][3] , \matrix_out[7][2] , 
        \matrix_out[7][1] , \matrix_out[7][0] }), .addr({\addr_a[7][5] , 
        \addr_a[7][4] , \addr_a[7][3] , \addr_a[7][2] , \addr_a[7][1] , 
        \addr_a[7][0] }), .wr_en(wr_en_a[7]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_24 \matrix[8]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[8][7] , \matrix_out[8][6] , \matrix_out[8][5] , 
        \matrix_out[8][4] , \matrix_out[8][3] , \matrix_out[8][2] , 
        \matrix_out[8][1] , \matrix_out[8][0] }), .addr({\addr_a[8][5] , 
        \addr_a[8][4] , \addr_a[8][3] , \addr_a[8][2] , \addr_a[8][1] , 
        \addr_a[8][0] }), .wr_en(wr_en_a[8]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_23 \matrix[9]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[9][7] , \matrix_out[9][6] , \matrix_out[9][5] , 
        \matrix_out[9][4] , \matrix_out[9][3] , \matrix_out[9][2] , 
        \matrix_out[9][1] , \matrix_out[9][0] }), .addr({\addr_a[9][5] , 
        \addr_a[9][4] , \addr_a[9][3] , \addr_a[9][2] , \addr_a[9][1] , 
        \addr_a[9][0] }), .wr_en(wr_en_a[9]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_22 \matrix[10]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[10][7] , \matrix_out[10][6] , 
        \matrix_out[10][5] , \matrix_out[10][4] , \matrix_out[10][3] , 
        \matrix_out[10][2] , \matrix_out[10][1] , \matrix_out[10][0] }), 
        .addr({\addr_a[10][5] , \addr_a[10][4] , \addr_a[10][3] , 
        \addr_a[10][2] , \addr_a[10][1] , \addr_a[10][0] }), .wr_en(
        wr_en_a[10]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_21 \matrix[11]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[11][7] , \matrix_out[11][6] , 
        \matrix_out[11][5] , \matrix_out[11][4] , \matrix_out[11][3] , 
        \matrix_out[11][2] , \matrix_out[11][1] , \matrix_out[11][0] }), 
        .addr({\addr_a[11][5] , \addr_a[11][4] , \addr_a[11][3] , 
        \addr_a[11][2] , \addr_a[11][1] , \addr_a[11][0] }), .wr_en(
        wr_en_a[11]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_20 \matrix[12]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[12][7] , \matrix_out[12][6] , 
        \matrix_out[12][5] , \matrix_out[12][4] , \matrix_out[12][3] , 
        \matrix_out[12][2] , \matrix_out[12][1] , \matrix_out[12][0] }), 
        .addr({\addr_a[12][5] , \addr_a[12][4] , \addr_a[12][3] , 
        \addr_a[12][2] , \addr_a[12][1] , \addr_a[12][0] }), .wr_en(
        wr_en_a[12]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_19 \matrix[13]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[13][7] , \matrix_out[13][6] , 
        \matrix_out[13][5] , \matrix_out[13][4] , \matrix_out[13][3] , 
        \matrix_out[13][2] , \matrix_out[13][1] , \matrix_out[13][0] }), 
        .addr({\addr_a[13][5] , \addr_a[13][4] , \addr_a[13][3] , 
        \addr_a[13][2] , \addr_a[13][1] , \addr_a[13][0] }), .wr_en(
        wr_en_a[13]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_18 \matrix[14]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[14][7] , \matrix_out[14][6] , 
        \matrix_out[14][5] , \matrix_out[14][4] , \matrix_out[14][3] , 
        \matrix_out[14][2] , \matrix_out[14][1] , \matrix_out[14][0] }), 
        .addr({\addr_a[14][5] , \addr_a[14][4] , \addr_a[14][3] , 
        \addr_a[14][2] , \addr_a[14][1] , \addr_a[14][0] }), .wr_en(
        wr_en_a[14]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_17 \matrix[15]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[15][7] , \matrix_out[15][6] , 
        \matrix_out[15][5] , \matrix_out[15][4] , \matrix_out[15][3] , 
        \matrix_out[15][2] , \matrix_out[15][1] , \matrix_out[15][0] }), 
        .addr({\addr_a[15][5] , \addr_a[15][4] , \addr_a[15][3] , 
        \addr_a[15][2] , \addr_a[15][1] , \addr_a[15][0] }), .wr_en(
        wr_en_a[15]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_16 \matrix[16]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[16][7] , \matrix_out[16][6] , 
        \matrix_out[16][5] , \matrix_out[16][4] , \matrix_out[16][3] , 
        \matrix_out[16][2] , \matrix_out[16][1] , \matrix_out[16][0] }), 
        .addr({\addr_a[16][5] , \addr_a[16][4] , \addr_a[16][3] , 
        \addr_a[16][2] , \addr_a[16][1] , \addr_a[16][0] }), .wr_en(
        wr_en_a[16]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_15 \matrix[17]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[17][7] , \matrix_out[17][6] , 
        \matrix_out[17][5] , \matrix_out[17][4] , \matrix_out[17][3] , 
        \matrix_out[17][2] , \matrix_out[17][1] , \matrix_out[17][0] }), 
        .addr({\addr_a[17][5] , \addr_a[17][4] , \addr_a[17][3] , 
        \addr_a[17][2] , \addr_a[17][1] , \addr_a[17][0] }), .wr_en(
        wr_en_a[17]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_14 \matrix[18]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[18][7] , \matrix_out[18][6] , 
        \matrix_out[18][5] , \matrix_out[18][4] , \matrix_out[18][3] , 
        \matrix_out[18][2] , \matrix_out[18][1] , \matrix_out[18][0] }), 
        .addr({\addr_a[18][5] , \addr_a[18][4] , \addr_a[18][3] , 
        \addr_a[18][2] , \addr_a[18][1] , \addr_a[18][0] }), .wr_en(
        wr_en_a[18]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_13 \matrix[19]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[19][7] , \matrix_out[19][6] , 
        \matrix_out[19][5] , \matrix_out[19][4] , \matrix_out[19][3] , 
        \matrix_out[19][2] , \matrix_out[19][1] , \matrix_out[19][0] }), 
        .addr({\addr_a[19][5] , \addr_a[19][4] , \addr_a[19][3] , 
        \addr_a[19][2] , \addr_a[19][1] , \addr_a[19][0] }), .wr_en(
        wr_en_a[19]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_12 \matrix[20]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[20][7] , \matrix_out[20][6] , 
        \matrix_out[20][5] , \matrix_out[20][4] , \matrix_out[20][3] , 
        \matrix_out[20][2] , \matrix_out[20][1] , \matrix_out[20][0] }), 
        .addr({\addr_a[20][5] , \addr_a[20][4] , \addr_a[20][3] , 
        \addr_a[20][2] , \addr_a[20][1] , \addr_a[20][0] }), .wr_en(
        wr_en_a[20]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_11 \matrix[21]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[21][7] , \matrix_out[21][6] , 
        \matrix_out[21][5] , \matrix_out[21][4] , \matrix_out[21][3] , 
        \matrix_out[21][2] , \matrix_out[21][1] , \matrix_out[21][0] }), 
        .addr({\addr_a[21][5] , \addr_a[21][4] , \addr_a[21][3] , 
        \addr_a[21][2] , \addr_a[21][1] , \addr_a[21][0] }), .wr_en(
        wr_en_a[21]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_10 \matrix[22]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[22][7] , \matrix_out[22][6] , 
        \matrix_out[22][5] , \matrix_out[22][4] , \matrix_out[22][3] , 
        \matrix_out[22][2] , \matrix_out[22][1] , \matrix_out[22][0] }), 
        .addr({\addr_a[22][5] , \addr_a[22][4] , \addr_a[22][3] , 
        \addr_a[22][2] , \addr_a[22][1] , \addr_a[22][0] }), .wr_en(
        wr_en_a[22]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_9 \matrix[23]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[23][7] , \matrix_out[23][6] , 
        \matrix_out[23][5] , \matrix_out[23][4] , \matrix_out[23][3] , 
        \matrix_out[23][2] , \matrix_out[23][1] , \matrix_out[23][0] }), 
        .addr({\addr_a[23][5] , \addr_a[23][4] , \addr_a[23][3] , 
        \addr_a[23][2] , \addr_a[23][1] , \addr_a[23][0] }), .wr_en(
        wr_en_a[23]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_8 \matrix[24]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[24][7] , \matrix_out[24][6] , 
        \matrix_out[24][5] , \matrix_out[24][4] , \matrix_out[24][3] , 
        \matrix_out[24][2] , \matrix_out[24][1] , \matrix_out[24][0] }), 
        .addr({\addr_a[24][5] , \addr_a[24][4] , \addr_a[24][3] , 
        \addr_a[24][2] , \addr_a[24][1] , \addr_a[24][0] }), .wr_en(
        wr_en_a[24]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_7 \matrix[25]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[25][7] , \matrix_out[25][6] , 
        \matrix_out[25][5] , \matrix_out[25][4] , \matrix_out[25][3] , 
        \matrix_out[25][2] , \matrix_out[25][1] , \matrix_out[25][0] }), 
        .addr({\addr_a[25][5] , \addr_a[25][4] , \addr_a[25][3] , 
        \addr_a[25][2] , \addr_a[25][1] , \addr_a[25][0] }), .wr_en(
        wr_en_a[25]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_6 \matrix[26]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[26][7] , \matrix_out[26][6] , 
        \matrix_out[26][5] , \matrix_out[26][4] , \matrix_out[26][3] , 
        \matrix_out[26][2] , \matrix_out[26][1] , \matrix_out[26][0] }), 
        .addr({\addr_a[26][5] , \addr_a[26][4] , \addr_a[26][3] , 
        \addr_a[26][2] , \addr_a[26][1] , \addr_a[26][0] }), .wr_en(
        wr_en_a[26]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_5 \matrix[27]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[27][7] , \matrix_out[27][6] , 
        \matrix_out[27][5] , \matrix_out[27][4] , \matrix_out[27][3] , 
        \matrix_out[27][2] , \matrix_out[27][1] , \matrix_out[27][0] }), 
        .addr({\addr_a[27][5] , \addr_a[27][4] , \addr_a[27][3] , 
        \addr_a[27][2] , \addr_a[27][1] , \addr_a[27][0] }), .wr_en(
        wr_en_a[27]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_4 \matrix[28]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[28][7] , \matrix_out[28][6] , 
        \matrix_out[28][5] , \matrix_out[28][4] , \matrix_out[28][3] , 
        \matrix_out[28][2] , \matrix_out[28][1] , \matrix_out[28][0] }), 
        .addr({\addr_a[28][5] , \addr_a[28][4] , \addr_a[28][3] , 
        \addr_a[28][2] , \addr_a[28][1] , \addr_a[28][0] }), .wr_en(
        wr_en_a[28]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_3 \matrix[29]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[29][7] , \matrix_out[29][6] , 
        \matrix_out[29][5] , \matrix_out[29][4] , \matrix_out[29][3] , 
        \matrix_out[29][2] , \matrix_out[29][1] , \matrix_out[29][0] }), 
        .addr({\addr_a[29][5] , \addr_a[29][4] , \addr_a[29][3] , 
        \addr_a[29][2] , \addr_a[29][1] , \addr_a[29][0] }), .wr_en(
        wr_en_a[29]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_2 \matrix[30]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[30][7] , \matrix_out[30][6] , 
        \matrix_out[30][5] , \matrix_out[30][4] , \matrix_out[30][3] , 
        \matrix_out[30][2] , \matrix_out[30][1] , \matrix_out[30][0] }), 
        .addr({\addr_a[30][5] , \addr_a[30][4] , \addr_a[30][3] , 
        \addr_a[30][2] , \addr_a[30][1] , \addr_a[30][0] }), .wr_en(
        wr_en_a[30]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_1 \matrix[31]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[31][7] , \matrix_out[31][6] , 
        \matrix_out[31][5] , \matrix_out[31][4] , \matrix_out[31][3] , 
        \matrix_out[31][2] , \matrix_out[31][1] , \matrix_out[31][0] }), 
        .addr({\addr_a[31][5] , \addr_a[31][4] , \addr_a[31][3] , 
        \addr_a[31][2] , \addr_a[31][1] , \addr_a[31][0] }), .wr_en(
        wr_en_a[31]) );
  memory_WIDTH8_SIZE32_LOGSIZE6_0 vector ( .clk(clk), .data_in(data_in), 
        .data_out(vector_out), .addr(addr_x), .wr_en(wr_en_x) );
  mac_31 \mac_mod[0]  ( .clk(clk), .clear_acc(n560), .a({\matrix_out[0][7] , 
        \matrix_out[0][6] , \matrix_out[0][5] , \matrix_out[0][4] , 
        \matrix_out[0][3] , \matrix_out[0][2] , \matrix_out[0][1] , 
        \matrix_out[0][0] }), .b({n556, n553, n1, n548, n545, n14, n529, n535}), .mac_out({\mac_out[0][15] , \mac_out[0][14] , \mac_out[0][13] , 
        \mac_out[0][12] , \mac_out[0][11] , \mac_out[0][10] , \mac_out[0][9] , 
        \mac_out[0][8] , \mac_out[0][7] , \mac_out[0][6] , \mac_out[0][5] , 
        \mac_out[0][4] , \mac_out[0][3] , \mac_out[0][2] , \mac_out[0][1] , 
        \mac_out[0][0] }) );
  mac_30 \mac_mod[1]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[1][7] , \matrix_out[1][6] , \matrix_out[1][5] , 
        \matrix_out[1][4] , \matrix_out[1][3] , \matrix_out[1][2] , 
        \matrix_out[1][1] , \matrix_out[1][0] }), .b({n554, n552, n551, n548, 
        n6, n540, n529, n534}), .mac_out({\mac_out[1][15] , \mac_out[1][14] , 
        \mac_out[1][13] , \mac_out[1][12] , \mac_out[1][11] , \mac_out[1][10] , 
        \mac_out[1][9] , \mac_out[1][8] , \mac_out[1][7] , \mac_out[1][6] , 
        \mac_out[1][5] , \mac_out[1][4] , \mac_out[1][3] , \mac_out[1][2] , 
        \mac_out[1][1] , \mac_out[1][0] }) );
  mac_29 \mac_mod[2]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[2][7] , \matrix_out[2][6] , \matrix_out[2][5] , 
        \matrix_out[2][4] , \matrix_out[2][3] , \matrix_out[2][2] , 
        \matrix_out[2][1] , \matrix_out[2][0] }), .b({n554, n8, n551, n2, n13, 
        n14, n533, n10}), .mac_out({\mac_out[2][15] , \mac_out[2][14] , 
        \mac_out[2][13] , \mac_out[2][12] , \mac_out[2][11] , \mac_out[2][10] , 
        \mac_out[2][9] , \mac_out[2][8] , \mac_out[2][7] , \mac_out[2][6] , 
        \mac_out[2][5] , \mac_out[2][4] , \mac_out[2][3] , \mac_out[2][2] , 
        \mac_out[2][1] , \mac_out[2][0] }) );
  mac_28 \mac_mod[3]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[3][7] , \matrix_out[3][6] , \matrix_out[3][5] , 
        \matrix_out[3][4] , \matrix_out[3][3] , \matrix_out[3][2] , 
        \matrix_out[3][1] , \matrix_out[3][0] }), .b({n554, n7, n551, n9, n12, 
        n4, n528, n535}), .mac_out({\mac_out[3][15] , \mac_out[3][14] , 
        \mac_out[3][13] , \mac_out[3][12] , \mac_out[3][11] , \mac_out[3][10] , 
        \mac_out[3][9] , \mac_out[3][8] , \mac_out[3][7] , \mac_out[3][6] , 
        \mac_out[3][5] , \mac_out[3][4] , \mac_out[3][3] , \mac_out[3][2] , 
        \mac_out[3][1] , \mac_out[3][0] }) );
  mac_27 \mac_mod[4]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[4][7] , \matrix_out[4][6] , \matrix_out[4][5] , 
        \matrix_out[4][4] , \matrix_out[4][3] , \matrix_out[4][2] , 
        \matrix_out[4][1] , \matrix_out[4][0] }), .b({n554, n552, n550, n2, 
        n19, n541, n528, n536}), .mac_out({\mac_out[4][15] , \mac_out[4][14] , 
        \mac_out[4][13] , \mac_out[4][12] , \mac_out[4][11] , \mac_out[4][10] , 
        \mac_out[4][9] , \mac_out[4][8] , \mac_out[4][7] , \mac_out[4][6] , 
        \mac_out[4][5] , \mac_out[4][4] , \mac_out[4][3] , \mac_out[4][2] , 
        \mac_out[4][1] , \mac_out[4][0] }) );
  mac_26 \mac_mod[5]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[5][7] , \matrix_out[5][6] , \matrix_out[5][5] , 
        \matrix_out[5][4] , \matrix_out[5][3] , \matrix_out[5][2] , 
        \matrix_out[5][1] , \matrix_out[5][0] }), .b({n554, n553, n1, n547, 
        n543, n4, n28, n535}), .mac_out({\mac_out[5][15] , \mac_out[5][14] , 
        \mac_out[5][13] , \mac_out[5][12] , \mac_out[5][11] , \mac_out[5][10] , 
        \mac_out[5][9] , \mac_out[5][8] , \mac_out[5][7] , \mac_out[5][6] , 
        \mac_out[5][5] , \mac_out[5][4] , \mac_out[5][3] , \mac_out[5][2] , 
        \mac_out[5][1] , \mac_out[5][0] }) );
  mac_25 \mac_mod[6]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[6][7] , \matrix_out[6][6] , \matrix_out[6][5] , 
        \matrix_out[6][4] , \matrix_out[6][3] , \matrix_out[6][2] , 
        \matrix_out[6][1] , \matrix_out[6][0] }), .b({n554, n7, n550, n546, 
        n545, n5, n531, n535}), .mac_out({\mac_out[6][15] , \mac_out[6][14] , 
        \mac_out[6][13] , \mac_out[6][12] , \mac_out[6][11] , \mac_out[6][10] , 
        \mac_out[6][9] , \mac_out[6][8] , \mac_out[6][7] , \mac_out[6][6] , 
        \mac_out[6][5] , \mac_out[6][4] , \mac_out[6][3] , \mac_out[6][2] , 
        \mac_out[6][1] , \mac_out[6][0] }) );
  mac_24 \mac_mod[7]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[7][7] , \matrix_out[7][6] , \matrix_out[7][5] , 
        \matrix_out[7][4] , \matrix_out[7][3] , \matrix_out[7][2] , 
        \matrix_out[7][1] , \matrix_out[7][0] }), .b({n554, n8, n550, n547, n6, 
        n15, n28, n10}), .mac_out({\mac_out[7][15] , \mac_out[7][14] , 
        \mac_out[7][13] , \mac_out[7][12] , \mac_out[7][11] , \mac_out[7][10] , 
        \mac_out[7][9] , \mac_out[7][8] , \mac_out[7][7] , \mac_out[7][6] , 
        \mac_out[7][5] , \mac_out[7][4] , \mac_out[7][3] , \mac_out[7][2] , 
        \mac_out[7][1] , \mac_out[7][0] }) );
  mac_23 \mac_mod[8]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[8][7] , \matrix_out[8][6] , \matrix_out[8][5] , 
        \matrix_out[8][4] , \matrix_out[8][3] , \matrix_out[8][2] , 
        \matrix_out[8][1] , \matrix_out[8][0] }), .b({n554, n8, n549, n547, 
        n19, n4, n16, n10}), .mac_out({\mac_out[8][15] , \mac_out[8][14] , 
        \mac_out[8][13] , \mac_out[8][12] , \mac_out[8][11] , \mac_out[8][10] , 
        \mac_out[8][9] , \mac_out[8][8] , \mac_out[8][7] , \mac_out[8][6] , 
        \mac_out[8][5] , \mac_out[8][4] , \mac_out[8][3] , \mac_out[8][2] , 
        \mac_out[8][1] , \mac_out[8][0] }) );
  mac_22 \mac_mod[9]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[9][7] , \matrix_out[9][6] , \matrix_out[9][5] , 
        \matrix_out[9][4] , \matrix_out[9][3] , \matrix_out[9][2] , 
        \matrix_out[9][1] , \matrix_out[9][0] }), .b({n554, n7, n549, n9, n20, 
        n15, n21, n10}), .mac_out({\mac_out[9][15] , \mac_out[9][14] , 
        \mac_out[9][13] , \mac_out[9][12] , \mac_out[9][11] , \mac_out[9][10] , 
        \mac_out[9][9] , \mac_out[9][8] , \mac_out[9][7] , \mac_out[9][6] , 
        \mac_out[9][5] , \mac_out[9][4] , \mac_out[9][3] , \mac_out[9][2] , 
        \mac_out[9][1] , \mac_out[9][0] }) );
  mac_21 \mac_mod[10]  ( .clk(clk), .clear_acc(n560), .a({\matrix_out[10][7] , 
        \matrix_out[10][6] , \matrix_out[10][5] , \matrix_out[10][4] , 
        \matrix_out[10][3] , \matrix_out[10][2] , \matrix_out[10][1] , 
        \matrix_out[10][0] }), .b({n554, n553, n550, n546, n543, n26, n25, 
        n536}), .mac_out({\mac_out[10][15] , \mac_out[10][14] , 
        \mac_out[10][13] , \mac_out[10][12] , \mac_out[10][11] , 
        \mac_out[10][10] , \mac_out[10][9] , \mac_out[10][8] , 
        \mac_out[10][7] , \mac_out[10][6] , \mac_out[10][5] , \mac_out[10][4] , 
        \mac_out[10][3] , \mac_out[10][2] , \mac_out[10][1] , \mac_out[10][0] }) );
  mac_20 \mac_mod[11]  ( .clk(clk), .clear_acc(n560), .a({\matrix_out[11][7] , 
        \matrix_out[11][6] , \matrix_out[11][5] , \matrix_out[11][4] , 
        \matrix_out[11][3] , \matrix_out[11][2] , \matrix_out[11][1] , 
        \matrix_out[11][0] }), .b({n554, n8, n550, n548, n6, n542, n532, n10}), 
        .mac_out({\mac_out[11][15] , \mac_out[11][14] , \mac_out[11][13] , 
        \mac_out[11][12] , \mac_out[11][11] , \mac_out[11][10] , 
        \mac_out[11][9] , \mac_out[11][8] , \mac_out[11][7] , \mac_out[11][6] , 
        \mac_out[11][5] , \mac_out[11][4] , \mac_out[11][3] , \mac_out[11][2] , 
        \mac_out[11][1] , \mac_out[11][0] }) );
  mac_19 \mac_mod[12]  ( .clk(clk), .clear_acc(n560), .a({\matrix_out[12][7] , 
        \matrix_out[12][6] , \matrix_out[12][5] , \matrix_out[12][4] , 
        \matrix_out[12][3] , \matrix_out[12][2] , \matrix_out[12][1] , 
        \matrix_out[12][0] }), .b({n554, n8, n550, n9, n19, n5, n16, n10}), 
        .mac_out({\mac_out[12][15] , \mac_out[12][14] , \mac_out[12][13] , 
        \mac_out[12][12] , \mac_out[12][11] , \mac_out[12][10] , 
        \mac_out[12][9] , \mac_out[12][8] , \mac_out[12][7] , \mac_out[12][6] , 
        \mac_out[12][5] , \mac_out[12][4] , \mac_out[12][3] , \mac_out[12][2] , 
        \mac_out[12][1] , \mac_out[12][0] }) );
  mac_18 \mac_mod[13]  ( .clk(clk), .clear_acc(n559), .a({\matrix_out[13][7] , 
        \matrix_out[13][6] , \matrix_out[13][5] , \matrix_out[13][4] , 
        \matrix_out[13][3] , \matrix_out[13][2] , \matrix_out[13][1] , 
        \matrix_out[13][0] }), .b({n555, n8, n1, n547, n19, n17, n24, n534}), 
        .mac_out({\mac_out[13][15] , \mac_out[13][14] , \mac_out[13][13] , 
        \mac_out[13][12] , \mac_out[13][11] , \mac_out[13][10] , 
        \mac_out[13][9] , \mac_out[13][8] , \mac_out[13][7] , \mac_out[13][6] , 
        \mac_out[13][5] , \mac_out[13][4] , \mac_out[13][3] , \mac_out[13][2] , 
        \mac_out[13][1] , \mac_out[13][0] }) );
  mac_17 \mac_mod[14]  ( .clk(clk), .clear_acc(n559), .a({\matrix_out[14][7] , 
        \matrix_out[14][6] , \matrix_out[14][5] , \matrix_out[14][4] , 
        \matrix_out[14][3] , \matrix_out[14][2] , \matrix_out[14][1] , 
        \matrix_out[14][0] }), .b({n555, n553, n550, n2, n19, n540, n530, n10}), .mac_out({\mac_out[14][15] , \mac_out[14][14] , \mac_out[14][13] , 
        \mac_out[14][12] , \mac_out[14][11] , \mac_out[14][10] , 
        \mac_out[14][9] , \mac_out[14][8] , \mac_out[14][7] , \mac_out[14][6] , 
        \mac_out[14][5] , \mac_out[14][4] , \mac_out[14][3] , \mac_out[14][2] , 
        \mac_out[14][1] , \mac_out[14][0] }) );
  mac_16 \mac_mod[15]  ( .clk(clk), .clear_acc(n559), .a({\matrix_out[15][7] , 
        \matrix_out[15][6] , \matrix_out[15][5] , \matrix_out[15][4] , 
        \matrix_out[15][3] , \matrix_out[15][2] , \matrix_out[15][1] , 
        \matrix_out[15][0] }), .b({n555, n552, n550, n547, n6, n18, n531, n10}), .mac_out({\mac_out[15][15] , \mac_out[15][14] , \mac_out[15][13] , 
        \mac_out[15][12] , \mac_out[15][11] , \mac_out[15][10] , 
        \mac_out[15][9] , \mac_out[15][8] , \mac_out[15][7] , \mac_out[15][6] , 
        \mac_out[15][5] , \mac_out[15][4] , \mac_out[15][3] , \mac_out[15][2] , 
        \mac_out[15][1] , \mac_out[15][0] }) );
  mac_15 \mac_mod[16]  ( .clk(clk), .clear_acc(n559), .a({\matrix_out[16][7] , 
        \matrix_out[16][6] , \matrix_out[16][5] , \matrix_out[16][4] , 
        \matrix_out[16][3] , \matrix_out[16][2] , \matrix_out[16][1] , 
        \matrix_out[16][0] }), .b({n555, n7, n549, n546, n545, n542, n23, n536}), .mac_out({\mac_out[16][15] , \mac_out[16][14] , \mac_out[16][13] , 
        \mac_out[16][12] , \mac_out[16][11] , \mac_out[16][10] , 
        \mac_out[16][9] , \mac_out[16][8] , \mac_out[16][7] , \mac_out[16][6] , 
        \mac_out[16][5] , \mac_out[16][4] , \mac_out[16][3] , \mac_out[16][2] , 
        \mac_out[16][1] , \mac_out[16][0] }) );
  mac_14 \mac_mod[17]  ( .clk(clk), .clear_acc(n559), .a({\matrix_out[17][7] , 
        \matrix_out[17][6] , \matrix_out[17][5] , \matrix_out[17][4] , 
        \matrix_out[17][3] , \matrix_out[17][2] , \matrix_out[17][1] , 
        \matrix_out[17][0] }), .b({n555, n552, n549, n548, n543, n26, n532, 
        n534}), .mac_out({\mac_out[17][15] , \mac_out[17][14] , 
        \mac_out[17][13] , \mac_out[17][12] , \mac_out[17][11] , 
        \mac_out[17][10] , \mac_out[17][9] , \mac_out[17][8] , 
        \mac_out[17][7] , \mac_out[17][6] , \mac_out[17][5] , \mac_out[17][4] , 
        \mac_out[17][3] , \mac_out[17][2] , \mac_out[17][1] , \mac_out[17][0] }) );
  mac_13 \mac_mod[18]  ( .clk(clk), .clear_acc(n559), .a({\matrix_out[18][7] , 
        \matrix_out[18][6] , \matrix_out[18][5] , \matrix_out[18][4] , 
        \matrix_out[18][3] , \matrix_out[18][2] , \matrix_out[18][1] , 
        \matrix_out[18][0] }), .b({n555, n7, n549, n2, n13, n541, n533, n536}), 
        .mac_out({\mac_out[18][15] , \mac_out[18][14] , \mac_out[18][13] , 
        \mac_out[18][12] , \mac_out[18][11] , \mac_out[18][10] , 
        \mac_out[18][9] , \mac_out[18][8] , \mac_out[18][7] , \mac_out[18][6] , 
        \mac_out[18][5] , \mac_out[18][4] , \mac_out[18][3] , \mac_out[18][2] , 
        \mac_out[18][1] , \mac_out[18][0] }) );
  mac_12 \mac_mod[19]  ( .clk(clk), .clear_acc(n559), .a({\matrix_out[19][7] , 
        \matrix_out[19][6] , \matrix_out[19][5] , \matrix_out[19][4] , 
        \matrix_out[19][3] , \matrix_out[19][2] , \matrix_out[19][1] , 
        \matrix_out[19][0] }), .b({n555, n552, n551, n546, n543, n17, n24, n10}), .mac_out({\mac_out[19][15] , \mac_out[19][14] , \mac_out[19][13] , 
        \mac_out[19][12] , \mac_out[19][11] , \mac_out[19][10] , 
        \mac_out[19][9] , \mac_out[19][8] , \mac_out[19][7] , \mac_out[19][6] , 
        \mac_out[19][5] , \mac_out[19][4] , \mac_out[19][3] , \mac_out[19][2] , 
        \mac_out[19][1] , \mac_out[19][0] }) );
  mac_11 \mac_mod[20]  ( .clk(clk), .clear_acc(n559), .a({\matrix_out[20][7] , 
        \matrix_out[20][6] , \matrix_out[20][5] , \matrix_out[20][4] , 
        \matrix_out[20][3] , \matrix_out[20][2] , \matrix_out[20][1] , 
        \matrix_out[20][0] }), .b({n555, n8, n550, n546, n12, n26, n533, n10}), 
        .mac_out({\mac_out[20][15] , \mac_out[20][14] , \mac_out[20][13] , 
        \mac_out[20][12] , \mac_out[20][11] , \mac_out[20][10] , 
        \mac_out[20][9] , \mac_out[20][8] , \mac_out[20][7] , \mac_out[20][6] , 
        \mac_out[20][5] , \mac_out[20][4] , \mac_out[20][3] , \mac_out[20][2] , 
        \mac_out[20][1] , \mac_out[20][0] }) );
  mac_10 \mac_mod[21]  ( .clk(clk), .clear_acc(n559), .a({\matrix_out[21][7] , 
        \matrix_out[21][6] , \matrix_out[21][5] , \matrix_out[21][4] , 
        \matrix_out[21][3] , \matrix_out[21][2] , \matrix_out[21][1] , 
        \matrix_out[21][0] }), .b({n555, n8, n1, n3, n11, n18, n21, n536}), 
        .mac_out({\mac_out[21][15] , \mac_out[21][14] , \mac_out[21][13] , 
        \mac_out[21][12] , \mac_out[21][11] , \mac_out[21][10] , 
        \mac_out[21][9] , \mac_out[21][8] , \mac_out[21][7] , \mac_out[21][6] , 
        \mac_out[21][5] , \mac_out[21][4] , \mac_out[21][3] , \mac_out[21][2] , 
        \mac_out[21][1] , \mac_out[21][0] }) );
  mac_9 \mac_mod[22]  ( .clk(clk), .clear_acc(n559), .a({\matrix_out[22][7] , 
        \matrix_out[22][6] , \matrix_out[22][5] , \matrix_out[22][4] , 
        \matrix_out[22][3] , \matrix_out[22][2] , \matrix_out[22][1] , 
        \matrix_out[22][0] }), .b({n555, n553, n1, n3, n20, n18, n23, n535}), 
        .mac_out({\mac_out[22][15] , \mac_out[22][14] , \mac_out[22][13] , 
        \mac_out[22][12] , \mac_out[22][11] , \mac_out[22][10] , 
        \mac_out[22][9] , \mac_out[22][8] , \mac_out[22][7] , \mac_out[22][6] , 
        \mac_out[22][5] , \mac_out[22][4] , \mac_out[22][3] , \mac_out[22][2] , 
        \mac_out[22][1] , \mac_out[22][0] }) );
  mac_8 \mac_mod[23]  ( .clk(clk), .clear_acc(n559), .a({\matrix_out[23][7] , 
        \matrix_out[23][6] , \matrix_out[23][5] , \matrix_out[23][4] , 
        \matrix_out[23][3] , \matrix_out[23][2] , \matrix_out[23][1] , 
        \matrix_out[23][0] }), .b({n555, n8, n551, n9, n543, n17, n22, n536}), 
        .mac_out({\mac_out[23][15] , \mac_out[23][14] , \mac_out[23][13] , 
        \mac_out[23][12] , \mac_out[23][11] , \mac_out[23][10] , 
        \mac_out[23][9] , \mac_out[23][8] , \mac_out[23][7] , \mac_out[23][6] , 
        \mac_out[23][5] , \mac_out[23][4] , \mac_out[23][3] , \mac_out[23][2] , 
        \mac_out[23][1] , \mac_out[23][0] }) );
  mac_7 \mac_mod[24]  ( .clk(clk), .clear_acc(n559), .a({\matrix_out[24][7] , 
        \matrix_out[24][6] , \matrix_out[24][5] , \matrix_out[24][4] , 
        \matrix_out[24][3] , \matrix_out[24][2] , \matrix_out[24][1] , 
        \matrix_out[24][0] }), .b({n555, n553, n549, n3, n12, n15, n27, n535}), 
        .mac_out({\mac_out[24][15] , \mac_out[24][14] , \mac_out[24][13] , 
        \mac_out[24][12] , \mac_out[24][11] , \mac_out[24][10] , 
        \mac_out[24][9] , \mac_out[24][8] , \mac_out[24][7] , \mac_out[24][6] , 
        \mac_out[24][5] , \mac_out[24][4] , \mac_out[24][3] , \mac_out[24][2] , 
        \mac_out[24][1] , \mac_out[24][0] }) );
  mac_6 \mac_mod[25]  ( .clk(clk), .clear_acc(n560), .a({\matrix_out[25][7] , 
        \matrix_out[25][6] , \matrix_out[25][5] , \matrix_out[25][4] , 
        \matrix_out[25][3] , \matrix_out[25][2] , \matrix_out[25][1] , 
        \matrix_out[25][0] }), .b({n556, n7, n1, n2, n545, n541, n531, n535}), 
        .mac_out({\mac_out[25][15] , \mac_out[25][14] , \mac_out[25][13] , 
        \mac_out[25][12] , \mac_out[25][11] , \mac_out[25][10] , 
        \mac_out[25][9] , \mac_out[25][8] , \mac_out[25][7] , \mac_out[25][6] , 
        \mac_out[25][5] , \mac_out[25][4] , \mac_out[25][3] , \mac_out[25][2] , 
        \mac_out[25][1] , \mac_out[25][0] }) );
  mac_5 \mac_mod[26]  ( .clk(clk), .clear_acc(n560), .a({\matrix_out[26][7] , 
        \matrix_out[26][6] , \matrix_out[26][5] , \matrix_out[26][4] , 
        \matrix_out[26][3] , \matrix_out[26][2] , \matrix_out[26][1] , 
        \matrix_out[26][0] }), .b({n556, n553, n1, n3, n13, n15, n27, n534}), 
        .mac_out({\mac_out[26][15] , \mac_out[26][14] , \mac_out[26][13] , 
        \mac_out[26][12] , \mac_out[26][11] , \mac_out[26][10] , 
        \mac_out[26][9] , \mac_out[26][8] , \mac_out[26][7] , \mac_out[26][6] , 
        \mac_out[26][5] , \mac_out[26][4] , \mac_out[26][3] , \mac_out[26][2] , 
        \mac_out[26][1] , \mac_out[26][0] }) );
  mac_4 \mac_mod[27]  ( .clk(clk), .clear_acc(n560), .a({\matrix_out[27][7] , 
        \matrix_out[27][6] , \matrix_out[27][5] , \matrix_out[27][4] , 
        \matrix_out[27][3] , \matrix_out[27][2] , \matrix_out[27][1] , 
        \matrix_out[27][0] }), .b({n556, n552, n1, n3, n20, n14, n528, n536}), 
        .mac_out({\mac_out[27][15] , \mac_out[27][14] , \mac_out[27][13] , 
        \mac_out[27][12] , \mac_out[27][11] , \mac_out[27][10] , 
        \mac_out[27][9] , \mac_out[27][8] , \mac_out[27][7] , \mac_out[27][6] , 
        \mac_out[27][5] , \mac_out[27][4] , \mac_out[27][3] , \mac_out[27][2] , 
        \mac_out[27][1] , \mac_out[27][0] }) );
  mac_3 \mac_mod[28]  ( .clk(clk), .clear_acc(n560), .a({\matrix_out[28][7] , 
        \matrix_out[28][6] , \matrix_out[28][5] , \matrix_out[28][4] , 
        \matrix_out[28][3] , \matrix_out[28][2] , \matrix_out[28][1] , 
        \matrix_out[28][0] }), .b({n556, n553, n1, n548, n545, n542, n529, 
        n536}), .mac_out({\mac_out[28][15] , \mac_out[28][14] , 
        \mac_out[28][13] , \mac_out[28][12] , \mac_out[28][11] , 
        \mac_out[28][10] , \mac_out[28][9] , \mac_out[28][8] , 
        \mac_out[28][7] , \mac_out[28][6] , \mac_out[28][5] , \mac_out[28][4] , 
        \mac_out[28][3] , \mac_out[28][2] , \mac_out[28][1] , \mac_out[28][0] }) );
  mac_2 \mac_mod[29]  ( .clk(clk), .clear_acc(n560), .a({\matrix_out[29][7] , 
        \matrix_out[29][6] , \matrix_out[29][5] , \matrix_out[29][4] , 
        \matrix_out[29][3] , \matrix_out[29][2] , \matrix_out[29][1] , 
        \matrix_out[29][0] }), .b({n556, n552, n551, n547, n20, n5, n530, n536}), .mac_out({\mac_out[29][15] , \mac_out[29][14] , \mac_out[29][13] , 
        \mac_out[29][12] , \mac_out[29][11] , \mac_out[29][10] , 
        \mac_out[29][9] , \mac_out[29][8] , \mac_out[29][7] , \mac_out[29][6] , 
        \mac_out[29][5] , \mac_out[29][4] , \mac_out[29][3] , \mac_out[29][2] , 
        \mac_out[29][1] , \mac_out[29][0] }) );
  mac_1 \mac_mod[30]  ( .clk(clk), .clear_acc(n560), .a({\matrix_out[30][7] , 
        \matrix_out[30][6] , \matrix_out[30][5] , \matrix_out[30][4] , 
        \matrix_out[30][3] , \matrix_out[30][2] , \matrix_out[30][1] , 
        \matrix_out[30][0] }), .b({n556, n7, n549, n548, n6, n540, n27, n534}), 
        .mac_out({\mac_out[30][15] , \mac_out[30][14] , \mac_out[30][13] , 
        \mac_out[30][12] , \mac_out[30][11] , \mac_out[30][10] , 
        \mac_out[30][9] , \mac_out[30][8] , \mac_out[30][7] , \mac_out[30][6] , 
        \mac_out[30][5] , \mac_out[30][4] , \mac_out[30][3] , \mac_out[30][2] , 
        \mac_out[30][1] , \mac_out[30][0] }) );
  mac_0 \mac_mod[31]  ( .clk(clk), .clear_acc(n560), .a({\matrix_out[31][7] , 
        \matrix_out[31][6] , \matrix_out[31][5] , \matrix_out[31][4] , 
        \matrix_out[31][3] , \matrix_out[31][2] , \matrix_out[31][1] , 
        \matrix_out[31][0] }), .b({n556, n7, n549, n2, n543, n542, n16, n535}), 
        .mac_out({\mac_out[31][15] , \mac_out[31][14] , \mac_out[31][13] , 
        \mac_out[31][12] , \mac_out[31][11] , \mac_out[31][10] , 
        \mac_out[31][9] , \mac_out[31][8] , \mac_out[31][7] , \mac_out[31][6] , 
        \mac_out[31][5] , \mac_out[31][4] , \mac_out[31][3] , \mac_out[31][2] , 
        \mac_out[31][1] , \mac_out[31][0] }) );
  memory_WIDTH16_SIZE1_LOGSIZE6_31 \y[0]  ( .clk(clk), .data_in({
        \mac_out[0][15] , \mac_out[0][14] , \mac_out[0][13] , \mac_out[0][12] , 
        \mac_out[0][11] , \mac_out[0][10] , \mac_out[0][9] , \mac_out[0][8] , 
        \mac_out[0][7] , \mac_out[0][6] , \mac_out[0][5] , \mac_out[0][4] , 
        \mac_out[0][3] , \mac_out[0][2] , \mac_out[0][1] , \mac_out[0][0] }), 
        .data_out({\mux[0][15] , \mux[0][14] , \mux[0][13] , \mux[0][12] , 
        \mux[0][11] , \mux[0][10] , \mux[0][9] , \mux[0][8] , \mux[0][7] , 
        \mux[0][6] , \mux[0][5] , \mux[0][4] , \mux[0][3] , \mux[0][2] , 
        \mux[0][1] , \mux[0][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_30 \y[1]  ( .clk(clk), .data_in({
        \mac_out[1][15] , \mac_out[1][14] , \mac_out[1][13] , \mac_out[1][12] , 
        \mac_out[1][11] , \mac_out[1][10] , \mac_out[1][9] , \mac_out[1][8] , 
        \mac_out[1][7] , \mac_out[1][6] , \mac_out[1][5] , \mac_out[1][4] , 
        \mac_out[1][3] , \mac_out[1][2] , \mac_out[1][1] , \mac_out[1][0] }), 
        .data_out({\mux[1][15] , \mux[1][14] , \mux[1][13] , \mux[1][12] , 
        \mux[1][11] , \mux[1][10] , \mux[1][9] , \mux[1][8] , \mux[1][7] , 
        \mux[1][6] , \mux[1][5] , \mux[1][4] , \mux[1][3] , \mux[1][2] , 
        \mux[1][1] , \mux[1][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_29 \y[2]  ( .clk(clk), .data_in({
        \mac_out[2][15] , \mac_out[2][14] , \mac_out[2][13] , \mac_out[2][12] , 
        \mac_out[2][11] , \mac_out[2][10] , \mac_out[2][9] , \mac_out[2][8] , 
        \mac_out[2][7] , \mac_out[2][6] , \mac_out[2][5] , \mac_out[2][4] , 
        \mac_out[2][3] , \mac_out[2][2] , \mac_out[2][1] , \mac_out[2][0] }), 
        .data_out({\mux[2][15] , \mux[2][14] , \mux[2][13] , \mux[2][12] , 
        \mux[2][11] , \mux[2][10] , \mux[2][9] , \mux[2][8] , \mux[2][7] , 
        \mux[2][6] , \mux[2][5] , \mux[2][4] , \mux[2][3] , \mux[2][2] , 
        \mux[2][1] , \mux[2][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_28 \y[3]  ( .clk(clk), .data_in({
        \mac_out[3][15] , \mac_out[3][14] , \mac_out[3][13] , \mac_out[3][12] , 
        \mac_out[3][11] , \mac_out[3][10] , \mac_out[3][9] , \mac_out[3][8] , 
        \mac_out[3][7] , \mac_out[3][6] , \mac_out[3][5] , \mac_out[3][4] , 
        \mac_out[3][3] , \mac_out[3][2] , \mac_out[3][1] , \mac_out[3][0] }), 
        .data_out({\mux[3][15] , \mux[3][14] , \mux[3][13] , \mux[3][12] , 
        \mux[3][11] , \mux[3][10] , \mux[3][9] , \mux[3][8] , \mux[3][7] , 
        \mux[3][6] , \mux[3][5] , \mux[3][4] , \mux[3][3] , \mux[3][2] , 
        \mux[3][1] , \mux[3][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_27 \y[4]  ( .clk(clk), .data_in({
        \mac_out[4][15] , \mac_out[4][14] , \mac_out[4][13] , \mac_out[4][12] , 
        \mac_out[4][11] , \mac_out[4][10] , \mac_out[4][9] , \mac_out[4][8] , 
        \mac_out[4][7] , \mac_out[4][6] , \mac_out[4][5] , \mac_out[4][4] , 
        \mac_out[4][3] , \mac_out[4][2] , \mac_out[4][1] , \mac_out[4][0] }), 
        .data_out({\mux[4][15] , \mux[4][14] , \mux[4][13] , \mux[4][12] , 
        \mux[4][11] , \mux[4][10] , \mux[4][9] , \mux[4][8] , \mux[4][7] , 
        \mux[4][6] , \mux[4][5] , \mux[4][4] , \mux[4][3] , \mux[4][2] , 
        \mux[4][1] , \mux[4][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_26 \y[5]  ( .clk(clk), .data_in({
        \mac_out[5][15] , \mac_out[5][14] , \mac_out[5][13] , \mac_out[5][12] , 
        \mac_out[5][11] , \mac_out[5][10] , \mac_out[5][9] , \mac_out[5][8] , 
        \mac_out[5][7] , \mac_out[5][6] , \mac_out[5][5] , \mac_out[5][4] , 
        \mac_out[5][3] , \mac_out[5][2] , \mac_out[5][1] , \mac_out[5][0] }), 
        .data_out({\mux[5][15] , \mux[5][14] , \mux[5][13] , \mux[5][12] , 
        \mux[5][11] , \mux[5][10] , \mux[5][9] , \mux[5][8] , \mux[5][7] , 
        \mux[5][6] , \mux[5][5] , \mux[5][4] , \mux[5][3] , \mux[5][2] , 
        \mux[5][1] , \mux[5][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_25 \y[6]  ( .clk(clk), .data_in({
        \mac_out[6][15] , \mac_out[6][14] , \mac_out[6][13] , \mac_out[6][12] , 
        \mac_out[6][11] , \mac_out[6][10] , \mac_out[6][9] , \mac_out[6][8] , 
        \mac_out[6][7] , \mac_out[6][6] , \mac_out[6][5] , \mac_out[6][4] , 
        \mac_out[6][3] , \mac_out[6][2] , \mac_out[6][1] , \mac_out[6][0] }), 
        .data_out({\mux[6][15] , \mux[6][14] , \mux[6][13] , \mux[6][12] , 
        \mux[6][11] , \mux[6][10] , \mux[6][9] , \mux[6][8] , \mux[6][7] , 
        \mux[6][6] , \mux[6][5] , \mux[6][4] , \mux[6][3] , \mux[6][2] , 
        \mux[6][1] , \mux[6][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_24 \y[7]  ( .clk(clk), .data_in({
        \mac_out[7][15] , \mac_out[7][14] , \mac_out[7][13] , \mac_out[7][12] , 
        \mac_out[7][11] , \mac_out[7][10] , \mac_out[7][9] , \mac_out[7][8] , 
        \mac_out[7][7] , \mac_out[7][6] , \mac_out[7][5] , \mac_out[7][4] , 
        \mac_out[7][3] , \mac_out[7][2] , \mac_out[7][1] , \mac_out[7][0] }), 
        .data_out({\mux[7][15] , \mux[7][14] , \mux[7][13] , \mux[7][12] , 
        \mux[7][11] , \mux[7][10] , \mux[7][9] , \mux[7][8] , \mux[7][7] , 
        \mux[7][6] , \mux[7][5] , \mux[7][4] , \mux[7][3] , \mux[7][2] , 
        \mux[7][1] , \mux[7][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_23 \y[8]  ( .clk(clk), .data_in({
        \mac_out[8][15] , \mac_out[8][14] , \mac_out[8][13] , \mac_out[8][12] , 
        \mac_out[8][11] , \mac_out[8][10] , \mac_out[8][9] , \mac_out[8][8] , 
        \mac_out[8][7] , \mac_out[8][6] , \mac_out[8][5] , \mac_out[8][4] , 
        \mac_out[8][3] , \mac_out[8][2] , \mac_out[8][1] , \mac_out[8][0] }), 
        .data_out({\mux[8][15] , \mux[8][14] , \mux[8][13] , \mux[8][12] , 
        \mux[8][11] , \mux[8][10] , \mux[8][9] , \mux[8][8] , \mux[8][7] , 
        \mux[8][6] , \mux[8][5] , \mux[8][4] , \mux[8][3] , \mux[8][2] , 
        \mux[8][1] , \mux[8][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_22 \y[9]  ( .clk(clk), .data_in({
        \mac_out[9][15] , \mac_out[9][14] , \mac_out[9][13] , \mac_out[9][12] , 
        \mac_out[9][11] , \mac_out[9][10] , \mac_out[9][9] , \mac_out[9][8] , 
        \mac_out[9][7] , \mac_out[9][6] , \mac_out[9][5] , \mac_out[9][4] , 
        \mac_out[9][3] , \mac_out[9][2] , \mac_out[9][1] , \mac_out[9][0] }), 
        .data_out({\mux[9][15] , \mux[9][14] , \mux[9][13] , \mux[9][12] , 
        \mux[9][11] , \mux[9][10] , \mux[9][9] , \mux[9][8] , \mux[9][7] , 
        \mux[9][6] , \mux[9][5] , \mux[9][4] , \mux[9][3] , \mux[9][2] , 
        \mux[9][1] , \mux[9][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_21 \y[10]  ( .clk(clk), .data_in({
        \mac_out[10][15] , \mac_out[10][14] , \mac_out[10][13] , 
        \mac_out[10][12] , \mac_out[10][11] , \mac_out[10][10] , 
        \mac_out[10][9] , \mac_out[10][8] , \mac_out[10][7] , \mac_out[10][6] , 
        \mac_out[10][5] , \mac_out[10][4] , \mac_out[10][3] , \mac_out[10][2] , 
        \mac_out[10][1] , \mac_out[10][0] }), .data_out({\mux[10][15] , 
        \mux[10][14] , \mux[10][13] , \mux[10][12] , \mux[10][11] , 
        \mux[10][10] , \mux[10][9] , \mux[10][8] , \mux[10][7] , \mux[10][6] , 
        \mux[10][5] , \mux[10][4] , \mux[10][3] , \mux[10][2] , \mux[10][1] , 
        \mux[10][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_20 \y[11]  ( .clk(clk), .data_in({
        \mac_out[11][15] , \mac_out[11][14] , \mac_out[11][13] , 
        \mac_out[11][12] , \mac_out[11][11] , \mac_out[11][10] , 
        \mac_out[11][9] , \mac_out[11][8] , \mac_out[11][7] , \mac_out[11][6] , 
        \mac_out[11][5] , \mac_out[11][4] , \mac_out[11][3] , \mac_out[11][2] , 
        \mac_out[11][1] , \mac_out[11][0] }), .data_out({\mux[11][15] , 
        \mux[11][14] , \mux[11][13] , \mux[11][12] , \mux[11][11] , 
        \mux[11][10] , \mux[11][9] , \mux[11][8] , \mux[11][7] , \mux[11][6] , 
        \mux[11][5] , \mux[11][4] , \mux[11][3] , \mux[11][2] , \mux[11][1] , 
        \mux[11][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_19 \y[12]  ( .clk(clk), .data_in({
        \mac_out[12][15] , \mac_out[12][14] , \mac_out[12][13] , 
        \mac_out[12][12] , \mac_out[12][11] , \mac_out[12][10] , 
        \mac_out[12][9] , \mac_out[12][8] , \mac_out[12][7] , \mac_out[12][6] , 
        \mac_out[12][5] , \mac_out[12][4] , \mac_out[12][3] , \mac_out[12][2] , 
        \mac_out[12][1] , \mac_out[12][0] }), .data_out({\mux[12][15] , 
        \mux[12][14] , \mux[12][13] , \mux[12][12] , \mux[12][11] , 
        \mux[12][10] , \mux[12][9] , \mux[12][8] , \mux[12][7] , \mux[12][6] , 
        \mux[12][5] , \mux[12][4] , \mux[12][3] , \mux[12][2] , \mux[12][1] , 
        \mux[12][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_18 \y[13]  ( .clk(clk), .data_in({
        \mac_out[13][15] , \mac_out[13][14] , \mac_out[13][13] , 
        \mac_out[13][12] , \mac_out[13][11] , \mac_out[13][10] , 
        \mac_out[13][9] , \mac_out[13][8] , \mac_out[13][7] , \mac_out[13][6] , 
        \mac_out[13][5] , \mac_out[13][4] , \mac_out[13][3] , \mac_out[13][2] , 
        \mac_out[13][1] , \mac_out[13][0] }), .data_out({\mux[13][15] , 
        \mux[13][14] , \mux[13][13] , \mux[13][12] , \mux[13][11] , 
        \mux[13][10] , \mux[13][9] , \mux[13][8] , \mux[13][7] , \mux[13][6] , 
        \mux[13][5] , \mux[13][4] , \mux[13][3] , \mux[13][2] , \mux[13][1] , 
        \mux[13][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_17 \y[14]  ( .clk(clk), .data_in({
        \mac_out[14][15] , \mac_out[14][14] , \mac_out[14][13] , 
        \mac_out[14][12] , \mac_out[14][11] , \mac_out[14][10] , 
        \mac_out[14][9] , \mac_out[14][8] , \mac_out[14][7] , \mac_out[14][6] , 
        \mac_out[14][5] , \mac_out[14][4] , \mac_out[14][3] , \mac_out[14][2] , 
        \mac_out[14][1] , \mac_out[14][0] }), .data_out({\mux[14][15] , 
        \mux[14][14] , \mux[14][13] , \mux[14][12] , \mux[14][11] , 
        \mux[14][10] , \mux[14][9] , \mux[14][8] , \mux[14][7] , \mux[14][6] , 
        \mux[14][5] , \mux[14][4] , \mux[14][3] , \mux[14][2] , \mux[14][1] , 
        \mux[14][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_16 \y[15]  ( .clk(clk), .data_in({
        \mac_out[15][15] , \mac_out[15][14] , \mac_out[15][13] , 
        \mac_out[15][12] , \mac_out[15][11] , \mac_out[15][10] , 
        \mac_out[15][9] , \mac_out[15][8] , \mac_out[15][7] , \mac_out[15][6] , 
        \mac_out[15][5] , \mac_out[15][4] , \mac_out[15][3] , \mac_out[15][2] , 
        \mac_out[15][1] , \mac_out[15][0] }), .data_out({\mux[15][15] , 
        \mux[15][14] , \mux[15][13] , \mux[15][12] , \mux[15][11] , 
        \mux[15][10] , \mux[15][9] , \mux[15][8] , \mux[15][7] , \mux[15][6] , 
        \mux[15][5] , \mux[15][4] , \mux[15][3] , \mux[15][2] , \mux[15][1] , 
        \mux[15][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_15 \y[16]  ( .clk(clk), .data_in({
        \mac_out[16][15] , \mac_out[16][14] , \mac_out[16][13] , 
        \mac_out[16][12] , \mac_out[16][11] , \mac_out[16][10] , 
        \mac_out[16][9] , \mac_out[16][8] , \mac_out[16][7] , \mac_out[16][6] , 
        \mac_out[16][5] , \mac_out[16][4] , \mac_out[16][3] , \mac_out[16][2] , 
        \mac_out[16][1] , \mac_out[16][0] }), .data_out({\mux[16][15] , 
        \mux[16][14] , \mux[16][13] , \mux[16][12] , \mux[16][11] , 
        \mux[16][10] , \mux[16][9] , \mux[16][8] , \mux[16][7] , \mux[16][6] , 
        \mux[16][5] , \mux[16][4] , \mux[16][3] , \mux[16][2] , \mux[16][1] , 
        \mux[16][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_14 \y[17]  ( .clk(clk), .data_in({
        \mac_out[17][15] , \mac_out[17][14] , \mac_out[17][13] , 
        \mac_out[17][12] , \mac_out[17][11] , \mac_out[17][10] , 
        \mac_out[17][9] , \mac_out[17][8] , \mac_out[17][7] , \mac_out[17][6] , 
        \mac_out[17][5] , \mac_out[17][4] , \mac_out[17][3] , \mac_out[17][2] , 
        \mac_out[17][1] , \mac_out[17][0] }), .data_out({\mux[17][15] , 
        \mux[17][14] , \mux[17][13] , \mux[17][12] , \mux[17][11] , 
        \mux[17][10] , \mux[17][9] , \mux[17][8] , \mux[17][7] , \mux[17][6] , 
        \mux[17][5] , \mux[17][4] , \mux[17][3] , \mux[17][2] , \mux[17][1] , 
        \mux[17][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_13 \y[18]  ( .clk(clk), .data_in({
        \mac_out[18][15] , \mac_out[18][14] , \mac_out[18][13] , 
        \mac_out[18][12] , \mac_out[18][11] , \mac_out[18][10] , 
        \mac_out[18][9] , \mac_out[18][8] , \mac_out[18][7] , \mac_out[18][6] , 
        \mac_out[18][5] , \mac_out[18][4] , \mac_out[18][3] , \mac_out[18][2] , 
        \mac_out[18][1] , \mac_out[18][0] }), .data_out({\mux[18][15] , 
        \mux[18][14] , \mux[18][13] , \mux[18][12] , \mux[18][11] , 
        \mux[18][10] , \mux[18][9] , \mux[18][8] , \mux[18][7] , \mux[18][6] , 
        \mux[18][5] , \mux[18][4] , \mux[18][3] , \mux[18][2] , \mux[18][1] , 
        \mux[18][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_12 \y[19]  ( .clk(clk), .data_in({
        \mac_out[19][15] , \mac_out[19][14] , \mac_out[19][13] , 
        \mac_out[19][12] , \mac_out[19][11] , \mac_out[19][10] , 
        \mac_out[19][9] , \mac_out[19][8] , \mac_out[19][7] , \mac_out[19][6] , 
        \mac_out[19][5] , \mac_out[19][4] , \mac_out[19][3] , \mac_out[19][2] , 
        \mac_out[19][1] , \mac_out[19][0] }), .data_out({\mux[19][15] , 
        \mux[19][14] , \mux[19][13] , \mux[19][12] , \mux[19][11] , 
        \mux[19][10] , \mux[19][9] , \mux[19][8] , \mux[19][7] , \mux[19][6] , 
        \mux[19][5] , \mux[19][4] , \mux[19][3] , \mux[19][2] , \mux[19][1] , 
        \mux[19][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_11 \y[20]  ( .clk(clk), .data_in({
        \mac_out[20][15] , \mac_out[20][14] , \mac_out[20][13] , 
        \mac_out[20][12] , \mac_out[20][11] , \mac_out[20][10] , 
        \mac_out[20][9] , \mac_out[20][8] , \mac_out[20][7] , \mac_out[20][6] , 
        \mac_out[20][5] , \mac_out[20][4] , \mac_out[20][3] , \mac_out[20][2] , 
        \mac_out[20][1] , \mac_out[20][0] }), .data_out({\mux[20][15] , 
        \mux[20][14] , \mux[20][13] , \mux[20][12] , \mux[20][11] , 
        \mux[20][10] , \mux[20][9] , \mux[20][8] , \mux[20][7] , \mux[20][6] , 
        \mux[20][5] , \mux[20][4] , \mux[20][3] , \mux[20][2] , \mux[20][1] , 
        \mux[20][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_10 \y[21]  ( .clk(clk), .data_in({
        \mac_out[21][15] , \mac_out[21][14] , \mac_out[21][13] , 
        \mac_out[21][12] , \mac_out[21][11] , \mac_out[21][10] , 
        \mac_out[21][9] , \mac_out[21][8] , \mac_out[21][7] , \mac_out[21][6] , 
        \mac_out[21][5] , \mac_out[21][4] , \mac_out[21][3] , \mac_out[21][2] , 
        \mac_out[21][1] , \mac_out[21][0] }), .data_out({\mux[21][15] , 
        \mux[21][14] , \mux[21][13] , \mux[21][12] , \mux[21][11] , 
        \mux[21][10] , \mux[21][9] , \mux[21][8] , \mux[21][7] , \mux[21][6] , 
        \mux[21][5] , \mux[21][4] , \mux[21][3] , \mux[21][2] , \mux[21][1] , 
        \mux[21][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_9 \y[22]  ( .clk(clk), .data_in({
        \mac_out[22][15] , \mac_out[22][14] , \mac_out[22][13] , 
        \mac_out[22][12] , \mac_out[22][11] , \mac_out[22][10] , 
        \mac_out[22][9] , \mac_out[22][8] , \mac_out[22][7] , \mac_out[22][6] , 
        \mac_out[22][5] , \mac_out[22][4] , \mac_out[22][3] , \mac_out[22][2] , 
        \mac_out[22][1] , \mac_out[22][0] }), .data_out({\mux[22][15] , 
        \mux[22][14] , \mux[22][13] , \mux[22][12] , \mux[22][11] , 
        \mux[22][10] , \mux[22][9] , \mux[22][8] , \mux[22][7] , \mux[22][6] , 
        \mux[22][5] , \mux[22][4] , \mux[22][3] , \mux[22][2] , \mux[22][1] , 
        \mux[22][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_8 \y[23]  ( .clk(clk), .data_in({
        \mac_out[23][15] , \mac_out[23][14] , \mac_out[23][13] , 
        \mac_out[23][12] , \mac_out[23][11] , \mac_out[23][10] , 
        \mac_out[23][9] , \mac_out[23][8] , \mac_out[23][7] , \mac_out[23][6] , 
        \mac_out[23][5] , \mac_out[23][4] , \mac_out[23][3] , \mac_out[23][2] , 
        \mac_out[23][1] , \mac_out[23][0] }), .data_out({\mux[23][15] , 
        \mux[23][14] , \mux[23][13] , \mux[23][12] , \mux[23][11] , 
        \mux[23][10] , \mux[23][9] , \mux[23][8] , \mux[23][7] , \mux[23][6] , 
        \mux[23][5] , \mux[23][4] , \mux[23][3] , \mux[23][2] , \mux[23][1] , 
        \mux[23][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_7 \y[24]  ( .clk(clk), .data_in({
        \mac_out[24][15] , \mac_out[24][14] , \mac_out[24][13] , 
        \mac_out[24][12] , \mac_out[24][11] , \mac_out[24][10] , 
        \mac_out[24][9] , \mac_out[24][8] , \mac_out[24][7] , \mac_out[24][6] , 
        \mac_out[24][5] , \mac_out[24][4] , \mac_out[24][3] , \mac_out[24][2] , 
        \mac_out[24][1] , \mac_out[24][0] }), .data_out({\mux[24][15] , 
        \mux[24][14] , \mux[24][13] , \mux[24][12] , \mux[24][11] , 
        \mux[24][10] , \mux[24][9] , \mux[24][8] , \mux[24][7] , \mux[24][6] , 
        \mux[24][5] , \mux[24][4] , \mux[24][3] , \mux[24][2] , \mux[24][1] , 
        \mux[24][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_6 \y[25]  ( .clk(clk), .data_in({
        \mac_out[25][15] , \mac_out[25][14] , \mac_out[25][13] , 
        \mac_out[25][12] , \mac_out[25][11] , \mac_out[25][10] , 
        \mac_out[25][9] , \mac_out[25][8] , \mac_out[25][7] , \mac_out[25][6] , 
        \mac_out[25][5] , \mac_out[25][4] , \mac_out[25][3] , \mac_out[25][2] , 
        \mac_out[25][1] , \mac_out[25][0] }), .data_out({\mux[25][15] , 
        \mux[25][14] , \mux[25][13] , \mux[25][12] , \mux[25][11] , 
        \mux[25][10] , \mux[25][9] , \mux[25][8] , \mux[25][7] , \mux[25][6] , 
        \mux[25][5] , \mux[25][4] , \mux[25][3] , \mux[25][2] , \mux[25][1] , 
        \mux[25][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        wr_en_y) );
  memory_WIDTH16_SIZE1_LOGSIZE6_5 \y[26]  ( .clk(clk), .data_in({
        \mac_out[26][15] , \mac_out[26][14] , \mac_out[26][13] , 
        \mac_out[26][12] , \mac_out[26][11] , \mac_out[26][10] , 
        \mac_out[26][9] , \mac_out[26][8] , \mac_out[26][7] , \mac_out[26][6] , 
        \mac_out[26][5] , \mac_out[26][4] , \mac_out[26][3] , \mac_out[26][2] , 
        \mac_out[26][1] , \mac_out[26][0] }), .data_out({\mux[26][15] , 
        \mux[26][14] , \mux[26][13] , \mux[26][12] , \mux[26][11] , 
        \mux[26][10] , \mux[26][9] , \mux[26][8] , \mux[26][7] , \mux[26][6] , 
        \mux[26][5] , \mux[26][4] , \mux[26][3] , \mux[26][2] , \mux[26][1] , 
        \mux[26][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        wr_en_y) );
  memory_WIDTH16_SIZE1_LOGSIZE6_4 \y[27]  ( .clk(clk), .data_in({
        \mac_out[27][15] , \mac_out[27][14] , \mac_out[27][13] , 
        \mac_out[27][12] , \mac_out[27][11] , \mac_out[27][10] , 
        \mac_out[27][9] , \mac_out[27][8] , \mac_out[27][7] , \mac_out[27][6] , 
        \mac_out[27][5] , \mac_out[27][4] , \mac_out[27][3] , \mac_out[27][2] , 
        \mac_out[27][1] , \mac_out[27][0] }), .data_out({\mux[27][15] , 
        \mux[27][14] , \mux[27][13] , \mux[27][12] , \mux[27][11] , 
        \mux[27][10] , \mux[27][9] , \mux[27][8] , \mux[27][7] , \mux[27][6] , 
        \mux[27][5] , \mux[27][4] , \mux[27][3] , \mux[27][2] , \mux[27][1] , 
        \mux[27][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_3 \y[28]  ( .clk(clk), .data_in({
        \mac_out[28][15] , \mac_out[28][14] , \mac_out[28][13] , 
        \mac_out[28][12] , \mac_out[28][11] , \mac_out[28][10] , 
        \mac_out[28][9] , \mac_out[28][8] , \mac_out[28][7] , \mac_out[28][6] , 
        \mac_out[28][5] , \mac_out[28][4] , \mac_out[28][3] , \mac_out[28][2] , 
        \mac_out[28][1] , \mac_out[28][0] }), .data_out({\mux[28][15] , 
        \mux[28][14] , \mux[28][13] , \mux[28][12] , \mux[28][11] , 
        \mux[28][10] , \mux[28][9] , \mux[28][8] , \mux[28][7] , \mux[28][6] , 
        \mux[28][5] , \mux[28][4] , \mux[28][3] , \mux[28][2] , \mux[28][1] , 
        \mux[28][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_2 \y[29]  ( .clk(clk), .data_in({
        \mac_out[29][15] , \mac_out[29][14] , \mac_out[29][13] , 
        \mac_out[29][12] , \mac_out[29][11] , \mac_out[29][10] , 
        \mac_out[29][9] , \mac_out[29][8] , \mac_out[29][7] , \mac_out[29][6] , 
        \mac_out[29][5] , \mac_out[29][4] , \mac_out[29][3] , \mac_out[29][2] , 
        \mac_out[29][1] , \mac_out[29][0] }), .data_out({\mux[29][15] , 
        \mux[29][14] , \mux[29][13] , \mux[29][12] , \mux[29][11] , 
        \mux[29][10] , \mux[29][9] , \mux[29][8] , \mux[29][7] , \mux[29][6] , 
        \mux[29][5] , \mux[29][4] , \mux[29][3] , \mux[29][2] , \mux[29][1] , 
        \mux[29][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  memory_WIDTH16_SIZE1_LOGSIZE6_1 \y[30]  ( .clk(clk), .data_in({
        \mac_out[30][15] , \mac_out[30][14] , \mac_out[30][13] , 
        \mac_out[30][12] , \mac_out[30][11] , \mac_out[30][10] , 
        \mac_out[30][9] , \mac_out[30][8] , \mac_out[30][7] , \mac_out[30][6] , 
        \mac_out[30][5] , \mac_out[30][4] , \mac_out[30][3] , \mac_out[30][2] , 
        \mac_out[30][1] , \mac_out[30][0] }), .data_out({\mux[30][15] , 
        \mux[30][14] , \mux[30][13] , \mux[30][12] , \mux[30][11] , 
        \mux[30][10] , \mux[30][9] , \mux[30][8] , \mux[30][7] , \mux[30][6] , 
        \mux[30][5] , \mux[30][4] , \mux[30][3] , \mux[30][2] , \mux[30][1] , 
        \mux[30][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n557) );
  memory_WIDTH16_SIZE1_LOGSIZE6_0 \y[31]  ( .clk(clk), .data_in({
        \mac_out[31][15] , \mac_out[31][14] , \mac_out[31][13] , 
        \mac_out[31][12] , \mac_out[31][11] , \mac_out[31][10] , 
        \mac_out[31][9] , \mac_out[31][8] , \mac_out[31][7] , \mac_out[31][6] , 
        \mac_out[31][5] , \mac_out[31][4] , \mac_out[31][3] , \mac_out[31][2] , 
        \mac_out[31][1] , \mac_out[31][0] }), .data_out({\mux[31][15] , 
        \mux[31][14] , \mux[31][13] , \mux[31][12] , \mux[31][11] , 
        \mux[31][10] , \mux[31][9] , \mux[31][8] , \mux[31][7] , \mux[31][6] , 
        \mux[31][5] , \mux[31][4] , \mux[31][3] , \mux[31][2] , \mux[31][1] , 
        \mux[31][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(
        n558) );
  BUF_X1 U2 ( .A(n537), .Z(n22) );
  CLKBUF_X3 U3 ( .A(vector_out[6]), .Z(n552) );
  CLKBUF_X3 U4 ( .A(vector_out[6]), .Z(n7) );
  CLKBUF_X3 U5 ( .A(vector_out[6]), .Z(n553) );
  BUF_X2 U6 ( .A(vector_out[2]), .Z(n18) );
  CLKBUF_X2 U7 ( .A(vector_out[2]), .Z(n14) );
  CLKBUF_X2 U8 ( .A(vector_out[2]), .Z(n540) );
  BUF_X2 U9 ( .A(vector_out[2]), .Z(n4) );
  BUF_X2 U10 ( .A(vector_out[2]), .Z(n26) );
  BUF_X2 U11 ( .A(vector_out[2]), .Z(n17) );
  BUF_X2 U12 ( .A(vector_out[2]), .Z(n541) );
  BUF_X1 U13 ( .A(n538), .Z(n21) );
  BUF_X2 U14 ( .A(n538), .Z(n27) );
  BUF_X2 U15 ( .A(n539), .Z(n23) );
  BUF_X2 U16 ( .A(vector_out[1]), .Z(n539) );
  BUF_X2 U17 ( .A(n537), .Z(n16) );
  BUF_X1 U18 ( .A(n539), .Z(n25) );
  CLKBUF_X3 U19 ( .A(n544), .Z(n12) );
  BUF_X1 U20 ( .A(vector_out[3]), .Z(n544) );
  CLKBUF_X3 U21 ( .A(n539), .Z(n533) );
  CLKBUF_X3 U22 ( .A(n538), .Z(n528) );
  BUF_X1 U23 ( .A(vector_out[1]), .Z(n537) );
  CLKBUF_X3 U24 ( .A(n538), .Z(n529) );
  BUF_X2 U25 ( .A(vector_out[1]), .Z(n538) );
  BUF_X2 U26 ( .A(vector_out[0]), .Z(n534) );
  BUF_X1 U27 ( .A(n539), .Z(n28) );
  CLKBUF_X2 U28 ( .A(vector_out[2]), .Z(n5) );
  BUF_X4 U29 ( .A(vector_out[4]), .Z(n546) );
  BUF_X4 U30 ( .A(vector_out[2]), .Z(n542) );
  BUF_X4 U31 ( .A(vector_out[5]), .Z(n1) );
  BUF_X4 U32 ( .A(vector_out[5]), .Z(n550) );
  BUF_X4 U33 ( .A(vector_out[4]), .Z(n2) );
  BUF_X4 U34 ( .A(vector_out[4]), .Z(n3) );
  CLKBUF_X3 U35 ( .A(vector_out[3]), .Z(n6) );
  BUF_X4 U36 ( .A(vector_out[6]), .Z(n8) );
  BUF_X4 U37 ( .A(vector_out[4]), .Z(n9) );
  BUF_X4 U38 ( .A(vector_out[4]), .Z(n547) );
  CLKBUF_X3 U39 ( .A(n538), .Z(n24) );
  BUF_X4 U40 ( .A(vector_out[4]), .Z(n548) );
  CLKBUF_X3 U41 ( .A(vector_out[0]), .Z(n10) );
  CLKBUF_X1 U42 ( .A(n544), .Z(n11) );
  CLKBUF_X3 U43 ( .A(n544), .Z(n13) );
  BUF_X4 U44 ( .A(vector_out[3]), .Z(n19) );
  BUF_X4 U45 ( .A(vector_out[2]), .Z(n15) );
  CLKBUF_X3 U46 ( .A(vector_out[3]), .Z(n545) );
  CLKBUF_X3 U47 ( .A(vector_out[3]), .Z(n20) );
  CLKBUF_X3 U48 ( .A(n538), .Z(n532) );
  CLKBUF_X3 U49 ( .A(n539), .Z(n531) );
  BUF_X4 U50 ( .A(vector_out[3]), .Z(n543) );
  CLKBUF_X3 U51 ( .A(vector_out[0]), .Z(n535) );
  CLKBUF_X3 U52 ( .A(n539), .Z(n530) );
  BUF_X1 U53 ( .A(n527), .Z(n522) );
  BUF_X1 U54 ( .A(n527), .Z(n524) );
  BUF_X1 U55 ( .A(n527), .Z(n523) );
  BUF_X1 U56 ( .A(n526), .Z(n518) );
  BUF_X1 U57 ( .A(n527), .Z(n520) );
  BUF_X1 U58 ( .A(n527), .Z(n519) );
  BUF_X1 U59 ( .A(n527), .Z(n521) );
  BUF_X1 U60 ( .A(n518), .Z(n517) );
  BUF_X1 U61 ( .A(n525), .Z(n526) );
  BUF_X1 U62 ( .A(n525), .Z(n527) );
  BUF_X1 U63 ( .A(addr_y[1]), .Z(n515) );
  BUF_X1 U64 ( .A(n512), .Z(n514) );
  BUF_X1 U65 ( .A(n516), .Z(n512) );
  BUF_X1 U66 ( .A(n516), .Z(n513) );
  BUF_X1 U67 ( .A(addr_y[0]), .Z(n525) );
  BUF_X1 U68 ( .A(clear_acc), .Z(n559) );
  BUF_X1 U69 ( .A(wr_en_y), .Z(n557) );
  BUF_X1 U70 ( .A(wr_en_y), .Z(n558) );
  BUF_X1 U71 ( .A(clear_acc), .Z(n560) );
  BUF_X1 U72 ( .A(addr_y[2]), .Z(n510) );
  BUF_X1 U73 ( .A(addr_y[2]), .Z(n511) );
  BUF_X1 U74 ( .A(addr_y[3]), .Z(n509) );
  BUF_X1 U75 ( .A(addr_y[1]), .Z(n516) );
  BUF_X4 U76 ( .A(vector_out[5]), .Z(n549) );
  BUF_X4 U77 ( .A(vector_out[7]), .Z(n555) );
  BUF_X4 U78 ( .A(vector_out[7]), .Z(n554) );
  MUX2_X1 U79 ( .A(\mux[30][0] ), .B(\mux[31][0] ), .S(n520), .Z(n29) );
  MUX2_X1 U80 ( .A(\mux[28][0] ), .B(\mux[29][0] ), .S(n519), .Z(n30) );
  MUX2_X1 U81 ( .A(n30), .B(n29), .S(n515), .Z(n31) );
  MUX2_X1 U82 ( .A(\mux[26][0] ), .B(\mux[27][0] ), .S(n521), .Z(n32) );
  MUX2_X1 U83 ( .A(\mux[24][0] ), .B(\mux[25][0] ), .S(n525), .Z(n33) );
  MUX2_X1 U84 ( .A(n33), .B(n32), .S(n514), .Z(n34) );
  MUX2_X1 U85 ( .A(n34), .B(n31), .S(n511), .Z(n35) );
  MUX2_X1 U86 ( .A(\mux[22][0] ), .B(\mux[23][0] ), .S(addr_y[0]), .Z(n36) );
  MUX2_X1 U87 ( .A(\mux[20][0] ), .B(\mux[21][0] ), .S(n525), .Z(n37) );
  MUX2_X1 U88 ( .A(n37), .B(n36), .S(addr_y[1]), .Z(n38) );
  MUX2_X1 U89 ( .A(\mux[18][0] ), .B(\mux[19][0] ), .S(addr_y[0]), .Z(n39) );
  MUX2_X1 U90 ( .A(\mux[16][0] ), .B(\mux[17][0] ), .S(n519), .Z(n40) );
  MUX2_X1 U91 ( .A(n40), .B(n39), .S(n516), .Z(n41) );
  MUX2_X1 U92 ( .A(n41), .B(n38), .S(n511), .Z(n42) );
  MUX2_X1 U93 ( .A(n42), .B(n35), .S(addr_y[3]), .Z(n43) );
  MUX2_X1 U94 ( .A(\mux[14][0] ), .B(\mux[15][0] ), .S(n518), .Z(n44) );
  MUX2_X1 U95 ( .A(\mux[12][0] ), .B(\mux[13][0] ), .S(n525), .Z(n45) );
  MUX2_X1 U96 ( .A(n45), .B(n44), .S(n512), .Z(n46) );
  MUX2_X1 U97 ( .A(\mux[10][0] ), .B(\mux[11][0] ), .S(addr_y[0]), .Z(n47) );
  MUX2_X1 U98 ( .A(\mux[8][0] ), .B(\mux[9][0] ), .S(n521), .Z(n48) );
  MUX2_X1 U99 ( .A(n48), .B(n47), .S(n513), .Z(n49) );
  MUX2_X1 U100 ( .A(n49), .B(n46), .S(addr_y[2]), .Z(n50) );
  MUX2_X1 U101 ( .A(\mux[6][0] ), .B(\mux[7][0] ), .S(n525), .Z(n51) );
  MUX2_X1 U102 ( .A(\mux[4][0] ), .B(\mux[5][0] ), .S(n525), .Z(n52) );
  MUX2_X1 U103 ( .A(n52), .B(n51), .S(addr_y[1]), .Z(n53) );
  MUX2_X1 U104 ( .A(\mux[2][0] ), .B(\mux[3][0] ), .S(addr_y[0]), .Z(n54) );
  MUX2_X1 U105 ( .A(\mux[0][0] ), .B(\mux[1][0] ), .S(n527), .Z(n55) );
  MUX2_X1 U106 ( .A(n55), .B(n54), .S(n515), .Z(n56) );
  MUX2_X1 U107 ( .A(n56), .B(n53), .S(n510), .Z(n57) );
  MUX2_X1 U108 ( .A(n57), .B(n50), .S(addr_y[3]), .Z(n58) );
  MUX2_X1 U109 ( .A(n58), .B(n43), .S(addr_y[4]), .Z(data_out[0]) );
  MUX2_X1 U110 ( .A(\mux[30][1] ), .B(\mux[31][1] ), .S(n517), .Z(n59) );
  MUX2_X1 U111 ( .A(\mux[28][1] ), .B(\mux[29][1] ), .S(n517), .Z(n60) );
  MUX2_X1 U112 ( .A(n60), .B(n59), .S(n512), .Z(n61) );
  MUX2_X1 U113 ( .A(\mux[26][1] ), .B(\mux[27][1] ), .S(n517), .Z(n62) );
  MUX2_X1 U114 ( .A(\mux[24][1] ), .B(\mux[25][1] ), .S(n517), .Z(n63) );
  MUX2_X1 U115 ( .A(n63), .B(n62), .S(n512), .Z(n64) );
  MUX2_X1 U116 ( .A(n64), .B(n61), .S(addr_y[2]), .Z(n65) );
  MUX2_X1 U117 ( .A(\mux[22][1] ), .B(\mux[23][1] ), .S(n517), .Z(n66) );
  MUX2_X1 U118 ( .A(\mux[20][1] ), .B(\mux[21][1] ), .S(n517), .Z(n67) );
  MUX2_X1 U119 ( .A(n67), .B(n66), .S(n512), .Z(n68) );
  MUX2_X1 U120 ( .A(\mux[18][1] ), .B(\mux[19][1] ), .S(n517), .Z(n69) );
  MUX2_X1 U121 ( .A(\mux[16][1] ), .B(\mux[17][1] ), .S(n517), .Z(n70) );
  MUX2_X1 U122 ( .A(n70), .B(n69), .S(n512), .Z(n71) );
  MUX2_X1 U123 ( .A(n71), .B(n68), .S(addr_y[2]), .Z(n72) );
  MUX2_X1 U124 ( .A(n72), .B(n65), .S(addr_y[3]), .Z(n73) );
  MUX2_X1 U125 ( .A(\mux[14][1] ), .B(\mux[15][1] ), .S(n517), .Z(n74) );
  MUX2_X1 U126 ( .A(\mux[12][1] ), .B(\mux[13][1] ), .S(n517), .Z(n75) );
  MUX2_X1 U127 ( .A(n75), .B(n74), .S(n512), .Z(n76) );
  MUX2_X1 U128 ( .A(\mux[10][1] ), .B(\mux[11][1] ), .S(n517), .Z(n77) );
  MUX2_X1 U129 ( .A(\mux[8][1] ), .B(\mux[9][1] ), .S(n517), .Z(n78) );
  MUX2_X1 U130 ( .A(n78), .B(n77), .S(n512), .Z(n79) );
  MUX2_X1 U131 ( .A(n79), .B(n76), .S(n511), .Z(n80) );
  MUX2_X1 U132 ( .A(\mux[6][1] ), .B(\mux[7][1] ), .S(n524), .Z(n81) );
  MUX2_X1 U133 ( .A(\mux[4][1] ), .B(\mux[5][1] ), .S(n523), .Z(n82) );
  MUX2_X1 U134 ( .A(n82), .B(n81), .S(n512), .Z(n83) );
  MUX2_X1 U135 ( .A(\mux[2][1] ), .B(\mux[3][1] ), .S(n520), .Z(n84) );
  MUX2_X1 U136 ( .A(\mux[0][1] ), .B(\mux[1][1] ), .S(n519), .Z(n85) );
  MUX2_X1 U137 ( .A(n85), .B(n84), .S(n512), .Z(n86) );
  MUX2_X1 U138 ( .A(n86), .B(n83), .S(addr_y[2]), .Z(n87) );
  MUX2_X1 U139 ( .A(n87), .B(n80), .S(addr_y[3]), .Z(n88) );
  MUX2_X1 U140 ( .A(n88), .B(n73), .S(addr_y[4]), .Z(data_out[1]) );
  MUX2_X1 U141 ( .A(\mux[30][2] ), .B(\mux[31][2] ), .S(n521), .Z(n89) );
  MUX2_X1 U142 ( .A(\mux[28][2] ), .B(\mux[29][2] ), .S(n525), .Z(n90) );
  MUX2_X1 U143 ( .A(n90), .B(n89), .S(n512), .Z(n91) );
  MUX2_X1 U144 ( .A(\mux[26][2] ), .B(\mux[27][2] ), .S(n518), .Z(n92) );
  MUX2_X1 U145 ( .A(\mux[24][2] ), .B(\mux[25][2] ), .S(n526), .Z(n93) );
  MUX2_X1 U146 ( .A(n93), .B(n92), .S(n512), .Z(n94) );
  MUX2_X1 U147 ( .A(n94), .B(n91), .S(addr_y[2]), .Z(n95) );
  MUX2_X1 U148 ( .A(\mux[22][2] ), .B(\mux[23][2] ), .S(addr_y[0]), .Z(n96) );
  MUX2_X1 U149 ( .A(\mux[20][2] ), .B(\mux[21][2] ), .S(n527), .Z(n97) );
  MUX2_X1 U150 ( .A(n97), .B(n96), .S(n512), .Z(n98) );
  MUX2_X1 U151 ( .A(\mux[18][2] ), .B(\mux[19][2] ), .S(n517), .Z(n99) );
  MUX2_X1 U152 ( .A(\mux[16][2] ), .B(\mux[17][2] ), .S(n522), .Z(n100) );
  MUX2_X1 U153 ( .A(n100), .B(n99), .S(n512), .Z(n101) );
  MUX2_X1 U154 ( .A(n101), .B(n98), .S(addr_y[2]), .Z(n102) );
  MUX2_X1 U155 ( .A(n102), .B(n95), .S(addr_y[3]), .Z(n103) );
  MUX2_X1 U156 ( .A(\mux[14][2] ), .B(\mux[15][2] ), .S(n519), .Z(n104) );
  MUX2_X1 U157 ( .A(\mux[12][2] ), .B(\mux[13][2] ), .S(n517), .Z(n105) );
  MUX2_X1 U158 ( .A(n105), .B(n104), .S(n513), .Z(n106) );
  MUX2_X1 U159 ( .A(\mux[10][2] ), .B(\mux[11][2] ), .S(addr_y[0]), .Z(n107)
         );
  MUX2_X1 U160 ( .A(\mux[8][2] ), .B(\mux[9][2] ), .S(n525), .Z(n108) );
  MUX2_X1 U161 ( .A(n108), .B(n107), .S(n513), .Z(n109) );
  MUX2_X1 U162 ( .A(n109), .B(n106), .S(n510), .Z(n110) );
  MUX2_X1 U163 ( .A(\mux[6][2] ), .B(\mux[7][2] ), .S(n521), .Z(n111) );
  MUX2_X1 U164 ( .A(\mux[4][2] ), .B(\mux[5][2] ), .S(n526), .Z(n112) );
  MUX2_X1 U165 ( .A(n112), .B(n111), .S(n513), .Z(n113) );
  MUX2_X1 U166 ( .A(\mux[2][2] ), .B(\mux[3][2] ), .S(n527), .Z(n114) );
  MUX2_X1 U167 ( .A(\mux[0][2] ), .B(\mux[1][2] ), .S(n524), .Z(n115) );
  MUX2_X1 U168 ( .A(n115), .B(n114), .S(n513), .Z(n116) );
  MUX2_X1 U169 ( .A(n116), .B(n113), .S(n511), .Z(n117) );
  MUX2_X1 U170 ( .A(n117), .B(n110), .S(addr_y[3]), .Z(n118) );
  MUX2_X1 U171 ( .A(n118), .B(n103), .S(addr_y[4]), .Z(data_out[2]) );
  MUX2_X1 U172 ( .A(\mux[30][3] ), .B(\mux[31][3] ), .S(n524), .Z(n119) );
  MUX2_X1 U173 ( .A(\mux[28][3] ), .B(\mux[29][3] ), .S(n522), .Z(n120) );
  MUX2_X1 U174 ( .A(n120), .B(n119), .S(n513), .Z(n121) );
  MUX2_X1 U175 ( .A(\mux[26][3] ), .B(\mux[27][3] ), .S(addr_y[0]), .Z(n122)
         );
  MUX2_X1 U176 ( .A(\mux[24][3] ), .B(\mux[25][3] ), .S(n525), .Z(n123) );
  MUX2_X1 U177 ( .A(n123), .B(n122), .S(n513), .Z(n124) );
  MUX2_X1 U178 ( .A(n124), .B(n121), .S(n511), .Z(n125) );
  MUX2_X1 U179 ( .A(\mux[22][3] ), .B(\mux[23][3] ), .S(addr_y[0]), .Z(n126)
         );
  MUX2_X1 U180 ( .A(\mux[20][3] ), .B(\mux[21][3] ), .S(n526), .Z(n127) );
  MUX2_X1 U181 ( .A(n127), .B(n126), .S(n513), .Z(n128) );
  MUX2_X1 U182 ( .A(\mux[18][3] ), .B(\mux[19][3] ), .S(n527), .Z(n129) );
  MUX2_X1 U183 ( .A(\mux[16][3] ), .B(\mux[17][3] ), .S(n518), .Z(n130) );
  MUX2_X1 U184 ( .A(n130), .B(n129), .S(n513), .Z(n131) );
  MUX2_X1 U185 ( .A(n131), .B(n128), .S(addr_y[2]), .Z(n132) );
  MUX2_X1 U186 ( .A(n132), .B(n125), .S(addr_y[3]), .Z(n133) );
  MUX2_X1 U187 ( .A(\mux[14][3] ), .B(\mux[15][3] ), .S(n519), .Z(n134) );
  MUX2_X1 U188 ( .A(\mux[12][3] ), .B(\mux[13][3] ), .S(n517), .Z(n135) );
  MUX2_X1 U189 ( .A(n135), .B(n134), .S(n513), .Z(n136) );
  MUX2_X1 U190 ( .A(\mux[10][3] ), .B(\mux[11][3] ), .S(n521), .Z(n137) );
  MUX2_X1 U191 ( .A(\mux[8][3] ), .B(\mux[9][3] ), .S(addr_y[0]), .Z(n138) );
  MUX2_X1 U192 ( .A(n138), .B(n137), .S(n513), .Z(n139) );
  MUX2_X1 U193 ( .A(n139), .B(n136), .S(addr_y[2]), .Z(n140) );
  MUX2_X1 U194 ( .A(\mux[6][3] ), .B(\mux[7][3] ), .S(n525), .Z(n141) );
  MUX2_X1 U195 ( .A(\mux[4][3] ), .B(\mux[5][3] ), .S(n526), .Z(n142) );
  MUX2_X1 U196 ( .A(n142), .B(n141), .S(n513), .Z(n143) );
  MUX2_X1 U197 ( .A(\mux[2][3] ), .B(\mux[3][3] ), .S(n527), .Z(n144) );
  MUX2_X1 U198 ( .A(\mux[0][3] ), .B(\mux[1][3] ), .S(n522), .Z(n145) );
  MUX2_X1 U199 ( .A(n145), .B(n144), .S(n513), .Z(n146) );
  MUX2_X1 U200 ( .A(n146), .B(n143), .S(n510), .Z(n147) );
  MUX2_X1 U201 ( .A(n147), .B(n140), .S(addr_y[3]), .Z(n148) );
  MUX2_X1 U202 ( .A(n148), .B(n133), .S(addr_y[4]), .Z(data_out[3]) );
  MUX2_X1 U203 ( .A(\mux[30][4] ), .B(\mux[31][4] ), .S(n526), .Z(n149) );
  MUX2_X1 U204 ( .A(\mux[28][4] ), .B(\mux[29][4] ), .S(n527), .Z(n150) );
  MUX2_X1 U205 ( .A(n150), .B(n149), .S(n516), .Z(n151) );
  MUX2_X1 U206 ( .A(\mux[26][4] ), .B(\mux[27][4] ), .S(n523), .Z(n152) );
  MUX2_X1 U207 ( .A(\mux[24][4] ), .B(\mux[25][4] ), .S(n522), .Z(n153) );
  MUX2_X1 U208 ( .A(n153), .B(n152), .S(n512), .Z(n154) );
  MUX2_X1 U209 ( .A(n154), .B(n151), .S(addr_y[2]), .Z(n155) );
  MUX2_X1 U210 ( .A(\mux[22][4] ), .B(\mux[23][4] ), .S(addr_y[0]), .Z(n156)
         );
  MUX2_X1 U211 ( .A(\mux[20][4] ), .B(\mux[21][4] ), .S(n524), .Z(n157) );
  MUX2_X1 U212 ( .A(n157), .B(n156), .S(n513), .Z(n158) );
  MUX2_X1 U213 ( .A(\mux[18][4] ), .B(\mux[19][4] ), .S(n525), .Z(n159) );
  MUX2_X1 U214 ( .A(\mux[16][4] ), .B(\mux[17][4] ), .S(addr_y[0]), .Z(n160)
         );
  MUX2_X1 U215 ( .A(n160), .B(n159), .S(n515), .Z(n161) );
  MUX2_X1 U216 ( .A(n161), .B(n158), .S(n510), .Z(n162) );
  MUX2_X1 U217 ( .A(n162), .B(n155), .S(n509), .Z(n163) );
  MUX2_X1 U218 ( .A(\mux[14][4] ), .B(\mux[15][4] ), .S(n526), .Z(n164) );
  MUX2_X1 U219 ( .A(\mux[12][4] ), .B(\mux[13][4] ), .S(n527), .Z(n165) );
  MUX2_X1 U220 ( .A(n165), .B(n164), .S(n514), .Z(n166) );
  MUX2_X1 U221 ( .A(\mux[10][4] ), .B(\mux[11][4] ), .S(n520), .Z(n167) );
  MUX2_X1 U222 ( .A(\mux[8][4] ), .B(\mux[9][4] ), .S(n523), .Z(n168) );
  MUX2_X1 U223 ( .A(n168), .B(n167), .S(n512), .Z(n169) );
  MUX2_X1 U224 ( .A(n169), .B(n166), .S(addr_y[2]), .Z(n170) );
  MUX2_X1 U225 ( .A(\mux[6][4] ), .B(\mux[7][4] ), .S(n526), .Z(n171) );
  MUX2_X1 U226 ( .A(\mux[4][4] ), .B(\mux[5][4] ), .S(n527), .Z(n172) );
  MUX2_X1 U227 ( .A(n172), .B(n171), .S(addr_y[1]), .Z(n173) );
  MUX2_X1 U228 ( .A(\mux[2][4] ), .B(\mux[3][4] ), .S(n525), .Z(n174) );
  MUX2_X1 U229 ( .A(\mux[0][4] ), .B(\mux[1][4] ), .S(addr_y[0]), .Z(n175) );
  MUX2_X1 U230 ( .A(n175), .B(n174), .S(n516), .Z(n176) );
  MUX2_X1 U231 ( .A(n176), .B(n173), .S(n511), .Z(n177) );
  MUX2_X1 U232 ( .A(n177), .B(n170), .S(n509), .Z(n178) );
  MUX2_X1 U233 ( .A(n178), .B(n163), .S(addr_y[4]), .Z(data_out[4]) );
  MUX2_X1 U234 ( .A(\mux[30][5] ), .B(\mux[31][5] ), .S(n517), .Z(n179) );
  MUX2_X1 U235 ( .A(\mux[28][5] ), .B(\mux[29][5] ), .S(addr_y[0]), .Z(n180)
         );
  MUX2_X1 U236 ( .A(n180), .B(n179), .S(n512), .Z(n181) );
  MUX2_X1 U237 ( .A(\mux[26][5] ), .B(\mux[27][5] ), .S(n525), .Z(n182) );
  MUX2_X1 U238 ( .A(\mux[24][5] ), .B(\mux[25][5] ), .S(n522), .Z(n183) );
  MUX2_X1 U239 ( .A(n183), .B(n182), .S(n513), .Z(n184) );
  MUX2_X1 U240 ( .A(n184), .B(n181), .S(addr_y[2]), .Z(n185) );
  MUX2_X1 U241 ( .A(\mux[22][5] ), .B(\mux[23][5] ), .S(n526), .Z(n186) );
  MUX2_X1 U242 ( .A(\mux[20][5] ), .B(\mux[21][5] ), .S(n527), .Z(n187) );
  MUX2_X1 U243 ( .A(n187), .B(n186), .S(n515), .Z(n188) );
  MUX2_X1 U244 ( .A(\mux[18][5] ), .B(\mux[19][5] ), .S(n526), .Z(n189) );
  MUX2_X1 U245 ( .A(\mux[16][5] ), .B(\mux[17][5] ), .S(n520), .Z(n190) );
  MUX2_X1 U246 ( .A(n190), .B(n189), .S(n514), .Z(n191) );
  MUX2_X1 U247 ( .A(n191), .B(n188), .S(n510), .Z(n192) );
  MUX2_X1 U248 ( .A(n192), .B(n185), .S(n509), .Z(n193) );
  MUX2_X1 U249 ( .A(\mux[14][5] ), .B(\mux[15][5] ), .S(n526), .Z(n194) );
  MUX2_X1 U250 ( .A(\mux[12][5] ), .B(\mux[13][5] ), .S(n526), .Z(n195) );
  MUX2_X1 U251 ( .A(n195), .B(n194), .S(n516), .Z(n196) );
  MUX2_X1 U252 ( .A(\mux[10][5] ), .B(\mux[11][5] ), .S(n520), .Z(n197) );
  MUX2_X1 U253 ( .A(\mux[8][5] ), .B(\mux[9][5] ), .S(n525), .Z(n198) );
  MUX2_X1 U254 ( .A(n198), .B(n197), .S(n514), .Z(n199) );
  MUX2_X1 U255 ( .A(n199), .B(n196), .S(addr_y[2]), .Z(n200) );
  MUX2_X1 U256 ( .A(\mux[6][5] ), .B(\mux[7][5] ), .S(addr_y[0]), .Z(n201) );
  MUX2_X1 U257 ( .A(\mux[4][5] ), .B(\mux[5][5] ), .S(n527), .Z(n202) );
  MUX2_X1 U258 ( .A(n202), .B(n201), .S(n515), .Z(n203) );
  MUX2_X1 U259 ( .A(\mux[2][5] ), .B(\mux[3][5] ), .S(n526), .Z(n204) );
  MUX2_X1 U260 ( .A(\mux[0][5] ), .B(\mux[1][5] ), .S(n526), .Z(n205) );
  MUX2_X1 U261 ( .A(n205), .B(n204), .S(n516), .Z(n206) );
  MUX2_X1 U262 ( .A(n206), .B(n203), .S(addr_y[2]), .Z(n207) );
  MUX2_X1 U263 ( .A(n207), .B(n200), .S(n509), .Z(n208) );
  MUX2_X1 U264 ( .A(n208), .B(n193), .S(addr_y[4]), .Z(data_out[5]) );
  MUX2_X1 U265 ( .A(\mux[30][6] ), .B(\mux[31][6] ), .S(n527), .Z(n209) );
  MUX2_X1 U266 ( .A(\mux[28][6] ), .B(\mux[29][6] ), .S(n527), .Z(n210) );
  MUX2_X1 U267 ( .A(n210), .B(n209), .S(addr_y[1]), .Z(n211) );
  MUX2_X1 U268 ( .A(\mux[26][6] ), .B(\mux[27][6] ), .S(n519), .Z(n212) );
  MUX2_X1 U269 ( .A(\mux[24][6] ), .B(\mux[25][6] ), .S(addr_y[0]), .Z(n213)
         );
  MUX2_X1 U270 ( .A(n213), .B(n212), .S(n512), .Z(n214) );
  MUX2_X1 U271 ( .A(n214), .B(n211), .S(addr_y[2]), .Z(n215) );
  MUX2_X1 U272 ( .A(\mux[22][6] ), .B(\mux[23][6] ), .S(addr_y[0]), .Z(n216)
         );
  MUX2_X1 U273 ( .A(\mux[20][6] ), .B(\mux[21][6] ), .S(n525), .Z(n217) );
  MUX2_X1 U274 ( .A(n217), .B(n216), .S(n513), .Z(n218) );
  MUX2_X1 U275 ( .A(\mux[18][6] ), .B(\mux[19][6] ), .S(n524), .Z(n219) );
  MUX2_X1 U276 ( .A(\mux[16][6] ), .B(\mux[17][6] ), .S(n526), .Z(n220) );
  MUX2_X1 U277 ( .A(n220), .B(n219), .S(n514), .Z(n221) );
  MUX2_X1 U278 ( .A(n221), .B(n218), .S(addr_y[2]), .Z(n222) );
  MUX2_X1 U279 ( .A(n222), .B(n215), .S(n509), .Z(n223) );
  MUX2_X1 U280 ( .A(\mux[14][6] ), .B(\mux[15][6] ), .S(n526), .Z(n224) );
  MUX2_X1 U281 ( .A(\mux[12][6] ), .B(\mux[13][6] ), .S(n527), .Z(n225) );
  MUX2_X1 U282 ( .A(n225), .B(n224), .S(n516), .Z(n226) );
  MUX2_X1 U283 ( .A(\mux[10][6] ), .B(\mux[11][6] ), .S(n518), .Z(n227) );
  MUX2_X1 U284 ( .A(\mux[8][6] ), .B(\mux[9][6] ), .S(n523), .Z(n228) );
  MUX2_X1 U285 ( .A(n228), .B(n227), .S(n515), .Z(n229) );
  MUX2_X1 U286 ( .A(n229), .B(n226), .S(n510), .Z(n230) );
  MUX2_X1 U287 ( .A(\mux[6][6] ), .B(\mux[7][6] ), .S(addr_y[0]), .Z(n231) );
  MUX2_X1 U288 ( .A(\mux[4][6] ), .B(\mux[5][6] ), .S(n525), .Z(n232) );
  MUX2_X1 U289 ( .A(n232), .B(n231), .S(n514), .Z(n233) );
  MUX2_X1 U290 ( .A(\mux[2][6] ), .B(\mux[3][6] ), .S(n525), .Z(n234) );
  MUX2_X1 U291 ( .A(\mux[0][6] ), .B(\mux[1][6] ), .S(n526), .Z(n235) );
  MUX2_X1 U292 ( .A(n235), .B(n234), .S(n513), .Z(n236) );
  MUX2_X1 U293 ( .A(n236), .B(n233), .S(addr_y[2]), .Z(n237) );
  MUX2_X1 U294 ( .A(n237), .B(n230), .S(n509), .Z(n238) );
  MUX2_X1 U295 ( .A(n238), .B(n223), .S(addr_y[4]), .Z(data_out[6]) );
  MUX2_X1 U296 ( .A(\mux[30][7] ), .B(\mux[31][7] ), .S(n526), .Z(n239) );
  MUX2_X1 U297 ( .A(\mux[28][7] ), .B(\mux[29][7] ), .S(n518), .Z(n240) );
  MUX2_X1 U298 ( .A(n240), .B(n239), .S(n514), .Z(n241) );
  MUX2_X1 U299 ( .A(\mux[26][7] ), .B(\mux[27][7] ), .S(n525), .Z(n242) );
  MUX2_X1 U300 ( .A(\mux[24][7] ), .B(\mux[25][7] ), .S(n527), .Z(n243) );
  MUX2_X1 U301 ( .A(n243), .B(n242), .S(n514), .Z(n244) );
  MUX2_X1 U302 ( .A(n244), .B(n241), .S(n510), .Z(n245) );
  MUX2_X1 U303 ( .A(\mux[22][7] ), .B(\mux[23][7] ), .S(n517), .Z(n246) );
  MUX2_X1 U304 ( .A(\mux[20][7] ), .B(\mux[21][7] ), .S(n521), .Z(n247) );
  MUX2_X1 U305 ( .A(n247), .B(n246), .S(n514), .Z(n248) );
  MUX2_X1 U306 ( .A(\mux[18][7] ), .B(\mux[19][7] ), .S(n527), .Z(n249) );
  MUX2_X1 U307 ( .A(\mux[16][7] ), .B(\mux[17][7] ), .S(n522), .Z(n250) );
  MUX2_X1 U308 ( .A(n250), .B(n249), .S(n514), .Z(n251) );
  MUX2_X1 U309 ( .A(n251), .B(n248), .S(n510), .Z(n252) );
  MUX2_X1 U310 ( .A(n252), .B(n245), .S(n509), .Z(n253) );
  MUX2_X1 U311 ( .A(\mux[14][7] ), .B(\mux[15][7] ), .S(n524), .Z(n254) );
  MUX2_X1 U312 ( .A(\mux[12][7] ), .B(\mux[13][7] ), .S(n523), .Z(n255) );
  MUX2_X1 U313 ( .A(n255), .B(n254), .S(n514), .Z(n256) );
  MUX2_X1 U314 ( .A(\mux[10][7] ), .B(\mux[11][7] ), .S(n520), .Z(n257) );
  MUX2_X1 U315 ( .A(\mux[8][7] ), .B(\mux[9][7] ), .S(n519), .Z(n258) );
  MUX2_X1 U316 ( .A(n258), .B(n257), .S(n514), .Z(n259) );
  MUX2_X1 U317 ( .A(n259), .B(n256), .S(n510), .Z(n260) );
  MUX2_X1 U318 ( .A(\mux[6][7] ), .B(\mux[7][7] ), .S(n517), .Z(n261) );
  MUX2_X1 U319 ( .A(\mux[4][7] ), .B(\mux[5][7] ), .S(n525), .Z(n262) );
  MUX2_X1 U320 ( .A(n262), .B(n261), .S(n514), .Z(n263) );
  MUX2_X1 U321 ( .A(\mux[2][7] ), .B(\mux[3][7] ), .S(n517), .Z(n264) );
  MUX2_X1 U322 ( .A(\mux[0][7] ), .B(\mux[1][7] ), .S(n522), .Z(n265) );
  MUX2_X1 U323 ( .A(n265), .B(n264), .S(n514), .Z(n266) );
  MUX2_X1 U324 ( .A(n266), .B(n263), .S(n510), .Z(n267) );
  MUX2_X1 U325 ( .A(n267), .B(n260), .S(n509), .Z(n268) );
  MUX2_X1 U326 ( .A(n268), .B(n253), .S(addr_y[4]), .Z(data_out[7]) );
  MUX2_X1 U327 ( .A(\mux[30][8] ), .B(\mux[31][8] ), .S(n524), .Z(n269) );
  MUX2_X1 U328 ( .A(\mux[28][8] ), .B(\mux[29][8] ), .S(n523), .Z(n270) );
  MUX2_X1 U329 ( .A(n270), .B(n269), .S(n514), .Z(n271) );
  MUX2_X1 U330 ( .A(\mux[26][8] ), .B(\mux[27][8] ), .S(n520), .Z(n272) );
  MUX2_X1 U331 ( .A(\mux[24][8] ), .B(\mux[25][8] ), .S(n519), .Z(n273) );
  MUX2_X1 U332 ( .A(n273), .B(n272), .S(n514), .Z(n274) );
  MUX2_X1 U333 ( .A(n274), .B(n271), .S(n510), .Z(n275) );
  MUX2_X1 U334 ( .A(\mux[22][8] ), .B(\mux[23][8] ), .S(n521), .Z(n276) );
  MUX2_X1 U335 ( .A(\mux[20][8] ), .B(\mux[21][8] ), .S(n521), .Z(n277) );
  MUX2_X1 U336 ( .A(n277), .B(n276), .S(n514), .Z(n278) );
  MUX2_X1 U337 ( .A(\mux[18][8] ), .B(\mux[19][8] ), .S(n520), .Z(n279) );
  MUX2_X1 U338 ( .A(\mux[16][8] ), .B(\mux[17][8] ), .S(n523), .Z(n280) );
  MUX2_X1 U339 ( .A(n280), .B(n279), .S(n514), .Z(n281) );
  MUX2_X1 U340 ( .A(n281), .B(n278), .S(n510), .Z(n282) );
  MUX2_X1 U341 ( .A(n282), .B(n275), .S(n509), .Z(n283) );
  MUX2_X1 U342 ( .A(\mux[14][8] ), .B(\mux[15][8] ), .S(n518), .Z(n284) );
  MUX2_X1 U343 ( .A(\mux[12][8] ), .B(\mux[13][8] ), .S(n518), .Z(n285) );
  MUX2_X1 U344 ( .A(n285), .B(n284), .S(n513), .Z(n286) );
  MUX2_X1 U345 ( .A(\mux[10][8] ), .B(\mux[11][8] ), .S(n518), .Z(n287) );
  MUX2_X1 U346 ( .A(\mux[8][8] ), .B(\mux[9][8] ), .S(n518), .Z(n288) );
  MUX2_X1 U347 ( .A(n288), .B(n287), .S(n516), .Z(n289) );
  MUX2_X1 U348 ( .A(n289), .B(n286), .S(n510), .Z(n290) );
  MUX2_X1 U349 ( .A(\mux[6][8] ), .B(\mux[7][8] ), .S(n518), .Z(n291) );
  MUX2_X1 U350 ( .A(\mux[4][8] ), .B(\mux[5][8] ), .S(n518), .Z(n292) );
  MUX2_X1 U351 ( .A(n292), .B(n291), .S(n512), .Z(n293) );
  MUX2_X1 U352 ( .A(\mux[2][8] ), .B(\mux[3][8] ), .S(n518), .Z(n294) );
  MUX2_X1 U353 ( .A(\mux[0][8] ), .B(\mux[1][8] ), .S(n518), .Z(n295) );
  MUX2_X1 U354 ( .A(n295), .B(n294), .S(n515), .Z(n296) );
  MUX2_X1 U355 ( .A(n296), .B(n293), .S(n510), .Z(n297) );
  MUX2_X1 U356 ( .A(n297), .B(n290), .S(n509), .Z(n298) );
  MUX2_X1 U357 ( .A(n298), .B(n283), .S(addr_y[4]), .Z(data_out[8]) );
  MUX2_X1 U358 ( .A(\mux[30][9] ), .B(\mux[31][9] ), .S(n518), .Z(n299) );
  MUX2_X1 U359 ( .A(\mux[28][9] ), .B(\mux[29][9] ), .S(n518), .Z(n300) );
  MUX2_X1 U360 ( .A(n300), .B(n299), .S(n514), .Z(n301) );
  MUX2_X1 U361 ( .A(\mux[26][9] ), .B(\mux[27][9] ), .S(n518), .Z(n302) );
  MUX2_X1 U362 ( .A(\mux[24][9] ), .B(\mux[25][9] ), .S(n518), .Z(n303) );
  MUX2_X1 U363 ( .A(n303), .B(n302), .S(n513), .Z(n304) );
  MUX2_X1 U364 ( .A(n304), .B(n301), .S(n510), .Z(n305) );
  MUX2_X1 U365 ( .A(\mux[22][9] ), .B(\mux[23][9] ), .S(n521), .Z(n306) );
  MUX2_X1 U366 ( .A(\mux[20][9] ), .B(\mux[21][9] ), .S(addr_y[0]), .Z(n307)
         );
  MUX2_X1 U367 ( .A(n307), .B(n306), .S(addr_y[1]), .Z(n308) );
  MUX2_X1 U368 ( .A(\mux[18][9] ), .B(\mux[19][9] ), .S(n518), .Z(n309) );
  MUX2_X1 U369 ( .A(\mux[16][9] ), .B(\mux[17][9] ), .S(n526), .Z(n310) );
  MUX2_X1 U370 ( .A(n310), .B(n309), .S(n516), .Z(n311) );
  MUX2_X1 U371 ( .A(n311), .B(n308), .S(n510), .Z(n312) );
  MUX2_X1 U372 ( .A(n312), .B(n305), .S(n509), .Z(n313) );
  MUX2_X1 U373 ( .A(\mux[14][9] ), .B(\mux[15][9] ), .S(n525), .Z(n314) );
  MUX2_X1 U374 ( .A(\mux[12][9] ), .B(\mux[13][9] ), .S(n527), .Z(n315) );
  MUX2_X1 U375 ( .A(n315), .B(n314), .S(n512), .Z(n316) );
  MUX2_X1 U376 ( .A(\mux[10][9] ), .B(\mux[11][9] ), .S(n517), .Z(n317) );
  MUX2_X1 U377 ( .A(\mux[8][9] ), .B(\mux[9][9] ), .S(n523), .Z(n318) );
  MUX2_X1 U378 ( .A(n318), .B(n317), .S(n515), .Z(n319) );
  MUX2_X1 U379 ( .A(n319), .B(n316), .S(n510), .Z(n320) );
  MUX2_X1 U380 ( .A(\mux[6][9] ), .B(\mux[7][9] ), .S(addr_y[0]), .Z(n321) );
  MUX2_X1 U381 ( .A(\mux[4][9] ), .B(\mux[5][9] ), .S(n522), .Z(n322) );
  MUX2_X1 U382 ( .A(n322), .B(n321), .S(n514), .Z(n323) );
  MUX2_X1 U383 ( .A(\mux[2][9] ), .B(\mux[3][9] ), .S(n524), .Z(n324) );
  MUX2_X1 U384 ( .A(\mux[0][9] ), .B(\mux[1][9] ), .S(n523), .Z(n325) );
  MUX2_X1 U385 ( .A(n325), .B(n324), .S(n513), .Z(n326) );
  MUX2_X1 U386 ( .A(n326), .B(n323), .S(n510), .Z(n327) );
  MUX2_X1 U387 ( .A(n327), .B(n320), .S(n509), .Z(n328) );
  MUX2_X1 U388 ( .A(n328), .B(n313), .S(addr_y[4]), .Z(data_out[9]) );
  MUX2_X1 U389 ( .A(\mux[30][10] ), .B(\mux[31][10] ), .S(n521), .Z(n329) );
  MUX2_X1 U390 ( .A(\mux[28][10] ), .B(\mux[29][10] ), .S(n520), .Z(n330) );
  MUX2_X1 U391 ( .A(n330), .B(n329), .S(addr_y[1]), .Z(n331) );
  MUX2_X1 U392 ( .A(\mux[26][10] ), .B(\mux[27][10] ), .S(addr_y[0]), .Z(n332)
         );
  MUX2_X1 U393 ( .A(\mux[24][10] ), .B(\mux[25][10] ), .S(n526), .Z(n333) );
  MUX2_X1 U394 ( .A(n333), .B(n332), .S(addr_y[1]), .Z(n334) );
  MUX2_X1 U395 ( .A(n334), .B(n331), .S(n511), .Z(n335) );
  MUX2_X1 U396 ( .A(\mux[22][10] ), .B(\mux[23][10] ), .S(n518), .Z(n336) );
  MUX2_X1 U397 ( .A(\mux[20][10] ), .B(\mux[21][10] ), .S(n525), .Z(n337) );
  MUX2_X1 U398 ( .A(n337), .B(n336), .S(n512), .Z(n338) );
  MUX2_X1 U399 ( .A(\mux[18][10] ), .B(\mux[19][10] ), .S(n527), .Z(n339) );
  MUX2_X1 U400 ( .A(\mux[16][10] ), .B(\mux[17][10] ), .S(n517), .Z(n340) );
  MUX2_X1 U401 ( .A(n340), .B(n339), .S(n513), .Z(n341) );
  MUX2_X1 U402 ( .A(n341), .B(n338), .S(n511), .Z(n342) );
  MUX2_X1 U403 ( .A(n342), .B(n335), .S(addr_y[3]), .Z(n343) );
  MUX2_X1 U404 ( .A(\mux[14][10] ), .B(\mux[15][10] ), .S(n520), .Z(n344) );
  MUX2_X1 U405 ( .A(\mux[12][10] ), .B(\mux[13][10] ), .S(n518), .Z(n345) );
  MUX2_X1 U406 ( .A(n345), .B(n344), .S(n516), .Z(n346) );
  MUX2_X1 U407 ( .A(\mux[10][10] ), .B(\mux[11][10] ), .S(n522), .Z(n347) );
  MUX2_X1 U408 ( .A(\mux[8][10] ), .B(\mux[9][10] ), .S(n524), .Z(n348) );
  MUX2_X1 U409 ( .A(n348), .B(n347), .S(n515), .Z(n349) );
  MUX2_X1 U410 ( .A(n349), .B(n346), .S(n511), .Z(n350) );
  MUX2_X1 U411 ( .A(\mux[6][10] ), .B(\mux[7][10] ), .S(n519), .Z(n351) );
  MUX2_X1 U412 ( .A(\mux[4][10] ), .B(\mux[5][10] ), .S(n523), .Z(n352) );
  MUX2_X1 U413 ( .A(n352), .B(n351), .S(n514), .Z(n353) );
  MUX2_X1 U414 ( .A(\mux[2][10] ), .B(\mux[3][10] ), .S(addr_y[0]), .Z(n354)
         );
  MUX2_X1 U415 ( .A(\mux[0][10] ), .B(\mux[1][10] ), .S(n518), .Z(n355) );
  MUX2_X1 U416 ( .A(n355), .B(n354), .S(n516), .Z(n356) );
  MUX2_X1 U417 ( .A(n356), .B(n353), .S(n511), .Z(n357) );
  MUX2_X1 U418 ( .A(n357), .B(n350), .S(addr_y[3]), .Z(n358) );
  MUX2_X1 U419 ( .A(n358), .B(n343), .S(addr_y[4]), .Z(data_out[10]) );
  MUX2_X1 U420 ( .A(\mux[30][11] ), .B(\mux[31][11] ), .S(n525), .Z(n359) );
  MUX2_X1 U421 ( .A(\mux[28][11] ), .B(\mux[29][11] ), .S(n527), .Z(n360) );
  MUX2_X1 U422 ( .A(n360), .B(n359), .S(addr_y[1]), .Z(n361) );
  MUX2_X1 U423 ( .A(\mux[26][11] ), .B(\mux[27][11] ), .S(n526), .Z(n362) );
  MUX2_X1 U424 ( .A(\mux[24][11] ), .B(\mux[25][11] ), .S(n517), .Z(n363) );
  MUX2_X1 U425 ( .A(n363), .B(n362), .S(addr_y[1]), .Z(n364) );
  MUX2_X1 U426 ( .A(n364), .B(n361), .S(n511), .Z(n365) );
  MUX2_X1 U427 ( .A(\mux[22][11] ), .B(\mux[23][11] ), .S(n519), .Z(n366) );
  MUX2_X1 U428 ( .A(\mux[20][11] ), .B(\mux[21][11] ), .S(n526), .Z(n367) );
  MUX2_X1 U429 ( .A(n367), .B(n366), .S(n512), .Z(n368) );
  MUX2_X1 U430 ( .A(\mux[18][11] ), .B(\mux[19][11] ), .S(n522), .Z(n369) );
  MUX2_X1 U431 ( .A(\mux[16][11] ), .B(\mux[17][11] ), .S(n524), .Z(n370) );
  MUX2_X1 U432 ( .A(n370), .B(n369), .S(n513), .Z(n371) );
  MUX2_X1 U433 ( .A(n371), .B(n368), .S(n511), .Z(n372) );
  MUX2_X1 U434 ( .A(n372), .B(n365), .S(addr_y[3]), .Z(n373) );
  MUX2_X1 U435 ( .A(\mux[14][11] ), .B(\mux[15][11] ), .S(n519), .Z(n374) );
  MUX2_X1 U436 ( .A(\mux[12][11] ), .B(\mux[13][11] ), .S(n519), .Z(n375) );
  MUX2_X1 U437 ( .A(n375), .B(n374), .S(addr_y[1]), .Z(n376) );
  MUX2_X1 U438 ( .A(\mux[10][11] ), .B(\mux[11][11] ), .S(n519), .Z(n377) );
  MUX2_X1 U439 ( .A(\mux[8][11] ), .B(\mux[9][11] ), .S(n519), .Z(n378) );
  MUX2_X1 U440 ( .A(n378), .B(n377), .S(addr_y[1]), .Z(n379) );
  MUX2_X1 U441 ( .A(n379), .B(n376), .S(n511), .Z(n380) );
  MUX2_X1 U442 ( .A(\mux[6][11] ), .B(\mux[7][11] ), .S(n519), .Z(n381) );
  MUX2_X1 U443 ( .A(\mux[4][11] ), .B(\mux[5][11] ), .S(n519), .Z(n382) );
  MUX2_X1 U444 ( .A(n382), .B(n381), .S(addr_y[1]), .Z(n383) );
  MUX2_X1 U445 ( .A(\mux[2][11] ), .B(\mux[3][11] ), .S(n519), .Z(n384) );
  MUX2_X1 U446 ( .A(\mux[0][11] ), .B(\mux[1][11] ), .S(n519), .Z(n385) );
  MUX2_X1 U447 ( .A(n385), .B(n384), .S(n516), .Z(n386) );
  MUX2_X1 U448 ( .A(n386), .B(n383), .S(n511), .Z(n387) );
  MUX2_X1 U449 ( .A(n387), .B(n380), .S(addr_y[3]), .Z(n388) );
  MUX2_X1 U450 ( .A(n388), .B(n373), .S(addr_y[4]), .Z(data_out[11]) );
  MUX2_X1 U451 ( .A(\mux[30][12] ), .B(\mux[31][12] ), .S(n519), .Z(n389) );
  MUX2_X1 U452 ( .A(\mux[28][12] ), .B(\mux[29][12] ), .S(n519), .Z(n390) );
  MUX2_X1 U453 ( .A(n390), .B(n389), .S(addr_y[1]), .Z(n391) );
  MUX2_X1 U454 ( .A(\mux[26][12] ), .B(\mux[27][12] ), .S(n519), .Z(n392) );
  MUX2_X1 U455 ( .A(\mux[24][12] ), .B(\mux[25][12] ), .S(n519), .Z(n393) );
  MUX2_X1 U456 ( .A(n393), .B(n392), .S(n516), .Z(n394) );
  MUX2_X1 U457 ( .A(n394), .B(n391), .S(n511), .Z(n395) );
  MUX2_X1 U458 ( .A(\mux[22][12] ), .B(\mux[23][12] ), .S(n520), .Z(n396) );
  MUX2_X1 U459 ( .A(\mux[20][12] ), .B(\mux[21][12] ), .S(n520), .Z(n397) );
  MUX2_X1 U460 ( .A(n397), .B(n396), .S(n516), .Z(n398) );
  MUX2_X1 U461 ( .A(\mux[18][12] ), .B(\mux[19][12] ), .S(n520), .Z(n399) );
  MUX2_X1 U462 ( .A(\mux[16][12] ), .B(\mux[17][12] ), .S(n520), .Z(n400) );
  MUX2_X1 U463 ( .A(n400), .B(n399), .S(n515), .Z(n401) );
  MUX2_X1 U464 ( .A(n401), .B(n398), .S(n511), .Z(n402) );
  MUX2_X1 U465 ( .A(n402), .B(n395), .S(n509), .Z(n403) );
  MUX2_X1 U466 ( .A(\mux[14][12] ), .B(\mux[15][12] ), .S(n520), .Z(n404) );
  MUX2_X1 U467 ( .A(\mux[12][12] ), .B(\mux[13][12] ), .S(n520), .Z(n405) );
  MUX2_X1 U468 ( .A(n405), .B(n404), .S(addr_y[1]), .Z(n406) );
  MUX2_X1 U469 ( .A(\mux[10][12] ), .B(\mux[11][12] ), .S(n520), .Z(n407) );
  MUX2_X1 U470 ( .A(\mux[8][12] ), .B(\mux[9][12] ), .S(n520), .Z(n408) );
  MUX2_X1 U471 ( .A(n408), .B(n407), .S(n516), .Z(n409) );
  MUX2_X1 U472 ( .A(n409), .B(n406), .S(n511), .Z(n410) );
  MUX2_X1 U473 ( .A(\mux[6][12] ), .B(\mux[7][12] ), .S(n520), .Z(n411) );
  MUX2_X1 U474 ( .A(\mux[4][12] ), .B(\mux[5][12] ), .S(n520), .Z(n412) );
  MUX2_X1 U475 ( .A(n412), .B(n411), .S(n516), .Z(n413) );
  MUX2_X1 U476 ( .A(\mux[2][12] ), .B(\mux[3][12] ), .S(n520), .Z(n414) );
  MUX2_X1 U477 ( .A(\mux[0][12] ), .B(\mux[1][12] ), .S(n520), .Z(n415) );
  MUX2_X1 U478 ( .A(n415), .B(n414), .S(n514), .Z(n416) );
  MUX2_X1 U479 ( .A(n416), .B(n413), .S(n511), .Z(n417) );
  MUX2_X1 U480 ( .A(n417), .B(n410), .S(addr_y[3]), .Z(n418) );
  MUX2_X1 U481 ( .A(n418), .B(n403), .S(addr_y[4]), .Z(data_out[12]) );
  MUX2_X1 U482 ( .A(\mux[30][13] ), .B(\mux[31][13] ), .S(n521), .Z(n419) );
  MUX2_X1 U483 ( .A(\mux[28][13] ), .B(\mux[29][13] ), .S(n521), .Z(n420) );
  MUX2_X1 U484 ( .A(n420), .B(n419), .S(addr_y[1]), .Z(n421) );
  MUX2_X1 U485 ( .A(\mux[26][13] ), .B(\mux[27][13] ), .S(n521), .Z(n422) );
  MUX2_X1 U486 ( .A(\mux[24][13] ), .B(\mux[25][13] ), .S(n521), .Z(n423) );
  MUX2_X1 U487 ( .A(n423), .B(n422), .S(addr_y[1]), .Z(n424) );
  MUX2_X1 U488 ( .A(n424), .B(n421), .S(addr_y[2]), .Z(n425) );
  MUX2_X1 U489 ( .A(\mux[22][13] ), .B(\mux[23][13] ), .S(n521), .Z(n426) );
  MUX2_X1 U490 ( .A(\mux[20][13] ), .B(\mux[21][13] ), .S(n521), .Z(n427) );
  MUX2_X1 U491 ( .A(n427), .B(n426), .S(n516), .Z(n428) );
  MUX2_X1 U492 ( .A(\mux[18][13] ), .B(\mux[19][13] ), .S(n521), .Z(n429) );
  MUX2_X1 U493 ( .A(\mux[16][13] ), .B(\mux[17][13] ), .S(n521), .Z(n430) );
  MUX2_X1 U494 ( .A(n430), .B(n429), .S(addr_y[1]), .Z(n431) );
  MUX2_X1 U495 ( .A(n431), .B(n428), .S(n510), .Z(n432) );
  MUX2_X1 U496 ( .A(n432), .B(n425), .S(n509), .Z(n433) );
  MUX2_X1 U497 ( .A(\mux[14][13] ), .B(\mux[15][13] ), .S(n521), .Z(n434) );
  MUX2_X1 U498 ( .A(\mux[12][13] ), .B(\mux[13][13] ), .S(n521), .Z(n435) );
  MUX2_X1 U499 ( .A(n435), .B(n434), .S(addr_y[1]), .Z(n436) );
  MUX2_X1 U500 ( .A(\mux[10][13] ), .B(\mux[11][13] ), .S(n521), .Z(n437) );
  MUX2_X1 U501 ( .A(\mux[8][13] ), .B(\mux[9][13] ), .S(n521), .Z(n438) );
  MUX2_X1 U502 ( .A(n438), .B(n437), .S(n516), .Z(n439) );
  MUX2_X1 U503 ( .A(n439), .B(n436), .S(n511), .Z(n440) );
  MUX2_X1 U504 ( .A(\mux[6][13] ), .B(\mux[7][13] ), .S(n522), .Z(n441) );
  MUX2_X1 U505 ( .A(\mux[4][13] ), .B(\mux[5][13] ), .S(n522), .Z(n442) );
  MUX2_X1 U506 ( .A(n442), .B(n441), .S(addr_y[1]), .Z(n443) );
  MUX2_X1 U507 ( .A(\mux[2][13] ), .B(\mux[3][13] ), .S(n522), .Z(n444) );
  MUX2_X1 U508 ( .A(\mux[0][13] ), .B(\mux[1][13] ), .S(n522), .Z(n445) );
  MUX2_X1 U509 ( .A(n445), .B(n444), .S(addr_y[1]), .Z(n446) );
  MUX2_X1 U510 ( .A(n446), .B(n443), .S(addr_y[2]), .Z(n447) );
  MUX2_X1 U511 ( .A(n447), .B(n440), .S(addr_y[3]), .Z(n448) );
  MUX2_X1 U512 ( .A(n448), .B(n433), .S(addr_y[4]), .Z(data_out[13]) );
  MUX2_X1 U513 ( .A(\mux[30][14] ), .B(\mux[31][14] ), .S(n522), .Z(n449) );
  MUX2_X1 U514 ( .A(\mux[28][14] ), .B(\mux[29][14] ), .S(n522), .Z(n450) );
  MUX2_X1 U515 ( .A(n450), .B(n449), .S(n516), .Z(n451) );
  MUX2_X1 U516 ( .A(\mux[26][14] ), .B(\mux[27][14] ), .S(n522), .Z(n452) );
  MUX2_X1 U517 ( .A(\mux[24][14] ), .B(\mux[25][14] ), .S(n522), .Z(n453) );
  MUX2_X1 U518 ( .A(n453), .B(n452), .S(n516), .Z(n454) );
  MUX2_X1 U519 ( .A(n454), .B(n451), .S(n510), .Z(n455) );
  MUX2_X1 U520 ( .A(\mux[22][14] ), .B(\mux[23][14] ), .S(n522), .Z(n456) );
  MUX2_X1 U521 ( .A(\mux[20][14] ), .B(\mux[21][14] ), .S(n522), .Z(n457) );
  MUX2_X1 U522 ( .A(n457), .B(n456), .S(addr_y[1]), .Z(n458) );
  MUX2_X1 U523 ( .A(\mux[18][14] ), .B(\mux[19][14] ), .S(n522), .Z(n459) );
  MUX2_X1 U524 ( .A(\mux[16][14] ), .B(\mux[17][14] ), .S(n522), .Z(n460) );
  MUX2_X1 U525 ( .A(n460), .B(n459), .S(n516), .Z(n461) );
  MUX2_X1 U526 ( .A(n461), .B(n458), .S(n511), .Z(n462) );
  MUX2_X1 U527 ( .A(n462), .B(n455), .S(n509), .Z(n463) );
  MUX2_X1 U528 ( .A(\mux[14][14] ), .B(\mux[15][14] ), .S(n523), .Z(n464) );
  MUX2_X1 U529 ( .A(\mux[12][14] ), .B(\mux[13][14] ), .S(n523), .Z(n465) );
  MUX2_X1 U530 ( .A(n465), .B(n464), .S(n515), .Z(n466) );
  MUX2_X1 U531 ( .A(\mux[10][14] ), .B(\mux[11][14] ), .S(n523), .Z(n467) );
  MUX2_X1 U532 ( .A(\mux[8][14] ), .B(\mux[9][14] ), .S(n523), .Z(n468) );
  MUX2_X1 U533 ( .A(n468), .B(n467), .S(n515), .Z(n469) );
  MUX2_X1 U534 ( .A(n469), .B(n466), .S(addr_y[2]), .Z(n470) );
  MUX2_X1 U535 ( .A(\mux[6][14] ), .B(\mux[7][14] ), .S(n523), .Z(n471) );
  MUX2_X1 U536 ( .A(\mux[4][14] ), .B(\mux[5][14] ), .S(n523), .Z(n472) );
  MUX2_X1 U537 ( .A(n472), .B(n471), .S(n515), .Z(n473) );
  MUX2_X1 U538 ( .A(\mux[2][14] ), .B(\mux[3][14] ), .S(n523), .Z(n474) );
  MUX2_X1 U539 ( .A(\mux[0][14] ), .B(\mux[1][14] ), .S(n523), .Z(n475) );
  MUX2_X1 U540 ( .A(n475), .B(n474), .S(n515), .Z(n476) );
  MUX2_X1 U541 ( .A(n476), .B(n473), .S(n510), .Z(n477) );
  MUX2_X1 U542 ( .A(n477), .B(n470), .S(addr_y[3]), .Z(n478) );
  MUX2_X1 U543 ( .A(n478), .B(n463), .S(addr_y[4]), .Z(data_out[14]) );
  MUX2_X1 U544 ( .A(\mux[30][15] ), .B(\mux[31][15] ), .S(n523), .Z(n479) );
  MUX2_X1 U545 ( .A(\mux[28][15] ), .B(\mux[29][15] ), .S(n523), .Z(n480) );
  MUX2_X1 U546 ( .A(n480), .B(n479), .S(n515), .Z(n481) );
  MUX2_X1 U547 ( .A(\mux[26][15] ), .B(\mux[27][15] ), .S(n523), .Z(n482) );
  MUX2_X1 U548 ( .A(\mux[24][15] ), .B(\mux[25][15] ), .S(n523), .Z(n483) );
  MUX2_X1 U549 ( .A(n483), .B(n482), .S(n515), .Z(n484) );
  MUX2_X1 U550 ( .A(n484), .B(n481), .S(n511), .Z(n485) );
  MUX2_X1 U551 ( .A(\mux[22][15] ), .B(\mux[23][15] ), .S(n524), .Z(n486) );
  MUX2_X1 U552 ( .A(\mux[20][15] ), .B(\mux[21][15] ), .S(n524), .Z(n487) );
  MUX2_X1 U553 ( .A(n487), .B(n486), .S(n515), .Z(n488) );
  MUX2_X1 U554 ( .A(\mux[18][15] ), .B(\mux[19][15] ), .S(n524), .Z(n489) );
  MUX2_X1 U555 ( .A(\mux[16][15] ), .B(\mux[17][15] ), .S(n524), .Z(n490) );
  MUX2_X1 U556 ( .A(n490), .B(n489), .S(n515), .Z(n491) );
  MUX2_X1 U557 ( .A(n491), .B(n488), .S(addr_y[2]), .Z(n492) );
  MUX2_X1 U558 ( .A(n492), .B(n485), .S(n509), .Z(n493) );
  MUX2_X1 U559 ( .A(\mux[14][15] ), .B(\mux[15][15] ), .S(n524), .Z(n494) );
  MUX2_X1 U560 ( .A(\mux[12][15] ), .B(\mux[13][15] ), .S(n524), .Z(n495) );
  MUX2_X1 U561 ( .A(n495), .B(n494), .S(n515), .Z(n496) );
  MUX2_X1 U562 ( .A(\mux[10][15] ), .B(\mux[11][15] ), .S(n524), .Z(n497) );
  MUX2_X1 U563 ( .A(\mux[8][15] ), .B(\mux[9][15] ), .S(n524), .Z(n498) );
  MUX2_X1 U564 ( .A(n498), .B(n497), .S(n515), .Z(n499) );
  MUX2_X1 U565 ( .A(n499), .B(n496), .S(n510), .Z(n500) );
  MUX2_X1 U566 ( .A(\mux[6][15] ), .B(\mux[7][15] ), .S(n524), .Z(n501) );
  MUX2_X1 U567 ( .A(\mux[4][15] ), .B(\mux[5][15] ), .S(n524), .Z(n502) );
  MUX2_X1 U568 ( .A(n502), .B(n501), .S(n515), .Z(n503) );
  MUX2_X1 U569 ( .A(\mux[2][15] ), .B(\mux[3][15] ), .S(n524), .Z(n504) );
  MUX2_X1 U570 ( .A(\mux[0][15] ), .B(\mux[1][15] ), .S(n524), .Z(n505) );
  MUX2_X1 U571 ( .A(n505), .B(n504), .S(n515), .Z(n506) );
  MUX2_X1 U572 ( .A(n506), .B(n503), .S(n511), .Z(n507) );
  MUX2_X1 U573 ( .A(n507), .B(n500), .S(addr_y[3]), .Z(n508) );
  MUX2_X1 U574 ( .A(n508), .B(n493), .S(addr_y[4]), .Z(data_out[15]) );
  CLKBUF_X3 U575 ( .A(vector_out[0]), .Z(n536) );
  CLKBUF_X3 U576 ( .A(vector_out[5]), .Z(n551) );
  CLKBUF_X3 U577 ( .A(vector_out[7]), .Z(n556) );
endmodule


module mvm_32_32_8_1 ( clk, reset, loadMatrix, loadVector, start, done, 
        data_in, data_out );
  input [7:0] data_in;
  output [15:0] data_out;
  input clk, reset, loadMatrix, loadVector, start;
  output done;
  wire   wr_en_x, clear_acc, wr_en_y, \addr_a[31][4] , \addr_a[31][3] ,
         \addr_a[31][2] , \addr_a[31][1] , \addr_a[31][0] , \addr_a[30][4] ,
         \addr_a[30][3] , \addr_a[30][2] , \addr_a[30][1] , \addr_a[30][0] ,
         \addr_a[29][4] , \addr_a[29][3] , \addr_a[29][2] , \addr_a[29][1] ,
         \addr_a[29][0] , \addr_a[28][4] , \addr_a[28][3] , \addr_a[28][2] ,
         \addr_a[28][1] , \addr_a[28][0] , \addr_a[27][4] , \addr_a[27][3] ,
         \addr_a[27][2] , \addr_a[27][1] , \addr_a[27][0] , \addr_a[26][4] ,
         \addr_a[26][3] , \addr_a[26][2] , \addr_a[26][1] , \addr_a[26][0] ,
         \addr_a[25][4] , \addr_a[25][3] , \addr_a[25][2] , \addr_a[25][1] ,
         \addr_a[25][0] , \addr_a[24][4] , \addr_a[24][3] , \addr_a[24][2] ,
         \addr_a[24][1] , \addr_a[24][0] , \addr_a[23][4] , \addr_a[23][3] ,
         \addr_a[23][2] , \addr_a[23][1] , \addr_a[23][0] , \addr_a[22][4] ,
         \addr_a[22][3] , \addr_a[22][2] , \addr_a[22][1] , \addr_a[22][0] ,
         \addr_a[21][4] , \addr_a[21][3] , \addr_a[21][2] , \addr_a[21][1] ,
         \addr_a[21][0] , \addr_a[20][4] , \addr_a[20][3] , \addr_a[20][2] ,
         \addr_a[20][1] , \addr_a[20][0] , \addr_a[19][4] , \addr_a[19][3] ,
         \addr_a[19][2] , \addr_a[19][1] , \addr_a[19][0] , \addr_a[18][4] ,
         \addr_a[18][3] , \addr_a[18][2] , \addr_a[18][1] , \addr_a[18][0] ,
         \addr_a[17][4] , \addr_a[17][3] , \addr_a[17][2] , \addr_a[17][1] ,
         \addr_a[17][0] , \addr_a[16][4] , \addr_a[16][3] , \addr_a[16][2] ,
         \addr_a[16][1] , \addr_a[16][0] , \addr_a[15][4] , \addr_a[15][3] ,
         \addr_a[15][2] , \addr_a[15][1] , \addr_a[15][0] , \addr_a[14][4] ,
         \addr_a[14][3] , \addr_a[14][2] , \addr_a[14][1] , \addr_a[14][0] ,
         \addr_a[13][4] , \addr_a[13][3] , \addr_a[13][2] , \addr_a[13][1] ,
         \addr_a[13][0] , \addr_a[12][4] , \addr_a[12][3] , \addr_a[12][2] ,
         \addr_a[12][1] , \addr_a[12][0] , \addr_a[11][4] , \addr_a[11][3] ,
         \addr_a[11][2] , \addr_a[11][1] , \addr_a[11][0] , \addr_a[10][4] ,
         \addr_a[10][3] , \addr_a[10][2] , \addr_a[10][1] , \addr_a[10][0] ,
         \addr_a[9][4] , \addr_a[9][3] , \addr_a[9][2] , \addr_a[9][1] ,
         \addr_a[9][0] , \addr_a[8][4] , \addr_a[8][3] , \addr_a[8][2] ,
         \addr_a[8][1] , \addr_a[8][0] , \addr_a[7][4] , \addr_a[7][3] ,
         \addr_a[7][2] , \addr_a[7][1] , \addr_a[7][0] , \addr_a[6][4] ,
         \addr_a[6][3] , \addr_a[6][2] , \addr_a[6][1] , \addr_a[6][0] ,
         \addr_a[5][4] , \addr_a[5][3] , \addr_a[5][2] , \addr_a[5][1] ,
         \addr_a[5][0] , \addr_a[4][4] , \addr_a[4][3] , \addr_a[4][2] ,
         \addr_a[4][1] , \addr_a[4][0] , \addr_a[3][4] , \addr_a[3][3] ,
         \addr_a[3][2] , \addr_a[3][1] , \addr_a[3][0] , \addr_a[2][4] ,
         \addr_a[2][3] , \addr_a[2][2] , \addr_a[2][1] , \addr_a[2][0] ,
         \addr_a[1][4] , \addr_a[1][3] , \addr_a[1][2] , \addr_a[1][1] ,
         \addr_a[1][0] , \addr_a[0][4] , \addr_a[0][3] , \addr_a[0][2] ,
         \addr_a[0][1] , \addr_a[0][0] ;
  wire   [5:0] addr_x;
  wire   [5:0] addr_y;
  wire   [31:0] wr_en_a;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32;

  controlpath c ( .clk(clk), .reset(reset), .start(start), .loadMatrix(
        loadMatrix), .loadVector(loadVector), .wr_en_x(wr_en_x), .clear_acc(
        clear_acc), .wr_en_y(wr_en_y), .done(done), .addr_x({
        SYNOPSYS_UNCONNECTED__0, addr_x[4:0]}), .addr_y(addr_y), .addr_a({
        SYNOPSYS_UNCONNECTED__1, \addr_a[31][4] , \addr_a[31][3] , 
        \addr_a[31][2] , \addr_a[31][1] , \addr_a[31][0] , 
        SYNOPSYS_UNCONNECTED__2, \addr_a[30][4] , \addr_a[30][3] , 
        \addr_a[30][2] , \addr_a[30][1] , \addr_a[30][0] , 
        SYNOPSYS_UNCONNECTED__3, \addr_a[29][4] , \addr_a[29][3] , 
        \addr_a[29][2] , \addr_a[29][1] , \addr_a[29][0] , 
        SYNOPSYS_UNCONNECTED__4, \addr_a[28][4] , \addr_a[28][3] , 
        \addr_a[28][2] , \addr_a[28][1] , \addr_a[28][0] , 
        SYNOPSYS_UNCONNECTED__5, \addr_a[27][4] , \addr_a[27][3] , 
        \addr_a[27][2] , \addr_a[27][1] , \addr_a[27][0] , 
        SYNOPSYS_UNCONNECTED__6, \addr_a[26][4] , \addr_a[26][3] , 
        \addr_a[26][2] , \addr_a[26][1] , \addr_a[26][0] , 
        SYNOPSYS_UNCONNECTED__7, \addr_a[25][4] , \addr_a[25][3] , 
        \addr_a[25][2] , \addr_a[25][1] , \addr_a[25][0] , 
        SYNOPSYS_UNCONNECTED__8, \addr_a[24][4] , \addr_a[24][3] , 
        \addr_a[24][2] , \addr_a[24][1] , \addr_a[24][0] , 
        SYNOPSYS_UNCONNECTED__9, \addr_a[23][4] , \addr_a[23][3] , 
        \addr_a[23][2] , \addr_a[23][1] , \addr_a[23][0] , 
        SYNOPSYS_UNCONNECTED__10, \addr_a[22][4] , \addr_a[22][3] , 
        \addr_a[22][2] , \addr_a[22][1] , \addr_a[22][0] , 
        SYNOPSYS_UNCONNECTED__11, \addr_a[21][4] , \addr_a[21][3] , 
        \addr_a[21][2] , \addr_a[21][1] , \addr_a[21][0] , 
        SYNOPSYS_UNCONNECTED__12, \addr_a[20][4] , \addr_a[20][3] , 
        \addr_a[20][2] , \addr_a[20][1] , \addr_a[20][0] , 
        SYNOPSYS_UNCONNECTED__13, \addr_a[19][4] , \addr_a[19][3] , 
        \addr_a[19][2] , \addr_a[19][1] , \addr_a[19][0] , 
        SYNOPSYS_UNCONNECTED__14, \addr_a[18][4] , \addr_a[18][3] , 
        \addr_a[18][2] , \addr_a[18][1] , \addr_a[18][0] , 
        SYNOPSYS_UNCONNECTED__15, \addr_a[17][4] , \addr_a[17][3] , 
        \addr_a[17][2] , \addr_a[17][1] , \addr_a[17][0] , 
        SYNOPSYS_UNCONNECTED__16, \addr_a[16][4] , \addr_a[16][3] , 
        \addr_a[16][2] , \addr_a[16][1] , \addr_a[16][0] , 
        SYNOPSYS_UNCONNECTED__17, \addr_a[15][4] , \addr_a[15][3] , 
        \addr_a[15][2] , \addr_a[15][1] , \addr_a[15][0] , 
        SYNOPSYS_UNCONNECTED__18, \addr_a[14][4] , \addr_a[14][3] , 
        \addr_a[14][2] , \addr_a[14][1] , \addr_a[14][0] , 
        SYNOPSYS_UNCONNECTED__19, \addr_a[13][4] , \addr_a[13][3] , 
        \addr_a[13][2] , \addr_a[13][1] , \addr_a[13][0] , 
        SYNOPSYS_UNCONNECTED__20, \addr_a[12][4] , \addr_a[12][3] , 
        \addr_a[12][2] , \addr_a[12][1] , \addr_a[12][0] , 
        SYNOPSYS_UNCONNECTED__21, \addr_a[11][4] , \addr_a[11][3] , 
        \addr_a[11][2] , \addr_a[11][1] , \addr_a[11][0] , 
        SYNOPSYS_UNCONNECTED__22, \addr_a[10][4] , \addr_a[10][3] , 
        \addr_a[10][2] , \addr_a[10][1] , \addr_a[10][0] , 
        SYNOPSYS_UNCONNECTED__23, \addr_a[9][4] , \addr_a[9][3] , 
        \addr_a[9][2] , \addr_a[9][1] , \addr_a[9][0] , 
        SYNOPSYS_UNCONNECTED__24, \addr_a[8][4] , \addr_a[8][3] , 
        \addr_a[8][2] , \addr_a[8][1] , \addr_a[8][0] , 
        SYNOPSYS_UNCONNECTED__25, \addr_a[7][4] , \addr_a[7][3] , 
        \addr_a[7][2] , \addr_a[7][1] , \addr_a[7][0] , 
        SYNOPSYS_UNCONNECTED__26, \addr_a[6][4] , \addr_a[6][3] , 
        \addr_a[6][2] , \addr_a[6][1] , \addr_a[6][0] , 
        SYNOPSYS_UNCONNECTED__27, \addr_a[5][4] , \addr_a[5][3] , 
        \addr_a[5][2] , \addr_a[5][1] , \addr_a[5][0] , 
        SYNOPSYS_UNCONNECTED__28, \addr_a[4][4] , \addr_a[4][3] , 
        \addr_a[4][2] , \addr_a[4][1] , \addr_a[4][0] , 
        SYNOPSYS_UNCONNECTED__29, \addr_a[3][4] , \addr_a[3][3] , 
        \addr_a[3][2] , \addr_a[3][1] , \addr_a[3][0] , 
        SYNOPSYS_UNCONNECTED__30, \addr_a[2][4] , \addr_a[2][3] , 
        \addr_a[2][2] , \addr_a[2][1] , \addr_a[2][0] , 
        SYNOPSYS_UNCONNECTED__31, \addr_a[1][4] , \addr_a[1][3] , 
        \addr_a[1][2] , \addr_a[1][1] , \addr_a[1][0] , 
        SYNOPSYS_UNCONNECTED__32, \addr_a[0][4] , \addr_a[0][3] , 
        \addr_a[0][2] , \addr_a[0][1] , \addr_a[0][0] }), .wr_en_a(wr_en_a) );
  datapath d ( .clk(clk), .wr_en_x(wr_en_x), .clear_acc(clear_acc), .wr_en_y(
        wr_en_y), .addr_x({1'b0, addr_x[4:0]}), .addr_y(addr_y), .addr_a({1'b0, 
        \addr_a[31][4] , \addr_a[31][3] , \addr_a[31][2] , \addr_a[31][1] , 
        \addr_a[31][0] , 1'b0, \addr_a[30][4] , \addr_a[30][3] , 
        \addr_a[30][2] , \addr_a[30][1] , \addr_a[30][0] , 1'b0, 
        \addr_a[29][4] , \addr_a[29][3] , \addr_a[29][2] , \addr_a[29][1] , 
        \addr_a[29][0] , 1'b0, \addr_a[28][4] , \addr_a[28][3] , 
        \addr_a[28][2] , \addr_a[28][1] , \addr_a[28][0] , 1'b0, 
        \addr_a[27][4] , \addr_a[27][3] , \addr_a[27][2] , \addr_a[27][1] , 
        \addr_a[27][0] , 1'b0, \addr_a[26][4] , \addr_a[26][3] , 
        \addr_a[26][2] , \addr_a[26][1] , \addr_a[26][0] , 1'b0, 
        \addr_a[25][4] , \addr_a[25][3] , \addr_a[25][2] , \addr_a[25][1] , 
        \addr_a[25][0] , 1'b0, \addr_a[24][4] , \addr_a[24][3] , 
        \addr_a[24][2] , \addr_a[24][1] , \addr_a[24][0] , 1'b0, 
        \addr_a[23][4] , \addr_a[23][3] , \addr_a[23][2] , \addr_a[23][1] , 
        \addr_a[23][0] , 1'b0, \addr_a[22][4] , \addr_a[22][3] , 
        \addr_a[22][2] , \addr_a[22][1] , \addr_a[22][0] , 1'b0, 
        \addr_a[21][4] , \addr_a[21][3] , \addr_a[21][2] , \addr_a[21][1] , 
        \addr_a[21][0] , 1'b0, \addr_a[20][4] , \addr_a[20][3] , 
        \addr_a[20][2] , \addr_a[20][1] , \addr_a[20][0] , 1'b0, 
        \addr_a[19][4] , \addr_a[19][3] , \addr_a[19][2] , \addr_a[19][1] , 
        \addr_a[19][0] , 1'b0, \addr_a[18][4] , \addr_a[18][3] , 
        \addr_a[18][2] , \addr_a[18][1] , \addr_a[18][0] , 1'b0, 
        \addr_a[17][4] , \addr_a[17][3] , \addr_a[17][2] , \addr_a[17][1] , 
        \addr_a[17][0] , 1'b0, \addr_a[16][4] , \addr_a[16][3] , 
        \addr_a[16][2] , \addr_a[16][1] , \addr_a[16][0] , 1'b0, 
        \addr_a[15][4] , \addr_a[15][3] , \addr_a[15][2] , \addr_a[15][1] , 
        \addr_a[15][0] , 1'b0, \addr_a[14][4] , \addr_a[14][3] , 
        \addr_a[14][2] , \addr_a[14][1] , \addr_a[14][0] , 1'b0, 
        \addr_a[13][4] , \addr_a[13][3] , \addr_a[13][2] , \addr_a[13][1] , 
        \addr_a[13][0] , 1'b0, \addr_a[12][4] , \addr_a[12][3] , 
        \addr_a[12][2] , \addr_a[12][1] , \addr_a[12][0] , 1'b0, 
        \addr_a[11][4] , \addr_a[11][3] , \addr_a[11][2] , \addr_a[11][1] , 
        \addr_a[11][0] , 1'b0, \addr_a[10][4] , \addr_a[10][3] , 
        \addr_a[10][2] , \addr_a[10][1] , \addr_a[10][0] , 1'b0, 
        \addr_a[9][4] , \addr_a[9][3] , \addr_a[9][2] , \addr_a[9][1] , 
        \addr_a[9][0] , 1'b0, \addr_a[8][4] , \addr_a[8][3] , \addr_a[8][2] , 
        \addr_a[8][1] , \addr_a[8][0] , 1'b0, \addr_a[7][4] , \addr_a[7][3] , 
        \addr_a[7][2] , \addr_a[7][1] , \addr_a[7][0] , 1'b0, \addr_a[6][4] , 
        \addr_a[6][3] , \addr_a[6][2] , \addr_a[6][1] , \addr_a[6][0] , 1'b0, 
        \addr_a[5][4] , \addr_a[5][3] , \addr_a[5][2] , \addr_a[5][1] , 
        \addr_a[5][0] , 1'b0, \addr_a[4][4] , \addr_a[4][3] , \addr_a[4][2] , 
        \addr_a[4][1] , \addr_a[4][0] , 1'b0, \addr_a[3][4] , \addr_a[3][3] , 
        \addr_a[3][2] , \addr_a[3][1] , \addr_a[3][0] , 1'b0, \addr_a[2][4] , 
        \addr_a[2][3] , \addr_a[2][2] , \addr_a[2][1] , \addr_a[2][0] , 1'b0, 
        \addr_a[1][4] , \addr_a[1][3] , \addr_a[1][2] , \addr_a[1][1] , 
        \addr_a[1][0] , 1'b0, \addr_a[0][4] , \addr_a[0][3] , \addr_a[0][2] , 
        \addr_a[0][1] , \addr_a[0][0] }), .data_in(data_in), .wr_en_a(wr_en_a), 
        .data_out(data_out) );
endmodule

