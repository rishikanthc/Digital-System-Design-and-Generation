
module controlpath ( clk, reset, start, loadMatrix, loadVector, wr_en_x, 
        clear_acc, wr_en_y, done, addr_x, addr_y, .addr_a({\addr_a[7][3] , 
        \addr_a[7][2] , \addr_a[7][1] , \addr_a[7][0] , \addr_a[6][3] , 
        \addr_a[6][2] , \addr_a[6][1] , \addr_a[6][0] , \addr_a[5][3] , 
        \addr_a[5][2] , \addr_a[5][1] , \addr_a[5][0] , \addr_a[4][3] , 
        \addr_a[4][2] , \addr_a[4][1] , \addr_a[4][0] , \addr_a[3][3] , 
        \addr_a[3][2] , \addr_a[3][1] , \addr_a[3][0] , \addr_a[2][3] , 
        \addr_a[2][2] , \addr_a[2][1] , \addr_a[2][0] , \addr_a[1][3] , 
        \addr_a[1][2] , \addr_a[1][1] , \addr_a[1][0] , \addr_a[0][3] , 
        \addr_a[0][2] , \addr_a[0][1] , \addr_a[0][0] }), wr_en_a );
  output [3:0] addr_x;
  output [3:0] addr_y;
  output [7:0] wr_en_a;
  input clk, reset, start, loadMatrix, loadVector;
  output wr_en_x, clear_acc, wr_en_y, done, \addr_a[7][3] , \addr_a[7][2] ,
         \addr_a[7][1] , \addr_a[7][0] , \addr_a[6][3] , \addr_a[6][2] ,
         \addr_a[6][1] , \addr_a[6][0] , \addr_a[5][3] , \addr_a[5][2] ,
         \addr_a[5][1] , \addr_a[5][0] , \addr_a[4][3] , \addr_a[4][2] ,
         \addr_a[4][1] , \addr_a[4][0] , \addr_a[3][3] , \addr_a[3][2] ,
         \addr_a[3][1] , \addr_a[3][0] , \addr_a[2][3] , \addr_a[2][2] ,
         \addr_a[2][1] , \addr_a[2][0] , \addr_a[1][3] , \addr_a[1][2] ,
         \addr_a[1][1] , \addr_a[1][0] , \addr_a[0][3] , \addr_a[0][2] ,
         \addr_a[0][1] , \addr_a[0][0] ;
  wire   N128, N129, N130, N136, N137, N138, N244, N245, N246, N247, N248, n23,
         n24, n26, n31, n38, n39, n40, n42, n43, n44, n46, n47, n48, n49, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n78, n79, n80,
         n81, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n25, n27, n28, n29, n30;
  wire   [2:0] state;
  wire   [3:0] counter;
  wire   [3:0] counter2;
  assign addr_y[3] = 1'b0;
  assign \addr_a[0][3]  = 1'b0;
  assign \addr_a[1][3]  = 1'b0;
  assign \addr_a[2][3]  = 1'b0;
  assign \addr_a[3][3]  = 1'b0;
  assign \addr_a[4][3]  = 1'b0;
  assign \addr_a[5][3]  = 1'b0;
  assign \addr_a[6][3]  = 1'b0;
  assign \addr_a[7][3]  = 1'b0;
  assign addr_x[3] = 1'b0;

  NOR4_X2 U6 ( .A1(n38), .A2(n39), .A3(n40), .A4(n11), .ZN(wr_en_y) );
  NAND3_X1 U137 ( .A1(n64), .A2(n6), .A3(n10), .ZN(n63) );
  NAND3_X1 U138 ( .A1(n72), .A2(n71), .A3(n73), .ZN(n66) );
  NAND3_X1 U139 ( .A1(state[1]), .A2(n23), .A3(state[0]), .ZN(n75) );
  NAND3_X1 U140 ( .A1(N244), .A2(n31), .A3(n86), .ZN(n53) );
  NAND3_X1 U142 ( .A1(n73), .A2(state[0]), .A3(n100), .ZN(n99) );
  NAND3_X1 U144 ( .A1(N244), .A2(n31), .A3(n91), .ZN(n42) );
  DFF_X1 \state_reg[1]  ( .D(N129), .CK(clk), .Q(state[1]), .QN(n24) );
  DFF_X1 \counter2_reg[2]  ( .D(N138), .CK(clk), .Q(counter2[2]), .QN(n12) );
  DFF_X1 \state_reg[2]  ( .D(N130), .CK(clk), .Q(state[2]), .QN(n23) );
  DFF_X1 \counter_reg[1]  ( .D(n102), .CK(clk), .Q(counter[1]), .QN(n31) );
  DFF_X1 \counter_reg[0]  ( .D(n104), .CK(clk), .Q(counter[0]), .QN(N244) );
  DFF_X1 \counter_reg[2]  ( .D(n101), .CK(clk), .Q(counter[2]), .QN(n6) );
  DFF_X1 \counter_reg[3]  ( .D(n103), .CK(clk), .Q(counter[3]), .QN(n26) );
  DFF_X1 \counter2_reg[1]  ( .D(N137), .CK(clk), .Q(counter2[1]), .QN(n11) );
  DFF_X1 \counter2_reg[0]  ( .D(N136), .CK(clk), .Q(counter2[0]), .QN(n7) );
  DFF_X1 \state_reg[0]  ( .D(N128), .CK(clk), .Q(state[0]) );
  NOR4_X1 U4 ( .A1(loadMatrix), .A2(loadVector), .A3(reset), .A4(start), .ZN(
        n73) );
  NOR2_X2 U5 ( .A1(n20), .A2(n12), .ZN(\addr_a[7][2] ) );
  NOR2_X2 U7 ( .A1(n13), .A2(n12), .ZN(\addr_a[0][2] ) );
  NOR2_X2 U8 ( .A1(n15), .A2(n12), .ZN(\addr_a[2][2] ) );
  NOR2_X2 U9 ( .A1(n16), .A2(n12), .ZN(\addr_a[3][2] ) );
  NOR2_X2 U10 ( .A1(n18), .A2(n12), .ZN(\addr_a[5][2] ) );
  NOR2_X2 U11 ( .A1(n19), .A2(n12), .ZN(\addr_a[6][2] ) );
  NOR2_X2 U12 ( .A1(n14), .A2(n12), .ZN(\addr_a[1][2] ) );
  NOR2_X2 U13 ( .A1(n17), .A2(n12), .ZN(\addr_a[4][2] ) );
  NOR2_X1 U14 ( .A1(n81), .A2(n12), .ZN(addr_x[2]) );
  INV_X1 U15 ( .A(n71), .ZN(n10) );
  NOR2_X1 U16 ( .A1(n95), .A2(n80), .ZN(N137) );
  NOR3_X1 U17 ( .A1(n1), .A2(n38), .A3(n59), .ZN(done) );
  OAI21_X1 U18 ( .B1(n64), .B2(n71), .A(n66), .ZN(n65) );
  NAND2_X1 U19 ( .A1(n55), .A2(n25), .ZN(n58) );
  INV_X1 U20 ( .A(N246), .ZN(n25) );
  NAND2_X1 U21 ( .A1(N246), .A2(n55), .ZN(n46) );
  INV_X1 U22 ( .A(n76), .ZN(n21) );
  NAND2_X1 U23 ( .A1(n68), .A2(n91), .ZN(n59) );
  NAND2_X1 U24 ( .A1(n91), .A2(n69), .ZN(n40) );
  AND2_X1 U25 ( .A1(n22), .A2(n38), .ZN(n81) );
  INV_X1 U26 ( .A(n93), .ZN(n14) );
  OAI21_X1 U27 ( .B1(n40), .B2(n43), .A(n38), .ZN(n93) );
  INV_X1 U28 ( .A(n85), .ZN(n20) );
  OAI21_X1 U29 ( .B1(n47), .B2(n43), .A(n38), .ZN(n85) );
  INV_X1 U30 ( .A(n94), .ZN(n13) );
  OAI21_X1 U31 ( .B1(n42), .B2(n43), .A(n38), .ZN(n94) );
  INV_X1 U32 ( .A(n92), .ZN(n15) );
  OAI21_X1 U33 ( .B1(n43), .B2(n59), .A(n38), .ZN(n92) );
  INV_X1 U34 ( .A(n90), .ZN(n16) );
  OAI21_X1 U35 ( .B1(n43), .B2(n56), .A(n38), .ZN(n90) );
  INV_X1 U36 ( .A(n89), .ZN(n17) );
  OAI21_X1 U37 ( .B1(n43), .B2(n53), .A(n38), .ZN(n89) );
  INV_X1 U38 ( .A(n88), .ZN(n18) );
  OAI21_X1 U39 ( .B1(n43), .B2(n51), .A(n38), .ZN(n88) );
  INV_X1 U40 ( .A(n87), .ZN(n19) );
  OAI21_X1 U41 ( .B1(n43), .B2(n48), .A(n38), .ZN(n87) );
  NAND2_X1 U42 ( .A1(n64), .A2(n91), .ZN(n56) );
  NAND2_X1 U43 ( .A1(n86), .A2(n69), .ZN(n51) );
  NAND2_X1 U44 ( .A1(n86), .A2(n64), .ZN(n47) );
  NOR2_X1 U45 ( .A1(n14), .A2(n11), .ZN(\addr_a[1][1] ) );
  NOR2_X1 U46 ( .A1(n15), .A2(n11), .ZN(\addr_a[2][1] ) );
  NOR2_X1 U47 ( .A1(n16), .A2(n11), .ZN(\addr_a[3][1] ) );
  NOR2_X1 U48 ( .A1(n17), .A2(n11), .ZN(\addr_a[4][1] ) );
  NOR2_X1 U49 ( .A1(n18), .A2(n11), .ZN(\addr_a[5][1] ) );
  NOR2_X1 U50 ( .A1(n19), .A2(n11), .ZN(\addr_a[6][1] ) );
  NOR2_X1 U51 ( .A1(n20), .A2(n11), .ZN(\addr_a[7][1] ) );
  NOR2_X1 U52 ( .A1(n81), .A2(n11), .ZN(addr_x[1]) );
  NOR2_X1 U53 ( .A1(n13), .A2(n11), .ZN(\addr_a[0][1] ) );
  NOR2_X1 U54 ( .A1(n14), .A2(n7), .ZN(\addr_a[1][0] ) );
  NOR2_X1 U55 ( .A1(n15), .A2(n7), .ZN(\addr_a[2][0] ) );
  NOR2_X1 U56 ( .A1(n16), .A2(n7), .ZN(\addr_a[3][0] ) );
  NOR2_X1 U57 ( .A1(n17), .A2(n7), .ZN(\addr_a[4][0] ) );
  NOR2_X1 U58 ( .A1(n18), .A2(n7), .ZN(\addr_a[5][0] ) );
  NOR2_X1 U59 ( .A1(n19), .A2(n7), .ZN(\addr_a[6][0] ) );
  NOR2_X1 U60 ( .A1(n20), .A2(n7), .ZN(\addr_a[7][0] ) );
  NOR2_X1 U61 ( .A1(n81), .A2(n7), .ZN(addr_x[0]) );
  NOR2_X1 U62 ( .A1(n13), .A2(n7), .ZN(\addr_a[0][0] ) );
  NAND2_X1 U63 ( .A1(n68), .A2(n86), .ZN(n48) );
  INV_X1 U64 ( .A(n84), .ZN(n22) );
  OR2_X1 U65 ( .A1(n28), .A2(n100), .ZN(n72) );
  NAND2_X1 U66 ( .A1(n73), .A2(n74), .ZN(n71) );
  OR2_X1 U67 ( .A1(n74), .A2(n28), .ZN(n95) );
  NAND2_X1 U68 ( .A1(n79), .A2(n96), .ZN(n80) );
  NOR2_X1 U69 ( .A1(n9), .A2(n75), .ZN(addr_y[1]) );
  INV_X1 U70 ( .A(n80), .ZN(n9) );
  INV_X1 U71 ( .A(n73), .ZN(n28) );
  OR2_X1 U72 ( .A1(counter2[0]), .A2(counter2[2]), .ZN(n39) );
  NAND2_X1 U73 ( .A1(n97), .A2(n23), .ZN(n38) );
  NAND3_X1 U74 ( .A1(n24), .A2(n23), .A3(state[0]), .ZN(n76) );
  OR2_X1 U75 ( .A1(n79), .A2(counter2[2]), .ZN(n1) );
  AOI221_X1 U76 ( .B1(n42), .B2(n84), .C1(n21), .C2(counter[3]), .A(done), 
        .ZN(n100) );
  NAND2_X1 U77 ( .A1(n21), .A2(n26), .ZN(n43) );
  NOR3_X1 U78 ( .A1(state[1]), .A2(state[2]), .A3(state[0]), .ZN(n84) );
  NOR2_X1 U79 ( .A1(counter[2]), .A2(counter[3]), .ZN(n91) );
  NOR2_X1 U80 ( .A1(n31), .A2(N244), .ZN(n64) );
  NOR2_X1 U81 ( .A1(n6), .A2(counter[3]), .ZN(n86) );
  NOR2_X1 U82 ( .A1(N244), .A2(counter[1]), .ZN(n69) );
  NOR2_X1 U83 ( .A1(n31), .A2(counter[0]), .ZN(n68) );
  OAI22_X1 U84 ( .A1(n70), .A2(n26), .B1(n47), .B2(n71), .ZN(n103) );
  AOI21_X1 U85 ( .B1(n10), .B2(n6), .A(n65), .ZN(n70) );
  NOR2_X1 U86 ( .A1(n24), .A2(state[0]), .ZN(n97) );
  NOR2_X1 U87 ( .A1(N248), .A2(N247), .ZN(n55) );
  INV_X1 U88 ( .A(n5), .ZN(N247) );
  INV_X1 U89 ( .A(n2), .ZN(N245) );
  NOR2_X1 U90 ( .A1(n42), .A2(n22), .ZN(wr_en_x) );
  OR2_X1 U91 ( .A1(counter2[1]), .A2(counter2[0]), .ZN(n79) );
  OAI21_X1 U92 ( .B1(n8), .B2(n6), .A(n63), .ZN(n101) );
  INV_X1 U93 ( .A(n65), .ZN(n8) );
  NOR3_X1 U94 ( .A1(n76), .A2(n61), .A3(n40), .ZN(wr_en_a[1]) );
  NOR4_X1 U95 ( .A1(N245), .A2(n1), .A3(counter[0]), .A4(n58), .ZN(n61) );
  NOR3_X1 U96 ( .A1(n76), .A2(n62), .A3(n42), .ZN(wr_en_a[0]) );
  NOR4_X1 U97 ( .A1(N245), .A2(N244), .A3(n1), .A4(n58), .ZN(n62) );
  NOR3_X1 U98 ( .A1(n59), .A2(n60), .A3(n76), .ZN(wr_en_a[2]) );
  NOR4_X1 U99 ( .A1(N244), .A2(n1), .A3(n2), .A4(n58), .ZN(n60) );
  NOR3_X1 U100 ( .A1(n56), .A2(n57), .A3(n76), .ZN(wr_en_a[3]) );
  NOR4_X1 U101 ( .A1(n1), .A2(counter[0]), .A3(n2), .A4(n58), .ZN(n57) );
  NOR3_X1 U102 ( .A1(n53), .A2(n54), .A3(n76), .ZN(wr_en_a[4]) );
  NOR4_X1 U103 ( .A1(N245), .A2(N244), .A3(n1), .A4(n46), .ZN(n54) );
  NOR3_X1 U104 ( .A1(n51), .A2(n52), .A3(n76), .ZN(wr_en_a[5]) );
  NOR4_X1 U105 ( .A1(N245), .A2(n1), .A3(n46), .A4(counter[0]), .ZN(n52) );
  NOR3_X1 U106 ( .A1(n48), .A2(n49), .A3(n76), .ZN(wr_en_a[6]) );
  NOR4_X1 U107 ( .A1(N244), .A2(n1), .A3(n46), .A4(n2), .ZN(n49) );
  NOR2_X1 U108 ( .A1(n43), .A2(n44), .ZN(wr_en_a[7]) );
  NOR4_X1 U109 ( .A1(n1), .A2(n46), .A3(counter[0]), .A4(n2), .ZN(n44) );
  NAND4_X1 U110 ( .A1(n75), .A2(n76), .A3(n22), .A4(n23), .ZN(clear_acc) );
  OAI221_X1 U111 ( .B1(n38), .B2(n72), .C1(reset), .C2(n29), .A(n99), .ZN(N128) );
  OAI221_X1 U112 ( .B1(n97), .B2(n72), .C1(n28), .C2(n23), .A(n27), .ZN(N130)
         );
  OAI22_X1 U113 ( .A1(N244), .A2(n66), .B1(counter[0]), .B2(n71), .ZN(n104) );
  OAI22_X1 U114 ( .A1(n12), .A2(n95), .B1(n96), .B2(n95), .ZN(N138) );
  NOR2_X1 U115 ( .A1(n96), .A2(n12), .ZN(n74) );
  NAND2_X1 U116 ( .A1(counter2[0]), .A2(counter2[1]), .ZN(n96) );
  OAI21_X1 U117 ( .B1(n31), .B2(n66), .A(n67), .ZN(n102) );
  OAI21_X1 U118 ( .B1(n68), .B2(n69), .A(n10), .ZN(n67) );
  OAI21_X1 U119 ( .B1(n24), .B2(n28), .A(n98), .ZN(N129) );
  NAND4_X1 U120 ( .A1(start), .A2(n29), .A3(n30), .A4(n27), .ZN(n98) );
  INV_X1 U121 ( .A(loadVector), .ZN(n30) );
  NOR2_X1 U122 ( .A1(counter2[0]), .A2(n95), .ZN(N136) );
  AOI21_X1 U123 ( .B1(n78), .B2(n1), .A(n75), .ZN(addr_y[2]) );
  NAND2_X1 U124 ( .A1(counter2[2]), .A2(n79), .ZN(n78) );
  NOR2_X1 U125 ( .A1(counter2[0]), .A2(n75), .ZN(addr_y[0]) );
  INV_X1 U126 ( .A(reset), .ZN(n27) );
  INV_X1 U127 ( .A(loadMatrix), .ZN(n29) );
  NOR2_X1 U128 ( .A1(counter[1]), .A2(counter[0]), .ZN(n3) );
  AOI21_X1 U129 ( .B1(counter[0]), .B2(counter[1]), .A(n3), .ZN(n2) );
  NAND2_X1 U130 ( .A1(n3), .A2(n6), .ZN(n4) );
  OAI21_X1 U131 ( .B1(n3), .B2(n6), .A(n4), .ZN(N246) );
  NOR2_X1 U132 ( .A1(n4), .A2(counter[3]), .ZN(N248) );
  AOI21_X1 U133 ( .B1(n4), .B2(counter[3]), .A(N248), .ZN(n5) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE4_8 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N13, N14, N15, N16, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N28, N29, N30, N31, N32, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[19]  ( .D(N13), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[17]  ( .D(N15), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N19), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N20), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N21), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N23), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N25), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N29), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N30), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N31), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N32), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n355), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n354), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n353), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n352), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n351), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n350), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n349), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n348), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n347), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n346), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n345), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n344), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n343), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n342), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n341), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n340), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n339), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n338), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n337), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n336), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n335), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n334), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n333), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n332), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n331), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n330), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n329), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n328), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n327), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n326), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n325), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n324), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n323), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n322), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n321), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n320), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n319), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n318), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n317), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n316), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n315), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n314), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n313), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n312), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n311), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n310), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n309), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n308), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n307), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n306), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n305), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n304), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n303), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n302), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n301), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n300), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n299), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n298), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n297), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n296), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n295), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n294), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n293), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n292), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n291), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n290), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n289), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n288), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n287), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n286), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n285), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n284), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n283), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n282), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n281), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n280), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n279), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n278), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n277), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n276), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n275), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n274), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n273), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n272), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n271), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n270), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n269), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n268), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n267), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n266), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n265), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n264), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n263), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n262), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n261), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n260), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n259), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n258), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n257), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n256), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n255), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n254), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n253), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n252), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n251), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n250), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n249), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n248), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n247), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n246), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n245), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n244), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n243), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n242), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n241), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n240), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n239), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n238), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n237), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n236), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n235), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n234), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n233), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n232), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n231), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n230), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n229), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n228), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n227), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n226), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n225), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n224), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n223), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n222), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n221), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n220), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n219), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n218), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n217), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n216), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n215), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n214), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n213), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n212), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n211), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n210), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n209), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n208), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n207), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n206), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n205), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n204), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n203), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n202), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n201), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n200), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n199), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n198), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n197), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n196), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U350 ( .A1(n466), .A2(n467), .A3(n46), .ZN(n25) );
  NAND3_X1 U351 ( .A1(n46), .A2(n467), .A3(N10), .ZN(n47) );
  NAND3_X1 U352 ( .A1(n46), .A2(n466), .A3(N11), .ZN(n68) );
  NAND3_X1 U353 ( .A1(N10), .A2(n46), .A3(N11), .ZN(n89) );
  NAND3_X1 U354 ( .A1(n466), .A2(n467), .A3(n132), .ZN(n111) );
  NAND3_X1 U355 ( .A1(N10), .A2(n467), .A3(n132), .ZN(n133) );
  NAND3_X1 U356 ( .A1(N11), .A2(n466), .A3(n132), .ZN(n154) );
  NAND3_X1 U357 ( .A1(N11), .A2(N10), .A3(n132), .ZN(n175) );
  SDFF_X1 \data_out_reg[5]  ( .D(n364), .SI(n367), .SE(n468), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n424), .SI(n427), .SE(n468), .CK(clk), .Q(
        data_out[15]) );
  BUF_X1 U3 ( .A(n25), .Z(n465) );
  BUF_X1 U4 ( .A(n68), .Z(n463) );
  BUF_X1 U5 ( .A(n133), .Z(n460) );
  BUF_X1 U6 ( .A(n453), .Z(n452) );
  BUF_X1 U7 ( .A(N10), .Z(n455) );
  BUF_X1 U8 ( .A(N10), .Z(n456) );
  BUF_X1 U9 ( .A(N10), .Z(n457) );
  BUF_X1 U10 ( .A(N10), .Z(n454) );
  BUF_X1 U11 ( .A(N11), .Z(n453) );
  BUF_X1 U12 ( .A(n89), .Z(n462) );
  BUF_X1 U13 ( .A(n47), .Z(n464) );
  BUF_X1 U14 ( .A(n175), .Z(n458) );
  BUF_X1 U15 ( .A(n111), .Z(n461) );
  BUF_X1 U16 ( .A(n154), .Z(n459) );
  NOR2_X1 U17 ( .A1(n110), .A2(N12), .ZN(n46) );
  NOR2_X1 U18 ( .A1(n468), .A2(n110), .ZN(n132) );
  INV_X1 U19 ( .A(N12), .ZN(n468) );
  INV_X1 U20 ( .A(N11), .ZN(n467) );
  INV_X1 U21 ( .A(N10), .ZN(n466) );
  OAI21_X1 U22 ( .B1(n477), .B2(n47), .A(n60), .ZN(n228) );
  NAND2_X1 U23 ( .A1(\mem[1][12] ), .A2(n47), .ZN(n60) );
  OAI21_X1 U24 ( .B1(n476), .B2(n47), .A(n61), .ZN(n229) );
  NAND2_X1 U25 ( .A1(\mem[1][13] ), .A2(n47), .ZN(n61) );
  OAI21_X1 U26 ( .B1(n475), .B2(n464), .A(n62), .ZN(n230) );
  NAND2_X1 U27 ( .A1(\mem[1][14] ), .A2(n47), .ZN(n62) );
  OAI21_X1 U28 ( .B1(n474), .B2(n464), .A(n63), .ZN(n231) );
  NAND2_X1 U29 ( .A1(\mem[1][15] ), .A2(n47), .ZN(n63) );
  OAI21_X1 U30 ( .B1(n473), .B2(n47), .A(n64), .ZN(n232) );
  NAND2_X1 U31 ( .A1(\mem[1][16] ), .A2(n47), .ZN(n64) );
  OAI21_X1 U32 ( .B1(n472), .B2(n47), .A(n65), .ZN(n233) );
  NAND2_X1 U33 ( .A1(\mem[1][17] ), .A2(n47), .ZN(n65) );
  OAI21_X1 U34 ( .B1(n471), .B2(n47), .A(n66), .ZN(n234) );
  NAND2_X1 U35 ( .A1(\mem[1][18] ), .A2(n47), .ZN(n66) );
  OAI21_X1 U36 ( .B1(n470), .B2(n47), .A(n67), .ZN(n235) );
  NAND2_X1 U37 ( .A1(\mem[1][19] ), .A2(n464), .ZN(n67) );
  OAI21_X1 U38 ( .B1(n477), .B2(n68), .A(n81), .ZN(n248) );
  NAND2_X1 U39 ( .A1(\mem[2][12] ), .A2(n68), .ZN(n81) );
  OAI21_X1 U40 ( .B1(n476), .B2(n68), .A(n82), .ZN(n249) );
  NAND2_X1 U41 ( .A1(\mem[2][13] ), .A2(n68), .ZN(n82) );
  OAI21_X1 U42 ( .B1(n475), .B2(n463), .A(n83), .ZN(n250) );
  NAND2_X1 U43 ( .A1(\mem[2][14] ), .A2(n68), .ZN(n83) );
  OAI21_X1 U44 ( .B1(n474), .B2(n463), .A(n84), .ZN(n251) );
  NAND2_X1 U45 ( .A1(\mem[2][15] ), .A2(n68), .ZN(n84) );
  OAI21_X1 U46 ( .B1(n473), .B2(n463), .A(n85), .ZN(n252) );
  NAND2_X1 U47 ( .A1(\mem[2][16] ), .A2(n68), .ZN(n85) );
  OAI21_X1 U48 ( .B1(n472), .B2(n463), .A(n86), .ZN(n253) );
  NAND2_X1 U49 ( .A1(\mem[2][17] ), .A2(n68), .ZN(n86) );
  OAI21_X1 U50 ( .B1(n471), .B2(n463), .A(n87), .ZN(n254) );
  NAND2_X1 U51 ( .A1(\mem[2][18] ), .A2(n68), .ZN(n87) );
  OAI21_X1 U52 ( .B1(n470), .B2(n68), .A(n88), .ZN(n255) );
  NAND2_X1 U53 ( .A1(\mem[2][19] ), .A2(n68), .ZN(n88) );
  OAI21_X1 U54 ( .B1(n477), .B2(n89), .A(n102), .ZN(n268) );
  NAND2_X1 U55 ( .A1(\mem[3][12] ), .A2(n89), .ZN(n102) );
  OAI21_X1 U56 ( .B1(n476), .B2(n89), .A(n103), .ZN(n269) );
  NAND2_X1 U57 ( .A1(\mem[3][13] ), .A2(n89), .ZN(n103) );
  OAI21_X1 U58 ( .B1(n475), .B2(n462), .A(n104), .ZN(n270) );
  NAND2_X1 U59 ( .A1(\mem[3][14] ), .A2(n89), .ZN(n104) );
  OAI21_X1 U60 ( .B1(n474), .B2(n462), .A(n105), .ZN(n271) );
  NAND2_X1 U61 ( .A1(\mem[3][15] ), .A2(n89), .ZN(n105) );
  OAI21_X1 U62 ( .B1(n473), .B2(n89), .A(n106), .ZN(n272) );
  NAND2_X1 U63 ( .A1(\mem[3][16] ), .A2(n89), .ZN(n106) );
  OAI21_X1 U64 ( .B1(n472), .B2(n89), .A(n107), .ZN(n273) );
  NAND2_X1 U65 ( .A1(\mem[3][17] ), .A2(n89), .ZN(n107) );
  OAI21_X1 U66 ( .B1(n471), .B2(n89), .A(n108), .ZN(n274) );
  NAND2_X1 U67 ( .A1(\mem[3][18] ), .A2(n89), .ZN(n108) );
  OAI21_X1 U68 ( .B1(n470), .B2(n89), .A(n109), .ZN(n275) );
  NAND2_X1 U69 ( .A1(\mem[3][19] ), .A2(n462), .ZN(n109) );
  OAI21_X1 U70 ( .B1(n489), .B2(n111), .A(n112), .ZN(n276) );
  NAND2_X1 U71 ( .A1(\mem[4][0] ), .A2(n461), .ZN(n112) );
  OAI21_X1 U72 ( .B1(n488), .B2(n111), .A(n113), .ZN(n277) );
  NAND2_X1 U73 ( .A1(\mem[4][1] ), .A2(n461), .ZN(n113) );
  OAI21_X1 U74 ( .B1(n487), .B2(n111), .A(n114), .ZN(n278) );
  NAND2_X1 U75 ( .A1(\mem[4][2] ), .A2(n461), .ZN(n114) );
  OAI21_X1 U76 ( .B1(n486), .B2(n111), .A(n115), .ZN(n279) );
  NAND2_X1 U77 ( .A1(\mem[4][3] ), .A2(n461), .ZN(n115) );
  OAI21_X1 U78 ( .B1(n485), .B2(n461), .A(n116), .ZN(n280) );
  NAND2_X1 U79 ( .A1(\mem[4][4] ), .A2(n461), .ZN(n116) );
  OAI21_X1 U80 ( .B1(n484), .B2(n111), .A(n117), .ZN(n281) );
  NAND2_X1 U81 ( .A1(\mem[4][5] ), .A2(n461), .ZN(n117) );
  OAI21_X1 U82 ( .B1(n483), .B2(n111), .A(n118), .ZN(n282) );
  NAND2_X1 U83 ( .A1(\mem[4][6] ), .A2(n461), .ZN(n118) );
  OAI21_X1 U84 ( .B1(n482), .B2(n111), .A(n119), .ZN(n283) );
  NAND2_X1 U85 ( .A1(\mem[4][7] ), .A2(n461), .ZN(n119) );
  OAI21_X1 U86 ( .B1(n481), .B2(n111), .A(n120), .ZN(n284) );
  NAND2_X1 U87 ( .A1(\mem[4][8] ), .A2(n461), .ZN(n120) );
  OAI21_X1 U88 ( .B1(n480), .B2(n111), .A(n121), .ZN(n285) );
  NAND2_X1 U89 ( .A1(\mem[4][9] ), .A2(n461), .ZN(n121) );
  OAI21_X1 U90 ( .B1(n479), .B2(n111), .A(n122), .ZN(n286) );
  NAND2_X1 U91 ( .A1(\mem[4][10] ), .A2(n461), .ZN(n122) );
  OAI21_X1 U92 ( .B1(n478), .B2(n111), .A(n123), .ZN(n287) );
  NAND2_X1 U93 ( .A1(\mem[4][11] ), .A2(n461), .ZN(n123) );
  OAI21_X1 U94 ( .B1(n477), .B2(n111), .A(n124), .ZN(n288) );
  NAND2_X1 U95 ( .A1(\mem[4][12] ), .A2(n111), .ZN(n124) );
  OAI21_X1 U96 ( .B1(n476), .B2(n461), .A(n125), .ZN(n289) );
  NAND2_X1 U97 ( .A1(\mem[4][13] ), .A2(n111), .ZN(n125) );
  OAI21_X1 U98 ( .B1(n475), .B2(n461), .A(n126), .ZN(n290) );
  NAND2_X1 U99 ( .A1(\mem[4][14] ), .A2(n111), .ZN(n126) );
  OAI21_X1 U100 ( .B1(n474), .B2(n111), .A(n127), .ZN(n291) );
  NAND2_X1 U101 ( .A1(\mem[4][15] ), .A2(n111), .ZN(n127) );
  OAI21_X1 U102 ( .B1(n473), .B2(n111), .A(n128), .ZN(n292) );
  NAND2_X1 U103 ( .A1(\mem[4][16] ), .A2(n111), .ZN(n128) );
  OAI21_X1 U104 ( .B1(n472), .B2(n111), .A(n129), .ZN(n293) );
  NAND2_X1 U105 ( .A1(\mem[4][17] ), .A2(n111), .ZN(n129) );
  OAI21_X1 U106 ( .B1(n471), .B2(n111), .A(n130), .ZN(n294) );
  NAND2_X1 U107 ( .A1(\mem[4][18] ), .A2(n111), .ZN(n130) );
  OAI21_X1 U108 ( .B1(n470), .B2(n111), .A(n131), .ZN(n295) );
  NAND2_X1 U109 ( .A1(\mem[4][19] ), .A2(n461), .ZN(n131) );
  OAI21_X1 U110 ( .B1(n489), .B2(n133), .A(n134), .ZN(n296) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n133), .ZN(n134) );
  OAI21_X1 U112 ( .B1(n488), .B2(n460), .A(n135), .ZN(n297) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n133), .ZN(n135) );
  OAI21_X1 U114 ( .B1(n487), .B2(n460), .A(n136), .ZN(n298) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n133), .ZN(n136) );
  OAI21_X1 U116 ( .B1(n486), .B2(n460), .A(n137), .ZN(n299) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n133), .ZN(n137) );
  OAI21_X1 U118 ( .B1(n485), .B2(n460), .A(n138), .ZN(n300) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n133), .ZN(n138) );
  OAI21_X1 U120 ( .B1(n484), .B2(n460), .A(n139), .ZN(n301) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n133), .ZN(n139) );
  OAI21_X1 U122 ( .B1(n483), .B2(n460), .A(n140), .ZN(n302) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n133), .ZN(n140) );
  OAI21_X1 U124 ( .B1(n482), .B2(n460), .A(n141), .ZN(n303) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n133), .ZN(n141) );
  OAI21_X1 U126 ( .B1(n481), .B2(n460), .A(n142), .ZN(n304) );
  NAND2_X1 U127 ( .A1(\mem[5][8] ), .A2(n133), .ZN(n142) );
  OAI21_X1 U128 ( .B1(n480), .B2(n133), .A(n143), .ZN(n305) );
  NAND2_X1 U129 ( .A1(\mem[5][9] ), .A2(n133), .ZN(n143) );
  OAI21_X1 U130 ( .B1(n479), .B2(n460), .A(n144), .ZN(n306) );
  NAND2_X1 U131 ( .A1(\mem[5][10] ), .A2(n133), .ZN(n144) );
  OAI21_X1 U132 ( .B1(n478), .B2(n460), .A(n145), .ZN(n307) );
  NAND2_X1 U133 ( .A1(\mem[5][11] ), .A2(n133), .ZN(n145) );
  OAI21_X1 U134 ( .B1(n477), .B2(n133), .A(n146), .ZN(n308) );
  NAND2_X1 U135 ( .A1(\mem[5][12] ), .A2(n133), .ZN(n146) );
  OAI21_X1 U136 ( .B1(n476), .B2(n460), .A(n147), .ZN(n309) );
  NAND2_X1 U137 ( .A1(\mem[5][13] ), .A2(n133), .ZN(n147) );
  OAI21_X1 U138 ( .B1(n475), .B2(n133), .A(n148), .ZN(n310) );
  NAND2_X1 U139 ( .A1(\mem[5][14] ), .A2(n133), .ZN(n148) );
  OAI21_X1 U140 ( .B1(n474), .B2(n460), .A(n149), .ZN(n311) );
  NAND2_X1 U141 ( .A1(\mem[5][15] ), .A2(n133), .ZN(n149) );
  OAI21_X1 U142 ( .B1(n473), .B2(n460), .A(n150), .ZN(n312) );
  NAND2_X1 U143 ( .A1(\mem[5][16] ), .A2(n133), .ZN(n150) );
  OAI21_X1 U144 ( .B1(n472), .B2(n460), .A(n151), .ZN(n313) );
  NAND2_X1 U145 ( .A1(\mem[5][17] ), .A2(n133), .ZN(n151) );
  OAI21_X1 U146 ( .B1(n471), .B2(n460), .A(n152), .ZN(n314) );
  NAND2_X1 U147 ( .A1(\mem[5][18] ), .A2(n133), .ZN(n152) );
  OAI21_X1 U148 ( .B1(n470), .B2(n460), .A(n153), .ZN(n315) );
  NAND2_X1 U149 ( .A1(\mem[5][19] ), .A2(n133), .ZN(n153) );
  OAI21_X1 U150 ( .B1(n489), .B2(n154), .A(n155), .ZN(n316) );
  NAND2_X1 U151 ( .A1(\mem[6][0] ), .A2(n459), .ZN(n155) );
  OAI21_X1 U152 ( .B1(n488), .B2(n154), .A(n156), .ZN(n317) );
  NAND2_X1 U153 ( .A1(\mem[6][1] ), .A2(n459), .ZN(n156) );
  OAI21_X1 U154 ( .B1(n487), .B2(n154), .A(n157), .ZN(n318) );
  NAND2_X1 U155 ( .A1(\mem[6][2] ), .A2(n459), .ZN(n157) );
  OAI21_X1 U156 ( .B1(n486), .B2(n154), .A(n158), .ZN(n319) );
  NAND2_X1 U157 ( .A1(\mem[6][3] ), .A2(n459), .ZN(n158) );
  OAI21_X1 U158 ( .B1(n485), .B2(n459), .A(n159), .ZN(n320) );
  NAND2_X1 U159 ( .A1(\mem[6][4] ), .A2(n459), .ZN(n159) );
  OAI21_X1 U160 ( .B1(n484), .B2(n154), .A(n160), .ZN(n321) );
  NAND2_X1 U161 ( .A1(\mem[6][5] ), .A2(n459), .ZN(n160) );
  OAI21_X1 U162 ( .B1(n483), .B2(n154), .A(n161), .ZN(n322) );
  NAND2_X1 U163 ( .A1(\mem[6][6] ), .A2(n459), .ZN(n161) );
  OAI21_X1 U164 ( .B1(n482), .B2(n154), .A(n162), .ZN(n323) );
  NAND2_X1 U165 ( .A1(\mem[6][7] ), .A2(n459), .ZN(n162) );
  OAI21_X1 U166 ( .B1(n481), .B2(n154), .A(n163), .ZN(n324) );
  NAND2_X1 U167 ( .A1(\mem[6][8] ), .A2(n459), .ZN(n163) );
  OAI21_X1 U168 ( .B1(n480), .B2(n154), .A(n164), .ZN(n325) );
  NAND2_X1 U169 ( .A1(\mem[6][9] ), .A2(n459), .ZN(n164) );
  OAI21_X1 U170 ( .B1(n479), .B2(n154), .A(n165), .ZN(n326) );
  NAND2_X1 U171 ( .A1(\mem[6][10] ), .A2(n459), .ZN(n165) );
  OAI21_X1 U172 ( .B1(n478), .B2(n154), .A(n166), .ZN(n327) );
  NAND2_X1 U173 ( .A1(\mem[6][11] ), .A2(n459), .ZN(n166) );
  OAI21_X1 U174 ( .B1(n477), .B2(n154), .A(n167), .ZN(n328) );
  NAND2_X1 U175 ( .A1(\mem[6][12] ), .A2(n154), .ZN(n167) );
  OAI21_X1 U176 ( .B1(n476), .B2(n459), .A(n168), .ZN(n329) );
  NAND2_X1 U177 ( .A1(\mem[6][13] ), .A2(n154), .ZN(n168) );
  OAI21_X1 U178 ( .B1(n475), .B2(n459), .A(n169), .ZN(n330) );
  NAND2_X1 U179 ( .A1(\mem[6][14] ), .A2(n154), .ZN(n169) );
  OAI21_X1 U180 ( .B1(n474), .B2(n154), .A(n170), .ZN(n331) );
  NAND2_X1 U181 ( .A1(\mem[6][15] ), .A2(n154), .ZN(n170) );
  OAI21_X1 U182 ( .B1(n473), .B2(n154), .A(n171), .ZN(n332) );
  NAND2_X1 U183 ( .A1(\mem[6][16] ), .A2(n154), .ZN(n171) );
  OAI21_X1 U184 ( .B1(n472), .B2(n154), .A(n172), .ZN(n333) );
  NAND2_X1 U185 ( .A1(\mem[6][17] ), .A2(n154), .ZN(n172) );
  OAI21_X1 U186 ( .B1(n471), .B2(n154), .A(n173), .ZN(n334) );
  NAND2_X1 U187 ( .A1(\mem[6][18] ), .A2(n154), .ZN(n173) );
  OAI21_X1 U188 ( .B1(n470), .B2(n154), .A(n174), .ZN(n335) );
  NAND2_X1 U189 ( .A1(\mem[6][19] ), .A2(n459), .ZN(n174) );
  OAI21_X1 U190 ( .B1(n489), .B2(n175), .A(n176), .ZN(n336) );
  NAND2_X1 U191 ( .A1(\mem[7][0] ), .A2(n458), .ZN(n176) );
  OAI21_X1 U192 ( .B1(n488), .B2(n175), .A(n177), .ZN(n337) );
  NAND2_X1 U193 ( .A1(\mem[7][1] ), .A2(n458), .ZN(n177) );
  OAI21_X1 U194 ( .B1(n487), .B2(n175), .A(n178), .ZN(n338) );
  NAND2_X1 U195 ( .A1(\mem[7][2] ), .A2(n458), .ZN(n178) );
  OAI21_X1 U196 ( .B1(n486), .B2(n175), .A(n179), .ZN(n339) );
  NAND2_X1 U197 ( .A1(\mem[7][3] ), .A2(n458), .ZN(n179) );
  OAI21_X1 U198 ( .B1(n485), .B2(n458), .A(n180), .ZN(n340) );
  NAND2_X1 U199 ( .A1(\mem[7][4] ), .A2(n458), .ZN(n180) );
  OAI21_X1 U200 ( .B1(n484), .B2(n175), .A(n181), .ZN(n341) );
  NAND2_X1 U201 ( .A1(\mem[7][5] ), .A2(n458), .ZN(n181) );
  OAI21_X1 U202 ( .B1(n483), .B2(n175), .A(n182), .ZN(n342) );
  NAND2_X1 U203 ( .A1(\mem[7][6] ), .A2(n458), .ZN(n182) );
  OAI21_X1 U204 ( .B1(n482), .B2(n175), .A(n183), .ZN(n343) );
  NAND2_X1 U205 ( .A1(\mem[7][7] ), .A2(n458), .ZN(n183) );
  OAI21_X1 U206 ( .B1(n481), .B2(n175), .A(n184), .ZN(n344) );
  NAND2_X1 U207 ( .A1(\mem[7][8] ), .A2(n458), .ZN(n184) );
  OAI21_X1 U208 ( .B1(n480), .B2(n175), .A(n185), .ZN(n345) );
  NAND2_X1 U209 ( .A1(\mem[7][9] ), .A2(n458), .ZN(n185) );
  OAI21_X1 U210 ( .B1(n479), .B2(n175), .A(n186), .ZN(n346) );
  NAND2_X1 U211 ( .A1(\mem[7][10] ), .A2(n458), .ZN(n186) );
  OAI21_X1 U212 ( .B1(n478), .B2(n175), .A(n187), .ZN(n347) );
  NAND2_X1 U213 ( .A1(\mem[7][11] ), .A2(n458), .ZN(n187) );
  OAI21_X1 U214 ( .B1(n477), .B2(n175), .A(n188), .ZN(n348) );
  NAND2_X1 U215 ( .A1(\mem[7][12] ), .A2(n175), .ZN(n188) );
  OAI21_X1 U216 ( .B1(n476), .B2(n458), .A(n189), .ZN(n349) );
  NAND2_X1 U217 ( .A1(\mem[7][13] ), .A2(n175), .ZN(n189) );
  OAI21_X1 U218 ( .B1(n475), .B2(n458), .A(n190), .ZN(n350) );
  NAND2_X1 U219 ( .A1(\mem[7][14] ), .A2(n175), .ZN(n190) );
  OAI21_X1 U220 ( .B1(n474), .B2(n175), .A(n191), .ZN(n351) );
  NAND2_X1 U221 ( .A1(\mem[7][15] ), .A2(n175), .ZN(n191) );
  OAI21_X1 U222 ( .B1(n473), .B2(n175), .A(n192), .ZN(n352) );
  NAND2_X1 U223 ( .A1(\mem[7][16] ), .A2(n175), .ZN(n192) );
  OAI21_X1 U224 ( .B1(n472), .B2(n175), .A(n193), .ZN(n353) );
  NAND2_X1 U225 ( .A1(\mem[7][17] ), .A2(n175), .ZN(n193) );
  OAI21_X1 U226 ( .B1(n471), .B2(n175), .A(n194), .ZN(n354) );
  NAND2_X1 U227 ( .A1(\mem[7][18] ), .A2(n175), .ZN(n194) );
  OAI21_X1 U228 ( .B1(n470), .B2(n175), .A(n195), .ZN(n355) );
  NAND2_X1 U229 ( .A1(\mem[7][19] ), .A2(n458), .ZN(n195) );
  NAND2_X1 U230 ( .A1(wr_en), .A2(n469), .ZN(n110) );
  INV_X1 U231 ( .A(addr[3]), .ZN(n469) );
  OAI21_X1 U232 ( .B1(n25), .B2(n489), .A(n26), .ZN(n196) );
  NAND2_X1 U233 ( .A1(\mem[0][0] ), .A2(n25), .ZN(n26) );
  OAI21_X1 U234 ( .B1(n25), .B2(n488), .A(n27), .ZN(n197) );
  NAND2_X1 U235 ( .A1(\mem[0][1] ), .A2(n25), .ZN(n27) );
  OAI21_X1 U236 ( .B1(n25), .B2(n487), .A(n28), .ZN(n198) );
  NAND2_X1 U237 ( .A1(\mem[0][2] ), .A2(n465), .ZN(n28) );
  OAI21_X1 U238 ( .B1(n25), .B2(n486), .A(n29), .ZN(n199) );
  NAND2_X1 U239 ( .A1(\mem[0][3] ), .A2(n465), .ZN(n29) );
  OAI21_X1 U240 ( .B1(n25), .B2(n485), .A(n30), .ZN(n200) );
  NAND2_X1 U241 ( .A1(\mem[0][4] ), .A2(n465), .ZN(n30) );
  OAI21_X1 U242 ( .B1(n25), .B2(n484), .A(n31), .ZN(n201) );
  NAND2_X1 U243 ( .A1(\mem[0][5] ), .A2(n465), .ZN(n31) );
  OAI21_X1 U244 ( .B1(n25), .B2(n483), .A(n32), .ZN(n202) );
  NAND2_X1 U245 ( .A1(\mem[0][6] ), .A2(n465), .ZN(n32) );
  OAI21_X1 U246 ( .B1(n25), .B2(n482), .A(n33), .ZN(n203) );
  NAND2_X1 U247 ( .A1(\mem[0][7] ), .A2(n25), .ZN(n33) );
  OAI21_X1 U248 ( .B1(n25), .B2(n481), .A(n34), .ZN(n204) );
  NAND2_X1 U249 ( .A1(\mem[0][8] ), .A2(n25), .ZN(n34) );
  OAI21_X1 U250 ( .B1(n465), .B2(n480), .A(n35), .ZN(n205) );
  NAND2_X1 U251 ( .A1(\mem[0][9] ), .A2(n25), .ZN(n35) );
  OAI21_X1 U252 ( .B1(n25), .B2(n479), .A(n36), .ZN(n206) );
  NAND2_X1 U253 ( .A1(\mem[0][10] ), .A2(n25), .ZN(n36) );
  OAI21_X1 U254 ( .B1(n25), .B2(n478), .A(n37), .ZN(n207) );
  NAND2_X1 U255 ( .A1(\mem[0][11] ), .A2(n25), .ZN(n37) );
  OAI21_X1 U256 ( .B1(n489), .B2(n47), .A(n48), .ZN(n216) );
  NAND2_X1 U257 ( .A1(\mem[1][0] ), .A2(n464), .ZN(n48) );
  OAI21_X1 U258 ( .B1(n488), .B2(n47), .A(n49), .ZN(n217) );
  NAND2_X1 U259 ( .A1(\mem[1][1] ), .A2(n464), .ZN(n49) );
  OAI21_X1 U260 ( .B1(n487), .B2(n47), .A(n50), .ZN(n218) );
  NAND2_X1 U261 ( .A1(\mem[1][2] ), .A2(n464), .ZN(n50) );
  OAI21_X1 U262 ( .B1(n486), .B2(n47), .A(n51), .ZN(n219) );
  NAND2_X1 U263 ( .A1(\mem[1][3] ), .A2(n464), .ZN(n51) );
  OAI21_X1 U264 ( .B1(n485), .B2(n47), .A(n52), .ZN(n220) );
  NAND2_X1 U265 ( .A1(\mem[1][4] ), .A2(n464), .ZN(n52) );
  OAI21_X1 U266 ( .B1(n484), .B2(n47), .A(n53), .ZN(n221) );
  NAND2_X1 U267 ( .A1(\mem[1][5] ), .A2(n464), .ZN(n53) );
  OAI21_X1 U268 ( .B1(n483), .B2(n47), .A(n54), .ZN(n222) );
  NAND2_X1 U269 ( .A1(\mem[1][6] ), .A2(n464), .ZN(n54) );
  OAI21_X1 U270 ( .B1(n482), .B2(n47), .A(n55), .ZN(n223) );
  NAND2_X1 U271 ( .A1(\mem[1][7] ), .A2(n464), .ZN(n55) );
  OAI21_X1 U272 ( .B1(n481), .B2(n47), .A(n56), .ZN(n224) );
  NAND2_X1 U273 ( .A1(\mem[1][8] ), .A2(n464), .ZN(n56) );
  OAI21_X1 U274 ( .B1(n480), .B2(n464), .A(n57), .ZN(n225) );
  NAND2_X1 U275 ( .A1(\mem[1][9] ), .A2(n464), .ZN(n57) );
  OAI21_X1 U276 ( .B1(n479), .B2(n47), .A(n58), .ZN(n226) );
  NAND2_X1 U277 ( .A1(\mem[1][10] ), .A2(n464), .ZN(n58) );
  OAI21_X1 U278 ( .B1(n478), .B2(n47), .A(n59), .ZN(n227) );
  NAND2_X1 U279 ( .A1(\mem[1][11] ), .A2(n464), .ZN(n59) );
  OAI21_X1 U280 ( .B1(n489), .B2(n463), .A(n69), .ZN(n236) );
  NAND2_X1 U281 ( .A1(\mem[2][0] ), .A2(n68), .ZN(n69) );
  OAI21_X1 U282 ( .B1(n488), .B2(n463), .A(n70), .ZN(n237) );
  NAND2_X1 U283 ( .A1(\mem[2][1] ), .A2(n68), .ZN(n70) );
  OAI21_X1 U284 ( .B1(n487), .B2(n463), .A(n71), .ZN(n238) );
  NAND2_X1 U285 ( .A1(\mem[2][2] ), .A2(n68), .ZN(n71) );
  OAI21_X1 U286 ( .B1(n486), .B2(n463), .A(n72), .ZN(n239) );
  NAND2_X1 U287 ( .A1(\mem[2][3] ), .A2(n68), .ZN(n72) );
  OAI21_X1 U288 ( .B1(n485), .B2(n463), .A(n73), .ZN(n240) );
  NAND2_X1 U289 ( .A1(\mem[2][4] ), .A2(n68), .ZN(n73) );
  OAI21_X1 U290 ( .B1(n484), .B2(n463), .A(n74), .ZN(n241) );
  NAND2_X1 U291 ( .A1(\mem[2][5] ), .A2(n68), .ZN(n74) );
  OAI21_X1 U292 ( .B1(n483), .B2(n463), .A(n75), .ZN(n242) );
  NAND2_X1 U293 ( .A1(\mem[2][6] ), .A2(n68), .ZN(n75) );
  OAI21_X1 U294 ( .B1(n482), .B2(n463), .A(n76), .ZN(n243) );
  NAND2_X1 U295 ( .A1(\mem[2][7] ), .A2(n68), .ZN(n76) );
  OAI21_X1 U296 ( .B1(n481), .B2(n463), .A(n77), .ZN(n244) );
  NAND2_X1 U297 ( .A1(\mem[2][8] ), .A2(n68), .ZN(n77) );
  OAI21_X1 U298 ( .B1(n480), .B2(n68), .A(n78), .ZN(n245) );
  NAND2_X1 U299 ( .A1(\mem[2][9] ), .A2(n68), .ZN(n78) );
  OAI21_X1 U300 ( .B1(n479), .B2(n463), .A(n79), .ZN(n246) );
  NAND2_X1 U301 ( .A1(\mem[2][10] ), .A2(n68), .ZN(n79) );
  OAI21_X1 U302 ( .B1(n478), .B2(n463), .A(n80), .ZN(n247) );
  NAND2_X1 U303 ( .A1(\mem[2][11] ), .A2(n68), .ZN(n80) );
  OAI21_X1 U304 ( .B1(n489), .B2(n89), .A(n90), .ZN(n256) );
  NAND2_X1 U305 ( .A1(\mem[3][0] ), .A2(n462), .ZN(n90) );
  OAI21_X1 U306 ( .B1(n488), .B2(n89), .A(n91), .ZN(n257) );
  NAND2_X1 U307 ( .A1(\mem[3][1] ), .A2(n462), .ZN(n91) );
  OAI21_X1 U308 ( .B1(n487), .B2(n89), .A(n92), .ZN(n258) );
  NAND2_X1 U309 ( .A1(\mem[3][2] ), .A2(n462), .ZN(n92) );
  OAI21_X1 U310 ( .B1(n486), .B2(n89), .A(n93), .ZN(n259) );
  NAND2_X1 U311 ( .A1(\mem[3][3] ), .A2(n462), .ZN(n93) );
  OAI21_X1 U312 ( .B1(n485), .B2(n89), .A(n94), .ZN(n260) );
  NAND2_X1 U313 ( .A1(\mem[3][4] ), .A2(n462), .ZN(n94) );
  OAI21_X1 U314 ( .B1(n484), .B2(n89), .A(n95), .ZN(n261) );
  NAND2_X1 U315 ( .A1(\mem[3][5] ), .A2(n462), .ZN(n95) );
  OAI21_X1 U316 ( .B1(n483), .B2(n89), .A(n96), .ZN(n262) );
  NAND2_X1 U317 ( .A1(\mem[3][6] ), .A2(n462), .ZN(n96) );
  OAI21_X1 U318 ( .B1(n482), .B2(n89), .A(n97), .ZN(n263) );
  NAND2_X1 U319 ( .A1(\mem[3][7] ), .A2(n462), .ZN(n97) );
  OAI21_X1 U320 ( .B1(n481), .B2(n89), .A(n98), .ZN(n264) );
  NAND2_X1 U321 ( .A1(\mem[3][8] ), .A2(n462), .ZN(n98) );
  OAI21_X1 U322 ( .B1(n480), .B2(n462), .A(n99), .ZN(n265) );
  NAND2_X1 U323 ( .A1(\mem[3][9] ), .A2(n462), .ZN(n99) );
  OAI21_X1 U324 ( .B1(n479), .B2(n89), .A(n100), .ZN(n266) );
  NAND2_X1 U325 ( .A1(\mem[3][10] ), .A2(n462), .ZN(n100) );
  OAI21_X1 U326 ( .B1(n478), .B2(n89), .A(n101), .ZN(n267) );
  NAND2_X1 U327 ( .A1(\mem[3][11] ), .A2(n462), .ZN(n101) );
  OAI21_X1 U328 ( .B1(n465), .B2(n477), .A(n38), .ZN(n208) );
  NAND2_X1 U329 ( .A1(\mem[0][12] ), .A2(n465), .ZN(n38) );
  OAI21_X1 U330 ( .B1(n465), .B2(n476), .A(n39), .ZN(n209) );
  NAND2_X1 U331 ( .A1(\mem[0][13] ), .A2(n465), .ZN(n39) );
  OAI21_X1 U332 ( .B1(n465), .B2(n475), .A(n40), .ZN(n210) );
  NAND2_X1 U333 ( .A1(\mem[0][14] ), .A2(n465), .ZN(n40) );
  OAI21_X1 U334 ( .B1(n25), .B2(n474), .A(n41), .ZN(n211) );
  NAND2_X1 U335 ( .A1(\mem[0][15] ), .A2(n465), .ZN(n41) );
  OAI21_X1 U336 ( .B1(n25), .B2(n473), .A(n42), .ZN(n212) );
  NAND2_X1 U337 ( .A1(\mem[0][16] ), .A2(n465), .ZN(n42) );
  OAI21_X1 U338 ( .B1(n25), .B2(n472), .A(n43), .ZN(n213) );
  NAND2_X1 U339 ( .A1(\mem[0][17] ), .A2(n465), .ZN(n43) );
  OAI21_X1 U340 ( .B1(n25), .B2(n471), .A(n44), .ZN(n214) );
  NAND2_X1 U341 ( .A1(\mem[0][18] ), .A2(n465), .ZN(n44) );
  OAI21_X1 U342 ( .B1(n25), .B2(n470), .A(n45), .ZN(n215) );
  NAND2_X1 U343 ( .A1(\mem[0][19] ), .A2(n465), .ZN(n45) );
  INV_X1 U344 ( .A(data_in[0]), .ZN(n489) );
  INV_X1 U345 ( .A(data_in[1]), .ZN(n488) );
  INV_X1 U346 ( .A(data_in[2]), .ZN(n487) );
  INV_X1 U347 ( .A(data_in[3]), .ZN(n486) );
  INV_X1 U348 ( .A(data_in[4]), .ZN(n485) );
  INV_X1 U349 ( .A(data_in[5]), .ZN(n484) );
  INV_X1 U358 ( .A(data_in[6]), .ZN(n483) );
  INV_X1 U359 ( .A(data_in[7]), .ZN(n482) );
  INV_X1 U360 ( .A(data_in[8]), .ZN(n481) );
  INV_X1 U361 ( .A(data_in[9]), .ZN(n480) );
  INV_X1 U362 ( .A(data_in[10]), .ZN(n479) );
  INV_X1 U363 ( .A(data_in[11]), .ZN(n478) );
  INV_X1 U364 ( .A(data_in[12]), .ZN(n477) );
  INV_X1 U365 ( .A(data_in[13]), .ZN(n476) );
  INV_X1 U366 ( .A(data_in[14]), .ZN(n475) );
  INV_X1 U367 ( .A(data_in[15]), .ZN(n474) );
  INV_X1 U368 ( .A(data_in[16]), .ZN(n473) );
  INV_X1 U369 ( .A(data_in[17]), .ZN(n472) );
  INV_X1 U370 ( .A(data_in[18]), .ZN(n471) );
  INV_X1 U371 ( .A(data_in[19]), .ZN(n470) );
  MUX2_X1 U372 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n457), .Z(n1) );
  MUX2_X1 U373 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n457), .Z(n2) );
  MUX2_X1 U374 ( .A(n2), .B(n1), .S(n452), .Z(n3) );
  MUX2_X1 U375 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n454), .Z(n4) );
  MUX2_X1 U376 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n454), .Z(n5) );
  MUX2_X1 U377 ( .A(n5), .B(n4), .S(n452), .Z(n6) );
  MUX2_X1 U378 ( .A(n6), .B(n3), .S(N12), .Z(N32) );
  MUX2_X1 U379 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n455), .Z(n7) );
  MUX2_X1 U380 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n455), .Z(n8) );
  MUX2_X1 U381 ( .A(n8), .B(n7), .S(n452), .Z(n9) );
  MUX2_X1 U382 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n456), .Z(n10) );
  MUX2_X1 U383 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n456), .Z(n11) );
  MUX2_X1 U384 ( .A(n11), .B(n10), .S(n452), .Z(n12) );
  MUX2_X1 U385 ( .A(n12), .B(n9), .S(N12), .Z(N31) );
  MUX2_X1 U386 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n454), .Z(n13) );
  MUX2_X1 U387 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n454), .Z(n14) );
  MUX2_X1 U388 ( .A(n14), .B(n13), .S(n453), .Z(n15) );
  MUX2_X1 U389 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n454), .Z(n16) );
  MUX2_X1 U390 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n454), .Z(n17) );
  MUX2_X1 U391 ( .A(n17), .B(n16), .S(n453), .Z(n18) );
  MUX2_X1 U392 ( .A(n18), .B(n15), .S(N12), .Z(N30) );
  MUX2_X1 U393 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n454), .Z(n19) );
  MUX2_X1 U394 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n454), .Z(n20) );
  MUX2_X1 U395 ( .A(n20), .B(n19), .S(n453), .Z(n21) );
  MUX2_X1 U396 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n454), .Z(n22) );
  MUX2_X1 U397 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n454), .Z(n23) );
  MUX2_X1 U398 ( .A(n23), .B(n22), .S(n453), .Z(n24) );
  MUX2_X1 U399 ( .A(n24), .B(n21), .S(N12), .Z(N29) );
  MUX2_X1 U400 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n454), .Z(n356) );
  MUX2_X1 U401 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n454), .Z(n357) );
  MUX2_X1 U402 ( .A(n357), .B(n356), .S(n453), .Z(n358) );
  MUX2_X1 U403 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n454), .Z(n359) );
  MUX2_X1 U404 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n454), .Z(n360) );
  MUX2_X1 U405 ( .A(n360), .B(n359), .S(n453), .Z(n361) );
  MUX2_X1 U406 ( .A(n361), .B(n358), .S(N12), .Z(N28) );
  MUX2_X1 U407 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n454), .Z(n362) );
  MUX2_X1 U408 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n455), .Z(n363) );
  MUX2_X1 U409 ( .A(n363), .B(n362), .S(n453), .Z(n364) );
  MUX2_X1 U410 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n457), .Z(n365) );
  MUX2_X1 U411 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n457), .Z(n366) );
  MUX2_X1 U412 ( .A(n366), .B(n365), .S(n453), .Z(n367) );
  MUX2_X1 U413 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n456), .Z(n368) );
  MUX2_X1 U414 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n456), .Z(n369) );
  MUX2_X1 U415 ( .A(n369), .B(n368), .S(n453), .Z(n370) );
  MUX2_X1 U416 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n454), .Z(n371) );
  MUX2_X1 U417 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n455), .Z(n372) );
  MUX2_X1 U418 ( .A(n372), .B(n371), .S(n453), .Z(n373) );
  MUX2_X1 U419 ( .A(n373), .B(n370), .S(N12), .Z(N26) );
  MUX2_X1 U420 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n457), .Z(n374) );
  MUX2_X1 U421 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n457), .Z(n375) );
  MUX2_X1 U422 ( .A(n375), .B(n374), .S(n453), .Z(n376) );
  MUX2_X1 U423 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n455), .Z(n377) );
  MUX2_X1 U424 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n456), .Z(n378) );
  MUX2_X1 U425 ( .A(n378), .B(n377), .S(n453), .Z(n379) );
  MUX2_X1 U426 ( .A(n379), .B(n376), .S(N12), .Z(N25) );
  MUX2_X1 U427 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n455), .Z(n380) );
  MUX2_X1 U428 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n454), .Z(n381) );
  MUX2_X1 U429 ( .A(n381), .B(n380), .S(n453), .Z(n382) );
  MUX2_X1 U430 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n455), .Z(n383) );
  MUX2_X1 U431 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n455), .Z(n384) );
  MUX2_X1 U432 ( .A(n384), .B(n383), .S(N11), .Z(n385) );
  MUX2_X1 U433 ( .A(n385), .B(n382), .S(N12), .Z(N24) );
  MUX2_X1 U434 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n454), .Z(n386) );
  MUX2_X1 U435 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n454), .Z(n387) );
  MUX2_X1 U436 ( .A(n387), .B(n386), .S(n453), .Z(n388) );
  MUX2_X1 U437 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n456), .Z(n389) );
  MUX2_X1 U438 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n456), .Z(n390) );
  MUX2_X1 U439 ( .A(n390), .B(n389), .S(N11), .Z(n391) );
  MUX2_X1 U440 ( .A(n391), .B(n388), .S(N12), .Z(N23) );
  MUX2_X1 U441 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n456), .Z(n392) );
  MUX2_X1 U442 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n454), .Z(n393) );
  MUX2_X1 U443 ( .A(n393), .B(n392), .S(n453), .Z(n394) );
  MUX2_X1 U444 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n457), .Z(n395) );
  MUX2_X1 U445 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n457), .Z(n396) );
  MUX2_X1 U446 ( .A(n396), .B(n395), .S(N11), .Z(n397) );
  MUX2_X1 U447 ( .A(n397), .B(n394), .S(N12), .Z(N22) );
  MUX2_X1 U448 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n455), .Z(n398) );
  MUX2_X1 U449 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n455), .Z(n399) );
  MUX2_X1 U450 ( .A(n399), .B(n398), .S(n453), .Z(n400) );
  MUX2_X1 U451 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n455), .Z(n401) );
  MUX2_X1 U452 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n455), .Z(n402) );
  MUX2_X1 U453 ( .A(n402), .B(n401), .S(N11), .Z(n403) );
  MUX2_X1 U454 ( .A(n403), .B(n400), .S(N12), .Z(N21) );
  MUX2_X1 U455 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n455), .Z(n404) );
  MUX2_X1 U456 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n455), .Z(n405) );
  MUX2_X1 U457 ( .A(n405), .B(n404), .S(n453), .Z(n406) );
  MUX2_X1 U458 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n455), .Z(n407) );
  MUX2_X1 U459 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n455), .Z(n408) );
  MUX2_X1 U460 ( .A(n408), .B(n407), .S(N11), .Z(n409) );
  MUX2_X1 U461 ( .A(n409), .B(n406), .S(N12), .Z(N20) );
  MUX2_X1 U462 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n455), .Z(n410) );
  MUX2_X1 U463 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n455), .Z(n411) );
  MUX2_X1 U464 ( .A(n411), .B(n410), .S(n453), .Z(n412) );
  MUX2_X1 U465 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n455), .Z(n413) );
  MUX2_X1 U466 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n455), .Z(n414) );
  MUX2_X1 U467 ( .A(n414), .B(n413), .S(N11), .Z(n415) );
  MUX2_X1 U468 ( .A(n415), .B(n412), .S(N12), .Z(N19) );
  MUX2_X1 U469 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n456), .Z(n416) );
  MUX2_X1 U470 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n456), .Z(n417) );
  MUX2_X1 U471 ( .A(n417), .B(n416), .S(n452), .Z(n418) );
  MUX2_X1 U472 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n456), .Z(n419) );
  MUX2_X1 U473 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n456), .Z(n420) );
  MUX2_X1 U474 ( .A(n420), .B(n419), .S(n452), .Z(n421) );
  MUX2_X1 U475 ( .A(n421), .B(n418), .S(N12), .Z(N18) );
  MUX2_X1 U476 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n456), .Z(n422) );
  MUX2_X1 U477 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n456), .Z(n423) );
  MUX2_X1 U478 ( .A(n423), .B(n422), .S(n453), .Z(n424) );
  MUX2_X1 U479 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n456), .Z(n425) );
  MUX2_X1 U480 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n456), .Z(n426) );
  MUX2_X1 U481 ( .A(n426), .B(n425), .S(n453), .Z(n427) );
  MUX2_X1 U482 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n456), .Z(n428) );
  MUX2_X1 U483 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n456), .Z(n429) );
  MUX2_X1 U484 ( .A(n429), .B(n428), .S(n452), .Z(n430) );
  MUX2_X1 U485 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n456), .Z(n431) );
  MUX2_X1 U486 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n456), .Z(n432) );
  MUX2_X1 U487 ( .A(n432), .B(n431), .S(n452), .Z(n433) );
  MUX2_X1 U488 ( .A(n433), .B(n430), .S(N12), .Z(N16) );
  MUX2_X1 U489 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n457), .Z(n434) );
  MUX2_X1 U490 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n457), .Z(n435) );
  MUX2_X1 U491 ( .A(n435), .B(n434), .S(n452), .Z(n436) );
  MUX2_X1 U492 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n457), .Z(n437) );
  MUX2_X1 U493 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n457), .Z(n438) );
  MUX2_X1 U494 ( .A(n438), .B(n437), .S(n452), .Z(n439) );
  MUX2_X1 U495 ( .A(n439), .B(n436), .S(N12), .Z(N15) );
  MUX2_X1 U496 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n457), .Z(n440) );
  MUX2_X1 U497 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n457), .Z(n441) );
  MUX2_X1 U498 ( .A(n441), .B(n440), .S(n452), .Z(n442) );
  MUX2_X1 U499 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n457), .Z(n443) );
  MUX2_X1 U500 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n457), .Z(n444) );
  MUX2_X1 U501 ( .A(n444), .B(n443), .S(n453), .Z(n445) );
  MUX2_X1 U502 ( .A(n445), .B(n442), .S(N12), .Z(N14) );
  MUX2_X1 U503 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n457), .Z(n446) );
  MUX2_X1 U504 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n457), .Z(n447) );
  MUX2_X1 U505 ( .A(n447), .B(n446), .S(n452), .Z(n448) );
  MUX2_X1 U506 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n457), .Z(n449) );
  MUX2_X1 U507 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n457), .Z(n450) );
  MUX2_X1 U508 ( .A(n450), .B(n449), .S(n453), .Z(n451) );
  MUX2_X1 U509 ( .A(n451), .B(n448), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE4_7 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N13, N14, N15, N16, N17, N18, N22, N24, N25, N26, N27,
         N28, N29, N30, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[19]  ( .D(N13), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[17]  ( .D(N15), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[15]  ( .D(N17), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N25), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N27), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N29), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N30), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N32), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n490), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n491), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n492), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n493), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n494), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n495), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n496), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n497), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n498), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n499), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n500), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n501), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n502), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n503), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n504), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n505), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n506), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n507), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n508), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n509), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n510), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n511), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n512), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n513), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n514), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n515), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n516), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n517), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n518), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n519), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n520), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n521), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n522), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n523), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n524), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n525), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n526), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n527), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n528), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n529), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n530), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n531), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n532), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n533), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n534), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n535), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n536), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n537), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n538), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n539), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n540), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n541), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n542), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n543), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n544), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n545), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n546), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n547), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n548), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n549), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n550), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n551), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n552), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n553), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n554), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n555), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n556), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n557), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n558), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n559), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n560), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n561), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n562), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n563), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n564), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n565), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n566), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n567), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n568), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n569), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n570), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n571), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n572), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n573), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n574), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n575), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n576), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n577), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n578), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n579), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n580), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n581), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n582), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n583), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n584), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n585), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n586), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n587), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n588), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n589), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n590), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n591), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n592), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n593), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n594), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n595), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n596), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n597), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n598), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n599), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n600), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n601), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n602), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n603), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n604), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n605), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n606), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n607), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n608), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n609), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n610), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n611), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n612), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n613), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n614), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n615), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n616), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n617), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n618), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n619), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n620), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n621), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n622), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n623), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n624), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n625), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n626), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n627), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n628), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n629), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n630), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n631), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n632), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n633), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n634), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n635), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n636), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n637), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n638), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n639), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n640), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n641), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n642), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n643), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n644), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n645), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n646), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n647), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n648), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n649), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U350 ( .A1(n466), .A2(n467), .A3(n799), .ZN(n820) );
  NAND3_X1 U351 ( .A1(n799), .A2(n467), .A3(N10), .ZN(n798) );
  NAND3_X1 U352 ( .A1(n799), .A2(n466), .A3(N11), .ZN(n777) );
  NAND3_X1 U353 ( .A1(N10), .A2(n799), .A3(N11), .ZN(n756) );
  NAND3_X1 U354 ( .A1(n466), .A2(n467), .A3(n713), .ZN(n734) );
  NAND3_X1 U355 ( .A1(N10), .A2(n467), .A3(n713), .ZN(n712) );
  NAND3_X1 U356 ( .A1(N11), .A2(n466), .A3(n713), .ZN(n691) );
  NAND3_X1 U357 ( .A1(N11), .A2(N10), .A3(n713), .ZN(n670) );
  SDFF_X1 \data_out_reg[13]  ( .D(n412), .SI(n415), .SE(n468), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n400), .SI(n403), .SE(n468), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[12]  ( .D(n406), .SI(n409), .SE(n468), .CK(clk), .Q(
        data_out[12]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n9), .SI(n12), .SE(n468), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n388), .SI(n391), .SE(n468), .CK(clk), .Q(
        data_out[9]) );
  BUF_X1 U3 ( .A(n777), .Z(n463) );
  BUF_X1 U4 ( .A(n712), .Z(n460) );
  BUF_X1 U5 ( .A(n670), .Z(n458) );
  BUF_X1 U6 ( .A(n453), .Z(n452) );
  BUF_X1 U7 ( .A(N10), .Z(n455) );
  BUF_X1 U8 ( .A(N10), .Z(n456) );
  BUF_X1 U9 ( .A(N10), .Z(n457) );
  BUF_X1 U10 ( .A(N10), .Z(n454) );
  BUF_X1 U11 ( .A(N11), .Z(n453) );
  BUF_X1 U12 ( .A(n820), .Z(n465) );
  BUF_X1 U13 ( .A(n756), .Z(n462) );
  BUF_X1 U14 ( .A(n798), .Z(n464) );
  BUF_X1 U15 ( .A(n734), .Z(n461) );
  BUF_X1 U16 ( .A(n691), .Z(n459) );
  NOR2_X1 U17 ( .A1(n735), .A2(N12), .ZN(n799) );
  NOR2_X1 U18 ( .A1(n468), .A2(n735), .ZN(n713) );
  INV_X1 U19 ( .A(N12), .ZN(n468) );
  INV_X1 U20 ( .A(N11), .ZN(n467) );
  INV_X1 U21 ( .A(N10), .ZN(n466) );
  OAI21_X1 U22 ( .B1(n477), .B2(n798), .A(n785), .ZN(n617) );
  NAND2_X1 U23 ( .A1(\mem[1][12] ), .A2(n798), .ZN(n785) );
  OAI21_X1 U24 ( .B1(n476), .B2(n798), .A(n784), .ZN(n616) );
  NAND2_X1 U25 ( .A1(\mem[1][13] ), .A2(n798), .ZN(n784) );
  OAI21_X1 U26 ( .B1(n475), .B2(n798), .A(n783), .ZN(n615) );
  NAND2_X1 U27 ( .A1(\mem[1][14] ), .A2(n798), .ZN(n783) );
  OAI21_X1 U28 ( .B1(n474), .B2(n464), .A(n782), .ZN(n614) );
  NAND2_X1 U29 ( .A1(\mem[1][15] ), .A2(n798), .ZN(n782) );
  OAI21_X1 U30 ( .B1(n473), .B2(n798), .A(n781), .ZN(n613) );
  NAND2_X1 U31 ( .A1(\mem[1][16] ), .A2(n464), .ZN(n781) );
  OAI21_X1 U32 ( .B1(n472), .B2(n798), .A(n780), .ZN(n612) );
  NAND2_X1 U33 ( .A1(\mem[1][17] ), .A2(n798), .ZN(n780) );
  OAI21_X1 U34 ( .B1(n471), .B2(n798), .A(n779), .ZN(n611) );
  NAND2_X1 U35 ( .A1(\mem[1][18] ), .A2(n798), .ZN(n779) );
  OAI21_X1 U36 ( .B1(n470), .B2(n798), .A(n778), .ZN(n610) );
  NAND2_X1 U37 ( .A1(\mem[1][19] ), .A2(n464), .ZN(n778) );
  OAI21_X1 U38 ( .B1(n477), .B2(n463), .A(n764), .ZN(n597) );
  NAND2_X1 U39 ( .A1(\mem[2][12] ), .A2(n463), .ZN(n764) );
  OAI21_X1 U40 ( .B1(n476), .B2(n463), .A(n763), .ZN(n596) );
  NAND2_X1 U41 ( .A1(\mem[2][13] ), .A2(n463), .ZN(n763) );
  OAI21_X1 U42 ( .B1(n475), .B2(n463), .A(n762), .ZN(n595) );
  NAND2_X1 U43 ( .A1(\mem[2][14] ), .A2(n463), .ZN(n762) );
  OAI21_X1 U44 ( .B1(n474), .B2(n777), .A(n761), .ZN(n594) );
  NAND2_X1 U45 ( .A1(\mem[2][15] ), .A2(n463), .ZN(n761) );
  OAI21_X1 U46 ( .B1(n473), .B2(n777), .A(n760), .ZN(n593) );
  NAND2_X1 U47 ( .A1(\mem[2][16] ), .A2(n463), .ZN(n760) );
  OAI21_X1 U48 ( .B1(n472), .B2(n777), .A(n759), .ZN(n592) );
  NAND2_X1 U49 ( .A1(\mem[2][17] ), .A2(n463), .ZN(n759) );
  OAI21_X1 U50 ( .B1(n471), .B2(n777), .A(n758), .ZN(n591) );
  NAND2_X1 U51 ( .A1(\mem[2][18] ), .A2(n463), .ZN(n758) );
  OAI21_X1 U52 ( .B1(n470), .B2(n777), .A(n757), .ZN(n590) );
  NAND2_X1 U53 ( .A1(\mem[2][19] ), .A2(n463), .ZN(n757) );
  OAI21_X1 U54 ( .B1(n477), .B2(n756), .A(n743), .ZN(n577) );
  NAND2_X1 U55 ( .A1(\mem[3][12] ), .A2(n756), .ZN(n743) );
  OAI21_X1 U56 ( .B1(n476), .B2(n756), .A(n742), .ZN(n576) );
  NAND2_X1 U57 ( .A1(\mem[3][13] ), .A2(n756), .ZN(n742) );
  OAI21_X1 U58 ( .B1(n475), .B2(n756), .A(n741), .ZN(n575) );
  NAND2_X1 U59 ( .A1(\mem[3][14] ), .A2(n756), .ZN(n741) );
  OAI21_X1 U60 ( .B1(n474), .B2(n462), .A(n740), .ZN(n574) );
  NAND2_X1 U61 ( .A1(\mem[3][15] ), .A2(n756), .ZN(n740) );
  OAI21_X1 U62 ( .B1(n473), .B2(n756), .A(n739), .ZN(n573) );
  NAND2_X1 U63 ( .A1(\mem[3][16] ), .A2(n462), .ZN(n739) );
  OAI21_X1 U64 ( .B1(n472), .B2(n756), .A(n738), .ZN(n572) );
  NAND2_X1 U65 ( .A1(\mem[3][17] ), .A2(n756), .ZN(n738) );
  OAI21_X1 U66 ( .B1(n471), .B2(n756), .A(n737), .ZN(n571) );
  NAND2_X1 U67 ( .A1(\mem[3][18] ), .A2(n756), .ZN(n737) );
  OAI21_X1 U68 ( .B1(n470), .B2(n756), .A(n736), .ZN(n570) );
  NAND2_X1 U69 ( .A1(\mem[3][19] ), .A2(n462), .ZN(n736) );
  OAI21_X1 U70 ( .B1(n489), .B2(n734), .A(n733), .ZN(n569) );
  NAND2_X1 U71 ( .A1(\mem[4][0] ), .A2(n461), .ZN(n733) );
  OAI21_X1 U72 ( .B1(n488), .B2(n734), .A(n732), .ZN(n568) );
  NAND2_X1 U73 ( .A1(\mem[4][1] ), .A2(n461), .ZN(n732) );
  OAI21_X1 U74 ( .B1(n487), .B2(n734), .A(n731), .ZN(n567) );
  NAND2_X1 U75 ( .A1(\mem[4][2] ), .A2(n461), .ZN(n731) );
  OAI21_X1 U76 ( .B1(n486), .B2(n734), .A(n730), .ZN(n566) );
  NAND2_X1 U77 ( .A1(\mem[4][3] ), .A2(n461), .ZN(n730) );
  OAI21_X1 U78 ( .B1(n485), .B2(n461), .A(n729), .ZN(n565) );
  NAND2_X1 U79 ( .A1(\mem[4][4] ), .A2(n461), .ZN(n729) );
  OAI21_X1 U80 ( .B1(n484), .B2(n734), .A(n728), .ZN(n564) );
  NAND2_X1 U81 ( .A1(\mem[4][5] ), .A2(n461), .ZN(n728) );
  OAI21_X1 U82 ( .B1(n483), .B2(n734), .A(n727), .ZN(n563) );
  NAND2_X1 U83 ( .A1(\mem[4][6] ), .A2(n461), .ZN(n727) );
  OAI21_X1 U84 ( .B1(n482), .B2(n734), .A(n726), .ZN(n562) );
  NAND2_X1 U85 ( .A1(\mem[4][7] ), .A2(n461), .ZN(n726) );
  OAI21_X1 U86 ( .B1(n481), .B2(n734), .A(n725), .ZN(n561) );
  NAND2_X1 U87 ( .A1(\mem[4][8] ), .A2(n461), .ZN(n725) );
  OAI21_X1 U88 ( .B1(n480), .B2(n734), .A(n724), .ZN(n560) );
  NAND2_X1 U89 ( .A1(\mem[4][9] ), .A2(n461), .ZN(n724) );
  OAI21_X1 U90 ( .B1(n479), .B2(n734), .A(n723), .ZN(n559) );
  NAND2_X1 U91 ( .A1(\mem[4][10] ), .A2(n461), .ZN(n723) );
  OAI21_X1 U92 ( .B1(n478), .B2(n734), .A(n722), .ZN(n558) );
  NAND2_X1 U93 ( .A1(\mem[4][11] ), .A2(n461), .ZN(n722) );
  OAI21_X1 U94 ( .B1(n477), .B2(n734), .A(n721), .ZN(n557) );
  NAND2_X1 U95 ( .A1(\mem[4][12] ), .A2(n734), .ZN(n721) );
  OAI21_X1 U96 ( .B1(n476), .B2(n461), .A(n720), .ZN(n556) );
  NAND2_X1 U97 ( .A1(\mem[4][13] ), .A2(n734), .ZN(n720) );
  OAI21_X1 U98 ( .B1(n475), .B2(n461), .A(n719), .ZN(n555) );
  NAND2_X1 U99 ( .A1(\mem[4][14] ), .A2(n734), .ZN(n719) );
  OAI21_X1 U100 ( .B1(n474), .B2(n734), .A(n718), .ZN(n554) );
  NAND2_X1 U101 ( .A1(\mem[4][15] ), .A2(n734), .ZN(n718) );
  OAI21_X1 U102 ( .B1(n473), .B2(n734), .A(n717), .ZN(n553) );
  NAND2_X1 U103 ( .A1(\mem[4][16] ), .A2(n734), .ZN(n717) );
  OAI21_X1 U104 ( .B1(n472), .B2(n734), .A(n716), .ZN(n552) );
  NAND2_X1 U105 ( .A1(\mem[4][17] ), .A2(n734), .ZN(n716) );
  OAI21_X1 U106 ( .B1(n471), .B2(n734), .A(n715), .ZN(n551) );
  NAND2_X1 U107 ( .A1(\mem[4][18] ), .A2(n734), .ZN(n715) );
  OAI21_X1 U108 ( .B1(n470), .B2(n734), .A(n714), .ZN(n550) );
  NAND2_X1 U109 ( .A1(\mem[4][19] ), .A2(n461), .ZN(n714) );
  OAI21_X1 U110 ( .B1(n489), .B2(n460), .A(n711), .ZN(n549) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n460), .ZN(n711) );
  OAI21_X1 U112 ( .B1(n488), .B2(n460), .A(n710), .ZN(n548) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n460), .ZN(n710) );
  OAI21_X1 U114 ( .B1(n487), .B2(n460), .A(n709), .ZN(n547) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n712), .ZN(n709) );
  OAI21_X1 U116 ( .B1(n486), .B2(n712), .A(n708), .ZN(n546) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n460), .ZN(n708) );
  OAI21_X1 U118 ( .B1(n485), .B2(n712), .A(n707), .ZN(n545) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n712), .ZN(n707) );
  OAI21_X1 U120 ( .B1(n484), .B2(n712), .A(n706), .ZN(n544) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n712), .ZN(n706) );
  OAI21_X1 U122 ( .B1(n483), .B2(n712), .A(n705), .ZN(n543) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n712), .ZN(n705) );
  OAI21_X1 U124 ( .B1(n482), .B2(n712), .A(n704), .ZN(n542) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n712), .ZN(n704) );
  OAI21_X1 U126 ( .B1(n481), .B2(n712), .A(n703), .ZN(n541) );
  NAND2_X1 U127 ( .A1(\mem[5][8] ), .A2(n712), .ZN(n703) );
  OAI21_X1 U128 ( .B1(n480), .B2(n460), .A(n702), .ZN(n540) );
  NAND2_X1 U129 ( .A1(\mem[5][9] ), .A2(n712), .ZN(n702) );
  OAI21_X1 U130 ( .B1(n479), .B2(n712), .A(n701), .ZN(n539) );
  NAND2_X1 U131 ( .A1(\mem[5][10] ), .A2(n712), .ZN(n701) );
  OAI21_X1 U132 ( .B1(n478), .B2(n712), .A(n700), .ZN(n538) );
  NAND2_X1 U133 ( .A1(\mem[5][11] ), .A2(n712), .ZN(n700) );
  OAI21_X1 U134 ( .B1(n477), .B2(n460), .A(n699), .ZN(n537) );
  NAND2_X1 U135 ( .A1(\mem[5][12] ), .A2(n460), .ZN(n699) );
  OAI21_X1 U136 ( .B1(n476), .B2(n460), .A(n698), .ZN(n536) );
  NAND2_X1 U137 ( .A1(\mem[5][13] ), .A2(n460), .ZN(n698) );
  OAI21_X1 U138 ( .B1(n475), .B2(n460), .A(n697), .ZN(n535) );
  NAND2_X1 U139 ( .A1(\mem[5][14] ), .A2(n460), .ZN(n697) );
  OAI21_X1 U140 ( .B1(n474), .B2(n712), .A(n696), .ZN(n534) );
  NAND2_X1 U141 ( .A1(\mem[5][15] ), .A2(n460), .ZN(n696) );
  OAI21_X1 U142 ( .B1(n473), .B2(n712), .A(n695), .ZN(n533) );
  NAND2_X1 U143 ( .A1(\mem[5][16] ), .A2(n460), .ZN(n695) );
  OAI21_X1 U144 ( .B1(n472), .B2(n712), .A(n694), .ZN(n532) );
  NAND2_X1 U145 ( .A1(\mem[5][17] ), .A2(n460), .ZN(n694) );
  OAI21_X1 U146 ( .B1(n471), .B2(n460), .A(n693), .ZN(n531) );
  NAND2_X1 U147 ( .A1(\mem[5][18] ), .A2(n460), .ZN(n693) );
  OAI21_X1 U148 ( .B1(n470), .B2(n460), .A(n692), .ZN(n530) );
  NAND2_X1 U149 ( .A1(\mem[5][19] ), .A2(n460), .ZN(n692) );
  OAI21_X1 U150 ( .B1(n489), .B2(n691), .A(n690), .ZN(n529) );
  NAND2_X1 U151 ( .A1(\mem[6][0] ), .A2(n459), .ZN(n690) );
  OAI21_X1 U152 ( .B1(n488), .B2(n691), .A(n689), .ZN(n528) );
  NAND2_X1 U153 ( .A1(\mem[6][1] ), .A2(n459), .ZN(n689) );
  OAI21_X1 U154 ( .B1(n487), .B2(n691), .A(n688), .ZN(n527) );
  NAND2_X1 U155 ( .A1(\mem[6][2] ), .A2(n459), .ZN(n688) );
  OAI21_X1 U156 ( .B1(n486), .B2(n691), .A(n687), .ZN(n526) );
  NAND2_X1 U157 ( .A1(\mem[6][3] ), .A2(n459), .ZN(n687) );
  OAI21_X1 U158 ( .B1(n485), .B2(n459), .A(n686), .ZN(n525) );
  NAND2_X1 U159 ( .A1(\mem[6][4] ), .A2(n459), .ZN(n686) );
  OAI21_X1 U160 ( .B1(n484), .B2(n691), .A(n685), .ZN(n524) );
  NAND2_X1 U161 ( .A1(\mem[6][5] ), .A2(n459), .ZN(n685) );
  OAI21_X1 U162 ( .B1(n483), .B2(n691), .A(n684), .ZN(n523) );
  NAND2_X1 U163 ( .A1(\mem[6][6] ), .A2(n459), .ZN(n684) );
  OAI21_X1 U164 ( .B1(n482), .B2(n691), .A(n683), .ZN(n522) );
  NAND2_X1 U165 ( .A1(\mem[6][7] ), .A2(n459), .ZN(n683) );
  OAI21_X1 U166 ( .B1(n481), .B2(n691), .A(n682), .ZN(n521) );
  NAND2_X1 U167 ( .A1(\mem[6][8] ), .A2(n459), .ZN(n682) );
  OAI21_X1 U168 ( .B1(n480), .B2(n691), .A(n681), .ZN(n520) );
  NAND2_X1 U169 ( .A1(\mem[6][9] ), .A2(n459), .ZN(n681) );
  OAI21_X1 U170 ( .B1(n479), .B2(n691), .A(n680), .ZN(n519) );
  NAND2_X1 U171 ( .A1(\mem[6][10] ), .A2(n459), .ZN(n680) );
  OAI21_X1 U172 ( .B1(n478), .B2(n691), .A(n679), .ZN(n518) );
  NAND2_X1 U173 ( .A1(\mem[6][11] ), .A2(n459), .ZN(n679) );
  OAI21_X1 U174 ( .B1(n477), .B2(n691), .A(n678), .ZN(n517) );
  NAND2_X1 U175 ( .A1(\mem[6][12] ), .A2(n691), .ZN(n678) );
  OAI21_X1 U176 ( .B1(n476), .B2(n459), .A(n677), .ZN(n516) );
  NAND2_X1 U177 ( .A1(\mem[6][13] ), .A2(n691), .ZN(n677) );
  OAI21_X1 U178 ( .B1(n475), .B2(n459), .A(n676), .ZN(n515) );
  NAND2_X1 U179 ( .A1(\mem[6][14] ), .A2(n691), .ZN(n676) );
  OAI21_X1 U180 ( .B1(n474), .B2(n691), .A(n675), .ZN(n514) );
  NAND2_X1 U181 ( .A1(\mem[6][15] ), .A2(n691), .ZN(n675) );
  OAI21_X1 U182 ( .B1(n473), .B2(n691), .A(n674), .ZN(n513) );
  NAND2_X1 U183 ( .A1(\mem[6][16] ), .A2(n691), .ZN(n674) );
  OAI21_X1 U184 ( .B1(n472), .B2(n691), .A(n673), .ZN(n512) );
  NAND2_X1 U185 ( .A1(\mem[6][17] ), .A2(n691), .ZN(n673) );
  OAI21_X1 U186 ( .B1(n471), .B2(n691), .A(n672), .ZN(n511) );
  NAND2_X1 U187 ( .A1(\mem[6][18] ), .A2(n691), .ZN(n672) );
  OAI21_X1 U188 ( .B1(n470), .B2(n691), .A(n671), .ZN(n510) );
  NAND2_X1 U189 ( .A1(\mem[6][19] ), .A2(n459), .ZN(n671) );
  OAI21_X1 U190 ( .B1(n489), .B2(n670), .A(n669), .ZN(n509) );
  NAND2_X1 U191 ( .A1(\mem[7][0] ), .A2(n670), .ZN(n669) );
  OAI21_X1 U192 ( .B1(n488), .B2(n458), .A(n668), .ZN(n508) );
  NAND2_X1 U193 ( .A1(\mem[7][1] ), .A2(n670), .ZN(n668) );
  OAI21_X1 U194 ( .B1(n487), .B2(n458), .A(n667), .ZN(n507) );
  NAND2_X1 U195 ( .A1(\mem[7][2] ), .A2(n670), .ZN(n667) );
  OAI21_X1 U196 ( .B1(n486), .B2(n458), .A(n666), .ZN(n506) );
  NAND2_X1 U197 ( .A1(\mem[7][3] ), .A2(n670), .ZN(n666) );
  OAI21_X1 U198 ( .B1(n485), .B2(n458), .A(n665), .ZN(n505) );
  NAND2_X1 U199 ( .A1(\mem[7][4] ), .A2(n670), .ZN(n665) );
  OAI21_X1 U200 ( .B1(n484), .B2(n458), .A(n664), .ZN(n504) );
  NAND2_X1 U201 ( .A1(\mem[7][5] ), .A2(n670), .ZN(n664) );
  OAI21_X1 U202 ( .B1(n483), .B2(n458), .A(n663), .ZN(n503) );
  NAND2_X1 U203 ( .A1(\mem[7][6] ), .A2(n670), .ZN(n663) );
  OAI21_X1 U204 ( .B1(n482), .B2(n458), .A(n662), .ZN(n502) );
  NAND2_X1 U205 ( .A1(\mem[7][7] ), .A2(n670), .ZN(n662) );
  OAI21_X1 U206 ( .B1(n481), .B2(n458), .A(n661), .ZN(n501) );
  NAND2_X1 U207 ( .A1(\mem[7][8] ), .A2(n670), .ZN(n661) );
  OAI21_X1 U208 ( .B1(n480), .B2(n670), .A(n660), .ZN(n500) );
  NAND2_X1 U209 ( .A1(\mem[7][9] ), .A2(n670), .ZN(n660) );
  OAI21_X1 U210 ( .B1(n479), .B2(n458), .A(n659), .ZN(n499) );
  NAND2_X1 U211 ( .A1(\mem[7][10] ), .A2(n670), .ZN(n659) );
  OAI21_X1 U212 ( .B1(n478), .B2(n458), .A(n658), .ZN(n498) );
  NAND2_X1 U213 ( .A1(\mem[7][11] ), .A2(n670), .ZN(n658) );
  OAI21_X1 U214 ( .B1(n477), .B2(n670), .A(n657), .ZN(n497) );
  NAND2_X1 U215 ( .A1(\mem[7][12] ), .A2(n670), .ZN(n657) );
  OAI21_X1 U216 ( .B1(n476), .B2(n458), .A(n656), .ZN(n496) );
  NAND2_X1 U217 ( .A1(\mem[7][13] ), .A2(n670), .ZN(n656) );
  OAI21_X1 U218 ( .B1(n475), .B2(n670), .A(n655), .ZN(n495) );
  NAND2_X1 U219 ( .A1(\mem[7][14] ), .A2(n670), .ZN(n655) );
  OAI21_X1 U220 ( .B1(n474), .B2(n458), .A(n654), .ZN(n494) );
  NAND2_X1 U221 ( .A1(\mem[7][15] ), .A2(n670), .ZN(n654) );
  OAI21_X1 U222 ( .B1(n473), .B2(n458), .A(n653), .ZN(n493) );
  NAND2_X1 U223 ( .A1(\mem[7][16] ), .A2(n670), .ZN(n653) );
  OAI21_X1 U224 ( .B1(n472), .B2(n458), .A(n652), .ZN(n492) );
  NAND2_X1 U225 ( .A1(\mem[7][17] ), .A2(n670), .ZN(n652) );
  OAI21_X1 U226 ( .B1(n471), .B2(n458), .A(n651), .ZN(n491) );
  NAND2_X1 U227 ( .A1(\mem[7][18] ), .A2(n670), .ZN(n651) );
  OAI21_X1 U228 ( .B1(n470), .B2(n458), .A(n650), .ZN(n490) );
  NAND2_X1 U229 ( .A1(\mem[7][19] ), .A2(n670), .ZN(n650) );
  NAND2_X1 U230 ( .A1(wr_en), .A2(n469), .ZN(n735) );
  INV_X1 U231 ( .A(addr[3]), .ZN(n469) );
  OAI21_X1 U232 ( .B1(n465), .B2(n489), .A(n819), .ZN(n649) );
  NAND2_X1 U233 ( .A1(\mem[0][0] ), .A2(n465), .ZN(n819) );
  OAI21_X1 U234 ( .B1(n820), .B2(n488), .A(n818), .ZN(n648) );
  NAND2_X1 U235 ( .A1(\mem[0][1] ), .A2(n465), .ZN(n818) );
  OAI21_X1 U236 ( .B1(n820), .B2(n487), .A(n817), .ZN(n647) );
  NAND2_X1 U237 ( .A1(\mem[0][2] ), .A2(n465), .ZN(n817) );
  OAI21_X1 U238 ( .B1(n820), .B2(n486), .A(n816), .ZN(n646) );
  NAND2_X1 U239 ( .A1(\mem[0][3] ), .A2(n465), .ZN(n816) );
  OAI21_X1 U240 ( .B1(n820), .B2(n485), .A(n815), .ZN(n645) );
  NAND2_X1 U241 ( .A1(\mem[0][4] ), .A2(n465), .ZN(n815) );
  OAI21_X1 U242 ( .B1(n820), .B2(n484), .A(n814), .ZN(n644) );
  NAND2_X1 U243 ( .A1(\mem[0][5] ), .A2(n465), .ZN(n814) );
  OAI21_X1 U244 ( .B1(n820), .B2(n483), .A(n813), .ZN(n643) );
  NAND2_X1 U245 ( .A1(\mem[0][6] ), .A2(n465), .ZN(n813) );
  OAI21_X1 U246 ( .B1(n820), .B2(n482), .A(n812), .ZN(n642) );
  NAND2_X1 U247 ( .A1(\mem[0][7] ), .A2(n465), .ZN(n812) );
  OAI21_X1 U248 ( .B1(n820), .B2(n481), .A(n811), .ZN(n641) );
  NAND2_X1 U249 ( .A1(\mem[0][8] ), .A2(n465), .ZN(n811) );
  OAI21_X1 U250 ( .B1(n820), .B2(n480), .A(n810), .ZN(n640) );
  NAND2_X1 U251 ( .A1(\mem[0][9] ), .A2(n465), .ZN(n810) );
  OAI21_X1 U252 ( .B1(n820), .B2(n479), .A(n809), .ZN(n639) );
  NAND2_X1 U253 ( .A1(\mem[0][10] ), .A2(n465), .ZN(n809) );
  OAI21_X1 U254 ( .B1(n820), .B2(n478), .A(n808), .ZN(n638) );
  NAND2_X1 U255 ( .A1(\mem[0][11] ), .A2(n465), .ZN(n808) );
  OAI21_X1 U256 ( .B1(n489), .B2(n798), .A(n797), .ZN(n629) );
  NAND2_X1 U257 ( .A1(\mem[1][0] ), .A2(n464), .ZN(n797) );
  OAI21_X1 U258 ( .B1(n488), .B2(n798), .A(n796), .ZN(n628) );
  NAND2_X1 U259 ( .A1(\mem[1][1] ), .A2(n464), .ZN(n796) );
  OAI21_X1 U260 ( .B1(n487), .B2(n798), .A(n795), .ZN(n627) );
  NAND2_X1 U261 ( .A1(\mem[1][2] ), .A2(n464), .ZN(n795) );
  OAI21_X1 U262 ( .B1(n486), .B2(n798), .A(n794), .ZN(n626) );
  NAND2_X1 U263 ( .A1(\mem[1][3] ), .A2(n464), .ZN(n794) );
  OAI21_X1 U264 ( .B1(n485), .B2(n798), .A(n793), .ZN(n625) );
  NAND2_X1 U265 ( .A1(\mem[1][4] ), .A2(n464), .ZN(n793) );
  OAI21_X1 U266 ( .B1(n484), .B2(n798), .A(n792), .ZN(n624) );
  NAND2_X1 U267 ( .A1(\mem[1][5] ), .A2(n464), .ZN(n792) );
  OAI21_X1 U268 ( .B1(n483), .B2(n798), .A(n791), .ZN(n623) );
  NAND2_X1 U269 ( .A1(\mem[1][6] ), .A2(n464), .ZN(n791) );
  OAI21_X1 U270 ( .B1(n482), .B2(n798), .A(n790), .ZN(n622) );
  NAND2_X1 U271 ( .A1(\mem[1][7] ), .A2(n464), .ZN(n790) );
  OAI21_X1 U272 ( .B1(n481), .B2(n798), .A(n789), .ZN(n621) );
  NAND2_X1 U273 ( .A1(\mem[1][8] ), .A2(n464), .ZN(n789) );
  OAI21_X1 U274 ( .B1(n480), .B2(n464), .A(n788), .ZN(n620) );
  NAND2_X1 U275 ( .A1(\mem[1][9] ), .A2(n464), .ZN(n788) );
  OAI21_X1 U276 ( .B1(n479), .B2(n798), .A(n787), .ZN(n619) );
  NAND2_X1 U277 ( .A1(\mem[1][10] ), .A2(n464), .ZN(n787) );
  OAI21_X1 U278 ( .B1(n478), .B2(n798), .A(n786), .ZN(n618) );
  NAND2_X1 U279 ( .A1(\mem[1][11] ), .A2(n464), .ZN(n786) );
  OAI21_X1 U280 ( .B1(n489), .B2(n777), .A(n776), .ZN(n609) );
  NAND2_X1 U281 ( .A1(\mem[2][0] ), .A2(n777), .ZN(n776) );
  OAI21_X1 U282 ( .B1(n488), .B2(n777), .A(n775), .ZN(n608) );
  NAND2_X1 U283 ( .A1(\mem[2][1] ), .A2(n777), .ZN(n775) );
  OAI21_X1 U284 ( .B1(n487), .B2(n777), .A(n774), .ZN(n607) );
  NAND2_X1 U285 ( .A1(\mem[2][2] ), .A2(n777), .ZN(n774) );
  OAI21_X1 U286 ( .B1(n486), .B2(n777), .A(n773), .ZN(n606) );
  NAND2_X1 U287 ( .A1(\mem[2][3] ), .A2(n463), .ZN(n773) );
  OAI21_X1 U288 ( .B1(n485), .B2(n777), .A(n772), .ZN(n605) );
  NAND2_X1 U289 ( .A1(\mem[2][4] ), .A2(n463), .ZN(n772) );
  OAI21_X1 U290 ( .B1(n484), .B2(n777), .A(n771), .ZN(n604) );
  NAND2_X1 U291 ( .A1(\mem[2][5] ), .A2(n463), .ZN(n771) );
  OAI21_X1 U292 ( .B1(n483), .B2(n777), .A(n770), .ZN(n603) );
  NAND2_X1 U293 ( .A1(\mem[2][6] ), .A2(n777), .ZN(n770) );
  OAI21_X1 U294 ( .B1(n482), .B2(n777), .A(n769), .ZN(n602) );
  NAND2_X1 U295 ( .A1(\mem[2][7] ), .A2(n777), .ZN(n769) );
  OAI21_X1 U296 ( .B1(n481), .B2(n777), .A(n768), .ZN(n601) );
  NAND2_X1 U297 ( .A1(\mem[2][8] ), .A2(n777), .ZN(n768) );
  OAI21_X1 U298 ( .B1(n480), .B2(n463), .A(n767), .ZN(n600) );
  NAND2_X1 U299 ( .A1(\mem[2][9] ), .A2(n463), .ZN(n767) );
  OAI21_X1 U300 ( .B1(n479), .B2(n777), .A(n766), .ZN(n599) );
  NAND2_X1 U301 ( .A1(\mem[2][10] ), .A2(n777), .ZN(n766) );
  OAI21_X1 U302 ( .B1(n478), .B2(n777), .A(n765), .ZN(n598) );
  NAND2_X1 U303 ( .A1(\mem[2][11] ), .A2(n777), .ZN(n765) );
  OAI21_X1 U304 ( .B1(n489), .B2(n756), .A(n755), .ZN(n589) );
  NAND2_X1 U305 ( .A1(\mem[3][0] ), .A2(n462), .ZN(n755) );
  OAI21_X1 U306 ( .B1(n488), .B2(n756), .A(n754), .ZN(n588) );
  NAND2_X1 U307 ( .A1(\mem[3][1] ), .A2(n462), .ZN(n754) );
  OAI21_X1 U308 ( .B1(n487), .B2(n756), .A(n753), .ZN(n587) );
  NAND2_X1 U309 ( .A1(\mem[3][2] ), .A2(n462), .ZN(n753) );
  OAI21_X1 U310 ( .B1(n486), .B2(n756), .A(n752), .ZN(n586) );
  NAND2_X1 U311 ( .A1(\mem[3][3] ), .A2(n462), .ZN(n752) );
  OAI21_X1 U312 ( .B1(n485), .B2(n756), .A(n751), .ZN(n585) );
  NAND2_X1 U313 ( .A1(\mem[3][4] ), .A2(n462), .ZN(n751) );
  OAI21_X1 U314 ( .B1(n484), .B2(n756), .A(n750), .ZN(n584) );
  NAND2_X1 U315 ( .A1(\mem[3][5] ), .A2(n462), .ZN(n750) );
  OAI21_X1 U316 ( .B1(n483), .B2(n756), .A(n749), .ZN(n583) );
  NAND2_X1 U317 ( .A1(\mem[3][6] ), .A2(n462), .ZN(n749) );
  OAI21_X1 U318 ( .B1(n482), .B2(n756), .A(n748), .ZN(n582) );
  NAND2_X1 U319 ( .A1(\mem[3][7] ), .A2(n462), .ZN(n748) );
  OAI21_X1 U320 ( .B1(n481), .B2(n756), .A(n747), .ZN(n581) );
  NAND2_X1 U321 ( .A1(\mem[3][8] ), .A2(n462), .ZN(n747) );
  OAI21_X1 U322 ( .B1(n480), .B2(n462), .A(n746), .ZN(n580) );
  NAND2_X1 U323 ( .A1(\mem[3][9] ), .A2(n462), .ZN(n746) );
  OAI21_X1 U324 ( .B1(n479), .B2(n756), .A(n745), .ZN(n579) );
  NAND2_X1 U325 ( .A1(\mem[3][10] ), .A2(n462), .ZN(n745) );
  OAI21_X1 U326 ( .B1(n478), .B2(n756), .A(n744), .ZN(n578) );
  NAND2_X1 U327 ( .A1(\mem[3][11] ), .A2(n462), .ZN(n744) );
  OAI21_X1 U328 ( .B1(n820), .B2(n477), .A(n807), .ZN(n637) );
  NAND2_X1 U329 ( .A1(\mem[0][12] ), .A2(n820), .ZN(n807) );
  OAI21_X1 U330 ( .B1(n820), .B2(n476), .A(n806), .ZN(n636) );
  NAND2_X1 U331 ( .A1(\mem[0][13] ), .A2(n820), .ZN(n806) );
  OAI21_X1 U332 ( .B1(n465), .B2(n475), .A(n805), .ZN(n635) );
  NAND2_X1 U333 ( .A1(\mem[0][14] ), .A2(n820), .ZN(n805) );
  OAI21_X1 U334 ( .B1(n820), .B2(n474), .A(n804), .ZN(n634) );
  NAND2_X1 U335 ( .A1(\mem[0][15] ), .A2(n465), .ZN(n804) );
  OAI21_X1 U336 ( .B1(n820), .B2(n473), .A(n803), .ZN(n633) );
  NAND2_X1 U337 ( .A1(\mem[0][16] ), .A2(n820), .ZN(n803) );
  OAI21_X1 U338 ( .B1(n820), .B2(n472), .A(n802), .ZN(n632) );
  NAND2_X1 U339 ( .A1(\mem[0][17] ), .A2(n820), .ZN(n802) );
  OAI21_X1 U340 ( .B1(n820), .B2(n471), .A(n801), .ZN(n631) );
  NAND2_X1 U341 ( .A1(\mem[0][18] ), .A2(n820), .ZN(n801) );
  OAI21_X1 U342 ( .B1(n820), .B2(n470), .A(n800), .ZN(n630) );
  NAND2_X1 U343 ( .A1(\mem[0][19] ), .A2(n465), .ZN(n800) );
  INV_X1 U344 ( .A(data_in[0]), .ZN(n489) );
  INV_X1 U345 ( .A(data_in[1]), .ZN(n488) );
  INV_X1 U346 ( .A(data_in[2]), .ZN(n487) );
  INV_X1 U347 ( .A(data_in[3]), .ZN(n486) );
  INV_X1 U348 ( .A(data_in[4]), .ZN(n485) );
  INV_X1 U349 ( .A(data_in[5]), .ZN(n484) );
  INV_X1 U358 ( .A(data_in[6]), .ZN(n483) );
  INV_X1 U359 ( .A(data_in[7]), .ZN(n482) );
  INV_X1 U360 ( .A(data_in[8]), .ZN(n481) );
  INV_X1 U361 ( .A(data_in[9]), .ZN(n480) );
  INV_X1 U362 ( .A(data_in[10]), .ZN(n479) );
  INV_X1 U363 ( .A(data_in[11]), .ZN(n478) );
  INV_X1 U364 ( .A(data_in[12]), .ZN(n477) );
  INV_X1 U365 ( .A(data_in[13]), .ZN(n476) );
  INV_X1 U366 ( .A(data_in[14]), .ZN(n475) );
  INV_X1 U367 ( .A(data_in[15]), .ZN(n474) );
  INV_X1 U368 ( .A(data_in[16]), .ZN(n473) );
  INV_X1 U369 ( .A(data_in[17]), .ZN(n472) );
  INV_X1 U370 ( .A(data_in[18]), .ZN(n471) );
  INV_X1 U371 ( .A(data_in[19]), .ZN(n470) );
  MUX2_X1 U372 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n456), .Z(n1) );
  MUX2_X1 U373 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n455), .Z(n2) );
  MUX2_X1 U374 ( .A(n2), .B(n1), .S(n453), .Z(n3) );
  MUX2_X1 U375 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n457), .Z(n4) );
  MUX2_X1 U376 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n455), .Z(n5) );
  MUX2_X1 U377 ( .A(n5), .B(n4), .S(n453), .Z(n6) );
  MUX2_X1 U378 ( .A(n6), .B(n3), .S(N12), .Z(N32) );
  MUX2_X1 U379 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n455), .Z(n7) );
  MUX2_X1 U380 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n454), .Z(n8) );
  MUX2_X1 U381 ( .A(n8), .B(n7), .S(n453), .Z(n9) );
  MUX2_X1 U382 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n457), .Z(n10) );
  MUX2_X1 U383 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n456), .Z(n11) );
  MUX2_X1 U384 ( .A(n11), .B(n10), .S(n453), .Z(n12) );
  MUX2_X1 U385 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n454), .Z(n13) );
  MUX2_X1 U386 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n454), .Z(n14) );
  MUX2_X1 U387 ( .A(n14), .B(n13), .S(n453), .Z(n15) );
  MUX2_X1 U388 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n454), .Z(n16) );
  MUX2_X1 U389 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n454), .Z(n17) );
  MUX2_X1 U390 ( .A(n17), .B(n16), .S(n453), .Z(n18) );
  MUX2_X1 U391 ( .A(n18), .B(n15), .S(N12), .Z(N30) );
  MUX2_X1 U392 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n454), .Z(n19) );
  MUX2_X1 U393 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n454), .Z(n20) );
  MUX2_X1 U394 ( .A(n20), .B(n19), .S(n453), .Z(n21) );
  MUX2_X1 U395 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n454), .Z(n22) );
  MUX2_X1 U396 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n454), .Z(n23) );
  MUX2_X1 U397 ( .A(n23), .B(n22), .S(n453), .Z(n24) );
  MUX2_X1 U398 ( .A(n24), .B(n21), .S(N12), .Z(N29) );
  MUX2_X1 U399 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n454), .Z(n356) );
  MUX2_X1 U400 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n454), .Z(n357) );
  MUX2_X1 U401 ( .A(n357), .B(n356), .S(n453), .Z(n358) );
  MUX2_X1 U402 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n454), .Z(n359) );
  MUX2_X1 U403 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n454), .Z(n360) );
  MUX2_X1 U404 ( .A(n360), .B(n359), .S(n453), .Z(n361) );
  MUX2_X1 U405 ( .A(n361), .B(n358), .S(N12), .Z(N28) );
  MUX2_X1 U406 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n455), .Z(n362) );
  MUX2_X1 U407 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n456), .Z(n363) );
  MUX2_X1 U408 ( .A(n363), .B(n362), .S(n453), .Z(n364) );
  MUX2_X1 U409 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n456), .Z(n365) );
  MUX2_X1 U410 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n455), .Z(n366) );
  MUX2_X1 U411 ( .A(n366), .B(n365), .S(n453), .Z(n367) );
  MUX2_X1 U412 ( .A(n367), .B(n364), .S(N12), .Z(N27) );
  MUX2_X1 U413 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n454), .Z(n368) );
  MUX2_X1 U414 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n457), .Z(n369) );
  MUX2_X1 U415 ( .A(n369), .B(n368), .S(n453), .Z(n370) );
  MUX2_X1 U416 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n457), .Z(n371) );
  MUX2_X1 U417 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n456), .Z(n372) );
  MUX2_X1 U418 ( .A(n372), .B(n371), .S(n453), .Z(n373) );
  MUX2_X1 U419 ( .A(n373), .B(n370), .S(N12), .Z(N26) );
  MUX2_X1 U420 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n455), .Z(n374) );
  MUX2_X1 U421 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n454), .Z(n375) );
  MUX2_X1 U422 ( .A(n375), .B(n374), .S(n453), .Z(n376) );
  MUX2_X1 U423 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n454), .Z(n377) );
  MUX2_X1 U424 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n456), .Z(n378) );
  MUX2_X1 U425 ( .A(n378), .B(n377), .S(n453), .Z(n379) );
  MUX2_X1 U426 ( .A(n379), .B(n376), .S(N12), .Z(N25) );
  MUX2_X1 U427 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n454), .Z(n380) );
  MUX2_X1 U428 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n456), .Z(n381) );
  MUX2_X1 U429 ( .A(n381), .B(n380), .S(n452), .Z(n382) );
  MUX2_X1 U430 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n454), .Z(n383) );
  MUX2_X1 U431 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n454), .Z(n384) );
  MUX2_X1 U432 ( .A(n384), .B(n383), .S(n452), .Z(n385) );
  MUX2_X1 U433 ( .A(n385), .B(n382), .S(N12), .Z(N24) );
  MUX2_X1 U434 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n457), .Z(n386) );
  MUX2_X1 U435 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n454), .Z(n387) );
  MUX2_X1 U436 ( .A(n387), .B(n386), .S(n452), .Z(n388) );
  MUX2_X1 U437 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n455), .Z(n389) );
  MUX2_X1 U438 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n456), .Z(n390) );
  MUX2_X1 U439 ( .A(n390), .B(n389), .S(n452), .Z(n391) );
  MUX2_X1 U440 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n457), .Z(n392) );
  MUX2_X1 U441 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n457), .Z(n393) );
  MUX2_X1 U442 ( .A(n393), .B(n392), .S(n452), .Z(n394) );
  MUX2_X1 U443 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n455), .Z(n395) );
  MUX2_X1 U444 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n457), .Z(n396) );
  MUX2_X1 U445 ( .A(n396), .B(n395), .S(n452), .Z(n397) );
  MUX2_X1 U446 ( .A(n397), .B(n394), .S(N12), .Z(N22) );
  MUX2_X1 U447 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n455), .Z(n398) );
  MUX2_X1 U448 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n455), .Z(n399) );
  MUX2_X1 U449 ( .A(n399), .B(n398), .S(n452), .Z(n400) );
  MUX2_X1 U450 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n455), .Z(n401) );
  MUX2_X1 U451 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n455), .Z(n402) );
  MUX2_X1 U452 ( .A(n402), .B(n401), .S(n452), .Z(n403) );
  MUX2_X1 U453 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n455), .Z(n404) );
  MUX2_X1 U454 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n455), .Z(n405) );
  MUX2_X1 U455 ( .A(n405), .B(n404), .S(n452), .Z(n406) );
  MUX2_X1 U456 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n455), .Z(n407) );
  MUX2_X1 U457 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n455), .Z(n408) );
  MUX2_X1 U458 ( .A(n408), .B(n407), .S(n452), .Z(n409) );
  MUX2_X1 U459 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n455), .Z(n410) );
  MUX2_X1 U460 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n455), .Z(n411) );
  MUX2_X1 U461 ( .A(n411), .B(n410), .S(n452), .Z(n412) );
  MUX2_X1 U462 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n455), .Z(n413) );
  MUX2_X1 U463 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n455), .Z(n414) );
  MUX2_X1 U464 ( .A(n414), .B(n413), .S(n452), .Z(n415) );
  MUX2_X1 U465 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n456), .Z(n416) );
  MUX2_X1 U466 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n456), .Z(n417) );
  MUX2_X1 U467 ( .A(n417), .B(n416), .S(n453), .Z(n418) );
  MUX2_X1 U468 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n456), .Z(n419) );
  MUX2_X1 U469 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n456), .Z(n420) );
  MUX2_X1 U470 ( .A(n420), .B(n419), .S(N11), .Z(n421) );
  MUX2_X1 U471 ( .A(n421), .B(n418), .S(N12), .Z(N18) );
  MUX2_X1 U472 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n456), .Z(n422) );
  MUX2_X1 U473 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n456), .Z(n423) );
  MUX2_X1 U474 ( .A(n423), .B(n422), .S(n453), .Z(n424) );
  MUX2_X1 U475 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n456), .Z(n425) );
  MUX2_X1 U476 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n456), .Z(n426) );
  MUX2_X1 U477 ( .A(n426), .B(n425), .S(N11), .Z(n427) );
  MUX2_X1 U478 ( .A(n427), .B(n424), .S(N12), .Z(N17) );
  MUX2_X1 U479 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n456), .Z(n428) );
  MUX2_X1 U480 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n456), .Z(n429) );
  MUX2_X1 U481 ( .A(n429), .B(n428), .S(n453), .Z(n430) );
  MUX2_X1 U482 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n456), .Z(n431) );
  MUX2_X1 U483 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n456), .Z(n432) );
  MUX2_X1 U484 ( .A(n432), .B(n431), .S(N11), .Z(n433) );
  MUX2_X1 U485 ( .A(n433), .B(n430), .S(N12), .Z(N16) );
  MUX2_X1 U486 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n457), .Z(n434) );
  MUX2_X1 U487 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n457), .Z(n435) );
  MUX2_X1 U488 ( .A(n435), .B(n434), .S(n453), .Z(n436) );
  MUX2_X1 U489 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n457), .Z(n437) );
  MUX2_X1 U490 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n457), .Z(n438) );
  MUX2_X1 U491 ( .A(n438), .B(n437), .S(N11), .Z(n439) );
  MUX2_X1 U492 ( .A(n439), .B(n436), .S(N12), .Z(N15) );
  MUX2_X1 U493 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n457), .Z(n440) );
  MUX2_X1 U494 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n457), .Z(n441) );
  MUX2_X1 U495 ( .A(n441), .B(n440), .S(n453), .Z(n442) );
  MUX2_X1 U496 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n457), .Z(n443) );
  MUX2_X1 U497 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n457), .Z(n444) );
  MUX2_X1 U498 ( .A(n444), .B(n443), .S(N11), .Z(n445) );
  MUX2_X1 U499 ( .A(n445), .B(n442), .S(N12), .Z(N14) );
  MUX2_X1 U500 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n457), .Z(n446) );
  MUX2_X1 U501 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n457), .Z(n447) );
  MUX2_X1 U502 ( .A(n447), .B(n446), .S(n453), .Z(n448) );
  MUX2_X1 U503 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n457), .Z(n449) );
  MUX2_X1 U504 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n457), .Z(n450) );
  MUX2_X1 U505 ( .A(n450), .B(n449), .S(N11), .Z(n451) );
  MUX2_X1 U506 ( .A(n451), .B(n448), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE4_6 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N13, N14, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N28, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[19]  ( .D(N13), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[15]  ( .D(N17), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N19), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N20), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N21), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N23), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N25), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[0]  ( .D(N32), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n490), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n491), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n492), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n493), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n494), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n495), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n496), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n497), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n498), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n499), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n500), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n501), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n502), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n503), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n504), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n505), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n506), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n507), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n508), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n509), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n510), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n511), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n512), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n513), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n514), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n515), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n516), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n517), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n518), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n519), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n520), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n521), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n522), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n523), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n524), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n525), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n526), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n527), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n528), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n529), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n530), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n531), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n532), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n533), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n534), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n535), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n536), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n537), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n538), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n539), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n540), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n541), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n542), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n543), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n544), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n545), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n546), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n547), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n548), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n549), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n550), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n551), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n552), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n553), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n554), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n555), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n556), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n557), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n558), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n559), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n560), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n561), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n562), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n563), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n564), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n565), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n566), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n567), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n568), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n569), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n570), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n571), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n572), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n573), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n574), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n575), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n576), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n577), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n578), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n579), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n580), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n581), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n582), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n583), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n584), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n585), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n586), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n587), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n588), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n589), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n590), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n591), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n592), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n593), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n594), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n595), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n596), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n597), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n598), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n599), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n600), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n601), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n602), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n603), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n604), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n605), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n606), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n607), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n608), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n609), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n610), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n611), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n612), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n613), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n614), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n615), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n616), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n617), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n618), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n619), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n620), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n621), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n622), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n623), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n624), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n625), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n626), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n627), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n628), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n629), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n630), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n631), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n632), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n633), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n634), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n635), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n636), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n637), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n638), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n639), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n640), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n641), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n642), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n643), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n644), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n645), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n646), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n647), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n648), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n649), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U350 ( .A1(n466), .A2(n467), .A3(n799), .ZN(n820) );
  NAND3_X1 U351 ( .A1(n799), .A2(n467), .A3(N10), .ZN(n798) );
  NAND3_X1 U352 ( .A1(n799), .A2(n466), .A3(N11), .ZN(n777) );
  NAND3_X1 U353 ( .A1(N10), .A2(n799), .A3(N11), .ZN(n756) );
  NAND3_X1 U354 ( .A1(n466), .A2(n467), .A3(n713), .ZN(n734) );
  NAND3_X1 U355 ( .A1(N10), .A2(n467), .A3(n713), .ZN(n712) );
  NAND3_X1 U356 ( .A1(N11), .A2(n466), .A3(n713), .ZN(n691) );
  NAND3_X1 U357 ( .A1(N11), .A2(N10), .A3(n713), .ZN(n670) );
  SDFF_X1 \data_out_reg[17]  ( .D(n436), .SI(n439), .SE(n468), .CK(clk), .Q(
        data_out[17]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n15), .SI(n18), .SE(n468), .CK(clk), .Q(
        data_out[2]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n9), .SI(n12), .SE(n468), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n364), .SI(n367), .SE(n468), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n21), .SI(n24), .SE(n468), .CK(clk), .Q(
        data_out[3]) );
  BUF_X1 U3 ( .A(n820), .Z(n465) );
  BUF_X1 U4 ( .A(n756), .Z(n462) );
  BUF_X1 U5 ( .A(n691), .Z(n459) );
  BUF_X1 U6 ( .A(n453), .Z(n452) );
  BUF_X1 U7 ( .A(N10), .Z(n454) );
  BUF_X1 U8 ( .A(N10), .Z(n455) );
  BUF_X1 U9 ( .A(N10), .Z(n456) );
  BUF_X1 U10 ( .A(N10), .Z(n457) );
  BUF_X1 U11 ( .A(N11), .Z(n453) );
  BUF_X1 U12 ( .A(n798), .Z(n464) );
  BUF_X1 U13 ( .A(n777), .Z(n463) );
  BUF_X1 U14 ( .A(n670), .Z(n458) );
  BUF_X1 U15 ( .A(n734), .Z(n461) );
  BUF_X1 U16 ( .A(n712), .Z(n460) );
  NOR2_X1 U17 ( .A1(n735), .A2(N12), .ZN(n799) );
  NOR2_X1 U18 ( .A1(n468), .A2(n735), .ZN(n713) );
  INV_X1 U19 ( .A(N12), .ZN(n468) );
  INV_X1 U20 ( .A(N11), .ZN(n467) );
  INV_X1 U21 ( .A(N10), .ZN(n466) );
  OAI21_X1 U22 ( .B1(n477), .B2(n798), .A(n785), .ZN(n617) );
  NAND2_X1 U23 ( .A1(\mem[1][12] ), .A2(n798), .ZN(n785) );
  OAI21_X1 U24 ( .B1(n476), .B2(n798), .A(n784), .ZN(n616) );
  NAND2_X1 U25 ( .A1(\mem[1][13] ), .A2(n798), .ZN(n784) );
  OAI21_X1 U26 ( .B1(n475), .B2(n798), .A(n783), .ZN(n615) );
  NAND2_X1 U27 ( .A1(\mem[1][14] ), .A2(n798), .ZN(n783) );
  OAI21_X1 U28 ( .B1(n474), .B2(n464), .A(n782), .ZN(n614) );
  NAND2_X1 U29 ( .A1(\mem[1][15] ), .A2(n798), .ZN(n782) );
  OAI21_X1 U30 ( .B1(n473), .B2(n798), .A(n781), .ZN(n613) );
  NAND2_X1 U31 ( .A1(\mem[1][16] ), .A2(n464), .ZN(n781) );
  OAI21_X1 U32 ( .B1(n472), .B2(n798), .A(n780), .ZN(n612) );
  NAND2_X1 U33 ( .A1(\mem[1][17] ), .A2(n798), .ZN(n780) );
  OAI21_X1 U34 ( .B1(n471), .B2(n798), .A(n779), .ZN(n611) );
  NAND2_X1 U35 ( .A1(\mem[1][18] ), .A2(n798), .ZN(n779) );
  OAI21_X1 U36 ( .B1(n470), .B2(n798), .A(n778), .ZN(n610) );
  NAND2_X1 U37 ( .A1(\mem[1][19] ), .A2(n464), .ZN(n778) );
  OAI21_X1 U38 ( .B1(n477), .B2(n777), .A(n764), .ZN(n597) );
  NAND2_X1 U39 ( .A1(\mem[2][12] ), .A2(n777), .ZN(n764) );
  OAI21_X1 U40 ( .B1(n476), .B2(n777), .A(n763), .ZN(n596) );
  NAND2_X1 U41 ( .A1(\mem[2][13] ), .A2(n777), .ZN(n763) );
  OAI21_X1 U42 ( .B1(n475), .B2(n777), .A(n762), .ZN(n595) );
  NAND2_X1 U43 ( .A1(\mem[2][14] ), .A2(n777), .ZN(n762) );
  OAI21_X1 U44 ( .B1(n474), .B2(n463), .A(n761), .ZN(n594) );
  NAND2_X1 U45 ( .A1(\mem[2][15] ), .A2(n777), .ZN(n761) );
  OAI21_X1 U46 ( .B1(n473), .B2(n777), .A(n760), .ZN(n593) );
  NAND2_X1 U47 ( .A1(\mem[2][16] ), .A2(n463), .ZN(n760) );
  OAI21_X1 U48 ( .B1(n472), .B2(n777), .A(n759), .ZN(n592) );
  NAND2_X1 U49 ( .A1(\mem[2][17] ), .A2(n777), .ZN(n759) );
  OAI21_X1 U50 ( .B1(n471), .B2(n777), .A(n758), .ZN(n591) );
  NAND2_X1 U51 ( .A1(\mem[2][18] ), .A2(n777), .ZN(n758) );
  OAI21_X1 U52 ( .B1(n470), .B2(n777), .A(n757), .ZN(n590) );
  NAND2_X1 U53 ( .A1(\mem[2][19] ), .A2(n463), .ZN(n757) );
  OAI21_X1 U54 ( .B1(n477), .B2(n462), .A(n743), .ZN(n577) );
  NAND2_X1 U55 ( .A1(\mem[3][12] ), .A2(n462), .ZN(n743) );
  OAI21_X1 U56 ( .B1(n476), .B2(n462), .A(n742), .ZN(n576) );
  NAND2_X1 U57 ( .A1(\mem[3][13] ), .A2(n462), .ZN(n742) );
  OAI21_X1 U58 ( .B1(n475), .B2(n462), .A(n741), .ZN(n575) );
  NAND2_X1 U59 ( .A1(\mem[3][14] ), .A2(n462), .ZN(n741) );
  OAI21_X1 U60 ( .B1(n474), .B2(n756), .A(n740), .ZN(n574) );
  NAND2_X1 U61 ( .A1(\mem[3][15] ), .A2(n462), .ZN(n740) );
  OAI21_X1 U62 ( .B1(n473), .B2(n756), .A(n739), .ZN(n573) );
  NAND2_X1 U63 ( .A1(\mem[3][16] ), .A2(n462), .ZN(n739) );
  OAI21_X1 U64 ( .B1(n472), .B2(n756), .A(n738), .ZN(n572) );
  NAND2_X1 U65 ( .A1(\mem[3][17] ), .A2(n462), .ZN(n738) );
  OAI21_X1 U66 ( .B1(n471), .B2(n756), .A(n737), .ZN(n571) );
  NAND2_X1 U67 ( .A1(\mem[3][18] ), .A2(n462), .ZN(n737) );
  OAI21_X1 U68 ( .B1(n470), .B2(n756), .A(n736), .ZN(n570) );
  NAND2_X1 U69 ( .A1(\mem[3][19] ), .A2(n462), .ZN(n736) );
  OAI21_X1 U70 ( .B1(n489), .B2(n734), .A(n733), .ZN(n569) );
  NAND2_X1 U71 ( .A1(\mem[4][0] ), .A2(n461), .ZN(n733) );
  OAI21_X1 U72 ( .B1(n488), .B2(n734), .A(n732), .ZN(n568) );
  NAND2_X1 U73 ( .A1(\mem[4][1] ), .A2(n461), .ZN(n732) );
  OAI21_X1 U74 ( .B1(n487), .B2(n734), .A(n731), .ZN(n567) );
  NAND2_X1 U75 ( .A1(\mem[4][2] ), .A2(n461), .ZN(n731) );
  OAI21_X1 U76 ( .B1(n486), .B2(n734), .A(n730), .ZN(n566) );
  NAND2_X1 U77 ( .A1(\mem[4][3] ), .A2(n461), .ZN(n730) );
  OAI21_X1 U78 ( .B1(n485), .B2(n461), .A(n729), .ZN(n565) );
  NAND2_X1 U79 ( .A1(\mem[4][4] ), .A2(n461), .ZN(n729) );
  OAI21_X1 U80 ( .B1(n484), .B2(n734), .A(n728), .ZN(n564) );
  NAND2_X1 U81 ( .A1(\mem[4][5] ), .A2(n461), .ZN(n728) );
  OAI21_X1 U82 ( .B1(n483), .B2(n734), .A(n727), .ZN(n563) );
  NAND2_X1 U83 ( .A1(\mem[4][6] ), .A2(n461), .ZN(n727) );
  OAI21_X1 U84 ( .B1(n482), .B2(n734), .A(n726), .ZN(n562) );
  NAND2_X1 U85 ( .A1(\mem[4][7] ), .A2(n461), .ZN(n726) );
  OAI21_X1 U86 ( .B1(n481), .B2(n734), .A(n725), .ZN(n561) );
  NAND2_X1 U87 ( .A1(\mem[4][8] ), .A2(n461), .ZN(n725) );
  OAI21_X1 U88 ( .B1(n480), .B2(n734), .A(n724), .ZN(n560) );
  NAND2_X1 U89 ( .A1(\mem[4][9] ), .A2(n461), .ZN(n724) );
  OAI21_X1 U90 ( .B1(n479), .B2(n734), .A(n723), .ZN(n559) );
  NAND2_X1 U91 ( .A1(\mem[4][10] ), .A2(n461), .ZN(n723) );
  OAI21_X1 U92 ( .B1(n478), .B2(n734), .A(n722), .ZN(n558) );
  NAND2_X1 U93 ( .A1(\mem[4][11] ), .A2(n461), .ZN(n722) );
  OAI21_X1 U94 ( .B1(n477), .B2(n734), .A(n721), .ZN(n557) );
  NAND2_X1 U95 ( .A1(\mem[4][12] ), .A2(n734), .ZN(n721) );
  OAI21_X1 U96 ( .B1(n476), .B2(n461), .A(n720), .ZN(n556) );
  NAND2_X1 U97 ( .A1(\mem[4][13] ), .A2(n734), .ZN(n720) );
  OAI21_X1 U98 ( .B1(n475), .B2(n461), .A(n719), .ZN(n555) );
  NAND2_X1 U99 ( .A1(\mem[4][14] ), .A2(n734), .ZN(n719) );
  OAI21_X1 U100 ( .B1(n474), .B2(n734), .A(n718), .ZN(n554) );
  NAND2_X1 U101 ( .A1(\mem[4][15] ), .A2(n734), .ZN(n718) );
  OAI21_X1 U102 ( .B1(n473), .B2(n734), .A(n717), .ZN(n553) );
  NAND2_X1 U103 ( .A1(\mem[4][16] ), .A2(n734), .ZN(n717) );
  OAI21_X1 U104 ( .B1(n472), .B2(n734), .A(n716), .ZN(n552) );
  NAND2_X1 U105 ( .A1(\mem[4][17] ), .A2(n734), .ZN(n716) );
  OAI21_X1 U106 ( .B1(n471), .B2(n734), .A(n715), .ZN(n551) );
  NAND2_X1 U107 ( .A1(\mem[4][18] ), .A2(n734), .ZN(n715) );
  OAI21_X1 U108 ( .B1(n470), .B2(n734), .A(n714), .ZN(n550) );
  NAND2_X1 U109 ( .A1(\mem[4][19] ), .A2(n461), .ZN(n714) );
  OAI21_X1 U110 ( .B1(n489), .B2(n712), .A(n711), .ZN(n549) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n460), .ZN(n711) );
  OAI21_X1 U112 ( .B1(n488), .B2(n712), .A(n710), .ZN(n548) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n460), .ZN(n710) );
  OAI21_X1 U114 ( .B1(n487), .B2(n712), .A(n709), .ZN(n547) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n460), .ZN(n709) );
  OAI21_X1 U116 ( .B1(n486), .B2(n712), .A(n708), .ZN(n546) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n460), .ZN(n708) );
  OAI21_X1 U118 ( .B1(n485), .B2(n460), .A(n707), .ZN(n545) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n460), .ZN(n707) );
  OAI21_X1 U120 ( .B1(n484), .B2(n712), .A(n706), .ZN(n544) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n460), .ZN(n706) );
  OAI21_X1 U122 ( .B1(n483), .B2(n712), .A(n705), .ZN(n543) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n460), .ZN(n705) );
  OAI21_X1 U124 ( .B1(n482), .B2(n712), .A(n704), .ZN(n542) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n460), .ZN(n704) );
  OAI21_X1 U126 ( .B1(n481), .B2(n712), .A(n703), .ZN(n541) );
  NAND2_X1 U127 ( .A1(\mem[5][8] ), .A2(n460), .ZN(n703) );
  OAI21_X1 U128 ( .B1(n480), .B2(n712), .A(n702), .ZN(n540) );
  NAND2_X1 U129 ( .A1(\mem[5][9] ), .A2(n460), .ZN(n702) );
  OAI21_X1 U130 ( .B1(n479), .B2(n712), .A(n701), .ZN(n539) );
  NAND2_X1 U131 ( .A1(\mem[5][10] ), .A2(n460), .ZN(n701) );
  OAI21_X1 U132 ( .B1(n478), .B2(n712), .A(n700), .ZN(n538) );
  NAND2_X1 U133 ( .A1(\mem[5][11] ), .A2(n460), .ZN(n700) );
  OAI21_X1 U134 ( .B1(n477), .B2(n712), .A(n699), .ZN(n537) );
  NAND2_X1 U135 ( .A1(\mem[5][12] ), .A2(n712), .ZN(n699) );
  OAI21_X1 U136 ( .B1(n476), .B2(n460), .A(n698), .ZN(n536) );
  NAND2_X1 U137 ( .A1(\mem[5][13] ), .A2(n712), .ZN(n698) );
  OAI21_X1 U138 ( .B1(n475), .B2(n460), .A(n697), .ZN(n535) );
  NAND2_X1 U139 ( .A1(\mem[5][14] ), .A2(n712), .ZN(n697) );
  OAI21_X1 U140 ( .B1(n474), .B2(n712), .A(n696), .ZN(n534) );
  NAND2_X1 U141 ( .A1(\mem[5][15] ), .A2(n712), .ZN(n696) );
  OAI21_X1 U142 ( .B1(n473), .B2(n712), .A(n695), .ZN(n533) );
  NAND2_X1 U143 ( .A1(\mem[5][16] ), .A2(n712), .ZN(n695) );
  OAI21_X1 U144 ( .B1(n472), .B2(n712), .A(n694), .ZN(n532) );
  NAND2_X1 U145 ( .A1(\mem[5][17] ), .A2(n712), .ZN(n694) );
  OAI21_X1 U146 ( .B1(n471), .B2(n712), .A(n693), .ZN(n531) );
  NAND2_X1 U147 ( .A1(\mem[5][18] ), .A2(n712), .ZN(n693) );
  OAI21_X1 U148 ( .B1(n470), .B2(n712), .A(n692), .ZN(n530) );
  NAND2_X1 U149 ( .A1(\mem[5][19] ), .A2(n460), .ZN(n692) );
  OAI21_X1 U150 ( .B1(n489), .B2(n459), .A(n690), .ZN(n529) );
  NAND2_X1 U151 ( .A1(\mem[6][0] ), .A2(n459), .ZN(n690) );
  OAI21_X1 U152 ( .B1(n488), .B2(n459), .A(n689), .ZN(n528) );
  NAND2_X1 U153 ( .A1(\mem[6][1] ), .A2(n459), .ZN(n689) );
  OAI21_X1 U154 ( .B1(n487), .B2(n459), .A(n688), .ZN(n527) );
  NAND2_X1 U155 ( .A1(\mem[6][2] ), .A2(n691), .ZN(n688) );
  OAI21_X1 U156 ( .B1(n486), .B2(n691), .A(n687), .ZN(n526) );
  NAND2_X1 U157 ( .A1(\mem[6][3] ), .A2(n459), .ZN(n687) );
  OAI21_X1 U158 ( .B1(n485), .B2(n691), .A(n686), .ZN(n525) );
  NAND2_X1 U159 ( .A1(\mem[6][4] ), .A2(n691), .ZN(n686) );
  OAI21_X1 U160 ( .B1(n484), .B2(n691), .A(n685), .ZN(n524) );
  NAND2_X1 U161 ( .A1(\mem[6][5] ), .A2(n691), .ZN(n685) );
  OAI21_X1 U162 ( .B1(n483), .B2(n691), .A(n684), .ZN(n523) );
  NAND2_X1 U163 ( .A1(\mem[6][6] ), .A2(n691), .ZN(n684) );
  OAI21_X1 U164 ( .B1(n482), .B2(n691), .A(n683), .ZN(n522) );
  NAND2_X1 U165 ( .A1(\mem[6][7] ), .A2(n691), .ZN(n683) );
  OAI21_X1 U166 ( .B1(n481), .B2(n691), .A(n682), .ZN(n521) );
  NAND2_X1 U167 ( .A1(\mem[6][8] ), .A2(n691), .ZN(n682) );
  OAI21_X1 U168 ( .B1(n480), .B2(n459), .A(n681), .ZN(n520) );
  NAND2_X1 U169 ( .A1(\mem[6][9] ), .A2(n691), .ZN(n681) );
  OAI21_X1 U170 ( .B1(n479), .B2(n691), .A(n680), .ZN(n519) );
  NAND2_X1 U171 ( .A1(\mem[6][10] ), .A2(n691), .ZN(n680) );
  OAI21_X1 U172 ( .B1(n478), .B2(n691), .A(n679), .ZN(n518) );
  NAND2_X1 U173 ( .A1(\mem[6][11] ), .A2(n691), .ZN(n679) );
  OAI21_X1 U174 ( .B1(n477), .B2(n459), .A(n678), .ZN(n517) );
  NAND2_X1 U175 ( .A1(\mem[6][12] ), .A2(n459), .ZN(n678) );
  OAI21_X1 U176 ( .B1(n476), .B2(n459), .A(n677), .ZN(n516) );
  NAND2_X1 U177 ( .A1(\mem[6][13] ), .A2(n459), .ZN(n677) );
  OAI21_X1 U178 ( .B1(n475), .B2(n459), .A(n676), .ZN(n515) );
  NAND2_X1 U179 ( .A1(\mem[6][14] ), .A2(n459), .ZN(n676) );
  OAI21_X1 U180 ( .B1(n474), .B2(n691), .A(n675), .ZN(n514) );
  NAND2_X1 U181 ( .A1(\mem[6][15] ), .A2(n459), .ZN(n675) );
  OAI21_X1 U182 ( .B1(n473), .B2(n691), .A(n674), .ZN(n513) );
  NAND2_X1 U183 ( .A1(\mem[6][16] ), .A2(n459), .ZN(n674) );
  OAI21_X1 U184 ( .B1(n472), .B2(n691), .A(n673), .ZN(n512) );
  NAND2_X1 U185 ( .A1(\mem[6][17] ), .A2(n459), .ZN(n673) );
  OAI21_X1 U186 ( .B1(n471), .B2(n459), .A(n672), .ZN(n511) );
  NAND2_X1 U187 ( .A1(\mem[6][18] ), .A2(n459), .ZN(n672) );
  OAI21_X1 U188 ( .B1(n470), .B2(n459), .A(n671), .ZN(n510) );
  NAND2_X1 U189 ( .A1(\mem[6][19] ), .A2(n459), .ZN(n671) );
  OAI21_X1 U190 ( .B1(n489), .B2(n670), .A(n669), .ZN(n509) );
  NAND2_X1 U191 ( .A1(\mem[7][0] ), .A2(n458), .ZN(n669) );
  OAI21_X1 U192 ( .B1(n488), .B2(n670), .A(n668), .ZN(n508) );
  NAND2_X1 U193 ( .A1(\mem[7][1] ), .A2(n458), .ZN(n668) );
  OAI21_X1 U194 ( .B1(n487), .B2(n670), .A(n667), .ZN(n507) );
  NAND2_X1 U195 ( .A1(\mem[7][2] ), .A2(n458), .ZN(n667) );
  OAI21_X1 U196 ( .B1(n486), .B2(n670), .A(n666), .ZN(n506) );
  NAND2_X1 U197 ( .A1(\mem[7][3] ), .A2(n458), .ZN(n666) );
  OAI21_X1 U198 ( .B1(n485), .B2(n458), .A(n665), .ZN(n505) );
  NAND2_X1 U199 ( .A1(\mem[7][4] ), .A2(n458), .ZN(n665) );
  OAI21_X1 U200 ( .B1(n484), .B2(n670), .A(n664), .ZN(n504) );
  NAND2_X1 U201 ( .A1(\mem[7][5] ), .A2(n458), .ZN(n664) );
  OAI21_X1 U202 ( .B1(n483), .B2(n670), .A(n663), .ZN(n503) );
  NAND2_X1 U203 ( .A1(\mem[7][6] ), .A2(n458), .ZN(n663) );
  OAI21_X1 U204 ( .B1(n482), .B2(n670), .A(n662), .ZN(n502) );
  NAND2_X1 U205 ( .A1(\mem[7][7] ), .A2(n458), .ZN(n662) );
  OAI21_X1 U206 ( .B1(n481), .B2(n670), .A(n661), .ZN(n501) );
  NAND2_X1 U207 ( .A1(\mem[7][8] ), .A2(n458), .ZN(n661) );
  OAI21_X1 U208 ( .B1(n480), .B2(n670), .A(n660), .ZN(n500) );
  NAND2_X1 U209 ( .A1(\mem[7][9] ), .A2(n458), .ZN(n660) );
  OAI21_X1 U210 ( .B1(n479), .B2(n670), .A(n659), .ZN(n499) );
  NAND2_X1 U211 ( .A1(\mem[7][10] ), .A2(n458), .ZN(n659) );
  OAI21_X1 U212 ( .B1(n478), .B2(n670), .A(n658), .ZN(n498) );
  NAND2_X1 U213 ( .A1(\mem[7][11] ), .A2(n458), .ZN(n658) );
  OAI21_X1 U214 ( .B1(n477), .B2(n670), .A(n657), .ZN(n497) );
  NAND2_X1 U215 ( .A1(\mem[7][12] ), .A2(n670), .ZN(n657) );
  OAI21_X1 U216 ( .B1(n476), .B2(n458), .A(n656), .ZN(n496) );
  NAND2_X1 U217 ( .A1(\mem[7][13] ), .A2(n670), .ZN(n656) );
  OAI21_X1 U218 ( .B1(n475), .B2(n458), .A(n655), .ZN(n495) );
  NAND2_X1 U219 ( .A1(\mem[7][14] ), .A2(n670), .ZN(n655) );
  OAI21_X1 U220 ( .B1(n474), .B2(n670), .A(n654), .ZN(n494) );
  NAND2_X1 U221 ( .A1(\mem[7][15] ), .A2(n670), .ZN(n654) );
  OAI21_X1 U222 ( .B1(n473), .B2(n670), .A(n653), .ZN(n493) );
  NAND2_X1 U223 ( .A1(\mem[7][16] ), .A2(n670), .ZN(n653) );
  OAI21_X1 U224 ( .B1(n472), .B2(n670), .A(n652), .ZN(n492) );
  NAND2_X1 U225 ( .A1(\mem[7][17] ), .A2(n670), .ZN(n652) );
  OAI21_X1 U226 ( .B1(n471), .B2(n670), .A(n651), .ZN(n491) );
  NAND2_X1 U227 ( .A1(\mem[7][18] ), .A2(n670), .ZN(n651) );
  OAI21_X1 U228 ( .B1(n470), .B2(n670), .A(n650), .ZN(n490) );
  NAND2_X1 U229 ( .A1(\mem[7][19] ), .A2(n458), .ZN(n650) );
  NAND2_X1 U230 ( .A1(wr_en), .A2(n469), .ZN(n735) );
  INV_X1 U231 ( .A(addr[3]), .ZN(n469) );
  OAI21_X1 U232 ( .B1(n820), .B2(n489), .A(n819), .ZN(n649) );
  NAND2_X1 U233 ( .A1(\mem[0][0] ), .A2(n820), .ZN(n819) );
  OAI21_X1 U234 ( .B1(n465), .B2(n488), .A(n818), .ZN(n648) );
  NAND2_X1 U235 ( .A1(\mem[0][1] ), .A2(n820), .ZN(n818) );
  OAI21_X1 U236 ( .B1(n465), .B2(n487), .A(n817), .ZN(n647) );
  NAND2_X1 U237 ( .A1(\mem[0][2] ), .A2(n820), .ZN(n817) );
  OAI21_X1 U238 ( .B1(n465), .B2(n486), .A(n816), .ZN(n646) );
  NAND2_X1 U239 ( .A1(\mem[0][3] ), .A2(n820), .ZN(n816) );
  OAI21_X1 U240 ( .B1(n465), .B2(n485), .A(n815), .ZN(n645) );
  NAND2_X1 U241 ( .A1(\mem[0][4] ), .A2(n820), .ZN(n815) );
  OAI21_X1 U242 ( .B1(n465), .B2(n484), .A(n814), .ZN(n644) );
  NAND2_X1 U243 ( .A1(\mem[0][5] ), .A2(n820), .ZN(n814) );
  OAI21_X1 U244 ( .B1(n465), .B2(n483), .A(n813), .ZN(n643) );
  NAND2_X1 U245 ( .A1(\mem[0][6] ), .A2(n820), .ZN(n813) );
  OAI21_X1 U246 ( .B1(n465), .B2(n482), .A(n812), .ZN(n642) );
  NAND2_X1 U247 ( .A1(\mem[0][7] ), .A2(n820), .ZN(n812) );
  OAI21_X1 U248 ( .B1(n465), .B2(n481), .A(n811), .ZN(n641) );
  NAND2_X1 U249 ( .A1(\mem[0][8] ), .A2(n820), .ZN(n811) );
  OAI21_X1 U250 ( .B1(n820), .B2(n480), .A(n810), .ZN(n640) );
  NAND2_X1 U251 ( .A1(\mem[0][9] ), .A2(n820), .ZN(n810) );
  OAI21_X1 U252 ( .B1(n465), .B2(n479), .A(n809), .ZN(n639) );
  NAND2_X1 U253 ( .A1(\mem[0][10] ), .A2(n820), .ZN(n809) );
  OAI21_X1 U254 ( .B1(n465), .B2(n478), .A(n808), .ZN(n638) );
  NAND2_X1 U255 ( .A1(\mem[0][11] ), .A2(n820), .ZN(n808) );
  OAI21_X1 U256 ( .B1(n489), .B2(n798), .A(n797), .ZN(n629) );
  NAND2_X1 U257 ( .A1(\mem[1][0] ), .A2(n464), .ZN(n797) );
  OAI21_X1 U258 ( .B1(n488), .B2(n798), .A(n796), .ZN(n628) );
  NAND2_X1 U259 ( .A1(\mem[1][1] ), .A2(n464), .ZN(n796) );
  OAI21_X1 U260 ( .B1(n487), .B2(n798), .A(n795), .ZN(n627) );
  NAND2_X1 U261 ( .A1(\mem[1][2] ), .A2(n464), .ZN(n795) );
  OAI21_X1 U262 ( .B1(n486), .B2(n798), .A(n794), .ZN(n626) );
  NAND2_X1 U263 ( .A1(\mem[1][3] ), .A2(n464), .ZN(n794) );
  OAI21_X1 U264 ( .B1(n485), .B2(n798), .A(n793), .ZN(n625) );
  NAND2_X1 U265 ( .A1(\mem[1][4] ), .A2(n464), .ZN(n793) );
  OAI21_X1 U266 ( .B1(n484), .B2(n798), .A(n792), .ZN(n624) );
  NAND2_X1 U267 ( .A1(\mem[1][5] ), .A2(n464), .ZN(n792) );
  OAI21_X1 U268 ( .B1(n483), .B2(n798), .A(n791), .ZN(n623) );
  NAND2_X1 U269 ( .A1(\mem[1][6] ), .A2(n464), .ZN(n791) );
  OAI21_X1 U270 ( .B1(n482), .B2(n798), .A(n790), .ZN(n622) );
  NAND2_X1 U271 ( .A1(\mem[1][7] ), .A2(n464), .ZN(n790) );
  OAI21_X1 U272 ( .B1(n481), .B2(n798), .A(n789), .ZN(n621) );
  NAND2_X1 U273 ( .A1(\mem[1][8] ), .A2(n464), .ZN(n789) );
  OAI21_X1 U274 ( .B1(n480), .B2(n464), .A(n788), .ZN(n620) );
  NAND2_X1 U275 ( .A1(\mem[1][9] ), .A2(n464), .ZN(n788) );
  OAI21_X1 U276 ( .B1(n479), .B2(n798), .A(n787), .ZN(n619) );
  NAND2_X1 U277 ( .A1(\mem[1][10] ), .A2(n464), .ZN(n787) );
  OAI21_X1 U278 ( .B1(n478), .B2(n798), .A(n786), .ZN(n618) );
  NAND2_X1 U279 ( .A1(\mem[1][11] ), .A2(n464), .ZN(n786) );
  OAI21_X1 U280 ( .B1(n489), .B2(n777), .A(n776), .ZN(n609) );
  NAND2_X1 U281 ( .A1(\mem[2][0] ), .A2(n463), .ZN(n776) );
  OAI21_X1 U282 ( .B1(n488), .B2(n777), .A(n775), .ZN(n608) );
  NAND2_X1 U283 ( .A1(\mem[2][1] ), .A2(n463), .ZN(n775) );
  OAI21_X1 U284 ( .B1(n487), .B2(n777), .A(n774), .ZN(n607) );
  NAND2_X1 U285 ( .A1(\mem[2][2] ), .A2(n463), .ZN(n774) );
  OAI21_X1 U286 ( .B1(n486), .B2(n777), .A(n773), .ZN(n606) );
  NAND2_X1 U287 ( .A1(\mem[2][3] ), .A2(n463), .ZN(n773) );
  OAI21_X1 U288 ( .B1(n485), .B2(n777), .A(n772), .ZN(n605) );
  NAND2_X1 U289 ( .A1(\mem[2][4] ), .A2(n463), .ZN(n772) );
  OAI21_X1 U290 ( .B1(n484), .B2(n777), .A(n771), .ZN(n604) );
  NAND2_X1 U291 ( .A1(\mem[2][5] ), .A2(n463), .ZN(n771) );
  OAI21_X1 U292 ( .B1(n483), .B2(n777), .A(n770), .ZN(n603) );
  NAND2_X1 U293 ( .A1(\mem[2][6] ), .A2(n463), .ZN(n770) );
  OAI21_X1 U294 ( .B1(n482), .B2(n777), .A(n769), .ZN(n602) );
  NAND2_X1 U295 ( .A1(\mem[2][7] ), .A2(n463), .ZN(n769) );
  OAI21_X1 U296 ( .B1(n481), .B2(n777), .A(n768), .ZN(n601) );
  NAND2_X1 U297 ( .A1(\mem[2][8] ), .A2(n463), .ZN(n768) );
  OAI21_X1 U298 ( .B1(n480), .B2(n463), .A(n767), .ZN(n600) );
  NAND2_X1 U299 ( .A1(\mem[2][9] ), .A2(n463), .ZN(n767) );
  OAI21_X1 U300 ( .B1(n479), .B2(n777), .A(n766), .ZN(n599) );
  NAND2_X1 U301 ( .A1(\mem[2][10] ), .A2(n463), .ZN(n766) );
  OAI21_X1 U302 ( .B1(n478), .B2(n777), .A(n765), .ZN(n598) );
  NAND2_X1 U303 ( .A1(\mem[2][11] ), .A2(n463), .ZN(n765) );
  OAI21_X1 U304 ( .B1(n489), .B2(n756), .A(n755), .ZN(n589) );
  NAND2_X1 U305 ( .A1(\mem[3][0] ), .A2(n756), .ZN(n755) );
  OAI21_X1 U306 ( .B1(n488), .B2(n756), .A(n754), .ZN(n588) );
  NAND2_X1 U307 ( .A1(\mem[3][1] ), .A2(n756), .ZN(n754) );
  OAI21_X1 U308 ( .B1(n487), .B2(n756), .A(n753), .ZN(n587) );
  NAND2_X1 U309 ( .A1(\mem[3][2] ), .A2(n756), .ZN(n753) );
  OAI21_X1 U310 ( .B1(n486), .B2(n756), .A(n752), .ZN(n586) );
  NAND2_X1 U311 ( .A1(\mem[3][3] ), .A2(n462), .ZN(n752) );
  OAI21_X1 U312 ( .B1(n485), .B2(n756), .A(n751), .ZN(n585) );
  NAND2_X1 U313 ( .A1(\mem[3][4] ), .A2(n462), .ZN(n751) );
  OAI21_X1 U314 ( .B1(n484), .B2(n756), .A(n750), .ZN(n584) );
  NAND2_X1 U315 ( .A1(\mem[3][5] ), .A2(n462), .ZN(n750) );
  OAI21_X1 U316 ( .B1(n483), .B2(n756), .A(n749), .ZN(n583) );
  NAND2_X1 U317 ( .A1(\mem[3][6] ), .A2(n756), .ZN(n749) );
  OAI21_X1 U318 ( .B1(n482), .B2(n756), .A(n748), .ZN(n582) );
  NAND2_X1 U319 ( .A1(\mem[3][7] ), .A2(n756), .ZN(n748) );
  OAI21_X1 U320 ( .B1(n481), .B2(n756), .A(n747), .ZN(n581) );
  NAND2_X1 U321 ( .A1(\mem[3][8] ), .A2(n756), .ZN(n747) );
  OAI21_X1 U322 ( .B1(n480), .B2(n462), .A(n746), .ZN(n580) );
  NAND2_X1 U323 ( .A1(\mem[3][9] ), .A2(n462), .ZN(n746) );
  OAI21_X1 U324 ( .B1(n479), .B2(n756), .A(n745), .ZN(n579) );
  NAND2_X1 U325 ( .A1(\mem[3][10] ), .A2(n756), .ZN(n745) );
  OAI21_X1 U326 ( .B1(n478), .B2(n756), .A(n744), .ZN(n578) );
  NAND2_X1 U327 ( .A1(\mem[3][11] ), .A2(n756), .ZN(n744) );
  OAI21_X1 U328 ( .B1(n820), .B2(n477), .A(n807), .ZN(n637) );
  NAND2_X1 U329 ( .A1(\mem[0][12] ), .A2(n820), .ZN(n807) );
  OAI21_X1 U330 ( .B1(n820), .B2(n476), .A(n806), .ZN(n636) );
  NAND2_X1 U331 ( .A1(\mem[0][13] ), .A2(n820), .ZN(n806) );
  OAI21_X1 U332 ( .B1(n465), .B2(n475), .A(n805), .ZN(n635) );
  NAND2_X1 U333 ( .A1(\mem[0][14] ), .A2(n820), .ZN(n805) );
  OAI21_X1 U334 ( .B1(n465), .B2(n474), .A(n804), .ZN(n634) );
  NAND2_X1 U335 ( .A1(\mem[0][15] ), .A2(n820), .ZN(n804) );
  OAI21_X1 U336 ( .B1(n465), .B2(n473), .A(n803), .ZN(n633) );
  NAND2_X1 U337 ( .A1(\mem[0][16] ), .A2(n820), .ZN(n803) );
  OAI21_X1 U338 ( .B1(n465), .B2(n472), .A(n802), .ZN(n632) );
  NAND2_X1 U339 ( .A1(\mem[0][17] ), .A2(n820), .ZN(n802) );
  OAI21_X1 U340 ( .B1(n465), .B2(n471), .A(n801), .ZN(n631) );
  NAND2_X1 U341 ( .A1(\mem[0][18] ), .A2(n820), .ZN(n801) );
  OAI21_X1 U342 ( .B1(n465), .B2(n470), .A(n800), .ZN(n630) );
  NAND2_X1 U343 ( .A1(\mem[0][19] ), .A2(n820), .ZN(n800) );
  INV_X1 U344 ( .A(data_in[0]), .ZN(n489) );
  INV_X1 U345 ( .A(data_in[1]), .ZN(n488) );
  INV_X1 U346 ( .A(data_in[2]), .ZN(n487) );
  INV_X1 U347 ( .A(data_in[3]), .ZN(n486) );
  INV_X1 U348 ( .A(data_in[4]), .ZN(n485) );
  INV_X1 U349 ( .A(data_in[5]), .ZN(n484) );
  INV_X1 U358 ( .A(data_in[6]), .ZN(n483) );
  INV_X1 U359 ( .A(data_in[7]), .ZN(n482) );
  INV_X1 U360 ( .A(data_in[8]), .ZN(n481) );
  INV_X1 U361 ( .A(data_in[9]), .ZN(n480) );
  INV_X1 U362 ( .A(data_in[10]), .ZN(n479) );
  INV_X1 U363 ( .A(data_in[11]), .ZN(n478) );
  INV_X1 U364 ( .A(data_in[12]), .ZN(n477) );
  INV_X1 U365 ( .A(data_in[13]), .ZN(n476) );
  INV_X1 U366 ( .A(data_in[14]), .ZN(n475) );
  INV_X1 U367 ( .A(data_in[15]), .ZN(n474) );
  INV_X1 U368 ( .A(data_in[16]), .ZN(n473) );
  INV_X1 U369 ( .A(data_in[17]), .ZN(n472) );
  INV_X1 U370 ( .A(data_in[18]), .ZN(n471) );
  INV_X1 U371 ( .A(data_in[19]), .ZN(n470) );
  MUX2_X1 U372 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n457), .Z(n1) );
  MUX2_X1 U373 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n454), .Z(n2) );
  MUX2_X1 U374 ( .A(n2), .B(n1), .S(n452), .Z(n3) );
  MUX2_X1 U375 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n455), .Z(n4) );
  MUX2_X1 U376 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n455), .Z(n5) );
  MUX2_X1 U377 ( .A(n5), .B(n4), .S(n452), .Z(n6) );
  MUX2_X1 U378 ( .A(n6), .B(n3), .S(N12), .Z(N32) );
  MUX2_X1 U379 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n457), .Z(n7) );
  MUX2_X1 U380 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n455), .Z(n8) );
  MUX2_X1 U381 ( .A(n8), .B(n7), .S(n452), .Z(n9) );
  MUX2_X1 U382 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n456), .Z(n10) );
  MUX2_X1 U383 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n455), .Z(n11) );
  MUX2_X1 U384 ( .A(n11), .B(n10), .S(n452), .Z(n12) );
  MUX2_X1 U385 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n454), .Z(n13) );
  MUX2_X1 U386 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n455), .Z(n14) );
  MUX2_X1 U387 ( .A(n14), .B(n13), .S(n453), .Z(n15) );
  MUX2_X1 U388 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n455), .Z(n16) );
  MUX2_X1 U389 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n456), .Z(n17) );
  MUX2_X1 U390 ( .A(n17), .B(n16), .S(n453), .Z(n18) );
  MUX2_X1 U391 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n454), .Z(n19) );
  MUX2_X1 U392 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n456), .Z(n20) );
  MUX2_X1 U393 ( .A(n20), .B(n19), .S(n453), .Z(n21) );
  MUX2_X1 U394 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n454), .Z(n22) );
  MUX2_X1 U395 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n457), .Z(n23) );
  MUX2_X1 U396 ( .A(n23), .B(n22), .S(n453), .Z(n24) );
  MUX2_X1 U397 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n454), .Z(n356) );
  MUX2_X1 U398 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n456), .Z(n357) );
  MUX2_X1 U399 ( .A(n357), .B(n356), .S(n453), .Z(n358) );
  MUX2_X1 U400 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n455), .Z(n359) );
  MUX2_X1 U401 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n457), .Z(n360) );
  MUX2_X1 U402 ( .A(n360), .B(n359), .S(n453), .Z(n361) );
  MUX2_X1 U403 ( .A(n361), .B(n358), .S(N12), .Z(N28) );
  MUX2_X1 U404 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n454), .Z(n362) );
  MUX2_X1 U405 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n454), .Z(n363) );
  MUX2_X1 U406 ( .A(n363), .B(n362), .S(n453), .Z(n364) );
  MUX2_X1 U407 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n454), .Z(n365) );
  MUX2_X1 U408 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n454), .Z(n366) );
  MUX2_X1 U409 ( .A(n366), .B(n365), .S(n453), .Z(n367) );
  MUX2_X1 U410 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n454), .Z(n368) );
  MUX2_X1 U411 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n454), .Z(n369) );
  MUX2_X1 U412 ( .A(n369), .B(n368), .S(n453), .Z(n370) );
  MUX2_X1 U413 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n454), .Z(n371) );
  MUX2_X1 U414 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n454), .Z(n372) );
  MUX2_X1 U415 ( .A(n372), .B(n371), .S(n453), .Z(n373) );
  MUX2_X1 U416 ( .A(n373), .B(n370), .S(N12), .Z(N26) );
  MUX2_X1 U417 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n454), .Z(n374) );
  MUX2_X1 U418 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n454), .Z(n375) );
  MUX2_X1 U419 ( .A(n375), .B(n374), .S(n453), .Z(n376) );
  MUX2_X1 U420 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n454), .Z(n377) );
  MUX2_X1 U421 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n454), .Z(n378) );
  MUX2_X1 U422 ( .A(n378), .B(n377), .S(n453), .Z(n379) );
  MUX2_X1 U423 ( .A(n379), .B(n376), .S(N12), .Z(N25) );
  MUX2_X1 U424 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n455), .Z(n380) );
  MUX2_X1 U425 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n455), .Z(n381) );
  MUX2_X1 U426 ( .A(n381), .B(n380), .S(n453), .Z(n382) );
  MUX2_X1 U427 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n455), .Z(n383) );
  MUX2_X1 U428 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n455), .Z(n384) );
  MUX2_X1 U429 ( .A(n384), .B(n383), .S(N11), .Z(n385) );
  MUX2_X1 U430 ( .A(n385), .B(n382), .S(N12), .Z(N24) );
  MUX2_X1 U431 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n455), .Z(n386) );
  MUX2_X1 U432 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n455), .Z(n387) );
  MUX2_X1 U433 ( .A(n387), .B(n386), .S(n453), .Z(n388) );
  MUX2_X1 U434 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n455), .Z(n389) );
  MUX2_X1 U435 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n455), .Z(n390) );
  MUX2_X1 U436 ( .A(n390), .B(n389), .S(N11), .Z(n391) );
  MUX2_X1 U437 ( .A(n391), .B(n388), .S(N12), .Z(N23) );
  MUX2_X1 U438 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n455), .Z(n392) );
  MUX2_X1 U439 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n455), .Z(n393) );
  MUX2_X1 U440 ( .A(n393), .B(n392), .S(n453), .Z(n394) );
  MUX2_X1 U441 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n455), .Z(n395) );
  MUX2_X1 U442 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n455), .Z(n396) );
  MUX2_X1 U443 ( .A(n396), .B(n395), .S(N11), .Z(n397) );
  MUX2_X1 U444 ( .A(n397), .B(n394), .S(N12), .Z(N22) );
  MUX2_X1 U445 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n456), .Z(n398) );
  MUX2_X1 U446 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n456), .Z(n399) );
  MUX2_X1 U447 ( .A(n399), .B(n398), .S(n453), .Z(n400) );
  MUX2_X1 U448 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n456), .Z(n401) );
  MUX2_X1 U449 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n456), .Z(n402) );
  MUX2_X1 U450 ( .A(n402), .B(n401), .S(N11), .Z(n403) );
  MUX2_X1 U451 ( .A(n403), .B(n400), .S(N12), .Z(N21) );
  MUX2_X1 U452 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n456), .Z(n404) );
  MUX2_X1 U453 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n456), .Z(n405) );
  MUX2_X1 U454 ( .A(n405), .B(n404), .S(n453), .Z(n406) );
  MUX2_X1 U455 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n456), .Z(n407) );
  MUX2_X1 U456 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n456), .Z(n408) );
  MUX2_X1 U457 ( .A(n408), .B(n407), .S(N11), .Z(n409) );
  MUX2_X1 U458 ( .A(n409), .B(n406), .S(N12), .Z(N20) );
  MUX2_X1 U459 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n456), .Z(n410) );
  MUX2_X1 U460 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n456), .Z(n411) );
  MUX2_X1 U461 ( .A(n411), .B(n410), .S(n453), .Z(n412) );
  MUX2_X1 U462 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n456), .Z(n413) );
  MUX2_X1 U463 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n456), .Z(n414) );
  MUX2_X1 U464 ( .A(n414), .B(n413), .S(N11), .Z(n415) );
  MUX2_X1 U465 ( .A(n415), .B(n412), .S(N12), .Z(N19) );
  MUX2_X1 U466 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n457), .Z(n416) );
  MUX2_X1 U467 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n457), .Z(n417) );
  MUX2_X1 U468 ( .A(n417), .B(n416), .S(n452), .Z(n418) );
  MUX2_X1 U469 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n457), .Z(n419) );
  MUX2_X1 U470 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n457), .Z(n420) );
  MUX2_X1 U471 ( .A(n420), .B(n419), .S(n452), .Z(n421) );
  MUX2_X1 U472 ( .A(n421), .B(n418), .S(N12), .Z(N18) );
  MUX2_X1 U473 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n457), .Z(n422) );
  MUX2_X1 U474 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n457), .Z(n423) );
  MUX2_X1 U475 ( .A(n423), .B(n422), .S(n452), .Z(n424) );
  MUX2_X1 U476 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n457), .Z(n425) );
  MUX2_X1 U477 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n457), .Z(n426) );
  MUX2_X1 U478 ( .A(n426), .B(n425), .S(n452), .Z(n427) );
  MUX2_X1 U479 ( .A(n427), .B(n424), .S(N12), .Z(N17) );
  MUX2_X1 U480 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n457), .Z(n428) );
  MUX2_X1 U481 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n457), .Z(n429) );
  MUX2_X1 U482 ( .A(n429), .B(n428), .S(n452), .Z(n430) );
  MUX2_X1 U483 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n457), .Z(n431) );
  MUX2_X1 U484 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n457), .Z(n432) );
  MUX2_X1 U485 ( .A(n432), .B(n431), .S(n452), .Z(n433) );
  MUX2_X1 U486 ( .A(n433), .B(n430), .S(N12), .Z(N16) );
  MUX2_X1 U487 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n457), .Z(n434) );
  MUX2_X1 U488 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n456), .Z(n435) );
  MUX2_X1 U489 ( .A(n435), .B(n434), .S(n453), .Z(n436) );
  MUX2_X1 U490 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n454), .Z(n437) );
  MUX2_X1 U491 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n456), .Z(n438) );
  MUX2_X1 U492 ( .A(n438), .B(n437), .S(n453), .Z(n439) );
  MUX2_X1 U493 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n455), .Z(n440) );
  MUX2_X1 U494 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n456), .Z(n441) );
  MUX2_X1 U495 ( .A(n441), .B(n440), .S(n452), .Z(n442) );
  MUX2_X1 U496 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n457), .Z(n443) );
  MUX2_X1 U497 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n457), .Z(n444) );
  MUX2_X1 U498 ( .A(n444), .B(n443), .S(n453), .Z(n445) );
  MUX2_X1 U499 ( .A(n445), .B(n442), .S(N12), .Z(N14) );
  MUX2_X1 U500 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n456), .Z(n446) );
  MUX2_X1 U501 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n457), .Z(n447) );
  MUX2_X1 U502 ( .A(n447), .B(n446), .S(n452), .Z(n448) );
  MUX2_X1 U503 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n454), .Z(n449) );
  MUX2_X1 U504 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n454), .Z(n450) );
  MUX2_X1 U505 ( .A(n450), .B(n449), .S(n453), .Z(n451) );
  MUX2_X1 U506 ( .A(n451), .B(n448), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE4_5 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N13, N14, N16, N17, N18, N19, N20, N22, N23, N24, N26,
         N27, N28, N30, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[19]  ( .D(N13), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[15]  ( .D(N17), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N19), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N20), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N23), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N27), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N30), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N32), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n490), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n491), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n492), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n493), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n494), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n495), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n496), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n497), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n498), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n499), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n500), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n501), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n502), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n503), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n504), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n505), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n506), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n507), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n508), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n509), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n510), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n511), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n512), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n513), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n514), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n515), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n516), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n517), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n518), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n519), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n520), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n521), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n522), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n523), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n524), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n525), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n526), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n527), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n528), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n529), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n530), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n531), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n532), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n533), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n534), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n535), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n536), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n537), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n538), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n539), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n540), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n541), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n542), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n543), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n544), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n545), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n546), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n547), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n548), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n549), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n550), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n551), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n552), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n553), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n554), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n555), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n556), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n557), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n558), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n559), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n560), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n561), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n562), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n563), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n564), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n565), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n566), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n567), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n568), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n569), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n570), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n571), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n572), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n573), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n574), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n575), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n576), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n577), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n578), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n579), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n580), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n581), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n582), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n583), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n584), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n585), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n586), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n587), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n588), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n589), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n590), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n591), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n592), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n593), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n594), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n595), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n596), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n597), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n598), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n599), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n600), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n601), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n602), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n603), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n604), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n605), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n606), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n607), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n608), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n609), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n610), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n611), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n612), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n613), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n614), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n615), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n616), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n617), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n618), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n619), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n620), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n621), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n622), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n623), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n624), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n625), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n626), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n627), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n628), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n629), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n630), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n631), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n632), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n633), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n634), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n635), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n636), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n637), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n638), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n639), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n640), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n641), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n642), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n643), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n644), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n645), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n646), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n647), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n648), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n649), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U350 ( .A1(n466), .A2(n467), .A3(n799), .ZN(n820) );
  NAND3_X1 U351 ( .A1(n799), .A2(n467), .A3(N10), .ZN(n798) );
  NAND3_X1 U352 ( .A1(n799), .A2(n466), .A3(N11), .ZN(n777) );
  NAND3_X1 U353 ( .A1(N10), .A2(n799), .A3(N11), .ZN(n756) );
  NAND3_X1 U354 ( .A1(n466), .A2(n467), .A3(n713), .ZN(n734) );
  NAND3_X1 U355 ( .A1(N10), .A2(n467), .A3(n713), .ZN(n712) );
  NAND3_X1 U356 ( .A1(N11), .A2(n466), .A3(n713), .ZN(n691) );
  NAND3_X1 U357 ( .A1(N11), .A2(N10), .A3(n713), .ZN(n670) );
  SDFF_X1 \data_out_reg[17]  ( .D(n436), .SI(n439), .SE(n468), .CK(clk), .Q(
        data_out[17]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n376), .SI(n379), .SE(n468), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n400), .SI(n403), .SE(n468), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n9), .SI(n12), .SE(n468), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n21), .SI(n24), .SE(n468), .CK(clk), .Q(
        data_out[3]) );
  BUF_X1 U3 ( .A(n798), .Z(n464) );
  BUF_X1 U4 ( .A(n734), .Z(n461) );
  BUF_X1 U5 ( .A(n756), .Z(n462) );
  BUF_X1 U6 ( .A(n691), .Z(n459) );
  BUF_X1 U7 ( .A(n453), .Z(n452) );
  BUF_X1 U8 ( .A(N10), .Z(n455) );
  BUF_X1 U9 ( .A(N10), .Z(n456) );
  BUF_X1 U10 ( .A(N10), .Z(n457) );
  BUF_X1 U11 ( .A(N10), .Z(n454) );
  BUF_X1 U12 ( .A(n820), .Z(n465) );
  BUF_X1 U13 ( .A(n777), .Z(n463) );
  BUF_X1 U14 ( .A(n670), .Z(n458) );
  BUF_X1 U15 ( .A(n712), .Z(n460) );
  BUF_X1 U16 ( .A(N11), .Z(n453) );
  NOR2_X1 U17 ( .A1(n735), .A2(N12), .ZN(n799) );
  NOR2_X1 U18 ( .A1(n468), .A2(n735), .ZN(n713) );
  INV_X1 U19 ( .A(N12), .ZN(n468) );
  INV_X1 U20 ( .A(N11), .ZN(n467) );
  INV_X1 U21 ( .A(N10), .ZN(n466) );
  OAI21_X1 U22 ( .B1(n477), .B2(n464), .A(n785), .ZN(n617) );
  NAND2_X1 U23 ( .A1(\mem[1][12] ), .A2(n464), .ZN(n785) );
  OAI21_X1 U24 ( .B1(n476), .B2(n464), .A(n784), .ZN(n616) );
  NAND2_X1 U25 ( .A1(\mem[1][13] ), .A2(n464), .ZN(n784) );
  OAI21_X1 U26 ( .B1(n475), .B2(n464), .A(n783), .ZN(n615) );
  NAND2_X1 U27 ( .A1(\mem[1][14] ), .A2(n464), .ZN(n783) );
  OAI21_X1 U28 ( .B1(n474), .B2(n798), .A(n782), .ZN(n614) );
  NAND2_X1 U29 ( .A1(\mem[1][15] ), .A2(n464), .ZN(n782) );
  OAI21_X1 U30 ( .B1(n473), .B2(n798), .A(n781), .ZN(n613) );
  NAND2_X1 U31 ( .A1(\mem[1][16] ), .A2(n464), .ZN(n781) );
  OAI21_X1 U32 ( .B1(n472), .B2(n798), .A(n780), .ZN(n612) );
  NAND2_X1 U33 ( .A1(\mem[1][17] ), .A2(n464), .ZN(n780) );
  OAI21_X1 U34 ( .B1(n471), .B2(n798), .A(n779), .ZN(n611) );
  NAND2_X1 U35 ( .A1(\mem[1][18] ), .A2(n464), .ZN(n779) );
  OAI21_X1 U36 ( .B1(n470), .B2(n798), .A(n778), .ZN(n610) );
  NAND2_X1 U37 ( .A1(\mem[1][19] ), .A2(n464), .ZN(n778) );
  OAI21_X1 U38 ( .B1(n477), .B2(n777), .A(n764), .ZN(n597) );
  NAND2_X1 U39 ( .A1(\mem[2][12] ), .A2(n777), .ZN(n764) );
  OAI21_X1 U40 ( .B1(n476), .B2(n777), .A(n763), .ZN(n596) );
  NAND2_X1 U41 ( .A1(\mem[2][13] ), .A2(n777), .ZN(n763) );
  OAI21_X1 U42 ( .B1(n475), .B2(n777), .A(n762), .ZN(n595) );
  NAND2_X1 U43 ( .A1(\mem[2][14] ), .A2(n777), .ZN(n762) );
  OAI21_X1 U44 ( .B1(n474), .B2(n463), .A(n761), .ZN(n594) );
  NAND2_X1 U45 ( .A1(\mem[2][15] ), .A2(n777), .ZN(n761) );
  OAI21_X1 U46 ( .B1(n473), .B2(n777), .A(n760), .ZN(n593) );
  NAND2_X1 U47 ( .A1(\mem[2][16] ), .A2(n463), .ZN(n760) );
  OAI21_X1 U48 ( .B1(n472), .B2(n777), .A(n759), .ZN(n592) );
  NAND2_X1 U49 ( .A1(\mem[2][17] ), .A2(n777), .ZN(n759) );
  OAI21_X1 U50 ( .B1(n471), .B2(n777), .A(n758), .ZN(n591) );
  NAND2_X1 U51 ( .A1(\mem[2][18] ), .A2(n777), .ZN(n758) );
  OAI21_X1 U52 ( .B1(n470), .B2(n777), .A(n757), .ZN(n590) );
  NAND2_X1 U53 ( .A1(\mem[2][19] ), .A2(n463), .ZN(n757) );
  OAI21_X1 U54 ( .B1(n477), .B2(n756), .A(n743), .ZN(n577) );
  NAND2_X1 U55 ( .A1(\mem[3][12] ), .A2(n756), .ZN(n743) );
  OAI21_X1 U56 ( .B1(n476), .B2(n756), .A(n742), .ZN(n576) );
  NAND2_X1 U57 ( .A1(\mem[3][13] ), .A2(n756), .ZN(n742) );
  OAI21_X1 U58 ( .B1(n475), .B2(n462), .A(n741), .ZN(n575) );
  NAND2_X1 U59 ( .A1(\mem[3][14] ), .A2(n756), .ZN(n741) );
  OAI21_X1 U60 ( .B1(n474), .B2(n462), .A(n740), .ZN(n574) );
  NAND2_X1 U61 ( .A1(\mem[3][15] ), .A2(n756), .ZN(n740) );
  OAI21_X1 U62 ( .B1(n473), .B2(n462), .A(n739), .ZN(n573) );
  NAND2_X1 U63 ( .A1(\mem[3][16] ), .A2(n756), .ZN(n739) );
  OAI21_X1 U64 ( .B1(n472), .B2(n462), .A(n738), .ZN(n572) );
  NAND2_X1 U65 ( .A1(\mem[3][17] ), .A2(n756), .ZN(n738) );
  OAI21_X1 U66 ( .B1(n471), .B2(n462), .A(n737), .ZN(n571) );
  NAND2_X1 U67 ( .A1(\mem[3][18] ), .A2(n756), .ZN(n737) );
  OAI21_X1 U68 ( .B1(n470), .B2(n756), .A(n736), .ZN(n570) );
  NAND2_X1 U69 ( .A1(\mem[3][19] ), .A2(n756), .ZN(n736) );
  OAI21_X1 U70 ( .B1(n489), .B2(n461), .A(n733), .ZN(n569) );
  NAND2_X1 U71 ( .A1(\mem[4][0] ), .A2(n461), .ZN(n733) );
  OAI21_X1 U72 ( .B1(n488), .B2(n461), .A(n732), .ZN(n568) );
  NAND2_X1 U73 ( .A1(\mem[4][1] ), .A2(n461), .ZN(n732) );
  OAI21_X1 U74 ( .B1(n487), .B2(n461), .A(n731), .ZN(n567) );
  NAND2_X1 U75 ( .A1(\mem[4][2] ), .A2(n734), .ZN(n731) );
  OAI21_X1 U76 ( .B1(n486), .B2(n734), .A(n730), .ZN(n566) );
  NAND2_X1 U77 ( .A1(\mem[4][3] ), .A2(n461), .ZN(n730) );
  OAI21_X1 U78 ( .B1(n485), .B2(n734), .A(n729), .ZN(n565) );
  NAND2_X1 U79 ( .A1(\mem[4][4] ), .A2(n734), .ZN(n729) );
  OAI21_X1 U80 ( .B1(n484), .B2(n734), .A(n728), .ZN(n564) );
  NAND2_X1 U81 ( .A1(\mem[4][5] ), .A2(n734), .ZN(n728) );
  OAI21_X1 U82 ( .B1(n483), .B2(n734), .A(n727), .ZN(n563) );
  NAND2_X1 U83 ( .A1(\mem[4][6] ), .A2(n734), .ZN(n727) );
  OAI21_X1 U84 ( .B1(n482), .B2(n734), .A(n726), .ZN(n562) );
  NAND2_X1 U85 ( .A1(\mem[4][7] ), .A2(n734), .ZN(n726) );
  OAI21_X1 U86 ( .B1(n481), .B2(n734), .A(n725), .ZN(n561) );
  NAND2_X1 U87 ( .A1(\mem[4][8] ), .A2(n734), .ZN(n725) );
  OAI21_X1 U88 ( .B1(n480), .B2(n461), .A(n724), .ZN(n560) );
  NAND2_X1 U89 ( .A1(\mem[4][9] ), .A2(n734), .ZN(n724) );
  OAI21_X1 U90 ( .B1(n479), .B2(n734), .A(n723), .ZN(n559) );
  NAND2_X1 U91 ( .A1(\mem[4][10] ), .A2(n734), .ZN(n723) );
  OAI21_X1 U92 ( .B1(n478), .B2(n734), .A(n722), .ZN(n558) );
  NAND2_X1 U93 ( .A1(\mem[4][11] ), .A2(n734), .ZN(n722) );
  OAI21_X1 U94 ( .B1(n477), .B2(n461), .A(n721), .ZN(n557) );
  NAND2_X1 U95 ( .A1(\mem[4][12] ), .A2(n461), .ZN(n721) );
  OAI21_X1 U96 ( .B1(n476), .B2(n461), .A(n720), .ZN(n556) );
  NAND2_X1 U97 ( .A1(\mem[4][13] ), .A2(n461), .ZN(n720) );
  OAI21_X1 U98 ( .B1(n475), .B2(n461), .A(n719), .ZN(n555) );
  NAND2_X1 U99 ( .A1(\mem[4][14] ), .A2(n461), .ZN(n719) );
  OAI21_X1 U100 ( .B1(n474), .B2(n734), .A(n718), .ZN(n554) );
  NAND2_X1 U101 ( .A1(\mem[4][15] ), .A2(n461), .ZN(n718) );
  OAI21_X1 U102 ( .B1(n473), .B2(n734), .A(n717), .ZN(n553) );
  NAND2_X1 U103 ( .A1(\mem[4][16] ), .A2(n461), .ZN(n717) );
  OAI21_X1 U104 ( .B1(n472), .B2(n734), .A(n716), .ZN(n552) );
  NAND2_X1 U105 ( .A1(\mem[4][17] ), .A2(n461), .ZN(n716) );
  OAI21_X1 U106 ( .B1(n471), .B2(n461), .A(n715), .ZN(n551) );
  NAND2_X1 U107 ( .A1(\mem[4][18] ), .A2(n461), .ZN(n715) );
  OAI21_X1 U108 ( .B1(n470), .B2(n461), .A(n714), .ZN(n550) );
  NAND2_X1 U109 ( .A1(\mem[4][19] ), .A2(n461), .ZN(n714) );
  OAI21_X1 U110 ( .B1(n489), .B2(n712), .A(n711), .ZN(n549) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n460), .ZN(n711) );
  OAI21_X1 U112 ( .B1(n488), .B2(n712), .A(n710), .ZN(n548) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n460), .ZN(n710) );
  OAI21_X1 U114 ( .B1(n487), .B2(n712), .A(n709), .ZN(n547) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n460), .ZN(n709) );
  OAI21_X1 U116 ( .B1(n486), .B2(n712), .A(n708), .ZN(n546) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n460), .ZN(n708) );
  OAI21_X1 U118 ( .B1(n485), .B2(n460), .A(n707), .ZN(n545) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n460), .ZN(n707) );
  OAI21_X1 U120 ( .B1(n484), .B2(n712), .A(n706), .ZN(n544) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n460), .ZN(n706) );
  OAI21_X1 U122 ( .B1(n483), .B2(n712), .A(n705), .ZN(n543) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n460), .ZN(n705) );
  OAI21_X1 U124 ( .B1(n482), .B2(n712), .A(n704), .ZN(n542) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n460), .ZN(n704) );
  OAI21_X1 U126 ( .B1(n481), .B2(n712), .A(n703), .ZN(n541) );
  NAND2_X1 U127 ( .A1(\mem[5][8] ), .A2(n460), .ZN(n703) );
  OAI21_X1 U128 ( .B1(n480), .B2(n712), .A(n702), .ZN(n540) );
  NAND2_X1 U129 ( .A1(\mem[5][9] ), .A2(n460), .ZN(n702) );
  OAI21_X1 U130 ( .B1(n479), .B2(n712), .A(n701), .ZN(n539) );
  NAND2_X1 U131 ( .A1(\mem[5][10] ), .A2(n460), .ZN(n701) );
  OAI21_X1 U132 ( .B1(n478), .B2(n712), .A(n700), .ZN(n538) );
  NAND2_X1 U133 ( .A1(\mem[5][11] ), .A2(n460), .ZN(n700) );
  OAI21_X1 U134 ( .B1(n477), .B2(n712), .A(n699), .ZN(n537) );
  NAND2_X1 U135 ( .A1(\mem[5][12] ), .A2(n712), .ZN(n699) );
  OAI21_X1 U136 ( .B1(n476), .B2(n460), .A(n698), .ZN(n536) );
  NAND2_X1 U137 ( .A1(\mem[5][13] ), .A2(n712), .ZN(n698) );
  OAI21_X1 U138 ( .B1(n475), .B2(n460), .A(n697), .ZN(n535) );
  NAND2_X1 U139 ( .A1(\mem[5][14] ), .A2(n712), .ZN(n697) );
  OAI21_X1 U140 ( .B1(n474), .B2(n712), .A(n696), .ZN(n534) );
  NAND2_X1 U141 ( .A1(\mem[5][15] ), .A2(n712), .ZN(n696) );
  OAI21_X1 U142 ( .B1(n473), .B2(n712), .A(n695), .ZN(n533) );
  NAND2_X1 U143 ( .A1(\mem[5][16] ), .A2(n712), .ZN(n695) );
  OAI21_X1 U144 ( .B1(n472), .B2(n712), .A(n694), .ZN(n532) );
  NAND2_X1 U145 ( .A1(\mem[5][17] ), .A2(n712), .ZN(n694) );
  OAI21_X1 U146 ( .B1(n471), .B2(n712), .A(n693), .ZN(n531) );
  NAND2_X1 U147 ( .A1(\mem[5][18] ), .A2(n712), .ZN(n693) );
  OAI21_X1 U148 ( .B1(n470), .B2(n712), .A(n692), .ZN(n530) );
  NAND2_X1 U149 ( .A1(\mem[5][19] ), .A2(n460), .ZN(n692) );
  OAI21_X1 U150 ( .B1(n489), .B2(n691), .A(n690), .ZN(n529) );
  NAND2_X1 U151 ( .A1(\mem[6][0] ), .A2(n691), .ZN(n690) );
  OAI21_X1 U152 ( .B1(n488), .B2(n459), .A(n689), .ZN(n528) );
  NAND2_X1 U153 ( .A1(\mem[6][1] ), .A2(n691), .ZN(n689) );
  OAI21_X1 U154 ( .B1(n487), .B2(n459), .A(n688), .ZN(n527) );
  NAND2_X1 U155 ( .A1(\mem[6][2] ), .A2(n691), .ZN(n688) );
  OAI21_X1 U156 ( .B1(n486), .B2(n459), .A(n687), .ZN(n526) );
  NAND2_X1 U157 ( .A1(\mem[6][3] ), .A2(n691), .ZN(n687) );
  OAI21_X1 U158 ( .B1(n485), .B2(n459), .A(n686), .ZN(n525) );
  NAND2_X1 U159 ( .A1(\mem[6][4] ), .A2(n691), .ZN(n686) );
  OAI21_X1 U160 ( .B1(n484), .B2(n459), .A(n685), .ZN(n524) );
  NAND2_X1 U161 ( .A1(\mem[6][5] ), .A2(n691), .ZN(n685) );
  OAI21_X1 U162 ( .B1(n483), .B2(n459), .A(n684), .ZN(n523) );
  NAND2_X1 U163 ( .A1(\mem[6][6] ), .A2(n691), .ZN(n684) );
  OAI21_X1 U164 ( .B1(n482), .B2(n459), .A(n683), .ZN(n522) );
  NAND2_X1 U165 ( .A1(\mem[6][7] ), .A2(n691), .ZN(n683) );
  OAI21_X1 U166 ( .B1(n481), .B2(n459), .A(n682), .ZN(n521) );
  NAND2_X1 U167 ( .A1(\mem[6][8] ), .A2(n691), .ZN(n682) );
  OAI21_X1 U168 ( .B1(n480), .B2(n691), .A(n681), .ZN(n520) );
  NAND2_X1 U169 ( .A1(\mem[6][9] ), .A2(n691), .ZN(n681) );
  OAI21_X1 U170 ( .B1(n479), .B2(n459), .A(n680), .ZN(n519) );
  NAND2_X1 U171 ( .A1(\mem[6][10] ), .A2(n691), .ZN(n680) );
  OAI21_X1 U172 ( .B1(n478), .B2(n459), .A(n679), .ZN(n518) );
  NAND2_X1 U173 ( .A1(\mem[6][11] ), .A2(n691), .ZN(n679) );
  OAI21_X1 U174 ( .B1(n477), .B2(n691), .A(n678), .ZN(n517) );
  NAND2_X1 U175 ( .A1(\mem[6][12] ), .A2(n691), .ZN(n678) );
  OAI21_X1 U176 ( .B1(n476), .B2(n459), .A(n677), .ZN(n516) );
  NAND2_X1 U177 ( .A1(\mem[6][13] ), .A2(n691), .ZN(n677) );
  OAI21_X1 U178 ( .B1(n475), .B2(n691), .A(n676), .ZN(n515) );
  NAND2_X1 U179 ( .A1(\mem[6][14] ), .A2(n691), .ZN(n676) );
  OAI21_X1 U180 ( .B1(n474), .B2(n459), .A(n675), .ZN(n514) );
  NAND2_X1 U181 ( .A1(\mem[6][15] ), .A2(n691), .ZN(n675) );
  OAI21_X1 U182 ( .B1(n473), .B2(n459), .A(n674), .ZN(n513) );
  NAND2_X1 U183 ( .A1(\mem[6][16] ), .A2(n691), .ZN(n674) );
  OAI21_X1 U184 ( .B1(n472), .B2(n459), .A(n673), .ZN(n512) );
  NAND2_X1 U185 ( .A1(\mem[6][17] ), .A2(n691), .ZN(n673) );
  OAI21_X1 U186 ( .B1(n471), .B2(n459), .A(n672), .ZN(n511) );
  NAND2_X1 U187 ( .A1(\mem[6][18] ), .A2(n691), .ZN(n672) );
  OAI21_X1 U188 ( .B1(n470), .B2(n459), .A(n671), .ZN(n510) );
  NAND2_X1 U189 ( .A1(\mem[6][19] ), .A2(n691), .ZN(n671) );
  OAI21_X1 U190 ( .B1(n489), .B2(n670), .A(n669), .ZN(n509) );
  NAND2_X1 U191 ( .A1(\mem[7][0] ), .A2(n458), .ZN(n669) );
  OAI21_X1 U192 ( .B1(n488), .B2(n670), .A(n668), .ZN(n508) );
  NAND2_X1 U193 ( .A1(\mem[7][1] ), .A2(n458), .ZN(n668) );
  OAI21_X1 U194 ( .B1(n487), .B2(n670), .A(n667), .ZN(n507) );
  NAND2_X1 U195 ( .A1(\mem[7][2] ), .A2(n458), .ZN(n667) );
  OAI21_X1 U196 ( .B1(n486), .B2(n670), .A(n666), .ZN(n506) );
  NAND2_X1 U197 ( .A1(\mem[7][3] ), .A2(n458), .ZN(n666) );
  OAI21_X1 U198 ( .B1(n485), .B2(n458), .A(n665), .ZN(n505) );
  NAND2_X1 U199 ( .A1(\mem[7][4] ), .A2(n458), .ZN(n665) );
  OAI21_X1 U200 ( .B1(n484), .B2(n670), .A(n664), .ZN(n504) );
  NAND2_X1 U201 ( .A1(\mem[7][5] ), .A2(n458), .ZN(n664) );
  OAI21_X1 U202 ( .B1(n483), .B2(n670), .A(n663), .ZN(n503) );
  NAND2_X1 U203 ( .A1(\mem[7][6] ), .A2(n458), .ZN(n663) );
  OAI21_X1 U204 ( .B1(n482), .B2(n670), .A(n662), .ZN(n502) );
  NAND2_X1 U205 ( .A1(\mem[7][7] ), .A2(n458), .ZN(n662) );
  OAI21_X1 U206 ( .B1(n481), .B2(n670), .A(n661), .ZN(n501) );
  NAND2_X1 U207 ( .A1(\mem[7][8] ), .A2(n458), .ZN(n661) );
  OAI21_X1 U208 ( .B1(n480), .B2(n670), .A(n660), .ZN(n500) );
  NAND2_X1 U209 ( .A1(\mem[7][9] ), .A2(n458), .ZN(n660) );
  OAI21_X1 U210 ( .B1(n479), .B2(n670), .A(n659), .ZN(n499) );
  NAND2_X1 U211 ( .A1(\mem[7][10] ), .A2(n458), .ZN(n659) );
  OAI21_X1 U212 ( .B1(n478), .B2(n670), .A(n658), .ZN(n498) );
  NAND2_X1 U213 ( .A1(\mem[7][11] ), .A2(n458), .ZN(n658) );
  OAI21_X1 U214 ( .B1(n477), .B2(n670), .A(n657), .ZN(n497) );
  NAND2_X1 U215 ( .A1(\mem[7][12] ), .A2(n670), .ZN(n657) );
  OAI21_X1 U216 ( .B1(n476), .B2(n458), .A(n656), .ZN(n496) );
  NAND2_X1 U217 ( .A1(\mem[7][13] ), .A2(n670), .ZN(n656) );
  OAI21_X1 U218 ( .B1(n475), .B2(n458), .A(n655), .ZN(n495) );
  NAND2_X1 U219 ( .A1(\mem[7][14] ), .A2(n670), .ZN(n655) );
  OAI21_X1 U220 ( .B1(n474), .B2(n670), .A(n654), .ZN(n494) );
  NAND2_X1 U221 ( .A1(\mem[7][15] ), .A2(n670), .ZN(n654) );
  OAI21_X1 U222 ( .B1(n473), .B2(n670), .A(n653), .ZN(n493) );
  NAND2_X1 U223 ( .A1(\mem[7][16] ), .A2(n670), .ZN(n653) );
  OAI21_X1 U224 ( .B1(n472), .B2(n670), .A(n652), .ZN(n492) );
  NAND2_X1 U225 ( .A1(\mem[7][17] ), .A2(n670), .ZN(n652) );
  OAI21_X1 U226 ( .B1(n471), .B2(n670), .A(n651), .ZN(n491) );
  NAND2_X1 U227 ( .A1(\mem[7][18] ), .A2(n670), .ZN(n651) );
  OAI21_X1 U228 ( .B1(n470), .B2(n670), .A(n650), .ZN(n490) );
  NAND2_X1 U229 ( .A1(\mem[7][19] ), .A2(n458), .ZN(n650) );
  NAND2_X1 U230 ( .A1(wr_en), .A2(n469), .ZN(n735) );
  INV_X1 U231 ( .A(addr[3]), .ZN(n469) );
  OAI21_X1 U232 ( .B1(n465), .B2(n489), .A(n819), .ZN(n649) );
  NAND2_X1 U233 ( .A1(\mem[0][0] ), .A2(n465), .ZN(n819) );
  OAI21_X1 U234 ( .B1(n820), .B2(n488), .A(n818), .ZN(n648) );
  NAND2_X1 U235 ( .A1(\mem[0][1] ), .A2(n465), .ZN(n818) );
  OAI21_X1 U236 ( .B1(n820), .B2(n487), .A(n817), .ZN(n647) );
  NAND2_X1 U237 ( .A1(\mem[0][2] ), .A2(n465), .ZN(n817) );
  OAI21_X1 U238 ( .B1(n820), .B2(n486), .A(n816), .ZN(n646) );
  NAND2_X1 U239 ( .A1(\mem[0][3] ), .A2(n465), .ZN(n816) );
  OAI21_X1 U240 ( .B1(n820), .B2(n485), .A(n815), .ZN(n645) );
  NAND2_X1 U241 ( .A1(\mem[0][4] ), .A2(n465), .ZN(n815) );
  OAI21_X1 U242 ( .B1(n820), .B2(n484), .A(n814), .ZN(n644) );
  NAND2_X1 U243 ( .A1(\mem[0][5] ), .A2(n465), .ZN(n814) );
  OAI21_X1 U244 ( .B1(n820), .B2(n483), .A(n813), .ZN(n643) );
  NAND2_X1 U245 ( .A1(\mem[0][6] ), .A2(n465), .ZN(n813) );
  OAI21_X1 U246 ( .B1(n820), .B2(n482), .A(n812), .ZN(n642) );
  NAND2_X1 U247 ( .A1(\mem[0][7] ), .A2(n465), .ZN(n812) );
  OAI21_X1 U248 ( .B1(n820), .B2(n481), .A(n811), .ZN(n641) );
  NAND2_X1 U249 ( .A1(\mem[0][8] ), .A2(n465), .ZN(n811) );
  OAI21_X1 U250 ( .B1(n820), .B2(n480), .A(n810), .ZN(n640) );
  NAND2_X1 U251 ( .A1(\mem[0][9] ), .A2(n465), .ZN(n810) );
  OAI21_X1 U252 ( .B1(n820), .B2(n479), .A(n809), .ZN(n639) );
  NAND2_X1 U253 ( .A1(\mem[0][10] ), .A2(n465), .ZN(n809) );
  OAI21_X1 U254 ( .B1(n820), .B2(n478), .A(n808), .ZN(n638) );
  NAND2_X1 U255 ( .A1(\mem[0][11] ), .A2(n465), .ZN(n808) );
  OAI21_X1 U256 ( .B1(n489), .B2(n798), .A(n797), .ZN(n629) );
  NAND2_X1 U257 ( .A1(\mem[1][0] ), .A2(n798), .ZN(n797) );
  OAI21_X1 U258 ( .B1(n488), .B2(n798), .A(n796), .ZN(n628) );
  NAND2_X1 U259 ( .A1(\mem[1][1] ), .A2(n798), .ZN(n796) );
  OAI21_X1 U260 ( .B1(n487), .B2(n798), .A(n795), .ZN(n627) );
  NAND2_X1 U261 ( .A1(\mem[1][2] ), .A2(n798), .ZN(n795) );
  OAI21_X1 U262 ( .B1(n486), .B2(n798), .A(n794), .ZN(n626) );
  NAND2_X1 U263 ( .A1(\mem[1][3] ), .A2(n464), .ZN(n794) );
  OAI21_X1 U264 ( .B1(n485), .B2(n798), .A(n793), .ZN(n625) );
  NAND2_X1 U265 ( .A1(\mem[1][4] ), .A2(n464), .ZN(n793) );
  OAI21_X1 U266 ( .B1(n484), .B2(n798), .A(n792), .ZN(n624) );
  NAND2_X1 U267 ( .A1(\mem[1][5] ), .A2(n464), .ZN(n792) );
  OAI21_X1 U268 ( .B1(n483), .B2(n798), .A(n791), .ZN(n623) );
  NAND2_X1 U269 ( .A1(\mem[1][6] ), .A2(n798), .ZN(n791) );
  OAI21_X1 U270 ( .B1(n482), .B2(n798), .A(n790), .ZN(n622) );
  NAND2_X1 U271 ( .A1(\mem[1][7] ), .A2(n798), .ZN(n790) );
  OAI21_X1 U272 ( .B1(n481), .B2(n798), .A(n789), .ZN(n621) );
  NAND2_X1 U273 ( .A1(\mem[1][8] ), .A2(n798), .ZN(n789) );
  OAI21_X1 U274 ( .B1(n480), .B2(n464), .A(n788), .ZN(n620) );
  NAND2_X1 U275 ( .A1(\mem[1][9] ), .A2(n464), .ZN(n788) );
  OAI21_X1 U276 ( .B1(n479), .B2(n798), .A(n787), .ZN(n619) );
  NAND2_X1 U277 ( .A1(\mem[1][10] ), .A2(n798), .ZN(n787) );
  OAI21_X1 U278 ( .B1(n478), .B2(n798), .A(n786), .ZN(n618) );
  NAND2_X1 U279 ( .A1(\mem[1][11] ), .A2(n798), .ZN(n786) );
  OAI21_X1 U280 ( .B1(n489), .B2(n777), .A(n776), .ZN(n609) );
  NAND2_X1 U281 ( .A1(\mem[2][0] ), .A2(n463), .ZN(n776) );
  OAI21_X1 U282 ( .B1(n488), .B2(n777), .A(n775), .ZN(n608) );
  NAND2_X1 U283 ( .A1(\mem[2][1] ), .A2(n463), .ZN(n775) );
  OAI21_X1 U284 ( .B1(n487), .B2(n777), .A(n774), .ZN(n607) );
  NAND2_X1 U285 ( .A1(\mem[2][2] ), .A2(n463), .ZN(n774) );
  OAI21_X1 U286 ( .B1(n486), .B2(n777), .A(n773), .ZN(n606) );
  NAND2_X1 U287 ( .A1(\mem[2][3] ), .A2(n463), .ZN(n773) );
  OAI21_X1 U288 ( .B1(n485), .B2(n777), .A(n772), .ZN(n605) );
  NAND2_X1 U289 ( .A1(\mem[2][4] ), .A2(n463), .ZN(n772) );
  OAI21_X1 U290 ( .B1(n484), .B2(n777), .A(n771), .ZN(n604) );
  NAND2_X1 U291 ( .A1(\mem[2][5] ), .A2(n463), .ZN(n771) );
  OAI21_X1 U292 ( .B1(n483), .B2(n777), .A(n770), .ZN(n603) );
  NAND2_X1 U293 ( .A1(\mem[2][6] ), .A2(n463), .ZN(n770) );
  OAI21_X1 U294 ( .B1(n482), .B2(n777), .A(n769), .ZN(n602) );
  NAND2_X1 U295 ( .A1(\mem[2][7] ), .A2(n463), .ZN(n769) );
  OAI21_X1 U296 ( .B1(n481), .B2(n777), .A(n768), .ZN(n601) );
  NAND2_X1 U297 ( .A1(\mem[2][8] ), .A2(n463), .ZN(n768) );
  OAI21_X1 U298 ( .B1(n480), .B2(n463), .A(n767), .ZN(n600) );
  NAND2_X1 U299 ( .A1(\mem[2][9] ), .A2(n463), .ZN(n767) );
  OAI21_X1 U300 ( .B1(n479), .B2(n777), .A(n766), .ZN(n599) );
  NAND2_X1 U301 ( .A1(\mem[2][10] ), .A2(n463), .ZN(n766) );
  OAI21_X1 U302 ( .B1(n478), .B2(n777), .A(n765), .ZN(n598) );
  NAND2_X1 U303 ( .A1(\mem[2][11] ), .A2(n463), .ZN(n765) );
  OAI21_X1 U304 ( .B1(n489), .B2(n462), .A(n755), .ZN(n589) );
  NAND2_X1 U305 ( .A1(\mem[3][0] ), .A2(n756), .ZN(n755) );
  OAI21_X1 U306 ( .B1(n488), .B2(n462), .A(n754), .ZN(n588) );
  NAND2_X1 U307 ( .A1(\mem[3][1] ), .A2(n756), .ZN(n754) );
  OAI21_X1 U308 ( .B1(n487), .B2(n462), .A(n753), .ZN(n587) );
  NAND2_X1 U309 ( .A1(\mem[3][2] ), .A2(n756), .ZN(n753) );
  OAI21_X1 U310 ( .B1(n486), .B2(n462), .A(n752), .ZN(n586) );
  NAND2_X1 U311 ( .A1(\mem[3][3] ), .A2(n756), .ZN(n752) );
  OAI21_X1 U312 ( .B1(n485), .B2(n462), .A(n751), .ZN(n585) );
  NAND2_X1 U313 ( .A1(\mem[3][4] ), .A2(n756), .ZN(n751) );
  OAI21_X1 U314 ( .B1(n484), .B2(n462), .A(n750), .ZN(n584) );
  NAND2_X1 U315 ( .A1(\mem[3][5] ), .A2(n756), .ZN(n750) );
  OAI21_X1 U316 ( .B1(n483), .B2(n462), .A(n749), .ZN(n583) );
  NAND2_X1 U317 ( .A1(\mem[3][6] ), .A2(n756), .ZN(n749) );
  OAI21_X1 U318 ( .B1(n482), .B2(n462), .A(n748), .ZN(n582) );
  NAND2_X1 U319 ( .A1(\mem[3][7] ), .A2(n756), .ZN(n748) );
  OAI21_X1 U320 ( .B1(n481), .B2(n462), .A(n747), .ZN(n581) );
  NAND2_X1 U321 ( .A1(\mem[3][8] ), .A2(n756), .ZN(n747) );
  OAI21_X1 U322 ( .B1(n480), .B2(n756), .A(n746), .ZN(n580) );
  NAND2_X1 U323 ( .A1(\mem[3][9] ), .A2(n756), .ZN(n746) );
  OAI21_X1 U324 ( .B1(n479), .B2(n462), .A(n745), .ZN(n579) );
  NAND2_X1 U325 ( .A1(\mem[3][10] ), .A2(n756), .ZN(n745) );
  OAI21_X1 U326 ( .B1(n478), .B2(n462), .A(n744), .ZN(n578) );
  NAND2_X1 U327 ( .A1(\mem[3][11] ), .A2(n756), .ZN(n744) );
  OAI21_X1 U328 ( .B1(n820), .B2(n477), .A(n807), .ZN(n637) );
  NAND2_X1 U329 ( .A1(\mem[0][12] ), .A2(n820), .ZN(n807) );
  OAI21_X1 U330 ( .B1(n820), .B2(n476), .A(n806), .ZN(n636) );
  NAND2_X1 U331 ( .A1(\mem[0][13] ), .A2(n820), .ZN(n806) );
  OAI21_X1 U332 ( .B1(n465), .B2(n475), .A(n805), .ZN(n635) );
  NAND2_X1 U333 ( .A1(\mem[0][14] ), .A2(n820), .ZN(n805) );
  OAI21_X1 U334 ( .B1(n820), .B2(n474), .A(n804), .ZN(n634) );
  NAND2_X1 U335 ( .A1(\mem[0][15] ), .A2(n465), .ZN(n804) );
  OAI21_X1 U336 ( .B1(n820), .B2(n473), .A(n803), .ZN(n633) );
  NAND2_X1 U337 ( .A1(\mem[0][16] ), .A2(n820), .ZN(n803) );
  OAI21_X1 U338 ( .B1(n820), .B2(n472), .A(n802), .ZN(n632) );
  NAND2_X1 U339 ( .A1(\mem[0][17] ), .A2(n820), .ZN(n802) );
  OAI21_X1 U340 ( .B1(n820), .B2(n471), .A(n801), .ZN(n631) );
  NAND2_X1 U341 ( .A1(\mem[0][18] ), .A2(n820), .ZN(n801) );
  OAI21_X1 U342 ( .B1(n820), .B2(n470), .A(n800), .ZN(n630) );
  NAND2_X1 U343 ( .A1(\mem[0][19] ), .A2(n465), .ZN(n800) );
  INV_X1 U344 ( .A(data_in[0]), .ZN(n489) );
  INV_X1 U345 ( .A(data_in[1]), .ZN(n488) );
  INV_X1 U346 ( .A(data_in[2]), .ZN(n487) );
  INV_X1 U347 ( .A(data_in[3]), .ZN(n486) );
  INV_X1 U348 ( .A(data_in[4]), .ZN(n485) );
  INV_X1 U349 ( .A(data_in[5]), .ZN(n484) );
  INV_X1 U358 ( .A(data_in[6]), .ZN(n483) );
  INV_X1 U359 ( .A(data_in[7]), .ZN(n482) );
  INV_X1 U360 ( .A(data_in[8]), .ZN(n481) );
  INV_X1 U361 ( .A(data_in[9]), .ZN(n480) );
  INV_X1 U362 ( .A(data_in[10]), .ZN(n479) );
  INV_X1 U363 ( .A(data_in[11]), .ZN(n478) );
  INV_X1 U364 ( .A(data_in[12]), .ZN(n477) );
  INV_X1 U365 ( .A(data_in[13]), .ZN(n476) );
  INV_X1 U366 ( .A(data_in[14]), .ZN(n475) );
  INV_X1 U367 ( .A(data_in[15]), .ZN(n474) );
  INV_X1 U368 ( .A(data_in[16]), .ZN(n473) );
  INV_X1 U369 ( .A(data_in[17]), .ZN(n472) );
  INV_X1 U370 ( .A(data_in[18]), .ZN(n471) );
  INV_X1 U371 ( .A(data_in[19]), .ZN(n470) );
  MUX2_X1 U372 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n456), .Z(n1) );
  MUX2_X1 U373 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n457), .Z(n2) );
  MUX2_X1 U374 ( .A(n2), .B(n1), .S(n453), .Z(n3) );
  MUX2_X1 U375 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n455), .Z(n4) );
  MUX2_X1 U376 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n454), .Z(n5) );
  MUX2_X1 U377 ( .A(n5), .B(n4), .S(n453), .Z(n6) );
  MUX2_X1 U378 ( .A(n6), .B(n3), .S(N12), .Z(N32) );
  MUX2_X1 U379 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n454), .Z(n7) );
  MUX2_X1 U380 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n456), .Z(n8) );
  MUX2_X1 U381 ( .A(n8), .B(n7), .S(n453), .Z(n9) );
  MUX2_X1 U382 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n456), .Z(n10) );
  MUX2_X1 U383 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n457), .Z(n11) );
  MUX2_X1 U384 ( .A(n11), .B(n10), .S(n453), .Z(n12) );
  MUX2_X1 U385 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n454), .Z(n13) );
  MUX2_X1 U386 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n454), .Z(n14) );
  MUX2_X1 U387 ( .A(n14), .B(n13), .S(n453), .Z(n15) );
  MUX2_X1 U388 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n454), .Z(n16) );
  MUX2_X1 U389 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n454), .Z(n17) );
  MUX2_X1 U390 ( .A(n17), .B(n16), .S(n453), .Z(n18) );
  MUX2_X1 U391 ( .A(n18), .B(n15), .S(N12), .Z(N30) );
  MUX2_X1 U392 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n454), .Z(n19) );
  MUX2_X1 U393 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n454), .Z(n20) );
  MUX2_X1 U394 ( .A(n20), .B(n19), .S(N11), .Z(n21) );
  MUX2_X1 U395 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n454), .Z(n22) );
  MUX2_X1 U396 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n454), .Z(n23) );
  MUX2_X1 U397 ( .A(n23), .B(n22), .S(N11), .Z(n24) );
  MUX2_X1 U398 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n454), .Z(n356) );
  MUX2_X1 U399 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n454), .Z(n357) );
  MUX2_X1 U400 ( .A(n357), .B(n356), .S(n453), .Z(n358) );
  MUX2_X1 U401 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n454), .Z(n359) );
  MUX2_X1 U402 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n454), .Z(n360) );
  MUX2_X1 U403 ( .A(n360), .B(n359), .S(n453), .Z(n361) );
  MUX2_X1 U404 ( .A(n361), .B(n358), .S(N12), .Z(N28) );
  MUX2_X1 U405 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n454), .Z(n362) );
  MUX2_X1 U406 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n457), .Z(n363) );
  MUX2_X1 U407 ( .A(n363), .B(n362), .S(n453), .Z(n364) );
  MUX2_X1 U408 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n454), .Z(n365) );
  MUX2_X1 U409 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n455), .Z(n366) );
  MUX2_X1 U410 ( .A(n366), .B(n365), .S(N11), .Z(n367) );
  MUX2_X1 U411 ( .A(n367), .B(n364), .S(N12), .Z(N27) );
  MUX2_X1 U412 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n456), .Z(n368) );
  MUX2_X1 U413 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n455), .Z(n369) );
  MUX2_X1 U414 ( .A(n369), .B(n368), .S(n453), .Z(n370) );
  MUX2_X1 U415 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n457), .Z(n371) );
  MUX2_X1 U416 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n456), .Z(n372) );
  MUX2_X1 U417 ( .A(n372), .B(n371), .S(N11), .Z(n373) );
  MUX2_X1 U418 ( .A(n373), .B(n370), .S(N12), .Z(N26) );
  MUX2_X1 U419 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n457), .Z(n374) );
  MUX2_X1 U420 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n455), .Z(n375) );
  MUX2_X1 U421 ( .A(n375), .B(n374), .S(N11), .Z(n376) );
  MUX2_X1 U422 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n454), .Z(n377) );
  MUX2_X1 U423 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n455), .Z(n378) );
  MUX2_X1 U424 ( .A(n378), .B(n377), .S(N11), .Z(n379) );
  MUX2_X1 U425 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n455), .Z(n380) );
  MUX2_X1 U426 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n457), .Z(n381) );
  MUX2_X1 U427 ( .A(n381), .B(n380), .S(n453), .Z(n382) );
  MUX2_X1 U428 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n455), .Z(n383) );
  MUX2_X1 U429 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n455), .Z(n384) );
  MUX2_X1 U430 ( .A(n384), .B(n383), .S(n453), .Z(n385) );
  MUX2_X1 U431 ( .A(n385), .B(n382), .S(N12), .Z(N24) );
  MUX2_X1 U432 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n457), .Z(n386) );
  MUX2_X1 U433 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n456), .Z(n387) );
  MUX2_X1 U434 ( .A(n387), .B(n386), .S(n453), .Z(n388) );
  MUX2_X1 U435 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n454), .Z(n389) );
  MUX2_X1 U436 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n454), .Z(n390) );
  MUX2_X1 U437 ( .A(n390), .B(n389), .S(n453), .Z(n391) );
  MUX2_X1 U438 ( .A(n391), .B(n388), .S(N12), .Z(N23) );
  MUX2_X1 U439 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n454), .Z(n392) );
  MUX2_X1 U440 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n457), .Z(n393) );
  MUX2_X1 U441 ( .A(n393), .B(n392), .S(n453), .Z(n394) );
  MUX2_X1 U442 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n456), .Z(n395) );
  MUX2_X1 U443 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n456), .Z(n396) );
  MUX2_X1 U444 ( .A(n396), .B(n395), .S(n453), .Z(n397) );
  MUX2_X1 U445 ( .A(n397), .B(n394), .S(N12), .Z(N22) );
  MUX2_X1 U446 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n455), .Z(n398) );
  MUX2_X1 U447 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n455), .Z(n399) );
  MUX2_X1 U448 ( .A(n399), .B(n398), .S(n453), .Z(n400) );
  MUX2_X1 U449 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n455), .Z(n401) );
  MUX2_X1 U450 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n455), .Z(n402) );
  MUX2_X1 U451 ( .A(n402), .B(n401), .S(n453), .Z(n403) );
  MUX2_X1 U452 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n455), .Z(n404) );
  MUX2_X1 U453 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n455), .Z(n405) );
  MUX2_X1 U454 ( .A(n405), .B(n404), .S(n453), .Z(n406) );
  MUX2_X1 U455 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n455), .Z(n407) );
  MUX2_X1 U456 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n455), .Z(n408) );
  MUX2_X1 U457 ( .A(n408), .B(n407), .S(n453), .Z(n409) );
  MUX2_X1 U458 ( .A(n409), .B(n406), .S(N12), .Z(N20) );
  MUX2_X1 U459 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n455), .Z(n410) );
  MUX2_X1 U460 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n455), .Z(n411) );
  MUX2_X1 U461 ( .A(n411), .B(n410), .S(n453), .Z(n412) );
  MUX2_X1 U462 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n455), .Z(n413) );
  MUX2_X1 U463 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n455), .Z(n414) );
  MUX2_X1 U464 ( .A(n414), .B(n413), .S(n453), .Z(n415) );
  MUX2_X1 U465 ( .A(n415), .B(n412), .S(N12), .Z(N19) );
  MUX2_X1 U466 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n456), .Z(n416) );
  MUX2_X1 U467 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n456), .Z(n417) );
  MUX2_X1 U468 ( .A(n417), .B(n416), .S(n452), .Z(n418) );
  MUX2_X1 U469 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n456), .Z(n419) );
  MUX2_X1 U470 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n456), .Z(n420) );
  MUX2_X1 U471 ( .A(n420), .B(n419), .S(n452), .Z(n421) );
  MUX2_X1 U472 ( .A(n421), .B(n418), .S(N12), .Z(N18) );
  MUX2_X1 U473 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n456), .Z(n422) );
  MUX2_X1 U474 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n456), .Z(n423) );
  MUX2_X1 U475 ( .A(n423), .B(n422), .S(n452), .Z(n424) );
  MUX2_X1 U476 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n456), .Z(n425) );
  MUX2_X1 U477 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n456), .Z(n426) );
  MUX2_X1 U478 ( .A(n426), .B(n425), .S(n452), .Z(n427) );
  MUX2_X1 U479 ( .A(n427), .B(n424), .S(N12), .Z(N17) );
  MUX2_X1 U480 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n456), .Z(n428) );
  MUX2_X1 U481 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n456), .Z(n429) );
  MUX2_X1 U482 ( .A(n429), .B(n428), .S(n452), .Z(n430) );
  MUX2_X1 U483 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n456), .Z(n431) );
  MUX2_X1 U484 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n456), .Z(n432) );
  MUX2_X1 U485 ( .A(n432), .B(n431), .S(n452), .Z(n433) );
  MUX2_X1 U486 ( .A(n433), .B(n430), .S(N12), .Z(N16) );
  MUX2_X1 U487 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n457), .Z(n434) );
  MUX2_X1 U488 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n457), .Z(n435) );
  MUX2_X1 U489 ( .A(n435), .B(n434), .S(n452), .Z(n436) );
  MUX2_X1 U490 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n457), .Z(n437) );
  MUX2_X1 U491 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n457), .Z(n438) );
  MUX2_X1 U492 ( .A(n438), .B(n437), .S(n452), .Z(n439) );
  MUX2_X1 U493 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n457), .Z(n440) );
  MUX2_X1 U494 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n457), .Z(n441) );
  MUX2_X1 U495 ( .A(n441), .B(n440), .S(n452), .Z(n442) );
  MUX2_X1 U496 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n457), .Z(n443) );
  MUX2_X1 U497 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n457), .Z(n444) );
  MUX2_X1 U498 ( .A(n444), .B(n443), .S(n452), .Z(n445) );
  MUX2_X1 U499 ( .A(n445), .B(n442), .S(N12), .Z(N14) );
  MUX2_X1 U500 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n457), .Z(n446) );
  MUX2_X1 U501 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n457), .Z(n447) );
  MUX2_X1 U502 ( .A(n447), .B(n446), .S(n452), .Z(n448) );
  MUX2_X1 U503 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n457), .Z(n449) );
  MUX2_X1 U504 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n457), .Z(n450) );
  MUX2_X1 U505 ( .A(n450), .B(n449), .S(n452), .Z(n451) );
  MUX2_X1 U506 ( .A(n451), .B(n448), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE4_4 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N13, N14, N16, N17, N18, N20, N22, N23, N24, N26, N27,
         N28, N30, N31, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[19]  ( .D(N13), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[15]  ( .D(N17), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N20), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N23), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N27), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N30), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N31), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n490), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n491), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n492), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n493), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n494), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n495), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n496), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n497), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n498), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n499), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n500), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n501), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n502), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n503), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n504), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n505), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n506), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n507), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n508), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n509), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n510), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n511), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n512), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n513), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n514), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n515), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n516), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n517), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n518), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n519), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n520), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n521), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n522), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n523), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n524), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n525), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n526), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n527), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n528), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n529), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n530), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n531), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n532), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n533), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n534), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n535), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n536), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n537), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n538), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n539), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n540), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n541), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n542), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n543), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n544), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n545), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n546), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n547), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n548), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n549), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n550), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n551), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n552), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n553), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n554), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n555), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n556), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n557), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n558), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n559), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n560), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n561), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n562), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n563), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n564), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n565), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n566), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n567), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n568), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n569), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n570), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n571), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n572), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n573), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n574), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n575), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n576), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n577), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n578), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n579), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n580), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n581), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n582), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n583), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n584), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n585), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n586), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n587), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n588), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n589), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n590), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n591), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n592), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n593), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n594), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n595), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n596), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n597), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n598), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n599), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n600), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n601), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n602), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n603), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n604), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n605), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n606), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n607), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n608), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n609), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n610), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n611), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n612), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n613), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n614), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n615), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n616), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n617), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n618), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n619), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n620), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n621), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n622), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n623), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n624), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n625), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n626), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n627), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n628), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n629), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n630), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n631), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n632), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n633), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n634), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n635), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n636), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n637), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n638), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n639), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n640), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n641), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n642), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n643), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n644), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n645), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n646), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n647), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n648), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n649), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U350 ( .A1(n466), .A2(n467), .A3(n799), .ZN(n820) );
  NAND3_X1 U351 ( .A1(n799), .A2(n467), .A3(N10), .ZN(n798) );
  NAND3_X1 U352 ( .A1(n799), .A2(n466), .A3(N11), .ZN(n777) );
  NAND3_X1 U353 ( .A1(N10), .A2(n799), .A3(N11), .ZN(n756) );
  NAND3_X1 U354 ( .A1(n466), .A2(n467), .A3(n713), .ZN(n734) );
  NAND3_X1 U355 ( .A1(N10), .A2(n467), .A3(n713), .ZN(n712) );
  NAND3_X1 U356 ( .A1(N11), .A2(n466), .A3(n713), .ZN(n691) );
  NAND3_X1 U357 ( .A1(N11), .A2(N10), .A3(n713), .ZN(n670) );
  SDFF_X1 \data_out_reg[13]  ( .D(n412), .SI(n415), .SE(n468), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n3), .SI(n6), .SE(n468), .CK(clk), .Q(
        data_out[0]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n21), .SI(n24), .SE(n468), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n376), .SI(n379), .SE(n468), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[17]  ( .D(n436), .SI(n439), .SE(n468), .CK(clk), .Q(
        data_out[17]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n400), .SI(n403), .SE(n468), .CK(clk), .Q(
        data_out[11]) );
  BUF_X1 U3 ( .A(n670), .Z(n458) );
  BUF_X1 U4 ( .A(n798), .Z(n464) );
  BUF_X1 U5 ( .A(n734), .Z(n461) );
  BUF_X1 U6 ( .A(n453), .Z(n452) );
  BUF_X1 U7 ( .A(N10), .Z(n455) );
  BUF_X1 U8 ( .A(N10), .Z(n456) );
  BUF_X1 U9 ( .A(N10), .Z(n457) );
  BUF_X1 U10 ( .A(N10), .Z(n454) );
  BUF_X1 U11 ( .A(n820), .Z(n465) );
  BUF_X1 U12 ( .A(n756), .Z(n462) );
  BUF_X1 U13 ( .A(n777), .Z(n463) );
  BUF_X1 U14 ( .A(n712), .Z(n460) );
  BUF_X1 U15 ( .A(n691), .Z(n459) );
  BUF_X1 U16 ( .A(N11), .Z(n453) );
  NOR2_X1 U17 ( .A1(n735), .A2(N12), .ZN(n799) );
  NOR2_X1 U18 ( .A1(n468), .A2(n735), .ZN(n713) );
  INV_X1 U19 ( .A(N12), .ZN(n468) );
  INV_X1 U20 ( .A(N11), .ZN(n467) );
  INV_X1 U21 ( .A(N10), .ZN(n466) );
  OAI21_X1 U22 ( .B1(n477), .B2(n798), .A(n785), .ZN(n617) );
  NAND2_X1 U23 ( .A1(\mem[1][12] ), .A2(n798), .ZN(n785) );
  OAI21_X1 U24 ( .B1(n476), .B2(n798), .A(n784), .ZN(n616) );
  NAND2_X1 U25 ( .A1(\mem[1][13] ), .A2(n798), .ZN(n784) );
  OAI21_X1 U26 ( .B1(n475), .B2(n464), .A(n783), .ZN(n615) );
  NAND2_X1 U27 ( .A1(\mem[1][14] ), .A2(n798), .ZN(n783) );
  OAI21_X1 U28 ( .B1(n474), .B2(n464), .A(n782), .ZN(n614) );
  NAND2_X1 U29 ( .A1(\mem[1][15] ), .A2(n798), .ZN(n782) );
  OAI21_X1 U30 ( .B1(n473), .B2(n464), .A(n781), .ZN(n613) );
  NAND2_X1 U31 ( .A1(\mem[1][16] ), .A2(n798), .ZN(n781) );
  OAI21_X1 U32 ( .B1(n472), .B2(n464), .A(n780), .ZN(n612) );
  NAND2_X1 U33 ( .A1(\mem[1][17] ), .A2(n798), .ZN(n780) );
  OAI21_X1 U34 ( .B1(n471), .B2(n464), .A(n779), .ZN(n611) );
  NAND2_X1 U35 ( .A1(\mem[1][18] ), .A2(n798), .ZN(n779) );
  OAI21_X1 U36 ( .B1(n470), .B2(n798), .A(n778), .ZN(n610) );
  NAND2_X1 U37 ( .A1(\mem[1][19] ), .A2(n798), .ZN(n778) );
  OAI21_X1 U38 ( .B1(n477), .B2(n777), .A(n764), .ZN(n597) );
  NAND2_X1 U39 ( .A1(\mem[2][12] ), .A2(n777), .ZN(n764) );
  OAI21_X1 U40 ( .B1(n476), .B2(n777), .A(n763), .ZN(n596) );
  NAND2_X1 U41 ( .A1(\mem[2][13] ), .A2(n777), .ZN(n763) );
  OAI21_X1 U42 ( .B1(n475), .B2(n777), .A(n762), .ZN(n595) );
  NAND2_X1 U43 ( .A1(\mem[2][14] ), .A2(n777), .ZN(n762) );
  OAI21_X1 U44 ( .B1(n474), .B2(n463), .A(n761), .ZN(n594) );
  NAND2_X1 U45 ( .A1(\mem[2][15] ), .A2(n777), .ZN(n761) );
  OAI21_X1 U46 ( .B1(n473), .B2(n777), .A(n760), .ZN(n593) );
  NAND2_X1 U47 ( .A1(\mem[2][16] ), .A2(n463), .ZN(n760) );
  OAI21_X1 U48 ( .B1(n472), .B2(n777), .A(n759), .ZN(n592) );
  NAND2_X1 U49 ( .A1(\mem[2][17] ), .A2(n777), .ZN(n759) );
  OAI21_X1 U50 ( .B1(n471), .B2(n777), .A(n758), .ZN(n591) );
  NAND2_X1 U51 ( .A1(\mem[2][18] ), .A2(n777), .ZN(n758) );
  OAI21_X1 U52 ( .B1(n470), .B2(n777), .A(n757), .ZN(n590) );
  NAND2_X1 U53 ( .A1(\mem[2][19] ), .A2(n463), .ZN(n757) );
  OAI21_X1 U54 ( .B1(n477), .B2(n756), .A(n743), .ZN(n577) );
  NAND2_X1 U55 ( .A1(\mem[3][12] ), .A2(n756), .ZN(n743) );
  OAI21_X1 U56 ( .B1(n476), .B2(n756), .A(n742), .ZN(n576) );
  NAND2_X1 U57 ( .A1(\mem[3][13] ), .A2(n756), .ZN(n742) );
  OAI21_X1 U58 ( .B1(n475), .B2(n756), .A(n741), .ZN(n575) );
  NAND2_X1 U59 ( .A1(\mem[3][14] ), .A2(n756), .ZN(n741) );
  OAI21_X1 U60 ( .B1(n474), .B2(n462), .A(n740), .ZN(n574) );
  NAND2_X1 U61 ( .A1(\mem[3][15] ), .A2(n756), .ZN(n740) );
  OAI21_X1 U62 ( .B1(n473), .B2(n756), .A(n739), .ZN(n573) );
  NAND2_X1 U63 ( .A1(\mem[3][16] ), .A2(n462), .ZN(n739) );
  OAI21_X1 U64 ( .B1(n472), .B2(n756), .A(n738), .ZN(n572) );
  NAND2_X1 U65 ( .A1(\mem[3][17] ), .A2(n756), .ZN(n738) );
  OAI21_X1 U66 ( .B1(n471), .B2(n756), .A(n737), .ZN(n571) );
  NAND2_X1 U67 ( .A1(\mem[3][18] ), .A2(n756), .ZN(n737) );
  OAI21_X1 U68 ( .B1(n470), .B2(n756), .A(n736), .ZN(n570) );
  NAND2_X1 U69 ( .A1(\mem[3][19] ), .A2(n462), .ZN(n736) );
  OAI21_X1 U70 ( .B1(n489), .B2(n734), .A(n733), .ZN(n569) );
  NAND2_X1 U71 ( .A1(\mem[4][0] ), .A2(n734), .ZN(n733) );
  OAI21_X1 U72 ( .B1(n488), .B2(n461), .A(n732), .ZN(n568) );
  NAND2_X1 U73 ( .A1(\mem[4][1] ), .A2(n734), .ZN(n732) );
  OAI21_X1 U74 ( .B1(n487), .B2(n461), .A(n731), .ZN(n567) );
  NAND2_X1 U75 ( .A1(\mem[4][2] ), .A2(n734), .ZN(n731) );
  OAI21_X1 U76 ( .B1(n486), .B2(n461), .A(n730), .ZN(n566) );
  NAND2_X1 U77 ( .A1(\mem[4][3] ), .A2(n734), .ZN(n730) );
  OAI21_X1 U78 ( .B1(n485), .B2(n461), .A(n729), .ZN(n565) );
  NAND2_X1 U79 ( .A1(\mem[4][4] ), .A2(n734), .ZN(n729) );
  OAI21_X1 U80 ( .B1(n484), .B2(n461), .A(n728), .ZN(n564) );
  NAND2_X1 U81 ( .A1(\mem[4][5] ), .A2(n734), .ZN(n728) );
  OAI21_X1 U82 ( .B1(n483), .B2(n461), .A(n727), .ZN(n563) );
  NAND2_X1 U83 ( .A1(\mem[4][6] ), .A2(n734), .ZN(n727) );
  OAI21_X1 U84 ( .B1(n482), .B2(n461), .A(n726), .ZN(n562) );
  NAND2_X1 U85 ( .A1(\mem[4][7] ), .A2(n734), .ZN(n726) );
  OAI21_X1 U86 ( .B1(n481), .B2(n461), .A(n725), .ZN(n561) );
  NAND2_X1 U87 ( .A1(\mem[4][8] ), .A2(n734), .ZN(n725) );
  OAI21_X1 U88 ( .B1(n480), .B2(n734), .A(n724), .ZN(n560) );
  NAND2_X1 U89 ( .A1(\mem[4][9] ), .A2(n734), .ZN(n724) );
  OAI21_X1 U90 ( .B1(n479), .B2(n461), .A(n723), .ZN(n559) );
  NAND2_X1 U91 ( .A1(\mem[4][10] ), .A2(n734), .ZN(n723) );
  OAI21_X1 U92 ( .B1(n478), .B2(n461), .A(n722), .ZN(n558) );
  NAND2_X1 U93 ( .A1(\mem[4][11] ), .A2(n734), .ZN(n722) );
  OAI21_X1 U94 ( .B1(n477), .B2(n734), .A(n721), .ZN(n557) );
  NAND2_X1 U95 ( .A1(\mem[4][12] ), .A2(n734), .ZN(n721) );
  OAI21_X1 U96 ( .B1(n476), .B2(n461), .A(n720), .ZN(n556) );
  NAND2_X1 U97 ( .A1(\mem[4][13] ), .A2(n734), .ZN(n720) );
  OAI21_X1 U98 ( .B1(n475), .B2(n734), .A(n719), .ZN(n555) );
  NAND2_X1 U99 ( .A1(\mem[4][14] ), .A2(n734), .ZN(n719) );
  OAI21_X1 U100 ( .B1(n474), .B2(n461), .A(n718), .ZN(n554) );
  NAND2_X1 U101 ( .A1(\mem[4][15] ), .A2(n734), .ZN(n718) );
  OAI21_X1 U102 ( .B1(n473), .B2(n461), .A(n717), .ZN(n553) );
  NAND2_X1 U103 ( .A1(\mem[4][16] ), .A2(n734), .ZN(n717) );
  OAI21_X1 U104 ( .B1(n472), .B2(n461), .A(n716), .ZN(n552) );
  NAND2_X1 U105 ( .A1(\mem[4][17] ), .A2(n734), .ZN(n716) );
  OAI21_X1 U106 ( .B1(n471), .B2(n461), .A(n715), .ZN(n551) );
  NAND2_X1 U107 ( .A1(\mem[4][18] ), .A2(n734), .ZN(n715) );
  OAI21_X1 U108 ( .B1(n470), .B2(n461), .A(n714), .ZN(n550) );
  NAND2_X1 U109 ( .A1(\mem[4][19] ), .A2(n734), .ZN(n714) );
  OAI21_X1 U110 ( .B1(n489), .B2(n712), .A(n711), .ZN(n549) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n460), .ZN(n711) );
  OAI21_X1 U112 ( .B1(n488), .B2(n712), .A(n710), .ZN(n548) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n460), .ZN(n710) );
  OAI21_X1 U114 ( .B1(n487), .B2(n712), .A(n709), .ZN(n547) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n460), .ZN(n709) );
  OAI21_X1 U116 ( .B1(n486), .B2(n712), .A(n708), .ZN(n546) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n460), .ZN(n708) );
  OAI21_X1 U118 ( .B1(n485), .B2(n460), .A(n707), .ZN(n545) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n460), .ZN(n707) );
  OAI21_X1 U120 ( .B1(n484), .B2(n712), .A(n706), .ZN(n544) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n460), .ZN(n706) );
  OAI21_X1 U122 ( .B1(n483), .B2(n712), .A(n705), .ZN(n543) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n460), .ZN(n705) );
  OAI21_X1 U124 ( .B1(n482), .B2(n712), .A(n704), .ZN(n542) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n460), .ZN(n704) );
  OAI21_X1 U126 ( .B1(n481), .B2(n712), .A(n703), .ZN(n541) );
  NAND2_X1 U127 ( .A1(\mem[5][8] ), .A2(n460), .ZN(n703) );
  OAI21_X1 U128 ( .B1(n480), .B2(n712), .A(n702), .ZN(n540) );
  NAND2_X1 U129 ( .A1(\mem[5][9] ), .A2(n460), .ZN(n702) );
  OAI21_X1 U130 ( .B1(n479), .B2(n712), .A(n701), .ZN(n539) );
  NAND2_X1 U131 ( .A1(\mem[5][10] ), .A2(n460), .ZN(n701) );
  OAI21_X1 U132 ( .B1(n478), .B2(n712), .A(n700), .ZN(n538) );
  NAND2_X1 U133 ( .A1(\mem[5][11] ), .A2(n460), .ZN(n700) );
  OAI21_X1 U134 ( .B1(n477), .B2(n712), .A(n699), .ZN(n537) );
  NAND2_X1 U135 ( .A1(\mem[5][12] ), .A2(n712), .ZN(n699) );
  OAI21_X1 U136 ( .B1(n476), .B2(n460), .A(n698), .ZN(n536) );
  NAND2_X1 U137 ( .A1(\mem[5][13] ), .A2(n712), .ZN(n698) );
  OAI21_X1 U138 ( .B1(n475), .B2(n460), .A(n697), .ZN(n535) );
  NAND2_X1 U139 ( .A1(\mem[5][14] ), .A2(n712), .ZN(n697) );
  OAI21_X1 U140 ( .B1(n474), .B2(n712), .A(n696), .ZN(n534) );
  NAND2_X1 U141 ( .A1(\mem[5][15] ), .A2(n712), .ZN(n696) );
  OAI21_X1 U142 ( .B1(n473), .B2(n712), .A(n695), .ZN(n533) );
  NAND2_X1 U143 ( .A1(\mem[5][16] ), .A2(n712), .ZN(n695) );
  OAI21_X1 U144 ( .B1(n472), .B2(n712), .A(n694), .ZN(n532) );
  NAND2_X1 U145 ( .A1(\mem[5][17] ), .A2(n712), .ZN(n694) );
  OAI21_X1 U146 ( .B1(n471), .B2(n712), .A(n693), .ZN(n531) );
  NAND2_X1 U147 ( .A1(\mem[5][18] ), .A2(n712), .ZN(n693) );
  OAI21_X1 U148 ( .B1(n470), .B2(n712), .A(n692), .ZN(n530) );
  NAND2_X1 U149 ( .A1(\mem[5][19] ), .A2(n460), .ZN(n692) );
  OAI21_X1 U150 ( .B1(n489), .B2(n691), .A(n690), .ZN(n529) );
  NAND2_X1 U151 ( .A1(\mem[6][0] ), .A2(n459), .ZN(n690) );
  OAI21_X1 U152 ( .B1(n488), .B2(n691), .A(n689), .ZN(n528) );
  NAND2_X1 U153 ( .A1(\mem[6][1] ), .A2(n459), .ZN(n689) );
  OAI21_X1 U154 ( .B1(n487), .B2(n691), .A(n688), .ZN(n527) );
  NAND2_X1 U155 ( .A1(\mem[6][2] ), .A2(n459), .ZN(n688) );
  OAI21_X1 U156 ( .B1(n486), .B2(n691), .A(n687), .ZN(n526) );
  NAND2_X1 U157 ( .A1(\mem[6][3] ), .A2(n459), .ZN(n687) );
  OAI21_X1 U158 ( .B1(n485), .B2(n459), .A(n686), .ZN(n525) );
  NAND2_X1 U159 ( .A1(\mem[6][4] ), .A2(n459), .ZN(n686) );
  OAI21_X1 U160 ( .B1(n484), .B2(n691), .A(n685), .ZN(n524) );
  NAND2_X1 U161 ( .A1(\mem[6][5] ), .A2(n459), .ZN(n685) );
  OAI21_X1 U162 ( .B1(n483), .B2(n691), .A(n684), .ZN(n523) );
  NAND2_X1 U163 ( .A1(\mem[6][6] ), .A2(n459), .ZN(n684) );
  OAI21_X1 U164 ( .B1(n482), .B2(n691), .A(n683), .ZN(n522) );
  NAND2_X1 U165 ( .A1(\mem[6][7] ), .A2(n459), .ZN(n683) );
  OAI21_X1 U166 ( .B1(n481), .B2(n691), .A(n682), .ZN(n521) );
  NAND2_X1 U167 ( .A1(\mem[6][8] ), .A2(n459), .ZN(n682) );
  OAI21_X1 U168 ( .B1(n480), .B2(n691), .A(n681), .ZN(n520) );
  NAND2_X1 U169 ( .A1(\mem[6][9] ), .A2(n459), .ZN(n681) );
  OAI21_X1 U170 ( .B1(n479), .B2(n691), .A(n680), .ZN(n519) );
  NAND2_X1 U171 ( .A1(\mem[6][10] ), .A2(n459), .ZN(n680) );
  OAI21_X1 U172 ( .B1(n478), .B2(n691), .A(n679), .ZN(n518) );
  NAND2_X1 U173 ( .A1(\mem[6][11] ), .A2(n459), .ZN(n679) );
  OAI21_X1 U174 ( .B1(n477), .B2(n691), .A(n678), .ZN(n517) );
  NAND2_X1 U175 ( .A1(\mem[6][12] ), .A2(n691), .ZN(n678) );
  OAI21_X1 U176 ( .B1(n476), .B2(n459), .A(n677), .ZN(n516) );
  NAND2_X1 U177 ( .A1(\mem[6][13] ), .A2(n691), .ZN(n677) );
  OAI21_X1 U178 ( .B1(n475), .B2(n459), .A(n676), .ZN(n515) );
  NAND2_X1 U179 ( .A1(\mem[6][14] ), .A2(n691), .ZN(n676) );
  OAI21_X1 U180 ( .B1(n474), .B2(n691), .A(n675), .ZN(n514) );
  NAND2_X1 U181 ( .A1(\mem[6][15] ), .A2(n691), .ZN(n675) );
  OAI21_X1 U182 ( .B1(n473), .B2(n691), .A(n674), .ZN(n513) );
  NAND2_X1 U183 ( .A1(\mem[6][16] ), .A2(n691), .ZN(n674) );
  OAI21_X1 U184 ( .B1(n472), .B2(n691), .A(n673), .ZN(n512) );
  NAND2_X1 U185 ( .A1(\mem[6][17] ), .A2(n691), .ZN(n673) );
  OAI21_X1 U186 ( .B1(n471), .B2(n691), .A(n672), .ZN(n511) );
  NAND2_X1 U187 ( .A1(\mem[6][18] ), .A2(n691), .ZN(n672) );
  OAI21_X1 U188 ( .B1(n470), .B2(n691), .A(n671), .ZN(n510) );
  NAND2_X1 U189 ( .A1(\mem[6][19] ), .A2(n459), .ZN(n671) );
  OAI21_X1 U190 ( .B1(n489), .B2(n458), .A(n669), .ZN(n509) );
  NAND2_X1 U191 ( .A1(\mem[7][0] ), .A2(n458), .ZN(n669) );
  OAI21_X1 U192 ( .B1(n488), .B2(n458), .A(n668), .ZN(n508) );
  NAND2_X1 U193 ( .A1(\mem[7][1] ), .A2(n458), .ZN(n668) );
  OAI21_X1 U194 ( .B1(n487), .B2(n458), .A(n667), .ZN(n507) );
  NAND2_X1 U195 ( .A1(\mem[7][2] ), .A2(n670), .ZN(n667) );
  OAI21_X1 U196 ( .B1(n486), .B2(n670), .A(n666), .ZN(n506) );
  NAND2_X1 U197 ( .A1(\mem[7][3] ), .A2(n458), .ZN(n666) );
  OAI21_X1 U198 ( .B1(n485), .B2(n670), .A(n665), .ZN(n505) );
  NAND2_X1 U199 ( .A1(\mem[7][4] ), .A2(n670), .ZN(n665) );
  OAI21_X1 U200 ( .B1(n484), .B2(n670), .A(n664), .ZN(n504) );
  NAND2_X1 U201 ( .A1(\mem[7][5] ), .A2(n670), .ZN(n664) );
  OAI21_X1 U202 ( .B1(n483), .B2(n670), .A(n663), .ZN(n503) );
  NAND2_X1 U203 ( .A1(\mem[7][6] ), .A2(n670), .ZN(n663) );
  OAI21_X1 U204 ( .B1(n482), .B2(n670), .A(n662), .ZN(n502) );
  NAND2_X1 U205 ( .A1(\mem[7][7] ), .A2(n670), .ZN(n662) );
  OAI21_X1 U206 ( .B1(n481), .B2(n670), .A(n661), .ZN(n501) );
  NAND2_X1 U207 ( .A1(\mem[7][8] ), .A2(n670), .ZN(n661) );
  OAI21_X1 U208 ( .B1(n480), .B2(n458), .A(n660), .ZN(n500) );
  NAND2_X1 U209 ( .A1(\mem[7][9] ), .A2(n670), .ZN(n660) );
  OAI21_X1 U210 ( .B1(n479), .B2(n670), .A(n659), .ZN(n499) );
  NAND2_X1 U211 ( .A1(\mem[7][10] ), .A2(n670), .ZN(n659) );
  OAI21_X1 U212 ( .B1(n478), .B2(n670), .A(n658), .ZN(n498) );
  NAND2_X1 U213 ( .A1(\mem[7][11] ), .A2(n670), .ZN(n658) );
  OAI21_X1 U214 ( .B1(n477), .B2(n458), .A(n657), .ZN(n497) );
  NAND2_X1 U215 ( .A1(\mem[7][12] ), .A2(n458), .ZN(n657) );
  OAI21_X1 U216 ( .B1(n476), .B2(n458), .A(n656), .ZN(n496) );
  NAND2_X1 U217 ( .A1(\mem[7][13] ), .A2(n458), .ZN(n656) );
  OAI21_X1 U218 ( .B1(n475), .B2(n458), .A(n655), .ZN(n495) );
  NAND2_X1 U219 ( .A1(\mem[7][14] ), .A2(n458), .ZN(n655) );
  OAI21_X1 U220 ( .B1(n474), .B2(n670), .A(n654), .ZN(n494) );
  NAND2_X1 U221 ( .A1(\mem[7][15] ), .A2(n458), .ZN(n654) );
  OAI21_X1 U222 ( .B1(n473), .B2(n670), .A(n653), .ZN(n493) );
  NAND2_X1 U223 ( .A1(\mem[7][16] ), .A2(n458), .ZN(n653) );
  OAI21_X1 U224 ( .B1(n472), .B2(n670), .A(n652), .ZN(n492) );
  NAND2_X1 U225 ( .A1(\mem[7][17] ), .A2(n458), .ZN(n652) );
  OAI21_X1 U226 ( .B1(n471), .B2(n458), .A(n651), .ZN(n491) );
  NAND2_X1 U227 ( .A1(\mem[7][18] ), .A2(n458), .ZN(n651) );
  OAI21_X1 U228 ( .B1(n470), .B2(n458), .A(n650), .ZN(n490) );
  NAND2_X1 U229 ( .A1(\mem[7][19] ), .A2(n458), .ZN(n650) );
  NAND2_X1 U230 ( .A1(wr_en), .A2(n469), .ZN(n735) );
  INV_X1 U231 ( .A(addr[3]), .ZN(n469) );
  OAI21_X1 U232 ( .B1(n465), .B2(n489), .A(n819), .ZN(n649) );
  NAND2_X1 U233 ( .A1(\mem[0][0] ), .A2(n465), .ZN(n819) );
  OAI21_X1 U234 ( .B1(n820), .B2(n488), .A(n818), .ZN(n648) );
  NAND2_X1 U235 ( .A1(\mem[0][1] ), .A2(n465), .ZN(n818) );
  OAI21_X1 U236 ( .B1(n820), .B2(n487), .A(n817), .ZN(n647) );
  NAND2_X1 U237 ( .A1(\mem[0][2] ), .A2(n465), .ZN(n817) );
  OAI21_X1 U238 ( .B1(n820), .B2(n486), .A(n816), .ZN(n646) );
  NAND2_X1 U239 ( .A1(\mem[0][3] ), .A2(n465), .ZN(n816) );
  OAI21_X1 U240 ( .B1(n820), .B2(n485), .A(n815), .ZN(n645) );
  NAND2_X1 U241 ( .A1(\mem[0][4] ), .A2(n465), .ZN(n815) );
  OAI21_X1 U242 ( .B1(n820), .B2(n484), .A(n814), .ZN(n644) );
  NAND2_X1 U243 ( .A1(\mem[0][5] ), .A2(n465), .ZN(n814) );
  OAI21_X1 U244 ( .B1(n820), .B2(n483), .A(n813), .ZN(n643) );
  NAND2_X1 U245 ( .A1(\mem[0][6] ), .A2(n465), .ZN(n813) );
  OAI21_X1 U246 ( .B1(n820), .B2(n482), .A(n812), .ZN(n642) );
  NAND2_X1 U247 ( .A1(\mem[0][7] ), .A2(n465), .ZN(n812) );
  OAI21_X1 U248 ( .B1(n820), .B2(n481), .A(n811), .ZN(n641) );
  NAND2_X1 U249 ( .A1(\mem[0][8] ), .A2(n465), .ZN(n811) );
  OAI21_X1 U250 ( .B1(n820), .B2(n480), .A(n810), .ZN(n640) );
  NAND2_X1 U251 ( .A1(\mem[0][9] ), .A2(n465), .ZN(n810) );
  OAI21_X1 U252 ( .B1(n820), .B2(n479), .A(n809), .ZN(n639) );
  NAND2_X1 U253 ( .A1(\mem[0][10] ), .A2(n465), .ZN(n809) );
  OAI21_X1 U254 ( .B1(n820), .B2(n478), .A(n808), .ZN(n638) );
  NAND2_X1 U255 ( .A1(\mem[0][11] ), .A2(n465), .ZN(n808) );
  OAI21_X1 U256 ( .B1(n489), .B2(n464), .A(n797), .ZN(n629) );
  NAND2_X1 U257 ( .A1(\mem[1][0] ), .A2(n798), .ZN(n797) );
  OAI21_X1 U258 ( .B1(n488), .B2(n464), .A(n796), .ZN(n628) );
  NAND2_X1 U259 ( .A1(\mem[1][1] ), .A2(n798), .ZN(n796) );
  OAI21_X1 U260 ( .B1(n487), .B2(n464), .A(n795), .ZN(n627) );
  NAND2_X1 U261 ( .A1(\mem[1][2] ), .A2(n798), .ZN(n795) );
  OAI21_X1 U262 ( .B1(n486), .B2(n464), .A(n794), .ZN(n626) );
  NAND2_X1 U263 ( .A1(\mem[1][3] ), .A2(n798), .ZN(n794) );
  OAI21_X1 U264 ( .B1(n485), .B2(n464), .A(n793), .ZN(n625) );
  NAND2_X1 U265 ( .A1(\mem[1][4] ), .A2(n798), .ZN(n793) );
  OAI21_X1 U266 ( .B1(n484), .B2(n464), .A(n792), .ZN(n624) );
  NAND2_X1 U267 ( .A1(\mem[1][5] ), .A2(n798), .ZN(n792) );
  OAI21_X1 U268 ( .B1(n483), .B2(n464), .A(n791), .ZN(n623) );
  NAND2_X1 U269 ( .A1(\mem[1][6] ), .A2(n798), .ZN(n791) );
  OAI21_X1 U270 ( .B1(n482), .B2(n464), .A(n790), .ZN(n622) );
  NAND2_X1 U271 ( .A1(\mem[1][7] ), .A2(n798), .ZN(n790) );
  OAI21_X1 U272 ( .B1(n481), .B2(n464), .A(n789), .ZN(n621) );
  NAND2_X1 U273 ( .A1(\mem[1][8] ), .A2(n798), .ZN(n789) );
  OAI21_X1 U274 ( .B1(n480), .B2(n798), .A(n788), .ZN(n620) );
  NAND2_X1 U275 ( .A1(\mem[1][9] ), .A2(n798), .ZN(n788) );
  OAI21_X1 U276 ( .B1(n479), .B2(n464), .A(n787), .ZN(n619) );
  NAND2_X1 U277 ( .A1(\mem[1][10] ), .A2(n798), .ZN(n787) );
  OAI21_X1 U278 ( .B1(n478), .B2(n464), .A(n786), .ZN(n618) );
  NAND2_X1 U279 ( .A1(\mem[1][11] ), .A2(n798), .ZN(n786) );
  OAI21_X1 U280 ( .B1(n489), .B2(n777), .A(n776), .ZN(n609) );
  NAND2_X1 U281 ( .A1(\mem[2][0] ), .A2(n463), .ZN(n776) );
  OAI21_X1 U282 ( .B1(n488), .B2(n777), .A(n775), .ZN(n608) );
  NAND2_X1 U283 ( .A1(\mem[2][1] ), .A2(n463), .ZN(n775) );
  OAI21_X1 U284 ( .B1(n487), .B2(n777), .A(n774), .ZN(n607) );
  NAND2_X1 U285 ( .A1(\mem[2][2] ), .A2(n463), .ZN(n774) );
  OAI21_X1 U286 ( .B1(n486), .B2(n777), .A(n773), .ZN(n606) );
  NAND2_X1 U287 ( .A1(\mem[2][3] ), .A2(n463), .ZN(n773) );
  OAI21_X1 U288 ( .B1(n485), .B2(n777), .A(n772), .ZN(n605) );
  NAND2_X1 U289 ( .A1(\mem[2][4] ), .A2(n463), .ZN(n772) );
  OAI21_X1 U290 ( .B1(n484), .B2(n777), .A(n771), .ZN(n604) );
  NAND2_X1 U291 ( .A1(\mem[2][5] ), .A2(n463), .ZN(n771) );
  OAI21_X1 U292 ( .B1(n483), .B2(n777), .A(n770), .ZN(n603) );
  NAND2_X1 U293 ( .A1(\mem[2][6] ), .A2(n463), .ZN(n770) );
  OAI21_X1 U294 ( .B1(n482), .B2(n777), .A(n769), .ZN(n602) );
  NAND2_X1 U295 ( .A1(\mem[2][7] ), .A2(n463), .ZN(n769) );
  OAI21_X1 U296 ( .B1(n481), .B2(n777), .A(n768), .ZN(n601) );
  NAND2_X1 U297 ( .A1(\mem[2][8] ), .A2(n463), .ZN(n768) );
  OAI21_X1 U298 ( .B1(n480), .B2(n463), .A(n767), .ZN(n600) );
  NAND2_X1 U299 ( .A1(\mem[2][9] ), .A2(n463), .ZN(n767) );
  OAI21_X1 U300 ( .B1(n479), .B2(n777), .A(n766), .ZN(n599) );
  NAND2_X1 U301 ( .A1(\mem[2][10] ), .A2(n463), .ZN(n766) );
  OAI21_X1 U302 ( .B1(n478), .B2(n777), .A(n765), .ZN(n598) );
  NAND2_X1 U303 ( .A1(\mem[2][11] ), .A2(n463), .ZN(n765) );
  OAI21_X1 U304 ( .B1(n489), .B2(n756), .A(n755), .ZN(n589) );
  NAND2_X1 U305 ( .A1(\mem[3][0] ), .A2(n462), .ZN(n755) );
  OAI21_X1 U306 ( .B1(n488), .B2(n756), .A(n754), .ZN(n588) );
  NAND2_X1 U307 ( .A1(\mem[3][1] ), .A2(n462), .ZN(n754) );
  OAI21_X1 U308 ( .B1(n487), .B2(n756), .A(n753), .ZN(n587) );
  NAND2_X1 U309 ( .A1(\mem[3][2] ), .A2(n462), .ZN(n753) );
  OAI21_X1 U310 ( .B1(n486), .B2(n756), .A(n752), .ZN(n586) );
  NAND2_X1 U311 ( .A1(\mem[3][3] ), .A2(n462), .ZN(n752) );
  OAI21_X1 U312 ( .B1(n485), .B2(n756), .A(n751), .ZN(n585) );
  NAND2_X1 U313 ( .A1(\mem[3][4] ), .A2(n462), .ZN(n751) );
  OAI21_X1 U314 ( .B1(n484), .B2(n756), .A(n750), .ZN(n584) );
  NAND2_X1 U315 ( .A1(\mem[3][5] ), .A2(n462), .ZN(n750) );
  OAI21_X1 U316 ( .B1(n483), .B2(n756), .A(n749), .ZN(n583) );
  NAND2_X1 U317 ( .A1(\mem[3][6] ), .A2(n462), .ZN(n749) );
  OAI21_X1 U318 ( .B1(n482), .B2(n756), .A(n748), .ZN(n582) );
  NAND2_X1 U319 ( .A1(\mem[3][7] ), .A2(n462), .ZN(n748) );
  OAI21_X1 U320 ( .B1(n481), .B2(n756), .A(n747), .ZN(n581) );
  NAND2_X1 U321 ( .A1(\mem[3][8] ), .A2(n462), .ZN(n747) );
  OAI21_X1 U322 ( .B1(n480), .B2(n462), .A(n746), .ZN(n580) );
  NAND2_X1 U323 ( .A1(\mem[3][9] ), .A2(n462), .ZN(n746) );
  OAI21_X1 U324 ( .B1(n479), .B2(n756), .A(n745), .ZN(n579) );
  NAND2_X1 U325 ( .A1(\mem[3][10] ), .A2(n462), .ZN(n745) );
  OAI21_X1 U326 ( .B1(n478), .B2(n756), .A(n744), .ZN(n578) );
  NAND2_X1 U327 ( .A1(\mem[3][11] ), .A2(n462), .ZN(n744) );
  OAI21_X1 U328 ( .B1(n820), .B2(n477), .A(n807), .ZN(n637) );
  NAND2_X1 U329 ( .A1(\mem[0][12] ), .A2(n820), .ZN(n807) );
  OAI21_X1 U330 ( .B1(n820), .B2(n476), .A(n806), .ZN(n636) );
  NAND2_X1 U331 ( .A1(\mem[0][13] ), .A2(n820), .ZN(n806) );
  OAI21_X1 U332 ( .B1(n465), .B2(n475), .A(n805), .ZN(n635) );
  NAND2_X1 U333 ( .A1(\mem[0][14] ), .A2(n820), .ZN(n805) );
  OAI21_X1 U334 ( .B1(n820), .B2(n474), .A(n804), .ZN(n634) );
  NAND2_X1 U335 ( .A1(\mem[0][15] ), .A2(n465), .ZN(n804) );
  OAI21_X1 U336 ( .B1(n820), .B2(n473), .A(n803), .ZN(n633) );
  NAND2_X1 U337 ( .A1(\mem[0][16] ), .A2(n820), .ZN(n803) );
  OAI21_X1 U338 ( .B1(n820), .B2(n472), .A(n802), .ZN(n632) );
  NAND2_X1 U339 ( .A1(\mem[0][17] ), .A2(n820), .ZN(n802) );
  OAI21_X1 U340 ( .B1(n820), .B2(n471), .A(n801), .ZN(n631) );
  NAND2_X1 U341 ( .A1(\mem[0][18] ), .A2(n820), .ZN(n801) );
  OAI21_X1 U342 ( .B1(n820), .B2(n470), .A(n800), .ZN(n630) );
  NAND2_X1 U343 ( .A1(\mem[0][19] ), .A2(n465), .ZN(n800) );
  INV_X1 U344 ( .A(data_in[0]), .ZN(n489) );
  INV_X1 U345 ( .A(data_in[1]), .ZN(n488) );
  INV_X1 U346 ( .A(data_in[2]), .ZN(n487) );
  INV_X1 U347 ( .A(data_in[3]), .ZN(n486) );
  INV_X1 U348 ( .A(data_in[4]), .ZN(n485) );
  INV_X1 U349 ( .A(data_in[5]), .ZN(n484) );
  INV_X1 U358 ( .A(data_in[6]), .ZN(n483) );
  INV_X1 U359 ( .A(data_in[7]), .ZN(n482) );
  INV_X1 U360 ( .A(data_in[8]), .ZN(n481) );
  INV_X1 U361 ( .A(data_in[9]), .ZN(n480) );
  INV_X1 U362 ( .A(data_in[10]), .ZN(n479) );
  INV_X1 U363 ( .A(data_in[11]), .ZN(n478) );
  INV_X1 U364 ( .A(data_in[12]), .ZN(n477) );
  INV_X1 U365 ( .A(data_in[13]), .ZN(n476) );
  INV_X1 U366 ( .A(data_in[14]), .ZN(n475) );
  INV_X1 U367 ( .A(data_in[15]), .ZN(n474) );
  INV_X1 U368 ( .A(data_in[16]), .ZN(n473) );
  INV_X1 U369 ( .A(data_in[17]), .ZN(n472) );
  INV_X1 U370 ( .A(data_in[18]), .ZN(n471) );
  INV_X1 U371 ( .A(data_in[19]), .ZN(n470) );
  MUX2_X1 U372 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n456), .Z(n1) );
  MUX2_X1 U373 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n457), .Z(n2) );
  MUX2_X1 U374 ( .A(n2), .B(n1), .S(n453), .Z(n3) );
  MUX2_X1 U375 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n457), .Z(n4) );
  MUX2_X1 U376 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n454), .Z(n5) );
  MUX2_X1 U377 ( .A(n5), .B(n4), .S(n453), .Z(n6) );
  MUX2_X1 U378 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n457), .Z(n7) );
  MUX2_X1 U379 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n454), .Z(n8) );
  MUX2_X1 U380 ( .A(n8), .B(n7), .S(n453), .Z(n9) );
  MUX2_X1 U381 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n455), .Z(n10) );
  MUX2_X1 U382 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n456), .Z(n11) );
  MUX2_X1 U383 ( .A(n11), .B(n10), .S(n453), .Z(n12) );
  MUX2_X1 U384 ( .A(n12), .B(n9), .S(N12), .Z(N31) );
  MUX2_X1 U385 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n454), .Z(n13) );
  MUX2_X1 U386 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n454), .Z(n14) );
  MUX2_X1 U387 ( .A(n14), .B(n13), .S(n453), .Z(n15) );
  MUX2_X1 U388 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n454), .Z(n16) );
  MUX2_X1 U389 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n454), .Z(n17) );
  MUX2_X1 U390 ( .A(n17), .B(n16), .S(n453), .Z(n18) );
  MUX2_X1 U391 ( .A(n18), .B(n15), .S(N12), .Z(N30) );
  MUX2_X1 U392 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n454), .Z(n19) );
  MUX2_X1 U393 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n454), .Z(n20) );
  MUX2_X1 U394 ( .A(n20), .B(n19), .S(n453), .Z(n21) );
  MUX2_X1 U395 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n454), .Z(n22) );
  MUX2_X1 U396 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n454), .Z(n23) );
  MUX2_X1 U397 ( .A(n23), .B(n22), .S(n453), .Z(n24) );
  MUX2_X1 U398 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n454), .Z(n356) );
  MUX2_X1 U399 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n454), .Z(n357) );
  MUX2_X1 U400 ( .A(n357), .B(n356), .S(n453), .Z(n358) );
  MUX2_X1 U401 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n454), .Z(n359) );
  MUX2_X1 U402 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n454), .Z(n360) );
  MUX2_X1 U403 ( .A(n360), .B(n359), .S(n453), .Z(n361) );
  MUX2_X1 U404 ( .A(n361), .B(n358), .S(N12), .Z(N28) );
  MUX2_X1 U405 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n456), .Z(n362) );
  MUX2_X1 U406 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n456), .Z(n363) );
  MUX2_X1 U407 ( .A(n363), .B(n362), .S(n453), .Z(n364) );
  MUX2_X1 U408 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n454), .Z(n365) );
  MUX2_X1 U409 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n455), .Z(n366) );
  MUX2_X1 U410 ( .A(n366), .B(n365), .S(n453), .Z(n367) );
  MUX2_X1 U411 ( .A(n367), .B(n364), .S(N12), .Z(N27) );
  MUX2_X1 U412 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n457), .Z(n368) );
  MUX2_X1 U413 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n457), .Z(n369) );
  MUX2_X1 U414 ( .A(n369), .B(n368), .S(n453), .Z(n370) );
  MUX2_X1 U415 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n455), .Z(n371) );
  MUX2_X1 U416 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n456), .Z(n372) );
  MUX2_X1 U417 ( .A(n372), .B(n371), .S(n453), .Z(n373) );
  MUX2_X1 U418 ( .A(n373), .B(n370), .S(N12), .Z(N26) );
  MUX2_X1 U419 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n454), .Z(n374) );
  MUX2_X1 U420 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n455), .Z(n375) );
  MUX2_X1 U421 ( .A(n375), .B(n374), .S(n453), .Z(n376) );
  MUX2_X1 U422 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n457), .Z(n377) );
  MUX2_X1 U423 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n455), .Z(n378) );
  MUX2_X1 U424 ( .A(n378), .B(n377), .S(n453), .Z(n379) );
  MUX2_X1 U425 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n455), .Z(n380) );
  MUX2_X1 U426 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n454), .Z(n381) );
  MUX2_X1 U427 ( .A(n381), .B(n380), .S(n453), .Z(n382) );
  MUX2_X1 U428 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n455), .Z(n383) );
  MUX2_X1 U429 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n455), .Z(n384) );
  MUX2_X1 U430 ( .A(n384), .B(n383), .S(n453), .Z(n385) );
  MUX2_X1 U431 ( .A(n385), .B(n382), .S(N12), .Z(N24) );
  MUX2_X1 U432 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n454), .Z(n386) );
  MUX2_X1 U433 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n454), .Z(n387) );
  MUX2_X1 U434 ( .A(n387), .B(n386), .S(n453), .Z(n388) );
  MUX2_X1 U435 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n456), .Z(n389) );
  MUX2_X1 U436 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n456), .Z(n390) );
  MUX2_X1 U437 ( .A(n390), .B(n389), .S(n453), .Z(n391) );
  MUX2_X1 U438 ( .A(n391), .B(n388), .S(N12), .Z(N23) );
  MUX2_X1 U439 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n456), .Z(n392) );
  MUX2_X1 U440 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n454), .Z(n393) );
  MUX2_X1 U441 ( .A(n393), .B(n392), .S(n453), .Z(n394) );
  MUX2_X1 U442 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n457), .Z(n395) );
  MUX2_X1 U443 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n457), .Z(n396) );
  MUX2_X1 U444 ( .A(n396), .B(n395), .S(N11), .Z(n397) );
  MUX2_X1 U445 ( .A(n397), .B(n394), .S(N12), .Z(N22) );
  MUX2_X1 U446 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n455), .Z(n398) );
  MUX2_X1 U447 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n455), .Z(n399) );
  MUX2_X1 U448 ( .A(n399), .B(n398), .S(N11), .Z(n400) );
  MUX2_X1 U449 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n455), .Z(n401) );
  MUX2_X1 U450 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n455), .Z(n402) );
  MUX2_X1 U451 ( .A(n402), .B(n401), .S(N11), .Z(n403) );
  MUX2_X1 U452 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n455), .Z(n404) );
  MUX2_X1 U453 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n455), .Z(n405) );
  MUX2_X1 U454 ( .A(n405), .B(n404), .S(n453), .Z(n406) );
  MUX2_X1 U455 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n455), .Z(n407) );
  MUX2_X1 U456 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n455), .Z(n408) );
  MUX2_X1 U457 ( .A(n408), .B(n407), .S(N11), .Z(n409) );
  MUX2_X1 U458 ( .A(n409), .B(n406), .S(N12), .Z(N20) );
  MUX2_X1 U459 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n455), .Z(n410) );
  MUX2_X1 U460 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n455), .Z(n411) );
  MUX2_X1 U461 ( .A(n411), .B(n410), .S(N11), .Z(n412) );
  MUX2_X1 U462 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n455), .Z(n413) );
  MUX2_X1 U463 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n455), .Z(n414) );
  MUX2_X1 U464 ( .A(n414), .B(n413), .S(N11), .Z(n415) );
  MUX2_X1 U465 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n456), .Z(n416) );
  MUX2_X1 U466 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n456), .Z(n417) );
  MUX2_X1 U467 ( .A(n417), .B(n416), .S(n452), .Z(n418) );
  MUX2_X1 U468 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n456), .Z(n419) );
  MUX2_X1 U469 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n456), .Z(n420) );
  MUX2_X1 U470 ( .A(n420), .B(n419), .S(n452), .Z(n421) );
  MUX2_X1 U471 ( .A(n421), .B(n418), .S(N12), .Z(N18) );
  MUX2_X1 U472 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n456), .Z(n422) );
  MUX2_X1 U473 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n456), .Z(n423) );
  MUX2_X1 U474 ( .A(n423), .B(n422), .S(n452), .Z(n424) );
  MUX2_X1 U475 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n456), .Z(n425) );
  MUX2_X1 U476 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n456), .Z(n426) );
  MUX2_X1 U477 ( .A(n426), .B(n425), .S(n452), .Z(n427) );
  MUX2_X1 U478 ( .A(n427), .B(n424), .S(N12), .Z(N17) );
  MUX2_X1 U479 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n456), .Z(n428) );
  MUX2_X1 U480 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n456), .Z(n429) );
  MUX2_X1 U481 ( .A(n429), .B(n428), .S(n452), .Z(n430) );
  MUX2_X1 U482 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n456), .Z(n431) );
  MUX2_X1 U483 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n456), .Z(n432) );
  MUX2_X1 U484 ( .A(n432), .B(n431), .S(n452), .Z(n433) );
  MUX2_X1 U485 ( .A(n433), .B(n430), .S(N12), .Z(N16) );
  MUX2_X1 U486 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n457), .Z(n434) );
  MUX2_X1 U487 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n457), .Z(n435) );
  MUX2_X1 U488 ( .A(n435), .B(n434), .S(n452), .Z(n436) );
  MUX2_X1 U489 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n457), .Z(n437) );
  MUX2_X1 U490 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n457), .Z(n438) );
  MUX2_X1 U491 ( .A(n438), .B(n437), .S(n452), .Z(n439) );
  MUX2_X1 U492 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n457), .Z(n440) );
  MUX2_X1 U493 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n457), .Z(n441) );
  MUX2_X1 U494 ( .A(n441), .B(n440), .S(n452), .Z(n442) );
  MUX2_X1 U495 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n457), .Z(n443) );
  MUX2_X1 U496 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n457), .Z(n444) );
  MUX2_X1 U497 ( .A(n444), .B(n443), .S(n452), .Z(n445) );
  MUX2_X1 U498 ( .A(n445), .B(n442), .S(N12), .Z(N14) );
  MUX2_X1 U499 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n457), .Z(n446) );
  MUX2_X1 U500 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n457), .Z(n447) );
  MUX2_X1 U501 ( .A(n447), .B(n446), .S(n452), .Z(n448) );
  MUX2_X1 U502 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n457), .Z(n449) );
  MUX2_X1 U503 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n457), .Z(n450) );
  MUX2_X1 U504 ( .A(n450), .B(n449), .S(n452), .Z(n451) );
  MUX2_X1 U505 ( .A(n451), .B(n448), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE4_3 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N13, N14, N16, N17, N18, N20, N22, N23, N24, N25, N26,
         N27, N28, N30, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[19]  ( .D(N13), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[15]  ( .D(N17), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N20), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N23), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N25), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N27), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N30), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N32), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n490), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n491), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n492), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n493), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n494), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n495), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n496), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n497), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n498), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n499), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n500), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n501), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n502), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n503), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n504), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n505), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n506), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n507), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n508), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n509), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n510), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n511), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n512), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n513), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n514), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n515), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n516), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n517), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n518), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n519), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n520), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n521), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n522), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n523), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n524), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n525), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n526), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n527), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n528), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n529), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n530), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n531), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n532), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n533), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n534), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n535), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n536), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n537), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n538), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n539), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n540), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n541), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n542), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n543), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n544), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n545), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n546), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n547), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n548), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n549), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n550), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n551), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n552), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n553), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n554), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n555), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n556), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n557), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n558), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n559), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n560), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n561), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n562), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n563), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n564), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n565), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n566), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n567), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n568), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n569), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n570), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n571), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n572), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n573), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n574), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n575), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n576), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n577), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n578), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n579), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n580), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n581), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n582), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n583), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n584), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n585), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n586), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n587), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n588), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n589), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n590), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n591), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n592), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n593), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n594), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n595), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n596), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n597), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n598), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n599), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n600), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n601), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n602), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n603), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n604), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n605), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n606), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n607), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n608), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n609), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n610), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n611), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n612), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n613), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n614), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n615), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n616), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n617), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n618), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n619), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n620), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n621), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n622), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n623), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n624), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n625), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n626), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n627), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n628), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n629), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n630), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n631), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n632), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n633), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n634), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n635), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n636), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n637), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n638), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n639), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n640), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n641), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n642), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n643), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n644), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n645), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n646), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n647), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n648), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n649), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U350 ( .A1(n466), .A2(n467), .A3(n799), .ZN(n820) );
  NAND3_X1 U351 ( .A1(n799), .A2(n467), .A3(N10), .ZN(n798) );
  NAND3_X1 U352 ( .A1(n799), .A2(n466), .A3(N11), .ZN(n777) );
  NAND3_X1 U353 ( .A1(N10), .A2(n799), .A3(N11), .ZN(n756) );
  NAND3_X1 U354 ( .A1(n466), .A2(n467), .A3(n713), .ZN(n734) );
  NAND3_X1 U355 ( .A1(N10), .A2(n467), .A3(n713), .ZN(n712) );
  NAND3_X1 U356 ( .A1(N11), .A2(n466), .A3(n713), .ZN(n691) );
  NAND3_X1 U357 ( .A1(N11), .A2(N10), .A3(n713), .ZN(n670) );
  SDFF_X1 \data_out_reg[17]  ( .D(n436), .SI(n439), .SE(n468), .CK(clk), .Q(
        data_out[17]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n400), .SI(n403), .SE(n468), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n412), .SI(n415), .SE(n468), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n9), .SI(n12), .SE(n468), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n21), .SI(n24), .SE(n468), .CK(clk), .Q(
        data_out[3]) );
  BUF_X1 U3 ( .A(n777), .Z(n463) );
  BUF_X1 U4 ( .A(n712), .Z(n460) );
  BUF_X1 U5 ( .A(n670), .Z(n458) );
  BUF_X1 U6 ( .A(n453), .Z(n452) );
  BUF_X1 U7 ( .A(N10), .Z(n454) );
  BUF_X1 U8 ( .A(N10), .Z(n455) );
  BUF_X1 U9 ( .A(N10), .Z(n456) );
  BUF_X1 U10 ( .A(N10), .Z(n457) );
  BUF_X1 U11 ( .A(N11), .Z(n453) );
  BUF_X1 U12 ( .A(n820), .Z(n465) );
  BUF_X1 U13 ( .A(n756), .Z(n462) );
  BUF_X1 U14 ( .A(n798), .Z(n464) );
  BUF_X1 U15 ( .A(n734), .Z(n461) );
  BUF_X1 U16 ( .A(n691), .Z(n459) );
  NOR2_X1 U17 ( .A1(n735), .A2(N12), .ZN(n799) );
  NOR2_X1 U18 ( .A1(n468), .A2(n735), .ZN(n713) );
  INV_X1 U19 ( .A(N12), .ZN(n468) );
  INV_X1 U20 ( .A(N11), .ZN(n467) );
  INV_X1 U21 ( .A(N10), .ZN(n466) );
  OAI21_X1 U22 ( .B1(n477), .B2(n798), .A(n785), .ZN(n617) );
  NAND2_X1 U23 ( .A1(\mem[1][12] ), .A2(n798), .ZN(n785) );
  OAI21_X1 U24 ( .B1(n476), .B2(n798), .A(n784), .ZN(n616) );
  NAND2_X1 U25 ( .A1(\mem[1][13] ), .A2(n798), .ZN(n784) );
  OAI21_X1 U26 ( .B1(n475), .B2(n798), .A(n783), .ZN(n615) );
  NAND2_X1 U27 ( .A1(\mem[1][14] ), .A2(n798), .ZN(n783) );
  OAI21_X1 U28 ( .B1(n474), .B2(n464), .A(n782), .ZN(n614) );
  NAND2_X1 U29 ( .A1(\mem[1][15] ), .A2(n798), .ZN(n782) );
  OAI21_X1 U30 ( .B1(n473), .B2(n798), .A(n781), .ZN(n613) );
  NAND2_X1 U31 ( .A1(\mem[1][16] ), .A2(n464), .ZN(n781) );
  OAI21_X1 U32 ( .B1(n472), .B2(n798), .A(n780), .ZN(n612) );
  NAND2_X1 U33 ( .A1(\mem[1][17] ), .A2(n798), .ZN(n780) );
  OAI21_X1 U34 ( .B1(n471), .B2(n798), .A(n779), .ZN(n611) );
  NAND2_X1 U35 ( .A1(\mem[1][18] ), .A2(n798), .ZN(n779) );
  OAI21_X1 U36 ( .B1(n470), .B2(n798), .A(n778), .ZN(n610) );
  NAND2_X1 U37 ( .A1(\mem[1][19] ), .A2(n464), .ZN(n778) );
  OAI21_X1 U38 ( .B1(n477), .B2(n463), .A(n764), .ZN(n597) );
  NAND2_X1 U39 ( .A1(\mem[2][12] ), .A2(n463), .ZN(n764) );
  OAI21_X1 U40 ( .B1(n476), .B2(n463), .A(n763), .ZN(n596) );
  NAND2_X1 U41 ( .A1(\mem[2][13] ), .A2(n463), .ZN(n763) );
  OAI21_X1 U42 ( .B1(n475), .B2(n463), .A(n762), .ZN(n595) );
  NAND2_X1 U43 ( .A1(\mem[2][14] ), .A2(n463), .ZN(n762) );
  OAI21_X1 U44 ( .B1(n474), .B2(n777), .A(n761), .ZN(n594) );
  NAND2_X1 U45 ( .A1(\mem[2][15] ), .A2(n463), .ZN(n761) );
  OAI21_X1 U46 ( .B1(n473), .B2(n777), .A(n760), .ZN(n593) );
  NAND2_X1 U47 ( .A1(\mem[2][16] ), .A2(n463), .ZN(n760) );
  OAI21_X1 U48 ( .B1(n472), .B2(n777), .A(n759), .ZN(n592) );
  NAND2_X1 U49 ( .A1(\mem[2][17] ), .A2(n463), .ZN(n759) );
  OAI21_X1 U50 ( .B1(n471), .B2(n777), .A(n758), .ZN(n591) );
  NAND2_X1 U51 ( .A1(\mem[2][18] ), .A2(n463), .ZN(n758) );
  OAI21_X1 U52 ( .B1(n470), .B2(n777), .A(n757), .ZN(n590) );
  NAND2_X1 U53 ( .A1(\mem[2][19] ), .A2(n463), .ZN(n757) );
  OAI21_X1 U54 ( .B1(n477), .B2(n756), .A(n743), .ZN(n577) );
  NAND2_X1 U55 ( .A1(\mem[3][12] ), .A2(n756), .ZN(n743) );
  OAI21_X1 U56 ( .B1(n476), .B2(n756), .A(n742), .ZN(n576) );
  NAND2_X1 U57 ( .A1(\mem[3][13] ), .A2(n756), .ZN(n742) );
  OAI21_X1 U58 ( .B1(n475), .B2(n756), .A(n741), .ZN(n575) );
  NAND2_X1 U59 ( .A1(\mem[3][14] ), .A2(n756), .ZN(n741) );
  OAI21_X1 U60 ( .B1(n474), .B2(n462), .A(n740), .ZN(n574) );
  NAND2_X1 U61 ( .A1(\mem[3][15] ), .A2(n756), .ZN(n740) );
  OAI21_X1 U62 ( .B1(n473), .B2(n756), .A(n739), .ZN(n573) );
  NAND2_X1 U63 ( .A1(\mem[3][16] ), .A2(n462), .ZN(n739) );
  OAI21_X1 U64 ( .B1(n472), .B2(n756), .A(n738), .ZN(n572) );
  NAND2_X1 U65 ( .A1(\mem[3][17] ), .A2(n756), .ZN(n738) );
  OAI21_X1 U66 ( .B1(n471), .B2(n756), .A(n737), .ZN(n571) );
  NAND2_X1 U67 ( .A1(\mem[3][18] ), .A2(n756), .ZN(n737) );
  OAI21_X1 U68 ( .B1(n470), .B2(n756), .A(n736), .ZN(n570) );
  NAND2_X1 U69 ( .A1(\mem[3][19] ), .A2(n462), .ZN(n736) );
  OAI21_X1 U70 ( .B1(n489), .B2(n734), .A(n733), .ZN(n569) );
  NAND2_X1 U71 ( .A1(\mem[4][0] ), .A2(n461), .ZN(n733) );
  OAI21_X1 U72 ( .B1(n488), .B2(n734), .A(n732), .ZN(n568) );
  NAND2_X1 U73 ( .A1(\mem[4][1] ), .A2(n461), .ZN(n732) );
  OAI21_X1 U74 ( .B1(n487), .B2(n734), .A(n731), .ZN(n567) );
  NAND2_X1 U75 ( .A1(\mem[4][2] ), .A2(n461), .ZN(n731) );
  OAI21_X1 U76 ( .B1(n486), .B2(n734), .A(n730), .ZN(n566) );
  NAND2_X1 U77 ( .A1(\mem[4][3] ), .A2(n461), .ZN(n730) );
  OAI21_X1 U78 ( .B1(n485), .B2(n461), .A(n729), .ZN(n565) );
  NAND2_X1 U79 ( .A1(\mem[4][4] ), .A2(n461), .ZN(n729) );
  OAI21_X1 U80 ( .B1(n484), .B2(n734), .A(n728), .ZN(n564) );
  NAND2_X1 U81 ( .A1(\mem[4][5] ), .A2(n461), .ZN(n728) );
  OAI21_X1 U82 ( .B1(n483), .B2(n734), .A(n727), .ZN(n563) );
  NAND2_X1 U83 ( .A1(\mem[4][6] ), .A2(n461), .ZN(n727) );
  OAI21_X1 U84 ( .B1(n482), .B2(n734), .A(n726), .ZN(n562) );
  NAND2_X1 U85 ( .A1(\mem[4][7] ), .A2(n461), .ZN(n726) );
  OAI21_X1 U86 ( .B1(n481), .B2(n734), .A(n725), .ZN(n561) );
  NAND2_X1 U87 ( .A1(\mem[4][8] ), .A2(n461), .ZN(n725) );
  OAI21_X1 U88 ( .B1(n480), .B2(n734), .A(n724), .ZN(n560) );
  NAND2_X1 U89 ( .A1(\mem[4][9] ), .A2(n461), .ZN(n724) );
  OAI21_X1 U90 ( .B1(n479), .B2(n734), .A(n723), .ZN(n559) );
  NAND2_X1 U91 ( .A1(\mem[4][10] ), .A2(n461), .ZN(n723) );
  OAI21_X1 U92 ( .B1(n478), .B2(n734), .A(n722), .ZN(n558) );
  NAND2_X1 U93 ( .A1(\mem[4][11] ), .A2(n461), .ZN(n722) );
  OAI21_X1 U94 ( .B1(n477), .B2(n734), .A(n721), .ZN(n557) );
  NAND2_X1 U95 ( .A1(\mem[4][12] ), .A2(n734), .ZN(n721) );
  OAI21_X1 U96 ( .B1(n476), .B2(n461), .A(n720), .ZN(n556) );
  NAND2_X1 U97 ( .A1(\mem[4][13] ), .A2(n734), .ZN(n720) );
  OAI21_X1 U98 ( .B1(n475), .B2(n461), .A(n719), .ZN(n555) );
  NAND2_X1 U99 ( .A1(\mem[4][14] ), .A2(n734), .ZN(n719) );
  OAI21_X1 U100 ( .B1(n474), .B2(n734), .A(n718), .ZN(n554) );
  NAND2_X1 U101 ( .A1(\mem[4][15] ), .A2(n734), .ZN(n718) );
  OAI21_X1 U102 ( .B1(n473), .B2(n734), .A(n717), .ZN(n553) );
  NAND2_X1 U103 ( .A1(\mem[4][16] ), .A2(n734), .ZN(n717) );
  OAI21_X1 U104 ( .B1(n472), .B2(n734), .A(n716), .ZN(n552) );
  NAND2_X1 U105 ( .A1(\mem[4][17] ), .A2(n734), .ZN(n716) );
  OAI21_X1 U106 ( .B1(n471), .B2(n734), .A(n715), .ZN(n551) );
  NAND2_X1 U107 ( .A1(\mem[4][18] ), .A2(n734), .ZN(n715) );
  OAI21_X1 U108 ( .B1(n470), .B2(n734), .A(n714), .ZN(n550) );
  NAND2_X1 U109 ( .A1(\mem[4][19] ), .A2(n461), .ZN(n714) );
  OAI21_X1 U110 ( .B1(n489), .B2(n460), .A(n711), .ZN(n549) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n460), .ZN(n711) );
  OAI21_X1 U112 ( .B1(n488), .B2(n460), .A(n710), .ZN(n548) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n460), .ZN(n710) );
  OAI21_X1 U114 ( .B1(n487), .B2(n460), .A(n709), .ZN(n547) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n712), .ZN(n709) );
  OAI21_X1 U116 ( .B1(n486), .B2(n712), .A(n708), .ZN(n546) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n460), .ZN(n708) );
  OAI21_X1 U118 ( .B1(n485), .B2(n712), .A(n707), .ZN(n545) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n712), .ZN(n707) );
  OAI21_X1 U120 ( .B1(n484), .B2(n712), .A(n706), .ZN(n544) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n712), .ZN(n706) );
  OAI21_X1 U122 ( .B1(n483), .B2(n712), .A(n705), .ZN(n543) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n712), .ZN(n705) );
  OAI21_X1 U124 ( .B1(n482), .B2(n712), .A(n704), .ZN(n542) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n712), .ZN(n704) );
  OAI21_X1 U126 ( .B1(n481), .B2(n712), .A(n703), .ZN(n541) );
  NAND2_X1 U127 ( .A1(\mem[5][8] ), .A2(n712), .ZN(n703) );
  OAI21_X1 U128 ( .B1(n480), .B2(n460), .A(n702), .ZN(n540) );
  NAND2_X1 U129 ( .A1(\mem[5][9] ), .A2(n712), .ZN(n702) );
  OAI21_X1 U130 ( .B1(n479), .B2(n712), .A(n701), .ZN(n539) );
  NAND2_X1 U131 ( .A1(\mem[5][10] ), .A2(n712), .ZN(n701) );
  OAI21_X1 U132 ( .B1(n478), .B2(n712), .A(n700), .ZN(n538) );
  NAND2_X1 U133 ( .A1(\mem[5][11] ), .A2(n712), .ZN(n700) );
  OAI21_X1 U134 ( .B1(n477), .B2(n460), .A(n699), .ZN(n537) );
  NAND2_X1 U135 ( .A1(\mem[5][12] ), .A2(n460), .ZN(n699) );
  OAI21_X1 U136 ( .B1(n476), .B2(n460), .A(n698), .ZN(n536) );
  NAND2_X1 U137 ( .A1(\mem[5][13] ), .A2(n460), .ZN(n698) );
  OAI21_X1 U138 ( .B1(n475), .B2(n460), .A(n697), .ZN(n535) );
  NAND2_X1 U139 ( .A1(\mem[5][14] ), .A2(n460), .ZN(n697) );
  OAI21_X1 U140 ( .B1(n474), .B2(n712), .A(n696), .ZN(n534) );
  NAND2_X1 U141 ( .A1(\mem[5][15] ), .A2(n460), .ZN(n696) );
  OAI21_X1 U142 ( .B1(n473), .B2(n712), .A(n695), .ZN(n533) );
  NAND2_X1 U143 ( .A1(\mem[5][16] ), .A2(n460), .ZN(n695) );
  OAI21_X1 U144 ( .B1(n472), .B2(n712), .A(n694), .ZN(n532) );
  NAND2_X1 U145 ( .A1(\mem[5][17] ), .A2(n460), .ZN(n694) );
  OAI21_X1 U146 ( .B1(n471), .B2(n460), .A(n693), .ZN(n531) );
  NAND2_X1 U147 ( .A1(\mem[5][18] ), .A2(n460), .ZN(n693) );
  OAI21_X1 U148 ( .B1(n470), .B2(n460), .A(n692), .ZN(n530) );
  NAND2_X1 U149 ( .A1(\mem[5][19] ), .A2(n460), .ZN(n692) );
  OAI21_X1 U150 ( .B1(n489), .B2(n691), .A(n690), .ZN(n529) );
  NAND2_X1 U151 ( .A1(\mem[6][0] ), .A2(n459), .ZN(n690) );
  OAI21_X1 U152 ( .B1(n488), .B2(n691), .A(n689), .ZN(n528) );
  NAND2_X1 U153 ( .A1(\mem[6][1] ), .A2(n459), .ZN(n689) );
  OAI21_X1 U154 ( .B1(n487), .B2(n691), .A(n688), .ZN(n527) );
  NAND2_X1 U155 ( .A1(\mem[6][2] ), .A2(n459), .ZN(n688) );
  OAI21_X1 U156 ( .B1(n486), .B2(n691), .A(n687), .ZN(n526) );
  NAND2_X1 U157 ( .A1(\mem[6][3] ), .A2(n459), .ZN(n687) );
  OAI21_X1 U158 ( .B1(n485), .B2(n459), .A(n686), .ZN(n525) );
  NAND2_X1 U159 ( .A1(\mem[6][4] ), .A2(n459), .ZN(n686) );
  OAI21_X1 U160 ( .B1(n484), .B2(n691), .A(n685), .ZN(n524) );
  NAND2_X1 U161 ( .A1(\mem[6][5] ), .A2(n459), .ZN(n685) );
  OAI21_X1 U162 ( .B1(n483), .B2(n691), .A(n684), .ZN(n523) );
  NAND2_X1 U163 ( .A1(\mem[6][6] ), .A2(n459), .ZN(n684) );
  OAI21_X1 U164 ( .B1(n482), .B2(n691), .A(n683), .ZN(n522) );
  NAND2_X1 U165 ( .A1(\mem[6][7] ), .A2(n459), .ZN(n683) );
  OAI21_X1 U166 ( .B1(n481), .B2(n691), .A(n682), .ZN(n521) );
  NAND2_X1 U167 ( .A1(\mem[6][8] ), .A2(n459), .ZN(n682) );
  OAI21_X1 U168 ( .B1(n480), .B2(n691), .A(n681), .ZN(n520) );
  NAND2_X1 U169 ( .A1(\mem[6][9] ), .A2(n459), .ZN(n681) );
  OAI21_X1 U170 ( .B1(n479), .B2(n691), .A(n680), .ZN(n519) );
  NAND2_X1 U171 ( .A1(\mem[6][10] ), .A2(n459), .ZN(n680) );
  OAI21_X1 U172 ( .B1(n478), .B2(n691), .A(n679), .ZN(n518) );
  NAND2_X1 U173 ( .A1(\mem[6][11] ), .A2(n459), .ZN(n679) );
  OAI21_X1 U174 ( .B1(n477), .B2(n691), .A(n678), .ZN(n517) );
  NAND2_X1 U175 ( .A1(\mem[6][12] ), .A2(n691), .ZN(n678) );
  OAI21_X1 U176 ( .B1(n476), .B2(n459), .A(n677), .ZN(n516) );
  NAND2_X1 U177 ( .A1(\mem[6][13] ), .A2(n691), .ZN(n677) );
  OAI21_X1 U178 ( .B1(n475), .B2(n459), .A(n676), .ZN(n515) );
  NAND2_X1 U179 ( .A1(\mem[6][14] ), .A2(n691), .ZN(n676) );
  OAI21_X1 U180 ( .B1(n474), .B2(n691), .A(n675), .ZN(n514) );
  NAND2_X1 U181 ( .A1(\mem[6][15] ), .A2(n691), .ZN(n675) );
  OAI21_X1 U182 ( .B1(n473), .B2(n691), .A(n674), .ZN(n513) );
  NAND2_X1 U183 ( .A1(\mem[6][16] ), .A2(n691), .ZN(n674) );
  OAI21_X1 U184 ( .B1(n472), .B2(n691), .A(n673), .ZN(n512) );
  NAND2_X1 U185 ( .A1(\mem[6][17] ), .A2(n691), .ZN(n673) );
  OAI21_X1 U186 ( .B1(n471), .B2(n691), .A(n672), .ZN(n511) );
  NAND2_X1 U187 ( .A1(\mem[6][18] ), .A2(n691), .ZN(n672) );
  OAI21_X1 U188 ( .B1(n470), .B2(n691), .A(n671), .ZN(n510) );
  NAND2_X1 U189 ( .A1(\mem[6][19] ), .A2(n459), .ZN(n671) );
  OAI21_X1 U190 ( .B1(n489), .B2(n670), .A(n669), .ZN(n509) );
  NAND2_X1 U191 ( .A1(\mem[7][0] ), .A2(n670), .ZN(n669) );
  OAI21_X1 U192 ( .B1(n488), .B2(n458), .A(n668), .ZN(n508) );
  NAND2_X1 U193 ( .A1(\mem[7][1] ), .A2(n670), .ZN(n668) );
  OAI21_X1 U194 ( .B1(n487), .B2(n458), .A(n667), .ZN(n507) );
  NAND2_X1 U195 ( .A1(\mem[7][2] ), .A2(n670), .ZN(n667) );
  OAI21_X1 U196 ( .B1(n486), .B2(n458), .A(n666), .ZN(n506) );
  NAND2_X1 U197 ( .A1(\mem[7][3] ), .A2(n670), .ZN(n666) );
  OAI21_X1 U198 ( .B1(n485), .B2(n458), .A(n665), .ZN(n505) );
  NAND2_X1 U199 ( .A1(\mem[7][4] ), .A2(n670), .ZN(n665) );
  OAI21_X1 U200 ( .B1(n484), .B2(n458), .A(n664), .ZN(n504) );
  NAND2_X1 U201 ( .A1(\mem[7][5] ), .A2(n670), .ZN(n664) );
  OAI21_X1 U202 ( .B1(n483), .B2(n458), .A(n663), .ZN(n503) );
  NAND2_X1 U203 ( .A1(\mem[7][6] ), .A2(n670), .ZN(n663) );
  OAI21_X1 U204 ( .B1(n482), .B2(n458), .A(n662), .ZN(n502) );
  NAND2_X1 U205 ( .A1(\mem[7][7] ), .A2(n670), .ZN(n662) );
  OAI21_X1 U206 ( .B1(n481), .B2(n458), .A(n661), .ZN(n501) );
  NAND2_X1 U207 ( .A1(\mem[7][8] ), .A2(n670), .ZN(n661) );
  OAI21_X1 U208 ( .B1(n480), .B2(n670), .A(n660), .ZN(n500) );
  NAND2_X1 U209 ( .A1(\mem[7][9] ), .A2(n670), .ZN(n660) );
  OAI21_X1 U210 ( .B1(n479), .B2(n458), .A(n659), .ZN(n499) );
  NAND2_X1 U211 ( .A1(\mem[7][10] ), .A2(n670), .ZN(n659) );
  OAI21_X1 U212 ( .B1(n478), .B2(n458), .A(n658), .ZN(n498) );
  NAND2_X1 U213 ( .A1(\mem[7][11] ), .A2(n670), .ZN(n658) );
  OAI21_X1 U214 ( .B1(n477), .B2(n670), .A(n657), .ZN(n497) );
  NAND2_X1 U215 ( .A1(\mem[7][12] ), .A2(n670), .ZN(n657) );
  OAI21_X1 U216 ( .B1(n476), .B2(n458), .A(n656), .ZN(n496) );
  NAND2_X1 U217 ( .A1(\mem[7][13] ), .A2(n670), .ZN(n656) );
  OAI21_X1 U218 ( .B1(n475), .B2(n670), .A(n655), .ZN(n495) );
  NAND2_X1 U219 ( .A1(\mem[7][14] ), .A2(n670), .ZN(n655) );
  OAI21_X1 U220 ( .B1(n474), .B2(n458), .A(n654), .ZN(n494) );
  NAND2_X1 U221 ( .A1(\mem[7][15] ), .A2(n670), .ZN(n654) );
  OAI21_X1 U222 ( .B1(n473), .B2(n458), .A(n653), .ZN(n493) );
  NAND2_X1 U223 ( .A1(\mem[7][16] ), .A2(n670), .ZN(n653) );
  OAI21_X1 U224 ( .B1(n472), .B2(n458), .A(n652), .ZN(n492) );
  NAND2_X1 U225 ( .A1(\mem[7][17] ), .A2(n670), .ZN(n652) );
  OAI21_X1 U226 ( .B1(n471), .B2(n458), .A(n651), .ZN(n491) );
  NAND2_X1 U227 ( .A1(\mem[7][18] ), .A2(n670), .ZN(n651) );
  OAI21_X1 U228 ( .B1(n470), .B2(n458), .A(n650), .ZN(n490) );
  NAND2_X1 U229 ( .A1(\mem[7][19] ), .A2(n670), .ZN(n650) );
  NAND2_X1 U230 ( .A1(wr_en), .A2(n469), .ZN(n735) );
  INV_X1 U231 ( .A(addr[3]), .ZN(n469) );
  OAI21_X1 U232 ( .B1(n465), .B2(n489), .A(n819), .ZN(n649) );
  NAND2_X1 U233 ( .A1(\mem[0][0] ), .A2(n465), .ZN(n819) );
  OAI21_X1 U234 ( .B1(n820), .B2(n488), .A(n818), .ZN(n648) );
  NAND2_X1 U235 ( .A1(\mem[0][1] ), .A2(n465), .ZN(n818) );
  OAI21_X1 U236 ( .B1(n820), .B2(n487), .A(n817), .ZN(n647) );
  NAND2_X1 U237 ( .A1(\mem[0][2] ), .A2(n465), .ZN(n817) );
  OAI21_X1 U238 ( .B1(n820), .B2(n486), .A(n816), .ZN(n646) );
  NAND2_X1 U239 ( .A1(\mem[0][3] ), .A2(n465), .ZN(n816) );
  OAI21_X1 U240 ( .B1(n820), .B2(n485), .A(n815), .ZN(n645) );
  NAND2_X1 U241 ( .A1(\mem[0][4] ), .A2(n465), .ZN(n815) );
  OAI21_X1 U242 ( .B1(n820), .B2(n484), .A(n814), .ZN(n644) );
  NAND2_X1 U243 ( .A1(\mem[0][5] ), .A2(n465), .ZN(n814) );
  OAI21_X1 U244 ( .B1(n820), .B2(n483), .A(n813), .ZN(n643) );
  NAND2_X1 U245 ( .A1(\mem[0][6] ), .A2(n465), .ZN(n813) );
  OAI21_X1 U246 ( .B1(n820), .B2(n482), .A(n812), .ZN(n642) );
  NAND2_X1 U247 ( .A1(\mem[0][7] ), .A2(n465), .ZN(n812) );
  OAI21_X1 U248 ( .B1(n820), .B2(n481), .A(n811), .ZN(n641) );
  NAND2_X1 U249 ( .A1(\mem[0][8] ), .A2(n465), .ZN(n811) );
  OAI21_X1 U250 ( .B1(n820), .B2(n480), .A(n810), .ZN(n640) );
  NAND2_X1 U251 ( .A1(\mem[0][9] ), .A2(n465), .ZN(n810) );
  OAI21_X1 U252 ( .B1(n820), .B2(n479), .A(n809), .ZN(n639) );
  NAND2_X1 U253 ( .A1(\mem[0][10] ), .A2(n465), .ZN(n809) );
  OAI21_X1 U254 ( .B1(n820), .B2(n478), .A(n808), .ZN(n638) );
  NAND2_X1 U255 ( .A1(\mem[0][11] ), .A2(n465), .ZN(n808) );
  OAI21_X1 U256 ( .B1(n489), .B2(n798), .A(n797), .ZN(n629) );
  NAND2_X1 U257 ( .A1(\mem[1][0] ), .A2(n464), .ZN(n797) );
  OAI21_X1 U258 ( .B1(n488), .B2(n798), .A(n796), .ZN(n628) );
  NAND2_X1 U259 ( .A1(\mem[1][1] ), .A2(n464), .ZN(n796) );
  OAI21_X1 U260 ( .B1(n487), .B2(n798), .A(n795), .ZN(n627) );
  NAND2_X1 U261 ( .A1(\mem[1][2] ), .A2(n464), .ZN(n795) );
  OAI21_X1 U262 ( .B1(n486), .B2(n798), .A(n794), .ZN(n626) );
  NAND2_X1 U263 ( .A1(\mem[1][3] ), .A2(n464), .ZN(n794) );
  OAI21_X1 U264 ( .B1(n485), .B2(n798), .A(n793), .ZN(n625) );
  NAND2_X1 U265 ( .A1(\mem[1][4] ), .A2(n464), .ZN(n793) );
  OAI21_X1 U266 ( .B1(n484), .B2(n798), .A(n792), .ZN(n624) );
  NAND2_X1 U267 ( .A1(\mem[1][5] ), .A2(n464), .ZN(n792) );
  OAI21_X1 U268 ( .B1(n483), .B2(n798), .A(n791), .ZN(n623) );
  NAND2_X1 U269 ( .A1(\mem[1][6] ), .A2(n464), .ZN(n791) );
  OAI21_X1 U270 ( .B1(n482), .B2(n798), .A(n790), .ZN(n622) );
  NAND2_X1 U271 ( .A1(\mem[1][7] ), .A2(n464), .ZN(n790) );
  OAI21_X1 U272 ( .B1(n481), .B2(n798), .A(n789), .ZN(n621) );
  NAND2_X1 U273 ( .A1(\mem[1][8] ), .A2(n464), .ZN(n789) );
  OAI21_X1 U274 ( .B1(n480), .B2(n464), .A(n788), .ZN(n620) );
  NAND2_X1 U275 ( .A1(\mem[1][9] ), .A2(n464), .ZN(n788) );
  OAI21_X1 U276 ( .B1(n479), .B2(n798), .A(n787), .ZN(n619) );
  NAND2_X1 U277 ( .A1(\mem[1][10] ), .A2(n464), .ZN(n787) );
  OAI21_X1 U278 ( .B1(n478), .B2(n798), .A(n786), .ZN(n618) );
  NAND2_X1 U279 ( .A1(\mem[1][11] ), .A2(n464), .ZN(n786) );
  OAI21_X1 U280 ( .B1(n489), .B2(n777), .A(n776), .ZN(n609) );
  NAND2_X1 U281 ( .A1(\mem[2][0] ), .A2(n777), .ZN(n776) );
  OAI21_X1 U282 ( .B1(n488), .B2(n777), .A(n775), .ZN(n608) );
  NAND2_X1 U283 ( .A1(\mem[2][1] ), .A2(n777), .ZN(n775) );
  OAI21_X1 U284 ( .B1(n487), .B2(n777), .A(n774), .ZN(n607) );
  NAND2_X1 U285 ( .A1(\mem[2][2] ), .A2(n777), .ZN(n774) );
  OAI21_X1 U286 ( .B1(n486), .B2(n777), .A(n773), .ZN(n606) );
  NAND2_X1 U287 ( .A1(\mem[2][3] ), .A2(n463), .ZN(n773) );
  OAI21_X1 U288 ( .B1(n485), .B2(n777), .A(n772), .ZN(n605) );
  NAND2_X1 U289 ( .A1(\mem[2][4] ), .A2(n463), .ZN(n772) );
  OAI21_X1 U290 ( .B1(n484), .B2(n777), .A(n771), .ZN(n604) );
  NAND2_X1 U291 ( .A1(\mem[2][5] ), .A2(n463), .ZN(n771) );
  OAI21_X1 U292 ( .B1(n483), .B2(n777), .A(n770), .ZN(n603) );
  NAND2_X1 U293 ( .A1(\mem[2][6] ), .A2(n777), .ZN(n770) );
  OAI21_X1 U294 ( .B1(n482), .B2(n777), .A(n769), .ZN(n602) );
  NAND2_X1 U295 ( .A1(\mem[2][7] ), .A2(n777), .ZN(n769) );
  OAI21_X1 U296 ( .B1(n481), .B2(n777), .A(n768), .ZN(n601) );
  NAND2_X1 U297 ( .A1(\mem[2][8] ), .A2(n777), .ZN(n768) );
  OAI21_X1 U298 ( .B1(n480), .B2(n463), .A(n767), .ZN(n600) );
  NAND2_X1 U299 ( .A1(\mem[2][9] ), .A2(n463), .ZN(n767) );
  OAI21_X1 U300 ( .B1(n479), .B2(n777), .A(n766), .ZN(n599) );
  NAND2_X1 U301 ( .A1(\mem[2][10] ), .A2(n777), .ZN(n766) );
  OAI21_X1 U302 ( .B1(n478), .B2(n777), .A(n765), .ZN(n598) );
  NAND2_X1 U303 ( .A1(\mem[2][11] ), .A2(n777), .ZN(n765) );
  OAI21_X1 U304 ( .B1(n489), .B2(n756), .A(n755), .ZN(n589) );
  NAND2_X1 U305 ( .A1(\mem[3][0] ), .A2(n462), .ZN(n755) );
  OAI21_X1 U306 ( .B1(n488), .B2(n756), .A(n754), .ZN(n588) );
  NAND2_X1 U307 ( .A1(\mem[3][1] ), .A2(n462), .ZN(n754) );
  OAI21_X1 U308 ( .B1(n487), .B2(n756), .A(n753), .ZN(n587) );
  NAND2_X1 U309 ( .A1(\mem[3][2] ), .A2(n462), .ZN(n753) );
  OAI21_X1 U310 ( .B1(n486), .B2(n756), .A(n752), .ZN(n586) );
  NAND2_X1 U311 ( .A1(\mem[3][3] ), .A2(n462), .ZN(n752) );
  OAI21_X1 U312 ( .B1(n485), .B2(n756), .A(n751), .ZN(n585) );
  NAND2_X1 U313 ( .A1(\mem[3][4] ), .A2(n462), .ZN(n751) );
  OAI21_X1 U314 ( .B1(n484), .B2(n756), .A(n750), .ZN(n584) );
  NAND2_X1 U315 ( .A1(\mem[3][5] ), .A2(n462), .ZN(n750) );
  OAI21_X1 U316 ( .B1(n483), .B2(n756), .A(n749), .ZN(n583) );
  NAND2_X1 U317 ( .A1(\mem[3][6] ), .A2(n462), .ZN(n749) );
  OAI21_X1 U318 ( .B1(n482), .B2(n756), .A(n748), .ZN(n582) );
  NAND2_X1 U319 ( .A1(\mem[3][7] ), .A2(n462), .ZN(n748) );
  OAI21_X1 U320 ( .B1(n481), .B2(n756), .A(n747), .ZN(n581) );
  NAND2_X1 U321 ( .A1(\mem[3][8] ), .A2(n462), .ZN(n747) );
  OAI21_X1 U322 ( .B1(n480), .B2(n462), .A(n746), .ZN(n580) );
  NAND2_X1 U323 ( .A1(\mem[3][9] ), .A2(n462), .ZN(n746) );
  OAI21_X1 U324 ( .B1(n479), .B2(n756), .A(n745), .ZN(n579) );
  NAND2_X1 U325 ( .A1(\mem[3][10] ), .A2(n462), .ZN(n745) );
  OAI21_X1 U326 ( .B1(n478), .B2(n756), .A(n744), .ZN(n578) );
  NAND2_X1 U327 ( .A1(\mem[3][11] ), .A2(n462), .ZN(n744) );
  OAI21_X1 U328 ( .B1(n820), .B2(n477), .A(n807), .ZN(n637) );
  NAND2_X1 U329 ( .A1(\mem[0][12] ), .A2(n820), .ZN(n807) );
  OAI21_X1 U330 ( .B1(n820), .B2(n476), .A(n806), .ZN(n636) );
  NAND2_X1 U331 ( .A1(\mem[0][13] ), .A2(n820), .ZN(n806) );
  OAI21_X1 U332 ( .B1(n465), .B2(n475), .A(n805), .ZN(n635) );
  NAND2_X1 U333 ( .A1(\mem[0][14] ), .A2(n820), .ZN(n805) );
  OAI21_X1 U334 ( .B1(n820), .B2(n474), .A(n804), .ZN(n634) );
  NAND2_X1 U335 ( .A1(\mem[0][15] ), .A2(n465), .ZN(n804) );
  OAI21_X1 U336 ( .B1(n820), .B2(n473), .A(n803), .ZN(n633) );
  NAND2_X1 U337 ( .A1(\mem[0][16] ), .A2(n820), .ZN(n803) );
  OAI21_X1 U338 ( .B1(n820), .B2(n472), .A(n802), .ZN(n632) );
  NAND2_X1 U339 ( .A1(\mem[0][17] ), .A2(n820), .ZN(n802) );
  OAI21_X1 U340 ( .B1(n820), .B2(n471), .A(n801), .ZN(n631) );
  NAND2_X1 U341 ( .A1(\mem[0][18] ), .A2(n820), .ZN(n801) );
  OAI21_X1 U342 ( .B1(n820), .B2(n470), .A(n800), .ZN(n630) );
  NAND2_X1 U343 ( .A1(\mem[0][19] ), .A2(n465), .ZN(n800) );
  INV_X1 U344 ( .A(data_in[0]), .ZN(n489) );
  INV_X1 U345 ( .A(data_in[1]), .ZN(n488) );
  INV_X1 U346 ( .A(data_in[2]), .ZN(n487) );
  INV_X1 U347 ( .A(data_in[3]), .ZN(n486) );
  INV_X1 U348 ( .A(data_in[4]), .ZN(n485) );
  INV_X1 U349 ( .A(data_in[5]), .ZN(n484) );
  INV_X1 U358 ( .A(data_in[6]), .ZN(n483) );
  INV_X1 U359 ( .A(data_in[7]), .ZN(n482) );
  INV_X1 U360 ( .A(data_in[8]), .ZN(n481) );
  INV_X1 U361 ( .A(data_in[9]), .ZN(n480) );
  INV_X1 U362 ( .A(data_in[10]), .ZN(n479) );
  INV_X1 U363 ( .A(data_in[11]), .ZN(n478) );
  INV_X1 U364 ( .A(data_in[12]), .ZN(n477) );
  INV_X1 U365 ( .A(data_in[13]), .ZN(n476) );
  INV_X1 U366 ( .A(data_in[14]), .ZN(n475) );
  INV_X1 U367 ( .A(data_in[15]), .ZN(n474) );
  INV_X1 U368 ( .A(data_in[16]), .ZN(n473) );
  INV_X1 U369 ( .A(data_in[17]), .ZN(n472) );
  INV_X1 U370 ( .A(data_in[18]), .ZN(n471) );
  INV_X1 U371 ( .A(data_in[19]), .ZN(n470) );
  MUX2_X1 U372 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n455), .Z(n1) );
  MUX2_X1 U373 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n454), .Z(n2) );
  MUX2_X1 U374 ( .A(n2), .B(n1), .S(n453), .Z(n3) );
  MUX2_X1 U375 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n456), .Z(n4) );
  MUX2_X1 U376 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n457), .Z(n5) );
  MUX2_X1 U377 ( .A(n5), .B(n4), .S(n453), .Z(n6) );
  MUX2_X1 U378 ( .A(n6), .B(n3), .S(N12), .Z(N32) );
  MUX2_X1 U379 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n455), .Z(n7) );
  MUX2_X1 U380 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n456), .Z(n8) );
  MUX2_X1 U381 ( .A(n8), .B(n7), .S(n453), .Z(n9) );
  MUX2_X1 U382 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n457), .Z(n10) );
  MUX2_X1 U383 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n454), .Z(n11) );
  MUX2_X1 U384 ( .A(n11), .B(n10), .S(n453), .Z(n12) );
  MUX2_X1 U385 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n454), .Z(n13) );
  MUX2_X1 U386 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n454), .Z(n14) );
  MUX2_X1 U387 ( .A(n14), .B(n13), .S(n453), .Z(n15) );
  MUX2_X1 U388 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n456), .Z(n16) );
  MUX2_X1 U389 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n454), .Z(n17) );
  MUX2_X1 U390 ( .A(n17), .B(n16), .S(n453), .Z(n18) );
  MUX2_X1 U391 ( .A(n18), .B(n15), .S(N12), .Z(N30) );
  MUX2_X1 U392 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n457), .Z(n19) );
  MUX2_X1 U393 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n455), .Z(n20) );
  MUX2_X1 U394 ( .A(n20), .B(n19), .S(n453), .Z(n21) );
  MUX2_X1 U395 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n456), .Z(n22) );
  MUX2_X1 U396 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n457), .Z(n23) );
  MUX2_X1 U397 ( .A(n23), .B(n22), .S(n453), .Z(n24) );
  MUX2_X1 U398 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n457), .Z(n356) );
  MUX2_X1 U399 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n457), .Z(n357) );
  MUX2_X1 U400 ( .A(n357), .B(n356), .S(n453), .Z(n358) );
  MUX2_X1 U401 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n456), .Z(n359) );
  MUX2_X1 U402 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n455), .Z(n360) );
  MUX2_X1 U403 ( .A(n360), .B(n359), .S(n453), .Z(n361) );
  MUX2_X1 U404 ( .A(n361), .B(n358), .S(N12), .Z(N28) );
  MUX2_X1 U405 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n454), .Z(n362) );
  MUX2_X1 U406 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n454), .Z(n363) );
  MUX2_X1 U407 ( .A(n363), .B(n362), .S(n453), .Z(n364) );
  MUX2_X1 U408 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n454), .Z(n365) );
  MUX2_X1 U409 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n454), .Z(n366) );
  MUX2_X1 U410 ( .A(n366), .B(n365), .S(n453), .Z(n367) );
  MUX2_X1 U411 ( .A(n367), .B(n364), .S(N12), .Z(N27) );
  MUX2_X1 U412 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n454), .Z(n368) );
  MUX2_X1 U413 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n454), .Z(n369) );
  MUX2_X1 U414 ( .A(n369), .B(n368), .S(n453), .Z(n370) );
  MUX2_X1 U415 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n454), .Z(n371) );
  MUX2_X1 U416 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n454), .Z(n372) );
  MUX2_X1 U417 ( .A(n372), .B(n371), .S(n453), .Z(n373) );
  MUX2_X1 U418 ( .A(n373), .B(n370), .S(N12), .Z(N26) );
  MUX2_X1 U419 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n454), .Z(n374) );
  MUX2_X1 U420 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n454), .Z(n375) );
  MUX2_X1 U421 ( .A(n375), .B(n374), .S(n453), .Z(n376) );
  MUX2_X1 U422 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n454), .Z(n377) );
  MUX2_X1 U423 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n454), .Z(n378) );
  MUX2_X1 U424 ( .A(n378), .B(n377), .S(n453), .Z(n379) );
  MUX2_X1 U425 ( .A(n379), .B(n376), .S(N12), .Z(N25) );
  MUX2_X1 U426 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n455), .Z(n380) );
  MUX2_X1 U427 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n455), .Z(n381) );
  MUX2_X1 U428 ( .A(n381), .B(n380), .S(n452), .Z(n382) );
  MUX2_X1 U429 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n455), .Z(n383) );
  MUX2_X1 U430 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n455), .Z(n384) );
  MUX2_X1 U431 ( .A(n384), .B(n383), .S(n452), .Z(n385) );
  MUX2_X1 U432 ( .A(n385), .B(n382), .S(N12), .Z(N24) );
  MUX2_X1 U433 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n455), .Z(n386) );
  MUX2_X1 U434 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n455), .Z(n387) );
  MUX2_X1 U435 ( .A(n387), .B(n386), .S(n452), .Z(n388) );
  MUX2_X1 U436 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n455), .Z(n389) );
  MUX2_X1 U437 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n455), .Z(n390) );
  MUX2_X1 U438 ( .A(n390), .B(n389), .S(n452), .Z(n391) );
  MUX2_X1 U439 ( .A(n391), .B(n388), .S(N12), .Z(N23) );
  MUX2_X1 U440 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n455), .Z(n392) );
  MUX2_X1 U441 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n455), .Z(n393) );
  MUX2_X1 U442 ( .A(n393), .B(n392), .S(n452), .Z(n394) );
  MUX2_X1 U443 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n455), .Z(n395) );
  MUX2_X1 U444 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n455), .Z(n396) );
  MUX2_X1 U445 ( .A(n396), .B(n395), .S(n452), .Z(n397) );
  MUX2_X1 U446 ( .A(n397), .B(n394), .S(N12), .Z(N22) );
  MUX2_X1 U447 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n456), .Z(n398) );
  MUX2_X1 U448 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n456), .Z(n399) );
  MUX2_X1 U449 ( .A(n399), .B(n398), .S(n452), .Z(n400) );
  MUX2_X1 U450 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n456), .Z(n401) );
  MUX2_X1 U451 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n456), .Z(n402) );
  MUX2_X1 U452 ( .A(n402), .B(n401), .S(n452), .Z(n403) );
  MUX2_X1 U453 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n456), .Z(n404) );
  MUX2_X1 U454 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n456), .Z(n405) );
  MUX2_X1 U455 ( .A(n405), .B(n404), .S(n452), .Z(n406) );
  MUX2_X1 U456 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n456), .Z(n407) );
  MUX2_X1 U457 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n456), .Z(n408) );
  MUX2_X1 U458 ( .A(n408), .B(n407), .S(n452), .Z(n409) );
  MUX2_X1 U459 ( .A(n409), .B(n406), .S(N12), .Z(N20) );
  MUX2_X1 U460 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n456), .Z(n410) );
  MUX2_X1 U461 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n456), .Z(n411) );
  MUX2_X1 U462 ( .A(n411), .B(n410), .S(n452), .Z(n412) );
  MUX2_X1 U463 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n456), .Z(n413) );
  MUX2_X1 U464 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n456), .Z(n414) );
  MUX2_X1 U465 ( .A(n414), .B(n413), .S(n452), .Z(n415) );
  MUX2_X1 U466 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n457), .Z(n416) );
  MUX2_X1 U467 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n457), .Z(n417) );
  MUX2_X1 U468 ( .A(n417), .B(n416), .S(n453), .Z(n418) );
  MUX2_X1 U469 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n457), .Z(n419) );
  MUX2_X1 U470 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n457), .Z(n420) );
  MUX2_X1 U471 ( .A(n420), .B(n419), .S(n453), .Z(n421) );
  MUX2_X1 U472 ( .A(n421), .B(n418), .S(N12), .Z(N18) );
  MUX2_X1 U473 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n457), .Z(n422) );
  MUX2_X1 U474 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n457), .Z(n423) );
  MUX2_X1 U475 ( .A(n423), .B(n422), .S(n453), .Z(n424) );
  MUX2_X1 U476 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n457), .Z(n425) );
  MUX2_X1 U477 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n457), .Z(n426) );
  MUX2_X1 U478 ( .A(n426), .B(n425), .S(N11), .Z(n427) );
  MUX2_X1 U479 ( .A(n427), .B(n424), .S(N12), .Z(N17) );
  MUX2_X1 U480 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n457), .Z(n428) );
  MUX2_X1 U481 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n457), .Z(n429) );
  MUX2_X1 U482 ( .A(n429), .B(n428), .S(n453), .Z(n430) );
  MUX2_X1 U483 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n457), .Z(n431) );
  MUX2_X1 U484 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n457), .Z(n432) );
  MUX2_X1 U485 ( .A(n432), .B(n431), .S(N11), .Z(n433) );
  MUX2_X1 U486 ( .A(n433), .B(n430), .S(N12), .Z(N16) );
  MUX2_X1 U487 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n454), .Z(n434) );
  MUX2_X1 U488 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n455), .Z(n435) );
  MUX2_X1 U489 ( .A(n435), .B(n434), .S(N11), .Z(n436) );
  MUX2_X1 U490 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n455), .Z(n437) );
  MUX2_X1 U491 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n456), .Z(n438) );
  MUX2_X1 U492 ( .A(n438), .B(n437), .S(N11), .Z(n439) );
  MUX2_X1 U493 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n454), .Z(n440) );
  MUX2_X1 U494 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n455), .Z(n441) );
  MUX2_X1 U495 ( .A(n441), .B(n440), .S(n453), .Z(n442) );
  MUX2_X1 U496 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n457), .Z(n443) );
  MUX2_X1 U497 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n456), .Z(n444) );
  MUX2_X1 U498 ( .A(n444), .B(n443), .S(N11), .Z(n445) );
  MUX2_X1 U499 ( .A(n445), .B(n442), .S(N12), .Z(N14) );
  MUX2_X1 U500 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n457), .Z(n446) );
  MUX2_X1 U501 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n456), .Z(n447) );
  MUX2_X1 U502 ( .A(n447), .B(n446), .S(n453), .Z(n448) );
  MUX2_X1 U503 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n455), .Z(n449) );
  MUX2_X1 U504 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n454), .Z(n450) );
  MUX2_X1 U505 ( .A(n450), .B(n449), .S(N11), .Z(n451) );
  MUX2_X1 U506 ( .A(n451), .B(n448), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE4_2 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N13, N14, N16, N18, N20, N21, N22, N23, N24, N26, N27,
         N28, N29, N30, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[19]  ( .D(N13), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N20), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N21), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N23), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N27), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N29), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N30), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N32), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n490), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n491), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n492), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n493), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n494), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n495), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n496), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n497), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n498), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n499), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n500), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n501), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n502), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n503), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n504), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n505), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n506), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n507), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n508), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n509), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n510), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n511), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n512), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n513), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n514), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n515), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n516), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n517), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n518), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n519), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n520), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n521), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n522), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n523), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n524), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n525), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n526), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n527), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n528), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n529), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n530), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n531), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n532), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n533), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n534), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n535), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n536), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n537), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n538), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n539), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n540), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n541), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n542), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n543), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n544), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n545), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n546), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n547), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n548), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n549), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n550), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n551), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n552), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n553), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n554), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n555), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n556), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n557), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n558), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n559), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n560), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n561), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n562), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n563), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n564), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n565), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n566), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n567), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n568), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n569), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n570), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n571), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n572), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n573), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n574), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n575), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n576), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n577), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n578), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n579), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n580), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n581), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n582), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n583), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n584), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n585), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n586), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n587), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n588), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n589), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n590), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n591), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n592), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n593), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n594), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n595), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n596), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n597), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n598), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n599), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n600), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n601), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n602), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n603), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n604), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n605), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n606), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n607), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n608), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n609), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n610), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n611), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n612), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n613), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n614), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n615), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n616), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n617), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n618), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n619), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n620), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n621), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n622), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n623), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n624), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n625), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n626), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n627), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n628), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n629), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n630), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n631), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n632), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n633), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n634), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n635), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n636), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n637), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n638), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n639), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n640), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n641), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n642), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n643), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n644), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n645), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n646), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n647), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n648), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n649), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U350 ( .A1(n466), .A2(n467), .A3(n799), .ZN(n820) );
  NAND3_X1 U351 ( .A1(n799), .A2(n467), .A3(N10), .ZN(n798) );
  NAND3_X1 U352 ( .A1(n799), .A2(n466), .A3(N11), .ZN(n777) );
  NAND3_X1 U353 ( .A1(N10), .A2(n799), .A3(N11), .ZN(n756) );
  NAND3_X1 U354 ( .A1(n466), .A2(n467), .A3(n713), .ZN(n734) );
  NAND3_X1 U355 ( .A1(N10), .A2(n467), .A3(n713), .ZN(n712) );
  NAND3_X1 U356 ( .A1(N11), .A2(n466), .A3(n713), .ZN(n691) );
  NAND3_X1 U357 ( .A1(N11), .A2(N10), .A3(n713), .ZN(n670) );
  SDFF_X1 \data_out_reg[15]  ( .D(n424), .SI(n427), .SE(n468), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n412), .SI(n415), .SE(n468), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[17]  ( .D(n436), .SI(n439), .SE(n468), .CK(clk), .Q(
        data_out[17]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n376), .SI(n379), .SE(n468), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n9), .SI(n12), .SE(n468), .CK(clk), .Q(
        data_out[1]) );
  BUF_X1 U3 ( .A(n820), .Z(n465) );
  BUF_X1 U4 ( .A(n777), .Z(n463) );
  BUF_X1 U5 ( .A(n712), .Z(n460) );
  BUF_X1 U6 ( .A(n453), .Z(n452) );
  BUF_X1 U7 ( .A(N10), .Z(n454) );
  BUF_X1 U8 ( .A(N10), .Z(n455) );
  BUF_X1 U9 ( .A(N10), .Z(n456) );
  BUF_X1 U10 ( .A(N10), .Z(n457) );
  BUF_X1 U11 ( .A(N11), .Z(n453) );
  BUF_X1 U12 ( .A(n756), .Z(n462) );
  BUF_X1 U13 ( .A(n798), .Z(n464) );
  BUF_X1 U14 ( .A(n670), .Z(n458) );
  BUF_X1 U15 ( .A(n734), .Z(n461) );
  BUF_X1 U16 ( .A(n691), .Z(n459) );
  NOR2_X1 U17 ( .A1(n735), .A2(N12), .ZN(n799) );
  NOR2_X1 U18 ( .A1(n468), .A2(n735), .ZN(n713) );
  INV_X1 U19 ( .A(N12), .ZN(n468) );
  INV_X1 U20 ( .A(N11), .ZN(n467) );
  INV_X1 U21 ( .A(N10), .ZN(n466) );
  OAI21_X1 U22 ( .B1(n477), .B2(n798), .A(n785), .ZN(n617) );
  NAND2_X1 U23 ( .A1(\mem[1][12] ), .A2(n798), .ZN(n785) );
  OAI21_X1 U24 ( .B1(n476), .B2(n798), .A(n784), .ZN(n616) );
  NAND2_X1 U25 ( .A1(\mem[1][13] ), .A2(n798), .ZN(n784) );
  OAI21_X1 U26 ( .B1(n475), .B2(n798), .A(n783), .ZN(n615) );
  NAND2_X1 U27 ( .A1(\mem[1][14] ), .A2(n798), .ZN(n783) );
  OAI21_X1 U28 ( .B1(n474), .B2(n464), .A(n782), .ZN(n614) );
  NAND2_X1 U29 ( .A1(\mem[1][15] ), .A2(n798), .ZN(n782) );
  OAI21_X1 U30 ( .B1(n473), .B2(n798), .A(n781), .ZN(n613) );
  NAND2_X1 U31 ( .A1(\mem[1][16] ), .A2(n464), .ZN(n781) );
  OAI21_X1 U32 ( .B1(n472), .B2(n798), .A(n780), .ZN(n612) );
  NAND2_X1 U33 ( .A1(\mem[1][17] ), .A2(n798), .ZN(n780) );
  OAI21_X1 U34 ( .B1(n471), .B2(n798), .A(n779), .ZN(n611) );
  NAND2_X1 U35 ( .A1(\mem[1][18] ), .A2(n798), .ZN(n779) );
  OAI21_X1 U36 ( .B1(n470), .B2(n798), .A(n778), .ZN(n610) );
  NAND2_X1 U37 ( .A1(\mem[1][19] ), .A2(n464), .ZN(n778) );
  OAI21_X1 U38 ( .B1(n477), .B2(n777), .A(n764), .ZN(n597) );
  NAND2_X1 U39 ( .A1(\mem[2][12] ), .A2(n777), .ZN(n764) );
  OAI21_X1 U40 ( .B1(n476), .B2(n777), .A(n763), .ZN(n596) );
  NAND2_X1 U41 ( .A1(\mem[2][13] ), .A2(n777), .ZN(n763) );
  OAI21_X1 U42 ( .B1(n475), .B2(n463), .A(n762), .ZN(n595) );
  NAND2_X1 U43 ( .A1(\mem[2][14] ), .A2(n777), .ZN(n762) );
  OAI21_X1 U44 ( .B1(n474), .B2(n463), .A(n761), .ZN(n594) );
  NAND2_X1 U45 ( .A1(\mem[2][15] ), .A2(n777), .ZN(n761) );
  OAI21_X1 U46 ( .B1(n473), .B2(n463), .A(n760), .ZN(n593) );
  NAND2_X1 U47 ( .A1(\mem[2][16] ), .A2(n777), .ZN(n760) );
  OAI21_X1 U48 ( .B1(n472), .B2(n463), .A(n759), .ZN(n592) );
  NAND2_X1 U49 ( .A1(\mem[2][17] ), .A2(n777), .ZN(n759) );
  OAI21_X1 U50 ( .B1(n471), .B2(n463), .A(n758), .ZN(n591) );
  NAND2_X1 U51 ( .A1(\mem[2][18] ), .A2(n777), .ZN(n758) );
  OAI21_X1 U52 ( .B1(n470), .B2(n777), .A(n757), .ZN(n590) );
  NAND2_X1 U53 ( .A1(\mem[2][19] ), .A2(n777), .ZN(n757) );
  OAI21_X1 U54 ( .B1(n477), .B2(n756), .A(n743), .ZN(n577) );
  NAND2_X1 U55 ( .A1(\mem[3][12] ), .A2(n756), .ZN(n743) );
  OAI21_X1 U56 ( .B1(n476), .B2(n756), .A(n742), .ZN(n576) );
  NAND2_X1 U57 ( .A1(\mem[3][13] ), .A2(n756), .ZN(n742) );
  OAI21_X1 U58 ( .B1(n475), .B2(n756), .A(n741), .ZN(n575) );
  NAND2_X1 U59 ( .A1(\mem[3][14] ), .A2(n756), .ZN(n741) );
  OAI21_X1 U60 ( .B1(n474), .B2(n462), .A(n740), .ZN(n574) );
  NAND2_X1 U61 ( .A1(\mem[3][15] ), .A2(n756), .ZN(n740) );
  OAI21_X1 U62 ( .B1(n473), .B2(n756), .A(n739), .ZN(n573) );
  NAND2_X1 U63 ( .A1(\mem[3][16] ), .A2(n462), .ZN(n739) );
  OAI21_X1 U64 ( .B1(n472), .B2(n756), .A(n738), .ZN(n572) );
  NAND2_X1 U65 ( .A1(\mem[3][17] ), .A2(n756), .ZN(n738) );
  OAI21_X1 U66 ( .B1(n471), .B2(n756), .A(n737), .ZN(n571) );
  NAND2_X1 U67 ( .A1(\mem[3][18] ), .A2(n756), .ZN(n737) );
  OAI21_X1 U68 ( .B1(n470), .B2(n756), .A(n736), .ZN(n570) );
  NAND2_X1 U69 ( .A1(\mem[3][19] ), .A2(n462), .ZN(n736) );
  OAI21_X1 U70 ( .B1(n489), .B2(n734), .A(n733), .ZN(n569) );
  NAND2_X1 U71 ( .A1(\mem[4][0] ), .A2(n461), .ZN(n733) );
  OAI21_X1 U72 ( .B1(n488), .B2(n734), .A(n732), .ZN(n568) );
  NAND2_X1 U73 ( .A1(\mem[4][1] ), .A2(n461), .ZN(n732) );
  OAI21_X1 U74 ( .B1(n487), .B2(n734), .A(n731), .ZN(n567) );
  NAND2_X1 U75 ( .A1(\mem[4][2] ), .A2(n461), .ZN(n731) );
  OAI21_X1 U76 ( .B1(n486), .B2(n734), .A(n730), .ZN(n566) );
  NAND2_X1 U77 ( .A1(\mem[4][3] ), .A2(n461), .ZN(n730) );
  OAI21_X1 U78 ( .B1(n485), .B2(n461), .A(n729), .ZN(n565) );
  NAND2_X1 U79 ( .A1(\mem[4][4] ), .A2(n461), .ZN(n729) );
  OAI21_X1 U80 ( .B1(n484), .B2(n734), .A(n728), .ZN(n564) );
  NAND2_X1 U81 ( .A1(\mem[4][5] ), .A2(n461), .ZN(n728) );
  OAI21_X1 U82 ( .B1(n483), .B2(n734), .A(n727), .ZN(n563) );
  NAND2_X1 U83 ( .A1(\mem[4][6] ), .A2(n461), .ZN(n727) );
  OAI21_X1 U84 ( .B1(n482), .B2(n734), .A(n726), .ZN(n562) );
  NAND2_X1 U85 ( .A1(\mem[4][7] ), .A2(n461), .ZN(n726) );
  OAI21_X1 U86 ( .B1(n481), .B2(n734), .A(n725), .ZN(n561) );
  NAND2_X1 U87 ( .A1(\mem[4][8] ), .A2(n461), .ZN(n725) );
  OAI21_X1 U88 ( .B1(n480), .B2(n734), .A(n724), .ZN(n560) );
  NAND2_X1 U89 ( .A1(\mem[4][9] ), .A2(n461), .ZN(n724) );
  OAI21_X1 U90 ( .B1(n479), .B2(n734), .A(n723), .ZN(n559) );
  NAND2_X1 U91 ( .A1(\mem[4][10] ), .A2(n461), .ZN(n723) );
  OAI21_X1 U92 ( .B1(n478), .B2(n734), .A(n722), .ZN(n558) );
  NAND2_X1 U93 ( .A1(\mem[4][11] ), .A2(n461), .ZN(n722) );
  OAI21_X1 U94 ( .B1(n477), .B2(n734), .A(n721), .ZN(n557) );
  NAND2_X1 U95 ( .A1(\mem[4][12] ), .A2(n734), .ZN(n721) );
  OAI21_X1 U96 ( .B1(n476), .B2(n461), .A(n720), .ZN(n556) );
  NAND2_X1 U97 ( .A1(\mem[4][13] ), .A2(n734), .ZN(n720) );
  OAI21_X1 U98 ( .B1(n475), .B2(n461), .A(n719), .ZN(n555) );
  NAND2_X1 U99 ( .A1(\mem[4][14] ), .A2(n734), .ZN(n719) );
  OAI21_X1 U100 ( .B1(n474), .B2(n734), .A(n718), .ZN(n554) );
  NAND2_X1 U101 ( .A1(\mem[4][15] ), .A2(n734), .ZN(n718) );
  OAI21_X1 U102 ( .B1(n473), .B2(n734), .A(n717), .ZN(n553) );
  NAND2_X1 U103 ( .A1(\mem[4][16] ), .A2(n734), .ZN(n717) );
  OAI21_X1 U104 ( .B1(n472), .B2(n734), .A(n716), .ZN(n552) );
  NAND2_X1 U105 ( .A1(\mem[4][17] ), .A2(n734), .ZN(n716) );
  OAI21_X1 U106 ( .B1(n471), .B2(n734), .A(n715), .ZN(n551) );
  NAND2_X1 U107 ( .A1(\mem[4][18] ), .A2(n734), .ZN(n715) );
  OAI21_X1 U108 ( .B1(n470), .B2(n734), .A(n714), .ZN(n550) );
  NAND2_X1 U109 ( .A1(\mem[4][19] ), .A2(n461), .ZN(n714) );
  OAI21_X1 U110 ( .B1(n489), .B2(n712), .A(n711), .ZN(n549) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n712), .ZN(n711) );
  OAI21_X1 U112 ( .B1(n488), .B2(n460), .A(n710), .ZN(n548) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n712), .ZN(n710) );
  OAI21_X1 U114 ( .B1(n487), .B2(n460), .A(n709), .ZN(n547) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n712), .ZN(n709) );
  OAI21_X1 U116 ( .B1(n486), .B2(n460), .A(n708), .ZN(n546) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n712), .ZN(n708) );
  OAI21_X1 U118 ( .B1(n485), .B2(n460), .A(n707), .ZN(n545) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n712), .ZN(n707) );
  OAI21_X1 U120 ( .B1(n484), .B2(n460), .A(n706), .ZN(n544) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n712), .ZN(n706) );
  OAI21_X1 U122 ( .B1(n483), .B2(n460), .A(n705), .ZN(n543) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n712), .ZN(n705) );
  OAI21_X1 U124 ( .B1(n482), .B2(n460), .A(n704), .ZN(n542) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n712), .ZN(n704) );
  OAI21_X1 U126 ( .B1(n481), .B2(n460), .A(n703), .ZN(n541) );
  NAND2_X1 U127 ( .A1(\mem[5][8] ), .A2(n712), .ZN(n703) );
  OAI21_X1 U128 ( .B1(n480), .B2(n712), .A(n702), .ZN(n540) );
  NAND2_X1 U129 ( .A1(\mem[5][9] ), .A2(n712), .ZN(n702) );
  OAI21_X1 U130 ( .B1(n479), .B2(n460), .A(n701), .ZN(n539) );
  NAND2_X1 U131 ( .A1(\mem[5][10] ), .A2(n712), .ZN(n701) );
  OAI21_X1 U132 ( .B1(n478), .B2(n460), .A(n700), .ZN(n538) );
  NAND2_X1 U133 ( .A1(\mem[5][11] ), .A2(n712), .ZN(n700) );
  OAI21_X1 U134 ( .B1(n477), .B2(n712), .A(n699), .ZN(n537) );
  NAND2_X1 U135 ( .A1(\mem[5][12] ), .A2(n712), .ZN(n699) );
  OAI21_X1 U136 ( .B1(n476), .B2(n460), .A(n698), .ZN(n536) );
  NAND2_X1 U137 ( .A1(\mem[5][13] ), .A2(n712), .ZN(n698) );
  OAI21_X1 U138 ( .B1(n475), .B2(n712), .A(n697), .ZN(n535) );
  NAND2_X1 U139 ( .A1(\mem[5][14] ), .A2(n712), .ZN(n697) );
  OAI21_X1 U140 ( .B1(n474), .B2(n460), .A(n696), .ZN(n534) );
  NAND2_X1 U141 ( .A1(\mem[5][15] ), .A2(n712), .ZN(n696) );
  OAI21_X1 U142 ( .B1(n473), .B2(n460), .A(n695), .ZN(n533) );
  NAND2_X1 U143 ( .A1(\mem[5][16] ), .A2(n712), .ZN(n695) );
  OAI21_X1 U144 ( .B1(n472), .B2(n460), .A(n694), .ZN(n532) );
  NAND2_X1 U145 ( .A1(\mem[5][17] ), .A2(n712), .ZN(n694) );
  OAI21_X1 U146 ( .B1(n471), .B2(n460), .A(n693), .ZN(n531) );
  NAND2_X1 U147 ( .A1(\mem[5][18] ), .A2(n712), .ZN(n693) );
  OAI21_X1 U148 ( .B1(n470), .B2(n460), .A(n692), .ZN(n530) );
  NAND2_X1 U149 ( .A1(\mem[5][19] ), .A2(n712), .ZN(n692) );
  OAI21_X1 U150 ( .B1(n489), .B2(n691), .A(n690), .ZN(n529) );
  NAND2_X1 U151 ( .A1(\mem[6][0] ), .A2(n459), .ZN(n690) );
  OAI21_X1 U152 ( .B1(n488), .B2(n691), .A(n689), .ZN(n528) );
  NAND2_X1 U153 ( .A1(\mem[6][1] ), .A2(n459), .ZN(n689) );
  OAI21_X1 U154 ( .B1(n487), .B2(n691), .A(n688), .ZN(n527) );
  NAND2_X1 U155 ( .A1(\mem[6][2] ), .A2(n459), .ZN(n688) );
  OAI21_X1 U156 ( .B1(n486), .B2(n691), .A(n687), .ZN(n526) );
  NAND2_X1 U157 ( .A1(\mem[6][3] ), .A2(n459), .ZN(n687) );
  OAI21_X1 U158 ( .B1(n485), .B2(n459), .A(n686), .ZN(n525) );
  NAND2_X1 U159 ( .A1(\mem[6][4] ), .A2(n459), .ZN(n686) );
  OAI21_X1 U160 ( .B1(n484), .B2(n691), .A(n685), .ZN(n524) );
  NAND2_X1 U161 ( .A1(\mem[6][5] ), .A2(n459), .ZN(n685) );
  OAI21_X1 U162 ( .B1(n483), .B2(n691), .A(n684), .ZN(n523) );
  NAND2_X1 U163 ( .A1(\mem[6][6] ), .A2(n459), .ZN(n684) );
  OAI21_X1 U164 ( .B1(n482), .B2(n691), .A(n683), .ZN(n522) );
  NAND2_X1 U165 ( .A1(\mem[6][7] ), .A2(n459), .ZN(n683) );
  OAI21_X1 U166 ( .B1(n481), .B2(n691), .A(n682), .ZN(n521) );
  NAND2_X1 U167 ( .A1(\mem[6][8] ), .A2(n459), .ZN(n682) );
  OAI21_X1 U168 ( .B1(n480), .B2(n691), .A(n681), .ZN(n520) );
  NAND2_X1 U169 ( .A1(\mem[6][9] ), .A2(n459), .ZN(n681) );
  OAI21_X1 U170 ( .B1(n479), .B2(n691), .A(n680), .ZN(n519) );
  NAND2_X1 U171 ( .A1(\mem[6][10] ), .A2(n459), .ZN(n680) );
  OAI21_X1 U172 ( .B1(n478), .B2(n691), .A(n679), .ZN(n518) );
  NAND2_X1 U173 ( .A1(\mem[6][11] ), .A2(n459), .ZN(n679) );
  OAI21_X1 U174 ( .B1(n477), .B2(n691), .A(n678), .ZN(n517) );
  NAND2_X1 U175 ( .A1(\mem[6][12] ), .A2(n691), .ZN(n678) );
  OAI21_X1 U176 ( .B1(n476), .B2(n459), .A(n677), .ZN(n516) );
  NAND2_X1 U177 ( .A1(\mem[6][13] ), .A2(n691), .ZN(n677) );
  OAI21_X1 U178 ( .B1(n475), .B2(n459), .A(n676), .ZN(n515) );
  NAND2_X1 U179 ( .A1(\mem[6][14] ), .A2(n691), .ZN(n676) );
  OAI21_X1 U180 ( .B1(n474), .B2(n691), .A(n675), .ZN(n514) );
  NAND2_X1 U181 ( .A1(\mem[6][15] ), .A2(n691), .ZN(n675) );
  OAI21_X1 U182 ( .B1(n473), .B2(n691), .A(n674), .ZN(n513) );
  NAND2_X1 U183 ( .A1(\mem[6][16] ), .A2(n691), .ZN(n674) );
  OAI21_X1 U184 ( .B1(n472), .B2(n691), .A(n673), .ZN(n512) );
  NAND2_X1 U185 ( .A1(\mem[6][17] ), .A2(n691), .ZN(n673) );
  OAI21_X1 U186 ( .B1(n471), .B2(n691), .A(n672), .ZN(n511) );
  NAND2_X1 U187 ( .A1(\mem[6][18] ), .A2(n691), .ZN(n672) );
  OAI21_X1 U188 ( .B1(n470), .B2(n691), .A(n671), .ZN(n510) );
  NAND2_X1 U189 ( .A1(\mem[6][19] ), .A2(n459), .ZN(n671) );
  OAI21_X1 U190 ( .B1(n489), .B2(n670), .A(n669), .ZN(n509) );
  NAND2_X1 U191 ( .A1(\mem[7][0] ), .A2(n458), .ZN(n669) );
  OAI21_X1 U192 ( .B1(n488), .B2(n670), .A(n668), .ZN(n508) );
  NAND2_X1 U193 ( .A1(\mem[7][1] ), .A2(n458), .ZN(n668) );
  OAI21_X1 U194 ( .B1(n487), .B2(n670), .A(n667), .ZN(n507) );
  NAND2_X1 U195 ( .A1(\mem[7][2] ), .A2(n458), .ZN(n667) );
  OAI21_X1 U196 ( .B1(n486), .B2(n670), .A(n666), .ZN(n506) );
  NAND2_X1 U197 ( .A1(\mem[7][3] ), .A2(n458), .ZN(n666) );
  OAI21_X1 U198 ( .B1(n485), .B2(n458), .A(n665), .ZN(n505) );
  NAND2_X1 U199 ( .A1(\mem[7][4] ), .A2(n458), .ZN(n665) );
  OAI21_X1 U200 ( .B1(n484), .B2(n670), .A(n664), .ZN(n504) );
  NAND2_X1 U201 ( .A1(\mem[7][5] ), .A2(n458), .ZN(n664) );
  OAI21_X1 U202 ( .B1(n483), .B2(n670), .A(n663), .ZN(n503) );
  NAND2_X1 U203 ( .A1(\mem[7][6] ), .A2(n458), .ZN(n663) );
  OAI21_X1 U204 ( .B1(n482), .B2(n670), .A(n662), .ZN(n502) );
  NAND2_X1 U205 ( .A1(\mem[7][7] ), .A2(n458), .ZN(n662) );
  OAI21_X1 U206 ( .B1(n481), .B2(n670), .A(n661), .ZN(n501) );
  NAND2_X1 U207 ( .A1(\mem[7][8] ), .A2(n458), .ZN(n661) );
  OAI21_X1 U208 ( .B1(n480), .B2(n670), .A(n660), .ZN(n500) );
  NAND2_X1 U209 ( .A1(\mem[7][9] ), .A2(n458), .ZN(n660) );
  OAI21_X1 U210 ( .B1(n479), .B2(n670), .A(n659), .ZN(n499) );
  NAND2_X1 U211 ( .A1(\mem[7][10] ), .A2(n458), .ZN(n659) );
  OAI21_X1 U212 ( .B1(n478), .B2(n670), .A(n658), .ZN(n498) );
  NAND2_X1 U213 ( .A1(\mem[7][11] ), .A2(n458), .ZN(n658) );
  OAI21_X1 U214 ( .B1(n477), .B2(n670), .A(n657), .ZN(n497) );
  NAND2_X1 U215 ( .A1(\mem[7][12] ), .A2(n670), .ZN(n657) );
  OAI21_X1 U216 ( .B1(n476), .B2(n458), .A(n656), .ZN(n496) );
  NAND2_X1 U217 ( .A1(\mem[7][13] ), .A2(n670), .ZN(n656) );
  OAI21_X1 U218 ( .B1(n475), .B2(n458), .A(n655), .ZN(n495) );
  NAND2_X1 U219 ( .A1(\mem[7][14] ), .A2(n670), .ZN(n655) );
  OAI21_X1 U220 ( .B1(n474), .B2(n670), .A(n654), .ZN(n494) );
  NAND2_X1 U221 ( .A1(\mem[7][15] ), .A2(n670), .ZN(n654) );
  OAI21_X1 U222 ( .B1(n473), .B2(n670), .A(n653), .ZN(n493) );
  NAND2_X1 U223 ( .A1(\mem[7][16] ), .A2(n670), .ZN(n653) );
  OAI21_X1 U224 ( .B1(n472), .B2(n670), .A(n652), .ZN(n492) );
  NAND2_X1 U225 ( .A1(\mem[7][17] ), .A2(n670), .ZN(n652) );
  OAI21_X1 U226 ( .B1(n471), .B2(n670), .A(n651), .ZN(n491) );
  NAND2_X1 U227 ( .A1(\mem[7][18] ), .A2(n670), .ZN(n651) );
  OAI21_X1 U228 ( .B1(n470), .B2(n670), .A(n650), .ZN(n490) );
  NAND2_X1 U229 ( .A1(\mem[7][19] ), .A2(n458), .ZN(n650) );
  NAND2_X1 U230 ( .A1(wr_en), .A2(n469), .ZN(n735) );
  INV_X1 U231 ( .A(addr[3]), .ZN(n469) );
  OAI21_X1 U232 ( .B1(n820), .B2(n489), .A(n819), .ZN(n649) );
  NAND2_X1 U233 ( .A1(\mem[0][0] ), .A2(n820), .ZN(n819) );
  OAI21_X1 U234 ( .B1(n820), .B2(n488), .A(n818), .ZN(n648) );
  NAND2_X1 U235 ( .A1(\mem[0][1] ), .A2(n820), .ZN(n818) );
  OAI21_X1 U236 ( .B1(n820), .B2(n487), .A(n817), .ZN(n647) );
  NAND2_X1 U237 ( .A1(\mem[0][2] ), .A2(n465), .ZN(n817) );
  OAI21_X1 U238 ( .B1(n820), .B2(n486), .A(n816), .ZN(n646) );
  NAND2_X1 U239 ( .A1(\mem[0][3] ), .A2(n465), .ZN(n816) );
  OAI21_X1 U240 ( .B1(n820), .B2(n485), .A(n815), .ZN(n645) );
  NAND2_X1 U241 ( .A1(\mem[0][4] ), .A2(n465), .ZN(n815) );
  OAI21_X1 U242 ( .B1(n820), .B2(n484), .A(n814), .ZN(n644) );
  NAND2_X1 U243 ( .A1(\mem[0][5] ), .A2(n465), .ZN(n814) );
  OAI21_X1 U244 ( .B1(n820), .B2(n483), .A(n813), .ZN(n643) );
  NAND2_X1 U245 ( .A1(\mem[0][6] ), .A2(n465), .ZN(n813) );
  OAI21_X1 U246 ( .B1(n820), .B2(n482), .A(n812), .ZN(n642) );
  NAND2_X1 U247 ( .A1(\mem[0][7] ), .A2(n820), .ZN(n812) );
  OAI21_X1 U248 ( .B1(n820), .B2(n481), .A(n811), .ZN(n641) );
  NAND2_X1 U249 ( .A1(\mem[0][8] ), .A2(n820), .ZN(n811) );
  OAI21_X1 U250 ( .B1(n465), .B2(n480), .A(n810), .ZN(n640) );
  NAND2_X1 U251 ( .A1(\mem[0][9] ), .A2(n820), .ZN(n810) );
  OAI21_X1 U252 ( .B1(n820), .B2(n479), .A(n809), .ZN(n639) );
  NAND2_X1 U253 ( .A1(\mem[0][10] ), .A2(n820), .ZN(n809) );
  OAI21_X1 U254 ( .B1(n820), .B2(n478), .A(n808), .ZN(n638) );
  NAND2_X1 U255 ( .A1(\mem[0][11] ), .A2(n820), .ZN(n808) );
  OAI21_X1 U256 ( .B1(n489), .B2(n798), .A(n797), .ZN(n629) );
  NAND2_X1 U257 ( .A1(\mem[1][0] ), .A2(n464), .ZN(n797) );
  OAI21_X1 U258 ( .B1(n488), .B2(n798), .A(n796), .ZN(n628) );
  NAND2_X1 U259 ( .A1(\mem[1][1] ), .A2(n464), .ZN(n796) );
  OAI21_X1 U260 ( .B1(n487), .B2(n798), .A(n795), .ZN(n627) );
  NAND2_X1 U261 ( .A1(\mem[1][2] ), .A2(n464), .ZN(n795) );
  OAI21_X1 U262 ( .B1(n486), .B2(n798), .A(n794), .ZN(n626) );
  NAND2_X1 U263 ( .A1(\mem[1][3] ), .A2(n464), .ZN(n794) );
  OAI21_X1 U264 ( .B1(n485), .B2(n798), .A(n793), .ZN(n625) );
  NAND2_X1 U265 ( .A1(\mem[1][4] ), .A2(n464), .ZN(n793) );
  OAI21_X1 U266 ( .B1(n484), .B2(n798), .A(n792), .ZN(n624) );
  NAND2_X1 U267 ( .A1(\mem[1][5] ), .A2(n464), .ZN(n792) );
  OAI21_X1 U268 ( .B1(n483), .B2(n798), .A(n791), .ZN(n623) );
  NAND2_X1 U269 ( .A1(\mem[1][6] ), .A2(n464), .ZN(n791) );
  OAI21_X1 U270 ( .B1(n482), .B2(n798), .A(n790), .ZN(n622) );
  NAND2_X1 U271 ( .A1(\mem[1][7] ), .A2(n464), .ZN(n790) );
  OAI21_X1 U272 ( .B1(n481), .B2(n798), .A(n789), .ZN(n621) );
  NAND2_X1 U273 ( .A1(\mem[1][8] ), .A2(n464), .ZN(n789) );
  OAI21_X1 U274 ( .B1(n480), .B2(n464), .A(n788), .ZN(n620) );
  NAND2_X1 U275 ( .A1(\mem[1][9] ), .A2(n464), .ZN(n788) );
  OAI21_X1 U276 ( .B1(n479), .B2(n798), .A(n787), .ZN(n619) );
  NAND2_X1 U277 ( .A1(\mem[1][10] ), .A2(n464), .ZN(n787) );
  OAI21_X1 U278 ( .B1(n478), .B2(n798), .A(n786), .ZN(n618) );
  NAND2_X1 U279 ( .A1(\mem[1][11] ), .A2(n464), .ZN(n786) );
  OAI21_X1 U280 ( .B1(n489), .B2(n463), .A(n776), .ZN(n609) );
  NAND2_X1 U281 ( .A1(\mem[2][0] ), .A2(n777), .ZN(n776) );
  OAI21_X1 U282 ( .B1(n488), .B2(n463), .A(n775), .ZN(n608) );
  NAND2_X1 U283 ( .A1(\mem[2][1] ), .A2(n777), .ZN(n775) );
  OAI21_X1 U284 ( .B1(n487), .B2(n463), .A(n774), .ZN(n607) );
  NAND2_X1 U285 ( .A1(\mem[2][2] ), .A2(n777), .ZN(n774) );
  OAI21_X1 U286 ( .B1(n486), .B2(n463), .A(n773), .ZN(n606) );
  NAND2_X1 U287 ( .A1(\mem[2][3] ), .A2(n777), .ZN(n773) );
  OAI21_X1 U288 ( .B1(n485), .B2(n463), .A(n772), .ZN(n605) );
  NAND2_X1 U289 ( .A1(\mem[2][4] ), .A2(n777), .ZN(n772) );
  OAI21_X1 U290 ( .B1(n484), .B2(n463), .A(n771), .ZN(n604) );
  NAND2_X1 U291 ( .A1(\mem[2][5] ), .A2(n777), .ZN(n771) );
  OAI21_X1 U292 ( .B1(n483), .B2(n463), .A(n770), .ZN(n603) );
  NAND2_X1 U293 ( .A1(\mem[2][6] ), .A2(n777), .ZN(n770) );
  OAI21_X1 U294 ( .B1(n482), .B2(n463), .A(n769), .ZN(n602) );
  NAND2_X1 U295 ( .A1(\mem[2][7] ), .A2(n777), .ZN(n769) );
  OAI21_X1 U296 ( .B1(n481), .B2(n463), .A(n768), .ZN(n601) );
  NAND2_X1 U297 ( .A1(\mem[2][8] ), .A2(n777), .ZN(n768) );
  OAI21_X1 U298 ( .B1(n480), .B2(n777), .A(n767), .ZN(n600) );
  NAND2_X1 U299 ( .A1(\mem[2][9] ), .A2(n777), .ZN(n767) );
  OAI21_X1 U300 ( .B1(n479), .B2(n463), .A(n766), .ZN(n599) );
  NAND2_X1 U301 ( .A1(\mem[2][10] ), .A2(n777), .ZN(n766) );
  OAI21_X1 U302 ( .B1(n478), .B2(n463), .A(n765), .ZN(n598) );
  NAND2_X1 U303 ( .A1(\mem[2][11] ), .A2(n777), .ZN(n765) );
  OAI21_X1 U304 ( .B1(n489), .B2(n756), .A(n755), .ZN(n589) );
  NAND2_X1 U305 ( .A1(\mem[3][0] ), .A2(n462), .ZN(n755) );
  OAI21_X1 U306 ( .B1(n488), .B2(n756), .A(n754), .ZN(n588) );
  NAND2_X1 U307 ( .A1(\mem[3][1] ), .A2(n462), .ZN(n754) );
  OAI21_X1 U308 ( .B1(n487), .B2(n756), .A(n753), .ZN(n587) );
  NAND2_X1 U309 ( .A1(\mem[3][2] ), .A2(n462), .ZN(n753) );
  OAI21_X1 U310 ( .B1(n486), .B2(n756), .A(n752), .ZN(n586) );
  NAND2_X1 U311 ( .A1(\mem[3][3] ), .A2(n462), .ZN(n752) );
  OAI21_X1 U312 ( .B1(n485), .B2(n756), .A(n751), .ZN(n585) );
  NAND2_X1 U313 ( .A1(\mem[3][4] ), .A2(n462), .ZN(n751) );
  OAI21_X1 U314 ( .B1(n484), .B2(n756), .A(n750), .ZN(n584) );
  NAND2_X1 U315 ( .A1(\mem[3][5] ), .A2(n462), .ZN(n750) );
  OAI21_X1 U316 ( .B1(n483), .B2(n756), .A(n749), .ZN(n583) );
  NAND2_X1 U317 ( .A1(\mem[3][6] ), .A2(n462), .ZN(n749) );
  OAI21_X1 U318 ( .B1(n482), .B2(n756), .A(n748), .ZN(n582) );
  NAND2_X1 U319 ( .A1(\mem[3][7] ), .A2(n462), .ZN(n748) );
  OAI21_X1 U320 ( .B1(n481), .B2(n756), .A(n747), .ZN(n581) );
  NAND2_X1 U321 ( .A1(\mem[3][8] ), .A2(n462), .ZN(n747) );
  OAI21_X1 U322 ( .B1(n480), .B2(n462), .A(n746), .ZN(n580) );
  NAND2_X1 U323 ( .A1(\mem[3][9] ), .A2(n462), .ZN(n746) );
  OAI21_X1 U324 ( .B1(n479), .B2(n756), .A(n745), .ZN(n579) );
  NAND2_X1 U325 ( .A1(\mem[3][10] ), .A2(n462), .ZN(n745) );
  OAI21_X1 U326 ( .B1(n478), .B2(n756), .A(n744), .ZN(n578) );
  NAND2_X1 U327 ( .A1(\mem[3][11] ), .A2(n462), .ZN(n744) );
  OAI21_X1 U328 ( .B1(n465), .B2(n477), .A(n807), .ZN(n637) );
  NAND2_X1 U329 ( .A1(\mem[0][12] ), .A2(n465), .ZN(n807) );
  OAI21_X1 U330 ( .B1(n465), .B2(n476), .A(n806), .ZN(n636) );
  NAND2_X1 U331 ( .A1(\mem[0][13] ), .A2(n465), .ZN(n806) );
  OAI21_X1 U332 ( .B1(n465), .B2(n475), .A(n805), .ZN(n635) );
  NAND2_X1 U333 ( .A1(\mem[0][14] ), .A2(n465), .ZN(n805) );
  OAI21_X1 U334 ( .B1(n820), .B2(n474), .A(n804), .ZN(n634) );
  NAND2_X1 U335 ( .A1(\mem[0][15] ), .A2(n465), .ZN(n804) );
  OAI21_X1 U336 ( .B1(n820), .B2(n473), .A(n803), .ZN(n633) );
  NAND2_X1 U337 ( .A1(\mem[0][16] ), .A2(n465), .ZN(n803) );
  OAI21_X1 U338 ( .B1(n820), .B2(n472), .A(n802), .ZN(n632) );
  NAND2_X1 U339 ( .A1(\mem[0][17] ), .A2(n465), .ZN(n802) );
  OAI21_X1 U340 ( .B1(n820), .B2(n471), .A(n801), .ZN(n631) );
  NAND2_X1 U341 ( .A1(\mem[0][18] ), .A2(n465), .ZN(n801) );
  OAI21_X1 U342 ( .B1(n820), .B2(n470), .A(n800), .ZN(n630) );
  NAND2_X1 U343 ( .A1(\mem[0][19] ), .A2(n465), .ZN(n800) );
  INV_X1 U344 ( .A(data_in[0]), .ZN(n489) );
  INV_X1 U345 ( .A(data_in[1]), .ZN(n488) );
  INV_X1 U346 ( .A(data_in[2]), .ZN(n487) );
  INV_X1 U347 ( .A(data_in[3]), .ZN(n486) );
  INV_X1 U348 ( .A(data_in[4]), .ZN(n485) );
  INV_X1 U349 ( .A(data_in[5]), .ZN(n484) );
  INV_X1 U358 ( .A(data_in[6]), .ZN(n483) );
  INV_X1 U359 ( .A(data_in[7]), .ZN(n482) );
  INV_X1 U360 ( .A(data_in[8]), .ZN(n481) );
  INV_X1 U361 ( .A(data_in[9]), .ZN(n480) );
  INV_X1 U362 ( .A(data_in[10]), .ZN(n479) );
  INV_X1 U363 ( .A(data_in[11]), .ZN(n478) );
  INV_X1 U364 ( .A(data_in[12]), .ZN(n477) );
  INV_X1 U365 ( .A(data_in[13]), .ZN(n476) );
  INV_X1 U366 ( .A(data_in[14]), .ZN(n475) );
  INV_X1 U367 ( .A(data_in[15]), .ZN(n474) );
  INV_X1 U368 ( .A(data_in[16]), .ZN(n473) );
  INV_X1 U369 ( .A(data_in[17]), .ZN(n472) );
  INV_X1 U370 ( .A(data_in[18]), .ZN(n471) );
  INV_X1 U371 ( .A(data_in[19]), .ZN(n470) );
  MUX2_X1 U372 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n455), .Z(n1) );
  MUX2_X1 U373 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n454), .Z(n2) );
  MUX2_X1 U374 ( .A(n2), .B(n1), .S(n453), .Z(n3) );
  MUX2_X1 U375 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n456), .Z(n4) );
  MUX2_X1 U376 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n457), .Z(n5) );
  MUX2_X1 U377 ( .A(n5), .B(n4), .S(n453), .Z(n6) );
  MUX2_X1 U378 ( .A(n6), .B(n3), .S(N12), .Z(N32) );
  MUX2_X1 U379 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n455), .Z(n7) );
  MUX2_X1 U380 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n456), .Z(n8) );
  MUX2_X1 U381 ( .A(n8), .B(n7), .S(n453), .Z(n9) );
  MUX2_X1 U382 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n455), .Z(n10) );
  MUX2_X1 U383 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n455), .Z(n11) );
  MUX2_X1 U384 ( .A(n11), .B(n10), .S(n453), .Z(n12) );
  MUX2_X1 U385 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n454), .Z(n13) );
  MUX2_X1 U386 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n457), .Z(n14) );
  MUX2_X1 U387 ( .A(n14), .B(n13), .S(n453), .Z(n15) );
  MUX2_X1 U388 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n456), .Z(n16) );
  MUX2_X1 U389 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n454), .Z(n17) );
  MUX2_X1 U390 ( .A(n17), .B(n16), .S(n453), .Z(n18) );
  MUX2_X1 U391 ( .A(n18), .B(n15), .S(N12), .Z(N30) );
  MUX2_X1 U392 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n457), .Z(n19) );
  MUX2_X1 U393 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n455), .Z(n20) );
  MUX2_X1 U394 ( .A(n20), .B(n19), .S(n453), .Z(n21) );
  MUX2_X1 U395 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n454), .Z(n22) );
  MUX2_X1 U396 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n457), .Z(n23) );
  MUX2_X1 U397 ( .A(n23), .B(n22), .S(n453), .Z(n24) );
  MUX2_X1 U398 ( .A(n24), .B(n21), .S(N12), .Z(N29) );
  MUX2_X1 U399 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n456), .Z(n356) );
  MUX2_X1 U400 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n456), .Z(n357) );
  MUX2_X1 U401 ( .A(n357), .B(n356), .S(n453), .Z(n358) );
  MUX2_X1 U402 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n457), .Z(n359) );
  MUX2_X1 U403 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n456), .Z(n360) );
  MUX2_X1 U404 ( .A(n360), .B(n359), .S(n453), .Z(n361) );
  MUX2_X1 U405 ( .A(n361), .B(n358), .S(N12), .Z(N28) );
  MUX2_X1 U406 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n454), .Z(n362) );
  MUX2_X1 U407 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n454), .Z(n363) );
  MUX2_X1 U408 ( .A(n363), .B(n362), .S(n453), .Z(n364) );
  MUX2_X1 U409 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n454), .Z(n365) );
  MUX2_X1 U410 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n454), .Z(n366) );
  MUX2_X1 U411 ( .A(n366), .B(n365), .S(n453), .Z(n367) );
  MUX2_X1 U412 ( .A(n367), .B(n364), .S(N12), .Z(N27) );
  MUX2_X1 U413 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n454), .Z(n368) );
  MUX2_X1 U414 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n454), .Z(n369) );
  MUX2_X1 U415 ( .A(n369), .B(n368), .S(n453), .Z(n370) );
  MUX2_X1 U416 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n454), .Z(n371) );
  MUX2_X1 U417 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n454), .Z(n372) );
  MUX2_X1 U418 ( .A(n372), .B(n371), .S(n453), .Z(n373) );
  MUX2_X1 U419 ( .A(n373), .B(n370), .S(N12), .Z(N26) );
  MUX2_X1 U420 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n454), .Z(n374) );
  MUX2_X1 U421 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n454), .Z(n375) );
  MUX2_X1 U422 ( .A(n375), .B(n374), .S(n453), .Z(n376) );
  MUX2_X1 U423 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n454), .Z(n377) );
  MUX2_X1 U424 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n454), .Z(n378) );
  MUX2_X1 U425 ( .A(n378), .B(n377), .S(n453), .Z(n379) );
  MUX2_X1 U426 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n455), .Z(n380) );
  MUX2_X1 U427 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n455), .Z(n381) );
  MUX2_X1 U428 ( .A(n381), .B(n380), .S(n452), .Z(n382) );
  MUX2_X1 U429 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n455), .Z(n383) );
  MUX2_X1 U430 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n455), .Z(n384) );
  MUX2_X1 U431 ( .A(n384), .B(n383), .S(n452), .Z(n385) );
  MUX2_X1 U432 ( .A(n385), .B(n382), .S(N12), .Z(N24) );
  MUX2_X1 U433 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n455), .Z(n386) );
  MUX2_X1 U434 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n455), .Z(n387) );
  MUX2_X1 U435 ( .A(n387), .B(n386), .S(n452), .Z(n388) );
  MUX2_X1 U436 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n455), .Z(n389) );
  MUX2_X1 U437 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n455), .Z(n390) );
  MUX2_X1 U438 ( .A(n390), .B(n389), .S(n452), .Z(n391) );
  MUX2_X1 U439 ( .A(n391), .B(n388), .S(N12), .Z(N23) );
  MUX2_X1 U440 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n455), .Z(n392) );
  MUX2_X1 U441 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n455), .Z(n393) );
  MUX2_X1 U442 ( .A(n393), .B(n392), .S(n452), .Z(n394) );
  MUX2_X1 U443 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n455), .Z(n395) );
  MUX2_X1 U444 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n455), .Z(n396) );
  MUX2_X1 U445 ( .A(n396), .B(n395), .S(n452), .Z(n397) );
  MUX2_X1 U446 ( .A(n397), .B(n394), .S(N12), .Z(N22) );
  MUX2_X1 U447 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n456), .Z(n398) );
  MUX2_X1 U448 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n456), .Z(n399) );
  MUX2_X1 U449 ( .A(n399), .B(n398), .S(n452), .Z(n400) );
  MUX2_X1 U450 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n456), .Z(n401) );
  MUX2_X1 U451 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n456), .Z(n402) );
  MUX2_X1 U452 ( .A(n402), .B(n401), .S(n452), .Z(n403) );
  MUX2_X1 U453 ( .A(n403), .B(n400), .S(N12), .Z(N21) );
  MUX2_X1 U454 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n456), .Z(n404) );
  MUX2_X1 U455 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n456), .Z(n405) );
  MUX2_X1 U456 ( .A(n405), .B(n404), .S(n452), .Z(n406) );
  MUX2_X1 U457 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n456), .Z(n407) );
  MUX2_X1 U458 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n456), .Z(n408) );
  MUX2_X1 U459 ( .A(n408), .B(n407), .S(n452), .Z(n409) );
  MUX2_X1 U460 ( .A(n409), .B(n406), .S(N12), .Z(N20) );
  MUX2_X1 U461 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n456), .Z(n410) );
  MUX2_X1 U462 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n456), .Z(n411) );
  MUX2_X1 U463 ( .A(n411), .B(n410), .S(n452), .Z(n412) );
  MUX2_X1 U464 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n456), .Z(n413) );
  MUX2_X1 U465 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n456), .Z(n414) );
  MUX2_X1 U466 ( .A(n414), .B(n413), .S(n452), .Z(n415) );
  MUX2_X1 U467 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n457), .Z(n416) );
  MUX2_X1 U468 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n457), .Z(n417) );
  MUX2_X1 U469 ( .A(n417), .B(n416), .S(n453), .Z(n418) );
  MUX2_X1 U470 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n457), .Z(n419) );
  MUX2_X1 U471 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n457), .Z(n420) );
  MUX2_X1 U472 ( .A(n420), .B(n419), .S(n453), .Z(n421) );
  MUX2_X1 U473 ( .A(n421), .B(n418), .S(N12), .Z(N18) );
  MUX2_X1 U474 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n457), .Z(n422) );
  MUX2_X1 U475 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n457), .Z(n423) );
  MUX2_X1 U476 ( .A(n423), .B(n422), .S(N11), .Z(n424) );
  MUX2_X1 U477 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n457), .Z(n425) );
  MUX2_X1 U478 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n457), .Z(n426) );
  MUX2_X1 U479 ( .A(n426), .B(n425), .S(N11), .Z(n427) );
  MUX2_X1 U480 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n457), .Z(n428) );
  MUX2_X1 U481 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n457), .Z(n429) );
  MUX2_X1 U482 ( .A(n429), .B(n428), .S(n453), .Z(n430) );
  MUX2_X1 U483 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n457), .Z(n431) );
  MUX2_X1 U484 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n457), .Z(n432) );
  MUX2_X1 U485 ( .A(n432), .B(n431), .S(n453), .Z(n433) );
  MUX2_X1 U486 ( .A(n433), .B(n430), .S(N12), .Z(N16) );
  MUX2_X1 U487 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n456), .Z(n434) );
  MUX2_X1 U488 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n455), .Z(n435) );
  MUX2_X1 U489 ( .A(n435), .B(n434), .S(N11), .Z(n436) );
  MUX2_X1 U490 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n454), .Z(n437) );
  MUX2_X1 U491 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n457), .Z(n438) );
  MUX2_X1 U492 ( .A(n438), .B(n437), .S(N11), .Z(n439) );
  MUX2_X1 U493 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n454), .Z(n440) );
  MUX2_X1 U494 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n455), .Z(n441) );
  MUX2_X1 U495 ( .A(n441), .B(n440), .S(n453), .Z(n442) );
  MUX2_X1 U496 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n455), .Z(n443) );
  MUX2_X1 U497 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n457), .Z(n444) );
  MUX2_X1 U498 ( .A(n444), .B(n443), .S(N11), .Z(n445) );
  MUX2_X1 U499 ( .A(n445), .B(n442), .S(N12), .Z(N14) );
  MUX2_X1 U500 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n457), .Z(n446) );
  MUX2_X1 U501 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n454), .Z(n447) );
  MUX2_X1 U502 ( .A(n447), .B(n446), .S(n453), .Z(n448) );
  MUX2_X1 U503 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n454), .Z(n449) );
  MUX2_X1 U504 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n456), .Z(n450) );
  MUX2_X1 U505 ( .A(n450), .B(n449), .S(N11), .Z(n451) );
  MUX2_X1 U506 ( .A(n451), .B(n448), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE4_1 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N13, N14, N15, N16, N18, N24, N26, N28, N30, N32, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[19]  ( .D(N13), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[17]  ( .D(N15), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N30), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N32), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n490), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n491), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n492), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n493), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n494), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n495), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n496), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n497), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n498), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n499), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n500), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n501), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n502), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n503), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n504), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n505), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n506), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n507), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n508), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n509), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n510), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n511), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n512), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n513), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n514), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n515), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n516), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n517), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n518), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n519), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n520), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n521), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n522), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n523), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n524), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n525), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n526), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n527), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n528), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n529), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n530), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n531), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n532), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n533), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n534), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n535), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n536), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n537), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n538), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n539), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n540), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n541), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n542), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n543), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n544), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n545), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n546), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n547), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n548), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n549), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n550), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n551), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n552), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n553), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n554), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n555), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n556), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n557), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n558), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n559), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n560), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n561), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n562), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n563), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n564), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n565), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n566), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n567), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n568), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n569), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n570), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n571), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n572), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n573), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n574), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n575), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n576), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n577), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n578), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n579), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n580), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n581), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n582), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n583), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n584), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n585), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n586), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n587), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n588), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n589), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n590), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n591), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n592), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n593), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n594), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n595), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n596), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n597), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n598), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n599), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n600), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n601), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n602), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n603), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n604), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n605), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n606), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n607), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n608), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n609), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n610), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n611), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n612), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n613), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n614), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n615), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n616), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n617), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n618), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n619), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n620), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n621), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n622), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n623), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n624), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n625), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n626), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n627), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n628), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n629), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n630), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n631), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n632), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n633), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n634), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n635), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n636), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n637), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n638), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n639), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n640), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n641), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n642), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n643), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n644), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n645), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n646), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n647), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n648), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n649), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U350 ( .A1(n466), .A2(n467), .A3(n799), .ZN(n820) );
  NAND3_X1 U351 ( .A1(n799), .A2(n467), .A3(N10), .ZN(n798) );
  NAND3_X1 U352 ( .A1(n799), .A2(n466), .A3(N11), .ZN(n777) );
  NAND3_X1 U353 ( .A1(N10), .A2(n799), .A3(N11), .ZN(n756) );
  NAND3_X1 U354 ( .A1(n466), .A2(n467), .A3(n713), .ZN(n734) );
  NAND3_X1 U355 ( .A1(N10), .A2(n467), .A3(n713), .ZN(n712) );
  NAND3_X1 U356 ( .A1(N11), .A2(n466), .A3(n713), .ZN(n691) );
  NAND3_X1 U357 ( .A1(N11), .A2(N10), .A3(n713), .ZN(n670) );
  SDFF_X1 \data_out_reg[13]  ( .D(n412), .SI(n415), .SE(n468), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n424), .SI(n427), .SE(n468), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[12]  ( .D(n406), .SI(n409), .SE(n468), .CK(clk), .Q(
        data_out[12]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n376), .SI(n379), .SE(n468), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n364), .SI(n367), .SE(n468), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[10]  ( .D(n394), .SI(n397), .SE(n468), .CK(clk), .Q(
        data_out[10]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n388), .SI(n391), .SE(n468), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n21), .SI(n24), .SE(n468), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n400), .SI(n403), .SE(n468), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n9), .SI(n12), .SE(n468), .CK(clk), .Q(
        data_out[1]) );
  BUF_X1 U3 ( .A(n820), .Z(n465) );
  BUF_X1 U4 ( .A(n777), .Z(n463) );
  BUF_X1 U5 ( .A(n712), .Z(n460) );
  BUF_X1 U6 ( .A(n453), .Z(n452) );
  BUF_X1 U7 ( .A(N10), .Z(n454) );
  BUF_X1 U8 ( .A(N10), .Z(n455) );
  BUF_X1 U9 ( .A(N10), .Z(n456) );
  BUF_X1 U10 ( .A(N10), .Z(n457) );
  BUF_X1 U11 ( .A(n756), .Z(n462) );
  BUF_X1 U12 ( .A(n798), .Z(n464) );
  BUF_X1 U13 ( .A(n670), .Z(n458) );
  BUF_X1 U14 ( .A(n734), .Z(n461) );
  BUF_X1 U15 ( .A(n691), .Z(n459) );
  BUF_X1 U16 ( .A(N11), .Z(n453) );
  NOR2_X1 U17 ( .A1(n735), .A2(N12), .ZN(n799) );
  NOR2_X1 U18 ( .A1(n468), .A2(n735), .ZN(n713) );
  INV_X1 U19 ( .A(N12), .ZN(n468) );
  INV_X1 U20 ( .A(N11), .ZN(n467) );
  INV_X1 U21 ( .A(N10), .ZN(n466) );
  OAI21_X1 U22 ( .B1(n477), .B2(n798), .A(n785), .ZN(n617) );
  NAND2_X1 U23 ( .A1(\mem[1][12] ), .A2(n798), .ZN(n785) );
  OAI21_X1 U24 ( .B1(n476), .B2(n798), .A(n784), .ZN(n616) );
  NAND2_X1 U25 ( .A1(\mem[1][13] ), .A2(n798), .ZN(n784) );
  OAI21_X1 U26 ( .B1(n475), .B2(n798), .A(n783), .ZN(n615) );
  NAND2_X1 U27 ( .A1(\mem[1][14] ), .A2(n798), .ZN(n783) );
  OAI21_X1 U28 ( .B1(n474), .B2(n464), .A(n782), .ZN(n614) );
  NAND2_X1 U29 ( .A1(\mem[1][15] ), .A2(n798), .ZN(n782) );
  OAI21_X1 U30 ( .B1(n473), .B2(n798), .A(n781), .ZN(n613) );
  NAND2_X1 U31 ( .A1(\mem[1][16] ), .A2(n464), .ZN(n781) );
  OAI21_X1 U32 ( .B1(n472), .B2(n798), .A(n780), .ZN(n612) );
  NAND2_X1 U33 ( .A1(\mem[1][17] ), .A2(n798), .ZN(n780) );
  OAI21_X1 U34 ( .B1(n471), .B2(n798), .A(n779), .ZN(n611) );
  NAND2_X1 U35 ( .A1(\mem[1][18] ), .A2(n798), .ZN(n779) );
  OAI21_X1 U36 ( .B1(n470), .B2(n798), .A(n778), .ZN(n610) );
  NAND2_X1 U37 ( .A1(\mem[1][19] ), .A2(n464), .ZN(n778) );
  OAI21_X1 U38 ( .B1(n477), .B2(n777), .A(n764), .ZN(n597) );
  NAND2_X1 U39 ( .A1(\mem[2][12] ), .A2(n777), .ZN(n764) );
  OAI21_X1 U40 ( .B1(n476), .B2(n777), .A(n763), .ZN(n596) );
  NAND2_X1 U41 ( .A1(\mem[2][13] ), .A2(n777), .ZN(n763) );
  OAI21_X1 U42 ( .B1(n475), .B2(n463), .A(n762), .ZN(n595) );
  NAND2_X1 U43 ( .A1(\mem[2][14] ), .A2(n777), .ZN(n762) );
  OAI21_X1 U44 ( .B1(n474), .B2(n463), .A(n761), .ZN(n594) );
  NAND2_X1 U45 ( .A1(\mem[2][15] ), .A2(n777), .ZN(n761) );
  OAI21_X1 U46 ( .B1(n473), .B2(n463), .A(n760), .ZN(n593) );
  NAND2_X1 U47 ( .A1(\mem[2][16] ), .A2(n777), .ZN(n760) );
  OAI21_X1 U48 ( .B1(n472), .B2(n463), .A(n759), .ZN(n592) );
  NAND2_X1 U49 ( .A1(\mem[2][17] ), .A2(n777), .ZN(n759) );
  OAI21_X1 U50 ( .B1(n471), .B2(n463), .A(n758), .ZN(n591) );
  NAND2_X1 U51 ( .A1(\mem[2][18] ), .A2(n777), .ZN(n758) );
  OAI21_X1 U52 ( .B1(n470), .B2(n777), .A(n757), .ZN(n590) );
  NAND2_X1 U53 ( .A1(\mem[2][19] ), .A2(n777), .ZN(n757) );
  OAI21_X1 U54 ( .B1(n477), .B2(n756), .A(n743), .ZN(n577) );
  NAND2_X1 U55 ( .A1(\mem[3][12] ), .A2(n756), .ZN(n743) );
  OAI21_X1 U56 ( .B1(n476), .B2(n756), .A(n742), .ZN(n576) );
  NAND2_X1 U57 ( .A1(\mem[3][13] ), .A2(n756), .ZN(n742) );
  OAI21_X1 U58 ( .B1(n475), .B2(n756), .A(n741), .ZN(n575) );
  NAND2_X1 U59 ( .A1(\mem[3][14] ), .A2(n756), .ZN(n741) );
  OAI21_X1 U60 ( .B1(n474), .B2(n462), .A(n740), .ZN(n574) );
  NAND2_X1 U61 ( .A1(\mem[3][15] ), .A2(n756), .ZN(n740) );
  OAI21_X1 U62 ( .B1(n473), .B2(n756), .A(n739), .ZN(n573) );
  NAND2_X1 U63 ( .A1(\mem[3][16] ), .A2(n462), .ZN(n739) );
  OAI21_X1 U64 ( .B1(n472), .B2(n756), .A(n738), .ZN(n572) );
  NAND2_X1 U65 ( .A1(\mem[3][17] ), .A2(n756), .ZN(n738) );
  OAI21_X1 U66 ( .B1(n471), .B2(n756), .A(n737), .ZN(n571) );
  NAND2_X1 U67 ( .A1(\mem[3][18] ), .A2(n756), .ZN(n737) );
  OAI21_X1 U68 ( .B1(n470), .B2(n756), .A(n736), .ZN(n570) );
  NAND2_X1 U69 ( .A1(\mem[3][19] ), .A2(n462), .ZN(n736) );
  OAI21_X1 U70 ( .B1(n489), .B2(n734), .A(n733), .ZN(n569) );
  NAND2_X1 U71 ( .A1(\mem[4][0] ), .A2(n461), .ZN(n733) );
  OAI21_X1 U72 ( .B1(n488), .B2(n734), .A(n732), .ZN(n568) );
  NAND2_X1 U73 ( .A1(\mem[4][1] ), .A2(n461), .ZN(n732) );
  OAI21_X1 U74 ( .B1(n487), .B2(n734), .A(n731), .ZN(n567) );
  NAND2_X1 U75 ( .A1(\mem[4][2] ), .A2(n461), .ZN(n731) );
  OAI21_X1 U76 ( .B1(n486), .B2(n734), .A(n730), .ZN(n566) );
  NAND2_X1 U77 ( .A1(\mem[4][3] ), .A2(n461), .ZN(n730) );
  OAI21_X1 U78 ( .B1(n485), .B2(n461), .A(n729), .ZN(n565) );
  NAND2_X1 U79 ( .A1(\mem[4][4] ), .A2(n461), .ZN(n729) );
  OAI21_X1 U80 ( .B1(n484), .B2(n734), .A(n728), .ZN(n564) );
  NAND2_X1 U81 ( .A1(\mem[4][5] ), .A2(n461), .ZN(n728) );
  OAI21_X1 U82 ( .B1(n483), .B2(n734), .A(n727), .ZN(n563) );
  NAND2_X1 U83 ( .A1(\mem[4][6] ), .A2(n461), .ZN(n727) );
  OAI21_X1 U84 ( .B1(n482), .B2(n734), .A(n726), .ZN(n562) );
  NAND2_X1 U85 ( .A1(\mem[4][7] ), .A2(n461), .ZN(n726) );
  OAI21_X1 U86 ( .B1(n481), .B2(n734), .A(n725), .ZN(n561) );
  NAND2_X1 U87 ( .A1(\mem[4][8] ), .A2(n461), .ZN(n725) );
  OAI21_X1 U88 ( .B1(n480), .B2(n734), .A(n724), .ZN(n560) );
  NAND2_X1 U89 ( .A1(\mem[4][9] ), .A2(n461), .ZN(n724) );
  OAI21_X1 U90 ( .B1(n479), .B2(n734), .A(n723), .ZN(n559) );
  NAND2_X1 U91 ( .A1(\mem[4][10] ), .A2(n461), .ZN(n723) );
  OAI21_X1 U92 ( .B1(n478), .B2(n734), .A(n722), .ZN(n558) );
  NAND2_X1 U93 ( .A1(\mem[4][11] ), .A2(n461), .ZN(n722) );
  OAI21_X1 U94 ( .B1(n477), .B2(n734), .A(n721), .ZN(n557) );
  NAND2_X1 U95 ( .A1(\mem[4][12] ), .A2(n734), .ZN(n721) );
  OAI21_X1 U96 ( .B1(n476), .B2(n461), .A(n720), .ZN(n556) );
  NAND2_X1 U97 ( .A1(\mem[4][13] ), .A2(n734), .ZN(n720) );
  OAI21_X1 U98 ( .B1(n475), .B2(n461), .A(n719), .ZN(n555) );
  NAND2_X1 U99 ( .A1(\mem[4][14] ), .A2(n734), .ZN(n719) );
  OAI21_X1 U100 ( .B1(n474), .B2(n734), .A(n718), .ZN(n554) );
  NAND2_X1 U101 ( .A1(\mem[4][15] ), .A2(n734), .ZN(n718) );
  OAI21_X1 U102 ( .B1(n473), .B2(n734), .A(n717), .ZN(n553) );
  NAND2_X1 U103 ( .A1(\mem[4][16] ), .A2(n734), .ZN(n717) );
  OAI21_X1 U104 ( .B1(n472), .B2(n734), .A(n716), .ZN(n552) );
  NAND2_X1 U105 ( .A1(\mem[4][17] ), .A2(n734), .ZN(n716) );
  OAI21_X1 U106 ( .B1(n471), .B2(n734), .A(n715), .ZN(n551) );
  NAND2_X1 U107 ( .A1(\mem[4][18] ), .A2(n734), .ZN(n715) );
  OAI21_X1 U108 ( .B1(n470), .B2(n734), .A(n714), .ZN(n550) );
  NAND2_X1 U109 ( .A1(\mem[4][19] ), .A2(n461), .ZN(n714) );
  OAI21_X1 U110 ( .B1(n489), .B2(n712), .A(n711), .ZN(n549) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n712), .ZN(n711) );
  OAI21_X1 U112 ( .B1(n488), .B2(n460), .A(n710), .ZN(n548) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n712), .ZN(n710) );
  OAI21_X1 U114 ( .B1(n487), .B2(n460), .A(n709), .ZN(n547) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n712), .ZN(n709) );
  OAI21_X1 U116 ( .B1(n486), .B2(n460), .A(n708), .ZN(n546) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n712), .ZN(n708) );
  OAI21_X1 U118 ( .B1(n485), .B2(n460), .A(n707), .ZN(n545) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n712), .ZN(n707) );
  OAI21_X1 U120 ( .B1(n484), .B2(n460), .A(n706), .ZN(n544) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n712), .ZN(n706) );
  OAI21_X1 U122 ( .B1(n483), .B2(n460), .A(n705), .ZN(n543) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n712), .ZN(n705) );
  OAI21_X1 U124 ( .B1(n482), .B2(n460), .A(n704), .ZN(n542) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n712), .ZN(n704) );
  OAI21_X1 U126 ( .B1(n481), .B2(n460), .A(n703), .ZN(n541) );
  NAND2_X1 U127 ( .A1(\mem[5][8] ), .A2(n712), .ZN(n703) );
  OAI21_X1 U128 ( .B1(n480), .B2(n712), .A(n702), .ZN(n540) );
  NAND2_X1 U129 ( .A1(\mem[5][9] ), .A2(n712), .ZN(n702) );
  OAI21_X1 U130 ( .B1(n479), .B2(n460), .A(n701), .ZN(n539) );
  NAND2_X1 U131 ( .A1(\mem[5][10] ), .A2(n712), .ZN(n701) );
  OAI21_X1 U132 ( .B1(n478), .B2(n460), .A(n700), .ZN(n538) );
  NAND2_X1 U133 ( .A1(\mem[5][11] ), .A2(n712), .ZN(n700) );
  OAI21_X1 U134 ( .B1(n477), .B2(n712), .A(n699), .ZN(n537) );
  NAND2_X1 U135 ( .A1(\mem[5][12] ), .A2(n712), .ZN(n699) );
  OAI21_X1 U136 ( .B1(n476), .B2(n460), .A(n698), .ZN(n536) );
  NAND2_X1 U137 ( .A1(\mem[5][13] ), .A2(n712), .ZN(n698) );
  OAI21_X1 U138 ( .B1(n475), .B2(n712), .A(n697), .ZN(n535) );
  NAND2_X1 U139 ( .A1(\mem[5][14] ), .A2(n712), .ZN(n697) );
  OAI21_X1 U140 ( .B1(n474), .B2(n460), .A(n696), .ZN(n534) );
  NAND2_X1 U141 ( .A1(\mem[5][15] ), .A2(n712), .ZN(n696) );
  OAI21_X1 U142 ( .B1(n473), .B2(n460), .A(n695), .ZN(n533) );
  NAND2_X1 U143 ( .A1(\mem[5][16] ), .A2(n712), .ZN(n695) );
  OAI21_X1 U144 ( .B1(n472), .B2(n460), .A(n694), .ZN(n532) );
  NAND2_X1 U145 ( .A1(\mem[5][17] ), .A2(n712), .ZN(n694) );
  OAI21_X1 U146 ( .B1(n471), .B2(n460), .A(n693), .ZN(n531) );
  NAND2_X1 U147 ( .A1(\mem[5][18] ), .A2(n712), .ZN(n693) );
  OAI21_X1 U148 ( .B1(n470), .B2(n460), .A(n692), .ZN(n530) );
  NAND2_X1 U149 ( .A1(\mem[5][19] ), .A2(n712), .ZN(n692) );
  OAI21_X1 U150 ( .B1(n489), .B2(n691), .A(n690), .ZN(n529) );
  NAND2_X1 U151 ( .A1(\mem[6][0] ), .A2(n459), .ZN(n690) );
  OAI21_X1 U152 ( .B1(n488), .B2(n691), .A(n689), .ZN(n528) );
  NAND2_X1 U153 ( .A1(\mem[6][1] ), .A2(n459), .ZN(n689) );
  OAI21_X1 U154 ( .B1(n487), .B2(n691), .A(n688), .ZN(n527) );
  NAND2_X1 U155 ( .A1(\mem[6][2] ), .A2(n459), .ZN(n688) );
  OAI21_X1 U156 ( .B1(n486), .B2(n691), .A(n687), .ZN(n526) );
  NAND2_X1 U157 ( .A1(\mem[6][3] ), .A2(n459), .ZN(n687) );
  OAI21_X1 U158 ( .B1(n485), .B2(n459), .A(n686), .ZN(n525) );
  NAND2_X1 U159 ( .A1(\mem[6][4] ), .A2(n459), .ZN(n686) );
  OAI21_X1 U160 ( .B1(n484), .B2(n691), .A(n685), .ZN(n524) );
  NAND2_X1 U161 ( .A1(\mem[6][5] ), .A2(n459), .ZN(n685) );
  OAI21_X1 U162 ( .B1(n483), .B2(n691), .A(n684), .ZN(n523) );
  NAND2_X1 U163 ( .A1(\mem[6][6] ), .A2(n459), .ZN(n684) );
  OAI21_X1 U164 ( .B1(n482), .B2(n691), .A(n683), .ZN(n522) );
  NAND2_X1 U165 ( .A1(\mem[6][7] ), .A2(n459), .ZN(n683) );
  OAI21_X1 U166 ( .B1(n481), .B2(n691), .A(n682), .ZN(n521) );
  NAND2_X1 U167 ( .A1(\mem[6][8] ), .A2(n459), .ZN(n682) );
  OAI21_X1 U168 ( .B1(n480), .B2(n691), .A(n681), .ZN(n520) );
  NAND2_X1 U169 ( .A1(\mem[6][9] ), .A2(n459), .ZN(n681) );
  OAI21_X1 U170 ( .B1(n479), .B2(n691), .A(n680), .ZN(n519) );
  NAND2_X1 U171 ( .A1(\mem[6][10] ), .A2(n459), .ZN(n680) );
  OAI21_X1 U172 ( .B1(n478), .B2(n691), .A(n679), .ZN(n518) );
  NAND2_X1 U173 ( .A1(\mem[6][11] ), .A2(n459), .ZN(n679) );
  OAI21_X1 U174 ( .B1(n477), .B2(n691), .A(n678), .ZN(n517) );
  NAND2_X1 U175 ( .A1(\mem[6][12] ), .A2(n691), .ZN(n678) );
  OAI21_X1 U176 ( .B1(n476), .B2(n459), .A(n677), .ZN(n516) );
  NAND2_X1 U177 ( .A1(\mem[6][13] ), .A2(n691), .ZN(n677) );
  OAI21_X1 U178 ( .B1(n475), .B2(n459), .A(n676), .ZN(n515) );
  NAND2_X1 U179 ( .A1(\mem[6][14] ), .A2(n691), .ZN(n676) );
  OAI21_X1 U180 ( .B1(n474), .B2(n691), .A(n675), .ZN(n514) );
  NAND2_X1 U181 ( .A1(\mem[6][15] ), .A2(n691), .ZN(n675) );
  OAI21_X1 U182 ( .B1(n473), .B2(n691), .A(n674), .ZN(n513) );
  NAND2_X1 U183 ( .A1(\mem[6][16] ), .A2(n691), .ZN(n674) );
  OAI21_X1 U184 ( .B1(n472), .B2(n691), .A(n673), .ZN(n512) );
  NAND2_X1 U185 ( .A1(\mem[6][17] ), .A2(n691), .ZN(n673) );
  OAI21_X1 U186 ( .B1(n471), .B2(n691), .A(n672), .ZN(n511) );
  NAND2_X1 U187 ( .A1(\mem[6][18] ), .A2(n691), .ZN(n672) );
  OAI21_X1 U188 ( .B1(n470), .B2(n691), .A(n671), .ZN(n510) );
  NAND2_X1 U189 ( .A1(\mem[6][19] ), .A2(n459), .ZN(n671) );
  OAI21_X1 U190 ( .B1(n489), .B2(n670), .A(n669), .ZN(n509) );
  NAND2_X1 U191 ( .A1(\mem[7][0] ), .A2(n458), .ZN(n669) );
  OAI21_X1 U192 ( .B1(n488), .B2(n670), .A(n668), .ZN(n508) );
  NAND2_X1 U193 ( .A1(\mem[7][1] ), .A2(n458), .ZN(n668) );
  OAI21_X1 U194 ( .B1(n487), .B2(n670), .A(n667), .ZN(n507) );
  NAND2_X1 U195 ( .A1(\mem[7][2] ), .A2(n458), .ZN(n667) );
  OAI21_X1 U196 ( .B1(n486), .B2(n670), .A(n666), .ZN(n506) );
  NAND2_X1 U197 ( .A1(\mem[7][3] ), .A2(n458), .ZN(n666) );
  OAI21_X1 U198 ( .B1(n485), .B2(n458), .A(n665), .ZN(n505) );
  NAND2_X1 U199 ( .A1(\mem[7][4] ), .A2(n458), .ZN(n665) );
  OAI21_X1 U200 ( .B1(n484), .B2(n670), .A(n664), .ZN(n504) );
  NAND2_X1 U201 ( .A1(\mem[7][5] ), .A2(n458), .ZN(n664) );
  OAI21_X1 U202 ( .B1(n483), .B2(n670), .A(n663), .ZN(n503) );
  NAND2_X1 U203 ( .A1(\mem[7][6] ), .A2(n458), .ZN(n663) );
  OAI21_X1 U204 ( .B1(n482), .B2(n670), .A(n662), .ZN(n502) );
  NAND2_X1 U205 ( .A1(\mem[7][7] ), .A2(n458), .ZN(n662) );
  OAI21_X1 U206 ( .B1(n481), .B2(n670), .A(n661), .ZN(n501) );
  NAND2_X1 U207 ( .A1(\mem[7][8] ), .A2(n458), .ZN(n661) );
  OAI21_X1 U208 ( .B1(n480), .B2(n670), .A(n660), .ZN(n500) );
  NAND2_X1 U209 ( .A1(\mem[7][9] ), .A2(n458), .ZN(n660) );
  OAI21_X1 U210 ( .B1(n479), .B2(n670), .A(n659), .ZN(n499) );
  NAND2_X1 U211 ( .A1(\mem[7][10] ), .A2(n458), .ZN(n659) );
  OAI21_X1 U212 ( .B1(n478), .B2(n670), .A(n658), .ZN(n498) );
  NAND2_X1 U213 ( .A1(\mem[7][11] ), .A2(n458), .ZN(n658) );
  OAI21_X1 U214 ( .B1(n477), .B2(n670), .A(n657), .ZN(n497) );
  NAND2_X1 U215 ( .A1(\mem[7][12] ), .A2(n670), .ZN(n657) );
  OAI21_X1 U216 ( .B1(n476), .B2(n458), .A(n656), .ZN(n496) );
  NAND2_X1 U217 ( .A1(\mem[7][13] ), .A2(n670), .ZN(n656) );
  OAI21_X1 U218 ( .B1(n475), .B2(n458), .A(n655), .ZN(n495) );
  NAND2_X1 U219 ( .A1(\mem[7][14] ), .A2(n670), .ZN(n655) );
  OAI21_X1 U220 ( .B1(n474), .B2(n670), .A(n654), .ZN(n494) );
  NAND2_X1 U221 ( .A1(\mem[7][15] ), .A2(n670), .ZN(n654) );
  OAI21_X1 U222 ( .B1(n473), .B2(n670), .A(n653), .ZN(n493) );
  NAND2_X1 U223 ( .A1(\mem[7][16] ), .A2(n670), .ZN(n653) );
  OAI21_X1 U224 ( .B1(n472), .B2(n670), .A(n652), .ZN(n492) );
  NAND2_X1 U225 ( .A1(\mem[7][17] ), .A2(n670), .ZN(n652) );
  OAI21_X1 U226 ( .B1(n471), .B2(n670), .A(n651), .ZN(n491) );
  NAND2_X1 U227 ( .A1(\mem[7][18] ), .A2(n670), .ZN(n651) );
  OAI21_X1 U228 ( .B1(n470), .B2(n670), .A(n650), .ZN(n490) );
  NAND2_X1 U229 ( .A1(\mem[7][19] ), .A2(n458), .ZN(n650) );
  NAND2_X1 U230 ( .A1(wr_en), .A2(n469), .ZN(n735) );
  INV_X1 U231 ( .A(addr[3]), .ZN(n469) );
  OAI21_X1 U232 ( .B1(n820), .B2(n489), .A(n819), .ZN(n649) );
  NAND2_X1 U233 ( .A1(\mem[0][0] ), .A2(n820), .ZN(n819) );
  OAI21_X1 U234 ( .B1(n820), .B2(n488), .A(n818), .ZN(n648) );
  NAND2_X1 U235 ( .A1(\mem[0][1] ), .A2(n820), .ZN(n818) );
  OAI21_X1 U236 ( .B1(n820), .B2(n487), .A(n817), .ZN(n647) );
  NAND2_X1 U237 ( .A1(\mem[0][2] ), .A2(n465), .ZN(n817) );
  OAI21_X1 U238 ( .B1(n820), .B2(n486), .A(n816), .ZN(n646) );
  NAND2_X1 U239 ( .A1(\mem[0][3] ), .A2(n465), .ZN(n816) );
  OAI21_X1 U240 ( .B1(n820), .B2(n485), .A(n815), .ZN(n645) );
  NAND2_X1 U241 ( .A1(\mem[0][4] ), .A2(n465), .ZN(n815) );
  OAI21_X1 U242 ( .B1(n820), .B2(n484), .A(n814), .ZN(n644) );
  NAND2_X1 U243 ( .A1(\mem[0][5] ), .A2(n465), .ZN(n814) );
  OAI21_X1 U244 ( .B1(n820), .B2(n483), .A(n813), .ZN(n643) );
  NAND2_X1 U245 ( .A1(\mem[0][6] ), .A2(n820), .ZN(n813) );
  OAI21_X1 U246 ( .B1(n820), .B2(n482), .A(n812), .ZN(n642) );
  NAND2_X1 U247 ( .A1(\mem[0][7] ), .A2(n820), .ZN(n812) );
  OAI21_X1 U248 ( .B1(n820), .B2(n481), .A(n811), .ZN(n641) );
  NAND2_X1 U249 ( .A1(\mem[0][8] ), .A2(n820), .ZN(n811) );
  OAI21_X1 U250 ( .B1(n465), .B2(n480), .A(n810), .ZN(n640) );
  NAND2_X1 U251 ( .A1(\mem[0][9] ), .A2(n820), .ZN(n810) );
  OAI21_X1 U252 ( .B1(n820), .B2(n479), .A(n809), .ZN(n639) );
  NAND2_X1 U253 ( .A1(\mem[0][10] ), .A2(n465), .ZN(n809) );
  OAI21_X1 U254 ( .B1(n820), .B2(n478), .A(n808), .ZN(n638) );
  NAND2_X1 U255 ( .A1(\mem[0][11] ), .A2(n820), .ZN(n808) );
  OAI21_X1 U256 ( .B1(n489), .B2(n798), .A(n797), .ZN(n629) );
  NAND2_X1 U257 ( .A1(\mem[1][0] ), .A2(n464), .ZN(n797) );
  OAI21_X1 U258 ( .B1(n488), .B2(n798), .A(n796), .ZN(n628) );
  NAND2_X1 U259 ( .A1(\mem[1][1] ), .A2(n464), .ZN(n796) );
  OAI21_X1 U260 ( .B1(n487), .B2(n798), .A(n795), .ZN(n627) );
  NAND2_X1 U261 ( .A1(\mem[1][2] ), .A2(n464), .ZN(n795) );
  OAI21_X1 U262 ( .B1(n486), .B2(n798), .A(n794), .ZN(n626) );
  NAND2_X1 U263 ( .A1(\mem[1][3] ), .A2(n464), .ZN(n794) );
  OAI21_X1 U264 ( .B1(n485), .B2(n798), .A(n793), .ZN(n625) );
  NAND2_X1 U265 ( .A1(\mem[1][4] ), .A2(n464), .ZN(n793) );
  OAI21_X1 U266 ( .B1(n484), .B2(n798), .A(n792), .ZN(n624) );
  NAND2_X1 U267 ( .A1(\mem[1][5] ), .A2(n464), .ZN(n792) );
  OAI21_X1 U268 ( .B1(n483), .B2(n798), .A(n791), .ZN(n623) );
  NAND2_X1 U269 ( .A1(\mem[1][6] ), .A2(n464), .ZN(n791) );
  OAI21_X1 U270 ( .B1(n482), .B2(n798), .A(n790), .ZN(n622) );
  NAND2_X1 U271 ( .A1(\mem[1][7] ), .A2(n464), .ZN(n790) );
  OAI21_X1 U272 ( .B1(n481), .B2(n798), .A(n789), .ZN(n621) );
  NAND2_X1 U273 ( .A1(\mem[1][8] ), .A2(n464), .ZN(n789) );
  OAI21_X1 U274 ( .B1(n480), .B2(n464), .A(n788), .ZN(n620) );
  NAND2_X1 U275 ( .A1(\mem[1][9] ), .A2(n464), .ZN(n788) );
  OAI21_X1 U276 ( .B1(n479), .B2(n798), .A(n787), .ZN(n619) );
  NAND2_X1 U277 ( .A1(\mem[1][10] ), .A2(n464), .ZN(n787) );
  OAI21_X1 U278 ( .B1(n478), .B2(n798), .A(n786), .ZN(n618) );
  NAND2_X1 U279 ( .A1(\mem[1][11] ), .A2(n464), .ZN(n786) );
  OAI21_X1 U280 ( .B1(n489), .B2(n463), .A(n776), .ZN(n609) );
  NAND2_X1 U281 ( .A1(\mem[2][0] ), .A2(n777), .ZN(n776) );
  OAI21_X1 U282 ( .B1(n488), .B2(n463), .A(n775), .ZN(n608) );
  NAND2_X1 U283 ( .A1(\mem[2][1] ), .A2(n777), .ZN(n775) );
  OAI21_X1 U284 ( .B1(n487), .B2(n463), .A(n774), .ZN(n607) );
  NAND2_X1 U285 ( .A1(\mem[2][2] ), .A2(n777), .ZN(n774) );
  OAI21_X1 U286 ( .B1(n486), .B2(n463), .A(n773), .ZN(n606) );
  NAND2_X1 U287 ( .A1(\mem[2][3] ), .A2(n777), .ZN(n773) );
  OAI21_X1 U288 ( .B1(n485), .B2(n463), .A(n772), .ZN(n605) );
  NAND2_X1 U289 ( .A1(\mem[2][4] ), .A2(n777), .ZN(n772) );
  OAI21_X1 U290 ( .B1(n484), .B2(n463), .A(n771), .ZN(n604) );
  NAND2_X1 U291 ( .A1(\mem[2][5] ), .A2(n777), .ZN(n771) );
  OAI21_X1 U292 ( .B1(n483), .B2(n463), .A(n770), .ZN(n603) );
  NAND2_X1 U293 ( .A1(\mem[2][6] ), .A2(n777), .ZN(n770) );
  OAI21_X1 U294 ( .B1(n482), .B2(n463), .A(n769), .ZN(n602) );
  NAND2_X1 U295 ( .A1(\mem[2][7] ), .A2(n777), .ZN(n769) );
  OAI21_X1 U296 ( .B1(n481), .B2(n463), .A(n768), .ZN(n601) );
  NAND2_X1 U297 ( .A1(\mem[2][8] ), .A2(n777), .ZN(n768) );
  OAI21_X1 U298 ( .B1(n480), .B2(n777), .A(n767), .ZN(n600) );
  NAND2_X1 U299 ( .A1(\mem[2][9] ), .A2(n777), .ZN(n767) );
  OAI21_X1 U300 ( .B1(n479), .B2(n463), .A(n766), .ZN(n599) );
  NAND2_X1 U301 ( .A1(\mem[2][10] ), .A2(n777), .ZN(n766) );
  OAI21_X1 U302 ( .B1(n478), .B2(n463), .A(n765), .ZN(n598) );
  NAND2_X1 U303 ( .A1(\mem[2][11] ), .A2(n777), .ZN(n765) );
  OAI21_X1 U304 ( .B1(n489), .B2(n756), .A(n755), .ZN(n589) );
  NAND2_X1 U305 ( .A1(\mem[3][0] ), .A2(n462), .ZN(n755) );
  OAI21_X1 U306 ( .B1(n488), .B2(n756), .A(n754), .ZN(n588) );
  NAND2_X1 U307 ( .A1(\mem[3][1] ), .A2(n462), .ZN(n754) );
  OAI21_X1 U308 ( .B1(n487), .B2(n756), .A(n753), .ZN(n587) );
  NAND2_X1 U309 ( .A1(\mem[3][2] ), .A2(n462), .ZN(n753) );
  OAI21_X1 U310 ( .B1(n486), .B2(n756), .A(n752), .ZN(n586) );
  NAND2_X1 U311 ( .A1(\mem[3][3] ), .A2(n462), .ZN(n752) );
  OAI21_X1 U312 ( .B1(n485), .B2(n756), .A(n751), .ZN(n585) );
  NAND2_X1 U313 ( .A1(\mem[3][4] ), .A2(n462), .ZN(n751) );
  OAI21_X1 U314 ( .B1(n484), .B2(n756), .A(n750), .ZN(n584) );
  NAND2_X1 U315 ( .A1(\mem[3][5] ), .A2(n462), .ZN(n750) );
  OAI21_X1 U316 ( .B1(n483), .B2(n756), .A(n749), .ZN(n583) );
  NAND2_X1 U317 ( .A1(\mem[3][6] ), .A2(n462), .ZN(n749) );
  OAI21_X1 U318 ( .B1(n482), .B2(n756), .A(n748), .ZN(n582) );
  NAND2_X1 U319 ( .A1(\mem[3][7] ), .A2(n462), .ZN(n748) );
  OAI21_X1 U320 ( .B1(n481), .B2(n756), .A(n747), .ZN(n581) );
  NAND2_X1 U321 ( .A1(\mem[3][8] ), .A2(n462), .ZN(n747) );
  OAI21_X1 U322 ( .B1(n480), .B2(n462), .A(n746), .ZN(n580) );
  NAND2_X1 U323 ( .A1(\mem[3][9] ), .A2(n462), .ZN(n746) );
  OAI21_X1 U324 ( .B1(n479), .B2(n756), .A(n745), .ZN(n579) );
  NAND2_X1 U325 ( .A1(\mem[3][10] ), .A2(n462), .ZN(n745) );
  OAI21_X1 U326 ( .B1(n478), .B2(n756), .A(n744), .ZN(n578) );
  NAND2_X1 U327 ( .A1(\mem[3][11] ), .A2(n462), .ZN(n744) );
  OAI21_X1 U328 ( .B1(n465), .B2(n477), .A(n807), .ZN(n637) );
  NAND2_X1 U329 ( .A1(\mem[0][12] ), .A2(n465), .ZN(n807) );
  OAI21_X1 U330 ( .B1(n465), .B2(n476), .A(n806), .ZN(n636) );
  NAND2_X1 U331 ( .A1(\mem[0][13] ), .A2(n465), .ZN(n806) );
  OAI21_X1 U332 ( .B1(n465), .B2(n475), .A(n805), .ZN(n635) );
  NAND2_X1 U333 ( .A1(\mem[0][14] ), .A2(n465), .ZN(n805) );
  OAI21_X1 U334 ( .B1(n820), .B2(n474), .A(n804), .ZN(n634) );
  NAND2_X1 U335 ( .A1(\mem[0][15] ), .A2(n465), .ZN(n804) );
  OAI21_X1 U336 ( .B1(n820), .B2(n473), .A(n803), .ZN(n633) );
  NAND2_X1 U337 ( .A1(\mem[0][16] ), .A2(n465), .ZN(n803) );
  OAI21_X1 U338 ( .B1(n820), .B2(n472), .A(n802), .ZN(n632) );
  NAND2_X1 U339 ( .A1(\mem[0][17] ), .A2(n465), .ZN(n802) );
  OAI21_X1 U340 ( .B1(n820), .B2(n471), .A(n801), .ZN(n631) );
  NAND2_X1 U341 ( .A1(\mem[0][18] ), .A2(n465), .ZN(n801) );
  OAI21_X1 U342 ( .B1(n820), .B2(n470), .A(n800), .ZN(n630) );
  NAND2_X1 U343 ( .A1(\mem[0][19] ), .A2(n465), .ZN(n800) );
  INV_X1 U344 ( .A(data_in[0]), .ZN(n489) );
  INV_X1 U345 ( .A(data_in[1]), .ZN(n488) );
  INV_X1 U346 ( .A(data_in[2]), .ZN(n487) );
  INV_X1 U347 ( .A(data_in[3]), .ZN(n486) );
  INV_X1 U348 ( .A(data_in[4]), .ZN(n485) );
  INV_X1 U349 ( .A(data_in[5]), .ZN(n484) );
  INV_X1 U358 ( .A(data_in[6]), .ZN(n483) );
  INV_X1 U359 ( .A(data_in[7]), .ZN(n482) );
  INV_X1 U360 ( .A(data_in[8]), .ZN(n481) );
  INV_X1 U361 ( .A(data_in[9]), .ZN(n480) );
  INV_X1 U362 ( .A(data_in[10]), .ZN(n479) );
  INV_X1 U363 ( .A(data_in[11]), .ZN(n478) );
  INV_X1 U364 ( .A(data_in[12]), .ZN(n477) );
  INV_X1 U365 ( .A(data_in[13]), .ZN(n476) );
  INV_X1 U366 ( .A(data_in[14]), .ZN(n475) );
  INV_X1 U367 ( .A(data_in[15]), .ZN(n474) );
  INV_X1 U368 ( .A(data_in[16]), .ZN(n473) );
  INV_X1 U369 ( .A(data_in[17]), .ZN(n472) );
  INV_X1 U370 ( .A(data_in[18]), .ZN(n471) );
  INV_X1 U371 ( .A(data_in[19]), .ZN(n470) );
  MUX2_X1 U372 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n456), .Z(n1) );
  MUX2_X1 U373 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n454), .Z(n2) );
  MUX2_X1 U374 ( .A(n2), .B(n1), .S(n453), .Z(n3) );
  MUX2_X1 U375 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n455), .Z(n4) );
  MUX2_X1 U376 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n457), .Z(n5) );
  MUX2_X1 U377 ( .A(n5), .B(n4), .S(n453), .Z(n6) );
  MUX2_X1 U378 ( .A(n6), .B(n3), .S(N12), .Z(N32) );
  MUX2_X1 U379 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n456), .Z(n7) );
  MUX2_X1 U380 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n455), .Z(n8) );
  MUX2_X1 U381 ( .A(n8), .B(n7), .S(n453), .Z(n9) );
  MUX2_X1 U382 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n455), .Z(n10) );
  MUX2_X1 U383 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n454), .Z(n11) );
  MUX2_X1 U384 ( .A(n11), .B(n10), .S(n453), .Z(n12) );
  MUX2_X1 U385 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n454), .Z(n13) );
  MUX2_X1 U386 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n454), .Z(n14) );
  MUX2_X1 U387 ( .A(n14), .B(n13), .S(n453), .Z(n15) );
  MUX2_X1 U388 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n456), .Z(n16) );
  MUX2_X1 U389 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n456), .Z(n17) );
  MUX2_X1 U390 ( .A(n17), .B(n16), .S(n453), .Z(n18) );
  MUX2_X1 U391 ( .A(n18), .B(n15), .S(N12), .Z(N30) );
  MUX2_X1 U392 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n456), .Z(n19) );
  MUX2_X1 U393 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n456), .Z(n20) );
  MUX2_X1 U394 ( .A(n20), .B(n19), .S(n453), .Z(n21) );
  MUX2_X1 U395 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n455), .Z(n22) );
  MUX2_X1 U396 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n457), .Z(n23) );
  MUX2_X1 U397 ( .A(n23), .B(n22), .S(n453), .Z(n24) );
  MUX2_X1 U398 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n457), .Z(n356) );
  MUX2_X1 U399 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n457), .Z(n357) );
  MUX2_X1 U400 ( .A(n357), .B(n356), .S(n453), .Z(n358) );
  MUX2_X1 U401 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n455), .Z(n359) );
  MUX2_X1 U402 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n456), .Z(n360) );
  MUX2_X1 U403 ( .A(n360), .B(n359), .S(n453), .Z(n361) );
  MUX2_X1 U404 ( .A(n361), .B(n358), .S(N12), .Z(N28) );
  MUX2_X1 U405 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n454), .Z(n362) );
  MUX2_X1 U406 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n454), .Z(n363) );
  MUX2_X1 U407 ( .A(n363), .B(n362), .S(n453), .Z(n364) );
  MUX2_X1 U408 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n454), .Z(n365) );
  MUX2_X1 U409 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n454), .Z(n366) );
  MUX2_X1 U410 ( .A(n366), .B(n365), .S(n453), .Z(n367) );
  MUX2_X1 U411 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n454), .Z(n368) );
  MUX2_X1 U412 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n454), .Z(n369) );
  MUX2_X1 U413 ( .A(n369), .B(n368), .S(n453), .Z(n370) );
  MUX2_X1 U414 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n454), .Z(n371) );
  MUX2_X1 U415 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n454), .Z(n372) );
  MUX2_X1 U416 ( .A(n372), .B(n371), .S(n453), .Z(n373) );
  MUX2_X1 U417 ( .A(n373), .B(n370), .S(N12), .Z(N26) );
  MUX2_X1 U418 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n454), .Z(n374) );
  MUX2_X1 U419 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n454), .Z(n375) );
  MUX2_X1 U420 ( .A(n375), .B(n374), .S(n453), .Z(n376) );
  MUX2_X1 U421 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n454), .Z(n377) );
  MUX2_X1 U422 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n454), .Z(n378) );
  MUX2_X1 U423 ( .A(n378), .B(n377), .S(n453), .Z(n379) );
  MUX2_X1 U424 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n455), .Z(n380) );
  MUX2_X1 U425 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n455), .Z(n381) );
  MUX2_X1 U426 ( .A(n381), .B(n380), .S(n452), .Z(n382) );
  MUX2_X1 U427 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n455), .Z(n383) );
  MUX2_X1 U428 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n455), .Z(n384) );
  MUX2_X1 U429 ( .A(n384), .B(n383), .S(n452), .Z(n385) );
  MUX2_X1 U430 ( .A(n385), .B(n382), .S(N12), .Z(N24) );
  MUX2_X1 U431 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n455), .Z(n386) );
  MUX2_X1 U432 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n455), .Z(n387) );
  MUX2_X1 U433 ( .A(n387), .B(n386), .S(n452), .Z(n388) );
  MUX2_X1 U434 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n455), .Z(n389) );
  MUX2_X1 U435 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n455), .Z(n390) );
  MUX2_X1 U436 ( .A(n390), .B(n389), .S(n452), .Z(n391) );
  MUX2_X1 U437 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n455), .Z(n392) );
  MUX2_X1 U438 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n455), .Z(n393) );
  MUX2_X1 U439 ( .A(n393), .B(n392), .S(n452), .Z(n394) );
  MUX2_X1 U440 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n455), .Z(n395) );
  MUX2_X1 U441 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n455), .Z(n396) );
  MUX2_X1 U442 ( .A(n396), .B(n395), .S(n452), .Z(n397) );
  MUX2_X1 U443 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n456), .Z(n398) );
  MUX2_X1 U444 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n456), .Z(n399) );
  MUX2_X1 U445 ( .A(n399), .B(n398), .S(n452), .Z(n400) );
  MUX2_X1 U446 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n456), .Z(n401) );
  MUX2_X1 U447 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n456), .Z(n402) );
  MUX2_X1 U448 ( .A(n402), .B(n401), .S(n452), .Z(n403) );
  MUX2_X1 U449 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n456), .Z(n404) );
  MUX2_X1 U450 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n456), .Z(n405) );
  MUX2_X1 U451 ( .A(n405), .B(n404), .S(n452), .Z(n406) );
  MUX2_X1 U452 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n456), .Z(n407) );
  MUX2_X1 U453 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n456), .Z(n408) );
  MUX2_X1 U454 ( .A(n408), .B(n407), .S(n452), .Z(n409) );
  MUX2_X1 U455 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n456), .Z(n410) );
  MUX2_X1 U456 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n456), .Z(n411) );
  MUX2_X1 U457 ( .A(n411), .B(n410), .S(n452), .Z(n412) );
  MUX2_X1 U458 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n456), .Z(n413) );
  MUX2_X1 U459 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n456), .Z(n414) );
  MUX2_X1 U460 ( .A(n414), .B(n413), .S(n452), .Z(n415) );
  MUX2_X1 U461 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n457), .Z(n416) );
  MUX2_X1 U462 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n457), .Z(n417) );
  MUX2_X1 U463 ( .A(n417), .B(n416), .S(n453), .Z(n418) );
  MUX2_X1 U464 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n457), .Z(n419) );
  MUX2_X1 U465 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n457), .Z(n420) );
  MUX2_X1 U466 ( .A(n420), .B(n419), .S(n453), .Z(n421) );
  MUX2_X1 U467 ( .A(n421), .B(n418), .S(N12), .Z(N18) );
  MUX2_X1 U468 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n457), .Z(n422) );
  MUX2_X1 U469 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n457), .Z(n423) );
  MUX2_X1 U470 ( .A(n423), .B(n422), .S(N11), .Z(n424) );
  MUX2_X1 U471 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n457), .Z(n425) );
  MUX2_X1 U472 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n457), .Z(n426) );
  MUX2_X1 U473 ( .A(n426), .B(n425), .S(N11), .Z(n427) );
  MUX2_X1 U474 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n457), .Z(n428) );
  MUX2_X1 U475 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n457), .Z(n429) );
  MUX2_X1 U476 ( .A(n429), .B(n428), .S(n453), .Z(n430) );
  MUX2_X1 U477 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n457), .Z(n431) );
  MUX2_X1 U478 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n457), .Z(n432) );
  MUX2_X1 U479 ( .A(n432), .B(n431), .S(N11), .Z(n433) );
  MUX2_X1 U480 ( .A(n433), .B(n430), .S(N12), .Z(N16) );
  MUX2_X1 U481 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n454), .Z(n434) );
  MUX2_X1 U482 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n454), .Z(n435) );
  MUX2_X1 U483 ( .A(n435), .B(n434), .S(n453), .Z(n436) );
  MUX2_X1 U484 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n454), .Z(n437) );
  MUX2_X1 U485 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n456), .Z(n438) );
  MUX2_X1 U486 ( .A(n438), .B(n437), .S(N11), .Z(n439) );
  MUX2_X1 U487 ( .A(n439), .B(n436), .S(N12), .Z(N15) );
  MUX2_X1 U488 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n457), .Z(n440) );
  MUX2_X1 U489 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n457), .Z(n441) );
  MUX2_X1 U490 ( .A(n441), .B(n440), .S(n453), .Z(n442) );
  MUX2_X1 U491 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n457), .Z(n443) );
  MUX2_X1 U492 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n454), .Z(n444) );
  MUX2_X1 U493 ( .A(n444), .B(n443), .S(N11), .Z(n445) );
  MUX2_X1 U494 ( .A(n445), .B(n442), .S(N12), .Z(N14) );
  MUX2_X1 U495 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n455), .Z(n446) );
  MUX2_X1 U496 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n455), .Z(n447) );
  MUX2_X1 U497 ( .A(n447), .B(n446), .S(n453), .Z(n448) );
  MUX2_X1 U498 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n455), .Z(n449) );
  MUX2_X1 U499 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n457), .Z(n450) );
  MUX2_X1 U500 ( .A(n450), .B(n449), .S(N11), .Z(n451) );
  MUX2_X1 U501 ( .A(n451), .B(n448), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE4_0 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N22, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n491), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n492), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n493), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n494), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n495), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n496), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n497), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n498), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n499), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n500), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n501), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n502), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n503), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n504), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n505), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n506), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n507), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n508), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n509), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n510), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n511), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n512), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n513), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n514), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n515), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n516), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n517), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n518), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n519), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n520), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n521), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n522), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n523), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n524), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n525), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n526), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n527), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n528), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n529), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n530), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n531), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n532), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n533), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n534), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n535), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n536), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n537), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n538), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n539), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n540), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n541), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n542), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n543), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n544), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n545), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n546), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n547), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n548), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n549), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n550), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n551), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n552), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n553), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n554), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n555), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n556), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n557), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n558), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n559), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n560), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n561), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n562), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n563), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n564), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n565), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n566), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n567), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n568), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n569), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n570), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n571), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n572), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n573), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n574), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n575), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n576), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n577), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n578), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n579), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n580), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n581), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n582), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n583), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n584), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n585), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n586), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n587), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n588), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n589), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n590), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n591), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n592), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n593), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n594), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n595), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n596), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n597), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n598), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n599), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n600), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n601), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n602), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n603), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n604), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n605), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n606), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n607), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n608), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n609), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n610), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n611), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n612), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n613), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n614), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n615), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n616), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n617), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n618), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n619), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n620), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n621), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n622), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n623), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n624), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n625), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n626), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n627), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n628), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n629), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n630), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n631), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n632), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n633), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n634), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n635), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n636), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n637), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n638), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n639), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n640), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n641), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n642), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n643), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n644), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n645), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n646), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n647), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n648), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n649), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n650), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U350 ( .A1(n467), .A2(n468), .A3(n800), .ZN(n821) );
  NAND3_X1 U351 ( .A1(n800), .A2(n468), .A3(N10), .ZN(n799) );
  NAND3_X1 U352 ( .A1(n800), .A2(n467), .A3(N11), .ZN(n778) );
  NAND3_X1 U353 ( .A1(N10), .A2(n800), .A3(N11), .ZN(n757) );
  NAND3_X1 U354 ( .A1(n467), .A2(n468), .A3(n714), .ZN(n735) );
  NAND3_X1 U355 ( .A1(N10), .A2(n468), .A3(n714), .ZN(n713) );
  NAND3_X1 U356 ( .A1(N11), .A2(n467), .A3(n714), .ZN(n692) );
  NAND3_X1 U357 ( .A1(N11), .A2(N10), .A3(n714), .ZN(n671) );
  SDFF_X1 \data_out_reg[19]  ( .D(n449), .SI(n452), .SE(n469), .CK(clk), .Q(
        data_out[19]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n389), .SI(n392), .SE(n469), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n4), .SI(n7), .SE(n469), .CK(clk), .Q(
        data_out[0]) );
  SDFF_X1 \data_out_reg[16]  ( .D(n431), .SI(n434), .SE(n469), .CK(clk), .Q(
        data_out[16]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n383), .SI(n386), .SE(n469), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[14]  ( .D(n419), .SI(n422), .SE(n469), .CK(clk), .Q(
        data_out[14]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n401), .SI(n404), .SE(n469), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n22), .SI(n356), .SE(n469), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n377), .SI(n380), .SE(n469), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n365), .SI(n368), .SE(n469), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[18]  ( .D(n443), .SI(n446), .SE(n469), .CK(clk), .Q(
        data_out[18]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n16), .SI(n19), .SE(n469), .CK(clk), .Q(
        data_out[2]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n10), .SI(n13), .SE(n469), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[12]  ( .D(n407), .SI(n410), .SE(n469), .CK(clk), .Q(
        data_out[12]) );
  SDFF_X1 \data_out_reg[4]  ( .D(n359), .SI(n362), .SE(n469), .CK(clk), .Q(
        data_out[4]) );
  SDFF_X1 \data_out_reg[17]  ( .D(n437), .SI(n440), .SE(n469), .CK(clk), .Q(
        data_out[17]) );
  SDFF_X1 \data_out_reg[6]  ( .D(n371), .SI(n374), .SE(n469), .CK(clk), .Q(
        data_out[6]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n425), .SI(n428), .SE(n469), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n413), .SI(n416), .SE(n469), .CK(clk), .Q(
        data_out[13]) );
  BUF_X1 U3 ( .A(n713), .Z(n461) );
  BUF_X1 U4 ( .A(n821), .Z(n466) );
  BUF_X1 U5 ( .A(n778), .Z(n464) );
  BUF_X1 U6 ( .A(n454), .Z(n453) );
  BUF_X1 U7 ( .A(N10), .Z(n457) );
  BUF_X1 U8 ( .A(N10), .Z(n458) );
  BUF_X1 U9 ( .A(N10), .Z(n456) );
  BUF_X1 U10 ( .A(n757), .Z(n463) );
  BUF_X1 U11 ( .A(n799), .Z(n465) );
  BUF_X1 U12 ( .A(n671), .Z(n459) );
  BUF_X1 U13 ( .A(n692), .Z(n460) );
  BUF_X1 U14 ( .A(N11), .Z(n454) );
  BUF_X1 U15 ( .A(n735), .Z(n462) );
  NOR2_X1 U16 ( .A1(n736), .A2(N12), .ZN(n800) );
  NOR2_X1 U17 ( .A1(n469), .A2(n736), .ZN(n714) );
  INV_X1 U18 ( .A(N12), .ZN(n469) );
  INV_X1 U19 ( .A(N11), .ZN(n468) );
  INV_X1 U20 ( .A(N10), .ZN(n467) );
  NAND2_X1 U21 ( .A1(wr_en), .A2(n470), .ZN(n736) );
  INV_X1 U22 ( .A(addr[3]), .ZN(n470) );
  OAI21_X1 U23 ( .B1(n478), .B2(n799), .A(n786), .ZN(n618) );
  NAND2_X1 U24 ( .A1(\mem[1][12] ), .A2(n799), .ZN(n786) );
  OAI21_X1 U25 ( .B1(n477), .B2(n799), .A(n785), .ZN(n617) );
  NAND2_X1 U26 ( .A1(\mem[1][13] ), .A2(n799), .ZN(n785) );
  OAI21_X1 U27 ( .B1(n476), .B2(n799), .A(n784), .ZN(n616) );
  NAND2_X1 U28 ( .A1(\mem[1][14] ), .A2(n799), .ZN(n784) );
  OAI21_X1 U29 ( .B1(n475), .B2(n465), .A(n783), .ZN(n615) );
  NAND2_X1 U30 ( .A1(\mem[1][15] ), .A2(n799), .ZN(n783) );
  OAI21_X1 U31 ( .B1(n474), .B2(n799), .A(n782), .ZN(n614) );
  NAND2_X1 U32 ( .A1(\mem[1][16] ), .A2(n465), .ZN(n782) );
  OAI21_X1 U33 ( .B1(n473), .B2(n799), .A(n781), .ZN(n613) );
  NAND2_X1 U34 ( .A1(\mem[1][17] ), .A2(n799), .ZN(n781) );
  OAI21_X1 U35 ( .B1(n472), .B2(n799), .A(n780), .ZN(n612) );
  NAND2_X1 U36 ( .A1(\mem[1][18] ), .A2(n799), .ZN(n780) );
  OAI21_X1 U37 ( .B1(n471), .B2(n799), .A(n779), .ZN(n611) );
  NAND2_X1 U38 ( .A1(\mem[1][19] ), .A2(n465), .ZN(n779) );
  OAI21_X1 U39 ( .B1(n478), .B2(n778), .A(n765), .ZN(n598) );
  NAND2_X1 U40 ( .A1(\mem[2][12] ), .A2(n778), .ZN(n765) );
  OAI21_X1 U41 ( .B1(n477), .B2(n778), .A(n764), .ZN(n597) );
  NAND2_X1 U42 ( .A1(\mem[2][13] ), .A2(n778), .ZN(n764) );
  OAI21_X1 U43 ( .B1(n476), .B2(n464), .A(n763), .ZN(n596) );
  NAND2_X1 U44 ( .A1(\mem[2][14] ), .A2(n778), .ZN(n763) );
  OAI21_X1 U45 ( .B1(n475), .B2(n464), .A(n762), .ZN(n595) );
  NAND2_X1 U46 ( .A1(\mem[2][15] ), .A2(n778), .ZN(n762) );
  OAI21_X1 U47 ( .B1(n474), .B2(n464), .A(n761), .ZN(n594) );
  NAND2_X1 U48 ( .A1(\mem[2][16] ), .A2(n778), .ZN(n761) );
  OAI21_X1 U49 ( .B1(n473), .B2(n464), .A(n760), .ZN(n593) );
  NAND2_X1 U50 ( .A1(\mem[2][17] ), .A2(n778), .ZN(n760) );
  OAI21_X1 U51 ( .B1(n472), .B2(n464), .A(n759), .ZN(n592) );
  NAND2_X1 U52 ( .A1(\mem[2][18] ), .A2(n778), .ZN(n759) );
  OAI21_X1 U53 ( .B1(n471), .B2(n778), .A(n758), .ZN(n591) );
  NAND2_X1 U54 ( .A1(\mem[2][19] ), .A2(n778), .ZN(n758) );
  OAI21_X1 U55 ( .B1(n478), .B2(n757), .A(n744), .ZN(n578) );
  NAND2_X1 U56 ( .A1(\mem[3][12] ), .A2(n757), .ZN(n744) );
  OAI21_X1 U57 ( .B1(n477), .B2(n757), .A(n743), .ZN(n577) );
  NAND2_X1 U58 ( .A1(\mem[3][13] ), .A2(n757), .ZN(n743) );
  OAI21_X1 U59 ( .B1(n476), .B2(n757), .A(n742), .ZN(n576) );
  NAND2_X1 U60 ( .A1(\mem[3][14] ), .A2(n757), .ZN(n742) );
  OAI21_X1 U61 ( .B1(n475), .B2(n757), .A(n741), .ZN(n575) );
  NAND2_X1 U62 ( .A1(\mem[3][15] ), .A2(n463), .ZN(n741) );
  OAI21_X1 U63 ( .B1(n474), .B2(n463), .A(n740), .ZN(n574) );
  NAND2_X1 U64 ( .A1(\mem[3][16] ), .A2(n757), .ZN(n740) );
  OAI21_X1 U65 ( .B1(n473), .B2(n463), .A(n739), .ZN(n573) );
  NAND2_X1 U66 ( .A1(\mem[3][17] ), .A2(n757), .ZN(n739) );
  OAI21_X1 U67 ( .B1(n472), .B2(n463), .A(n738), .ZN(n572) );
  NAND2_X1 U68 ( .A1(\mem[3][18] ), .A2(n757), .ZN(n738) );
  OAI21_X1 U69 ( .B1(n471), .B2(n757), .A(n737), .ZN(n571) );
  NAND2_X1 U70 ( .A1(\mem[3][19] ), .A2(n463), .ZN(n737) );
  OAI21_X1 U71 ( .B1(n490), .B2(n462), .A(n734), .ZN(n570) );
  NAND2_X1 U72 ( .A1(\mem[4][0] ), .A2(n735), .ZN(n734) );
  OAI21_X1 U73 ( .B1(n489), .B2(n735), .A(n733), .ZN(n569) );
  NAND2_X1 U74 ( .A1(\mem[4][1] ), .A2(n735), .ZN(n733) );
  OAI21_X1 U75 ( .B1(n488), .B2(n735), .A(n732), .ZN(n568) );
  NAND2_X1 U76 ( .A1(\mem[4][2] ), .A2(n735), .ZN(n732) );
  OAI21_X1 U77 ( .B1(n487), .B2(n735), .A(n731), .ZN(n567) );
  NAND2_X1 U78 ( .A1(\mem[4][3] ), .A2(n735), .ZN(n731) );
  OAI21_X1 U79 ( .B1(n486), .B2(n735), .A(n730), .ZN(n566) );
  NAND2_X1 U80 ( .A1(\mem[4][4] ), .A2(n735), .ZN(n730) );
  OAI21_X1 U81 ( .B1(n485), .B2(n735), .A(n729), .ZN(n565) );
  NAND2_X1 U82 ( .A1(\mem[4][5] ), .A2(n735), .ZN(n729) );
  OAI21_X1 U83 ( .B1(n484), .B2(n735), .A(n728), .ZN(n564) );
  NAND2_X1 U84 ( .A1(\mem[4][6] ), .A2(n735), .ZN(n728) );
  OAI21_X1 U85 ( .B1(n483), .B2(n462), .A(n727), .ZN(n563) );
  NAND2_X1 U86 ( .A1(\mem[4][7] ), .A2(n735), .ZN(n727) );
  OAI21_X1 U87 ( .B1(n482), .B2(n462), .A(n726), .ZN(n562) );
  NAND2_X1 U88 ( .A1(\mem[4][8] ), .A2(n735), .ZN(n726) );
  OAI21_X1 U89 ( .B1(n481), .B2(n735), .A(n725), .ZN(n561) );
  NAND2_X1 U90 ( .A1(\mem[4][9] ), .A2(n735), .ZN(n725) );
  OAI21_X1 U91 ( .B1(n480), .B2(n462), .A(n724), .ZN(n560) );
  NAND2_X1 U92 ( .A1(\mem[4][10] ), .A2(n735), .ZN(n724) );
  OAI21_X1 U93 ( .B1(n479), .B2(n462), .A(n723), .ZN(n559) );
  NAND2_X1 U94 ( .A1(\mem[4][11] ), .A2(n735), .ZN(n723) );
  OAI21_X1 U95 ( .B1(n478), .B2(n735), .A(n722), .ZN(n558) );
  NAND2_X1 U96 ( .A1(\mem[4][12] ), .A2(n462), .ZN(n722) );
  OAI21_X1 U97 ( .B1(n477), .B2(n735), .A(n721), .ZN(n557) );
  NAND2_X1 U98 ( .A1(\mem[4][13] ), .A2(n462), .ZN(n721) );
  OAI21_X1 U99 ( .B1(n476), .B2(n462), .A(n720), .ZN(n556) );
  NAND2_X1 U100 ( .A1(\mem[4][14] ), .A2(n462), .ZN(n720) );
  OAI21_X1 U101 ( .B1(n475), .B2(n462), .A(n719), .ZN(n555) );
  NAND2_X1 U102 ( .A1(\mem[4][15] ), .A2(n462), .ZN(n719) );
  OAI21_X1 U103 ( .B1(n474), .B2(n462), .A(n718), .ZN(n554) );
  NAND2_X1 U104 ( .A1(\mem[4][16] ), .A2(n462), .ZN(n718) );
  OAI21_X1 U105 ( .B1(n473), .B2(n462), .A(n717), .ZN(n553) );
  NAND2_X1 U106 ( .A1(\mem[4][17] ), .A2(n462), .ZN(n717) );
  OAI21_X1 U107 ( .B1(n472), .B2(n735), .A(n716), .ZN(n552) );
  NAND2_X1 U108 ( .A1(\mem[4][18] ), .A2(n462), .ZN(n716) );
  OAI21_X1 U109 ( .B1(n471), .B2(n735), .A(n715), .ZN(n551) );
  NAND2_X1 U110 ( .A1(\mem[4][19] ), .A2(n735), .ZN(n715) );
  OAI21_X1 U111 ( .B1(n490), .B2(n461), .A(n712), .ZN(n550) );
  NAND2_X1 U112 ( .A1(\mem[5][0] ), .A2(n713), .ZN(n712) );
  OAI21_X1 U113 ( .B1(n489), .B2(n461), .A(n711), .ZN(n549) );
  NAND2_X1 U114 ( .A1(\mem[5][1] ), .A2(n713), .ZN(n711) );
  OAI21_X1 U115 ( .B1(n488), .B2(n461), .A(n710), .ZN(n548) );
  NAND2_X1 U116 ( .A1(\mem[5][2] ), .A2(n713), .ZN(n710) );
  OAI21_X1 U117 ( .B1(n487), .B2(n713), .A(n709), .ZN(n547) );
  NAND2_X1 U118 ( .A1(\mem[5][3] ), .A2(n713), .ZN(n709) );
  OAI21_X1 U119 ( .B1(n486), .B2(n713), .A(n708), .ZN(n546) );
  NAND2_X1 U120 ( .A1(\mem[5][4] ), .A2(n713), .ZN(n708) );
  OAI21_X1 U121 ( .B1(n485), .B2(n713), .A(n707), .ZN(n545) );
  NAND2_X1 U122 ( .A1(\mem[5][5] ), .A2(n713), .ZN(n707) );
  OAI21_X1 U123 ( .B1(n484), .B2(n713), .A(n706), .ZN(n544) );
  NAND2_X1 U124 ( .A1(\mem[5][6] ), .A2(n461), .ZN(n706) );
  OAI21_X1 U125 ( .B1(n483), .B2(n713), .A(n705), .ZN(n543) );
  NAND2_X1 U126 ( .A1(\mem[5][7] ), .A2(n461), .ZN(n705) );
  OAI21_X1 U127 ( .B1(n482), .B2(n713), .A(n704), .ZN(n542) );
  NAND2_X1 U128 ( .A1(\mem[5][8] ), .A2(n713), .ZN(n704) );
  OAI21_X1 U129 ( .B1(n481), .B2(n461), .A(n703), .ZN(n541) );
  NAND2_X1 U130 ( .A1(\mem[5][9] ), .A2(n461), .ZN(n703) );
  OAI21_X1 U131 ( .B1(n480), .B2(n713), .A(n702), .ZN(n540) );
  NAND2_X1 U132 ( .A1(\mem[5][10] ), .A2(n713), .ZN(n702) );
  OAI21_X1 U133 ( .B1(n479), .B2(n713), .A(n701), .ZN(n539) );
  NAND2_X1 U134 ( .A1(\mem[5][11] ), .A2(n713), .ZN(n701) );
  OAI21_X1 U135 ( .B1(n478), .B2(n461), .A(n700), .ZN(n538) );
  NAND2_X1 U136 ( .A1(\mem[5][12] ), .A2(n461), .ZN(n700) );
  OAI21_X1 U137 ( .B1(n477), .B2(n461), .A(n699), .ZN(n537) );
  NAND2_X1 U138 ( .A1(\mem[5][13] ), .A2(n461), .ZN(n699) );
  OAI21_X1 U139 ( .B1(n476), .B2(n461), .A(n698), .ZN(n536) );
  NAND2_X1 U140 ( .A1(\mem[5][14] ), .A2(n461), .ZN(n698) );
  OAI21_X1 U141 ( .B1(n475), .B2(n713), .A(n697), .ZN(n535) );
  NAND2_X1 U142 ( .A1(\mem[5][15] ), .A2(n461), .ZN(n697) );
  OAI21_X1 U143 ( .B1(n474), .B2(n713), .A(n696), .ZN(n534) );
  NAND2_X1 U144 ( .A1(\mem[5][16] ), .A2(n461), .ZN(n696) );
  OAI21_X1 U145 ( .B1(n473), .B2(n713), .A(n695), .ZN(n533) );
  NAND2_X1 U146 ( .A1(\mem[5][17] ), .A2(n461), .ZN(n695) );
  OAI21_X1 U147 ( .B1(n472), .B2(n713), .A(n694), .ZN(n532) );
  NAND2_X1 U148 ( .A1(\mem[5][18] ), .A2(n461), .ZN(n694) );
  OAI21_X1 U149 ( .B1(n471), .B2(n461), .A(n693), .ZN(n531) );
  NAND2_X1 U150 ( .A1(\mem[5][19] ), .A2(n461), .ZN(n693) );
  OAI21_X1 U151 ( .B1(n490), .B2(n692), .A(n691), .ZN(n530) );
  NAND2_X1 U152 ( .A1(\mem[6][0] ), .A2(n460), .ZN(n691) );
  OAI21_X1 U153 ( .B1(n489), .B2(n692), .A(n690), .ZN(n529) );
  NAND2_X1 U154 ( .A1(\mem[6][1] ), .A2(n460), .ZN(n690) );
  OAI21_X1 U155 ( .B1(n488), .B2(n692), .A(n689), .ZN(n528) );
  NAND2_X1 U156 ( .A1(\mem[6][2] ), .A2(n460), .ZN(n689) );
  OAI21_X1 U157 ( .B1(n487), .B2(n692), .A(n688), .ZN(n527) );
  NAND2_X1 U158 ( .A1(\mem[6][3] ), .A2(n460), .ZN(n688) );
  OAI21_X1 U159 ( .B1(n486), .B2(n460), .A(n687), .ZN(n526) );
  NAND2_X1 U160 ( .A1(\mem[6][4] ), .A2(n460), .ZN(n687) );
  OAI21_X1 U161 ( .B1(n485), .B2(n692), .A(n686), .ZN(n525) );
  NAND2_X1 U162 ( .A1(\mem[6][5] ), .A2(n460), .ZN(n686) );
  OAI21_X1 U163 ( .B1(n484), .B2(n692), .A(n685), .ZN(n524) );
  NAND2_X1 U164 ( .A1(\mem[6][6] ), .A2(n460), .ZN(n685) );
  OAI21_X1 U165 ( .B1(n483), .B2(n692), .A(n684), .ZN(n523) );
  NAND2_X1 U166 ( .A1(\mem[6][7] ), .A2(n460), .ZN(n684) );
  OAI21_X1 U167 ( .B1(n482), .B2(n692), .A(n683), .ZN(n522) );
  NAND2_X1 U168 ( .A1(\mem[6][8] ), .A2(n460), .ZN(n683) );
  OAI21_X1 U169 ( .B1(n481), .B2(n692), .A(n682), .ZN(n521) );
  NAND2_X1 U170 ( .A1(\mem[6][9] ), .A2(n460), .ZN(n682) );
  OAI21_X1 U171 ( .B1(n480), .B2(n692), .A(n681), .ZN(n520) );
  NAND2_X1 U172 ( .A1(\mem[6][10] ), .A2(n460), .ZN(n681) );
  OAI21_X1 U173 ( .B1(n479), .B2(n692), .A(n680), .ZN(n519) );
  NAND2_X1 U174 ( .A1(\mem[6][11] ), .A2(n460), .ZN(n680) );
  OAI21_X1 U175 ( .B1(n478), .B2(n692), .A(n679), .ZN(n518) );
  NAND2_X1 U176 ( .A1(\mem[6][12] ), .A2(n692), .ZN(n679) );
  OAI21_X1 U177 ( .B1(n477), .B2(n460), .A(n678), .ZN(n517) );
  NAND2_X1 U178 ( .A1(\mem[6][13] ), .A2(n692), .ZN(n678) );
  OAI21_X1 U179 ( .B1(n476), .B2(n460), .A(n677), .ZN(n516) );
  NAND2_X1 U180 ( .A1(\mem[6][14] ), .A2(n692), .ZN(n677) );
  OAI21_X1 U181 ( .B1(n475), .B2(n692), .A(n676), .ZN(n515) );
  NAND2_X1 U182 ( .A1(\mem[6][15] ), .A2(n692), .ZN(n676) );
  OAI21_X1 U183 ( .B1(n474), .B2(n692), .A(n675), .ZN(n514) );
  NAND2_X1 U184 ( .A1(\mem[6][16] ), .A2(n692), .ZN(n675) );
  OAI21_X1 U185 ( .B1(n473), .B2(n692), .A(n674), .ZN(n513) );
  NAND2_X1 U186 ( .A1(\mem[6][17] ), .A2(n692), .ZN(n674) );
  OAI21_X1 U187 ( .B1(n472), .B2(n692), .A(n673), .ZN(n512) );
  NAND2_X1 U188 ( .A1(\mem[6][18] ), .A2(n692), .ZN(n673) );
  OAI21_X1 U189 ( .B1(n471), .B2(n692), .A(n672), .ZN(n511) );
  NAND2_X1 U190 ( .A1(\mem[6][19] ), .A2(n460), .ZN(n672) );
  OAI21_X1 U191 ( .B1(n490), .B2(n671), .A(n670), .ZN(n510) );
  NAND2_X1 U192 ( .A1(\mem[7][0] ), .A2(n459), .ZN(n670) );
  OAI21_X1 U193 ( .B1(n489), .B2(n671), .A(n669), .ZN(n509) );
  NAND2_X1 U194 ( .A1(\mem[7][1] ), .A2(n459), .ZN(n669) );
  OAI21_X1 U195 ( .B1(n488), .B2(n671), .A(n668), .ZN(n508) );
  NAND2_X1 U196 ( .A1(\mem[7][2] ), .A2(n459), .ZN(n668) );
  OAI21_X1 U197 ( .B1(n487), .B2(n671), .A(n667), .ZN(n507) );
  NAND2_X1 U198 ( .A1(\mem[7][3] ), .A2(n459), .ZN(n667) );
  OAI21_X1 U199 ( .B1(n486), .B2(n459), .A(n666), .ZN(n506) );
  NAND2_X1 U200 ( .A1(\mem[7][4] ), .A2(n459), .ZN(n666) );
  OAI21_X1 U201 ( .B1(n485), .B2(n671), .A(n665), .ZN(n505) );
  NAND2_X1 U202 ( .A1(\mem[7][5] ), .A2(n459), .ZN(n665) );
  OAI21_X1 U203 ( .B1(n484), .B2(n671), .A(n664), .ZN(n504) );
  NAND2_X1 U204 ( .A1(\mem[7][6] ), .A2(n459), .ZN(n664) );
  OAI21_X1 U205 ( .B1(n483), .B2(n671), .A(n663), .ZN(n503) );
  NAND2_X1 U206 ( .A1(\mem[7][7] ), .A2(n459), .ZN(n663) );
  OAI21_X1 U207 ( .B1(n482), .B2(n671), .A(n662), .ZN(n502) );
  NAND2_X1 U208 ( .A1(\mem[7][8] ), .A2(n459), .ZN(n662) );
  OAI21_X1 U209 ( .B1(n481), .B2(n671), .A(n661), .ZN(n501) );
  NAND2_X1 U210 ( .A1(\mem[7][9] ), .A2(n459), .ZN(n661) );
  OAI21_X1 U211 ( .B1(n480), .B2(n671), .A(n660), .ZN(n500) );
  NAND2_X1 U212 ( .A1(\mem[7][10] ), .A2(n459), .ZN(n660) );
  OAI21_X1 U213 ( .B1(n479), .B2(n671), .A(n659), .ZN(n499) );
  NAND2_X1 U214 ( .A1(\mem[7][11] ), .A2(n459), .ZN(n659) );
  OAI21_X1 U215 ( .B1(n478), .B2(n671), .A(n658), .ZN(n498) );
  NAND2_X1 U216 ( .A1(\mem[7][12] ), .A2(n671), .ZN(n658) );
  OAI21_X1 U217 ( .B1(n477), .B2(n459), .A(n657), .ZN(n497) );
  NAND2_X1 U218 ( .A1(\mem[7][13] ), .A2(n671), .ZN(n657) );
  OAI21_X1 U219 ( .B1(n476), .B2(n459), .A(n656), .ZN(n496) );
  NAND2_X1 U220 ( .A1(\mem[7][14] ), .A2(n671), .ZN(n656) );
  OAI21_X1 U221 ( .B1(n475), .B2(n671), .A(n655), .ZN(n495) );
  NAND2_X1 U222 ( .A1(\mem[7][15] ), .A2(n671), .ZN(n655) );
  OAI21_X1 U223 ( .B1(n474), .B2(n671), .A(n654), .ZN(n494) );
  NAND2_X1 U224 ( .A1(\mem[7][16] ), .A2(n671), .ZN(n654) );
  OAI21_X1 U225 ( .B1(n473), .B2(n671), .A(n653), .ZN(n493) );
  NAND2_X1 U226 ( .A1(\mem[7][17] ), .A2(n671), .ZN(n653) );
  OAI21_X1 U227 ( .B1(n472), .B2(n671), .A(n652), .ZN(n492) );
  NAND2_X1 U228 ( .A1(\mem[7][18] ), .A2(n671), .ZN(n652) );
  OAI21_X1 U229 ( .B1(n471), .B2(n671), .A(n651), .ZN(n491) );
  NAND2_X1 U230 ( .A1(\mem[7][19] ), .A2(n459), .ZN(n651) );
  OAI21_X1 U231 ( .B1(n821), .B2(n490), .A(n820), .ZN(n650) );
  NAND2_X1 U232 ( .A1(\mem[0][0] ), .A2(n821), .ZN(n820) );
  OAI21_X1 U233 ( .B1(n821), .B2(n489), .A(n819), .ZN(n649) );
  NAND2_X1 U234 ( .A1(\mem[0][1] ), .A2(n821), .ZN(n819) );
  OAI21_X1 U235 ( .B1(n821), .B2(n488), .A(n818), .ZN(n648) );
  NAND2_X1 U236 ( .A1(\mem[0][2] ), .A2(n466), .ZN(n818) );
  OAI21_X1 U237 ( .B1(n821), .B2(n487), .A(n817), .ZN(n647) );
  NAND2_X1 U238 ( .A1(\mem[0][3] ), .A2(n466), .ZN(n817) );
  OAI21_X1 U239 ( .B1(n821), .B2(n486), .A(n816), .ZN(n646) );
  NAND2_X1 U240 ( .A1(\mem[0][4] ), .A2(n466), .ZN(n816) );
  OAI21_X1 U241 ( .B1(n821), .B2(n485), .A(n815), .ZN(n645) );
  NAND2_X1 U242 ( .A1(\mem[0][5] ), .A2(n466), .ZN(n815) );
  OAI21_X1 U243 ( .B1(n821), .B2(n484), .A(n814), .ZN(n644) );
  NAND2_X1 U244 ( .A1(\mem[0][6] ), .A2(n466), .ZN(n814) );
  OAI21_X1 U245 ( .B1(n821), .B2(n483), .A(n813), .ZN(n643) );
  NAND2_X1 U246 ( .A1(\mem[0][7] ), .A2(n821), .ZN(n813) );
  OAI21_X1 U247 ( .B1(n821), .B2(n482), .A(n812), .ZN(n642) );
  NAND2_X1 U248 ( .A1(\mem[0][8] ), .A2(n821), .ZN(n812) );
  OAI21_X1 U249 ( .B1(n466), .B2(n481), .A(n811), .ZN(n641) );
  NAND2_X1 U250 ( .A1(\mem[0][9] ), .A2(n821), .ZN(n811) );
  OAI21_X1 U251 ( .B1(n821), .B2(n480), .A(n810), .ZN(n640) );
  NAND2_X1 U252 ( .A1(\mem[0][10] ), .A2(n821), .ZN(n810) );
  OAI21_X1 U253 ( .B1(n821), .B2(n479), .A(n809), .ZN(n639) );
  NAND2_X1 U254 ( .A1(\mem[0][11] ), .A2(n821), .ZN(n809) );
  OAI21_X1 U255 ( .B1(n490), .B2(n799), .A(n798), .ZN(n630) );
  NAND2_X1 U256 ( .A1(\mem[1][0] ), .A2(n465), .ZN(n798) );
  OAI21_X1 U257 ( .B1(n489), .B2(n799), .A(n797), .ZN(n629) );
  NAND2_X1 U258 ( .A1(\mem[1][1] ), .A2(n465), .ZN(n797) );
  OAI21_X1 U259 ( .B1(n488), .B2(n799), .A(n796), .ZN(n628) );
  NAND2_X1 U260 ( .A1(\mem[1][2] ), .A2(n465), .ZN(n796) );
  OAI21_X1 U261 ( .B1(n487), .B2(n799), .A(n795), .ZN(n627) );
  NAND2_X1 U262 ( .A1(\mem[1][3] ), .A2(n465), .ZN(n795) );
  OAI21_X1 U263 ( .B1(n486), .B2(n799), .A(n794), .ZN(n626) );
  NAND2_X1 U264 ( .A1(\mem[1][4] ), .A2(n465), .ZN(n794) );
  OAI21_X1 U265 ( .B1(n485), .B2(n799), .A(n793), .ZN(n625) );
  NAND2_X1 U266 ( .A1(\mem[1][5] ), .A2(n465), .ZN(n793) );
  OAI21_X1 U267 ( .B1(n484), .B2(n799), .A(n792), .ZN(n624) );
  NAND2_X1 U268 ( .A1(\mem[1][6] ), .A2(n465), .ZN(n792) );
  OAI21_X1 U269 ( .B1(n483), .B2(n799), .A(n791), .ZN(n623) );
  NAND2_X1 U270 ( .A1(\mem[1][7] ), .A2(n465), .ZN(n791) );
  OAI21_X1 U271 ( .B1(n482), .B2(n799), .A(n790), .ZN(n622) );
  NAND2_X1 U272 ( .A1(\mem[1][8] ), .A2(n465), .ZN(n790) );
  OAI21_X1 U273 ( .B1(n481), .B2(n465), .A(n789), .ZN(n621) );
  NAND2_X1 U274 ( .A1(\mem[1][9] ), .A2(n465), .ZN(n789) );
  OAI21_X1 U275 ( .B1(n480), .B2(n799), .A(n788), .ZN(n620) );
  NAND2_X1 U276 ( .A1(\mem[1][10] ), .A2(n465), .ZN(n788) );
  OAI21_X1 U277 ( .B1(n479), .B2(n799), .A(n787), .ZN(n619) );
  NAND2_X1 U278 ( .A1(\mem[1][11] ), .A2(n465), .ZN(n787) );
  OAI21_X1 U279 ( .B1(n490), .B2(n464), .A(n777), .ZN(n610) );
  NAND2_X1 U280 ( .A1(\mem[2][0] ), .A2(n778), .ZN(n777) );
  OAI21_X1 U281 ( .B1(n489), .B2(n464), .A(n776), .ZN(n609) );
  NAND2_X1 U282 ( .A1(\mem[2][1] ), .A2(n778), .ZN(n776) );
  OAI21_X1 U283 ( .B1(n488), .B2(n464), .A(n775), .ZN(n608) );
  NAND2_X1 U284 ( .A1(\mem[2][2] ), .A2(n778), .ZN(n775) );
  OAI21_X1 U285 ( .B1(n487), .B2(n464), .A(n774), .ZN(n607) );
  NAND2_X1 U286 ( .A1(\mem[2][3] ), .A2(n778), .ZN(n774) );
  OAI21_X1 U287 ( .B1(n486), .B2(n464), .A(n773), .ZN(n606) );
  NAND2_X1 U288 ( .A1(\mem[2][4] ), .A2(n778), .ZN(n773) );
  OAI21_X1 U289 ( .B1(n485), .B2(n464), .A(n772), .ZN(n605) );
  NAND2_X1 U290 ( .A1(\mem[2][5] ), .A2(n778), .ZN(n772) );
  OAI21_X1 U291 ( .B1(n484), .B2(n464), .A(n771), .ZN(n604) );
  NAND2_X1 U292 ( .A1(\mem[2][6] ), .A2(n778), .ZN(n771) );
  OAI21_X1 U293 ( .B1(n483), .B2(n464), .A(n770), .ZN(n603) );
  NAND2_X1 U294 ( .A1(\mem[2][7] ), .A2(n778), .ZN(n770) );
  OAI21_X1 U295 ( .B1(n482), .B2(n464), .A(n769), .ZN(n602) );
  NAND2_X1 U296 ( .A1(\mem[2][8] ), .A2(n778), .ZN(n769) );
  OAI21_X1 U297 ( .B1(n481), .B2(n778), .A(n768), .ZN(n601) );
  NAND2_X1 U298 ( .A1(\mem[2][9] ), .A2(n778), .ZN(n768) );
  OAI21_X1 U299 ( .B1(n480), .B2(n464), .A(n767), .ZN(n600) );
  NAND2_X1 U300 ( .A1(\mem[2][10] ), .A2(n778), .ZN(n767) );
  OAI21_X1 U301 ( .B1(n479), .B2(n464), .A(n766), .ZN(n599) );
  NAND2_X1 U302 ( .A1(\mem[2][11] ), .A2(n778), .ZN(n766) );
  OAI21_X1 U303 ( .B1(n490), .B2(n757), .A(n756), .ZN(n590) );
  NAND2_X1 U304 ( .A1(\mem[3][0] ), .A2(n757), .ZN(n756) );
  OAI21_X1 U305 ( .B1(n489), .B2(n757), .A(n755), .ZN(n589) );
  NAND2_X1 U306 ( .A1(\mem[3][1] ), .A2(n463), .ZN(n755) );
  OAI21_X1 U307 ( .B1(n488), .B2(n757), .A(n754), .ZN(n588) );
  NAND2_X1 U308 ( .A1(\mem[3][2] ), .A2(n463), .ZN(n754) );
  OAI21_X1 U309 ( .B1(n487), .B2(n757), .A(n753), .ZN(n587) );
  NAND2_X1 U310 ( .A1(\mem[3][3] ), .A2(n463), .ZN(n753) );
  OAI21_X1 U311 ( .B1(n486), .B2(n757), .A(n752), .ZN(n586) );
  NAND2_X1 U312 ( .A1(\mem[3][4] ), .A2(n463), .ZN(n752) );
  OAI21_X1 U313 ( .B1(n485), .B2(n757), .A(n751), .ZN(n585) );
  NAND2_X1 U314 ( .A1(\mem[3][5] ), .A2(n463), .ZN(n751) );
  OAI21_X1 U315 ( .B1(n484), .B2(n757), .A(n750), .ZN(n584) );
  NAND2_X1 U316 ( .A1(\mem[3][6] ), .A2(n463), .ZN(n750) );
  OAI21_X1 U317 ( .B1(n483), .B2(n757), .A(n749), .ZN(n583) );
  NAND2_X1 U318 ( .A1(\mem[3][7] ), .A2(n463), .ZN(n749) );
  OAI21_X1 U319 ( .B1(n482), .B2(n757), .A(n748), .ZN(n582) );
  NAND2_X1 U320 ( .A1(\mem[3][8] ), .A2(n463), .ZN(n748) );
  OAI21_X1 U321 ( .B1(n481), .B2(n757), .A(n747), .ZN(n581) );
  NAND2_X1 U322 ( .A1(\mem[3][9] ), .A2(n463), .ZN(n747) );
  OAI21_X1 U323 ( .B1(n480), .B2(n757), .A(n746), .ZN(n580) );
  NAND2_X1 U324 ( .A1(\mem[3][10] ), .A2(n463), .ZN(n746) );
  OAI21_X1 U325 ( .B1(n479), .B2(n757), .A(n745), .ZN(n579) );
  NAND2_X1 U326 ( .A1(\mem[3][11] ), .A2(n463), .ZN(n745) );
  OAI21_X1 U327 ( .B1(n466), .B2(n478), .A(n808), .ZN(n638) );
  NAND2_X1 U328 ( .A1(\mem[0][12] ), .A2(n466), .ZN(n808) );
  OAI21_X1 U329 ( .B1(n466), .B2(n477), .A(n807), .ZN(n637) );
  NAND2_X1 U330 ( .A1(\mem[0][13] ), .A2(n466), .ZN(n807) );
  OAI21_X1 U331 ( .B1(n466), .B2(n476), .A(n806), .ZN(n636) );
  NAND2_X1 U332 ( .A1(\mem[0][14] ), .A2(n466), .ZN(n806) );
  OAI21_X1 U333 ( .B1(n821), .B2(n475), .A(n805), .ZN(n635) );
  NAND2_X1 U334 ( .A1(\mem[0][15] ), .A2(n466), .ZN(n805) );
  OAI21_X1 U335 ( .B1(n821), .B2(n474), .A(n804), .ZN(n634) );
  NAND2_X1 U336 ( .A1(\mem[0][16] ), .A2(n466), .ZN(n804) );
  OAI21_X1 U337 ( .B1(n821), .B2(n473), .A(n803), .ZN(n633) );
  NAND2_X1 U338 ( .A1(\mem[0][17] ), .A2(n466), .ZN(n803) );
  OAI21_X1 U339 ( .B1(n821), .B2(n472), .A(n802), .ZN(n632) );
  NAND2_X1 U340 ( .A1(\mem[0][18] ), .A2(n466), .ZN(n802) );
  OAI21_X1 U341 ( .B1(n821), .B2(n471), .A(n801), .ZN(n631) );
  NAND2_X1 U342 ( .A1(\mem[0][19] ), .A2(n466), .ZN(n801) );
  INV_X1 U343 ( .A(data_in[0]), .ZN(n490) );
  INV_X1 U344 ( .A(data_in[1]), .ZN(n489) );
  INV_X1 U345 ( .A(data_in[2]), .ZN(n488) );
  INV_X1 U346 ( .A(data_in[3]), .ZN(n487) );
  INV_X1 U347 ( .A(data_in[4]), .ZN(n486) );
  INV_X1 U348 ( .A(data_in[5]), .ZN(n485) );
  INV_X1 U349 ( .A(data_in[6]), .ZN(n484) );
  INV_X1 U358 ( .A(data_in[7]), .ZN(n483) );
  INV_X1 U359 ( .A(data_in[8]), .ZN(n482) );
  INV_X1 U360 ( .A(data_in[9]), .ZN(n481) );
  INV_X1 U361 ( .A(data_in[10]), .ZN(n480) );
  INV_X1 U362 ( .A(data_in[11]), .ZN(n479) );
  INV_X1 U363 ( .A(data_in[12]), .ZN(n478) );
  INV_X1 U364 ( .A(data_in[13]), .ZN(n477) );
  INV_X1 U365 ( .A(data_in[14]), .ZN(n476) );
  INV_X1 U366 ( .A(data_in[15]), .ZN(n475) );
  INV_X1 U367 ( .A(data_in[16]), .ZN(n474) );
  INV_X1 U368 ( .A(data_in[17]), .ZN(n473) );
  INV_X1 U369 ( .A(data_in[18]), .ZN(n472) );
  INV_X1 U370 ( .A(data_in[19]), .ZN(n471) );
  MUX2_X1 U371 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n455), .Z(n2) );
  MUX2_X1 U372 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n455), .Z(n3) );
  MUX2_X1 U373 ( .A(n3), .B(n2), .S(n454), .Z(n4) );
  MUX2_X1 U374 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n455), .Z(n5) );
  MUX2_X1 U375 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n455), .Z(n6) );
  MUX2_X1 U376 ( .A(n6), .B(n5), .S(n454), .Z(n7) );
  MUX2_X1 U377 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n455), .Z(n8) );
  MUX2_X1 U378 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n455), .Z(n9) );
  MUX2_X1 U379 ( .A(n9), .B(n8), .S(n454), .Z(n10) );
  MUX2_X1 U380 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n455), .Z(n11) );
  MUX2_X1 U381 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n455), .Z(n12) );
  MUX2_X1 U382 ( .A(n12), .B(n11), .S(n454), .Z(n13) );
  MUX2_X1 U383 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n456), .Z(n14) );
  MUX2_X1 U384 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n456), .Z(n15) );
  MUX2_X1 U385 ( .A(n15), .B(n14), .S(n454), .Z(n16) );
  MUX2_X1 U386 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n456), .Z(n17) );
  MUX2_X1 U387 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n456), .Z(n18) );
  MUX2_X1 U388 ( .A(n18), .B(n17), .S(n454), .Z(n19) );
  MUX2_X1 U389 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n456), .Z(n20) );
  MUX2_X1 U390 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n456), .Z(n21) );
  MUX2_X1 U391 ( .A(n21), .B(n20), .S(n453), .Z(n22) );
  MUX2_X1 U392 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n456), .Z(n23) );
  MUX2_X1 U393 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n456), .Z(n24) );
  MUX2_X1 U394 ( .A(n24), .B(n23), .S(n454), .Z(n356) );
  MUX2_X1 U395 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n456), .Z(n357) );
  MUX2_X1 U396 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n456), .Z(n358) );
  MUX2_X1 U397 ( .A(n358), .B(n357), .S(n453), .Z(n359) );
  MUX2_X1 U398 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n456), .Z(n360) );
  MUX2_X1 U399 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n456), .Z(n361) );
  MUX2_X1 U400 ( .A(n361), .B(n360), .S(n454), .Z(n362) );
  MUX2_X1 U401 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n455), .Z(n363) );
  MUX2_X1 U402 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n455), .Z(n364) );
  MUX2_X1 U403 ( .A(n364), .B(n363), .S(n453), .Z(n365) );
  MUX2_X1 U404 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n456), .Z(n366) );
  MUX2_X1 U405 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n456), .Z(n367) );
  MUX2_X1 U406 ( .A(n367), .B(n366), .S(n454), .Z(n368) );
  MUX2_X1 U407 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n456), .Z(n369) );
  MUX2_X1 U408 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n456), .Z(n370) );
  MUX2_X1 U409 ( .A(n370), .B(n369), .S(N11), .Z(n371) );
  MUX2_X1 U410 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n458), .Z(n372) );
  MUX2_X1 U411 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n458), .Z(n373) );
  MUX2_X1 U412 ( .A(n373), .B(n372), .S(n454), .Z(n374) );
  MUX2_X1 U413 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n458), .Z(n375) );
  MUX2_X1 U414 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n458), .Z(n376) );
  MUX2_X1 U415 ( .A(n376), .B(n375), .S(N11), .Z(n377) );
  MUX2_X1 U416 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n457), .Z(n378) );
  MUX2_X1 U417 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n457), .Z(n379) );
  MUX2_X1 U418 ( .A(n379), .B(n378), .S(n454), .Z(n380) );
  MUX2_X1 U419 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n458), .Z(n381) );
  MUX2_X1 U420 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n457), .Z(n382) );
  MUX2_X1 U421 ( .A(n382), .B(n381), .S(n454), .Z(n383) );
  MUX2_X1 U422 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n456), .Z(n384) );
  MUX2_X1 U423 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n456), .Z(n385) );
  MUX2_X1 U424 ( .A(n385), .B(n384), .S(n453), .Z(n386) );
  MUX2_X1 U425 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n457), .Z(n387) );
  MUX2_X1 U426 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n455), .Z(n388) );
  MUX2_X1 U427 ( .A(n388), .B(n387), .S(n454), .Z(n389) );
  MUX2_X1 U428 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n456), .Z(n390) );
  MUX2_X1 U429 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n456), .Z(n391) );
  MUX2_X1 U430 ( .A(n391), .B(n390), .S(n454), .Z(n392) );
  MUX2_X1 U431 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n455), .Z(n393) );
  MUX2_X1 U432 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n457), .Z(n394) );
  MUX2_X1 U433 ( .A(n394), .B(n393), .S(n454), .Z(n395) );
  MUX2_X1 U434 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n455), .Z(n396) );
  MUX2_X1 U435 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n458), .Z(n397) );
  MUX2_X1 U436 ( .A(n397), .B(n396), .S(n454), .Z(n398) );
  MUX2_X1 U437 ( .A(n398), .B(n395), .S(N12), .Z(N22) );
  MUX2_X1 U438 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n457), .Z(n399) );
  MUX2_X1 U439 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n456), .Z(n400) );
  MUX2_X1 U440 ( .A(n400), .B(n399), .S(n454), .Z(n401) );
  MUX2_X1 U441 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n455), .Z(n402) );
  MUX2_X1 U442 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n457), .Z(n403) );
  MUX2_X1 U443 ( .A(n403), .B(n402), .S(n454), .Z(n404) );
  MUX2_X1 U444 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n457), .Z(n405) );
  MUX2_X1 U445 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n455), .Z(n406) );
  MUX2_X1 U446 ( .A(n406), .B(n405), .S(n454), .Z(n407) );
  MUX2_X1 U447 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n455), .Z(n408) );
  MUX2_X1 U448 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n458), .Z(n409) );
  MUX2_X1 U449 ( .A(n409), .B(n408), .S(n454), .Z(n410) );
  MUX2_X1 U450 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n458), .Z(n411) );
  MUX2_X1 U451 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n455), .Z(n412) );
  MUX2_X1 U452 ( .A(n412), .B(n411), .S(n454), .Z(n413) );
  MUX2_X1 U453 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n455), .Z(n414) );
  MUX2_X1 U454 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n456), .Z(n415) );
  MUX2_X1 U455 ( .A(n415), .B(n414), .S(n454), .Z(n416) );
  MUX2_X1 U456 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n457), .Z(n417) );
  MUX2_X1 U457 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n457), .Z(n418) );
  MUX2_X1 U458 ( .A(n418), .B(n417), .S(n453), .Z(n419) );
  MUX2_X1 U459 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n457), .Z(n420) );
  MUX2_X1 U460 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n457), .Z(n421) );
  MUX2_X1 U461 ( .A(n421), .B(n420), .S(n453), .Z(n422) );
  MUX2_X1 U462 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n457), .Z(n423) );
  MUX2_X1 U463 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n457), .Z(n424) );
  MUX2_X1 U464 ( .A(n424), .B(n423), .S(n453), .Z(n425) );
  MUX2_X1 U465 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n457), .Z(n426) );
  MUX2_X1 U466 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n457), .Z(n427) );
  MUX2_X1 U467 ( .A(n427), .B(n426), .S(n453), .Z(n428) );
  MUX2_X1 U468 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n457), .Z(n429) );
  MUX2_X1 U469 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n457), .Z(n430) );
  MUX2_X1 U470 ( .A(n430), .B(n429), .S(n453), .Z(n431) );
  MUX2_X1 U471 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n457), .Z(n432) );
  MUX2_X1 U472 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n457), .Z(n433) );
  MUX2_X1 U473 ( .A(n433), .B(n432), .S(n453), .Z(n434) );
  MUX2_X1 U474 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n458), .Z(n435) );
  MUX2_X1 U475 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n458), .Z(n436) );
  MUX2_X1 U476 ( .A(n436), .B(n435), .S(n453), .Z(n437) );
  MUX2_X1 U477 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n458), .Z(n438) );
  MUX2_X1 U478 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n458), .Z(n439) );
  MUX2_X1 U479 ( .A(n439), .B(n438), .S(n453), .Z(n440) );
  MUX2_X1 U480 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n458), .Z(n441) );
  MUX2_X1 U481 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n458), .Z(n442) );
  MUX2_X1 U482 ( .A(n442), .B(n441), .S(n453), .Z(n443) );
  MUX2_X1 U483 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n458), .Z(n444) );
  MUX2_X1 U484 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n458), .Z(n445) );
  MUX2_X1 U485 ( .A(n445), .B(n444), .S(n453), .Z(n446) );
  MUX2_X1 U486 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n458), .Z(n447) );
  MUX2_X1 U487 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n458), .Z(n448) );
  MUX2_X1 U488 ( .A(n448), .B(n447), .S(n453), .Z(n449) );
  MUX2_X1 U489 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n458), .Z(n450) );
  MUX2_X1 U490 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n458), .Z(n451) );
  MUX2_X1 U491 ( .A(n451), .B(n450), .S(n453), .Z(n452) );
  CLKBUF_X1 U492 ( .A(N10), .Z(n455) );
endmodule


module mac_7_DW_mult_tc_1 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n4, n6, n7, n9, n12, n13, n16, n18, n19, n22, n25, n28, n30, n31,
         n34, n36, n37, n40, n42, n43, n46, n48, n49, n52, n55, n58, n60, n61,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n97, n98, n99, n100, n101, n103, n105, n106, n107,
         n108, n109, n111, n113, n114, n115, n116, n117, n119, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n139, n140, n141, n142, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n183, n185, n186, n187, n188, n193, n194, n195, n196, n198,
         n200, n201, n202, n203, n204, n205, n206, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n227, n228, n230, n232, n233, n234, n236, n238, n239, n240,
         n241, n242, n244, n246, n247, n248, n249, n250, n252, n254, n255,
         n256, n257, n258, n259, n260, n261, n263, n264, n266, n268, n270,
         n271, n272, n273, n274, n275, n277, n278, n279, n280, n282, n285,
         n286, n287, n291, n293, n295, n296, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n643, n644, n646, n647, n649,
         n650, n652, n653, n655, n656, n658, n659, n661, n662, n664, n665,
         n667, n668, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1116, n1119, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n37 = a[13];
  assign n43 = a[15];
  assign n49 = a[17];
  assign n55 = a[19];
  assign n61 = b[0];
  assign n668 = a[0];
  assign n1090 = b[19];
  assign n1091 = b[18];
  assign n1092 = b[17];
  assign n1093 = b[16];
  assign n1094 = b[15];
  assign n1095 = b[14];
  assign n1096 = b[13];
  assign n1097 = b[12];
  assign n1098 = b[11];
  assign n1099 = b[10];
  assign n1100 = b[9];
  assign n1101 = b[8];
  assign n1102 = b[7];
  assign n1103 = b[6];
  assign n1104 = b[5];
  assign n1105 = b[4];
  assign n1106 = b[3];
  assign n1107 = b[2];
  assign n1108 = b[1];

  FA_X1 U333 ( .A(n681), .B(n304), .CI(n700), .CO(n300), .S(n301) );
  FA_X1 U334 ( .A(n305), .B(n682), .CI(n308), .CO(n302), .S(n303) );
  FA_X1 U336 ( .A(n312), .B(n683), .CI(n309), .CO(n306), .S(n307) );
  FA_X1 U337 ( .A(n701), .B(n314), .CI(n720), .CO(n308), .S(n309) );
  FA_X1 U338 ( .A(n313), .B(n320), .CI(n318), .CO(n310), .S(n311) );
  FA_X1 U339 ( .A(n684), .B(n702), .CI(n315), .CO(n312), .S(n313) );
  FA_X1 U341 ( .A(n324), .B(n321), .CI(n319), .CO(n316), .S(n317) );
  FA_X1 U342 ( .A(n328), .B(n721), .CI(n326), .CO(n318), .S(n319) );
  FA_X1 U343 ( .A(n703), .B(n685), .CI(n740), .CO(n320), .S(n321) );
  FA_X1 U344 ( .A(n325), .B(n327), .CI(n332), .CO(n322), .S(n323) );
  FA_X1 U345 ( .A(n336), .B(n329), .CI(n334), .CO(n324), .S(n325) );
  FA_X1 U346 ( .A(n686), .B(n704), .CI(n722), .CO(n326), .S(n327) );
  FA_X1 U348 ( .A(n340), .B(n342), .CI(n333), .CO(n330), .S(n331) );
  FA_X1 U349 ( .A(n335), .B(n344), .CI(n337), .CO(n332), .S(n333) );
  FA_X1 U350 ( .A(n705), .B(n346), .CI(n723), .CO(n334), .S(n335) );
  FA_X1 U351 ( .A(n741), .B(n687), .CI(n760), .CO(n336), .S(n337) );
  FA_X1 U352 ( .A(n350), .B(n343), .CI(n341), .CO(n338), .S(n339) );
  FA_X1 U353 ( .A(n345), .B(n354), .CI(n352), .CO(n340), .S(n341) );
  FA_X1 U354 ( .A(n347), .B(n724), .CI(n356), .CO(n342), .S(n343) );
  FA_X1 U355 ( .A(n742), .B(n706), .CI(n688), .CO(n344), .S(n345) );
  FA_X1 U357 ( .A(n360), .B(n353), .CI(n351), .CO(n348), .S(n349) );
  FA_X1 U358 ( .A(n357), .B(n355), .CI(n362), .CO(n350), .S(n351) );
  FA_X1 U359 ( .A(n366), .B(n743), .CI(n364), .CO(n352), .S(n353) );
  FA_X1 U360 ( .A(n707), .B(n761), .CI(n725), .CO(n354), .S(n355) );
  FA_X1 U361 ( .A(n368), .B(n689), .CI(n780), .CO(n356), .S(n357) );
  FA_X1 U362 ( .A(n372), .B(n363), .CI(n361), .CO(n358), .S(n359) );
  FA_X1 U363 ( .A(n376), .B(n365), .CI(n374), .CO(n360), .S(n361) );
  FA_X1 U364 ( .A(n378), .B(n380), .CI(n367), .CO(n362), .S(n363) );
  FA_X1 U365 ( .A(n690), .B(n708), .CI(n369), .CO(n364), .S(n365) );
  FA_X1 U366 ( .A(n762), .B(n726), .CI(n744), .CO(n366), .S(n367) );
  FA_X1 U368 ( .A(n384), .B(n375), .CI(n373), .CO(n370), .S(n371) );
  FA_X1 U369 ( .A(n377), .B(n388), .CI(n386), .CO(n372), .S(n373) );
  FA_X1 U370 ( .A(n379), .B(n390), .CI(n381), .CO(n374), .S(n375) );
  FA_X1 U371 ( .A(n727), .B(n745), .CI(n392), .CO(n376), .S(n377) );
  FA_X1 U372 ( .A(n709), .B(n781), .CI(n763), .CO(n378), .S(n379) );
  FA_X1 U373 ( .A(n394), .B(n691), .CI(n800), .CO(n380), .S(n381) );
  FA_X1 U374 ( .A(n398), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U376 ( .A(n391), .B(n404), .CI(n393), .CO(n386), .S(n387) );
  FA_X1 U377 ( .A(n408), .B(n395), .CI(n406), .CO(n388), .S(n389) );
  FA_X1 U378 ( .A(n746), .B(n782), .CI(n764), .CO(n390), .S(n391) );
  FA_X1 U379 ( .A(n692), .B(n728), .CI(n710), .CO(n392), .S(n393) );
  FA_X1 U381 ( .A(n412), .B(n401), .CI(n399), .CO(n396), .S(n397) );
  FA_X1 U382 ( .A(n403), .B(n416), .CI(n414), .CO(n398), .S(n399) );
  FA_X1 U383 ( .A(n409), .B(n407), .CI(n418), .CO(n400), .S(n401) );
  FA_X1 U384 ( .A(n420), .B(n422), .CI(n405), .CO(n402), .S(n403) );
  FA_X1 U385 ( .A(n729), .B(n765), .CI(n747), .CO(n404), .S(n405) );
  FA_X1 U386 ( .A(n711), .B(n801), .CI(n783), .CO(n406), .S(n407) );
  FA_X1 U387 ( .A(n820), .B(n424), .CI(n693), .CO(n408), .S(n409) );
  FA_X1 U390 ( .A(n419), .B(n423), .CI(n434), .CO(n414), .S(n415) );
  FA_X1 U391 ( .A(n436), .B(n438), .CI(n421), .CO(n416), .S(n417) );
  FA_X1 U393 ( .A(n694), .B(n766), .CI(n712), .CO(n420), .S(n421) );
  FA_X1 U394 ( .A(n802), .B(n730), .CI(n784), .CO(n422), .S(n423) );
  FA_X1 U398 ( .A(n450), .B(n441), .CI(n435), .CO(n430), .S(n431) );
  FA_X1 U399 ( .A(n437), .B(n452), .CI(n439), .CO(n432), .S(n433) );
  FA_X1 U400 ( .A(n456), .B(n767), .CI(n454), .CO(n434), .S(n435) );
  FA_X1 U401 ( .A(n731), .B(n785), .CI(n749), .CO(n436), .S(n437) );
  FA_X1 U402 ( .A(n458), .B(n803), .CI(n713), .CO(n438), .S(n439) );
  FA_X1 U404 ( .A(n462), .B(n447), .CI(n445), .CO(n442), .S(n443) );
  FA_X1 U405 ( .A(n449), .B(n466), .CI(n464), .CO(n444), .S(n445) );
  FA_X1 U406 ( .A(n468), .B(n453), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U407 ( .A(n455), .B(n470), .CI(n457), .CO(n448), .S(n449) );
  FA_X1 U408 ( .A(n474), .B(n476), .CI(n472), .CO(n450), .S(n451) );
  FA_X1 U409 ( .A(n768), .B(n786), .CI(n459), .CO(n452), .S(n453) );
  FA_X1 U410 ( .A(n732), .B(n804), .CI(n714), .CO(n454), .S(n455) );
  FA_X1 U411 ( .A(n822), .B(n750), .CI(n696), .CO(n456), .S(n457) );
  FA_X1 U416 ( .A(n473), .B(n488), .CI(n475), .CO(n466), .S(n467) );
  FA_X1 U417 ( .A(n477), .B(n490), .CI(n492), .CO(n468), .S(n469) );
  FA_X1 U419 ( .A(n841), .B(n733), .CI(n751), .CO(n472), .S(n473) );
  FA_X1 U420 ( .A(n860), .B(n769), .CI(n697), .CO(n474), .S(n475) );
  FA_X1 U423 ( .A(n498), .B(n483), .CI(n481), .CO(n478), .S(n479) );
  FA_X1 U425 ( .A(n504), .B(n493), .CI(n502), .CO(n482), .S(n483) );
  FA_X1 U426 ( .A(n489), .B(n506), .CI(n491), .CO(n484), .S(n485) );
  FA_X1 U427 ( .A(n510), .B(n495), .CI(n508), .CO(n486), .S(n487) );
  FA_X1 U428 ( .A(n770), .B(n824), .CI(n842), .CO(n488), .S(n489) );
  FA_X1 U429 ( .A(n752), .B(n806), .CI(n861), .CO(n490), .S(n491) );
  FA_X1 U430 ( .A(n670), .B(n734), .CI(n788), .CO(n492), .S(n493) );
  HA_X1 U431 ( .A(n716), .B(n698), .CO(n494), .S(n495) );
  FA_X1 U433 ( .A(n516), .B(n505), .CI(n503), .CO(n498), .S(n499) );
  FA_X1 U435 ( .A(n511), .B(n522), .CI(n507), .CO(n502), .S(n503) );
  FA_X1 U436 ( .A(n526), .B(n807), .CI(n524), .CO(n504), .S(n505) );
  FA_X1 U437 ( .A(n771), .B(n825), .CI(n789), .CO(n506), .S(n507) );
  FA_X1 U438 ( .A(n753), .B(n843), .CI(n717), .CO(n508), .S(n509) );
  FA_X1 U439 ( .A(n862), .B(n699), .CI(n735), .CO(n510), .S(n511) );
  FA_X1 U442 ( .A(n525), .B(n523), .CI(n534), .CO(n516), .S(n517) );
  FA_X1 U443 ( .A(n536), .B(n540), .CI(n538), .CO(n518), .S(n519) );
  FA_X1 U444 ( .A(n826), .B(n844), .CI(n527), .CO(n520), .S(n521) );
  FA_X1 U445 ( .A(n754), .B(n772), .CI(n808), .CO(n522), .S(n523) );
  FA_X1 U446 ( .A(n863), .B(n790), .CI(n671), .CO(n524), .S(n525) );
  HA_X1 U447 ( .A(n718), .B(n736), .CO(n526), .S(n527) );
  FA_X1 U450 ( .A(n537), .B(n541), .CI(n539), .CO(n532), .S(n533) );
  FA_X1 U451 ( .A(n552), .B(n554), .CI(n550), .CO(n534), .S(n535) );
  FA_X1 U452 ( .A(n809), .B(n827), .CI(n791), .CO(n536), .S(n537) );
  FA_X1 U453 ( .A(n773), .B(n845), .CI(n737), .CO(n538), .S(n539) );
  FA_X1 U454 ( .A(n864), .B(n719), .CI(n755), .CO(n540), .S(n541) );
  FA_X1 U455 ( .A(n547), .B(n558), .CI(n545), .CO(n542), .S(n543) );
  FA_X1 U456 ( .A(n549), .B(n553), .CI(n560), .CO(n544), .S(n545) );
  FA_X1 U457 ( .A(n562), .B(n564), .CI(n551), .CO(n546), .S(n547) );
  FA_X1 U458 ( .A(n555), .B(n846), .CI(n566), .CO(n548), .S(n549) );
  FA_X1 U459 ( .A(n865), .B(n792), .CI(n828), .CO(n550), .S(n551) );
  FA_X1 U460 ( .A(n774), .B(n810), .CI(n672), .CO(n552), .S(n553) );
  HA_X1 U461 ( .A(n756), .B(n738), .CO(n554), .S(n555) );
  FA_X1 U463 ( .A(n563), .B(n565), .CI(n572), .CO(n558), .S(n559) );
  FA_X1 U464 ( .A(n574), .B(n576), .CI(n567), .CO(n560), .S(n561) );
  FA_X1 U465 ( .A(n811), .B(n829), .CI(n578), .CO(n562), .S(n563) );
  FA_X1 U466 ( .A(n757), .B(n847), .CI(n793), .CO(n564), .S(n565) );
  FA_X1 U467 ( .A(n775), .B(n739), .CI(n866), .CO(n566), .S(n567) );
  FA_X1 U468 ( .A(n582), .B(n573), .CI(n571), .CO(n568), .S(n569) );
  FA_X1 U469 ( .A(n577), .B(n575), .CI(n584), .CO(n570), .S(n571) );
  FA_X1 U470 ( .A(n588), .B(n579), .CI(n586), .CO(n572), .S(n573) );
  FA_X1 U471 ( .A(n794), .B(n848), .CI(n830), .CO(n574), .S(n575) );
  FA_X1 U472 ( .A(n867), .B(n812), .CI(n673), .CO(n576), .S(n577) );
  HA_X1 U473 ( .A(n758), .B(n776), .CO(n578), .S(n579) );
  FA_X1 U476 ( .A(n598), .B(n831), .CI(n596), .CO(n584), .S(n585) );
  FA_X1 U477 ( .A(n777), .B(n849), .CI(n813), .CO(n586), .S(n587) );
  FA_X1 U478 ( .A(n795), .B(n759), .CI(n868), .CO(n588), .S(n589) );
  FA_X1 U479 ( .A(n602), .B(n595), .CI(n593), .CO(n590), .S(n591) );
  FA_X1 U480 ( .A(n604), .B(n606), .CI(n597), .CO(n592), .S(n593) );
  FA_X1 U481 ( .A(n814), .B(n850), .CI(n599), .CO(n594), .S(n595) );
  FA_X1 U482 ( .A(n869), .B(n832), .CI(n674), .CO(n596), .S(n597) );
  HA_X1 U483 ( .A(n796), .B(n778), .CO(n598), .S(n599) );
  FA_X1 U484 ( .A(n610), .B(n605), .CI(n603), .CO(n600), .S(n601) );
  FA_X1 U485 ( .A(n612), .B(n614), .CI(n607), .CO(n602), .S(n603) );
  FA_X1 U486 ( .A(n797), .B(n851), .CI(n833), .CO(n604), .S(n605) );
  FA_X1 U487 ( .A(n779), .B(n815), .CI(n870), .CO(n606), .S(n607) );
  FA_X1 U488 ( .A(n613), .B(n618), .CI(n611), .CO(n608), .S(n609) );
  FA_X1 U489 ( .A(n615), .B(n871), .CI(n620), .CO(n610), .S(n611) );
  FA_X1 U490 ( .A(n675), .B(n834), .CI(n852), .CO(n612), .S(n613) );
  HA_X1 U491 ( .A(n798), .B(n816), .CO(n614), .S(n615) );
  FA_X1 U492 ( .A(n621), .B(n624), .CI(n619), .CO(n616), .S(n617) );
  FA_X1 U493 ( .A(n817), .B(n853), .CI(n626), .CO(n618), .S(n619) );
  FA_X1 U494 ( .A(n835), .B(n799), .CI(n872), .CO(n620), .S(n621) );
  FA_X1 U495 ( .A(n630), .B(n627), .CI(n625), .CO(n622), .S(n623) );
  FA_X1 U496 ( .A(n854), .B(n873), .CI(n676), .CO(n624), .S(n625) );
  HA_X1 U497 ( .A(n818), .B(n836), .CO(n626), .S(n627) );
  FA_X1 U498 ( .A(n634), .B(n837), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U499 ( .A(n874), .B(n819), .CI(n855), .CO(n630), .S(n631) );
  FA_X1 U500 ( .A(n677), .B(n856), .CI(n635), .CO(n632), .S(n633) );
  HA_X1 U501 ( .A(n838), .B(n875), .CO(n634), .S(n635) );
  FA_X1 U502 ( .A(n876), .B(n839), .CI(n857), .CO(n636), .S(n637) );
  HA_X1 U503 ( .A(n877), .B(n858), .CO(n638), .S(n639) );
  NAND2_X1 U1025 ( .A1(n52), .A2(n1490), .ZN(n1233) );
  NAND2_X1 U1026 ( .A1(n52), .A2(n1490), .ZN(n1234) );
  AND2_X1 U1027 ( .A1(n601), .A2(n608), .ZN(n1271) );
  BUF_X1 U1028 ( .A(n1108), .Z(n1529) );
  BUF_X2 U1029 ( .A(n1102), .Z(n1535) );
  BUF_X1 U1030 ( .A(n1097), .Z(n1310) );
  CLKBUF_X3 U1031 ( .A(n37), .Z(n1352) );
  BUF_X2 U1032 ( .A(n1095), .Z(n1541) );
  BUF_X2 U1033 ( .A(n13), .Z(n1524) );
  BUF_X2 U1034 ( .A(n13), .Z(n1340) );
  BUF_X2 U1035 ( .A(n1100), .Z(n1537) );
  BUF_X1 U1036 ( .A(n1097), .Z(n1311) );
  BUF_X2 U1037 ( .A(n16), .Z(n1409) );
  BUF_X2 U1038 ( .A(n22), .Z(n1509) );
  BUF_X2 U1039 ( .A(n1094), .Z(n1542) );
  BUF_X2 U1040 ( .A(n43), .Z(n1431) );
  BUF_X1 U1041 ( .A(n43), .Z(n1526) );
  BUF_X2 U1042 ( .A(n1092), .Z(n1544) );
  BUF_X2 U1043 ( .A(n1), .Z(n1383) );
  BUF_X2 U1044 ( .A(n1511), .Z(n1357) );
  BUF_X2 U1045 ( .A(n22), .Z(n1510) );
  CLKBUF_X3 U1046 ( .A(n61), .Z(n1527) );
  BUF_X2 U1047 ( .A(n1), .Z(n1305) );
  AND2_X1 U1048 ( .A1(n529), .A2(n542), .ZN(n1416) );
  INV_X1 U1049 ( .A(n1416), .ZN(n188) );
  INV_X1 U1050 ( .A(n1271), .ZN(n227) );
  BUF_X1 U1051 ( .A(n9), .Z(n1511) );
  CLKBUF_X1 U1052 ( .A(n242), .Z(n1235) );
  AOI21_X1 U1053 ( .B1(n1499), .B2(n255), .A(n252), .ZN(n1236) );
  BUF_X2 U1054 ( .A(n1091), .Z(n1545) );
  OR2_X1 U1055 ( .A1(n557), .A2(n568), .ZN(n1237) );
  OR2_X1 U1056 ( .A1(n427), .A2(n442), .ZN(n1238) );
  OR2_X1 U1057 ( .A1(n679), .A2(n879), .ZN(n1239) );
  AND2_X1 U1058 ( .A1(n1239), .A2(n263), .ZN(product[1]) );
  BUF_X2 U1059 ( .A(n12), .Z(n1244) );
  XNOR2_X1 U1060 ( .A(n446), .B(n1241), .ZN(n429) );
  XNOR2_X1 U1061 ( .A(n433), .B(n448), .ZN(n1241) );
  BUF_X1 U1062 ( .A(n1106), .Z(n1359) );
  OAI22_X1 U1063 ( .A1(n1404), .A2(n993), .B1(n992), .B2(n1413), .ZN(n1242) );
  BUF_X1 U1064 ( .A(n30), .Z(n1404) );
  BUF_X1 U1065 ( .A(n12), .Z(n1364) );
  CLKBUF_X1 U1066 ( .A(n430), .Z(n1243) );
  NAND2_X1 U1067 ( .A1(n1116), .A2(n1303), .ZN(n1406) );
  BUF_X2 U1068 ( .A(n30), .Z(n1405) );
  BUF_X2 U1069 ( .A(n28), .Z(n1414) );
  XNOR2_X1 U1070 ( .A(n1245), .B(n1246), .ZN(n419) );
  XOR2_X1 U1071 ( .A(n425), .B(n748), .Z(n1245) );
  AND3_X1 U1072 ( .A1(n1475), .A2(n1476), .A3(n1477), .ZN(n1246) );
  XNOR2_X1 U1073 ( .A(n1538), .B(n1305), .ZN(n1247) );
  CLKBUF_X3 U1074 ( .A(n7), .Z(n1523) );
  CLKBUF_X3 U1075 ( .A(n7), .Z(n1319) );
  INV_X1 U1076 ( .A(n1331), .ZN(n1248) );
  BUF_X2 U1077 ( .A(n4), .Z(n1331) );
  NAND3_X1 U1078 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1249) );
  BUF_X2 U1079 ( .A(n49), .Z(n1401) );
  XNOR2_X1 U1080 ( .A(n1250), .B(n482), .ZN(n463) );
  XNOR2_X1 U1081 ( .A(n467), .B(n484), .ZN(n1250) );
  CLKBUF_X1 U1082 ( .A(n28), .Z(n1413) );
  CLKBUF_X3 U1083 ( .A(n49), .Z(n1402) );
  INV_X1 U1084 ( .A(n641), .ZN(n1251) );
  CLKBUF_X3 U1085 ( .A(n58), .Z(n1503) );
  NAND2_X1 U1086 ( .A1(n1302), .A2(n1410), .ZN(n1335) );
  CLKBUF_X3 U1087 ( .A(n1099), .Z(n1538) );
  CLKBUF_X3 U1088 ( .A(n40), .Z(n1507) );
  BUF_X1 U1089 ( .A(n19), .Z(n1525) );
  CLKBUF_X2 U1090 ( .A(n19), .Z(n1337) );
  XNOR2_X1 U1091 ( .A(n1252), .B(n471), .ZN(n465) );
  XNOR2_X1 U1092 ( .A(n486), .B(n469), .ZN(n1252) );
  NAND2_X1 U1093 ( .A1(n446), .A2(n433), .ZN(n1253) );
  NAND2_X1 U1094 ( .A1(n446), .A2(n448), .ZN(n1254) );
  NAND2_X1 U1095 ( .A1(n433), .A2(n448), .ZN(n1255) );
  NAND3_X1 U1096 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n428) );
  CLKBUF_X2 U1097 ( .A(n1104), .Z(n1533) );
  BUF_X2 U1098 ( .A(n1108), .Z(n1256) );
  AOI21_X1 U1099 ( .B1(n1501), .B2(n247), .A(n244), .ZN(n242) );
  BUF_X1 U1100 ( .A(n1105), .Z(n1324) );
  NAND3_X1 U1101 ( .A1(n1475), .A2(n1476), .A3(n1477), .ZN(n1257) );
  OAI22_X1 U1102 ( .A1(n1379), .A2(n896), .B1(n895), .B2(n1503), .ZN(n1258) );
  XOR2_X1 U1103 ( .A(n417), .B(n432), .Z(n1259) );
  XOR2_X1 U1104 ( .A(n1243), .B(n1259), .Z(n413) );
  NAND2_X1 U1105 ( .A1(n430), .A2(n417), .ZN(n1260) );
  NAND2_X1 U1106 ( .A1(n430), .A2(n432), .ZN(n1261) );
  NAND2_X1 U1107 ( .A1(n417), .A2(n432), .ZN(n1262) );
  NAND3_X1 U1108 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n412) );
  CLKBUF_X1 U1109 ( .A(n176), .Z(n1263) );
  BUF_X1 U1110 ( .A(n42), .Z(n1375) );
  XOR2_X1 U1111 ( .A(n805), .B(n823), .Z(n1264) );
  XOR2_X1 U1112 ( .A(n1264), .B(n494), .Z(n471) );
  NAND2_X1 U1113 ( .A1(n805), .A2(n823), .ZN(n1265) );
  NAND2_X1 U1114 ( .A1(n805), .A2(n494), .ZN(n1266) );
  NAND2_X1 U1115 ( .A1(n823), .A2(n494), .ZN(n1267) );
  NAND3_X1 U1116 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n470) );
  NAND2_X1 U1117 ( .A1(n486), .A2(n469), .ZN(n1268) );
  NAND2_X1 U1118 ( .A1(n486), .A2(n471), .ZN(n1269) );
  NAND2_X1 U1119 ( .A1(n469), .A2(n471), .ZN(n1270) );
  NAND3_X1 U1120 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n464) );
  BUF_X1 U1121 ( .A(n46), .Z(n1508) );
  NAND2_X1 U1122 ( .A1(n1486), .A2(n46), .ZN(n1272) );
  NAND2_X1 U1123 ( .A1(n1486), .A2(n46), .ZN(n48) );
  BUF_X1 U1124 ( .A(n9), .Z(n1395) );
  BUF_X1 U1125 ( .A(n12), .Z(n1349) );
  BUF_X1 U1126 ( .A(n60), .Z(n1273) );
  CLKBUF_X1 U1127 ( .A(n1335), .Z(n1274) );
  BUF_X1 U1128 ( .A(n30), .Z(n1403) );
  BUF_X1 U1129 ( .A(n48), .Z(n1314) );
  CLKBUF_X2 U1130 ( .A(n25), .Z(n1451) );
  CLKBUF_X2 U1131 ( .A(n25), .Z(n1450) );
  CLKBUF_X1 U1132 ( .A(n1106), .Z(n1531) );
  INV_X1 U1133 ( .A(n193), .ZN(n1275) );
  OR2_X1 U1134 ( .A1(n150), .A2(n1481), .ZN(n1276) );
  CLKBUF_X1 U1135 ( .A(n1472), .Z(n1277) );
  CLKBUF_X1 U1136 ( .A(n16), .Z(n1415) );
  BUF_X2 U1137 ( .A(n1354), .Z(n1351) );
  BUF_X2 U1138 ( .A(n16), .Z(n1504) );
  XNOR2_X1 U1139 ( .A(n517), .B(n1278), .ZN(n1436) );
  AND3_X1 U1140 ( .A1(n1444), .A2(n1445), .A3(n1446), .ZN(n1278) );
  XOR2_X1 U1141 ( .A(n587), .B(n589), .Z(n1279) );
  XOR2_X1 U1142 ( .A(n1279), .B(n594), .Z(n583) );
  XOR2_X1 U1143 ( .A(n585), .B(n592), .Z(n1280) );
  XOR2_X1 U1144 ( .A(n1280), .B(n583), .Z(n581) );
  NAND2_X1 U1145 ( .A1(n587), .A2(n589), .ZN(n1281) );
  NAND2_X1 U1146 ( .A1(n587), .A2(n594), .ZN(n1282) );
  NAND2_X1 U1147 ( .A1(n589), .A2(n594), .ZN(n1283) );
  NAND3_X1 U1148 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n582) );
  NAND2_X1 U1149 ( .A1(n585), .A2(n592), .ZN(n1284) );
  NAND2_X1 U1150 ( .A1(n585), .A2(n583), .ZN(n1285) );
  NAND2_X1 U1151 ( .A1(n592), .A2(n583), .ZN(n1286) );
  NAND3_X1 U1152 ( .A1(n1284), .A2(n1285), .A3(n1286), .ZN(n580) );
  XNOR2_X1 U1153 ( .A(n1537), .B(n1352), .ZN(n1287) );
  CLKBUF_X3 U1154 ( .A(n36), .Z(n1394) );
  BUF_X2 U1155 ( .A(n36), .Z(n1393) );
  NOR2_X1 U1156 ( .A1(n1399), .A2(n209), .ZN(n1288) );
  XOR2_X1 U1157 ( .A(n570), .B(n561), .Z(n1289) );
  XOR2_X1 U1158 ( .A(n559), .B(n1289), .Z(n557) );
  NAND2_X1 U1159 ( .A1(n559), .A2(n570), .ZN(n1290) );
  NAND2_X1 U1160 ( .A1(n559), .A2(n561), .ZN(n1291) );
  NAND2_X1 U1161 ( .A1(n570), .A2(n561), .ZN(n1292) );
  NAND3_X1 U1162 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n556) );
  OR2_X2 U1163 ( .A1(n543), .A2(n556), .ZN(n1492) );
  XNOR2_X1 U1164 ( .A(n400), .B(n1293), .ZN(n385) );
  XNOR2_X1 U1165 ( .A(n402), .B(n389), .ZN(n1293) );
  CLKBUF_X1 U1166 ( .A(n148), .Z(n1294) );
  CLKBUF_X1 U1167 ( .A(n161), .Z(n1295) );
  NOR2_X1 U1168 ( .A1(n443), .A2(n460), .ZN(n161) );
  INV_X1 U1169 ( .A(n668), .ZN(n1296) );
  INV_X1 U1170 ( .A(n1528), .ZN(n1297) );
  INV_X1 U1171 ( .A(n1297), .ZN(n1298) );
  XNOR2_X1 U1172 ( .A(n1545), .B(n1383), .ZN(n1299) );
  CLKBUF_X1 U1173 ( .A(n1543), .Z(n1300) );
  CLKBUF_X3 U1174 ( .A(n1093), .Z(n1543) );
  XNOR2_X1 U1175 ( .A(n1436), .B(n1301), .ZN(n513) );
  XOR2_X1 U1176 ( .A(n1408), .B(n532), .Z(n1301) );
  CLKBUF_X3 U1177 ( .A(n31), .Z(n1323) );
  BUF_X2 U1178 ( .A(n40), .Z(n1506) );
  XOR2_X1 U1179 ( .A(n13), .B(a[4]), .Z(n1302) );
  XNOR2_X1 U1180 ( .A(n13), .B(a[6]), .ZN(n1303) );
  NAND3_X1 U1181 ( .A1(n1516), .A2(n1515), .A3(n1517), .ZN(n1304) );
  BUF_X2 U1182 ( .A(n1315), .Z(n1505) );
  XNOR2_X2 U1183 ( .A(n1526), .B(a[16]), .ZN(n1315) );
  BUF_X1 U1184 ( .A(n1098), .Z(n1306) );
  CLKBUF_X1 U1185 ( .A(n1383), .Z(n1307) );
  CLKBUF_X1 U1186 ( .A(n212), .Z(n1308) );
  BUF_X2 U1187 ( .A(n46), .Z(n1309) );
  BUF_X1 U1188 ( .A(n1107), .Z(n1312) );
  BUF_X2 U1189 ( .A(n1107), .Z(n1313) );
  CLKBUF_X1 U1190 ( .A(n1107), .Z(n1530) );
  AOI21_X1 U1191 ( .B1(n175), .B2(n1275), .A(n1263), .ZN(n1316) );
  XOR2_X1 U1192 ( .A(n37), .B(a[12]), .Z(n1487) );
  XNOR2_X1 U1193 ( .A(n1408), .B(n532), .ZN(n1317) );
  NOR2_X1 U1194 ( .A1(n371), .A2(n382), .ZN(n1318) );
  XNOR2_X1 U1195 ( .A(n1546), .B(n1305), .ZN(n1320) );
  XNOR2_X1 U1196 ( .A(n1358), .B(n1525), .ZN(n1321) );
  BUF_X2 U1197 ( .A(n1106), .Z(n1358) );
  XNOR2_X1 U1198 ( .A(n1), .B(n1296), .ZN(n1119) );
  NAND2_X1 U1199 ( .A1(n40), .A2(n1487), .ZN(n1472) );
  CLKBUF_X3 U1200 ( .A(n31), .Z(n1322) );
  BUF_X1 U1201 ( .A(n1233), .Z(n1325) );
  BUF_X2 U1202 ( .A(n61), .Z(n1528) );
  CLKBUF_X1 U1203 ( .A(n1309), .Z(n1326) );
  CLKBUF_X1 U1204 ( .A(n1542), .Z(n1327) );
  CLKBUF_X3 U1205 ( .A(n37), .Z(n1328) );
  CLKBUF_X1 U1206 ( .A(n221), .Z(n1329) );
  CLKBUF_X1 U1207 ( .A(n1541), .Z(n1330) );
  BUF_X2 U1208 ( .A(n4), .Z(n1332) );
  INV_X1 U1209 ( .A(n668), .ZN(n4) );
  CLKBUF_X1 U1210 ( .A(n162), .Z(n1333) );
  CLKBUF_X1 U1211 ( .A(n1453), .Z(n1334) );
  NAND2_X1 U1212 ( .A1(n1302), .A2(n1410), .ZN(n18) );
  CLKBUF_X2 U1213 ( .A(n19), .Z(n1336) );
  INV_X1 U1214 ( .A(n1314), .ZN(n1338) );
  INV_X1 U1215 ( .A(n1338), .ZN(n1339) );
  BUF_X1 U1216 ( .A(n1103), .Z(n1341) );
  BUF_X1 U1217 ( .A(n1103), .Z(n1342) );
  NAND2_X1 U1218 ( .A1(n1116), .A2(n1303), .ZN(n1343) );
  NAND2_X1 U1219 ( .A1(n1116), .A2(n1303), .ZN(n1412) );
  XNOR2_X1 U1220 ( .A(n1344), .B(n463), .ZN(n461) );
  XNOR2_X1 U1221 ( .A(n480), .B(n465), .ZN(n1344) );
  NOR2_X1 U1222 ( .A1(n581), .A2(n590), .ZN(n1345) );
  BUF_X1 U1223 ( .A(n1101), .Z(n1346) );
  BUF_X1 U1224 ( .A(n1101), .Z(n1347) );
  BUF_X2 U1225 ( .A(n1511), .Z(n1356) );
  AOI21_X1 U1226 ( .B1(n1381), .B2(n133), .A(n134), .ZN(n1348) );
  BUF_X2 U1227 ( .A(n1354), .Z(n1350) );
  CLKBUF_X1 U1228 ( .A(n1339), .Z(n1353) );
  XNOR2_X1 U1229 ( .A(n25), .B(a[10]), .ZN(n1354) );
  CLKBUF_X3 U1230 ( .A(n1096), .Z(n1540) );
  NAND2_X1 U1231 ( .A1(n1382), .A2(n1332), .ZN(n1355) );
  AOI21_X1 U1232 ( .B1(n221), .B2(n213), .A(n214), .ZN(n212) );
  CLKBUF_X1 U1233 ( .A(n1544), .Z(n1360) );
  BUF_X1 U1234 ( .A(n6), .Z(n1361) );
  BUF_X2 U1235 ( .A(n6), .Z(n1362) );
  CLKBUF_X1 U1236 ( .A(n12), .Z(n1363) );
  NAND2_X1 U1237 ( .A1(n1485), .A2(n9), .ZN(n12) );
  CLKBUF_X1 U1238 ( .A(n1546), .Z(n1365) );
  BUF_X2 U1239 ( .A(n1090), .Z(n1546) );
  AOI21_X1 U1240 ( .B1(n1493), .B2(n1416), .A(n183), .ZN(n1366) );
  CLKBUF_X3 U1241 ( .A(n55), .Z(n1367) );
  CLKBUF_X3 U1242 ( .A(n55), .Z(n1368) );
  CLKBUF_X1 U1243 ( .A(n1389), .Z(n1369) );
  CLKBUF_X1 U1244 ( .A(n1277), .Z(n1370) );
  XNOR2_X1 U1245 ( .A(n1371), .B(n535), .ZN(n531) );
  XNOR2_X1 U1246 ( .A(n546), .B(n548), .ZN(n1371) );
  OR2_X1 U1247 ( .A1(n195), .A2(n212), .ZN(n1372) );
  NAND2_X1 U1248 ( .A1(n1372), .A2(n196), .ZN(n194) );
  NAND2_X1 U1249 ( .A1(n1491), .A2(n58), .ZN(n60) );
  CLKBUF_X1 U1250 ( .A(n1452), .Z(n1373) );
  BUF_X1 U1251 ( .A(n42), .Z(n1374) );
  CLKBUF_X1 U1252 ( .A(n127), .Z(n1376) );
  CLKBUF_X1 U1253 ( .A(n264), .Z(n1377) );
  INV_X1 U1254 ( .A(n60), .ZN(n1378) );
  INV_X2 U1255 ( .A(n1378), .ZN(n1379) );
  INV_X1 U1256 ( .A(n1378), .ZN(n1380) );
  CLKBUF_X1 U1257 ( .A(n146), .Z(n1381) );
  XOR2_X1 U1258 ( .A(n1), .B(n668), .Z(n1382) );
  NAND3_X1 U1259 ( .A1(n1388), .A2(n1389), .A3(n1390), .ZN(n1384) );
  NAND3_X1 U1260 ( .A1(n1388), .A2(n1369), .A3(n1390), .ZN(n1385) );
  AOI21_X1 U1261 ( .B1(n1522), .B2(n126), .A(n1376), .ZN(n1386) );
  AOI21_X1 U1262 ( .B1(n153), .B2(n126), .A(n127), .ZN(n125) );
  NAND2_X1 U1263 ( .A1(n1382), .A2(n1332), .ZN(n1454) );
  NAND2_X1 U1264 ( .A1(n1119), .A2(n4), .ZN(n6) );
  NAND2_X1 U1265 ( .A1(n1487), .A2(n40), .ZN(n42) );
  XOR2_X1 U1266 ( .A(n310), .B(n307), .Z(n1387) );
  XOR2_X1 U1267 ( .A(n1377), .B(n1387), .Z(product[34]) );
  NAND2_X1 U1268 ( .A1(n264), .A2(n310), .ZN(n1388) );
  NAND2_X1 U1269 ( .A1(n264), .A2(n307), .ZN(n1389) );
  NAND2_X1 U1270 ( .A1(n310), .A2(n307), .ZN(n1390) );
  NAND3_X1 U1271 ( .A1(n1388), .A2(n1389), .A3(n1390), .ZN(n100) );
  CLKBUF_X1 U1272 ( .A(n106), .Z(n1391) );
  CLKBUF_X1 U1273 ( .A(n114), .Z(n1392) );
  NAND2_X1 U1274 ( .A1(n1489), .A2(n34), .ZN(n36) );
  NAND2_X1 U1275 ( .A1(n400), .A2(n402), .ZN(n1396) );
  NAND2_X1 U1276 ( .A1(n400), .A2(n389), .ZN(n1397) );
  NAND2_X1 U1277 ( .A1(n402), .A2(n389), .ZN(n1398) );
  NAND3_X1 U1278 ( .A1(n1396), .A2(n1397), .A3(n1398), .ZN(n384) );
  NOR2_X1 U1279 ( .A1(n557), .A2(n568), .ZN(n1399) );
  NOR2_X1 U1280 ( .A1(n557), .A2(n568), .ZN(n204) );
  NAND3_X1 U1281 ( .A1(n1444), .A2(n1445), .A3(n1446), .ZN(n1400) );
  NAND2_X1 U1282 ( .A1(n1488), .A2(n28), .ZN(n30) );
  CLKBUF_X1 U1283 ( .A(n840), .Z(n1407) );
  XNOR2_X1 U1284 ( .A(n519), .B(n521), .ZN(n1408) );
  XNOR2_X1 U1285 ( .A(n7), .B(a[4]), .ZN(n1410) );
  XNOR2_X1 U1286 ( .A(n1411), .B(n500), .ZN(n481) );
  XNOR2_X1 U1287 ( .A(n485), .B(n487), .ZN(n1411) );
  XOR2_X1 U1288 ( .A(n514), .B(n501), .Z(n1417) );
  XOR2_X1 U1289 ( .A(n499), .B(n1417), .Z(n497) );
  NAND2_X1 U1290 ( .A1(n499), .A2(n514), .ZN(n1418) );
  NAND2_X1 U1291 ( .A1(n499), .A2(n501), .ZN(n1419) );
  NAND2_X1 U1292 ( .A1(n514), .A2(n501), .ZN(n1420) );
  NAND3_X1 U1293 ( .A1(n1418), .A2(n1419), .A3(n1420), .ZN(n496) );
  XNOR2_X1 U1294 ( .A(n37), .B(a[14]), .ZN(n46) );
  XNOR2_X1 U1295 ( .A(n429), .B(n1421), .ZN(n427) );
  XNOR2_X1 U1296 ( .A(n444), .B(n431), .ZN(n1421) );
  XNOR2_X1 U1297 ( .A(n1422), .B(n413), .ZN(n411) );
  XNOR2_X1 U1298 ( .A(n428), .B(n415), .ZN(n1422) );
  XOR2_X1 U1299 ( .A(n520), .B(n509), .Z(n1423) );
  XOR2_X1 U1300 ( .A(n1423), .B(n518), .Z(n501) );
  NAND2_X1 U1301 ( .A1(n520), .A2(n509), .ZN(n1424) );
  NAND2_X1 U1302 ( .A1(n520), .A2(n518), .ZN(n1425) );
  NAND2_X1 U1303 ( .A1(n509), .A2(n518), .ZN(n1426) );
  NAND3_X1 U1304 ( .A1(n1424), .A2(n1425), .A3(n1426), .ZN(n500) );
  NAND2_X1 U1305 ( .A1(n487), .A2(n485), .ZN(n1427) );
  NAND2_X1 U1306 ( .A1(n487), .A2(n500), .ZN(n1428) );
  NAND2_X1 U1307 ( .A1(n485), .A2(n500), .ZN(n1429) );
  NAND3_X1 U1308 ( .A1(n1427), .A2(n1428), .A3(n1429), .ZN(n480) );
  CLKBUF_X2 U1309 ( .A(n43), .Z(n1430) );
  NAND2_X1 U1310 ( .A1(n413), .A2(n1249), .ZN(n1432) );
  NAND2_X1 U1311 ( .A1(n413), .A2(n415), .ZN(n1433) );
  NAND2_X1 U1312 ( .A1(n1249), .A2(n415), .ZN(n1434) );
  NAND3_X1 U1313 ( .A1(n1432), .A2(n1433), .A3(n1434), .ZN(n410) );
  CLKBUF_X1 U1314 ( .A(n151), .Z(n1435) );
  NAND2_X1 U1315 ( .A1(n519), .A2(n521), .ZN(n1437) );
  NAND2_X1 U1316 ( .A1(n519), .A2(n532), .ZN(n1438) );
  NAND2_X1 U1317 ( .A1(n521), .A2(n532), .ZN(n1439) );
  NAND3_X1 U1318 ( .A1(n1437), .A2(n1438), .A3(n1439), .ZN(n514) );
  NAND2_X1 U1319 ( .A1(n517), .A2(n1400), .ZN(n1440) );
  NAND2_X1 U1320 ( .A1(n517), .A2(n1317), .ZN(n1441) );
  NAND2_X1 U1321 ( .A1(n1400), .A2(n1317), .ZN(n1442) );
  NAND3_X1 U1322 ( .A1(n1440), .A2(n1441), .A3(n1442), .ZN(n512) );
  XOR2_X1 U1323 ( .A(n544), .B(n533), .Z(n1443) );
  XOR2_X1 U1324 ( .A(n531), .B(n1443), .Z(n529) );
  NAND2_X1 U1325 ( .A1(n546), .A2(n548), .ZN(n1444) );
  NAND2_X1 U1326 ( .A1(n546), .A2(n535), .ZN(n1445) );
  NAND2_X1 U1327 ( .A1(n548), .A2(n535), .ZN(n1446) );
  NAND2_X1 U1328 ( .A1(n544), .A2(n533), .ZN(n1447) );
  NAND2_X1 U1329 ( .A1(n531), .A2(n544), .ZN(n1448) );
  NAND2_X1 U1330 ( .A1(n531), .A2(n533), .ZN(n1449) );
  NAND3_X1 U1331 ( .A1(n1447), .A2(n1448), .A3(n1449), .ZN(n528) );
  NAND3_X1 U1332 ( .A1(n1457), .A2(n1458), .A3(n1456), .ZN(n1452) );
  NAND3_X1 U1333 ( .A1(n1461), .A2(n1462), .A3(n1460), .ZN(n1453) );
  XOR2_X1 U1334 ( .A(n303), .B(n306), .Z(n1455) );
  XOR2_X1 U1335 ( .A(n1455), .B(n1385), .Z(product[35]) );
  NAND2_X1 U1336 ( .A1(n303), .A2(n306), .ZN(n1456) );
  NAND2_X1 U1337 ( .A1(n303), .A2(n1384), .ZN(n1457) );
  NAND2_X1 U1338 ( .A1(n100), .A2(n306), .ZN(n1458) );
  NAND3_X1 U1339 ( .A1(n1458), .A2(n1457), .A3(n1456), .ZN(n99) );
  XOR2_X1 U1340 ( .A(n302), .B(n301), .Z(n1459) );
  XOR2_X1 U1341 ( .A(n1373), .B(n1459), .Z(product[36]) );
  NAND2_X1 U1342 ( .A1(n302), .A2(n301), .ZN(n1460) );
  NAND2_X1 U1343 ( .A1(n1452), .A2(n302), .ZN(n1461) );
  NAND2_X1 U1344 ( .A1(n301), .A2(n99), .ZN(n1462) );
  NAND3_X1 U1345 ( .A1(n1461), .A2(n1460), .A3(n1462), .ZN(n98) );
  NAND2_X1 U1346 ( .A1(n467), .A2(n484), .ZN(n1463) );
  NAND2_X1 U1347 ( .A1(n467), .A2(n482), .ZN(n1464) );
  NAND2_X1 U1348 ( .A1(n484), .A2(n482), .ZN(n1465) );
  NAND3_X1 U1349 ( .A1(n1463), .A2(n1464), .A3(n1465), .ZN(n462) );
  NAND2_X1 U1350 ( .A1(n480), .A2(n465), .ZN(n1466) );
  NAND2_X1 U1351 ( .A1(n480), .A2(n463), .ZN(n1467) );
  NAND2_X1 U1352 ( .A1(n465), .A2(n463), .ZN(n1468) );
  NAND3_X1 U1353 ( .A1(n1466), .A2(n1467), .A3(n1468), .ZN(n460) );
  NAND2_X1 U1354 ( .A1(n429), .A2(n444), .ZN(n1469) );
  NAND2_X1 U1355 ( .A1(n429), .A2(n431), .ZN(n1470) );
  NAND2_X1 U1356 ( .A1(n444), .A2(n431), .ZN(n1471) );
  NAND3_X1 U1357 ( .A1(n1469), .A2(n1470), .A3(n1471), .ZN(n426) );
  NOR2_X1 U1358 ( .A1(n427), .A2(n442), .ZN(n1473) );
  NOR2_X1 U1359 ( .A1(n427), .A2(n442), .ZN(n158) );
  XOR2_X1 U1360 ( .A(n821), .B(n1258), .Z(n1474) );
  XOR2_X1 U1361 ( .A(n1474), .B(n1407), .Z(n441) );
  NAND2_X1 U1362 ( .A1(n821), .A2(n695), .ZN(n1475) );
  NAND2_X1 U1363 ( .A1(n821), .A2(n840), .ZN(n1476) );
  NAND2_X1 U1364 ( .A1(n695), .A2(n840), .ZN(n1477) );
  NAND2_X1 U1365 ( .A1(n425), .A2(n748), .ZN(n1478) );
  NAND2_X1 U1366 ( .A1(n425), .A2(n1257), .ZN(n1479) );
  NAND2_X1 U1367 ( .A1(n748), .A2(n1257), .ZN(n1480) );
  NAND3_X1 U1368 ( .A1(n1480), .A2(n1479), .A3(n1478), .ZN(n418) );
  NOR2_X1 U1369 ( .A1(n410), .A2(n397), .ZN(n1481) );
  NOR2_X1 U1370 ( .A1(n397), .A2(n410), .ZN(n147) );
  NOR2_X2 U1371 ( .A1(n461), .A2(n478), .ZN(n166) );
  AOI21_X1 U1372 ( .B1(n114), .B2(n1497), .A(n111), .ZN(n1482) );
  NOR2_X1 U1373 ( .A1(n497), .A2(n512), .ZN(n1483) );
  NOR2_X1 U1374 ( .A1(n497), .A2(n512), .ZN(n177) );
  OR2_X1 U1375 ( .A1(n513), .A2(n528), .ZN(n1493) );
  NOR2_X1 U1376 ( .A1(n581), .A2(n590), .ZN(n215) );
  NOR2_X1 U1377 ( .A1(n591), .A2(n600), .ZN(n218) );
  NOR2_X1 U1378 ( .A1(n349), .A2(n358), .ZN(n123) );
  NAND2_X1 U1379 ( .A1(n591), .A2(n600), .ZN(n219) );
  NAND2_X1 U1380 ( .A1(n581), .A2(n590), .ZN(n216) );
  OR2_X1 U1381 ( .A1(n617), .A2(n622), .ZN(n1484) );
  OR2_X1 U1382 ( .A1(n339), .A2(n348), .ZN(n1496) );
  OR2_X1 U1383 ( .A1(n609), .A2(n616), .ZN(n1494) );
  BUF_X2 U1384 ( .A(n1105), .Z(n1532) );
  XOR2_X1 U1385 ( .A(n7), .B(a[2]), .Z(n1485) );
  XOR2_X1 U1386 ( .A(n1526), .B(a[14]), .Z(n1486) );
  XOR2_X1 U1387 ( .A(n25), .B(a[8]), .Z(n1488) );
  XOR2_X1 U1388 ( .A(n31), .B(a[10]), .Z(n1489) );
  XOR2_X1 U1389 ( .A(n49), .B(a[16]), .Z(n1490) );
  XOR2_X1 U1390 ( .A(n55), .B(a[18]), .Z(n1491) );
  OAI21_X1 U1391 ( .B1(n152), .B2(n1276), .A(n144), .ZN(n142) );
  INV_X1 U1392 ( .A(n1381), .ZN(n144) );
  NOR2_X1 U1393 ( .A1(n1483), .A2(n180), .ZN(n175) );
  INV_X1 U1394 ( .A(n200), .ZN(n198) );
  NOR2_X1 U1395 ( .A1(n131), .A2(n128), .ZN(n126) );
  INV_X1 U1396 ( .A(n1308), .ZN(n211) );
  AOI21_X1 U1397 ( .B1(n1493), .B2(n1416), .A(n183), .ZN(n181) );
  INV_X1 U1398 ( .A(n185), .ZN(n183) );
  INV_X1 U1399 ( .A(n171), .ZN(n279) );
  XOR2_X1 U1400 ( .A(n168), .B(n76), .Z(product[20]) );
  NAND2_X1 U1401 ( .A1(n278), .A2(n167), .ZN(n76) );
  AOI21_X1 U1402 ( .B1(n173), .B2(n279), .A(n170), .ZN(n168) );
  XOR2_X1 U1403 ( .A(n137), .B(n70), .Z(product[26]) );
  NAND2_X1 U1404 ( .A1(n272), .A2(n136), .ZN(n70) );
  AOI21_X1 U1405 ( .B1(n142), .B2(n273), .A(n139), .ZN(n137) );
  INV_X1 U1406 ( .A(n1318), .ZN(n272) );
  XOR2_X1 U1407 ( .A(n206), .B(n82), .Z(product[14]) );
  NAND2_X1 U1408 ( .A1(n1237), .A2(n205), .ZN(n82) );
  AOI21_X1 U1409 ( .B1(n211), .B2(n285), .A(n208), .ZN(n206) );
  XOR2_X1 U1410 ( .A(n201), .B(n81), .Z(product[15]) );
  NAND2_X1 U1411 ( .A1(n1492), .A2(n200), .ZN(n81) );
  AOI21_X1 U1412 ( .B1(n211), .B2(n1288), .A(n203), .ZN(n201) );
  XOR2_X1 U1413 ( .A(n163), .B(n75), .Z(product[21]) );
  NAND2_X1 U1414 ( .A1(n277), .A2(n1333), .ZN(n75) );
  XOR2_X1 U1415 ( .A(n152), .B(n73), .Z(product[23]) );
  NAND2_X1 U1416 ( .A1(n275), .A2(n1435), .ZN(n73) );
  XOR2_X1 U1417 ( .A(n193), .B(n80), .Z(product[16]) );
  NAND2_X1 U1418 ( .A1(n282), .A2(n188), .ZN(n80) );
  INV_X1 U1419 ( .A(n1329), .ZN(n220) );
  NAND2_X1 U1420 ( .A1(n1493), .A2(n282), .ZN(n180) );
  XNOR2_X1 U1421 ( .A(n160), .B(n74), .ZN(product[22]) );
  NAND2_X1 U1422 ( .A1(n1238), .A2(n159), .ZN(n74) );
  XNOR2_X1 U1423 ( .A(n173), .B(n77), .ZN(product[19]) );
  NAND2_X1 U1424 ( .A1(n279), .A2(n172), .ZN(n77) );
  XNOR2_X1 U1425 ( .A(n149), .B(n72), .ZN(product[24]) );
  NAND2_X1 U1426 ( .A1(n274), .A2(n1294), .ZN(n72) );
  INV_X1 U1427 ( .A(n1481), .ZN(n274) );
  XNOR2_X1 U1428 ( .A(n130), .B(n69), .ZN(product[27]) );
  NAND2_X1 U1429 ( .A1(n271), .A2(n129), .ZN(n69) );
  INV_X1 U1430 ( .A(n128), .ZN(n271) );
  XNOR2_X1 U1431 ( .A(n186), .B(n79), .ZN(product[17]) );
  XNOR2_X1 U1432 ( .A(n142), .B(n71), .ZN(product[25]) );
  NAND2_X1 U1433 ( .A1(n273), .A2(n141), .ZN(n71) );
  XNOR2_X1 U1434 ( .A(n179), .B(n78), .ZN(product[18]) );
  NAND2_X1 U1435 ( .A1(n280), .A2(n178), .ZN(n78) );
  INV_X1 U1436 ( .A(n177), .ZN(n280) );
  INV_X1 U1437 ( .A(n172), .ZN(n170) );
  INV_X1 U1438 ( .A(n141), .ZN(n139) );
  NOR2_X1 U1439 ( .A1(n1345), .A2(n218), .ZN(n213) );
  OAI21_X1 U1440 ( .B1(n215), .B2(n219), .A(n216), .ZN(n214) );
  INV_X1 U1441 ( .A(n113), .ZN(n111) );
  INV_X1 U1442 ( .A(n238), .ZN(n236) );
  NOR2_X1 U1443 ( .A1(n371), .A2(n382), .ZN(n135) );
  NOR2_X1 U1444 ( .A1(n359), .A2(n370), .ZN(n128) );
  NAND2_X1 U1445 ( .A1(n270), .A2(n124), .ZN(n68) );
  INV_X1 U1446 ( .A(n123), .ZN(n270) );
  NAND2_X1 U1447 ( .A1(n268), .A2(n116), .ZN(n66) );
  INV_X1 U1448 ( .A(n115), .ZN(n268) );
  NAND2_X1 U1449 ( .A1(n266), .A2(n108), .ZN(n64) );
  INV_X1 U1450 ( .A(n107), .ZN(n266) );
  INV_X1 U1451 ( .A(n209), .ZN(n285) );
  NAND2_X1 U1452 ( .A1(n411), .A2(n426), .ZN(n151) );
  NAND2_X1 U1453 ( .A1(n1498), .A2(n105), .ZN(n63) );
  NAND2_X1 U1454 ( .A1(n1496), .A2(n121), .ZN(n67) );
  NAND2_X1 U1455 ( .A1(n1497), .A2(n113), .ZN(n65) );
  XOR2_X1 U1456 ( .A(n220), .B(n85), .Z(product[11]) );
  NAND2_X1 U1457 ( .A1(n287), .A2(n219), .ZN(n85) );
  INV_X1 U1458 ( .A(n218), .ZN(n287) );
  XOR2_X1 U1459 ( .A(n228), .B(n86), .Z(product[10]) );
  NAND2_X1 U1460 ( .A1(n1495), .A2(n227), .ZN(n86) );
  AOI21_X1 U1461 ( .B1(n233), .B2(n1494), .A(n230), .ZN(n228) );
  NOR2_X1 U1462 ( .A1(n479), .A2(n496), .ZN(n171) );
  NAND2_X1 U1463 ( .A1(n479), .A2(n496), .ZN(n172) );
  XNOR2_X1 U1464 ( .A(n239), .B(n88), .ZN(product[8]) );
  NAND2_X1 U1465 ( .A1(n1484), .A2(n238), .ZN(n88) );
  XNOR2_X1 U1466 ( .A(n211), .B(n83), .ZN(product[13]) );
  NAND2_X1 U1467 ( .A1(n285), .A2(n210), .ZN(n83) );
  XNOR2_X1 U1468 ( .A(n233), .B(n87), .ZN(product[9]) );
  NAND2_X1 U1469 ( .A1(n1494), .A2(n232), .ZN(n87) );
  XNOR2_X1 U1470 ( .A(n217), .B(n84), .ZN(product[12]) );
  NAND2_X1 U1471 ( .A1(n286), .A2(n216), .ZN(n84) );
  OAI21_X1 U1472 ( .B1(n220), .B2(n218), .A(n219), .ZN(n217) );
  INV_X1 U1473 ( .A(n1345), .ZN(n286) );
  NAND2_X1 U1474 ( .A1(n383), .A2(n396), .ZN(n141) );
  NAND2_X1 U1475 ( .A1(n497), .A2(n512), .ZN(n178) );
  NAND2_X1 U1476 ( .A1(n397), .A2(n410), .ZN(n148) );
  NAND2_X1 U1477 ( .A1(n359), .A2(n370), .ZN(n129) );
  NAND2_X1 U1478 ( .A1(n443), .A2(n460), .ZN(n162) );
  NAND2_X1 U1479 ( .A1(n543), .A2(n556), .ZN(n200) );
  INV_X1 U1480 ( .A(n232), .ZN(n230) );
  NAND2_X1 U1481 ( .A1(n371), .A2(n382), .ZN(n136) );
  INV_X1 U1482 ( .A(n210), .ZN(n208) );
  INV_X1 U1483 ( .A(n121), .ZN(n119) );
  NAND2_X1 U1484 ( .A1(n1495), .A2(n1494), .ZN(n222) );
  INV_X1 U1485 ( .A(n246), .ZN(n244) );
  AOI21_X1 U1486 ( .B1(n1499), .B2(n255), .A(n252), .ZN(n250) );
  INV_X1 U1487 ( .A(n254), .ZN(n252) );
  OAI21_X1 U1488 ( .B1(n256), .B2(n258), .A(n257), .ZN(n255) );
  OR2_X2 U1489 ( .A1(n601), .A2(n608), .ZN(n1495) );
  NAND2_X1 U1490 ( .A1(n291), .A2(n241), .ZN(n89) );
  INV_X1 U1491 ( .A(n240), .ZN(n291) );
  OAI21_X1 U1492 ( .B1(n248), .B2(n250), .A(n249), .ZN(n247) );
  XOR2_X1 U1493 ( .A(n91), .B(n1236), .Z(product[5]) );
  NAND2_X1 U1494 ( .A1(n293), .A2(n249), .ZN(n91) );
  INV_X1 U1495 ( .A(n248), .ZN(n293) );
  NOR2_X1 U1496 ( .A1(n569), .A2(n580), .ZN(n209) );
  NOR2_X1 U1497 ( .A1(n317), .A2(n322), .ZN(n107) );
  NOR2_X1 U1498 ( .A1(n331), .A2(n338), .ZN(n115) );
  INV_X1 U1499 ( .A(n259), .ZN(n258) );
  OAI21_X1 U1500 ( .B1(n260), .B2(n263), .A(n261), .ZN(n259) );
  NAND2_X1 U1501 ( .A1(n569), .A2(n580), .ZN(n210) );
  NAND2_X1 U1502 ( .A1(n349), .A2(n358), .ZN(n124) );
  XNOR2_X1 U1503 ( .A(n92), .B(n255), .ZN(product[4]) );
  NAND2_X1 U1504 ( .A1(n1499), .A2(n254), .ZN(n92) );
  XNOR2_X1 U1505 ( .A(n90), .B(n247), .ZN(product[6]) );
  NAND2_X1 U1506 ( .A1(n1501), .A2(n246), .ZN(n90) );
  NAND2_X1 U1507 ( .A1(n609), .A2(n616), .ZN(n232) );
  NAND2_X1 U1508 ( .A1(n323), .A2(n330), .ZN(n113) );
  NAND2_X1 U1509 ( .A1(n339), .A2(n348), .ZN(n121) );
  NAND2_X1 U1510 ( .A1(n617), .A2(n622), .ZN(n238) );
  NAND2_X1 U1511 ( .A1(n311), .A2(n316), .ZN(n105) );
  NAND2_X1 U1512 ( .A1(n317), .A2(n322), .ZN(n108) );
  NAND2_X1 U1513 ( .A1(n331), .A2(n338), .ZN(n116) );
  OR2_X1 U1514 ( .A1(n323), .A2(n330), .ZN(n1497) );
  OR2_X1 U1515 ( .A1(n311), .A2(n316), .ZN(n1498) );
  XOR2_X1 U1516 ( .A(n93), .B(n258), .Z(product[3]) );
  NAND2_X1 U1517 ( .A1(n295), .A2(n257), .ZN(n93) );
  INV_X1 U1518 ( .A(n256), .ZN(n295) );
  XOR2_X1 U1519 ( .A(n94), .B(n263), .Z(product[2]) );
  NAND2_X1 U1520 ( .A1(n296), .A2(n261), .ZN(n94) );
  INV_X1 U1521 ( .A(n260), .ZN(n296) );
  NAND2_X1 U1522 ( .A1(n639), .A2(n678), .ZN(n257) );
  NOR2_X1 U1523 ( .A1(n639), .A2(n678), .ZN(n256) );
  NOR2_X1 U1524 ( .A1(n633), .A2(n636), .ZN(n248) );
  NOR2_X1 U1525 ( .A1(n878), .A2(n859), .ZN(n260) );
  NAND2_X1 U1526 ( .A1(n679), .A2(n879), .ZN(n263) );
  NAND2_X1 U1527 ( .A1(n878), .A2(n859), .ZN(n261) );
  INV_X1 U1528 ( .A(n298), .ZN(n299) );
  OR2_X1 U1529 ( .A1(n637), .A2(n638), .ZN(n1499) );
  INV_X1 U1530 ( .A(n328), .ZN(n329) );
  INV_X1 U1531 ( .A(n394), .ZN(n395) );
  NOR2_X1 U1532 ( .A1(n623), .A2(n628), .ZN(n240) );
  NAND2_X1 U1533 ( .A1(n633), .A2(n636), .ZN(n249) );
  INV_X1 U1534 ( .A(n105), .ZN(n103) );
  NAND2_X1 U1535 ( .A1(n629), .A2(n632), .ZN(n246) );
  XNOR2_X1 U1536 ( .A(n1500), .B(n1512), .ZN(product[38]) );
  XNOR2_X1 U1537 ( .A(n680), .B(n298), .ZN(n1500) );
  NAND2_X1 U1538 ( .A1(n623), .A2(n628), .ZN(n241) );
  NAND2_X1 U1539 ( .A1(n637), .A2(n638), .ZN(n254) );
  OR2_X1 U1540 ( .A1(n629), .A2(n632), .ZN(n1501) );
  AND3_X1 U1541 ( .A1(n1520), .A2(n1519), .A3(n1518), .ZN(product[39]) );
  OR2_X1 U1542 ( .A1(n1298), .A2(n1148), .ZN(n1068) );
  OAI22_X1 U1543 ( .A1(n1362), .A2(n1086), .B1(n1085), .B2(n1332), .ZN(n877)
         );
  OAI22_X1 U1544 ( .A1(n1454), .A2(n1088), .B1(n1087), .B2(n1331), .ZN(n879)
         );
  OAI22_X1 U1545 ( .A1(n1355), .A2(n1149), .B1(n1089), .B2(n1332), .ZN(n679)
         );
  OR2_X1 U1546 ( .A1(n1528), .A2(n1149), .ZN(n1089) );
  OAI22_X1 U1547 ( .A1(n1362), .A2(n1087), .B1(n1086), .B2(n1331), .ZN(n878)
         );
  OAI22_X1 U1548 ( .A1(n1362), .A2(n1081), .B1(n1080), .B2(n1331), .ZN(n872)
         );
  AND2_X1 U1549 ( .A1(n1298), .A2(n656), .ZN(n799) );
  XNOR2_X1 U1550 ( .A(n1527), .B(n1402), .ZN(n920) );
  OAI22_X1 U1551 ( .A1(n1362), .A2(n1074), .B1(n1073), .B2(n1331), .ZN(n865)
         );
  XNOR2_X1 U1552 ( .A(n1527), .B(n1450), .ZN(n1004) );
  OAI22_X1 U1553 ( .A1(n1454), .A2(n1084), .B1(n1083), .B2(n1332), .ZN(n875)
         );
  XNOR2_X1 U1554 ( .A(n1527), .B(n1340), .ZN(n1046) );
  OAI22_X1 U1555 ( .A1(n1069), .A2(n1361), .B1(n1069), .B2(n1332), .ZN(n667)
         );
  OAI22_X1 U1556 ( .A1(n1355), .A2(n1082), .B1(n1081), .B2(n1332), .ZN(n873)
         );
  OAI22_X1 U1557 ( .A1(n1362), .A2(n1072), .B1(n1071), .B2(n1332), .ZN(n863)
         );
  OR2_X1 U1558 ( .A1(n1298), .A2(n1147), .ZN(n1047) );
  AND2_X1 U1559 ( .A1(n1298), .A2(n662), .ZN(n839) );
  OAI22_X1 U1560 ( .A1(n1362), .A2(n1085), .B1(n1084), .B2(n1332), .ZN(n876)
         );
  XNOR2_X1 U1561 ( .A(n1528), .B(n1431), .ZN(n941) );
  XNOR2_X1 U1562 ( .A(n1546), .B(n1524), .ZN(n1027) );
  XNOR2_X1 U1563 ( .A(n1365), .B(n1328), .ZN(n943) );
  XNOR2_X1 U1564 ( .A(n1365), .B(n1401), .ZN(n901) );
  XNOR2_X1 U1565 ( .A(n1365), .B(n1431), .ZN(n922) );
  XNOR2_X1 U1566 ( .A(n1365), .B(n1450), .ZN(n985) );
  BUF_X1 U1567 ( .A(n1101), .Z(n1536) );
  BUF_X1 U1568 ( .A(n1103), .Z(n1534) );
  BUF_X1 U1569 ( .A(n1098), .Z(n1539) );
  XNOR2_X1 U1570 ( .A(n1545), .B(n1352), .ZN(n944) );
  XNOR2_X1 U1571 ( .A(n1327), .B(n1431), .ZN(n926) );
  XNOR2_X1 U1572 ( .A(n1330), .B(n1402), .ZN(n906) );
  XNOR2_X1 U1573 ( .A(n1300), .B(n1430), .ZN(n925) );
  XNOR2_X1 U1574 ( .A(n1330), .B(n1431), .ZN(n927) );
  XNOR2_X1 U1575 ( .A(n1532), .B(n1524), .ZN(n1042) );
  XNOR2_X1 U1576 ( .A(n1360), .B(n1352), .ZN(n945) );
  XNOR2_X1 U1577 ( .A(n1300), .B(n1328), .ZN(n946) );
  XNOR2_X1 U1578 ( .A(n1310), .B(n1340), .ZN(n1034) );
  XNOR2_X1 U1579 ( .A(n1540), .B(n1401), .ZN(n907) );
  XNOR2_X1 U1580 ( .A(n1358), .B(n1340), .ZN(n1043) );
  XNOR2_X1 U1581 ( .A(n1533), .B(n1340), .ZN(n1041) );
  XNOR2_X1 U1582 ( .A(n1540), .B(n1340), .ZN(n1033) );
  XNOR2_X1 U1583 ( .A(n1324), .B(n1328), .ZN(n958) );
  XNOR2_X1 U1584 ( .A(n1359), .B(n1352), .ZN(n959) );
  XNOR2_X1 U1585 ( .A(n1539), .B(n1340), .ZN(n1035) );
  XNOR2_X1 U1586 ( .A(n1529), .B(n1430), .ZN(n940) );
  XNOR2_X1 U1587 ( .A(n1533), .B(n1352), .ZN(n957) );
  XNOR2_X1 U1588 ( .A(n1324), .B(n1401), .ZN(n916) );
  XNOR2_X1 U1589 ( .A(n1324), .B(n1431), .ZN(n937) );
  XNOR2_X1 U1590 ( .A(n1541), .B(n1524), .ZN(n1032) );
  XNOR2_X1 U1591 ( .A(n1359), .B(n1401), .ZN(n917) );
  XNOR2_X1 U1592 ( .A(n1535), .B(n1340), .ZN(n1039) );
  XNOR2_X1 U1593 ( .A(n1536), .B(n1340), .ZN(n1038) );
  XNOR2_X1 U1594 ( .A(n1543), .B(n1524), .ZN(n1030) );
  XNOR2_X1 U1595 ( .A(n1542), .B(n1340), .ZN(n1031) );
  XNOR2_X1 U1596 ( .A(n1313), .B(n1431), .ZN(n939) );
  XNOR2_X1 U1597 ( .A(n1538), .B(n1340), .ZN(n1036) );
  XNOR2_X1 U1598 ( .A(n1311), .B(n1402), .ZN(n908) );
  XNOR2_X1 U1599 ( .A(n1534), .B(n1352), .ZN(n956) );
  XNOR2_X1 U1600 ( .A(n1531), .B(n1430), .ZN(n938) );
  XNOR2_X1 U1601 ( .A(n1312), .B(n1524), .ZN(n1044) );
  XNOR2_X1 U1602 ( .A(n1256), .B(n1402), .ZN(n919) );
  XNOR2_X1 U1603 ( .A(n1533), .B(n1431), .ZN(n936) );
  XNOR2_X1 U1604 ( .A(n1342), .B(n1340), .ZN(n1040) );
  XNOR2_X1 U1605 ( .A(n1312), .B(n1402), .ZN(n918) );
  XNOR2_X1 U1606 ( .A(n1535), .B(n1328), .ZN(n955) );
  XNOR2_X1 U1607 ( .A(n1530), .B(n1352), .ZN(n960) );
  XNOR2_X1 U1608 ( .A(n1536), .B(n1352), .ZN(n954) );
  XNOR2_X1 U1609 ( .A(n1534), .B(n1430), .ZN(n935) );
  XNOR2_X1 U1610 ( .A(n1540), .B(n1328), .ZN(n949) );
  XNOR2_X1 U1611 ( .A(n1538), .B(n1402), .ZN(n910) );
  XNOR2_X1 U1612 ( .A(n1537), .B(n1340), .ZN(n1037) );
  XNOR2_X1 U1613 ( .A(n1256), .B(n1340), .ZN(n1045) );
  XNOR2_X1 U1614 ( .A(n1306), .B(n1430), .ZN(n930) );
  XNOR2_X1 U1615 ( .A(n1529), .B(n1328), .ZN(n961) );
  XNOR2_X1 U1616 ( .A(n1544), .B(n1524), .ZN(n1029) );
  XNOR2_X1 U1617 ( .A(n1310), .B(n1431), .ZN(n929) );
  XNOR2_X1 U1618 ( .A(n1330), .B(n1352), .ZN(n948) );
  XNOR2_X1 U1619 ( .A(n1537), .B(n1402), .ZN(n911) );
  XNOR2_X1 U1620 ( .A(n1533), .B(n1402), .ZN(n915) );
  XNOR2_X1 U1621 ( .A(n1537), .B(n1352), .ZN(n953) );
  XNOR2_X1 U1622 ( .A(n1535), .B(n1431), .ZN(n934) );
  XNOR2_X1 U1623 ( .A(n1545), .B(n1524), .ZN(n1028) );
  XNOR2_X1 U1624 ( .A(n1311), .B(n1328), .ZN(n950) );
  XNOR2_X1 U1625 ( .A(n1542), .B(n1328), .ZN(n947) );
  XNOR2_X1 U1626 ( .A(n1538), .B(n1431), .ZN(n931) );
  XNOR2_X1 U1627 ( .A(n1306), .B(n1401), .ZN(n909) );
  XNOR2_X1 U1628 ( .A(n1341), .B(n1401), .ZN(n914) );
  XNOR2_X1 U1629 ( .A(n1540), .B(n1430), .ZN(n928) );
  XNOR2_X1 U1630 ( .A(n1346), .B(n1401), .ZN(n912) );
  XNOR2_X1 U1631 ( .A(n1346), .B(n1430), .ZN(n933) );
  XNOR2_X1 U1632 ( .A(n1538), .B(n1352), .ZN(n952) );
  XNOR2_X1 U1633 ( .A(n1537), .B(n1430), .ZN(n932) );
  XNOR2_X1 U1634 ( .A(n1306), .B(n1328), .ZN(n951) );
  XNOR2_X1 U1635 ( .A(n1535), .B(n1401), .ZN(n913) );
  XNOR2_X1 U1636 ( .A(n1360), .B(n1430), .ZN(n924) );
  XNOR2_X1 U1637 ( .A(n1545), .B(n1430), .ZN(n923) );
  XNOR2_X1 U1638 ( .A(n1327), .B(n1401), .ZN(n905) );
  XNOR2_X1 U1639 ( .A(n1300), .B(n1402), .ZN(n904) );
  XNOR2_X1 U1640 ( .A(n1360), .B(n1401), .ZN(n903) );
  XNOR2_X1 U1641 ( .A(n1545), .B(n1402), .ZN(n902) );
  XNOR2_X1 U1642 ( .A(n1256), .B(n1451), .ZN(n1003) );
  XNOR2_X1 U1643 ( .A(n1536), .B(n1450), .ZN(n996) );
  XNOR2_X1 U1644 ( .A(n1535), .B(n1451), .ZN(n997) );
  XNOR2_X1 U1645 ( .A(n1313), .B(n1451), .ZN(n1002) );
  XNOR2_X1 U1646 ( .A(n1539), .B(n1451), .ZN(n993) );
  XNOR2_X1 U1647 ( .A(n1311), .B(n1450), .ZN(n992) );
  XNOR2_X1 U1648 ( .A(n1538), .B(n1450), .ZN(n994) );
  XNOR2_X1 U1649 ( .A(n1537), .B(n1451), .ZN(n995) );
  XNOR2_X1 U1650 ( .A(n1341), .B(n1451), .ZN(n998) );
  XNOR2_X1 U1651 ( .A(n1531), .B(n1450), .ZN(n1001) );
  XNOR2_X1 U1652 ( .A(n1544), .B(n1450), .ZN(n987) );
  XNOR2_X1 U1653 ( .A(n1540), .B(n1451), .ZN(n991) );
  XNOR2_X1 U1654 ( .A(n1532), .B(n1451), .ZN(n1000) );
  XNOR2_X1 U1655 ( .A(n1533), .B(n1451), .ZN(n999) );
  XNOR2_X1 U1656 ( .A(n1545), .B(n1451), .ZN(n986) );
  XNOR2_X1 U1657 ( .A(n1543), .B(n1450), .ZN(n988) );
  XNOR2_X1 U1658 ( .A(n1541), .B(n1450), .ZN(n990) );
  XNOR2_X1 U1659 ( .A(n1542), .B(n1450), .ZN(n989) );
  XNOR2_X1 U1660 ( .A(n1306), .B(n1367), .ZN(n888) );
  XNOR2_X1 U1661 ( .A(n1538), .B(n1368), .ZN(n889) );
  XNOR2_X1 U1662 ( .A(n1529), .B(n1367), .ZN(n898) );
  XNOR2_X1 U1663 ( .A(n1313), .B(n1368), .ZN(n897) );
  XNOR2_X1 U1664 ( .A(n1535), .B(n1368), .ZN(n892) );
  XNOR2_X1 U1665 ( .A(n1536), .B(n1368), .ZN(n891) );
  XNOR2_X1 U1666 ( .A(n1531), .B(n1368), .ZN(n896) );
  XNOR2_X1 U1667 ( .A(n1532), .B(n1367), .ZN(n895) );
  XNOR2_X1 U1668 ( .A(n1342), .B(n1368), .ZN(n893) );
  XNOR2_X1 U1669 ( .A(n1537), .B(n1367), .ZN(n890) );
  XNOR2_X1 U1670 ( .A(n1533), .B(n1367), .ZN(n894) );
  XNOR2_X1 U1671 ( .A(n1310), .B(n1368), .ZN(n887) );
  XNOR2_X1 U1672 ( .A(n1540), .B(n1367), .ZN(n886) );
  XNOR2_X1 U1673 ( .A(n1330), .B(n1368), .ZN(n885) );
  XNOR2_X1 U1674 ( .A(n1327), .B(n1367), .ZN(n884) );
  XNOR2_X1 U1675 ( .A(n1360), .B(n1367), .ZN(n882) );
  XNOR2_X1 U1676 ( .A(n1545), .B(n1368), .ZN(n881) );
  XNOR2_X1 U1677 ( .A(n1300), .B(n1368), .ZN(n883) );
  AND2_X1 U1678 ( .A1(n1298), .A2(n665), .ZN(n859) );
  INV_X1 U1679 ( .A(n314), .ZN(n315) );
  INV_X1 U1680 ( .A(n304), .ZN(n305) );
  OAI22_X1 U1681 ( .A1(n1355), .A2(n1071), .B1(n1299), .B2(n1331), .ZN(n862)
         );
  AND2_X1 U1682 ( .A1(n1528), .A2(n641), .ZN(n699) );
  INV_X1 U1683 ( .A(n649), .ZN(n740) );
  INV_X1 U1684 ( .A(n643), .ZN(n700) );
  INV_X1 U1685 ( .A(n346), .ZN(n347) );
  OAI22_X1 U1686 ( .A1(n1355), .A2(n1073), .B1(n1072), .B2(n1331), .ZN(n864)
         );
  AND2_X1 U1687 ( .A1(n1298), .A2(n644), .ZN(n719) );
  AND2_X1 U1688 ( .A1(n1528), .A2(n650), .ZN(n759) );
  OAI22_X1 U1689 ( .A1(n1355), .A2(n1077), .B1(n1076), .B2(n1332), .ZN(n868)
         );
  INV_X1 U1690 ( .A(n667), .ZN(n860) );
  INV_X1 U1691 ( .A(n652), .ZN(n760) );
  INV_X1 U1692 ( .A(n646), .ZN(n720) );
  OAI22_X1 U1693 ( .A1(n1362), .A2(n1080), .B1(n1079), .B2(n1331), .ZN(n871)
         );
  INV_X1 U1694 ( .A(n424), .ZN(n425) );
  AND2_X1 U1695 ( .A1(n1528), .A2(n653), .ZN(n779) );
  OAI22_X1 U1696 ( .A1(n1361), .A2(n1079), .B1(n1078), .B2(n1331), .ZN(n870)
         );
  AND2_X1 U1697 ( .A1(n1528), .A2(n647), .ZN(n739) );
  OAI22_X1 U1698 ( .A1(n1362), .A2(n1075), .B1(n1074), .B2(n1331), .ZN(n866)
         );
  AND2_X1 U1699 ( .A1(n1528), .A2(n659), .ZN(n819) );
  OAI22_X1 U1700 ( .A1(n1454), .A2(n1083), .B1(n1082), .B2(n1331), .ZN(n874)
         );
  OAI22_X1 U1701 ( .A1(n1454), .A2(n1247), .B1(n1077), .B2(n1332), .ZN(n869)
         );
  OAI22_X1 U1702 ( .A1(n1362), .A2(n1076), .B1(n1075), .B2(n1331), .ZN(n867)
         );
  INV_X1 U1703 ( .A(n458), .ZN(n459) );
  INV_X1 U1704 ( .A(n1430), .ZN(n1142) );
  INV_X1 U1705 ( .A(n1402), .ZN(n1141) );
  INV_X1 U1706 ( .A(n1328), .ZN(n1143) );
  INV_X1 U1707 ( .A(n1524), .ZN(n1147) );
  OAI22_X1 U1708 ( .A1(n1454), .A2(n1070), .B1(n1320), .B2(n1331), .ZN(n861)
         );
  INV_X1 U1709 ( .A(n368), .ZN(n369) );
  INV_X1 U1710 ( .A(n640), .ZN(n680) );
  XNOR2_X1 U1711 ( .A(n1527), .B(n1328), .ZN(n962) );
  XNOR2_X1 U1712 ( .A(n1527), .B(n1367), .ZN(n899) );
  INV_X1 U1713 ( .A(n658), .ZN(n800) );
  INV_X1 U1714 ( .A(n655), .ZN(n780) );
  INV_X1 U1715 ( .A(n1451), .ZN(n1145) );
  INV_X1 U1716 ( .A(n1367), .ZN(n1140) );
  OR2_X1 U1717 ( .A1(n1527), .A2(n1145), .ZN(n1005) );
  OR2_X1 U1718 ( .A1(n1527), .A2(n1142), .ZN(n942) );
  OR2_X1 U1719 ( .A1(n1527), .A2(n1141), .ZN(n921) );
  OR2_X1 U1720 ( .A1(n1528), .A2(n1146), .ZN(n1026) );
  OR2_X1 U1721 ( .A1(n1528), .A2(n1140), .ZN(n900) );
  OR2_X1 U1722 ( .A1(n1528), .A2(n1143), .ZN(n963) );
  OR2_X1 U1723 ( .A1(n1528), .A2(n1144), .ZN(n984) );
  XNOR2_X1 U1724 ( .A(n1365), .B(n1367), .ZN(n880) );
  AND2_X1 U1725 ( .A1(n1298), .A2(n1248), .ZN(product[0]) );
  XNOR2_X1 U1726 ( .A(n49), .B(a[18]), .ZN(n58) );
  XNOR2_X1 U1727 ( .A(n7), .B(a[4]), .ZN(n16) );
  XNOR2_X1 U1728 ( .A(n19), .B(a[8]), .ZN(n28) );
  XNOR2_X1 U1729 ( .A(n1526), .B(a[16]), .ZN(n52) );
  XNOR2_X1 U1730 ( .A(n31), .B(a[12]), .ZN(n40) );
  XNOR2_X1 U1731 ( .A(n25), .B(a[10]), .ZN(n34) );
  XNOR2_X1 U1732 ( .A(n13), .B(a[6]), .ZN(n22) );
  XNOR2_X1 U1733 ( .A(n1), .B(a[2]), .ZN(n9) );
  NOR2_X1 U1734 ( .A1(n1399), .A2(n209), .ZN(n202) );
  OAI21_X1 U1735 ( .B1(n204), .B2(n210), .A(n205), .ZN(n203) );
  NAND2_X1 U1736 ( .A1(n557), .A2(n568), .ZN(n205) );
  XNOR2_X1 U1737 ( .A(n1533), .B(n1319), .ZN(n1062) );
  XNOR2_X1 U1738 ( .A(n1347), .B(n1319), .ZN(n1059) );
  INV_X1 U1739 ( .A(n1319), .ZN(n1148) );
  XNOR2_X1 U1740 ( .A(n1542), .B(n1523), .ZN(n1052) );
  XNOR2_X1 U1741 ( .A(n1543), .B(n1523), .ZN(n1051) );
  XNOR2_X1 U1742 ( .A(n1544), .B(n1523), .ZN(n1050) );
  XNOR2_X1 U1743 ( .A(n1545), .B(n1523), .ZN(n1049) );
  XNOR2_X1 U1744 ( .A(n1341), .B(n1523), .ZN(n1061) );
  XNOR2_X1 U1745 ( .A(n1535), .B(n1523), .ZN(n1060) );
  XNOR2_X1 U1746 ( .A(n1310), .B(n1319), .ZN(n1055) );
  XNOR2_X1 U1747 ( .A(n1539), .B(n1319), .ZN(n1056) );
  XNOR2_X1 U1748 ( .A(n1359), .B(n1319), .ZN(n1064) );
  XNOR2_X1 U1749 ( .A(n1324), .B(n1523), .ZN(n1063) );
  XNOR2_X1 U1750 ( .A(n1527), .B(n1319), .ZN(n1067) );
  XNOR2_X1 U1751 ( .A(n1540), .B(n1319), .ZN(n1054) );
  XNOR2_X1 U1752 ( .A(n1537), .B(n1319), .ZN(n1058) );
  XNOR2_X1 U1753 ( .A(n1538), .B(n1319), .ZN(n1057) );
  XNOR2_X1 U1754 ( .A(n1541), .B(n1319), .ZN(n1053) );
  XNOR2_X1 U1755 ( .A(n1546), .B(n1523), .ZN(n1048) );
  XNOR2_X1 U1756 ( .A(n1256), .B(n1319), .ZN(n1066) );
  XNOR2_X1 U1757 ( .A(n1312), .B(n1319), .ZN(n1065) );
  XNOR2_X1 U1758 ( .A(n1546), .B(n1336), .ZN(n1006) );
  INV_X1 U1759 ( .A(n1337), .ZN(n1146) );
  XNOR2_X1 U1760 ( .A(n1545), .B(n1336), .ZN(n1007) );
  XNOR2_X1 U1761 ( .A(n1527), .B(n1336), .ZN(n1025) );
  XNOR2_X1 U1762 ( .A(n1543), .B(n1337), .ZN(n1009) );
  XNOR2_X1 U1763 ( .A(n1544), .B(n1337), .ZN(n1008) );
  XNOR2_X1 U1764 ( .A(n1256), .B(n1336), .ZN(n1024) );
  XNOR2_X1 U1765 ( .A(n1097), .B(n1525), .ZN(n1013) );
  XNOR2_X1 U1766 ( .A(n1306), .B(n1337), .ZN(n1014) );
  XNOR2_X1 U1767 ( .A(n1540), .B(n1525), .ZN(n1012) );
  XNOR2_X1 U1768 ( .A(n1313), .B(n1337), .ZN(n1023) );
  XNOR2_X1 U1769 ( .A(n1535), .B(n1336), .ZN(n1018) );
  XNOR2_X1 U1770 ( .A(n1542), .B(n1336), .ZN(n1010) );
  XNOR2_X1 U1771 ( .A(n1541), .B(n1337), .ZN(n1011) );
  XNOR2_X1 U1772 ( .A(n1533), .B(n1336), .ZN(n1020) );
  XNOR2_X1 U1773 ( .A(n1341), .B(n1337), .ZN(n1019) );
  XNOR2_X1 U1774 ( .A(n1532), .B(n1525), .ZN(n1021) );
  XNOR2_X1 U1775 ( .A(n1537), .B(n1336), .ZN(n1016) );
  XNOR2_X1 U1776 ( .A(n1347), .B(n1337), .ZN(n1017) );
  XNOR2_X1 U1777 ( .A(n1538), .B(n1337), .ZN(n1015) );
  XOR2_X1 U1778 ( .A(n19), .B(a[6]), .Z(n1116) );
  XNOR2_X1 U1779 ( .A(n1365), .B(n1322), .ZN(n964) );
  XNOR2_X1 U1780 ( .A(n1545), .B(n1323), .ZN(n965) );
  XNOR2_X1 U1781 ( .A(n1360), .B(n1322), .ZN(n966) );
  XNOR2_X1 U1782 ( .A(n1543), .B(n1323), .ZN(n967) );
  XNOR2_X1 U1783 ( .A(n1306), .B(n1322), .ZN(n972) );
  XNOR2_X1 U1784 ( .A(n1542), .B(n1322), .ZN(n968) );
  XNOR2_X1 U1785 ( .A(n1311), .B(n1323), .ZN(n971) );
  XNOR2_X1 U1786 ( .A(n1541), .B(n1322), .ZN(n969) );
  XNOR2_X1 U1787 ( .A(n1540), .B(n1323), .ZN(n970) );
  XNOR2_X1 U1788 ( .A(n1346), .B(n1322), .ZN(n975) );
  XNOR2_X1 U1789 ( .A(n1535), .B(n1322), .ZN(n976) );
  XNOR2_X1 U1790 ( .A(n1538), .B(n1323), .ZN(n973) );
  XNOR2_X1 U1791 ( .A(n1537), .B(n1323), .ZN(n974) );
  INV_X1 U1792 ( .A(n1323), .ZN(n1144) );
  XNOR2_X1 U1793 ( .A(n1527), .B(n1323), .ZN(n983) );
  XNOR2_X1 U1794 ( .A(n1342), .B(n1322), .ZN(n977) );
  XNOR2_X1 U1795 ( .A(n1256), .B(n1322), .ZN(n982) );
  XNOR2_X1 U1796 ( .A(n1533), .B(n1322), .ZN(n978) );
  XNOR2_X1 U1797 ( .A(n1324), .B(n1323), .ZN(n979) );
  XNOR2_X1 U1798 ( .A(n1530), .B(n1323), .ZN(n981) );
  XNOR2_X1 U1799 ( .A(n1358), .B(n1322), .ZN(n980) );
  OAI21_X1 U1800 ( .B1(n141), .B2(n135), .A(n136), .ZN(n134) );
  INV_X1 U1801 ( .A(n661), .ZN(n820) );
  INV_X1 U1802 ( .A(n187), .ZN(n282) );
  OAI21_X1 U1803 ( .B1(n193), .B2(n187), .A(n188), .ZN(n186) );
  NOR2_X1 U1804 ( .A1(n529), .A2(n542), .ZN(n187) );
  AOI21_X1 U1805 ( .B1(n1495), .B2(n230), .A(n1271), .ZN(n223) );
  INV_X1 U1806 ( .A(n664), .ZN(n840) );
  NAND2_X1 U1807 ( .A1(n145), .A2(n133), .ZN(n131) );
  INV_X1 U1808 ( .A(n140), .ZN(n273) );
  NOR2_X1 U1809 ( .A1(n140), .A2(n1318), .ZN(n133) );
  NOR2_X1 U1810 ( .A1(n383), .A2(n396), .ZN(n140) );
  OAI21_X1 U1811 ( .B1(n147), .B2(n151), .A(n148), .ZN(n146) );
  AOI21_X1 U1812 ( .B1(n146), .B2(n133), .A(n134), .ZN(n132) );
  INV_X1 U1813 ( .A(n234), .ZN(n233) );
  OAI21_X1 U1814 ( .B1(n222), .B2(n234), .A(n223), .ZN(n221) );
  AOI21_X1 U1815 ( .B1(n239), .B2(n1484), .A(n236), .ZN(n234) );
  OAI21_X1 U1816 ( .B1(n242), .B2(n240), .A(n241), .ZN(n239) );
  XOR2_X1 U1817 ( .A(n1235), .B(n89), .Z(product[7]) );
  XNOR2_X1 U1818 ( .A(n1544), .B(n1305), .ZN(n1071) );
  XNOR2_X1 U1819 ( .A(n1545), .B(n1383), .ZN(n1070) );
  XNOR2_X1 U1820 ( .A(n1540), .B(n1305), .ZN(n1075) );
  XNOR2_X1 U1821 ( .A(n1311), .B(n1305), .ZN(n1076) );
  XNOR2_X1 U1822 ( .A(n1539), .B(n1383), .ZN(n1077) );
  XNOR2_X1 U1823 ( .A(n1347), .B(n1383), .ZN(n1080) );
  XNOR2_X1 U1824 ( .A(n1535), .B(n1305), .ZN(n1081) );
  XNOR2_X1 U1825 ( .A(n1543), .B(n1383), .ZN(n1072) );
  XNOR2_X1 U1826 ( .A(n1541), .B(n1383), .ZN(n1074) );
  XNOR2_X1 U1827 ( .A(n1542), .B(n1383), .ZN(n1073) );
  XNOR2_X1 U1828 ( .A(n1537), .B(n1383), .ZN(n1079) );
  XNOR2_X1 U1829 ( .A(n1538), .B(n1305), .ZN(n1078) );
  XNOR2_X1 U1830 ( .A(n1534), .B(n1383), .ZN(n1082) );
  XNOR2_X1 U1831 ( .A(n1533), .B(n1305), .ZN(n1083) );
  XNOR2_X1 U1832 ( .A(n1305), .B(n1546), .ZN(n1069) );
  XNOR2_X1 U1833 ( .A(n1312), .B(n1307), .ZN(n1086) );
  XNOR2_X1 U1834 ( .A(n1358), .B(n1383), .ZN(n1085) );
  XNOR2_X1 U1835 ( .A(n1527), .B(n1307), .ZN(n1088) );
  XNOR2_X1 U1836 ( .A(n1532), .B(n1305), .ZN(n1084) );
  XNOR2_X1 U1837 ( .A(n1256), .B(n1305), .ZN(n1087) );
  INV_X1 U1838 ( .A(n1383), .ZN(n1149) );
  NAND2_X1 U1839 ( .A1(n156), .A2(n164), .ZN(n154) );
  NAND2_X1 U1840 ( .A1(n461), .A2(n478), .ZN(n167) );
  OAI21_X1 U1841 ( .B1(n158), .B2(n162), .A(n159), .ZN(n157) );
  NAND2_X1 U1842 ( .A1(n427), .A2(n442), .ZN(n159) );
  OAI21_X1 U1843 ( .B1(n193), .B2(n180), .A(n1366), .ZN(n179) );
  NAND2_X1 U1844 ( .A1(n513), .A2(n528), .ZN(n185) );
  OAI21_X1 U1845 ( .B1(n152), .B2(n150), .A(n1435), .ZN(n149) );
  INV_X1 U1846 ( .A(n150), .ZN(n275) );
  NOR2_X1 U1847 ( .A1(n150), .A2(n1481), .ZN(n145) );
  NOR2_X1 U1848 ( .A1(n411), .A2(n426), .ZN(n150) );
  OAI21_X1 U1849 ( .B1(n163), .B2(n1295), .A(n1333), .ZN(n160) );
  INV_X1 U1850 ( .A(n1295), .ZN(n277) );
  NOR2_X1 U1851 ( .A1(n161), .A2(n1473), .ZN(n156) );
  XNOR2_X1 U1852 ( .A(n715), .B(n1242), .ZN(n477) );
  OR2_X1 U1853 ( .A1(n787), .A2(n715), .ZN(n476) );
  NAND2_X1 U1854 ( .A1(n1493), .A2(n185), .ZN(n79) );
  OAI22_X1 U1855 ( .A1(n1394), .A2(n965), .B1(n964), .B2(n1351), .ZN(n346) );
  OAI22_X1 U1856 ( .A1(n964), .A2(n1393), .B1(n964), .B2(n1350), .ZN(n652) );
  OAI22_X1 U1857 ( .A1(n1393), .A2(n966), .B1(n965), .B2(n1350), .ZN(n761) );
  OAI22_X1 U1858 ( .A1(n1394), .A2(n967), .B1(n966), .B2(n1351), .ZN(n762) );
  OAI22_X1 U1859 ( .A1(n1393), .A2(n968), .B1(n967), .B2(n1350), .ZN(n763) );
  OAI22_X1 U1860 ( .A1(n1393), .A2(n975), .B1(n974), .B2(n1351), .ZN(n770) );
  OAI22_X1 U1861 ( .A1(n1393), .A2(n973), .B1(n972), .B2(n1350), .ZN(n768) );
  OAI22_X1 U1862 ( .A1(n1394), .A2(n972), .B1(n971), .B2(n1351), .ZN(n767) );
  OAI22_X1 U1863 ( .A1(n1394), .A2(n1144), .B1(n984), .B2(n1350), .ZN(n674) );
  OAI22_X1 U1864 ( .A1(n1393), .A2(n977), .B1(n976), .B2(n1351), .ZN(n772) );
  OAI22_X1 U1865 ( .A1(n1394), .A2(n969), .B1(n968), .B2(n1351), .ZN(n764) );
  OAI22_X1 U1866 ( .A1(n1393), .A2(n982), .B1(n981), .B2(n1351), .ZN(n777) );
  OAI22_X1 U1867 ( .A1(n1393), .A2(n976), .B1(n975), .B2(n1351), .ZN(n771) );
  OAI22_X1 U1868 ( .A1(n1393), .A2(n983), .B1(n982), .B2(n1350), .ZN(n778) );
  OAI22_X1 U1869 ( .A1(n1394), .A2(n971), .B1(n970), .B2(n1351), .ZN(n766) );
  OAI22_X1 U1870 ( .A1(n1393), .A2(n970), .B1(n969), .B2(n1351), .ZN(n765) );
  OAI22_X1 U1871 ( .A1(n1393), .A2(n980), .B1(n979), .B2(n1351), .ZN(n775) );
  OAI22_X1 U1872 ( .A1(n1394), .A2(n978), .B1(n977), .B2(n1350), .ZN(n773) );
  OAI22_X1 U1873 ( .A1(n1394), .A2(n979), .B1(n978), .B2(n1350), .ZN(n774) );
  OAI22_X1 U1874 ( .A1(n1394), .A2(n974), .B1(n973), .B2(n1350), .ZN(n769) );
  INV_X1 U1875 ( .A(n1354), .ZN(n653) );
  OAI22_X1 U1876 ( .A1(n1394), .A2(n981), .B1(n980), .B2(n1350), .ZN(n776) );
  OAI22_X1 U1877 ( .A1(n943), .A2(n1374), .B1(n943), .B2(n1507), .ZN(n649) );
  OAI22_X1 U1878 ( .A1(n1370), .A2(n944), .B1(n943), .B2(n1507), .ZN(n328) );
  OAI22_X1 U1879 ( .A1(n1375), .A2(n945), .B1(n944), .B2(n1507), .ZN(n741) );
  OAI22_X1 U1880 ( .A1(n1370), .A2(n947), .B1(n946), .B2(n1507), .ZN(n743) );
  OAI22_X1 U1881 ( .A1(n1374), .A2(n946), .B1(n945), .B2(n1507), .ZN(n742) );
  OAI22_X1 U1882 ( .A1(n1370), .A2(n948), .B1(n947), .B2(n1507), .ZN(n744) );
  OAI22_X1 U1883 ( .A1(n1375), .A2(n949), .B1(n948), .B2(n1507), .ZN(n745) );
  OAI22_X1 U1884 ( .A1(n1472), .A2(n952), .B1(n951), .B2(n1507), .ZN(n748) );
  OAI22_X1 U1885 ( .A1(n1472), .A2(n958), .B1(n957), .B2(n1507), .ZN(n754) );
  OAI22_X1 U1886 ( .A1(n1374), .A2(n1143), .B1(n963), .B2(n1507), .ZN(n673) );
  OAI22_X1 U1887 ( .A1(n1472), .A2(n957), .B1(n956), .B2(n1507), .ZN(n753) );
  OAI22_X1 U1888 ( .A1(n1374), .A2(n950), .B1(n949), .B2(n1507), .ZN(n746) );
  OAI22_X1 U1889 ( .A1(n1277), .A2(n1287), .B1(n952), .B2(n1507), .ZN(n749) );
  OAI22_X1 U1890 ( .A1(n1375), .A2(n951), .B1(n950), .B2(n1507), .ZN(n747) );
  OAI22_X1 U1891 ( .A1(n1472), .A2(n956), .B1(n955), .B2(n1506), .ZN(n752) );
  OAI22_X1 U1892 ( .A1(n1472), .A2(n960), .B1(n959), .B2(n1506), .ZN(n756) );
  INV_X1 U1893 ( .A(n1506), .ZN(n650) );
  OAI22_X1 U1894 ( .A1(n1277), .A2(n961), .B1(n960), .B2(n1507), .ZN(n757) );
  OAI22_X1 U1895 ( .A1(n1375), .A2(n955), .B1(n954), .B2(n1506), .ZN(n751) );
  OAI22_X1 U1896 ( .A1(n1374), .A2(n959), .B1(n958), .B2(n1507), .ZN(n755) );
  OAI22_X1 U1897 ( .A1(n1375), .A2(n962), .B1(n961), .B2(n1506), .ZN(n758) );
  OAI22_X1 U1898 ( .A1(n954), .A2(n42), .B1(n953), .B2(n1506), .ZN(n750) );
  INV_X1 U1899 ( .A(n166), .ZN(n278) );
  AOI21_X1 U1900 ( .B1(n173), .B2(n164), .A(n165), .ZN(n163) );
  AOI21_X1 U1901 ( .B1(n156), .B2(n165), .A(n157), .ZN(n155) );
  NOR2_X1 U1902 ( .A1(n166), .A2(n171), .ZN(n164) );
  OAI21_X1 U1903 ( .B1(n166), .B2(n172), .A(n167), .ZN(n165) );
  INV_X1 U1904 ( .A(n1508), .ZN(n647) );
  INV_X1 U1905 ( .A(n194), .ZN(n193) );
  INV_X1 U1906 ( .A(n1316), .ZN(n173) );
  OAI21_X1 U1907 ( .B1(n152), .B2(n131), .A(n1348), .ZN(n130) );
  OAI22_X1 U1908 ( .A1(n901), .A2(n1325), .B1(n901), .B2(n1505), .ZN(n643) );
  OAI22_X1 U1909 ( .A1(n1234), .A2(n902), .B1(n901), .B2(n1505), .ZN(n304) );
  OAI22_X1 U1910 ( .A1(n1325), .A2(n903), .B1(n902), .B2(n1505), .ZN(n701) );
  OAI21_X1 U1911 ( .B1(n132), .B2(n128), .A(n129), .ZN(n127) );
  OAI22_X1 U1912 ( .A1(n1325), .A2(n905), .B1(n904), .B2(n1505), .ZN(n703) );
  OAI22_X1 U1913 ( .A1(n1325), .A2(n904), .B1(n903), .B2(n1505), .ZN(n702) );
  OAI22_X1 U1914 ( .A1(n1325), .A2(n906), .B1(n905), .B2(n1505), .ZN(n704) );
  OAI22_X1 U1915 ( .A1(n1325), .A2(n907), .B1(n906), .B2(n1505), .ZN(n705) );
  OAI22_X1 U1916 ( .A1(n1325), .A2(n909), .B1(n908), .B2(n1505), .ZN(n707) );
  OAI22_X1 U1917 ( .A1(n1234), .A2(n908), .B1(n907), .B2(n1505), .ZN(n706) );
  OAI22_X1 U1918 ( .A1(n1325), .A2(n910), .B1(n909), .B2(n1505), .ZN(n708) );
  OAI22_X1 U1919 ( .A1(n1325), .A2(n911), .B1(n910), .B2(n1505), .ZN(n709) );
  OAI22_X1 U1920 ( .A1(n1234), .A2(n915), .B1(n914), .B2(n1505), .ZN(n713) );
  OAI22_X1 U1921 ( .A1(n1233), .A2(n912), .B1(n911), .B2(n1315), .ZN(n710) );
  OAI22_X1 U1922 ( .A1(n1234), .A2(n913), .B1(n912), .B2(n1315), .ZN(n711) );
  OAI22_X1 U1923 ( .A1(n1234), .A2(n914), .B1(n913), .B2(n1315), .ZN(n712) );
  OAI22_X1 U1924 ( .A1(n1233), .A2(n1141), .B1(n921), .B2(n1315), .ZN(n671) );
  OAI22_X1 U1925 ( .A1(n1234), .A2(n918), .B1(n917), .B2(n1315), .ZN(n716) );
  OAI22_X1 U1926 ( .A1(n1233), .A2(n919), .B1(n918), .B2(n1315), .ZN(n717) );
  OAI22_X1 U1927 ( .A1(n1234), .A2(n920), .B1(n919), .B2(n1315), .ZN(n718) );
  OAI22_X1 U1928 ( .A1(n1234), .A2(n917), .B1(n916), .B2(n1315), .ZN(n715) );
  OAI22_X1 U1929 ( .A1(n1233), .A2(n916), .B1(n915), .B2(n1315), .ZN(n714) );
  INV_X1 U1930 ( .A(n1315), .ZN(n644) );
  NAND2_X1 U1931 ( .A1(n202), .A2(n1492), .ZN(n195) );
  AOI21_X1 U1932 ( .B1(n203), .B2(n1492), .A(n198), .ZN(n196) );
  AOI21_X1 U1933 ( .B1(n194), .B2(n175), .A(n176), .ZN(n174) );
  OAI21_X1 U1934 ( .B1(n181), .B2(n177), .A(n178), .ZN(n176) );
  OAI22_X1 U1935 ( .A1(n922), .A2(n1353), .B1(n922), .B2(n1326), .ZN(n646) );
  OAI22_X1 U1936 ( .A1(n1353), .A2(n924), .B1(n923), .B2(n1326), .ZN(n721) );
  OAI22_X1 U1937 ( .A1(n1353), .A2(n923), .B1(n922), .B2(n1326), .ZN(n314) );
  OAI22_X1 U1938 ( .A1(n1353), .A2(n925), .B1(n924), .B2(n1326), .ZN(n722) );
  OAI22_X1 U1939 ( .A1(n1339), .A2(n927), .B1(n926), .B2(n1326), .ZN(n724) );
  OAI22_X1 U1940 ( .A1(n1339), .A2(n926), .B1(n925), .B2(n1326), .ZN(n723) );
  OAI22_X1 U1941 ( .A1(n1339), .A2(n928), .B1(n927), .B2(n1326), .ZN(n725) );
  OAI22_X1 U1942 ( .A1(n1339), .A2(n929), .B1(n928), .B2(n1326), .ZN(n726) );
  OAI22_X1 U1943 ( .A1(n1339), .A2(n930), .B1(n929), .B2(n1326), .ZN(n727) );
  OAI22_X1 U1944 ( .A1(n1272), .A2(n931), .B1(n930), .B2(n1309), .ZN(n728) );
  OAI22_X1 U1945 ( .A1(n1314), .A2(n933), .B1(n932), .B2(n1309), .ZN(n730) );
  OAI22_X1 U1946 ( .A1(n1272), .A2(n934), .B1(n933), .B2(n1309), .ZN(n731) );
  OAI22_X1 U1947 ( .A1(n48), .A2(n941), .B1(n940), .B2(n1508), .ZN(n738) );
  OAI22_X1 U1948 ( .A1(n1272), .A2(n932), .B1(n931), .B2(n1309), .ZN(n729) );
  OAI22_X1 U1949 ( .A1(n1272), .A2(n1142), .B1(n942), .B2(n1309), .ZN(n672) );
  OAI22_X1 U1950 ( .A1(n1272), .A2(n936), .B1(n935), .B2(n1309), .ZN(n733) );
  OAI22_X1 U1951 ( .A1(n1272), .A2(n937), .B1(n936), .B2(n1508), .ZN(n734) );
  OAI22_X1 U1952 ( .A1(n1272), .A2(n939), .B1(n938), .B2(n1309), .ZN(n736) );
  OAI22_X1 U1953 ( .A1(n48), .A2(n935), .B1(n934), .B2(n1309), .ZN(n732) );
  OAI22_X1 U1954 ( .A1(n1314), .A2(n940), .B1(n939), .B2(n1309), .ZN(n737) );
  OAI22_X1 U1955 ( .A1(n48), .A2(n938), .B1(n937), .B2(n1309), .ZN(n735) );
  NAND3_X1 U1956 ( .A1(n1516), .A2(n1515), .A3(n1517), .ZN(n1512) );
  OAI21_X1 U1957 ( .B1(n1386), .B2(n123), .A(n124), .ZN(n1513) );
  OAI22_X1 U1958 ( .A1(n880), .A2(n1379), .B1(n880), .B2(n1251), .ZN(n640) );
  OAI22_X1 U1959 ( .A1(n1379), .A2(n881), .B1(n880), .B2(n1251), .ZN(n298) );
  OAI22_X1 U1960 ( .A1(n1379), .A2(n882), .B1(n881), .B2(n1251), .ZN(n681) );
  OAI22_X1 U1961 ( .A1(n1379), .A2(n883), .B1(n882), .B2(n1251), .ZN(n682) );
  OAI22_X1 U1962 ( .A1(n1379), .A2(n884), .B1(n883), .B2(n1251), .ZN(n683) );
  OAI22_X1 U1963 ( .A1(n1379), .A2(n886), .B1(n885), .B2(n1251), .ZN(n685) );
  OAI22_X1 U1964 ( .A1(n1379), .A2(n885), .B1(n884), .B2(n1251), .ZN(n684) );
  OAI22_X1 U1965 ( .A1(n1379), .A2(n887), .B1(n886), .B2(n1251), .ZN(n686) );
  OAI22_X1 U1966 ( .A1(n1379), .A2(n888), .B1(n887), .B2(n1251), .ZN(n687) );
  OAI22_X1 U1967 ( .A1(n1379), .A2(n889), .B1(n888), .B2(n1251), .ZN(n688) );
  OAI22_X1 U1968 ( .A1(n1379), .A2(n890), .B1(n889), .B2(n1251), .ZN(n689) );
  OAI22_X1 U1969 ( .A1(n1379), .A2(n891), .B1(n890), .B2(n1503), .ZN(n690) );
  OAI22_X1 U1970 ( .A1(n1379), .A2(n892), .B1(n891), .B2(n1503), .ZN(n691) );
  OAI22_X1 U1971 ( .A1(n1380), .A2(n894), .B1(n893), .B2(n1503), .ZN(n693) );
  OAI22_X1 U1972 ( .A1(n1380), .A2(n893), .B1(n892), .B2(n1503), .ZN(n692) );
  OAI22_X1 U1973 ( .A1(n1273), .A2(n899), .B1(n898), .B2(n1503), .ZN(n698) );
  OAI22_X1 U1974 ( .A1(n1380), .A2(n895), .B1(n894), .B2(n1503), .ZN(n694) );
  OAI22_X1 U1975 ( .A1(n1273), .A2(n1140), .B1(n900), .B2(n1503), .ZN(n670) );
  INV_X1 U1976 ( .A(n1503), .ZN(n641) );
  OAI22_X1 U1977 ( .A1(n1273), .A2(n898), .B1(n897), .B2(n1503), .ZN(n697) );
  OAI22_X1 U1978 ( .A1(n1380), .A2(n896), .B1(n895), .B2(n1503), .ZN(n695) );
  OAI22_X1 U1979 ( .A1(n1273), .A2(n897), .B1(n896), .B2(n1503), .ZN(n696) );
  OAI22_X1 U1980 ( .A1(n985), .A2(n1403), .B1(n985), .B2(n1414), .ZN(n655) );
  OAI22_X1 U1981 ( .A1(n1405), .A2(n986), .B1(n985), .B2(n1414), .ZN(n368) );
  OAI22_X1 U1982 ( .A1(n1405), .A2(n987), .B1(n986), .B2(n1414), .ZN(n781) );
  OAI22_X1 U1983 ( .A1(n1403), .A2(n1003), .B1(n1002), .B2(n1413), .ZN(n797)
         );
  OAI22_X1 U1984 ( .A1(n1403), .A2(n992), .B1(n991), .B2(n1414), .ZN(n786) );
  OAI22_X1 U1985 ( .A1(n1405), .A2(n989), .B1(n988), .B2(n1414), .ZN(n783) );
  OAI22_X1 U1986 ( .A1(n1405), .A2(n990), .B1(n989), .B2(n1414), .ZN(n784) );
  OAI22_X1 U1987 ( .A1(n1405), .A2(n999), .B1(n998), .B2(n1414), .ZN(n793) );
  OAI22_X1 U1988 ( .A1(n1405), .A2(n996), .B1(n995), .B2(n1414), .ZN(n790) );
  OAI22_X1 U1989 ( .A1(n1405), .A2(n991), .B1(n990), .B2(n1413), .ZN(n785) );
  OAI22_X1 U1990 ( .A1(n1405), .A2(n1000), .B1(n999), .B2(n1414), .ZN(n794) );
  OAI22_X1 U1991 ( .A1(n1403), .A2(n988), .B1(n987), .B2(n1414), .ZN(n782) );
  OAI22_X1 U1992 ( .A1(n1403), .A2(n1145), .B1(n1005), .B2(n1414), .ZN(n675)
         );
  OAI22_X1 U1993 ( .A1(n1404), .A2(n1002), .B1(n1001), .B2(n1414), .ZN(n796)
         );
  OAI22_X1 U1994 ( .A1(n1404), .A2(n993), .B1(n992), .B2(n1413), .ZN(n787) );
  OAI22_X1 U1995 ( .A1(n1405), .A2(n1004), .B1(n1003), .B2(n1414), .ZN(n798)
         );
  INV_X1 U1996 ( .A(n1413), .ZN(n656) );
  OAI22_X1 U1997 ( .A1(n1404), .A2(n994), .B1(n993), .B2(n1413), .ZN(n788) );
  OAI22_X1 U1998 ( .A1(n1405), .A2(n995), .B1(n994), .B2(n1414), .ZN(n789) );
  OAI22_X1 U1999 ( .A1(n1404), .A2(n1001), .B1(n1000), .B2(n1413), .ZN(n795)
         );
  OAI22_X1 U2000 ( .A1(n1404), .A2(n998), .B1(n997), .B2(n1414), .ZN(n792) );
  OAI22_X1 U2001 ( .A1(n1403), .A2(n997), .B1(n996), .B2(n1414), .ZN(n791) );
  XOR2_X1 U2002 ( .A(n300), .B(n299), .Z(n1514) );
  XOR2_X1 U2003 ( .A(n1334), .B(n1514), .Z(product[37]) );
  NAND2_X1 U2004 ( .A1(n300), .A2(n299), .ZN(n1515) );
  NAND2_X1 U2005 ( .A1(n1453), .A2(n300), .ZN(n1516) );
  NAND2_X1 U2006 ( .A1(n299), .A2(n98), .ZN(n1517) );
  NAND3_X1 U2007 ( .A1(n1516), .A2(n1515), .A3(n1517), .ZN(n97) );
  NAND2_X1 U2008 ( .A1(n680), .A2(n298), .ZN(n1518) );
  NAND2_X1 U2009 ( .A1(n1304), .A2(n680), .ZN(n1519) );
  NAND2_X1 U2010 ( .A1(n298), .A2(n97), .ZN(n1520) );
  AOI21_X1 U2011 ( .B1(n1513), .B2(n1496), .A(n119), .ZN(n1521) );
  CLKBUF_X1 U2012 ( .A(n153), .Z(n1522) );
  OAI21_X1 U2013 ( .B1(n125), .B2(n123), .A(n124), .ZN(n122) );
  INV_X1 U2014 ( .A(n1522), .ZN(n152) );
  OAI22_X1 U2015 ( .A1(n1406), .A2(n1014), .B1(n1013), .B2(n1509), .ZN(n807)
         );
  OAI22_X1 U2016 ( .A1(n1406), .A2(n1007), .B1(n1006), .B2(n1510), .ZN(n394)
         );
  OAI22_X1 U2017 ( .A1(n1006), .A2(n1406), .B1(n1006), .B2(n1509), .ZN(n658)
         );
  OAI22_X1 U2018 ( .A1(n1406), .A2(n1012), .B1(n1011), .B2(n1510), .ZN(n805)
         );
  OAI22_X1 U2019 ( .A1(n1406), .A2(n1021), .B1(n1020), .B2(n1510), .ZN(n814)
         );
  OAI22_X1 U2020 ( .A1(n1343), .A2(n1024), .B1(n1023), .B2(n1510), .ZN(n817)
         );
  OAI22_X1 U2021 ( .A1(n1343), .A2(n1010), .B1(n1009), .B2(n1509), .ZN(n803)
         );
  OAI22_X1 U2022 ( .A1(n1406), .A2(n1008), .B1(n1007), .B2(n1510), .ZN(n801)
         );
  OAI22_X1 U2023 ( .A1(n1406), .A2(n1009), .B1(n1008), .B2(n1509), .ZN(n802)
         );
  OAI22_X1 U2024 ( .A1(n1406), .A2(n1015), .B1(n1014), .B2(n1509), .ZN(n808)
         );
  OAI22_X1 U2025 ( .A1(n1406), .A2(n1146), .B1(n1026), .B2(n1509), .ZN(n676)
         );
  OAI22_X1 U2026 ( .A1(n1013), .A2(n1412), .B1(n1012), .B2(n1510), .ZN(n806)
         );
  OAI22_X1 U2027 ( .A1(n1343), .A2(n1025), .B1(n1024), .B2(n1509), .ZN(n818)
         );
  OAI22_X1 U2028 ( .A1(n1406), .A2(n1019), .B1(n1018), .B2(n1510), .ZN(n812)
         );
  OAI22_X1 U2029 ( .A1(n1406), .A2(n1020), .B1(n1019), .B2(n1510), .ZN(n813)
         );
  OAI22_X1 U2030 ( .A1(n1406), .A2(n1018), .B1(n1017), .B2(n1509), .ZN(n811)
         );
  OAI22_X1 U2031 ( .A1(n1412), .A2(n1011), .B1(n1010), .B2(n1509), .ZN(n804)
         );
  OAI22_X1 U2032 ( .A1(n1343), .A2(n1017), .B1(n1016), .B2(n1509), .ZN(n810)
         );
  OAI22_X1 U2033 ( .A1(n1343), .A2(n1023), .B1(n1321), .B2(n1510), .ZN(n816)
         );
  OAI22_X1 U2034 ( .A1(n1343), .A2(n1016), .B1(n1015), .B2(n1509), .ZN(n809)
         );
  OAI22_X1 U2035 ( .A1(n1412), .A2(n1321), .B1(n1021), .B2(n1510), .ZN(n815)
         );
  INV_X1 U2036 ( .A(n1510), .ZN(n659) );
  OAI21_X1 U2037 ( .B1(n174), .B2(n154), .A(n155), .ZN(n153) );
  INV_X1 U2038 ( .A(n101), .ZN(n264) );
  XNOR2_X1 U2039 ( .A(n1513), .B(n67), .ZN(product[29]) );
  XNOR2_X1 U2040 ( .A(n1392), .B(n65), .ZN(product[31]) );
  AOI21_X1 U2041 ( .B1(n1392), .B2(n1497), .A(n111), .ZN(n109) );
  AOI21_X1 U2042 ( .B1(n122), .B2(n1496), .A(n119), .ZN(n117) );
  OAI22_X1 U2043 ( .A1(n1274), .A2(n1039), .B1(n1038), .B2(n1409), .ZN(n831)
         );
  OAI22_X1 U2044 ( .A1(n1335), .A2(n1031), .B1(n1030), .B2(n1409), .ZN(n823)
         );
  OAI22_X1 U2045 ( .A1(n1335), .A2(n1032), .B1(n1031), .B2(n1415), .ZN(n824)
         );
  OAI22_X1 U2046 ( .A1(n1274), .A2(n1041), .B1(n1040), .B2(n1504), .ZN(n833)
         );
  OAI22_X1 U2047 ( .A1(n1274), .A2(n1034), .B1(n1033), .B2(n1504), .ZN(n826)
         );
  OAI22_X1 U2048 ( .A1(n1274), .A2(n1045), .B1(n1044), .B2(n1504), .ZN(n837)
         );
  OAI22_X1 U2049 ( .A1(n18), .A2(n1028), .B1(n1027), .B2(n1409), .ZN(n424) );
  OAI22_X1 U2050 ( .A1(n1027), .A2(n18), .B1(n1027), .B2(n1409), .ZN(n661) );
  OAI22_X1 U2051 ( .A1(n1335), .A2(n1038), .B1(n1037), .B2(n1504), .ZN(n830)
         );
  OAI22_X1 U2052 ( .A1(n1335), .A2(n1044), .B1(n1043), .B2(n1504), .ZN(n836)
         );
  OAI22_X1 U2053 ( .A1(n18), .A2(n1030), .B1(n1029), .B2(n1409), .ZN(n822) );
  OAI22_X1 U2054 ( .A1(n1335), .A2(n1029), .B1(n1028), .B2(n1415), .ZN(n821)
         );
  OAI22_X1 U2055 ( .A1(n18), .A2(n1033), .B1(n1032), .B2(n1415), .ZN(n825) );
  OAI22_X1 U2056 ( .A1(n1335), .A2(n1040), .B1(n1039), .B2(n1409), .ZN(n832)
         );
  OAI22_X1 U2057 ( .A1(n1335), .A2(n1037), .B1(n1036), .B2(n1504), .ZN(n829)
         );
  OAI22_X1 U2058 ( .A1(n1274), .A2(n1147), .B1(n1047), .B2(n1415), .ZN(n677)
         );
  OAI22_X1 U2059 ( .A1(n1335), .A2(n1036), .B1(n1035), .B2(n1415), .ZN(n828)
         );
  OAI22_X1 U2060 ( .A1(n1335), .A2(n1043), .B1(n1042), .B2(n1504), .ZN(n835)
         );
  OAI22_X1 U2061 ( .A1(n18), .A2(n1042), .B1(n1041), .B2(n1504), .ZN(n834) );
  OAI22_X1 U2062 ( .A1(n1335), .A2(n1035), .B1(n1034), .B2(n1504), .ZN(n827)
         );
  OAI22_X1 U2063 ( .A1(n18), .A2(n1046), .B1(n1045), .B2(n1415), .ZN(n838) );
  INV_X1 U2064 ( .A(n1504), .ZN(n662) );
  XNOR2_X1 U2065 ( .A(n1391), .B(n63), .ZN(product[33]) );
  XOR2_X1 U2066 ( .A(n109), .B(n64), .Z(product[32]) );
  XOR2_X1 U2067 ( .A(n1521), .B(n66), .Z(product[30]) );
  XOR2_X1 U2068 ( .A(n1386), .B(n68), .Z(product[28]) );
  AOI21_X1 U2069 ( .B1(n106), .B2(n1498), .A(n103), .ZN(n101) );
  OAI21_X1 U2070 ( .B1(n1482), .B2(n107), .A(n108), .ZN(n106) );
  OAI21_X1 U2071 ( .B1(n117), .B2(n115), .A(n116), .ZN(n114) );
  OAI22_X1 U2072 ( .A1(n1363), .A2(n1055), .B1(n1054), .B2(n1357), .ZN(n846)
         );
  OAI22_X1 U2073 ( .A1(n1244), .A2(n1051), .B1(n1050), .B2(n1356), .ZN(n842)
         );
  OAI22_X1 U2074 ( .A1(n1349), .A2(n1062), .B1(n1061), .B2(n1395), .ZN(n853)
         );
  OAI22_X1 U2075 ( .A1(n1349), .A2(n1059), .B1(n1058), .B2(n1395), .ZN(n850)
         );
  OAI22_X1 U2076 ( .A1(n1244), .A2(n1060), .B1(n1059), .B2(n1357), .ZN(n851)
         );
  OAI22_X1 U2077 ( .A1(n1363), .A2(n1053), .B1(n1052), .B2(n1395), .ZN(n844)
         );
  OAI22_X1 U2078 ( .A1(n1364), .A2(n1049), .B1(n1048), .B2(n1357), .ZN(n458)
         );
  OAI22_X1 U2079 ( .A1(n1349), .A2(n1052), .B1(n1051), .B2(n1395), .ZN(n843)
         );
  OAI22_X1 U2080 ( .A1(n1349), .A2(n1063), .B1(n1062), .B2(n1395), .ZN(n854)
         );
  OAI22_X1 U2081 ( .A1(n1363), .A2(n1050), .B1(n1049), .B2(n1357), .ZN(n841)
         );
  OAI22_X1 U2082 ( .A1(n1364), .A2(n1057), .B1(n1056), .B2(n1395), .ZN(n848)
         );
  OAI22_X1 U2083 ( .A1(n1244), .A2(n1065), .B1(n1064), .B2(n1357), .ZN(n856)
         );
  OAI22_X1 U2084 ( .A1(n1349), .A2(n1056), .B1(n1055), .B2(n1395), .ZN(n847)
         );
  OAI22_X1 U2085 ( .A1(n1363), .A2(n1058), .B1(n1057), .B2(n1395), .ZN(n849)
         );
  OAI22_X1 U2086 ( .A1(n1244), .A2(n1148), .B1(n1068), .B2(n1395), .ZN(n678)
         );
  OAI22_X1 U2087 ( .A1(n1244), .A2(n1054), .B1(n1053), .B2(n1395), .ZN(n845)
         );
  OAI22_X1 U2088 ( .A1(n1363), .A2(n1061), .B1(n1060), .B2(n1356), .ZN(n852)
         );
  OAI22_X1 U2089 ( .A1(n1048), .A2(n1364), .B1(n1048), .B2(n1356), .ZN(n664)
         );
  OAI22_X1 U2090 ( .A1(n1364), .A2(n1064), .B1(n1063), .B2(n1356), .ZN(n855)
         );
  OAI22_X1 U2091 ( .A1(n1244), .A2(n1067), .B1(n1066), .B2(n1395), .ZN(n858)
         );
  OAI22_X1 U2092 ( .A1(n1349), .A2(n1066), .B1(n1065), .B2(n1357), .ZN(n857)
         );
  INV_X1 U2093 ( .A(n1357), .ZN(n665) );
endmodule


module mac_7_DW01_add_1 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n34, n35, n36, n37, n38, n39, n40, n41, n43, n45, n46, n47,
         n48, n49, n51, n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65,
         n67, n69, n70, n71, n72, n73, n75, n77, n78, n79, n80, n81, n83, n85,
         n86, n87, n88, n89, n91, n93, n94, n95, n96, n97, n99, n101, n102,
         n103, n104, n105, n107, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n119, n121, n122, n124, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n184, n185, n187, n189, n191,
         n193, n195, n197, n199, n201, n203, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407;

  FA_X1 U8 ( .A(B[33]), .B(A[33]), .CI(n40), .CO(n39), .S(SUM[33]) );
  FA_X1 U9 ( .A(B[32]), .B(A[32]), .CI(n185), .CO(n40), .S(SUM[32]) );
  CLKBUF_X1 U254 ( .A(n115), .Z(n344) );
  OR2_X1 U255 ( .A1(B[0]), .A2(A[0]), .ZN(n345) );
  NAND3_X1 U256 ( .A1(n373), .A2(n374), .A3(n375), .ZN(n346) );
  CLKBUF_X1 U257 ( .A(n39), .Z(n347) );
  CLKBUF_X1 U258 ( .A(n361), .Z(n348) );
  NAND3_X1 U259 ( .A1(n353), .A2(n354), .A3(n355), .ZN(n349) );
  NAND3_X1 U260 ( .A1(n369), .A2(n370), .A3(n371), .ZN(n350) );
  NAND3_X1 U261 ( .A1(n369), .A2(n370), .A3(n371), .ZN(n351) );
  XOR2_X1 U262 ( .A(B[36]), .B(A[36]), .Z(n352) );
  XOR2_X1 U263 ( .A(n351), .B(n352), .Z(SUM[36]) );
  NAND2_X1 U264 ( .A1(n350), .A2(B[36]), .ZN(n353) );
  NAND2_X1 U265 ( .A1(n37), .A2(A[36]), .ZN(n354) );
  NAND2_X1 U266 ( .A1(B[36]), .A2(A[36]), .ZN(n355) );
  NAND3_X1 U267 ( .A1(n353), .A2(n354), .A3(n355), .ZN(n36) );
  CLKBUF_X1 U268 ( .A(n110), .Z(n356) );
  CLKBUF_X1 U269 ( .A(n102), .Z(n357) );
  CLKBUF_X1 U270 ( .A(n62), .Z(n358) );
  CLKBUF_X1 U271 ( .A(n36), .Z(n359) );
  CLKBUF_X1 U272 ( .A(n346), .Z(n360) );
  NAND3_X1 U273 ( .A1(n377), .A2(n378), .A3(n379), .ZN(n361) );
  AOI21_X1 U274 ( .B1(n356), .B2(n395), .A(n107), .ZN(n362) );
  AOI21_X1 U275 ( .B1(n110), .B2(n395), .A(n107), .ZN(n105) );
  AOI21_X1 U276 ( .B1(n357), .B2(n396), .A(n99), .ZN(n363) );
  AOI21_X1 U277 ( .B1(n102), .B2(n396), .A(n99), .ZN(n97) );
  AOI21_X1 U278 ( .B1(n358), .B2(n404), .A(n59), .ZN(n364) );
  AOI21_X1 U279 ( .B1(n62), .B2(n404), .A(n59), .ZN(n57) );
  AOI21_X1 U280 ( .B1(n150), .B2(n114), .A(n344), .ZN(n365) );
  AOI21_X1 U281 ( .B1(n150), .B2(n114), .A(n115), .ZN(n113) );
  NOR2_X1 U282 ( .A1(B[3]), .A2(A[3]), .ZN(n366) );
  AOI21_X1 U283 ( .B1(n130), .B2(n143), .A(n131), .ZN(n367) );
  XOR2_X1 U284 ( .A(B[35]), .B(A[35]), .Z(n368) );
  XOR2_X1 U285 ( .A(n360), .B(n368), .Z(SUM[35]) );
  NAND2_X1 U286 ( .A1(n346), .A2(B[35]), .ZN(n369) );
  NAND2_X1 U287 ( .A1(n38), .A2(A[35]), .ZN(n370) );
  NAND2_X1 U288 ( .A1(B[35]), .A2(A[35]), .ZN(n371) );
  NAND3_X1 U289 ( .A1(n369), .A2(n370), .A3(n371), .ZN(n37) );
  XOR2_X1 U290 ( .A(B[34]), .B(A[34]), .Z(n372) );
  XOR2_X1 U291 ( .A(n347), .B(n372), .Z(SUM[34]) );
  NAND2_X1 U292 ( .A1(n39), .A2(B[34]), .ZN(n373) );
  NAND2_X1 U293 ( .A1(n39), .A2(A[34]), .ZN(n374) );
  NAND2_X1 U294 ( .A1(B[34]), .A2(A[34]), .ZN(n375) );
  NAND3_X1 U295 ( .A1(n373), .A2(n374), .A3(n375), .ZN(n38) );
  XOR2_X1 U296 ( .A(B[37]), .B(A[37]), .Z(n376) );
  XOR2_X1 U297 ( .A(n376), .B(n359), .Z(SUM[37]) );
  NAND2_X1 U298 ( .A1(B[37]), .A2(A[37]), .ZN(n377) );
  NAND2_X1 U299 ( .A1(B[37]), .A2(n349), .ZN(n378) );
  NAND2_X1 U300 ( .A1(A[37]), .A2(n36), .ZN(n379) );
  NAND3_X1 U301 ( .A1(n377), .A2(n378), .A3(n379), .ZN(n35) );
  XOR2_X1 U302 ( .A(B[38]), .B(A[38]), .Z(n380) );
  XOR2_X1 U303 ( .A(n380), .B(n348), .Z(SUM[38]) );
  NAND2_X1 U304 ( .A1(B[38]), .A2(A[38]), .ZN(n381) );
  NAND2_X1 U305 ( .A1(B[38]), .A2(n361), .ZN(n382) );
  NAND2_X1 U306 ( .A1(A[38]), .A2(n35), .ZN(n383) );
  NAND3_X1 U307 ( .A1(n381), .A2(n382), .A3(n383), .ZN(n34) );
  CLKBUF_X1 U308 ( .A(n54), .Z(n384) );
  CLKBUF_X1 U309 ( .A(n94), .Z(n385) );
  CLKBUF_X1 U310 ( .A(n86), .Z(n386) );
  CLKBUF_X1 U311 ( .A(n70), .Z(n387) );
  AOI21_X1 U312 ( .B1(n386), .B2(n401), .A(n83), .ZN(n388) );
  AOI21_X1 U313 ( .B1(n385), .B2(n400), .A(n91), .ZN(n389) );
  NOR2_X2 U314 ( .A1(B[9]), .A2(A[9]), .ZN(n144) );
  CLKBUF_X1 U315 ( .A(n46), .Z(n390) );
  AOI21_X1 U316 ( .B1(n384), .B2(n405), .A(n51), .ZN(n391) );
  CLKBUF_X1 U317 ( .A(n78), .Z(n392) );
  AOI21_X1 U318 ( .B1(n387), .B2(n403), .A(n67), .ZN(n393) );
  AOI21_X1 U319 ( .B1(n392), .B2(n402), .A(n75), .ZN(n394) );
  NOR2_X2 U320 ( .A1(B[11]), .A2(A[11]), .ZN(n132) );
  NOR2_X1 U321 ( .A1(B[7]), .A2(A[7]), .ZN(n155) );
  NOR2_X1 U322 ( .A1(B[8]), .A2(A[8]), .ZN(n147) );
  OR2_X1 U323 ( .A1(B[15]), .A2(A[15]), .ZN(n395) );
  OR2_X1 U324 ( .A1(B[17]), .A2(A[17]), .ZN(n396) );
  OR2_X1 U325 ( .A1(B[13]), .A2(A[13]), .ZN(n399) );
  OR2_X1 U326 ( .A1(B[12]), .A2(A[12]), .ZN(n398) );
  INV_X1 U327 ( .A(n150), .ZN(n149) );
  OAI21_X1 U328 ( .B1(n149), .B2(n140), .A(n141), .ZN(n139) );
  INV_X1 U329 ( .A(n143), .ZN(n141) );
  INV_X1 U330 ( .A(n142), .ZN(n140) );
  NAND2_X1 U331 ( .A1(n142), .A2(n130), .ZN(n128) );
  AOI21_X1 U332 ( .B1(n170), .B2(n161), .A(n162), .ZN(n160) );
  INV_X1 U333 ( .A(n171), .ZN(n170) );
  INV_X1 U334 ( .A(n180), .ZN(n179) );
  INV_X1 U335 ( .A(n85), .ZN(n83) );
  INV_X1 U336 ( .A(n77), .ZN(n75) );
  INV_X1 U337 ( .A(n109), .ZN(n107) );
  INV_X1 U338 ( .A(n101), .ZN(n99) );
  INV_X1 U339 ( .A(n53), .ZN(n51) );
  AOI21_X1 U340 ( .B1(n70), .B2(n403), .A(n67), .ZN(n65) );
  INV_X1 U341 ( .A(n69), .ZN(n67) );
  AOI21_X1 U342 ( .B1(n94), .B2(n400), .A(n91), .ZN(n89) );
  INV_X1 U343 ( .A(n93), .ZN(n91) );
  OAI21_X1 U344 ( .B1(n163), .B2(n169), .A(n164), .ZN(n162) );
  AOI21_X1 U345 ( .B1(n172), .B2(n180), .A(n173), .ZN(n171) );
  NOR2_X1 U346 ( .A1(n177), .A2(n366), .ZN(n172) );
  OAI21_X1 U347 ( .B1(n174), .B2(n178), .A(n175), .ZN(n173) );
  NOR2_X1 U348 ( .A1(n128), .A2(n116), .ZN(n114) );
  NAND2_X1 U349 ( .A1(n398), .A2(n399), .ZN(n116) );
  INV_X1 U350 ( .A(n61), .ZN(n59) );
  OAI21_X1 U351 ( .B1(n144), .B2(n148), .A(n145), .ZN(n143) );
  NOR2_X1 U352 ( .A1(n168), .A2(n163), .ZN(n161) );
  OAI21_X1 U353 ( .B1(n181), .B2(n184), .A(n182), .ZN(n180) );
  NOR2_X1 U354 ( .A1(n137), .A2(n132), .ZN(n130) );
  NAND2_X1 U355 ( .A1(n195), .A2(n80), .ZN(n11) );
  INV_X1 U356 ( .A(n79), .ZN(n195) );
  NAND2_X1 U357 ( .A1(n199), .A2(n96), .ZN(n15) );
  INV_X1 U358 ( .A(n95), .ZN(n199) );
  NAND2_X1 U359 ( .A1(n201), .A2(n104), .ZN(n17) );
  INV_X1 U360 ( .A(n103), .ZN(n201) );
  NOR2_X1 U361 ( .A1(n147), .A2(n144), .ZN(n142) );
  OAI21_X1 U362 ( .B1(n171), .B2(n151), .A(n152), .ZN(n150) );
  NAND2_X1 U363 ( .A1(n161), .A2(n153), .ZN(n151) );
  AOI21_X1 U364 ( .B1(n153), .B2(n162), .A(n154), .ZN(n152) );
  NOR2_X1 U365 ( .A1(n158), .A2(n155), .ZN(n153) );
  AOI21_X1 U366 ( .B1(n130), .B2(n143), .A(n131), .ZN(n129) );
  OAI21_X1 U367 ( .B1(n132), .B2(n138), .A(n133), .ZN(n131) );
  INV_X1 U368 ( .A(n126), .ZN(n124) );
  OAI21_X1 U369 ( .B1(n155), .B2(n159), .A(n156), .ZN(n154) );
  NAND2_X1 U370 ( .A1(n405), .A2(n53), .ZN(n4) );
  AOI21_X1 U371 ( .B1(n399), .B2(n124), .A(n119), .ZN(n117) );
  INV_X1 U372 ( .A(n121), .ZN(n119) );
  NAND2_X1 U373 ( .A1(n187), .A2(n48), .ZN(n3) );
  INV_X1 U374 ( .A(n47), .ZN(n187) );
  NAND2_X1 U375 ( .A1(n189), .A2(n56), .ZN(n5) );
  INV_X1 U376 ( .A(n55), .ZN(n189) );
  NAND2_X1 U377 ( .A1(n193), .A2(n72), .ZN(n9) );
  INV_X1 U378 ( .A(n71), .ZN(n193) );
  NAND2_X1 U379 ( .A1(n406), .A2(n45), .ZN(n2) );
  NAND2_X1 U380 ( .A1(n404), .A2(n61), .ZN(n6) );
  XOR2_X1 U381 ( .A(n393), .B(n7), .Z(SUM[26]) );
  NAND2_X1 U382 ( .A1(n191), .A2(n64), .ZN(n7) );
  INV_X1 U383 ( .A(n63), .ZN(n191) );
  NAND2_X1 U384 ( .A1(n403), .A2(n69), .ZN(n8) );
  NAND2_X1 U385 ( .A1(n402), .A2(n77), .ZN(n10) );
  NAND2_X1 U386 ( .A1(n401), .A2(n85), .ZN(n12) );
  XOR2_X1 U387 ( .A(n389), .B(n13), .Z(SUM[20]) );
  NAND2_X1 U388 ( .A1(n197), .A2(n88), .ZN(n13) );
  INV_X1 U389 ( .A(n87), .ZN(n197) );
  XNOR2_X1 U390 ( .A(n385), .B(n14), .ZN(SUM[19]) );
  NAND2_X1 U391 ( .A1(n400), .A2(n93), .ZN(n14) );
  NAND2_X1 U392 ( .A1(n396), .A2(n101), .ZN(n16) );
  XOR2_X1 U393 ( .A(n122), .B(n20), .Z(SUM[13]) );
  NAND2_X1 U394 ( .A1(n399), .A2(n121), .ZN(n20) );
  AOI21_X1 U395 ( .B1(n127), .B2(n398), .A(n124), .ZN(n122) );
  XNOR2_X1 U396 ( .A(n127), .B(n21), .ZN(SUM[12]) );
  NAND2_X1 U397 ( .A1(n398), .A2(n126), .ZN(n21) );
  XOR2_X1 U398 ( .A(n134), .B(n22), .Z(SUM[11]) );
  NAND2_X1 U399 ( .A1(n206), .A2(n133), .ZN(n22) );
  AOI21_X1 U400 ( .B1(n139), .B2(n207), .A(n136), .ZN(n134) );
  INV_X1 U401 ( .A(n137), .ZN(n207) );
  INV_X1 U402 ( .A(n168), .ZN(n213) );
  XOR2_X1 U403 ( .A(n160), .B(n27), .Z(SUM[6]) );
  NAND2_X1 U404 ( .A1(n211), .A2(n159), .ZN(n27) );
  INV_X1 U405 ( .A(n158), .ZN(n211) );
  XNOR2_X1 U406 ( .A(n146), .B(n24), .ZN(SUM[9]) );
  NAND2_X1 U407 ( .A1(n208), .A2(n145), .ZN(n24) );
  OAI21_X1 U408 ( .B1(n149), .B2(n147), .A(n148), .ZN(n146) );
  INV_X1 U409 ( .A(n138), .ZN(n136) );
  INV_X1 U410 ( .A(n169), .ZN(n167) );
  INV_X1 U411 ( .A(n132), .ZN(n206) );
  INV_X1 U412 ( .A(n144), .ZN(n208) );
  INV_X1 U413 ( .A(n155), .ZN(n210) );
  INV_X1 U414 ( .A(n163), .ZN(n212) );
  INV_X1 U415 ( .A(n366), .ZN(n214) );
  XOR2_X1 U416 ( .A(n165), .B(n28), .Z(SUM[5]) );
  NAND2_X1 U417 ( .A1(n212), .A2(n164), .ZN(n28) );
  AOI21_X1 U418 ( .B1(n170), .B2(n213), .A(n167), .ZN(n165) );
  XNOR2_X1 U419 ( .A(n170), .B(n29), .ZN(SUM[4]) );
  NAND2_X1 U420 ( .A1(n213), .A2(n169), .ZN(n29) );
  XNOR2_X1 U421 ( .A(n176), .B(n30), .ZN(SUM[3]) );
  NAND2_X1 U422 ( .A1(n214), .A2(n175), .ZN(n30) );
  OAI21_X1 U423 ( .B1(n179), .B2(n177), .A(n178), .ZN(n176) );
  XOR2_X1 U424 ( .A(n179), .B(n31), .Z(SUM[2]) );
  NAND2_X1 U425 ( .A1(n215), .A2(n178), .ZN(n31) );
  INV_X1 U426 ( .A(n177), .ZN(n215) );
  XOR2_X1 U427 ( .A(n32), .B(n184), .Z(SUM[1]) );
  NAND2_X1 U428 ( .A1(n216), .A2(n182), .ZN(n32) );
  INV_X1 U429 ( .A(n181), .ZN(n216) );
  AND2_X1 U430 ( .A1(n345), .A2(n184), .ZN(SUM[0]) );
  NAND2_X1 U431 ( .A1(n203), .A2(n112), .ZN(n19) );
  INV_X1 U432 ( .A(n111), .ZN(n203) );
  NAND2_X1 U433 ( .A1(n395), .A2(n109), .ZN(n18) );
  XNOR2_X1 U434 ( .A(n139), .B(n23), .ZN(SUM[10]) );
  NAND2_X1 U435 ( .A1(n207), .A2(n138), .ZN(n23) );
  XOR2_X1 U436 ( .A(n149), .B(n25), .Z(SUM[8]) );
  NAND2_X1 U437 ( .A1(n209), .A2(n148), .ZN(n25) );
  INV_X1 U438 ( .A(n147), .ZN(n209) );
  XNOR2_X1 U439 ( .A(n157), .B(n26), .ZN(SUM[7]) );
  NAND2_X1 U440 ( .A1(n210), .A2(n156), .ZN(n26) );
  OAI21_X1 U441 ( .B1(n160), .B2(n158), .A(n159), .ZN(n157) );
  NOR2_X1 U442 ( .A1(B[6]), .A2(A[6]), .ZN(n158) );
  NOR2_X1 U443 ( .A1(B[2]), .A2(A[2]), .ZN(n177) );
  NOR2_X1 U444 ( .A1(B[5]), .A2(A[5]), .ZN(n163) );
  NOR2_X1 U445 ( .A1(B[3]), .A2(A[3]), .ZN(n174) );
  NOR2_X1 U446 ( .A1(B[10]), .A2(A[10]), .ZN(n137) );
  NOR2_X1 U447 ( .A1(B[4]), .A2(A[4]), .ZN(n168) );
  NOR2_X1 U448 ( .A1(B[1]), .A2(A[1]), .ZN(n181) );
  NAND2_X1 U449 ( .A1(B[8]), .A2(A[8]), .ZN(n148) );
  NAND2_X1 U450 ( .A1(B[6]), .A2(A[6]), .ZN(n159) );
  NAND2_X1 U451 ( .A1(B[2]), .A2(A[2]), .ZN(n178) );
  NAND2_X1 U452 ( .A1(B[0]), .A2(A[0]), .ZN(n184) );
  NAND2_X1 U453 ( .A1(B[10]), .A2(A[10]), .ZN(n138) );
  NAND2_X1 U454 ( .A1(B[4]), .A2(A[4]), .ZN(n169) );
  NAND2_X1 U455 ( .A1(B[11]), .A2(A[11]), .ZN(n133) );
  NAND2_X1 U456 ( .A1(B[9]), .A2(A[9]), .ZN(n145) );
  NAND2_X1 U457 ( .A1(B[5]), .A2(A[5]), .ZN(n164) );
  NAND2_X1 U458 ( .A1(B[7]), .A2(A[7]), .ZN(n156) );
  NAND2_X1 U459 ( .A1(B[3]), .A2(A[3]), .ZN(n175) );
  NAND2_X1 U460 ( .A1(B[1]), .A2(A[1]), .ZN(n182) );
  INV_X1 U461 ( .A(n41), .ZN(n185) );
  INV_X1 U462 ( .A(n45), .ZN(n43) );
  NOR2_X1 U463 ( .A1(B[20]), .A2(A[20]), .ZN(n87) );
  NOR2_X1 U464 ( .A1(B[18]), .A2(A[18]), .ZN(n95) );
  NOR2_X1 U465 ( .A1(B[14]), .A2(A[14]), .ZN(n111) );
  NOR2_X1 U466 ( .A1(B[16]), .A2(A[16]), .ZN(n103) );
  NOR2_X1 U467 ( .A1(B[30]), .A2(A[30]), .ZN(n47) );
  NOR2_X1 U468 ( .A1(B[28]), .A2(A[28]), .ZN(n55) );
  NOR2_X1 U469 ( .A1(B[26]), .A2(A[26]), .ZN(n63) );
  NOR2_X1 U470 ( .A1(B[24]), .A2(A[24]), .ZN(n71) );
  NOR2_X1 U471 ( .A1(B[22]), .A2(A[22]), .ZN(n79) );
  OR2_X1 U472 ( .A1(B[19]), .A2(A[19]), .ZN(n400) );
  NAND2_X1 U473 ( .A1(B[21]), .A2(A[21]), .ZN(n85) );
  NAND2_X1 U474 ( .A1(B[15]), .A2(A[15]), .ZN(n109) );
  NAND2_X1 U475 ( .A1(B[17]), .A2(A[17]), .ZN(n101) );
  NAND2_X1 U476 ( .A1(B[12]), .A2(A[12]), .ZN(n126) );
  NAND2_X1 U477 ( .A1(B[13]), .A2(A[13]), .ZN(n121) );
  NAND2_X1 U478 ( .A1(B[19]), .A2(A[19]), .ZN(n93) );
  NAND2_X1 U479 ( .A1(B[23]), .A2(A[23]), .ZN(n77) );
  NAND2_X1 U480 ( .A1(B[25]), .A2(A[25]), .ZN(n69) );
  NAND2_X1 U481 ( .A1(B[27]), .A2(A[27]), .ZN(n61) );
  NAND2_X1 U482 ( .A1(B[29]), .A2(A[29]), .ZN(n53) );
  NAND2_X1 U483 ( .A1(B[31]), .A2(A[31]), .ZN(n45) );
  NAND2_X1 U484 ( .A1(B[20]), .A2(A[20]), .ZN(n88) );
  NAND2_X1 U485 ( .A1(B[18]), .A2(A[18]), .ZN(n96) );
  NAND2_X1 U486 ( .A1(B[14]), .A2(A[14]), .ZN(n112) );
  NAND2_X1 U487 ( .A1(B[16]), .A2(A[16]), .ZN(n104) );
  NAND2_X1 U488 ( .A1(B[30]), .A2(A[30]), .ZN(n48) );
  NAND2_X1 U489 ( .A1(B[28]), .A2(A[28]), .ZN(n56) );
  NAND2_X1 U490 ( .A1(B[26]), .A2(A[26]), .ZN(n64) );
  NAND2_X1 U491 ( .A1(B[24]), .A2(A[24]), .ZN(n72) );
  NAND2_X1 U492 ( .A1(B[22]), .A2(A[22]), .ZN(n80) );
  OR2_X1 U493 ( .A1(B[21]), .A2(A[21]), .ZN(n401) );
  OR2_X1 U494 ( .A1(B[23]), .A2(A[23]), .ZN(n402) );
  OR2_X1 U495 ( .A1(B[25]), .A2(A[25]), .ZN(n403) );
  OR2_X1 U496 ( .A1(B[27]), .A2(A[27]), .ZN(n404) );
  OR2_X1 U497 ( .A1(B[29]), .A2(A[29]), .ZN(n405) );
  OR2_X1 U498 ( .A1(B[31]), .A2(A[31]), .ZN(n406) );
  XNOR2_X1 U499 ( .A(n34), .B(n407), .ZN(SUM[39]) );
  XNOR2_X1 U500 ( .A(A[39]), .B(B[39]), .ZN(n407) );
  OAI21_X1 U501 ( .B1(n97), .B2(n95), .A(n96), .ZN(n94) );
  XOR2_X1 U502 ( .A(n363), .B(n15), .Z(SUM[18]) );
  XNOR2_X1 U503 ( .A(n357), .B(n16), .ZN(SUM[17]) );
  XNOR2_X1 U504 ( .A(n386), .B(n12), .ZN(SUM[21]) );
  AOI21_X1 U505 ( .B1(n86), .B2(n401), .A(n83), .ZN(n81) );
  AOI21_X1 U506 ( .B1(n78), .B2(n402), .A(n75), .ZN(n73) );
  XNOR2_X1 U507 ( .A(n392), .B(n10), .ZN(SUM[23]) );
  OAI21_X1 U508 ( .B1(n89), .B2(n87), .A(n88), .ZN(n86) );
  OAI21_X1 U509 ( .B1(n113), .B2(n111), .A(n112), .ZN(n110) );
  XNOR2_X1 U510 ( .A(n356), .B(n18), .ZN(SUM[15]) );
  XNOR2_X1 U511 ( .A(n387), .B(n8), .ZN(SUM[25]) );
  XOR2_X1 U512 ( .A(n364), .B(n5), .Z(SUM[28]) );
  OAI21_X1 U513 ( .B1(n149), .B2(n128), .A(n367), .ZN(n127) );
  OAI21_X1 U514 ( .B1(n129), .B2(n116), .A(n117), .ZN(n115) );
  XNOR2_X1 U515 ( .A(n384), .B(n4), .ZN(SUM[29]) );
  XNOR2_X1 U516 ( .A(n358), .B(n6), .ZN(SUM[27]) );
  XOR2_X1 U517 ( .A(n362), .B(n17), .Z(SUM[16]) );
  XOR2_X1 U518 ( .A(n394), .B(n9), .Z(SUM[24]) );
  OAI21_X1 U519 ( .B1(n73), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U520 ( .B1(n65), .B2(n63), .A(n64), .ZN(n62) );
  OAI21_X1 U521 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  OAI21_X1 U522 ( .B1(n105), .B2(n103), .A(n104), .ZN(n102) );
  AOI21_X1 U523 ( .B1(n54), .B2(n405), .A(n51), .ZN(n49) );
  XNOR2_X1 U524 ( .A(n390), .B(n2), .ZN(SUM[31]) );
  XOR2_X1 U525 ( .A(n365), .B(n19), .Z(SUM[14]) );
  XOR2_X1 U526 ( .A(n388), .B(n11), .Z(SUM[22]) );
  XOR2_X1 U527 ( .A(n391), .B(n3), .Z(SUM[30]) );
  AOI21_X1 U528 ( .B1(n46), .B2(n406), .A(n43), .ZN(n41) );
  OAI21_X1 U529 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  OAI21_X1 U530 ( .B1(n81), .B2(n79), .A(n80), .ZN(n78) );
endmodule


module mac_7 ( clk, clear_acc, a, b, mac_out );
  input [19:0] a;
  input [19:0] b;
  output [39:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, n2, n3;
  wire   [39:0] mul;
  wire   [39:0] pipeline;
  wire   [39:0] sum;

  DFF_X1 \pipeline_reg[39]  ( .D(mul[39]), .CK(clk), .Q(pipeline[39]) );
  DFF_X1 \pipeline_reg[38]  ( .D(mul[38]), .CK(clk), .Q(pipeline[38]) );
  DFF_X1 \pipeline_reg[37]  ( .D(mul[37]), .CK(clk), .Q(pipeline[37]) );
  DFF_X1 \pipeline_reg[36]  ( .D(mul[36]), .CK(clk), .Q(pipeline[36]) );
  DFF_X1 \pipeline_reg[35]  ( .D(mul[35]), .CK(clk), .Q(pipeline[35]) );
  DFF_X1 \pipeline_reg[34]  ( .D(mul[34]), .CK(clk), .Q(pipeline[34]) );
  DFF_X1 \pipeline_reg[33]  ( .D(mul[33]), .CK(clk), .Q(pipeline[33]) );
  DFF_X1 \pipeline_reg[32]  ( .D(mul[32]), .CK(clk), .Q(pipeline[32]) );
  DFF_X1 \pipeline_reg[31]  ( .D(mul[31]), .CK(clk), .Q(pipeline[31]) );
  DFF_X1 \pipeline_reg[30]  ( .D(mul[30]), .CK(clk), .Q(pipeline[30]) );
  DFF_X1 \pipeline_reg[29]  ( .D(mul[29]), .CK(clk), .Q(pipeline[29]) );
  DFF_X1 \pipeline_reg[28]  ( .D(mul[28]), .CK(clk), .Q(pipeline[28]) );
  DFF_X1 \pipeline_reg[27]  ( .D(mul[27]), .CK(clk), .Q(pipeline[27]) );
  DFF_X1 \pipeline_reg[26]  ( .D(mul[26]), .CK(clk), .Q(pipeline[26]) );
  DFF_X1 \pipeline_reg[25]  ( .D(mul[25]), .CK(clk), .Q(pipeline[25]) );
  DFF_X1 \pipeline_reg[24]  ( .D(mul[24]), .CK(clk), .Q(pipeline[24]) );
  DFF_X1 \pipeline_reg[23]  ( .D(mul[23]), .CK(clk), .Q(pipeline[23]) );
  DFF_X1 \pipeline_reg[22]  ( .D(mul[22]), .CK(clk), .Q(pipeline[22]) );
  DFF_X1 \pipeline_reg[21]  ( .D(mul[21]), .CK(clk), .Q(pipeline[21]) );
  DFF_X1 \pipeline_reg[20]  ( .D(mul[20]), .CK(clk), .Q(pipeline[20]) );
  DFF_X1 \pipeline_reg[19]  ( .D(mul[19]), .CK(clk), .Q(pipeline[19]) );
  DFF_X1 \pipeline_reg[18]  ( .D(mul[18]), .CK(clk), .Q(pipeline[18]) );
  DFF_X1 \pipeline_reg[17]  ( .D(mul[17]), .CK(clk), .Q(pipeline[17]) );
  DFF_X1 \pipeline_reg[16]  ( .D(mul[16]), .CK(clk), .Q(pipeline[16]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \mac_out_reg[17]  ( .D(N20), .CK(clk), .Q(mac_out[17]) );
  DFF_X1 \mac_out_reg[18]  ( .D(N21), .CK(clk), .Q(mac_out[18]) );
  DFF_X1 \mac_out_reg[19]  ( .D(N22), .CK(clk), .Q(mac_out[19]) );
  DFF_X1 \mac_out_reg[20]  ( .D(N23), .CK(clk), .Q(mac_out[20]) );
  DFF_X1 \mac_out_reg[21]  ( .D(N24), .CK(clk), .Q(mac_out[21]) );
  DFF_X1 \mac_out_reg[22]  ( .D(N25), .CK(clk), .Q(mac_out[22]) );
  DFF_X1 \mac_out_reg[23]  ( .D(N26), .CK(clk), .Q(mac_out[23]) );
  DFF_X1 \mac_out_reg[24]  ( .D(N27), .CK(clk), .Q(mac_out[24]) );
  DFF_X1 \mac_out_reg[25]  ( .D(N28), .CK(clk), .Q(mac_out[25]) );
  DFF_X1 \mac_out_reg[26]  ( .D(N29), .CK(clk), .Q(mac_out[26]) );
  DFF_X1 \mac_out_reg[27]  ( .D(N30), .CK(clk), .Q(mac_out[27]) );
  DFF_X1 \mac_out_reg[28]  ( .D(N31), .CK(clk), .Q(mac_out[28]) );
  DFF_X1 \mac_out_reg[29]  ( .D(N32), .CK(clk), .Q(mac_out[29]) );
  DFF_X1 \mac_out_reg[30]  ( .D(N33), .CK(clk), .Q(mac_out[30]) );
  DFF_X1 \mac_out_reg[31]  ( .D(N34), .CK(clk), .Q(mac_out[31]) );
  DFF_X1 \mac_out_reg[32]  ( .D(N35), .CK(clk), .Q(mac_out[32]) );
  DFF_X1 \mac_out_reg[33]  ( .D(N36), .CK(clk), .Q(mac_out[33]) );
  DFF_X1 \mac_out_reg[34]  ( .D(N37), .CK(clk), .Q(mac_out[34]) );
  DFF_X1 \mac_out_reg[35]  ( .D(N38), .CK(clk), .Q(mac_out[35]) );
  DFF_X1 \mac_out_reg[36]  ( .D(N39), .CK(clk), .Q(mac_out[36]) );
  DFF_X1 \mac_out_reg[37]  ( .D(N40), .CK(clk), .Q(mac_out[37]) );
  DFF_X1 \mac_out_reg[38]  ( .D(N41), .CK(clk), .Q(mac_out[38]) );
  DFF_X1 \mac_out_reg[39]  ( .D(N42), .CK(clk), .Q(mac_out[39]) );
  mac_7_DW_mult_tc_1 mult_355 ( .a(a), .b(b), .product(mul) );
  mac_7_DW01_add_1 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \mac_out_reg[16]  ( .D(N19), .CK(clk), .Q(mac_out[16]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  BUF_X1 U3 ( .A(n3), .Z(n2) );
  INV_X1 U4 ( .A(clear_acc), .ZN(n3) );
  AND2_X1 U6 ( .A1(sum[39]), .A2(n2), .ZN(N42) );
  AND2_X1 U7 ( .A1(sum[38]), .A2(n2), .ZN(N41) );
  AND2_X1 U8 ( .A1(sum[37]), .A2(n2), .ZN(N40) );
  AND2_X1 U9 ( .A1(sum[36]), .A2(n2), .ZN(N39) );
  AND2_X1 U10 ( .A1(sum[35]), .A2(n2), .ZN(N38) );
  AND2_X1 U11 ( .A1(sum[34]), .A2(n2), .ZN(N37) );
  AND2_X1 U12 ( .A1(sum[33]), .A2(n2), .ZN(N36) );
  AND2_X1 U13 ( .A1(sum[32]), .A2(n2), .ZN(N35) );
  AND2_X1 U14 ( .A1(sum[31]), .A2(n2), .ZN(N34) );
  AND2_X1 U15 ( .A1(sum[30]), .A2(n2), .ZN(N33) );
  AND2_X1 U16 ( .A1(sum[29]), .A2(n2), .ZN(N32) );
  AND2_X1 U17 ( .A1(sum[28]), .A2(n3), .ZN(N31) );
  AND2_X1 U18 ( .A1(sum[27]), .A2(n3), .ZN(N30) );
  AND2_X1 U19 ( .A1(sum[26]), .A2(n3), .ZN(N29) );
  AND2_X1 U20 ( .A1(sum[25]), .A2(n3), .ZN(N28) );
  AND2_X1 U21 ( .A1(sum[24]), .A2(n3), .ZN(N27) );
  AND2_X1 U22 ( .A1(sum[23]), .A2(n3), .ZN(N26) );
  AND2_X1 U23 ( .A1(sum[22]), .A2(n3), .ZN(N25) );
  AND2_X1 U24 ( .A1(sum[21]), .A2(n3), .ZN(N24) );
  AND2_X1 U25 ( .A1(sum[20]), .A2(n3), .ZN(N23) );
  AND2_X1 U26 ( .A1(sum[19]), .A2(n3), .ZN(N22) );
  AND2_X1 U27 ( .A1(sum[18]), .A2(n3), .ZN(N21) );
  AND2_X1 U28 ( .A1(sum[17]), .A2(n3), .ZN(N20) );
  AND2_X1 U29 ( .A1(sum[16]), .A2(n3), .ZN(N19) );
  AND2_X1 U30 ( .A1(sum[15]), .A2(n3), .ZN(N18) );
  AND2_X1 U31 ( .A1(sum[14]), .A2(n3), .ZN(N17) );
  AND2_X1 U32 ( .A1(sum[13]), .A2(n3), .ZN(N16) );
  AND2_X1 U33 ( .A1(sum[12]), .A2(n3), .ZN(N15) );
  AND2_X1 U34 ( .A1(sum[11]), .A2(n3), .ZN(N14) );
  AND2_X1 U35 ( .A1(sum[10]), .A2(n3), .ZN(N13) );
  AND2_X1 U36 ( .A1(sum[9]), .A2(n3), .ZN(N12) );
  AND2_X1 U37 ( .A1(sum[8]), .A2(n3), .ZN(N11) );
  AND2_X1 U38 ( .A1(sum[7]), .A2(n3), .ZN(N10) );
  AND2_X1 U39 ( .A1(sum[6]), .A2(n3), .ZN(N9) );
  AND2_X1 U40 ( .A1(sum[5]), .A2(n3), .ZN(N8) );
  AND2_X1 U41 ( .A1(sum[4]), .A2(n3), .ZN(N7) );
  AND2_X1 U42 ( .A1(sum[3]), .A2(n3), .ZN(N6) );
  AND2_X1 U43 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U44 ( .A1(sum[1]), .A2(n3), .ZN(N4) );
  AND2_X1 U45 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
endmodule


module mac_6_DW_mult_tc_1 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n6, n7, n9, n12, n13, n18, n19, n22, n24, n25, n28, n30, n31, n34,
         n36, n37, n40, n43, n46, n48, n49, n52, n54, n55, n60, n61, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n97, n98, n99, n100, n101, n103, n105, n106, n107, n108,
         n109, n111, n113, n114, n115, n116, n117, n119, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n185, n186, n187, n188, n193, n194, n195, n196, n200, n201,
         n202, n203, n204, n205, n206, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n225,
         n227, n228, n230, n232, n233, n234, n236, n238, n239, n240, n241,
         n242, n244, n246, n247, n248, n249, n250, n252, n254, n255, n256,
         n257, n258, n259, n260, n261, n263, n264, n266, n268, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n284, n285,
         n286, n287, n291, n293, n295, n296, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n643, n646,
         n647, n649, n650, n652, n653, n655, n656, n658, n659, n661, n662,
         n664, n665, n667, n668, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1113, n1140, n1141, n1142, n1143, n1144, n1145, n1147,
         n1148, n1149, n1233, n1234, n1235, n1236, n1237, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n37 = a[13];
  assign n43 = a[15];
  assign n49 = a[17];
  assign n55 = a[19];
  assign n61 = b[0];
  assign n668 = a[0];
  assign n1090 = b[19];
  assign n1091 = b[18];
  assign n1092 = b[17];
  assign n1093 = b[16];
  assign n1094 = b[15];
  assign n1095 = b[14];
  assign n1096 = b[13];
  assign n1097 = b[12];
  assign n1098 = b[11];
  assign n1099 = b[10];
  assign n1100 = b[9];
  assign n1101 = b[8];
  assign n1102 = b[7];
  assign n1103 = b[6];
  assign n1104 = b[5];
  assign n1105 = b[4];
  assign n1106 = b[3];
  assign n1107 = b[2];
  assign n1108 = b[1];

  FA_X1 U333 ( .A(n681), .B(n304), .CI(n700), .CO(n300), .S(n301) );
  FA_X1 U334 ( .A(n305), .B(n682), .CI(n308), .CO(n302), .S(n303) );
  FA_X1 U336 ( .A(n312), .B(n683), .CI(n309), .CO(n306), .S(n307) );
  FA_X1 U337 ( .A(n701), .B(n314), .CI(n720), .CO(n308), .S(n309) );
  FA_X1 U338 ( .A(n313), .B(n320), .CI(n318), .CO(n310), .S(n311) );
  FA_X1 U339 ( .A(n684), .B(n702), .CI(n315), .CO(n312), .S(n313) );
  FA_X1 U341 ( .A(n324), .B(n321), .CI(n319), .CO(n316), .S(n317) );
  FA_X1 U342 ( .A(n328), .B(n721), .CI(n326), .CO(n318), .S(n319) );
  FA_X1 U343 ( .A(n703), .B(n685), .CI(n740), .CO(n320), .S(n321) );
  FA_X1 U344 ( .A(n325), .B(n327), .CI(n332), .CO(n322), .S(n323) );
  FA_X1 U345 ( .A(n336), .B(n329), .CI(n334), .CO(n324), .S(n325) );
  FA_X1 U346 ( .A(n686), .B(n704), .CI(n722), .CO(n326), .S(n327) );
  FA_X1 U348 ( .A(n340), .B(n342), .CI(n333), .CO(n330), .S(n331) );
  FA_X1 U349 ( .A(n335), .B(n344), .CI(n337), .CO(n332), .S(n333) );
  FA_X1 U350 ( .A(n705), .B(n346), .CI(n723), .CO(n334), .S(n335) );
  FA_X1 U351 ( .A(n741), .B(n687), .CI(n760), .CO(n336), .S(n337) );
  FA_X1 U352 ( .A(n350), .B(n343), .CI(n341), .CO(n338), .S(n339) );
  FA_X1 U353 ( .A(n345), .B(n354), .CI(n352), .CO(n340), .S(n341) );
  FA_X1 U354 ( .A(n347), .B(n724), .CI(n356), .CO(n342), .S(n343) );
  FA_X1 U355 ( .A(n742), .B(n706), .CI(n688), .CO(n344), .S(n345) );
  FA_X1 U357 ( .A(n360), .B(n353), .CI(n351), .CO(n348), .S(n349) );
  FA_X1 U358 ( .A(n357), .B(n355), .CI(n362), .CO(n350), .S(n351) );
  FA_X1 U359 ( .A(n366), .B(n743), .CI(n364), .CO(n352), .S(n353) );
  FA_X1 U360 ( .A(n707), .B(n761), .CI(n725), .CO(n354), .S(n355) );
  FA_X1 U361 ( .A(n368), .B(n689), .CI(n780), .CO(n356), .S(n357) );
  FA_X1 U362 ( .A(n372), .B(n363), .CI(n361), .CO(n358), .S(n359) );
  FA_X1 U363 ( .A(n376), .B(n365), .CI(n374), .CO(n360), .S(n361) );
  FA_X1 U364 ( .A(n378), .B(n380), .CI(n367), .CO(n362), .S(n363) );
  FA_X1 U365 ( .A(n690), .B(n708), .CI(n369), .CO(n364), .S(n365) );
  FA_X1 U366 ( .A(n762), .B(n726), .CI(n744), .CO(n366), .S(n367) );
  FA_X1 U368 ( .A(n384), .B(n375), .CI(n373), .CO(n370), .S(n371) );
  FA_X1 U369 ( .A(n377), .B(n388), .CI(n386), .CO(n372), .S(n373) );
  FA_X1 U370 ( .A(n379), .B(n390), .CI(n381), .CO(n374), .S(n375) );
  FA_X1 U371 ( .A(n727), .B(n745), .CI(n392), .CO(n376), .S(n377) );
  FA_X1 U372 ( .A(n709), .B(n781), .CI(n763), .CO(n378), .S(n379) );
  FA_X1 U373 ( .A(n394), .B(n691), .CI(n800), .CO(n380), .S(n381) );
  FA_X1 U374 ( .A(n398), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U375 ( .A(n389), .B(n402), .CI(n400), .CO(n384), .S(n385) );
  FA_X1 U376 ( .A(n393), .B(n404), .CI(n391), .CO(n386), .S(n387) );
  FA_X1 U377 ( .A(n408), .B(n395), .CI(n406), .CO(n388), .S(n389) );
  FA_X1 U378 ( .A(n746), .B(n782), .CI(n764), .CO(n390), .S(n391) );
  FA_X1 U379 ( .A(n692), .B(n728), .CI(n710), .CO(n392), .S(n393) );
  FA_X1 U381 ( .A(n401), .B(n412), .CI(n399), .CO(n396), .S(n397) );
  FA_X1 U382 ( .A(n414), .B(n416), .CI(n403), .CO(n398), .S(n399) );
  FA_X1 U384 ( .A(n420), .B(n422), .CI(n405), .CO(n402), .S(n403) );
  FA_X1 U385 ( .A(n729), .B(n765), .CI(n747), .CO(n404), .S(n405) );
  FA_X1 U386 ( .A(n711), .B(n783), .CI(n801), .CO(n406), .S(n407) );
  FA_X1 U388 ( .A(n428), .B(n415), .CI(n413), .CO(n410), .S(n411) );
  FA_X1 U389 ( .A(n417), .B(n432), .CI(n430), .CO(n412), .S(n413) );
  FA_X1 U391 ( .A(n436), .B(n438), .CI(n421), .CO(n416), .S(n417) );
  FA_X1 U393 ( .A(n694), .B(n766), .CI(n712), .CO(n420), .S(n421) );
  FA_X1 U394 ( .A(n802), .B(n730), .CI(n784), .CO(n422), .S(n423) );
  FA_X1 U397 ( .A(n433), .B(n448), .CI(n446), .CO(n428), .S(n429) );
  FA_X1 U399 ( .A(n437), .B(n452), .CI(n439), .CO(n432), .S(n433) );
  FA_X1 U400 ( .A(n767), .B(n456), .CI(n454), .CO(n434), .S(n435) );
  FA_X1 U401 ( .A(n731), .B(n785), .CI(n749), .CO(n436), .S(n437) );
  FA_X1 U402 ( .A(n713), .B(n803), .CI(n458), .CO(n438), .S(n439) );
  FA_X1 U403 ( .A(n821), .B(n695), .CI(n840), .CO(n440), .S(n441) );
  FA_X1 U404 ( .A(n462), .B(n447), .CI(n445), .CO(n442), .S(n443) );
  FA_X1 U405 ( .A(n449), .B(n466), .CI(n464), .CO(n444), .S(n445) );
  FA_X1 U406 ( .A(n468), .B(n453), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U407 ( .A(n455), .B(n470), .CI(n457), .CO(n448), .S(n449) );
  FA_X1 U408 ( .A(n474), .B(n476), .CI(n472), .CO(n450), .S(n451) );
  FA_X1 U409 ( .A(n768), .B(n786), .CI(n459), .CO(n452), .S(n453) );
  FA_X1 U410 ( .A(n804), .B(n732), .CI(n714), .CO(n454), .S(n455) );
  FA_X1 U411 ( .A(n750), .B(n696), .CI(n822), .CO(n456), .S(n457) );
  FA_X1 U416 ( .A(n473), .B(n488), .CI(n475), .CO(n466), .S(n467) );
  FA_X1 U417 ( .A(n490), .B(n477), .CI(n492), .CO(n468), .S(n469) );
  FA_X1 U418 ( .A(n805), .B(n823), .CI(n494), .CO(n470), .S(n471) );
  FA_X1 U419 ( .A(n751), .B(n841), .CI(n733), .CO(n472), .S(n473) );
  FA_X1 U423 ( .A(n498), .B(n483), .CI(n481), .CO(n478), .S(n479) );
  FA_X1 U424 ( .A(n500), .B(n487), .CI(n485), .CO(n480), .S(n481) );
  FA_X1 U426 ( .A(n489), .B(n506), .CI(n491), .CO(n484), .S(n485) );
  FA_X1 U428 ( .A(n770), .B(n824), .CI(n842), .CO(n488), .S(n489) );
  FA_X1 U429 ( .A(n861), .B(n752), .CI(n806), .CO(n490), .S(n491) );
  FA_X1 U430 ( .A(n788), .B(n670), .CI(n734), .CO(n492), .S(n493) );
  HA_X1 U431 ( .A(n716), .B(n698), .CO(n494), .S(n495) );
  FA_X1 U433 ( .A(n516), .B(n505), .CI(n503), .CO(n498), .S(n499) );
  FA_X1 U434 ( .A(n520), .B(n509), .CI(n518), .CO(n500), .S(n501) );
  FA_X1 U436 ( .A(n526), .B(n807), .CI(n524), .CO(n504), .S(n505) );
  FA_X1 U437 ( .A(n771), .B(n825), .CI(n789), .CO(n506), .S(n507) );
  FA_X1 U438 ( .A(n717), .B(n753), .CI(n843), .CO(n508), .S(n509) );
  FA_X1 U439 ( .A(n735), .B(n699), .CI(n862), .CO(n510), .S(n511) );
  FA_X1 U440 ( .A(n517), .B(n530), .CI(n515), .CO(n512), .S(n513) );
  FA_X1 U441 ( .A(n519), .B(n521), .CI(n532), .CO(n514), .S(n515) );
  FA_X1 U443 ( .A(n536), .B(n540), .CI(n538), .CO(n518), .S(n519) );
  FA_X1 U444 ( .A(n826), .B(n844), .CI(n527), .CO(n520), .S(n521) );
  FA_X1 U445 ( .A(n754), .B(n772), .CI(n808), .CO(n522), .S(n523) );
  FA_X1 U446 ( .A(n863), .B(n790), .CI(n671), .CO(n524), .S(n525) );
  HA_X1 U447 ( .A(n718), .B(n736), .CO(n526), .S(n527) );
  FA_X1 U449 ( .A(n535), .B(n548), .CI(n546), .CO(n530), .S(n531) );
  FA_X1 U451 ( .A(n552), .B(n554), .CI(n550), .CO(n534), .S(n535) );
  FA_X1 U453 ( .A(n737), .B(n773), .CI(n845), .CO(n538), .S(n539) );
  FA_X1 U454 ( .A(n755), .B(n719), .CI(n864), .CO(n540), .S(n541) );
  FA_X1 U456 ( .A(n560), .B(n553), .CI(n549), .CO(n544), .S(n545) );
  FA_X1 U458 ( .A(n555), .B(n846), .CI(n566), .CO(n548), .S(n549) );
  FA_X1 U459 ( .A(n865), .B(n828), .CI(n792), .CO(n550), .S(n551) );
  HA_X1 U461 ( .A(n738), .B(n756), .CO(n554), .S(n555) );
  FA_X1 U462 ( .A(n561), .B(n570), .CI(n559), .CO(n556), .S(n557) );
  FA_X1 U463 ( .A(n563), .B(n565), .CI(n572), .CO(n558), .S(n559) );
  FA_X1 U466 ( .A(n757), .B(n847), .CI(n793), .CO(n564), .S(n565) );
  FA_X1 U467 ( .A(n866), .B(n739), .CI(n775), .CO(n566), .S(n567) );
  FA_X1 U468 ( .A(n582), .B(n573), .CI(n571), .CO(n568), .S(n569) );
  FA_X1 U469 ( .A(n577), .B(n575), .CI(n584), .CO(n570), .S(n571) );
  FA_X1 U470 ( .A(n588), .B(n579), .CI(n586), .CO(n572), .S(n573) );
  FA_X1 U471 ( .A(n848), .B(n830), .CI(n794), .CO(n574), .S(n575) );
  FA_X1 U472 ( .A(n867), .B(n812), .CI(n673), .CO(n576), .S(n577) );
  HA_X1 U473 ( .A(n758), .B(n776), .CO(n578), .S(n579) );
  FA_X1 U474 ( .A(n585), .B(n592), .CI(n583), .CO(n580), .S(n581) );
  FA_X1 U475 ( .A(n587), .B(n589), .CI(n594), .CO(n582), .S(n583) );
  FA_X1 U476 ( .A(n598), .B(n831), .CI(n596), .CO(n584), .S(n585) );
  FA_X1 U477 ( .A(n777), .B(n849), .CI(n813), .CO(n586), .S(n587) );
  FA_X1 U478 ( .A(n868), .B(n759), .CI(n795), .CO(n588), .S(n589) );
  FA_X1 U479 ( .A(n602), .B(n595), .CI(n593), .CO(n590), .S(n591) );
  FA_X1 U480 ( .A(n604), .B(n606), .CI(n597), .CO(n592), .S(n593) );
  FA_X1 U481 ( .A(n814), .B(n850), .CI(n599), .CO(n594), .S(n595) );
  FA_X1 U482 ( .A(n869), .B(n832), .CI(n674), .CO(n596), .S(n597) );
  HA_X1 U483 ( .A(n796), .B(n778), .CO(n598), .S(n599) );
  FA_X1 U485 ( .A(n612), .B(n614), .CI(n607), .CO(n602), .S(n603) );
  FA_X1 U486 ( .A(n797), .B(n851), .CI(n833), .CO(n604), .S(n605) );
  FA_X1 U487 ( .A(n815), .B(n870), .CI(n779), .CO(n606), .S(n607) );
  FA_X1 U488 ( .A(n613), .B(n618), .CI(n611), .CO(n608), .S(n609) );
  FA_X1 U489 ( .A(n615), .B(n871), .CI(n620), .CO(n610), .S(n611) );
  FA_X1 U490 ( .A(n852), .B(n834), .CI(n675), .CO(n612), .S(n613) );
  HA_X1 U491 ( .A(n816), .B(n798), .CO(n614), .S(n615) );
  FA_X1 U492 ( .A(n621), .B(n624), .CI(n619), .CO(n616), .S(n617) );
  FA_X1 U493 ( .A(n817), .B(n853), .CI(n626), .CO(n618), .S(n619) );
  FA_X1 U494 ( .A(n835), .B(n799), .CI(n872), .CO(n620), .S(n621) );
  FA_X1 U495 ( .A(n630), .B(n627), .CI(n625), .CO(n622), .S(n623) );
  FA_X1 U496 ( .A(n854), .B(n873), .CI(n676), .CO(n624), .S(n625) );
  HA_X1 U497 ( .A(n818), .B(n836), .CO(n626), .S(n627) );
  FA_X1 U498 ( .A(n634), .B(n837), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U499 ( .A(n874), .B(n819), .CI(n855), .CO(n630), .S(n631) );
  FA_X1 U500 ( .A(n677), .B(n856), .CI(n635), .CO(n632), .S(n633) );
  HA_X1 U501 ( .A(n838), .B(n875), .CO(n634), .S(n635) );
  FA_X1 U502 ( .A(n876), .B(n839), .CI(n857), .CO(n636), .S(n637) );
  HA_X1 U503 ( .A(n858), .B(n877), .CO(n638), .S(n639) );
  CLKBUF_X3 U1025 ( .A(n1356), .Z(n1528) );
  CLKBUF_X3 U1026 ( .A(n1356), .Z(n1334) );
  CLKBUF_X3 U1027 ( .A(n48), .Z(n1370) );
  CLKBUF_X1 U1028 ( .A(n465), .Z(n1233) );
  BUF_X2 U1029 ( .A(n25), .Z(n1544) );
  BUF_X2 U1030 ( .A(n46), .Z(n1524) );
  BUF_X2 U1031 ( .A(n28), .Z(n1428) );
  CLKBUF_X2 U1032 ( .A(n1097), .Z(n1560) );
  BUF_X2 U1033 ( .A(n37), .Z(n1303) );
  XNOR2_X1 U1034 ( .A(n1345), .B(n1303), .ZN(n1234) );
  BUF_X2 U1035 ( .A(n1105), .Z(n1552) );
  CLKBUF_X1 U1036 ( .A(n165), .Z(n1235) );
  AND2_X1 U1037 ( .A1(n529), .A2(n542), .ZN(n1440) );
  INV_X1 U1038 ( .A(n1440), .ZN(n188) );
  BUF_X1 U1039 ( .A(n1102), .Z(n1345) );
  BUF_X2 U1040 ( .A(n13), .Z(n1418) );
  BUF_X2 U1041 ( .A(n1103), .Z(n1554) );
  BUF_X1 U1042 ( .A(n1099), .Z(n1311) );
  BUF_X2 U1043 ( .A(n1103), .Z(n1305) );
  BUF_X1 U1044 ( .A(n1102), .Z(n1555) );
  BUF_X2 U1045 ( .A(n1098), .Z(n1559) );
  BUF_X1 U1046 ( .A(n48), .Z(n1369) );
  BUF_X2 U1047 ( .A(n1101), .Z(n1556) );
  BUF_X2 U1048 ( .A(n1494), .Z(n1338) );
  BUF_X2 U1049 ( .A(n1107), .Z(n1550) );
  NAND3_X1 U1050 ( .A1(n1411), .A2(n1412), .A3(n1413), .ZN(n562) );
  NAND3_X1 U1051 ( .A1(n1377), .A2(n1378), .A3(n1379), .ZN(n486) );
  BUF_X2 U1052 ( .A(n30), .Z(n1463) );
  BUF_X2 U1053 ( .A(n1464), .Z(n1445) );
  BUF_X2 U1054 ( .A(n1095), .Z(n1562) );
  BUF_X1 U1055 ( .A(n1093), .Z(n1564) );
  BUF_X1 U1056 ( .A(n49), .Z(n1546) );
  BUF_X1 U1057 ( .A(n1091), .Z(n1566) );
  BUF_X2 U1058 ( .A(n1), .Z(n1335) );
  BUF_X2 U1059 ( .A(n7), .Z(n1293) );
  XOR2_X1 U1060 ( .A(n1384), .B(n537), .Z(n533) );
  BUF_X2 U1061 ( .A(n1094), .Z(n1563) );
  BUF_X2 U1062 ( .A(n1), .Z(n1543) );
  INV_X1 U1063 ( .A(n298), .ZN(n299) );
  INV_X1 U1064 ( .A(n1459), .ZN(n200) );
  INV_X1 U1065 ( .A(n1295), .ZN(n185) );
  CLKBUF_X1 U1066 ( .A(n133), .Z(n1236) );
  BUF_X2 U1067 ( .A(n1106), .Z(n1551) );
  OR2_X1 U1068 ( .A1(n679), .A2(n879), .ZN(n1237) );
  AND2_X1 U1069 ( .A1(n1237), .A2(n263), .ZN(product[1]) );
  XNOR2_X1 U1070 ( .A(n1311), .B(n1365), .ZN(n1239) );
  XNOR2_X1 U1071 ( .A(n482), .B(n1240), .ZN(n463) );
  XNOR2_X1 U1072 ( .A(n484), .B(n467), .ZN(n1240) );
  CLKBUF_X1 U1073 ( .A(n434), .Z(n1241) );
  XNOR2_X1 U1074 ( .A(a[14]), .B(n37), .ZN(n46) );
  OAI22_X1 U1075 ( .A1(n1318), .A2(n898), .B1(n897), .B2(n1321), .ZN(n1242) );
  CLKBUF_X2 U1076 ( .A(n43), .Z(n1492) );
  CLKBUF_X1 U1077 ( .A(n469), .Z(n1243) );
  XOR2_X1 U1078 ( .A(n525), .B(n523), .Z(n1244) );
  XOR2_X1 U1079 ( .A(n534), .B(n1244), .Z(n517) );
  NAND2_X1 U1080 ( .A1(n534), .A2(n525), .ZN(n1245) );
  NAND2_X1 U1081 ( .A1(n534), .A2(n523), .ZN(n1246) );
  NAND2_X1 U1082 ( .A1(n525), .A2(n523), .ZN(n1247) );
  NAND3_X1 U1083 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n516) );
  CLKBUF_X1 U1084 ( .A(n164), .Z(n1248) );
  XNOR2_X1 U1085 ( .A(n1249), .B(n486), .ZN(n465) );
  XNOR2_X1 U1086 ( .A(n1243), .B(n471), .ZN(n1249) );
  XOR2_X1 U1087 ( .A(n610), .B(n605), .Z(n1250) );
  XOR2_X1 U1088 ( .A(n603), .B(n1250), .Z(n601) );
  NAND2_X1 U1089 ( .A1(n603), .A2(n610), .ZN(n1251) );
  NAND2_X1 U1090 ( .A1(n603), .A2(n605), .ZN(n1252) );
  NAND2_X1 U1091 ( .A1(n610), .A2(n605), .ZN(n1253) );
  NAND3_X1 U1092 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n600) );
  XOR2_X1 U1093 ( .A(n450), .B(n441), .Z(n1254) );
  XOR2_X1 U1094 ( .A(n435), .B(n1254), .Z(n431) );
  NAND2_X1 U1095 ( .A1(n435), .A2(n450), .ZN(n1255) );
  NAND2_X1 U1096 ( .A1(n435), .A2(n441), .ZN(n1256) );
  NAND2_X1 U1097 ( .A1(n450), .A2(n441), .ZN(n1257) );
  NAND3_X1 U1098 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n430) );
  CLKBUF_X3 U1099 ( .A(n43), .Z(n1493) );
  XNOR2_X1 U1100 ( .A(n1554), .B(n1303), .ZN(n1258) );
  CLKBUF_X1 U1101 ( .A(n1096), .Z(n1349) );
  CLKBUF_X1 U1102 ( .A(n544), .Z(n1259) );
  CLKBUF_X1 U1103 ( .A(n150), .Z(n1260) );
  NOR2_X1 U1104 ( .A1(n557), .A2(n568), .ZN(n1261) );
  NOR2_X1 U1105 ( .A1(n557), .A2(n568), .ZN(n204) );
  OR2_X2 U1106 ( .A1(n543), .A2(n556), .ZN(n1511) );
  INV_X1 U1107 ( .A(n665), .ZN(n1262) );
  CLKBUF_X3 U1108 ( .A(n9), .Z(n1530) );
  CLKBUF_X1 U1109 ( .A(n953), .Z(n1263) );
  CLKBUF_X3 U1110 ( .A(n61), .Z(n1300) );
  CLKBUF_X1 U1111 ( .A(n61), .Z(n1548) );
  CLKBUF_X1 U1112 ( .A(n46), .Z(n1343) );
  BUF_X2 U1113 ( .A(n40), .Z(n1526) );
  BUF_X2 U1114 ( .A(n1108), .Z(n1337) );
  XOR2_X1 U1115 ( .A(n544), .B(n533), .Z(n1264) );
  XOR2_X1 U1116 ( .A(n531), .B(n1264), .Z(n529) );
  NAND2_X1 U1117 ( .A1(n531), .A2(n1259), .ZN(n1265) );
  NAND2_X1 U1118 ( .A1(n531), .A2(n533), .ZN(n1266) );
  NAND2_X1 U1119 ( .A1(n1259), .A2(n533), .ZN(n1267) );
  NAND3_X1 U1120 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n528) );
  AND2_X1 U1121 ( .A1(n513), .A2(n528), .ZN(n1295) );
  NOR2_X1 U1122 ( .A1(n397), .A2(n410), .ZN(n1268) );
  NOR2_X1 U1123 ( .A1(n397), .A2(n410), .ZN(n147) );
  OR2_X2 U1124 ( .A1(n513), .A2(n528), .ZN(n1512) );
  XOR2_X1 U1125 ( .A(n1242), .B(n860), .Z(n1269) );
  XOR2_X1 U1126 ( .A(n1269), .B(n769), .Z(n475) );
  NAND2_X1 U1127 ( .A1(n769), .A2(n1242), .ZN(n1270) );
  NAND2_X1 U1128 ( .A1(n769), .A2(n860), .ZN(n1271) );
  NAND2_X1 U1129 ( .A1(n1242), .A2(n860), .ZN(n1272) );
  NAND3_X1 U1130 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n474) );
  CLKBUF_X3 U1131 ( .A(n7), .Z(n1470) );
  NOR2_X2 U1132 ( .A1(n581), .A2(n590), .ZN(n215) );
  BUF_X1 U1133 ( .A(n1100), .Z(n1557) );
  CLKBUF_X1 U1134 ( .A(n161), .Z(n1273) );
  NOR2_X1 U1135 ( .A1(n443), .A2(n460), .ZN(n161) );
  NOR2_X1 U1136 ( .A1(n371), .A2(n382), .ZN(n1274) );
  OAI22_X1 U1137 ( .A1(n1438), .A2(n1028), .B1(n1027), .B2(n1528), .ZN(n1275)
         );
  NOR2_X1 U1138 ( .A1(n371), .A2(n382), .ZN(n135) );
  XNOR2_X1 U1139 ( .A(n1556), .B(n1494), .ZN(n1276) );
  CLKBUF_X1 U1140 ( .A(n1106), .Z(n1336) );
  BUF_X2 U1141 ( .A(n1100), .Z(n1359) );
  XOR2_X1 U1142 ( .A(n418), .B(n407), .Z(n1277) );
  XOR2_X1 U1143 ( .A(n409), .B(n1277), .Z(n401) );
  NAND2_X1 U1144 ( .A1(n409), .A2(n418), .ZN(n1278) );
  NAND2_X1 U1145 ( .A1(n409), .A2(n407), .ZN(n1279) );
  NAND2_X1 U1146 ( .A1(n418), .A2(n407), .ZN(n1280) );
  NAND3_X1 U1147 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n400) );
  XOR2_X1 U1148 ( .A(n693), .B(n820), .Z(n1281) );
  XOR2_X1 U1149 ( .A(n1281), .B(n424), .Z(n409) );
  NAND2_X1 U1150 ( .A1(n424), .A2(n693), .ZN(n1282) );
  NAND2_X1 U1151 ( .A1(n424), .A2(n820), .ZN(n1283) );
  NAND2_X1 U1152 ( .A1(n693), .A2(n820), .ZN(n1284) );
  NAND3_X1 U1153 ( .A1(n1282), .A2(n1283), .A3(n1284), .ZN(n408) );
  XNOR2_X1 U1154 ( .A(n429), .B(n1285), .ZN(n427) );
  XNOR2_X1 U1155 ( .A(n444), .B(n431), .ZN(n1285) );
  BUF_X2 U1156 ( .A(n1553), .Z(n1332) );
  CLKBUF_X1 U1157 ( .A(n162), .Z(n1286) );
  XNOR2_X1 U1158 ( .A(n1287), .B(n440), .ZN(n419) );
  XNOR2_X1 U1159 ( .A(n425), .B(n748), .ZN(n1287) );
  CLKBUF_X3 U1160 ( .A(n13), .Z(n1288) );
  CLKBUF_X1 U1161 ( .A(n140), .Z(n1289) );
  OR2_X2 U1162 ( .A1(n1290), .A2(n1291), .ZN(n54) );
  XNOR2_X1 U1163 ( .A(n1546), .B(a[16]), .ZN(n1290) );
  XOR2_X1 U1164 ( .A(n43), .B(a[16]), .Z(n1291) );
  CLKBUF_X1 U1165 ( .A(n141), .Z(n1292) );
  CLKBUF_X1 U1166 ( .A(n172), .Z(n1294) );
  XOR2_X1 U1167 ( .A(n567), .B(n576), .Z(n1296) );
  XOR2_X1 U1168 ( .A(n574), .B(n1296), .Z(n561) );
  NAND2_X1 U1169 ( .A1(n574), .A2(n567), .ZN(n1297) );
  NAND2_X1 U1170 ( .A1(n574), .A2(n576), .ZN(n1298) );
  NAND2_X1 U1171 ( .A1(n567), .A2(n576), .ZN(n1299) );
  NAND3_X1 U1172 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n560) );
  NOR2_X1 U1173 ( .A1(n411), .A2(n426), .ZN(n150) );
  CLKBUF_X1 U1174 ( .A(n126), .Z(n1301) );
  CLKBUF_X1 U1175 ( .A(n1538), .Z(n1302) );
  CLKBUF_X1 U1176 ( .A(n1367), .Z(n1304) );
  BUF_X1 U1177 ( .A(n1553), .Z(n1330) );
  CLKBUF_X1 U1178 ( .A(n176), .Z(n1306) );
  BUF_X4 U1179 ( .A(n25), .Z(n1307) );
  AOI21_X1 U1180 ( .B1(n1398), .B2(n175), .A(n1306), .ZN(n1308) );
  BUF_X1 U1181 ( .A(n12), .Z(n1366) );
  CLKBUF_X1 U1182 ( .A(n12), .Z(n1368) );
  CLKBUF_X1 U1183 ( .A(n1542), .Z(n1309) );
  CLKBUF_X1 U1184 ( .A(n1099), .Z(n1310) );
  CLKBUF_X1 U1185 ( .A(n1099), .Z(n1340) );
  BUF_X1 U1186 ( .A(n1548), .Z(n1312) );
  NAND2_X1 U1187 ( .A1(n1327), .A2(n300), .ZN(n1313) );
  NAND3_X1 U1188 ( .A1(n1474), .A2(n1313), .A3(n1475), .ZN(n1314) );
  CLKBUF_X1 U1189 ( .A(n1467), .Z(n1315) );
  CLKBUF_X1 U1190 ( .A(n1539), .Z(n1316) );
  NAND2_X1 U1191 ( .A1(n1347), .A2(n1348), .ZN(n1317) );
  NAND2_X1 U1192 ( .A1(n1347), .A2(n1348), .ZN(n1318) );
  NAND2_X1 U1193 ( .A1(n1347), .A2(n1348), .ZN(n60) );
  BUF_X2 U1194 ( .A(n55), .Z(n1319) );
  XNOR2_X1 U1195 ( .A(n1373), .B(a[6]), .ZN(n1507) );
  BUF_X2 U1196 ( .A(n1482), .Z(n1320) );
  BUF_X1 U1197 ( .A(n1482), .Z(n1321) );
  CLKBUF_X1 U1198 ( .A(n1368), .Z(n1322) );
  BUF_X2 U1199 ( .A(n1368), .Z(n1323) );
  BUF_X1 U1200 ( .A(n1471), .Z(n1324) );
  XNOR2_X1 U1201 ( .A(n1325), .B(n791), .ZN(n537) );
  XNOR2_X1 U1202 ( .A(n809), .B(n827), .ZN(n1325) );
  CLKBUF_X1 U1203 ( .A(n1541), .Z(n1326) );
  NAND3_X1 U1204 ( .A1(n1542), .A2(n1541), .A3(n1540), .ZN(n1327) );
  NAND3_X1 U1205 ( .A1(n1309), .A2(n1326), .A3(n1540), .ZN(n1328) );
  OAI22_X1 U1206 ( .A1(n1465), .A2(n1017), .B1(n1016), .B2(n1445), .ZN(n1329)
         );
  CLKBUF_X1 U1207 ( .A(n1553), .Z(n1331) );
  CLKBUF_X1 U1208 ( .A(n1550), .Z(n1333) );
  XNOR2_X1 U1209 ( .A(n1450), .B(a[12]), .ZN(n1113) );
  XNOR2_X1 U1210 ( .A(n1336), .B(n1319), .ZN(n1339) );
  BUF_X2 U1211 ( .A(n1105), .Z(n1341) );
  XNOR2_X1 U1212 ( .A(n19), .B(a[8]), .ZN(n28) );
  CLKBUF_X1 U1213 ( .A(n1504), .Z(n1342) );
  CLKBUF_X1 U1214 ( .A(n1465), .Z(n1344) );
  CLKBUF_X1 U1215 ( .A(n1565), .Z(n1346) );
  BUF_X2 U1216 ( .A(n1092), .Z(n1565) );
  XOR2_X1 U1217 ( .A(n55), .B(a[18]), .Z(n1347) );
  XNOR2_X1 U1218 ( .A(n1546), .B(a[18]), .ZN(n1348) );
  CLKBUF_X1 U1219 ( .A(n1370), .Z(n1350) );
  OAI22_X1 U1220 ( .A1(n24), .A2(n1016), .B1(n1015), .B2(n1527), .ZN(n1351) );
  INV_X1 U1221 ( .A(n1564), .ZN(n1352) );
  INV_X1 U1222 ( .A(n1352), .ZN(n1353) );
  CLKBUF_X3 U1223 ( .A(n19), .Z(n1354) );
  CLKBUF_X1 U1224 ( .A(n1566), .Z(n1355) );
  XNOR2_X1 U1225 ( .A(n7), .B(a[4]), .ZN(n1356) );
  BUF_X2 U1226 ( .A(n52), .Z(n1357) );
  CLKBUF_X2 U1227 ( .A(n52), .Z(n1358) );
  OR2_X1 U1228 ( .A1(n1360), .A2(n668), .ZN(n6) );
  XNOR2_X1 U1229 ( .A(n1), .B(n668), .ZN(n1360) );
  OR2_X2 U1230 ( .A1(n1360), .A2(n668), .ZN(n1361) );
  XNOR2_X1 U1231 ( .A(n1362), .B(n463), .ZN(n461) );
  XNOR2_X1 U1232 ( .A(n480), .B(n465), .ZN(n1362) );
  OAI22_X1 U1233 ( .A1(n1437), .A2(n1035), .B1(n1034), .B2(n1334), .ZN(n1363)
         );
  CLKBUF_X1 U1234 ( .A(n1567), .Z(n1364) );
  BUF_X2 U1235 ( .A(n1090), .Z(n1567) );
  BUF_X2 U1236 ( .A(n19), .Z(n1365) );
  CLKBUF_X3 U1237 ( .A(n12), .Z(n1367) );
  NAND2_X1 U1238 ( .A1(n9), .A2(n1510), .ZN(n12) );
  NAND2_X1 U1239 ( .A1(n1505), .A2(n46), .ZN(n48) );
  INV_X2 U1240 ( .A(n668), .ZN(n1371) );
  CLKBUF_X3 U1241 ( .A(n34), .Z(n1372) );
  INV_X1 U1242 ( .A(n19), .ZN(n1373) );
  CLKBUF_X1 U1243 ( .A(n221), .Z(n1374) );
  AOI21_X1 U1244 ( .B1(n1374), .B2(n213), .A(n214), .ZN(n1375) );
  XOR2_X1 U1245 ( .A(n510), .B(n495), .Z(n1376) );
  XOR2_X1 U1246 ( .A(n1376), .B(n508), .Z(n487) );
  NAND2_X1 U1247 ( .A1(n510), .A2(n495), .ZN(n1377) );
  NAND2_X1 U1248 ( .A1(n510), .A2(n508), .ZN(n1378) );
  NAND2_X1 U1249 ( .A1(n495), .A2(n508), .ZN(n1379) );
  NAND2_X1 U1250 ( .A1(n469), .A2(n471), .ZN(n1380) );
  NAND2_X1 U1251 ( .A1(n471), .A2(n486), .ZN(n1381) );
  NAND2_X1 U1252 ( .A1(n469), .A2(n486), .ZN(n1382) );
  NAND3_X1 U1253 ( .A1(n1380), .A2(n1381), .A3(n1382), .ZN(n464) );
  INV_X1 U1254 ( .A(n1419), .ZN(n187) );
  CLKBUF_X1 U1255 ( .A(n28), .Z(n1529) );
  INV_X1 U1256 ( .A(n1450), .ZN(n1494) );
  CLKBUF_X1 U1257 ( .A(n203), .Z(n1383) );
  XOR2_X1 U1258 ( .A(n541), .B(n539), .Z(n1384) );
  NAND2_X1 U1259 ( .A1(n1351), .A2(n1363), .ZN(n1385) );
  NAND2_X1 U1260 ( .A1(n1351), .A2(n791), .ZN(n1386) );
  NAND2_X1 U1261 ( .A1(n791), .A2(n1363), .ZN(n1387) );
  NAND3_X1 U1262 ( .A1(n1387), .A2(n1386), .A3(n1385), .ZN(n536) );
  NAND2_X1 U1263 ( .A1(n541), .A2(n539), .ZN(n1388) );
  NAND2_X1 U1264 ( .A1(n541), .A2(n537), .ZN(n1389) );
  NAND2_X1 U1265 ( .A1(n539), .A2(n537), .ZN(n1390) );
  NAND3_X1 U1266 ( .A1(n1388), .A2(n1389), .A3(n1390), .ZN(n532) );
  BUF_X2 U1267 ( .A(n36), .Z(n1452) );
  XOR2_X1 U1268 ( .A(n547), .B(n558), .Z(n1391) );
  XOR2_X1 U1269 ( .A(n545), .B(n1391), .Z(n543) );
  NAND2_X1 U1270 ( .A1(n545), .A2(n547), .ZN(n1392) );
  NAND2_X1 U1271 ( .A1(n545), .A2(n558), .ZN(n1393) );
  NAND2_X1 U1272 ( .A1(n547), .A2(n558), .ZN(n1394) );
  NAND3_X1 U1273 ( .A1(n1392), .A2(n1393), .A3(n1394), .ZN(n542) );
  OR2_X1 U1274 ( .A1(n529), .A2(n542), .ZN(n1419) );
  NAND2_X1 U1275 ( .A1(n429), .A2(n444), .ZN(n1395) );
  NAND2_X1 U1276 ( .A1(n429), .A2(n431), .ZN(n1396) );
  NAND2_X1 U1277 ( .A1(n444), .A2(n431), .ZN(n1397) );
  NAND3_X1 U1278 ( .A1(n1395), .A2(n1396), .A3(n1397), .ZN(n426) );
  CLKBUF_X1 U1279 ( .A(n194), .Z(n1398) );
  XOR2_X1 U1280 ( .A(n511), .B(n522), .Z(n1399) );
  XOR2_X1 U1281 ( .A(n1399), .B(n507), .Z(n503) );
  NAND2_X1 U1282 ( .A1(n511), .A2(n522), .ZN(n1400) );
  NAND2_X1 U1283 ( .A1(n511), .A2(n507), .ZN(n1401) );
  NAND2_X1 U1284 ( .A1(n522), .A2(n507), .ZN(n1402) );
  NAND3_X1 U1285 ( .A1(n1400), .A2(n1401), .A3(n1402), .ZN(n502) );
  XOR2_X1 U1286 ( .A(n504), .B(n493), .Z(n1403) );
  XOR2_X1 U1287 ( .A(n1403), .B(n502), .Z(n483) );
  NAND2_X1 U1288 ( .A1(n504), .A2(n493), .ZN(n1404) );
  NAND2_X1 U1289 ( .A1(n504), .A2(n502), .ZN(n1405) );
  NAND2_X1 U1290 ( .A1(n493), .A2(n502), .ZN(n1406) );
  NAND3_X1 U1291 ( .A1(n1404), .A2(n1405), .A3(n1406), .ZN(n482) );
  NAND2_X1 U1292 ( .A1(n482), .A2(n484), .ZN(n1407) );
  NAND2_X1 U1293 ( .A1(n482), .A2(n467), .ZN(n1408) );
  NAND2_X1 U1294 ( .A1(n484), .A2(n467), .ZN(n1409) );
  NAND3_X1 U1295 ( .A1(n1407), .A2(n1408), .A3(n1409), .ZN(n462) );
  BUF_X1 U1296 ( .A(n30), .Z(n1462) );
  XOR2_X1 U1297 ( .A(n811), .B(n829), .Z(n1410) );
  XOR2_X1 U1298 ( .A(n1410), .B(n578), .Z(n563) );
  NAND2_X1 U1299 ( .A1(n811), .A2(n829), .ZN(n1411) );
  NAND2_X1 U1300 ( .A1(n811), .A2(n578), .ZN(n1412) );
  NAND2_X1 U1301 ( .A1(n829), .A2(n578), .ZN(n1413) );
  XOR2_X1 U1302 ( .A(n564), .B(n551), .Z(n1414) );
  XOR2_X1 U1303 ( .A(n1414), .B(n562), .Z(n547) );
  NAND2_X1 U1304 ( .A1(n564), .A2(n551), .ZN(n1415) );
  NAND2_X1 U1305 ( .A1(n564), .A2(n562), .ZN(n1416) );
  NAND2_X1 U1306 ( .A1(n551), .A2(n562), .ZN(n1417) );
  NAND3_X1 U1307 ( .A1(n1415), .A2(n1416), .A3(n1417), .ZN(n546) );
  BUF_X1 U1308 ( .A(n18), .Z(n1437) );
  XOR2_X1 U1309 ( .A(n1329), .B(n672), .Z(n1420) );
  XOR2_X1 U1310 ( .A(n774), .B(n1420), .Z(n553) );
  NAND2_X1 U1311 ( .A1(n774), .A2(n1329), .ZN(n1421) );
  NAND2_X1 U1312 ( .A1(n774), .A2(n672), .ZN(n1422) );
  NAND2_X1 U1313 ( .A1(n810), .A2(n672), .ZN(n1423) );
  NAND3_X1 U1314 ( .A1(n1421), .A2(n1422), .A3(n1423), .ZN(n552) );
  XOR2_X1 U1315 ( .A(n514), .B(n501), .Z(n1424) );
  XOR2_X1 U1316 ( .A(n499), .B(n1424), .Z(n497) );
  NAND2_X1 U1317 ( .A1(n499), .A2(n514), .ZN(n1425) );
  NAND2_X1 U1318 ( .A1(n499), .A2(n501), .ZN(n1426) );
  NAND2_X1 U1319 ( .A1(n514), .A2(n501), .ZN(n1427) );
  NAND3_X1 U1320 ( .A1(n1425), .A2(n1426), .A3(n1427), .ZN(n496) );
  CLKBUF_X1 U1321 ( .A(n264), .Z(n1429) );
  NAND2_X1 U1322 ( .A1(n1507), .A2(n22), .ZN(n24) );
  NAND2_X2 U1323 ( .A1(n1507), .A2(n22), .ZN(n1465) );
  XOR2_X1 U1324 ( .A(n1241), .B(n423), .Z(n1430) );
  XOR2_X1 U1325 ( .A(n1430), .B(n419), .Z(n415) );
  NAND2_X1 U1326 ( .A1(n425), .A2(n748), .ZN(n1431) );
  NAND2_X1 U1327 ( .A1(n425), .A2(n440), .ZN(n1432) );
  NAND2_X1 U1328 ( .A1(n748), .A2(n440), .ZN(n1433) );
  NAND3_X1 U1329 ( .A1(n1431), .A2(n1432), .A3(n1433), .ZN(n418) );
  NAND2_X1 U1330 ( .A1(n434), .A2(n423), .ZN(n1434) );
  NAND2_X1 U1331 ( .A1(n434), .A2(n419), .ZN(n1435) );
  NAND2_X1 U1332 ( .A1(n423), .A2(n419), .ZN(n1436) );
  NAND3_X1 U1333 ( .A1(n1434), .A2(n1435), .A3(n1436), .ZN(n414) );
  BUF_X2 U1334 ( .A(n18), .Z(n1438) );
  NAND2_X1 U1335 ( .A1(n1509), .A2(n1356), .ZN(n18) );
  BUF_X4 U1336 ( .A(n49), .Z(n1439) );
  NAND2_X1 U1337 ( .A1(n13), .A2(a[6]), .ZN(n1443) );
  NAND2_X1 U1338 ( .A1(n1441), .A2(n1442), .ZN(n1444) );
  NAND2_X1 U1339 ( .A1(n1443), .A2(n1444), .ZN(n1464) );
  INV_X1 U1340 ( .A(n13), .ZN(n1441) );
  INV_X1 U1341 ( .A(a[6]), .ZN(n1442) );
  BUF_X2 U1342 ( .A(n1464), .Z(n1527) );
  CLKBUF_X1 U1343 ( .A(n151), .Z(n1446) );
  CLKBUF_X1 U1344 ( .A(n54), .Z(n1447) );
  NAND2_X1 U1345 ( .A1(n1356), .A2(n1509), .ZN(n1471) );
  NOR2_X1 U1346 ( .A1(n497), .A2(n512), .ZN(n1448) );
  CLKBUF_X1 U1347 ( .A(n1372), .Z(n1449) );
  NOR2_X1 U1348 ( .A1(n497), .A2(n512), .ZN(n177) );
  INV_X1 U1349 ( .A(n37), .ZN(n1450) );
  AOI21_X1 U1350 ( .B1(n1512), .B2(n1440), .A(n1295), .ZN(n1451) );
  BUF_X2 U1351 ( .A(n36), .Z(n1453) );
  NAND2_X1 U1352 ( .A1(n1506), .A2(n34), .ZN(n36) );
  CLKBUF_X1 U1353 ( .A(n146), .Z(n1454) );
  CLKBUF_X1 U1354 ( .A(n1321), .Z(n1455) );
  AOI21_X1 U1355 ( .B1(n1454), .B2(n1236), .A(n134), .ZN(n1456) );
  OR2_X1 U1356 ( .A1(n60), .A2(n897), .ZN(n1457) );
  OR2_X1 U1357 ( .A1(n1339), .A2(n1482), .ZN(n1458) );
  NAND2_X1 U1358 ( .A1(n1457), .A2(n1458), .ZN(n696) );
  AND2_X1 U1359 ( .A1(n543), .A2(n556), .ZN(n1459) );
  NOR2_X1 U1360 ( .A1(n427), .A2(n442), .ZN(n1460) );
  NOR2_X1 U1361 ( .A1(n427), .A2(n442), .ZN(n158) );
  CLKBUF_X1 U1362 ( .A(n30), .Z(n1461) );
  NAND2_X1 U1363 ( .A1(n28), .A2(n1508), .ZN(n30) );
  NAND3_X1 U1364 ( .A1(n1474), .A2(n1473), .A3(n1475), .ZN(n1466) );
  NAND3_X1 U1365 ( .A1(n1477), .A2(n1478), .A3(n1479), .ZN(n1467) );
  CLKBUF_X1 U1366 ( .A(n106), .Z(n1468) );
  CLKBUF_X1 U1367 ( .A(n114), .Z(n1469) );
  XOR2_X1 U1368 ( .A(n300), .B(n299), .Z(n1472) );
  XOR2_X1 U1369 ( .A(n1328), .B(n1472), .Z(product[37]) );
  NAND2_X1 U1370 ( .A1(n1327), .A2(n300), .ZN(n1473) );
  NAND2_X1 U1371 ( .A1(n98), .A2(n299), .ZN(n1474) );
  NAND2_X1 U1372 ( .A1(n300), .A2(n299), .ZN(n1475) );
  NAND3_X1 U1373 ( .A1(n1313), .A2(n1474), .A3(n1475), .ZN(n97) );
  XOR2_X1 U1374 ( .A(n310), .B(n307), .Z(n1476) );
  XOR2_X1 U1375 ( .A(n1429), .B(n1476), .Z(product[34]) );
  NAND2_X1 U1376 ( .A1(n264), .A2(n310), .ZN(n1477) );
  NAND2_X1 U1377 ( .A1(n264), .A2(n307), .ZN(n1478) );
  NAND2_X1 U1378 ( .A1(n310), .A2(n307), .ZN(n1479) );
  NAND3_X1 U1379 ( .A1(n1478), .A2(n1477), .A3(n1479), .ZN(n100) );
  AOI21_X1 U1380 ( .B1(n1469), .B2(n1516), .A(n111), .ZN(n1480) );
  CLKBUF_X1 U1381 ( .A(n122), .Z(n1481) );
  XNOR2_X1 U1382 ( .A(n1546), .B(a[18]), .ZN(n1482) );
  CLKBUF_X1 U1383 ( .A(n1317), .Z(n1483) );
  NAND2_X1 U1384 ( .A1(n463), .A2(n480), .ZN(n1484) );
  NAND2_X1 U1385 ( .A1(n463), .A2(n1233), .ZN(n1485) );
  NAND2_X1 U1386 ( .A1(n480), .A2(n1233), .ZN(n1486) );
  NAND3_X1 U1387 ( .A1(n1484), .A2(n1485), .A3(n1486), .ZN(n460) );
  NOR2_X1 U1388 ( .A1(n461), .A2(n478), .ZN(n1487) );
  NAND2_X1 U1389 ( .A1(n43), .A2(n1489), .ZN(n1490) );
  NAND2_X1 U1390 ( .A1(n1488), .A2(a[14]), .ZN(n1491) );
  NAND2_X1 U1391 ( .A1(n1490), .A2(n1491), .ZN(n1505) );
  INV_X1 U1392 ( .A(n43), .ZN(n1488) );
  INV_X1 U1393 ( .A(a[14]), .ZN(n1489) );
  NOR2_X1 U1394 ( .A1(n461), .A2(n478), .ZN(n166) );
  CLKBUF_X1 U1395 ( .A(n127), .Z(n1495) );
  NAND2_X1 U1396 ( .A1(n7), .A2(n1497), .ZN(n1498) );
  NAND2_X1 U1397 ( .A1(n1496), .A2(a[2]), .ZN(n1499) );
  NAND2_X1 U1398 ( .A1(n1499), .A2(n1498), .ZN(n1510) );
  INV_X1 U1399 ( .A(n7), .ZN(n1496) );
  INV_X1 U1400 ( .A(a[2]), .ZN(n1497) );
  AOI21_X1 U1401 ( .B1(n122), .B2(n1517), .A(n119), .ZN(n1500) );
  CLKBUF_X1 U1402 ( .A(n153), .Z(n1501) );
  AOI21_X1 U1403 ( .B1(n153), .B2(n126), .A(n127), .ZN(n1502) );
  NAND2_X1 U1404 ( .A1(n1113), .A2(n40), .ZN(n1503) );
  NAND2_X2 U1405 ( .A1(n1113), .A2(n40), .ZN(n1504) );
  NOR2_X1 U1406 ( .A1(n359), .A2(n370), .ZN(n128) );
  NAND2_X1 U1407 ( .A1(n443), .A2(n460), .ZN(n162) );
  OR2_X1 U1408 ( .A1(n339), .A2(n348), .ZN(n1517) );
  XOR2_X1 U1409 ( .A(n31), .B(a[10]), .Z(n1506) );
  XOR2_X1 U1410 ( .A(n25), .B(a[8]), .Z(n1508) );
  XOR2_X1 U1411 ( .A(n13), .B(a[4]), .Z(n1509) );
  OAI21_X1 U1412 ( .B1(n152), .B2(n143), .A(n144), .ZN(n142) );
  INV_X1 U1413 ( .A(n145), .ZN(n143) );
  INV_X1 U1414 ( .A(n1501), .ZN(n152) );
  NAND2_X1 U1415 ( .A1(n145), .A2(n133), .ZN(n131) );
  XNOR2_X1 U1416 ( .A(n179), .B(n78), .ZN(product[18]) );
  NAND2_X1 U1417 ( .A1(n280), .A2(n178), .ZN(n78) );
  INV_X1 U1418 ( .A(n1448), .ZN(n280) );
  INV_X1 U1419 ( .A(n171), .ZN(n279) );
  INV_X1 U1420 ( .A(n1289), .ZN(n273) );
  XOR2_X1 U1421 ( .A(n168), .B(n76), .Z(product[20]) );
  NAND2_X1 U1422 ( .A1(n278), .A2(n167), .ZN(n76) );
  AOI21_X1 U1423 ( .B1(n173), .B2(n279), .A(n170), .ZN(n168) );
  XOR2_X1 U1424 ( .A(n137), .B(n70), .Z(product[26]) );
  NAND2_X1 U1425 ( .A1(n272), .A2(n136), .ZN(n70) );
  AOI21_X1 U1426 ( .B1(n142), .B2(n273), .A(n139), .ZN(n137) );
  XOR2_X1 U1427 ( .A(n206), .B(n82), .Z(product[14]) );
  NAND2_X1 U1428 ( .A1(n284), .A2(n205), .ZN(n82) );
  AOI21_X1 U1429 ( .B1(n211), .B2(n285), .A(n208), .ZN(n206) );
  XOR2_X1 U1430 ( .A(n201), .B(n81), .Z(product[15]) );
  AOI21_X1 U1431 ( .B1(n211), .B2(n202), .A(n1383), .ZN(n201) );
  XOR2_X1 U1432 ( .A(n163), .B(n75), .Z(product[21]) );
  NAND2_X1 U1433 ( .A1(n277), .A2(n1286), .ZN(n75) );
  INV_X1 U1434 ( .A(n1273), .ZN(n277) );
  XOR2_X1 U1435 ( .A(n152), .B(n73), .Z(product[23]) );
  NAND2_X1 U1436 ( .A1(n275), .A2(n1446), .ZN(n73) );
  XOR2_X1 U1437 ( .A(n193), .B(n80), .Z(product[16]) );
  NAND2_X1 U1438 ( .A1(n1419), .A2(n188), .ZN(n80) );
  XNOR2_X1 U1439 ( .A(n173), .B(n77), .ZN(product[19]) );
  NAND2_X1 U1440 ( .A1(n279), .A2(n1294), .ZN(n77) );
  XNOR2_X1 U1441 ( .A(n160), .B(n74), .ZN(product[22]) );
  NAND2_X1 U1442 ( .A1(n276), .A2(n159), .ZN(n74) );
  OAI21_X1 U1443 ( .B1(n163), .B2(n1273), .A(n1286), .ZN(n160) );
  XNOR2_X1 U1444 ( .A(n130), .B(n69), .ZN(product[27]) );
  NAND2_X1 U1445 ( .A1(n271), .A2(n129), .ZN(n69) );
  INV_X1 U1446 ( .A(n128), .ZN(n271) );
  XNOR2_X1 U1447 ( .A(n149), .B(n72), .ZN(product[24]) );
  NAND2_X1 U1448 ( .A1(n274), .A2(n148), .ZN(n72) );
  INV_X1 U1449 ( .A(n1268), .ZN(n274) );
  XNOR2_X1 U1450 ( .A(n186), .B(n79), .ZN(product[17]) );
  OAI21_X1 U1451 ( .B1(n193), .B2(n187), .A(n188), .ZN(n186) );
  XNOR2_X1 U1452 ( .A(n142), .B(n71), .ZN(product[25]) );
  NAND2_X1 U1453 ( .A1(n273), .A2(n1292), .ZN(n71) );
  INV_X1 U1454 ( .A(n1294), .ZN(n170) );
  INV_X1 U1455 ( .A(n1292), .ZN(n139) );
  INV_X1 U1456 ( .A(n121), .ZN(n119) );
  INV_X1 U1457 ( .A(n113), .ZN(n111) );
  NOR2_X1 U1458 ( .A1(n215), .A2(n218), .ZN(n213) );
  OAI21_X1 U1459 ( .B1(n215), .B2(n219), .A(n216), .ZN(n214) );
  OAI21_X1 U1460 ( .B1(n204), .B2(n210), .A(n205), .ZN(n203) );
  NAND2_X1 U1461 ( .A1(n1514), .A2(n1513), .ZN(n222) );
  NAND2_X1 U1462 ( .A1(n268), .A2(n116), .ZN(n66) );
  INV_X1 U1463 ( .A(n115), .ZN(n268) );
  NAND2_X1 U1464 ( .A1(n266), .A2(n108), .ZN(n64) );
  INV_X1 U1465 ( .A(n107), .ZN(n266) );
  NAND2_X1 U1466 ( .A1(n270), .A2(n124), .ZN(n68) );
  INV_X1 U1467 ( .A(n123), .ZN(n270) );
  NAND2_X1 U1468 ( .A1(n411), .A2(n426), .ZN(n151) );
  AOI21_X1 U1469 ( .B1(n239), .B2(n1515), .A(n236), .ZN(n234) );
  INV_X1 U1470 ( .A(n238), .ZN(n236) );
  INV_X1 U1471 ( .A(n209), .ZN(n285) );
  NAND2_X1 U1472 ( .A1(n1517), .A2(n121), .ZN(n67) );
  NAND2_X1 U1473 ( .A1(n1516), .A2(n113), .ZN(n65) );
  NAND2_X1 U1474 ( .A1(n1518), .A2(n105), .ZN(n63) );
  XOR2_X1 U1475 ( .A(n228), .B(n86), .Z(product[10]) );
  NAND2_X1 U1476 ( .A1(n1514), .A2(n227), .ZN(n86) );
  AOI21_X1 U1477 ( .B1(n233), .B2(n1513), .A(n230), .ZN(n228) );
  XOR2_X1 U1478 ( .A(n220), .B(n85), .Z(product[11]) );
  NAND2_X1 U1479 ( .A1(n287), .A2(n219), .ZN(n85) );
  INV_X1 U1480 ( .A(n218), .ZN(n287) );
  NOR2_X1 U1481 ( .A1(n383), .A2(n396), .ZN(n140) );
  NOR2_X1 U1482 ( .A1(n479), .A2(n496), .ZN(n171) );
  XNOR2_X1 U1483 ( .A(n239), .B(n88), .ZN(product[8]) );
  NAND2_X1 U1484 ( .A1(n1515), .A2(n238), .ZN(n88) );
  XNOR2_X1 U1485 ( .A(n211), .B(n83), .ZN(product[13]) );
  NAND2_X1 U1486 ( .A1(n285), .A2(n210), .ZN(n83) );
  NAND2_X1 U1487 ( .A1(n383), .A2(n396), .ZN(n141) );
  NAND2_X1 U1488 ( .A1(n479), .A2(n496), .ZN(n172) );
  XNOR2_X1 U1489 ( .A(n233), .B(n87), .ZN(product[9]) );
  NAND2_X1 U1490 ( .A1(n1513), .A2(n232), .ZN(n87) );
  XNOR2_X1 U1491 ( .A(n217), .B(n84), .ZN(product[12]) );
  NAND2_X1 U1492 ( .A1(n286), .A2(n216), .ZN(n84) );
  OAI21_X1 U1493 ( .B1(n220), .B2(n218), .A(n219), .ZN(n217) );
  INV_X1 U1494 ( .A(n215), .ZN(n286) );
  NAND2_X1 U1495 ( .A1(n359), .A2(n370), .ZN(n129) );
  NAND2_X1 U1496 ( .A1(n427), .A2(n442), .ZN(n159) );
  NAND2_X1 U1497 ( .A1(n497), .A2(n512), .ZN(n178) );
  NAND2_X1 U1498 ( .A1(n397), .A2(n410), .ZN(n148) );
  INV_X1 U1499 ( .A(n210), .ZN(n208) );
  INV_X1 U1500 ( .A(n246), .ZN(n244) );
  OAI21_X1 U1501 ( .B1(n256), .B2(n258), .A(n257), .ZN(n255) );
  AOI21_X1 U1502 ( .B1(n1521), .B2(n255), .A(n252), .ZN(n250) );
  NOR2_X1 U1503 ( .A1(n591), .A2(n600), .ZN(n218) );
  OR2_X1 U1504 ( .A1(n609), .A2(n616), .ZN(n1513) );
  NAND2_X1 U1505 ( .A1(n291), .A2(n241), .ZN(n89) );
  INV_X1 U1506 ( .A(n240), .ZN(n291) );
  OR2_X1 U1507 ( .A1(n601), .A2(n608), .ZN(n1514) );
  NAND2_X1 U1508 ( .A1(n591), .A2(n600), .ZN(n219) );
  OR2_X1 U1509 ( .A1(n617), .A2(n622), .ZN(n1515) );
  XOR2_X1 U1510 ( .A(n91), .B(n250), .Z(product[5]) );
  NAND2_X1 U1511 ( .A1(n293), .A2(n249), .ZN(n91) );
  INV_X1 U1512 ( .A(n248), .ZN(n293) );
  NOR2_X1 U1513 ( .A1(n569), .A2(n580), .ZN(n209) );
  NOR2_X1 U1514 ( .A1(n331), .A2(n338), .ZN(n115) );
  NOR2_X1 U1515 ( .A1(n317), .A2(n322), .ZN(n107) );
  NOR2_X1 U1516 ( .A1(n349), .A2(n358), .ZN(n123) );
  NAND2_X1 U1517 ( .A1(n569), .A2(n580), .ZN(n210) );
  NAND2_X1 U1518 ( .A1(n581), .A2(n590), .ZN(n216) );
  XNOR2_X1 U1519 ( .A(n90), .B(n247), .ZN(product[6]) );
  NAND2_X1 U1520 ( .A1(n1522), .A2(n246), .ZN(n90) );
  XNOR2_X1 U1521 ( .A(n92), .B(n255), .ZN(product[4]) );
  NAND2_X1 U1522 ( .A1(n1521), .A2(n254), .ZN(n92) );
  NAND2_X1 U1523 ( .A1(n323), .A2(n330), .ZN(n113) );
  NAND2_X1 U1524 ( .A1(n339), .A2(n348), .ZN(n121) );
  NAND2_X1 U1525 ( .A1(n311), .A2(n316), .ZN(n105) );
  NAND2_X1 U1526 ( .A1(n617), .A2(n622), .ZN(n238) );
  NAND2_X1 U1527 ( .A1(n609), .A2(n616), .ZN(n232) );
  NAND2_X1 U1528 ( .A1(n331), .A2(n338), .ZN(n116) );
  NAND2_X1 U1529 ( .A1(n317), .A2(n322), .ZN(n108) );
  NAND2_X1 U1530 ( .A1(n349), .A2(n358), .ZN(n124) );
  INV_X1 U1531 ( .A(n259), .ZN(n258) );
  OAI21_X1 U1532 ( .B1(n260), .B2(n263), .A(n261), .ZN(n259) );
  OR2_X1 U1533 ( .A1(n323), .A2(n330), .ZN(n1516) );
  OR2_X1 U1534 ( .A1(n311), .A2(n316), .ZN(n1518) );
  NAND2_X1 U1535 ( .A1(n601), .A2(n608), .ZN(n227) );
  XOR2_X1 U1536 ( .A(n93), .B(n258), .Z(product[3]) );
  NAND2_X1 U1537 ( .A1(n295), .A2(n257), .ZN(n93) );
  INV_X1 U1538 ( .A(n256), .ZN(n295) );
  XOR2_X1 U1539 ( .A(n94), .B(n263), .Z(product[2]) );
  NAND2_X1 U1540 ( .A1(n296), .A2(n261), .ZN(n94) );
  INV_X1 U1541 ( .A(n260), .ZN(n296) );
  INV_X1 U1542 ( .A(n105), .ZN(n103) );
  NAND2_X1 U1543 ( .A1(n639), .A2(n678), .ZN(n257) );
  NOR2_X1 U1544 ( .A1(n878), .A2(n859), .ZN(n260) );
  XNOR2_X1 U1545 ( .A(n1519), .B(n1535), .ZN(product[36]) );
  XNOR2_X1 U1546 ( .A(n302), .B(n301), .ZN(n1519) );
  XNOR2_X1 U1547 ( .A(n1314), .B(n1520), .ZN(product[38]) );
  XNOR2_X1 U1548 ( .A(n680), .B(n298), .ZN(n1520) );
  NAND2_X1 U1549 ( .A1(n679), .A2(n879), .ZN(n263) );
  NOR2_X1 U1550 ( .A1(n639), .A2(n678), .ZN(n256) );
  NAND2_X1 U1551 ( .A1(n878), .A2(n859), .ZN(n261) );
  INV_X1 U1552 ( .A(n394), .ZN(n395) );
  INV_X1 U1553 ( .A(n328), .ZN(n329) );
  NOR2_X1 U1554 ( .A1(n633), .A2(n636), .ZN(n248) );
  NOR2_X1 U1555 ( .A1(n623), .A2(n628), .ZN(n240) );
  NAND2_X1 U1556 ( .A1(n629), .A2(n632), .ZN(n246) );
  OR2_X1 U1557 ( .A1(n637), .A2(n638), .ZN(n1521) );
  NAND2_X1 U1558 ( .A1(n633), .A2(n636), .ZN(n249) );
  NAND2_X1 U1559 ( .A1(n623), .A2(n628), .ZN(n241) );
  NAND2_X1 U1560 ( .A1(n637), .A2(n638), .ZN(n254) );
  OR2_X1 U1561 ( .A1(n629), .A2(n632), .ZN(n1522) );
  AND3_X1 U1562 ( .A1(n1532), .A2(n1531), .A3(n1533), .ZN(product[39]) );
  OR2_X1 U1563 ( .A1(n1312), .A2(n1148), .ZN(n1068) );
  OAI22_X1 U1564 ( .A1(n1361), .A2(n1086), .B1(n1085), .B2(n1371), .ZN(n877)
         );
  OAI22_X1 U1565 ( .A1(n1361), .A2(n1088), .B1(n1087), .B2(n1371), .ZN(n879)
         );
  OAI22_X1 U1566 ( .A1(n1361), .A2(n1149), .B1(n1089), .B2(n1371), .ZN(n679)
         );
  OR2_X1 U1567 ( .A1(n1300), .A2(n1149), .ZN(n1089) );
  OAI22_X1 U1568 ( .A1(n1361), .A2(n1087), .B1(n1086), .B2(n1371), .ZN(n878)
         );
  OAI22_X1 U1569 ( .A1(n1361), .A2(n1072), .B1(n1071), .B2(n1371), .ZN(n863)
         );
  OAI22_X1 U1570 ( .A1(n1361), .A2(n1078), .B1(n1077), .B2(n1371), .ZN(n869)
         );
  XNOR2_X1 U1571 ( .A(n1548), .B(n1439), .ZN(n920) );
  OAI22_X1 U1572 ( .A1(n1361), .A2(n1084), .B1(n1083), .B2(n1371), .ZN(n875)
         );
  OAI22_X1 U1573 ( .A1(n1069), .A2(n6), .B1(n1069), .B2(n1371), .ZN(n667) );
  OR2_X1 U1574 ( .A1(n1312), .A2(n1147), .ZN(n1047) );
  AND2_X1 U1575 ( .A1(n1312), .A2(n662), .ZN(n839) );
  OAI22_X1 U1576 ( .A1(n1361), .A2(n1085), .B1(n1084), .B2(n1371), .ZN(n876)
         );
  XNOR2_X1 U1577 ( .A(n1364), .B(n1439), .ZN(n901) );
  INV_X1 U1578 ( .A(n643), .ZN(n700) );
  INV_X1 U1579 ( .A(n304), .ZN(n305) );
  BUF_X2 U1580 ( .A(n40), .Z(n1525) );
  BUF_X1 U1581 ( .A(n1096), .Z(n1561) );
  BUF_X1 U1582 ( .A(n1099), .Z(n1558) );
  BUF_X1 U1583 ( .A(n1104), .Z(n1553) );
  BUF_X1 U1584 ( .A(n1108), .Z(n1549) );
  XNOR2_X1 U1585 ( .A(n1341), .B(n1439), .ZN(n916) );
  XNOR2_X1 U1586 ( .A(n1551), .B(n1439), .ZN(n917) );
  XNOR2_X1 U1587 ( .A(n1562), .B(n1439), .ZN(n906) );
  XNOR2_X1 U1588 ( .A(n1330), .B(n1439), .ZN(n915) );
  XNOR2_X1 U1589 ( .A(n1561), .B(n1439), .ZN(n907) );
  XNOR2_X1 U1590 ( .A(n1550), .B(n1439), .ZN(n918) );
  XNOR2_X1 U1591 ( .A(n1560), .B(n1439), .ZN(n908) );
  XNOR2_X1 U1592 ( .A(n1305), .B(n1439), .ZN(n914) );
  XNOR2_X1 U1593 ( .A(n1549), .B(n1439), .ZN(n919) );
  XNOR2_X1 U1594 ( .A(n1555), .B(n1439), .ZN(n913) );
  XNOR2_X1 U1595 ( .A(n1556), .B(n1439), .ZN(n912) );
  XNOR2_X1 U1596 ( .A(n1359), .B(n1439), .ZN(n911) );
  XNOR2_X1 U1597 ( .A(n1310), .B(n1439), .ZN(n910) );
  XNOR2_X1 U1598 ( .A(n1559), .B(n1439), .ZN(n909) );
  XNOR2_X1 U1599 ( .A(n1563), .B(n1439), .ZN(n905) );
  XNOR2_X1 U1600 ( .A(n1355), .B(n1439), .ZN(n902) );
  XNOR2_X1 U1601 ( .A(n1353), .B(n1439), .ZN(n904) );
  XNOR2_X1 U1602 ( .A(n1346), .B(n1439), .ZN(n903) );
  XNOR2_X1 U1603 ( .A(n1551), .B(n1319), .ZN(n896) );
  XNOR2_X1 U1604 ( .A(n1559), .B(n1547), .ZN(n888) );
  XNOR2_X1 U1605 ( .A(n1552), .B(n1547), .ZN(n895) );
  XNOR2_X1 U1606 ( .A(n1558), .B(n1547), .ZN(n889) );
  XNOR2_X1 U1607 ( .A(n1555), .B(n1547), .ZN(n892) );
  XNOR2_X1 U1608 ( .A(n1107), .B(n1319), .ZN(n897) );
  XNOR2_X1 U1609 ( .A(n1331), .B(n1547), .ZN(n894) );
  XNOR2_X1 U1610 ( .A(n1554), .B(n1547), .ZN(n893) );
  XNOR2_X1 U1611 ( .A(n1549), .B(n1547), .ZN(n898) );
  XNOR2_X1 U1612 ( .A(n1556), .B(n1547), .ZN(n891) );
  XNOR2_X1 U1613 ( .A(n1359), .B(n1547), .ZN(n890) );
  XNOR2_X1 U1614 ( .A(n1560), .B(n1547), .ZN(n887) );
  XNOR2_X1 U1615 ( .A(n1349), .B(n1547), .ZN(n886) );
  XNOR2_X1 U1616 ( .A(n1562), .B(n1547), .ZN(n885) );
  XNOR2_X1 U1617 ( .A(n1563), .B(n1547), .ZN(n884) );
  XNOR2_X1 U1618 ( .A(n1353), .B(n1547), .ZN(n883) );
  XNOR2_X1 U1619 ( .A(n1346), .B(n1547), .ZN(n882) );
  XNOR2_X1 U1620 ( .A(n1355), .B(n1547), .ZN(n881) );
  AND2_X1 U1621 ( .A1(n1312), .A2(n665), .ZN(n859) );
  INV_X1 U1622 ( .A(n655), .ZN(n780) );
  INV_X1 U1623 ( .A(n314), .ZN(n315) );
  AND2_X1 U1624 ( .A1(n1312), .A2(n641), .ZN(n699) );
  OAI22_X1 U1625 ( .A1(n1361), .A2(n1071), .B1(n1070), .B2(n1371), .ZN(n862)
         );
  INV_X1 U1626 ( .A(n649), .ZN(n740) );
  INV_X1 U1627 ( .A(n346), .ZN(n347) );
  AND2_X1 U1628 ( .A1(n1300), .A2(n1291), .ZN(n719) );
  OAI22_X1 U1629 ( .A1(n6), .A2(n1073), .B1(n1072), .B2(n1371), .ZN(n864) );
  AND2_X1 U1630 ( .A1(n1312), .A2(n650), .ZN(n759) );
  OAI22_X1 U1631 ( .A1(n6), .A2(n1077), .B1(n1076), .B2(n1371), .ZN(n868) );
  INV_X1 U1632 ( .A(n667), .ZN(n860) );
  INV_X1 U1633 ( .A(n652), .ZN(n760) );
  INV_X1 U1634 ( .A(n646), .ZN(n720) );
  INV_X1 U1635 ( .A(n1275), .ZN(n425) );
  OAI22_X1 U1636 ( .A1(n1361), .A2(n1080), .B1(n1079), .B2(n1371), .ZN(n871)
         );
  AND2_X1 U1637 ( .A1(n1312), .A2(n647), .ZN(n739) );
  OAI22_X1 U1638 ( .A1(n1361), .A2(n1075), .B1(n1074), .B2(n1371), .ZN(n866)
         );
  AND2_X1 U1639 ( .A1(n1300), .A2(n653), .ZN(n779) );
  OAI22_X1 U1640 ( .A1(n1361), .A2(n1079), .B1(n1078), .B2(n1371), .ZN(n870)
         );
  OAI22_X1 U1641 ( .A1(n1361), .A2(n1074), .B1(n1073), .B2(n1371), .ZN(n865)
         );
  OAI22_X1 U1642 ( .A1(n1361), .A2(n1082), .B1(n1081), .B2(n1371), .ZN(n873)
         );
  AND2_X1 U1643 ( .A1(n61), .A2(n659), .ZN(n819) );
  OAI22_X1 U1644 ( .A1(n1361), .A2(n1083), .B1(n1082), .B2(n1371), .ZN(n874)
         );
  OAI22_X1 U1645 ( .A1(n1361), .A2(n1076), .B1(n1075), .B2(n1371), .ZN(n867)
         );
  OAI22_X1 U1646 ( .A1(n6), .A2(n1070), .B1(n1069), .B2(n1371), .ZN(n861) );
  OAI22_X1 U1647 ( .A1(n1361), .A2(n1081), .B1(n1080), .B2(n1371), .ZN(n872)
         );
  AND2_X1 U1648 ( .A1(n1312), .A2(n656), .ZN(n799) );
  INV_X1 U1649 ( .A(n458), .ZN(n459) );
  INV_X1 U1650 ( .A(n368), .ZN(n369) );
  XNOR2_X1 U1651 ( .A(n1300), .B(n1547), .ZN(n899) );
  INV_X1 U1652 ( .A(n658), .ZN(n800) );
  INV_X1 U1653 ( .A(n661), .ZN(n820) );
  INV_X1 U1654 ( .A(n1439), .ZN(n1141) );
  INV_X1 U1655 ( .A(n1319), .ZN(n1140) );
  OR2_X1 U1656 ( .A1(n1548), .A2(n1140), .ZN(n900) );
  OR2_X1 U1657 ( .A1(n1312), .A2(n1144), .ZN(n984) );
  OR2_X1 U1658 ( .A1(n1300), .A2(n1143), .ZN(n963) );
  OR2_X1 U1659 ( .A1(n1312), .A2(n1373), .ZN(n1026) );
  OR2_X1 U1660 ( .A1(n1548), .A2(n1142), .ZN(n942) );
  OR2_X1 U1661 ( .A1(n1300), .A2(n1141), .ZN(n921) );
  OR2_X1 U1662 ( .A1(n61), .A2(n1145), .ZN(n1005) );
  XNOR2_X1 U1663 ( .A(n1364), .B(n1547), .ZN(n880) );
  BUF_X4 U1664 ( .A(n55), .Z(n1547) );
  AND2_X1 U1665 ( .A1(n1312), .A2(n668), .ZN(product[0]) );
  XNOR2_X1 U1666 ( .A(n43), .B(a[16]), .ZN(n52) );
  XNOR2_X1 U1667 ( .A(n31), .B(a[12]), .ZN(n40) );
  XNOR2_X1 U1668 ( .A(n25), .B(a[10]), .ZN(n34) );
  XNOR2_X1 U1669 ( .A(n13), .B(a[6]), .ZN(n22) );
  XNOR2_X1 U1670 ( .A(n1), .B(a[2]), .ZN(n9) );
  NAND2_X1 U1671 ( .A1(n1466), .A2(n680), .ZN(n1531) );
  NAND2_X1 U1672 ( .A1(n97), .A2(n298), .ZN(n1532) );
  NAND2_X1 U1673 ( .A1(n680), .A2(n298), .ZN(n1533) );
  INV_X1 U1674 ( .A(n640), .ZN(n680) );
  NAND3_X1 U1675 ( .A1(n1539), .A2(n1538), .A3(n1537), .ZN(n1534) );
  NAND3_X1 U1676 ( .A1(n1316), .A2(n1302), .A3(n1537), .ZN(n1535) );
  AOI21_X1 U1677 ( .B1(n1522), .B2(n247), .A(n244), .ZN(n242) );
  XOR2_X1 U1678 ( .A(n303), .B(n306), .Z(n1536) );
  XOR2_X1 U1679 ( .A(n1536), .B(n1315), .Z(product[35]) );
  NAND2_X1 U1680 ( .A1(n303), .A2(n306), .ZN(n1537) );
  NAND2_X1 U1681 ( .A1(n303), .A2(n100), .ZN(n1538) );
  NAND2_X1 U1682 ( .A1(n1467), .A2(n306), .ZN(n1539) );
  NAND3_X1 U1683 ( .A1(n1539), .A2(n1538), .A3(n1537), .ZN(n99) );
  NAND2_X1 U1684 ( .A1(n302), .A2(n301), .ZN(n1540) );
  NAND2_X1 U1685 ( .A1(n1534), .A2(n302), .ZN(n1541) );
  NAND2_X1 U1686 ( .A1(n301), .A2(n99), .ZN(n1542) );
  NAND3_X1 U1687 ( .A1(n1542), .A2(n1541), .A3(n1540), .ZN(n98) );
  XNOR2_X1 U1688 ( .A(n1549), .B(n1338), .ZN(n961) );
  XNOR2_X1 U1689 ( .A(n1300), .B(n1338), .ZN(n962) );
  XNOR2_X1 U1690 ( .A(n1556), .B(n1494), .ZN(n954) );
  XNOR2_X1 U1691 ( .A(n1550), .B(n1338), .ZN(n960) );
  XNOR2_X1 U1692 ( .A(n1554), .B(n1303), .ZN(n956) );
  XNOR2_X1 U1693 ( .A(n1332), .B(n1303), .ZN(n957) );
  XNOR2_X1 U1694 ( .A(n1560), .B(n1338), .ZN(n950) );
  XNOR2_X1 U1695 ( .A(n1349), .B(n1303), .ZN(n949) );
  XNOR2_X1 U1696 ( .A(n1563), .B(n1303), .ZN(n947) );
  XNOR2_X1 U1697 ( .A(n1353), .B(n1303), .ZN(n946) );
  XNOR2_X1 U1698 ( .A(n1364), .B(n1303), .ZN(n943) );
  XNOR2_X1 U1699 ( .A(n1355), .B(n1338), .ZN(n944) );
  XNOR2_X1 U1700 ( .A(n1346), .B(n1338), .ZN(n945) );
  XNOR2_X1 U1701 ( .A(n1562), .B(n1338), .ZN(n948) );
  XNOR2_X1 U1702 ( .A(n1559), .B(n1338), .ZN(n951) );
  XNOR2_X1 U1703 ( .A(n1558), .B(n1303), .ZN(n952) );
  INV_X1 U1704 ( .A(n1303), .ZN(n1143) );
  XNOR2_X1 U1705 ( .A(n1345), .B(n1303), .ZN(n955) );
  XNOR2_X1 U1706 ( .A(n1557), .B(n1303), .ZN(n953) );
  XNOR2_X1 U1707 ( .A(n1336), .B(n1303), .ZN(n959) );
  XNOR2_X1 U1708 ( .A(n1552), .B(n1303), .ZN(n958) );
  INV_X1 U1709 ( .A(n1543), .ZN(n1149) );
  XNOR2_X1 U1710 ( .A(n1563), .B(n1543), .ZN(n1073) );
  XNOR2_X1 U1711 ( .A(n1341), .B(n1335), .ZN(n1084) );
  XNOR2_X1 U1712 ( .A(n1562), .B(n1335), .ZN(n1074) );
  XNOR2_X1 U1713 ( .A(n1305), .B(n1543), .ZN(n1082) );
  XNOR2_X1 U1714 ( .A(n1560), .B(n1543), .ZN(n1076) );
  XNOR2_X1 U1715 ( .A(n1349), .B(n1543), .ZN(n1075) );
  XNOR2_X1 U1716 ( .A(n1558), .B(n1335), .ZN(n1078) );
  XNOR2_X1 U1717 ( .A(n1565), .B(n1335), .ZN(n1071) );
  XNOR2_X1 U1718 ( .A(n1555), .B(n1335), .ZN(n1081) );
  XNOR2_X1 U1719 ( .A(n1556), .B(n1543), .ZN(n1080) );
  XNOR2_X1 U1720 ( .A(n1359), .B(n1543), .ZN(n1079) );
  XNOR2_X1 U1721 ( .A(n1559), .B(n1335), .ZN(n1077) );
  XNOR2_X1 U1722 ( .A(n1566), .B(n1543), .ZN(n1070) );
  XNOR2_X1 U1723 ( .A(n1333), .B(n1335), .ZN(n1086) );
  XNOR2_X1 U1724 ( .A(n1551), .B(n1543), .ZN(n1085) );
  XNOR2_X1 U1725 ( .A(n1300), .B(n1543), .ZN(n1088) );
  XNOR2_X1 U1726 ( .A(n1331), .B(n1335), .ZN(n1083) );
  XNOR2_X1 U1727 ( .A(n1564), .B(n1335), .ZN(n1072) );
  XNOR2_X1 U1728 ( .A(n1337), .B(n1335), .ZN(n1087) );
  XNOR2_X1 U1729 ( .A(n1567), .B(n1543), .ZN(n1069) );
  AOI21_X1 U1730 ( .B1(n146), .B2(n133), .A(n134), .ZN(n132) );
  INV_X1 U1731 ( .A(n1454), .ZN(n144) );
  AOI21_X1 U1732 ( .B1(n1514), .B2(n230), .A(n225), .ZN(n223) );
  INV_X1 U1733 ( .A(n227), .ZN(n225) );
  INV_X1 U1734 ( .A(n232), .ZN(n230) );
  AOI21_X1 U1735 ( .B1(n173), .B2(n1248), .A(n1235), .ZN(n163) );
  XNOR2_X1 U1736 ( .A(n1567), .B(n1354), .ZN(n1006) );
  XNOR2_X1 U1737 ( .A(n1565), .B(n1354), .ZN(n1008) );
  XNOR2_X1 U1738 ( .A(n1300), .B(n1354), .ZN(n1025) );
  XNOR2_X1 U1739 ( .A(n1566), .B(n1354), .ZN(n1007) );
  XNOR2_X1 U1740 ( .A(n1564), .B(n1354), .ZN(n1009) );
  XNOR2_X1 U1741 ( .A(n1337), .B(n1354), .ZN(n1024) );
  XNOR2_X1 U1742 ( .A(n1559), .B(n1354), .ZN(n1014) );
  XNOR2_X1 U1743 ( .A(n1562), .B(n1365), .ZN(n1011) );
  XNOR2_X1 U1744 ( .A(n1333), .B(n1354), .ZN(n1023) );
  XNOR2_X1 U1745 ( .A(n1563), .B(n1365), .ZN(n1010) );
  XNOR2_X1 U1746 ( .A(n1560), .B(n1365), .ZN(n1013) );
  XNOR2_X1 U1747 ( .A(n1332), .B(n1354), .ZN(n1020) );
  XNOR2_X1 U1748 ( .A(n1561), .B(n1365), .ZN(n1012) );
  XNOR2_X1 U1749 ( .A(n1305), .B(n1354), .ZN(n1019) );
  XNOR2_X1 U1750 ( .A(n1555), .B(n1354), .ZN(n1018) );
  XNOR2_X1 U1751 ( .A(n1556), .B(n1354), .ZN(n1017) );
  XNOR2_X1 U1752 ( .A(n1557), .B(n1365), .ZN(n1016) );
  XNOR2_X1 U1753 ( .A(n1311), .B(n1365), .ZN(n1015) );
  XNOR2_X1 U1754 ( .A(n1551), .B(n1354), .ZN(n1022) );
  XNOR2_X1 U1755 ( .A(n1341), .B(n1365), .ZN(n1021) );
  NAND2_X1 U1756 ( .A1(n156), .A2(n164), .ZN(n154) );
  XNOR2_X1 U1757 ( .A(n1355), .B(n1493), .ZN(n923) );
  XNOR2_X1 U1758 ( .A(n1364), .B(n1493), .ZN(n922) );
  XNOR2_X1 U1759 ( .A(n1346), .B(n1493), .ZN(n924) );
  XNOR2_X1 U1760 ( .A(n1563), .B(n1493), .ZN(n926) );
  XNOR2_X1 U1761 ( .A(n1353), .B(n1493), .ZN(n925) );
  XNOR2_X1 U1762 ( .A(n1562), .B(n1493), .ZN(n927) );
  XNOR2_X1 U1763 ( .A(n1349), .B(n1493), .ZN(n928) );
  XNOR2_X1 U1764 ( .A(n1560), .B(n1493), .ZN(n929) );
  OR2_X1 U1765 ( .A1(n787), .A2(n715), .ZN(n476) );
  XNOR2_X1 U1766 ( .A(n787), .B(n715), .ZN(n477) );
  XNOR2_X1 U1767 ( .A(n1559), .B(n1493), .ZN(n930) );
  XNOR2_X1 U1768 ( .A(n1359), .B(n1492), .ZN(n932) );
  XNOR2_X1 U1769 ( .A(n1311), .B(n1493), .ZN(n931) );
  XNOR2_X1 U1770 ( .A(n1345), .B(n1492), .ZN(n934) );
  XNOR2_X1 U1771 ( .A(n1556), .B(n1493), .ZN(n933) );
  XNOR2_X1 U1772 ( .A(n1548), .B(n1493), .ZN(n941) );
  XNOR2_X1 U1773 ( .A(n1554), .B(n1492), .ZN(n935) );
  XNOR2_X1 U1774 ( .A(n1551), .B(n1492), .ZN(n938) );
  INV_X1 U1775 ( .A(n1492), .ZN(n1142) );
  XNOR2_X1 U1776 ( .A(n1549), .B(n1492), .ZN(n940) );
  XNOR2_X1 U1777 ( .A(n1332), .B(n1493), .ZN(n936) );
  XNOR2_X1 U1778 ( .A(n1552), .B(n1493), .ZN(n937) );
  XNOR2_X1 U1779 ( .A(n1550), .B(n1492), .ZN(n939) );
  INV_X1 U1780 ( .A(n1274), .ZN(n272) );
  NOR2_X1 U1781 ( .A1(n140), .A2(n1274), .ZN(n133) );
  OAI21_X1 U1782 ( .B1(n141), .B2(n135), .A(n136), .ZN(n134) );
  NAND2_X1 U1783 ( .A1(n371), .A2(n382), .ZN(n136) );
  XNOR2_X1 U1784 ( .A(n1331), .B(n1470), .ZN(n1062) );
  INV_X1 U1785 ( .A(n1293), .ZN(n1148) );
  XNOR2_X1 U1786 ( .A(n1556), .B(n1293), .ZN(n1059) );
  XNOR2_X1 U1787 ( .A(n1300), .B(n1293), .ZN(n1067) );
  XNOR2_X1 U1788 ( .A(n1564), .B(n1470), .ZN(n1051) );
  XNOR2_X1 U1789 ( .A(n1563), .B(n1470), .ZN(n1052) );
  XNOR2_X1 U1790 ( .A(n1565), .B(n1470), .ZN(n1050) );
  XNOR2_X1 U1791 ( .A(n1359), .B(n1470), .ZN(n1058) );
  XNOR2_X1 U1792 ( .A(n1566), .B(n1293), .ZN(n1049) );
  XNOR2_X1 U1793 ( .A(n1337), .B(n1293), .ZN(n1066) );
  XNOR2_X1 U1794 ( .A(n1551), .B(n1293), .ZN(n1064) );
  XNOR2_X1 U1795 ( .A(n1310), .B(n1470), .ZN(n1057) );
  XNOR2_X1 U1796 ( .A(n1560), .B(n1470), .ZN(n1055) );
  XNOR2_X1 U1797 ( .A(n1559), .B(n1470), .ZN(n1056) );
  XNOR2_X1 U1798 ( .A(n1550), .B(n1293), .ZN(n1065) );
  XNOR2_X1 U1799 ( .A(n1341), .B(n1293), .ZN(n1063) );
  XNOR2_X1 U1800 ( .A(n1555), .B(n1470), .ZN(n1060) );
  XNOR2_X1 U1801 ( .A(n1305), .B(n1470), .ZN(n1061) );
  XNOR2_X1 U1802 ( .A(n1349), .B(n1470), .ZN(n1054) );
  XNOR2_X1 U1803 ( .A(n1562), .B(n1470), .ZN(n1053) );
  XNOR2_X1 U1804 ( .A(n1567), .B(n1293), .ZN(n1048) );
  XNOR2_X1 U1805 ( .A(n1364), .B(n1545), .ZN(n964) );
  XNOR2_X1 U1806 ( .A(n1355), .B(n1545), .ZN(n965) );
  XNOR2_X1 U1807 ( .A(n1346), .B(n1545), .ZN(n966) );
  XNOR2_X1 U1808 ( .A(n1353), .B(n1545), .ZN(n967) );
  XNOR2_X1 U1809 ( .A(n1559), .B(n1545), .ZN(n972) );
  XNOR2_X1 U1810 ( .A(n1560), .B(n1545), .ZN(n971) );
  XNOR2_X1 U1811 ( .A(n1561), .B(n1545), .ZN(n970) );
  XNOR2_X1 U1812 ( .A(n1562), .B(n1545), .ZN(n969) );
  INV_X1 U1813 ( .A(n1545), .ZN(n1144) );
  XNOR2_X1 U1814 ( .A(n1563), .B(n1545), .ZN(n968) );
  XNOR2_X1 U1815 ( .A(n1555), .B(n1545), .ZN(n976) );
  XNOR2_X1 U1816 ( .A(n1556), .B(n1545), .ZN(n975) );
  XNOR2_X1 U1817 ( .A(n1300), .B(n1545), .ZN(n983) );
  XNOR2_X1 U1818 ( .A(n1310), .B(n1545), .ZN(n973) );
  XNOR2_X1 U1819 ( .A(n1557), .B(n1545), .ZN(n974) );
  XNOR2_X1 U1820 ( .A(n1337), .B(n1545), .ZN(n982) );
  XNOR2_X1 U1821 ( .A(n1330), .B(n1545), .ZN(n978) );
  XNOR2_X1 U1822 ( .A(n1341), .B(n1545), .ZN(n979) );
  XNOR2_X1 U1823 ( .A(n1305), .B(n1545), .ZN(n977) );
  XNOR2_X1 U1824 ( .A(n1551), .B(n1545), .ZN(n980) );
  XNOR2_X1 U1825 ( .A(n1550), .B(n1545), .ZN(n981) );
  NOR2_X1 U1826 ( .A1(n1448), .A2(n180), .ZN(n175) );
  NAND2_X1 U1827 ( .A1(n1511), .A2(n200), .ZN(n81) );
  NAND2_X1 U1828 ( .A1(n202), .A2(n1511), .ZN(n195) );
  AOI21_X1 U1829 ( .B1(n203), .B2(n1511), .A(n1459), .ZN(n196) );
  XNOR2_X1 U1830 ( .A(n1364), .B(n1307), .ZN(n985) );
  XNOR2_X1 U1831 ( .A(n1566), .B(n1307), .ZN(n986) );
  XNOR2_X1 U1832 ( .A(n1563), .B(n1307), .ZN(n989) );
  XNOR2_X1 U1833 ( .A(n1561), .B(n1307), .ZN(n991) );
  XNOR2_X1 U1834 ( .A(n1562), .B(n1307), .ZN(n990) );
  XNOR2_X1 U1835 ( .A(n1300), .B(n1307), .ZN(n1004) );
  XNOR2_X1 U1836 ( .A(n1359), .B(n1307), .ZN(n995) );
  XNOR2_X1 U1837 ( .A(n1337), .B(n1307), .ZN(n1003) );
  XNOR2_X1 U1838 ( .A(n1564), .B(n1307), .ZN(n988) );
  XNOR2_X1 U1839 ( .A(n1565), .B(n1544), .ZN(n987) );
  INV_X1 U1840 ( .A(n1307), .ZN(n1145) );
  XNOR2_X1 U1841 ( .A(n1340), .B(n1544), .ZN(n994) );
  XNOR2_X1 U1842 ( .A(n1551), .B(n1544), .ZN(n1001) );
  XNOR2_X1 U1843 ( .A(n1550), .B(n1307), .ZN(n1002) );
  XNOR2_X1 U1844 ( .A(n1559), .B(n1544), .ZN(n993) );
  XNOR2_X1 U1845 ( .A(n1560), .B(n1544), .ZN(n992) );
  XNOR2_X1 U1846 ( .A(n1332), .B(n1307), .ZN(n999) );
  XNOR2_X1 U1847 ( .A(n1341), .B(n1307), .ZN(n1000) );
  XNOR2_X1 U1848 ( .A(n1554), .B(n1307), .ZN(n998) );
  XNOR2_X1 U1849 ( .A(n1556), .B(n25), .ZN(n996) );
  XNOR2_X1 U1850 ( .A(n1345), .B(n1544), .ZN(n997) );
  INV_X1 U1851 ( .A(n1261), .ZN(n284) );
  NOR2_X1 U1852 ( .A1(n1261), .A2(n209), .ZN(n202) );
  NAND2_X1 U1853 ( .A1(n557), .A2(n568), .ZN(n205) );
  OAI21_X1 U1854 ( .B1(n152), .B2(n1260), .A(n1446), .ZN(n149) );
  OAI21_X1 U1855 ( .B1(n152), .B2(n131), .A(n1456), .ZN(n130) );
  INV_X1 U1856 ( .A(n1260), .ZN(n275) );
  NOR2_X1 U1857 ( .A1(n131), .A2(n128), .ZN(n126) );
  NOR2_X1 U1858 ( .A1(n150), .A2(n1268), .ZN(n145) );
  INV_X1 U1859 ( .A(n1374), .ZN(n220) );
  AOI21_X1 U1860 ( .B1(n221), .B2(n213), .A(n214), .ZN(n212) );
  INV_X1 U1861 ( .A(n1288), .ZN(n1147) );
  XNOR2_X1 U1862 ( .A(n1563), .B(n1288), .ZN(n1031) );
  XNOR2_X1 U1863 ( .A(n1333), .B(n1288), .ZN(n1044) );
  XNOR2_X1 U1864 ( .A(n1561), .B(n1288), .ZN(n1033) );
  XNOR2_X1 U1865 ( .A(n1562), .B(n1288), .ZN(n1032) );
  XNOR2_X1 U1866 ( .A(n1300), .B(n1288), .ZN(n1046) );
  XNOR2_X1 U1867 ( .A(n1556), .B(n1288), .ZN(n1038) );
  XNOR2_X1 U1868 ( .A(n1337), .B(n1288), .ZN(n1045) );
  XNOR2_X1 U1869 ( .A(n1336), .B(n1288), .ZN(n1043) );
  XNOR2_X1 U1870 ( .A(n1359), .B(n1288), .ZN(n1037) );
  XNOR2_X1 U1871 ( .A(n1555), .B(n1288), .ZN(n1039) );
  XNOR2_X1 U1872 ( .A(n1554), .B(n1288), .ZN(n1040) );
  XNOR2_X1 U1873 ( .A(n1331), .B(n1288), .ZN(n1041) );
  XNOR2_X1 U1874 ( .A(n1341), .B(n1288), .ZN(n1042) );
  XNOR2_X1 U1875 ( .A(n1311), .B(n1288), .ZN(n1036) );
  XNOR2_X1 U1876 ( .A(n1559), .B(n1418), .ZN(n1035) );
  XNOR2_X1 U1877 ( .A(n1565), .B(n1418), .ZN(n1029) );
  XNOR2_X1 U1878 ( .A(n1564), .B(n1418), .ZN(n1030) );
  XNOR2_X1 U1879 ( .A(n1560), .B(n1418), .ZN(n1034) );
  XNOR2_X1 U1880 ( .A(n1566), .B(n1418), .ZN(n1028) );
  XNOR2_X1 U1881 ( .A(n1567), .B(n1418), .ZN(n1027) );
  INV_X1 U1882 ( .A(n1487), .ZN(n278) );
  NOR2_X1 U1883 ( .A1(n1487), .A2(n171), .ZN(n164) );
  OAI21_X1 U1884 ( .B1(n166), .B2(n172), .A(n167), .ZN(n165) );
  NAND2_X1 U1885 ( .A1(n461), .A2(n478), .ZN(n167) );
  XOR2_X1 U1886 ( .A(n242), .B(n89), .Z(product[7]) );
  INV_X1 U1887 ( .A(n1398), .ZN(n193) );
  INV_X1 U1888 ( .A(n234), .ZN(n233) );
  AOI21_X1 U1889 ( .B1(n194), .B2(n175), .A(n176), .ZN(n174) );
  OAI21_X1 U1890 ( .B1(n222), .B2(n234), .A(n223), .ZN(n221) );
  OAI21_X1 U1891 ( .B1(n242), .B2(n240), .A(n241), .ZN(n239) );
  INV_X1 U1892 ( .A(n664), .ZN(n840) );
  NAND2_X1 U1893 ( .A1(n1512), .A2(n185), .ZN(n79) );
  OAI21_X1 U1894 ( .B1(n193), .B2(n180), .A(n1451), .ZN(n179) );
  OAI21_X1 U1895 ( .B1(n181), .B2(n177), .A(n178), .ZN(n176) );
  NAND2_X1 U1896 ( .A1(n1512), .A2(n1419), .ZN(n180) );
  AOI21_X1 U1897 ( .B1(n1512), .B2(n1440), .A(n1295), .ZN(n181) );
  INV_X1 U1898 ( .A(n1460), .ZN(n276) );
  OAI22_X1 U1899 ( .A1(n880), .A2(n1483), .B1(n880), .B2(n1455), .ZN(n640) );
  OAI22_X1 U1900 ( .A1(n1483), .A2(n881), .B1(n880), .B2(n1455), .ZN(n298) );
  OAI22_X1 U1901 ( .A1(n1483), .A2(n882), .B1(n881), .B2(n1455), .ZN(n681) );
  OAI22_X1 U1902 ( .A1(n1483), .A2(n883), .B1(n882), .B2(n1455), .ZN(n682) );
  OAI22_X1 U1903 ( .A1(n1483), .A2(n884), .B1(n883), .B2(n1455), .ZN(n683) );
  AOI21_X1 U1904 ( .B1(n156), .B2(n165), .A(n157), .ZN(n155) );
  NOR2_X1 U1905 ( .A1(n161), .A2(n1460), .ZN(n156) );
  OAI21_X1 U1906 ( .B1(n162), .B2(n158), .A(n159), .ZN(n157) );
  OAI22_X1 U1907 ( .A1(n1483), .A2(n886), .B1(n885), .B2(n1455), .ZN(n685) );
  OAI22_X1 U1908 ( .A1(n1483), .A2(n885), .B1(n884), .B2(n1455), .ZN(n684) );
  OAI22_X1 U1909 ( .A1(n1483), .A2(n887), .B1(n886), .B2(n1455), .ZN(n686) );
  OAI22_X1 U1910 ( .A1(n1483), .A2(n888), .B1(n887), .B2(n1455), .ZN(n687) );
  OAI22_X1 U1911 ( .A1(n1483), .A2(n889), .B1(n888), .B2(n1455), .ZN(n688) );
  OAI22_X1 U1912 ( .A1(n1483), .A2(n890), .B1(n889), .B2(n1455), .ZN(n689) );
  OAI22_X1 U1913 ( .A1(n1317), .A2(n891), .B1(n890), .B2(n1455), .ZN(n690) );
  OAI22_X1 U1914 ( .A1(n1318), .A2(n892), .B1(n891), .B2(n1320), .ZN(n691) );
  OAI22_X1 U1915 ( .A1(n1317), .A2(n894), .B1(n893), .B2(n1321), .ZN(n693) );
  OAI22_X1 U1916 ( .A1(n1318), .A2(n893), .B1(n892), .B2(n1320), .ZN(n692) );
  OAI22_X1 U1917 ( .A1(n1317), .A2(n895), .B1(n894), .B2(n1321), .ZN(n694) );
  OAI22_X1 U1918 ( .A1(n1318), .A2(n899), .B1(n898), .B2(n1320), .ZN(n698) );
  OAI22_X1 U1919 ( .A1(n1317), .A2(n1140), .B1(n900), .B2(n1320), .ZN(n670) );
  OAI22_X1 U1920 ( .A1(n1317), .A2(n896), .B1(n895), .B2(n1321), .ZN(n695) );
  INV_X1 U1921 ( .A(n1320), .ZN(n641) );
  INV_X1 U1922 ( .A(n1375), .ZN(n211) );
  INV_X1 U1923 ( .A(n1308), .ZN(n173) );
  OAI21_X1 U1924 ( .B1(n212), .B2(n195), .A(n196), .ZN(n194) );
  OAI22_X1 U1925 ( .A1(n1323), .A2(n1055), .B1(n1054), .B2(n1262), .ZN(n846)
         );
  OAI22_X1 U1926 ( .A1(n1304), .A2(n1062), .B1(n1061), .B2(n1262), .ZN(n853)
         );
  OAI22_X1 U1927 ( .A1(n1304), .A2(n1059), .B1(n1058), .B2(n1262), .ZN(n850)
         );
  OAI22_X1 U1928 ( .A1(n1323), .A2(n1060), .B1(n1059), .B2(n1262), .ZN(n851)
         );
  OAI22_X1 U1929 ( .A1(n1367), .A2(n1053), .B1(n1052), .B2(n1530), .ZN(n844)
         );
  OAI22_X1 U1930 ( .A1(n1322), .A2(n1051), .B1(n1050), .B2(n1530), .ZN(n842)
         );
  OAI22_X1 U1931 ( .A1(n1304), .A2(n1148), .B1(n1068), .B2(n1262), .ZN(n678)
         );
  OAI22_X1 U1932 ( .A1(n1367), .A2(n1063), .B1(n1062), .B2(n1262), .ZN(n854)
         );
  OAI22_X1 U1933 ( .A1(n1323), .A2(n1065), .B1(n1064), .B2(n1262), .ZN(n856)
         );
  OAI22_X1 U1934 ( .A1(n1322), .A2(n1049), .B1(n1048), .B2(n1530), .ZN(n458)
         );
  OAI22_X1 U1935 ( .A1(n1367), .A2(n1052), .B1(n1051), .B2(n1530), .ZN(n843)
         );
  OAI22_X1 U1936 ( .A1(n1050), .A2(n1366), .B1(n1049), .B2(n1530), .ZN(n841)
         );
  OAI22_X1 U1937 ( .A1(n1323), .A2(n1057), .B1(n1056), .B2(n1530), .ZN(n848)
         );
  OAI22_X1 U1938 ( .A1(n1323), .A2(n1056), .B1(n1055), .B2(n1530), .ZN(n847)
         );
  OAI22_X1 U1939 ( .A1(n1367), .A2(n1058), .B1(n1057), .B2(n1530), .ZN(n849)
         );
  OAI22_X1 U1940 ( .A1(n1367), .A2(n1054), .B1(n1053), .B2(n1530), .ZN(n845)
         );
  OAI22_X1 U1941 ( .A1(n1323), .A2(n1067), .B1(n1066), .B2(n1530), .ZN(n858)
         );
  OAI22_X1 U1942 ( .A1(n1367), .A2(n1061), .B1(n1060), .B2(n1530), .ZN(n852)
         );
  OAI22_X1 U1943 ( .A1(n1048), .A2(n1366), .B1(n1048), .B2(n1530), .ZN(n664)
         );
  OAI22_X1 U1944 ( .A1(n1367), .A2(n1066), .B1(n1065), .B2(n1530), .ZN(n857)
         );
  OAI22_X1 U1945 ( .A1(n1367), .A2(n1064), .B1(n1063), .B2(n1530), .ZN(n855)
         );
  INV_X1 U1946 ( .A(n1530), .ZN(n665) );
  OAI21_X1 U1947 ( .B1(n248), .B2(n250), .A(n249), .ZN(n247) );
  INV_X1 U1948 ( .A(n254), .ZN(n252) );
  AOI21_X1 U1949 ( .B1(n1501), .B2(n1301), .A(n1495), .ZN(n125) );
  OAI21_X1 U1950 ( .B1(n132), .B2(n128), .A(n129), .ZN(n127) );
  OAI21_X1 U1951 ( .B1(n174), .B2(n154), .A(n155), .ZN(n153) );
  OAI21_X1 U1952 ( .B1(n151), .B2(n147), .A(n148), .ZN(n146) );
  OAI22_X1 U1953 ( .A1(n901), .A2(n1447), .B1(n901), .B2(n1357), .ZN(n643) );
  OAI22_X1 U1954 ( .A1(n1447), .A2(n902), .B1(n901), .B2(n1358), .ZN(n304) );
  OAI22_X1 U1955 ( .A1(n1447), .A2(n903), .B1(n902), .B2(n1357), .ZN(n701) );
  OAI22_X1 U1956 ( .A1(n1447), .A2(n905), .B1(n904), .B2(n1357), .ZN(n703) );
  OAI22_X1 U1957 ( .A1(n1447), .A2(n904), .B1(n903), .B2(n1358), .ZN(n702) );
  OAI22_X1 U1958 ( .A1(n1447), .A2(n906), .B1(n905), .B2(n1358), .ZN(n704) );
  OAI22_X1 U1959 ( .A1(n1447), .A2(n907), .B1(n906), .B2(n1357), .ZN(n705) );
  OAI22_X1 U1960 ( .A1(n1447), .A2(n908), .B1(n907), .B2(n1358), .ZN(n706) );
  OAI22_X1 U1961 ( .A1(n1447), .A2(n909), .B1(n908), .B2(n1357), .ZN(n707) );
  OAI22_X1 U1962 ( .A1(n54), .A2(n910), .B1(n909), .B2(n1358), .ZN(n708) );
  OAI22_X1 U1963 ( .A1(n54), .A2(n911), .B1(n910), .B2(n1357), .ZN(n709) );
  OAI22_X1 U1964 ( .A1(n54), .A2(n915), .B1(n914), .B2(n1357), .ZN(n713) );
  OAI22_X1 U1965 ( .A1(n54), .A2(n912), .B1(n911), .B2(n1358), .ZN(n710) );
  OAI22_X1 U1966 ( .A1(n54), .A2(n913), .B1(n912), .B2(n1358), .ZN(n711) );
  OAI22_X1 U1967 ( .A1(n54), .A2(n914), .B1(n913), .B2(n1357), .ZN(n712) );
  OAI22_X1 U1968 ( .A1(n54), .A2(n1141), .B1(n921), .B2(n1358), .ZN(n671) );
  OAI22_X1 U1969 ( .A1(n54), .A2(n918), .B1(n917), .B2(n1357), .ZN(n716) );
  OAI22_X1 U1970 ( .A1(n54), .A2(n919), .B1(n918), .B2(n1357), .ZN(n717) );
  OAI22_X1 U1971 ( .A1(n54), .A2(n917), .B1(n916), .B2(n1358), .ZN(n715) );
  OAI22_X1 U1972 ( .A1(n916), .A2(n54), .B1(n915), .B2(n1358), .ZN(n714) );
  OAI22_X1 U1973 ( .A1(n54), .A2(n920), .B1(n919), .B2(n1357), .ZN(n718) );
  OAI22_X1 U1974 ( .A1(n1452), .A2(n965), .B1(n964), .B2(n1449), .ZN(n346) );
  OAI22_X1 U1975 ( .A1(n964), .A2(n1452), .B1(n964), .B2(n1449), .ZN(n652) );
  OAI22_X1 U1976 ( .A1(n1452), .A2(n966), .B1(n965), .B2(n1449), .ZN(n761) );
  OAI22_X1 U1977 ( .A1(n1452), .A2(n967), .B1(n966), .B2(n1449), .ZN(n762) );
  OAI22_X1 U1978 ( .A1(n1452), .A2(n968), .B1(n967), .B2(n1449), .ZN(n763) );
  OAI22_X1 U1979 ( .A1(n1452), .A2(n973), .B1(n972), .B2(n1372), .ZN(n768) );
  OAI22_X1 U1980 ( .A1(n1452), .A2(n972), .B1(n971), .B2(n1372), .ZN(n767) );
  OAI22_X1 U1981 ( .A1(n1452), .A2(n975), .B1(n974), .B2(n1372), .ZN(n770) );
  OAI22_X1 U1982 ( .A1(n1452), .A2(n969), .B1(n968), .B2(n1372), .ZN(n764) );
  OAI22_X1 U1983 ( .A1(n1452), .A2(n971), .B1(n970), .B2(n1372), .ZN(n766) );
  OAI22_X1 U1984 ( .A1(n1452), .A2(n977), .B1(n976), .B2(n1372), .ZN(n772) );
  OAI22_X1 U1985 ( .A1(n1453), .A2(n970), .B1(n969), .B2(n1372), .ZN(n765) );
  OAI22_X1 U1986 ( .A1(n1452), .A2(n1144), .B1(n984), .B2(n1372), .ZN(n674) );
  OAI22_X1 U1987 ( .A1(n1453), .A2(n983), .B1(n982), .B2(n1372), .ZN(n778) );
  OAI22_X1 U1988 ( .A1(n1453), .A2(n976), .B1(n975), .B2(n1372), .ZN(n771) );
  OAI22_X1 U1989 ( .A1(n1453), .A2(n974), .B1(n973), .B2(n1372), .ZN(n769) );
  OAI22_X1 U1990 ( .A1(n1453), .A2(n982), .B1(n981), .B2(n1372), .ZN(n777) );
  OAI22_X1 U1991 ( .A1(n1453), .A2(n979), .B1(n978), .B2(n1372), .ZN(n774) );
  OAI22_X1 U1992 ( .A1(n1453), .A2(n980), .B1(n979), .B2(n1372), .ZN(n775) );
  OAI22_X1 U1993 ( .A1(n1453), .A2(n978), .B1(n977), .B2(n1372), .ZN(n773) );
  OAI22_X1 U1994 ( .A1(n1453), .A2(n981), .B1(n980), .B2(n1372), .ZN(n776) );
  INV_X1 U1995 ( .A(n1372), .ZN(n653) );
  OAI22_X1 U1996 ( .A1(n922), .A2(n1350), .B1(n922), .B2(n1343), .ZN(n646) );
  OAI22_X1 U1997 ( .A1(n1350), .A2(n924), .B1(n923), .B2(n1524), .ZN(n721) );
  OAI22_X1 U1998 ( .A1(n1350), .A2(n923), .B1(n922), .B2(n1524), .ZN(n314) );
  OAI22_X1 U1999 ( .A1(n1350), .A2(n925), .B1(n924), .B2(n1524), .ZN(n722) );
  OAI22_X1 U2000 ( .A1(n1350), .A2(n927), .B1(n926), .B2(n1524), .ZN(n724) );
  OAI22_X1 U2001 ( .A1(n1350), .A2(n926), .B1(n925), .B2(n1343), .ZN(n723) );
  OAI22_X1 U2002 ( .A1(n1350), .A2(n928), .B1(n927), .B2(n1524), .ZN(n725) );
  OAI22_X1 U2003 ( .A1(n1350), .A2(n929), .B1(n928), .B2(n1343), .ZN(n726) );
  OAI22_X1 U2004 ( .A1(n1370), .A2(n930), .B1(n929), .B2(n1524), .ZN(n727) );
  OAI22_X1 U2005 ( .A1(n1370), .A2(n931), .B1(n930), .B2(n1524), .ZN(n728) );
  OAI22_X1 U2006 ( .A1(n1370), .A2(n933), .B1(n932), .B2(n1524), .ZN(n730) );
  OAI22_X1 U2007 ( .A1(n1370), .A2(n934), .B1(n933), .B2(n1524), .ZN(n731) );
  OAI22_X1 U2008 ( .A1(n1370), .A2(n932), .B1(n931), .B2(n1524), .ZN(n729) );
  OAI22_X1 U2009 ( .A1(n936), .A2(n1370), .B1(n935), .B2(n1343), .ZN(n733) );
  OAI22_X1 U2010 ( .A1(n1370), .A2(n937), .B1(n936), .B2(n1524), .ZN(n734) );
  OAI22_X1 U2011 ( .A1(n1370), .A2(n1142), .B1(n942), .B2(n1524), .ZN(n672) );
  OAI22_X1 U2012 ( .A1(n1369), .A2(n935), .B1(n934), .B2(n46), .ZN(n732) );
  OAI22_X1 U2013 ( .A1(n1370), .A2(n941), .B1(n940), .B2(n1343), .ZN(n738) );
  OAI22_X1 U2014 ( .A1(n1370), .A2(n938), .B1(n937), .B2(n1524), .ZN(n735) );
  INV_X1 U2015 ( .A(n1524), .ZN(n647) );
  OAI22_X1 U2016 ( .A1(n1369), .A2(n939), .B1(n938), .B2(n1343), .ZN(n736) );
  OAI22_X1 U2017 ( .A1(n1369), .A2(n940), .B1(n939), .B2(n46), .ZN(n737) );
  OAI22_X1 U2018 ( .A1(n985), .A2(n1461), .B1(n985), .B2(n1428), .ZN(n655) );
  OAI22_X1 U2019 ( .A1(n1463), .A2(n986), .B1(n985), .B2(n1428), .ZN(n368) );
  OAI22_X1 U2020 ( .A1(n1463), .A2(n987), .B1(n986), .B2(n1428), .ZN(n781) );
  OAI22_X1 U2021 ( .A1(n1463), .A2(n992), .B1(n991), .B2(n1428), .ZN(n786) );
  OAI22_X1 U2022 ( .A1(n1461), .A2(n1003), .B1(n1002), .B2(n1428), .ZN(n797)
         );
  OAI22_X1 U2023 ( .A1(n1463), .A2(n989), .B1(n988), .B2(n1428), .ZN(n783) );
  OAI22_X1 U2024 ( .A1(n1461), .A2(n990), .B1(n989), .B2(n1428), .ZN(n784) );
  OAI22_X1 U2025 ( .A1(n1463), .A2(n991), .B1(n990), .B2(n1428), .ZN(n785) );
  OAI22_X1 U2026 ( .A1(n1463), .A2(n996), .B1(n995), .B2(n1428), .ZN(n790) );
  OAI22_X1 U2027 ( .A1(n1463), .A2(n988), .B1(n987), .B2(n1529), .ZN(n782) );
  OAI22_X1 U2028 ( .A1(n1461), .A2(n999), .B1(n998), .B2(n1428), .ZN(n793) );
  OAI22_X1 U2029 ( .A1(n1462), .A2(n994), .B1(n1529), .B2(n993), .ZN(n788) );
  OAI22_X1 U2030 ( .A1(n1462), .A2(n993), .B1(n992), .B2(n1529), .ZN(n787) );
  OAI22_X1 U2031 ( .A1(n1461), .A2(n1000), .B1(n999), .B2(n1428), .ZN(n794) );
  OAI22_X1 U2032 ( .A1(n1463), .A2(n995), .B1(n994), .B2(n1529), .ZN(n789) );
  OAI22_X1 U2033 ( .A1(n1461), .A2(n1002), .B1(n1001), .B2(n1428), .ZN(n796)
         );
  OAI22_X1 U2034 ( .A1(n1463), .A2(n1004), .B1(n1003), .B2(n1428), .ZN(n798)
         );
  INV_X1 U2035 ( .A(n1428), .ZN(n656) );
  OAI22_X1 U2036 ( .A1(n1463), .A2(n1145), .B1(n1005), .B2(n1428), .ZN(n675)
         );
  OAI22_X1 U2037 ( .A1(n1463), .A2(n1001), .B1(n1000), .B2(n1428), .ZN(n795)
         );
  OAI22_X1 U2038 ( .A1(n1463), .A2(n998), .B1(n997), .B2(n1529), .ZN(n792) );
  OAI22_X1 U2039 ( .A1(n1462), .A2(n997), .B1(n996), .B2(n1529), .ZN(n791) );
  OAI22_X1 U2040 ( .A1(n943), .A2(n1342), .B1(n943), .B2(n1525), .ZN(n649) );
  OAI22_X1 U2041 ( .A1(n1342), .A2(n944), .B1(n943), .B2(n1526), .ZN(n328) );
  OAI22_X1 U2042 ( .A1(n1342), .A2(n945), .B1(n944), .B2(n1525), .ZN(n741) );
  OAI22_X1 U2043 ( .A1(n1342), .A2(n947), .B1(n946), .B2(n1526), .ZN(n743) );
  OAI22_X1 U2044 ( .A1(n1342), .A2(n946), .B1(n945), .B2(n1525), .ZN(n742) );
  OAI22_X1 U2045 ( .A1(n1342), .A2(n948), .B1(n947), .B2(n1526), .ZN(n744) );
  OAI22_X1 U2046 ( .A1(n1504), .A2(n949), .B1(n948), .B2(n1525), .ZN(n745) );
  OAI22_X1 U2047 ( .A1(n1504), .A2(n957), .B1(n1258), .B2(n1525), .ZN(n753) );
  OAI22_X1 U2048 ( .A1(n1504), .A2(n952), .B1(n951), .B2(n1526), .ZN(n748) );
  OAI22_X1 U2049 ( .A1(n1504), .A2(n1263), .B1(n952), .B2(n1525), .ZN(n749) );
  OAI22_X1 U2050 ( .A1(n956), .A2(n1504), .B1(n1234), .B2(n1525), .ZN(n752) );
  OAI22_X1 U2051 ( .A1(n951), .A2(n1504), .B1(n950), .B2(n1526), .ZN(n747) );
  OAI22_X1 U2052 ( .A1(n950), .A2(n1504), .B1(n949), .B2(n1525), .ZN(n746) );
  OAI22_X1 U2053 ( .A1(n1503), .A2(n958), .B1(n957), .B2(n1526), .ZN(n754) );
  OAI22_X1 U2054 ( .A1(n1504), .A2(n1143), .B1(n963), .B2(n1526), .ZN(n673) );
  OAI22_X1 U2055 ( .A1(n1503), .A2(n955), .B1(n1276), .B2(n1526), .ZN(n751) );
  OAI22_X1 U2056 ( .A1(n1504), .A2(n961), .B1(n960), .B2(n1525), .ZN(n757) );
  OAI22_X1 U2057 ( .A1(n1504), .A2(n960), .B1(n959), .B2(n1526), .ZN(n756) );
  OAI22_X1 U2058 ( .A1(n1503), .A2(n954), .B1(n953), .B2(n1525), .ZN(n750) );
  INV_X1 U2059 ( .A(n1525), .ZN(n650) );
  OAI22_X1 U2060 ( .A1(n1503), .A2(n962), .B1(n961), .B2(n1526), .ZN(n758) );
  OAI22_X1 U2061 ( .A1(n1503), .A2(n959), .B1(n958), .B2(n1526), .ZN(n755) );
  BUF_X4 U2062 ( .A(n31), .Z(n1545) );
  XNOR2_X1 U2063 ( .A(n1469), .B(n65), .ZN(product[31]) );
  XNOR2_X1 U2064 ( .A(n1481), .B(n67), .ZN(product[29]) );
  INV_X1 U2065 ( .A(n101), .ZN(n264) );
  AOI21_X1 U2066 ( .B1(n114), .B2(n1516), .A(n111), .ZN(n109) );
  AOI21_X1 U2067 ( .B1(n1481), .B2(n1517), .A(n119), .ZN(n117) );
  OAI22_X1 U2068 ( .A1(n1344), .A2(n1014), .B1(n1013), .B2(n1445), .ZN(n807)
         );
  OAI22_X1 U2069 ( .A1(n1465), .A2(n1007), .B1(n1006), .B2(n1445), .ZN(n394)
         );
  OAI22_X1 U2070 ( .A1(n1465), .A2(n1012), .B1(n1011), .B2(n1445), .ZN(n805)
         );
  OAI22_X1 U2071 ( .A1(n1006), .A2(n1344), .B1(n1006), .B2(n1445), .ZN(n658)
         );
  OAI22_X1 U2072 ( .A1(n1465), .A2(n1021), .B1(n1020), .B2(n1445), .ZN(n814)
         );
  OAI22_X1 U2073 ( .A1(n1344), .A2(n1024), .B1(n1023), .B2(n1445), .ZN(n817)
         );
  OAI22_X1 U2074 ( .A1(n1465), .A2(n1010), .B1(n1009), .B2(n1445), .ZN(n803)
         );
  OAI22_X1 U2075 ( .A1(n1465), .A2(n1008), .B1(n1007), .B2(n1445), .ZN(n801)
         );
  OAI22_X1 U2076 ( .A1(n1465), .A2(n1239), .B1(n1014), .B2(n1445), .ZN(n808)
         );
  OAI22_X1 U2077 ( .A1(n1465), .A2(n1009), .B1(n1008), .B2(n1445), .ZN(n802)
         );
  OAI22_X1 U2078 ( .A1(n1344), .A2(n1373), .B1(n1026), .B2(n1445), .ZN(n676)
         );
  OAI22_X1 U2079 ( .A1(n24), .A2(n1013), .B1(n1012), .B2(n1527), .ZN(n806) );
  OAI22_X1 U2080 ( .A1(n1465), .A2(n1025), .B1(n1024), .B2(n1445), .ZN(n818)
         );
  OAI22_X1 U2081 ( .A1(n1465), .A2(n1019), .B1(n1018), .B2(n1445), .ZN(n812)
         );
  OAI22_X1 U2082 ( .A1(n1465), .A2(n1020), .B1(n1019), .B2(n1527), .ZN(n813)
         );
  OAI22_X1 U2083 ( .A1(n1465), .A2(n1018), .B1(n1017), .B2(n1445), .ZN(n811)
         );
  OAI22_X1 U2084 ( .A1(n24), .A2(n1011), .B1(n1010), .B2(n1527), .ZN(n804) );
  OAI22_X1 U2085 ( .A1(n1465), .A2(n1017), .B1(n1016), .B2(n1445), .ZN(n810)
         );
  OAI22_X1 U2086 ( .A1(n1465), .A2(n1023), .B1(n1022), .B2(n1445), .ZN(n816)
         );
  OAI22_X1 U2087 ( .A1(n24), .A2(n1016), .B1(n1239), .B2(n1445), .ZN(n809) );
  OAI22_X1 U2088 ( .A1(n24), .A2(n1022), .B1(n1021), .B2(n1527), .ZN(n815) );
  INV_X1 U2089 ( .A(n1527), .ZN(n659) );
  XNOR2_X1 U2090 ( .A(n1468), .B(n63), .ZN(product[33]) );
  XOR2_X1 U2091 ( .A(n1480), .B(n64), .Z(product[32]) );
  XOR2_X1 U2092 ( .A(n117), .B(n66), .Z(product[30]) );
  XOR2_X1 U2093 ( .A(n125), .B(n68), .Z(product[28]) );
  AOI21_X1 U2094 ( .B1(n106), .B2(n1518), .A(n103), .ZN(n101) );
  OAI21_X1 U2095 ( .B1(n1500), .B2(n115), .A(n116), .ZN(n114) );
  OAI21_X1 U2096 ( .B1(n1502), .B2(n123), .A(n124), .ZN(n122) );
  OAI22_X1 U2097 ( .A1(n1324), .A2(n1039), .B1(n1038), .B2(n1334), .ZN(n831)
         );
  OAI22_X1 U2098 ( .A1(n1438), .A2(n1031), .B1(n1030), .B2(n1334), .ZN(n823)
         );
  OAI22_X1 U2099 ( .A1(n1324), .A2(n1041), .B1(n1040), .B2(n1334), .ZN(n833)
         );
  OAI22_X1 U2100 ( .A1(n1437), .A2(n1032), .B1(n1031), .B2(n1528), .ZN(n824)
         );
  OAI22_X1 U2101 ( .A1(n1324), .A2(n1034), .B1(n1033), .B2(n1528), .ZN(n826)
         );
  OAI22_X1 U2102 ( .A1(n1438), .A2(n1045), .B1(n1044), .B2(n1528), .ZN(n837)
         );
  OAI22_X1 U2103 ( .A1(n1438), .A2(n1038), .B1(n1037), .B2(n1334), .ZN(n830)
         );
  OAI22_X1 U2104 ( .A1(n1438), .A2(n1044), .B1(n1043), .B2(n1528), .ZN(n836)
         );
  OAI22_X1 U2105 ( .A1(n1471), .A2(n1040), .B1(n1039), .B2(n1334), .ZN(n832)
         );
  OAI22_X1 U2106 ( .A1(n1438), .A2(n1028), .B1(n1027), .B2(n1528), .ZN(n424)
         );
  OAI22_X1 U2107 ( .A1(n1438), .A2(n1037), .B1(n1036), .B2(n1528), .ZN(n829)
         );
  OAI22_X1 U2108 ( .A1(n1471), .A2(n1030), .B1(n1029), .B2(n1334), .ZN(n822)
         );
  OAI22_X1 U2109 ( .A1(n1471), .A2(n1033), .B1(n1032), .B2(n1528), .ZN(n825)
         );
  OAI22_X1 U2110 ( .A1(n1438), .A2(n1147), .B1(n1047), .B2(n1528), .ZN(n677)
         );
  OAI22_X1 U2111 ( .A1(n1027), .A2(n1471), .B1(n1027), .B2(n1334), .ZN(n661)
         );
  OAI22_X1 U2112 ( .A1(n1324), .A2(n1043), .B1(n1042), .B2(n1528), .ZN(n835)
         );
  OAI22_X1 U2113 ( .A1(n1437), .A2(n1029), .B1(n1028), .B2(n1528), .ZN(n821)
         );
  OAI22_X1 U2114 ( .A1(n1471), .A2(n1036), .B1(n1035), .B2(n1334), .ZN(n828)
         );
  OAI22_X1 U2115 ( .A1(n1438), .A2(n1042), .B1(n1041), .B2(n1334), .ZN(n834)
         );
  OAI22_X1 U2116 ( .A1(n1438), .A2(n1035), .B1(n1034), .B2(n1528), .ZN(n827)
         );
  OAI22_X1 U2117 ( .A1(n1324), .A2(n1046), .B1(n1045), .B2(n1334), .ZN(n838)
         );
  INV_X1 U2118 ( .A(n1528), .ZN(n662) );
  OAI21_X1 U2119 ( .B1(n109), .B2(n107), .A(n108), .ZN(n106) );
endmodule


module mac_6_DW01_add_1 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n34, n35, n36, n37, n38, n39, n40, n41, n43, n45, n46, n47,
         n48, n49, n51, n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65,
         n67, n69, n70, n71, n72, n73, n75, n77, n78, n79, n80, n81, n83, n85,
         n86, n87, n88, n89, n91, n93, n94, n95, n96, n97, n99, n101, n102,
         n103, n104, n105, n107, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n119, n121, n122, n124, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n184, n185, n187, n189, n191,
         n193, n195, n197, n199, n201, n203, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409;

  FA_X1 U3 ( .A(B[38]), .B(A[38]), .CI(n35), .CO(n34), .S(SUM[38]) );
  FA_X1 U8 ( .A(B[33]), .B(A[33]), .CI(n40), .CO(n39), .S(SUM[33]) );
  FA_X1 U9 ( .A(B[32]), .B(A[32]), .CI(n185), .CO(n40), .S(SUM[32]) );
  NAND2_X1 U254 ( .A1(B[36]), .A2(A[36]), .ZN(n379) );
  NAND2_X1 U255 ( .A1(B[2]), .A2(A[2]), .ZN(n178) );
  INV_X1 U256 ( .A(n149), .ZN(n344) );
  OR2_X1 U257 ( .A1(B[11]), .A2(A[11]), .ZN(n345) );
  OR2_X1 U258 ( .A1(B[0]), .A2(A[0]), .ZN(n346) );
  CLKBUF_X1 U259 ( .A(n39), .Z(n347) );
  NAND3_X1 U260 ( .A1(n351), .A2(n352), .A3(n353), .ZN(n348) );
  NAND3_X1 U261 ( .A1(n351), .A2(n352), .A3(n353), .ZN(n349) );
  XOR2_X1 U262 ( .A(B[34]), .B(A[34]), .Z(n350) );
  XOR2_X1 U263 ( .A(n347), .B(n350), .Z(SUM[34]) );
  NAND2_X1 U264 ( .A1(n39), .A2(B[34]), .ZN(n351) );
  NAND2_X1 U265 ( .A1(n39), .A2(A[34]), .ZN(n352) );
  NAND2_X1 U266 ( .A1(B[34]), .A2(A[34]), .ZN(n353) );
  NAND3_X1 U267 ( .A1(n351), .A2(n352), .A3(n353), .ZN(n38) );
  NAND3_X1 U268 ( .A1(n356), .A2(n357), .A3(n358), .ZN(n354) );
  XOR2_X1 U269 ( .A(B[35]), .B(A[35]), .Z(n355) );
  XOR2_X1 U270 ( .A(n349), .B(n355), .Z(SUM[35]) );
  NAND2_X1 U271 ( .A1(n348), .A2(B[35]), .ZN(n356) );
  NAND2_X1 U272 ( .A1(n38), .A2(A[35]), .ZN(n357) );
  NAND2_X1 U273 ( .A1(B[35]), .A2(A[35]), .ZN(n358) );
  NAND3_X1 U274 ( .A1(n356), .A2(n357), .A3(n358), .ZN(n37) );
  CLKBUF_X1 U275 ( .A(n94), .Z(n359) );
  CLKBUF_X1 U276 ( .A(n70), .Z(n360) );
  CLKBUF_X1 U277 ( .A(n115), .Z(n361) );
  NOR2_X1 U278 ( .A1(B[7]), .A2(A[7]), .ZN(n362) );
  NOR2_X1 U279 ( .A1(B[7]), .A2(A[7]), .ZN(n155) );
  CLKBUF_X1 U280 ( .A(n380), .Z(n363) );
  CLKBUF_X1 U281 ( .A(n37), .Z(n364) );
  AOI21_X1 U282 ( .B1(n359), .B2(n400), .A(n91), .ZN(n365) );
  AOI21_X1 U283 ( .B1(n94), .B2(n400), .A(n91), .ZN(n89) );
  AOI21_X1 U284 ( .B1(n360), .B2(n406), .A(n67), .ZN(n366) );
  AOI21_X1 U285 ( .B1(n70), .B2(n406), .A(n67), .ZN(n65) );
  CLKBUF_X1 U286 ( .A(n171), .Z(n367) );
  AOI21_X1 U287 ( .B1(n344), .B2(n114), .A(n361), .ZN(n368) );
  AOI21_X1 U288 ( .B1(n150), .B2(n114), .A(n115), .ZN(n113) );
  AOI21_X1 U289 ( .B1(n143), .B2(n130), .A(n131), .ZN(n369) );
  CLKBUF_X1 U290 ( .A(n62), .Z(n370) );
  NOR2_X1 U291 ( .A1(B[5]), .A2(A[5]), .ZN(n371) );
  CLKBUF_X1 U292 ( .A(n110), .Z(n372) );
  NAND3_X1 U293 ( .A1(n380), .A2(n381), .A3(n379), .ZN(n373) );
  NAND3_X1 U294 ( .A1(n379), .A2(n363), .A3(n381), .ZN(n374) );
  CLKBUF_X1 U295 ( .A(n54), .Z(n375) );
  CLKBUF_X1 U296 ( .A(n102), .Z(n376) );
  NOR2_X1 U297 ( .A1(B[9]), .A2(A[9]), .ZN(n377) );
  NOR2_X1 U298 ( .A1(B[9]), .A2(A[9]), .ZN(n144) );
  XOR2_X1 U299 ( .A(B[36]), .B(A[36]), .Z(n378) );
  XOR2_X1 U300 ( .A(n378), .B(n364), .Z(SUM[36]) );
  NAND2_X1 U301 ( .A1(B[36]), .A2(n37), .ZN(n380) );
  NAND2_X1 U302 ( .A1(A[36]), .A2(n354), .ZN(n381) );
  NAND3_X1 U303 ( .A1(n380), .A2(n381), .A3(n379), .ZN(n36) );
  XOR2_X1 U304 ( .A(B[37]), .B(A[37]), .Z(n382) );
  XOR2_X1 U305 ( .A(n382), .B(n374), .Z(SUM[37]) );
  NAND2_X1 U306 ( .A1(B[37]), .A2(A[37]), .ZN(n383) );
  NAND2_X1 U307 ( .A1(B[37]), .A2(n373), .ZN(n384) );
  NAND2_X1 U308 ( .A1(A[37]), .A2(n36), .ZN(n385) );
  NAND3_X1 U309 ( .A1(n383), .A2(n384), .A3(n385), .ZN(n35) );
  NOR2_X1 U310 ( .A1(B[3]), .A2(A[3]), .ZN(n386) );
  NOR2_X1 U311 ( .A1(B[3]), .A2(A[3]), .ZN(n174) );
  NOR2_X1 U312 ( .A1(B[11]), .A2(A[11]), .ZN(n387) );
  AOI21_X1 U313 ( .B1(n372), .B2(n401), .A(n107), .ZN(n388) );
  NOR2_X1 U314 ( .A1(B[11]), .A2(A[11]), .ZN(n132) );
  AOI21_X1 U315 ( .B1(n110), .B2(n401), .A(n107), .ZN(n105) );
  CLKBUF_X1 U316 ( .A(n46), .Z(n389) );
  AOI21_X1 U317 ( .B1(n375), .B2(n407), .A(n51), .ZN(n390) );
  CLKBUF_X1 U318 ( .A(n86), .Z(n391) );
  CLKBUF_X1 U319 ( .A(n78), .Z(n392) );
  AOI21_X1 U320 ( .B1(n376), .B2(n402), .A(n99), .ZN(n393) );
  AOI21_X1 U321 ( .B1(n392), .B2(n404), .A(n75), .ZN(n394) );
  AOI21_X1 U322 ( .B1(n370), .B2(n405), .A(n59), .ZN(n395) );
  AOI21_X1 U323 ( .B1(n391), .B2(n403), .A(n83), .ZN(n396) );
  OAI21_X1 U324 ( .B1(n149), .B2(n140), .A(n141), .ZN(n139) );
  INV_X1 U325 ( .A(n143), .ZN(n141) );
  INV_X1 U326 ( .A(n142), .ZN(n140) );
  NAND2_X1 U327 ( .A1(n142), .A2(n130), .ZN(n128) );
  AOI21_X1 U328 ( .B1(n170), .B2(n161), .A(n162), .ZN(n160) );
  INV_X1 U329 ( .A(n367), .ZN(n170) );
  INV_X1 U330 ( .A(n180), .ZN(n179) );
  INV_X1 U331 ( .A(n85), .ZN(n83) );
  INV_X1 U332 ( .A(n77), .ZN(n75) );
  INV_X1 U333 ( .A(n69), .ZN(n67) );
  INV_X1 U334 ( .A(n53), .ZN(n51) );
  NAND2_X1 U335 ( .A1(n161), .A2(n153), .ZN(n151) );
  AOI21_X1 U336 ( .B1(n153), .B2(n162), .A(n154), .ZN(n152) );
  NOR2_X1 U337 ( .A1(n158), .A2(n362), .ZN(n153) );
  AOI21_X1 U338 ( .B1(n62), .B2(n405), .A(n59), .ZN(n57) );
  INV_X1 U339 ( .A(n61), .ZN(n59) );
  OAI21_X1 U340 ( .B1(n163), .B2(n169), .A(n164), .ZN(n162) );
  INV_X1 U341 ( .A(n109), .ZN(n107) );
  AOI21_X1 U342 ( .B1(n102), .B2(n402), .A(n99), .ZN(n97) );
  INV_X1 U343 ( .A(n101), .ZN(n99) );
  OAI21_X1 U344 ( .B1(n144), .B2(n148), .A(n145), .ZN(n143) );
  NOR2_X1 U345 ( .A1(n168), .A2(n371), .ZN(n161) );
  OAI21_X1 U346 ( .B1(n181), .B2(n184), .A(n182), .ZN(n180) );
  NOR2_X1 U347 ( .A1(n137), .A2(n387), .ZN(n130) );
  INV_X1 U348 ( .A(n93), .ZN(n91) );
  AOI21_X1 U349 ( .B1(n172), .B2(n180), .A(n173), .ZN(n171) );
  NOR2_X1 U350 ( .A1(n177), .A2(n386), .ZN(n172) );
  OAI21_X1 U351 ( .B1(n174), .B2(n178), .A(n175), .ZN(n173) );
  NOR2_X1 U352 ( .A1(n128), .A2(n116), .ZN(n114) );
  NAND2_X1 U353 ( .A1(n398), .A2(n399), .ZN(n116) );
  NAND2_X1 U354 ( .A1(n199), .A2(n96), .ZN(n15) );
  INV_X1 U355 ( .A(n95), .ZN(n199) );
  NOR2_X1 U356 ( .A1(n147), .A2(n377), .ZN(n142) );
  AOI21_X1 U357 ( .B1(n143), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U358 ( .B1(n132), .B2(n138), .A(n133), .ZN(n131) );
  INV_X1 U359 ( .A(n126), .ZN(n124) );
  OAI21_X1 U360 ( .B1(n155), .B2(n159), .A(n156), .ZN(n154) );
  AOI21_X1 U361 ( .B1(n399), .B2(n124), .A(n119), .ZN(n117) );
  INV_X1 U362 ( .A(n121), .ZN(n119) );
  NAND2_X1 U363 ( .A1(n187), .A2(n48), .ZN(n3) );
  INV_X1 U364 ( .A(n47), .ZN(n187) );
  NAND2_X1 U365 ( .A1(n191), .A2(n64), .ZN(n7) );
  INV_X1 U366 ( .A(n63), .ZN(n191) );
  NAND2_X1 U367 ( .A1(n193), .A2(n72), .ZN(n9) );
  INV_X1 U368 ( .A(n71), .ZN(n193) );
  NAND2_X1 U369 ( .A1(n195), .A2(n80), .ZN(n11) );
  INV_X1 U370 ( .A(n79), .ZN(n195) );
  NAND2_X1 U371 ( .A1(n408), .A2(n45), .ZN(n2) );
  XNOR2_X1 U372 ( .A(n375), .B(n4), .ZN(SUM[29]) );
  NAND2_X1 U373 ( .A1(n407), .A2(n53), .ZN(n4) );
  XOR2_X1 U374 ( .A(n395), .B(n5), .Z(SUM[28]) );
  NAND2_X1 U375 ( .A1(n189), .A2(n56), .ZN(n5) );
  INV_X1 U376 ( .A(n55), .ZN(n189) );
  NAND2_X1 U377 ( .A1(n405), .A2(n61), .ZN(n6) );
  NAND2_X1 U378 ( .A1(n406), .A2(n69), .ZN(n8) );
  NAND2_X1 U379 ( .A1(n404), .A2(n77), .ZN(n10) );
  NAND2_X1 U380 ( .A1(n403), .A2(n85), .ZN(n12) );
  XOR2_X1 U381 ( .A(n365), .B(n13), .Z(SUM[20]) );
  NAND2_X1 U382 ( .A1(n197), .A2(n88), .ZN(n13) );
  INV_X1 U383 ( .A(n87), .ZN(n197) );
  XNOR2_X1 U384 ( .A(n359), .B(n14), .ZN(SUM[19]) );
  NAND2_X1 U385 ( .A1(n400), .A2(n93), .ZN(n14) );
  NAND2_X1 U386 ( .A1(n402), .A2(n101), .ZN(n16) );
  XOR2_X1 U387 ( .A(n122), .B(n20), .Z(SUM[13]) );
  NAND2_X1 U388 ( .A1(n399), .A2(n121), .ZN(n20) );
  AOI21_X1 U389 ( .B1(n127), .B2(n398), .A(n124), .ZN(n122) );
  XOR2_X1 U390 ( .A(n134), .B(n22), .Z(SUM[11]) );
  NAND2_X1 U391 ( .A1(n345), .A2(n133), .ZN(n22) );
  AOI21_X1 U392 ( .B1(n139), .B2(n207), .A(n136), .ZN(n134) );
  NAND2_X1 U393 ( .A1(n201), .A2(n104), .ZN(n17) );
  INV_X1 U394 ( .A(n103), .ZN(n201) );
  INV_X1 U395 ( .A(n137), .ZN(n207) );
  INV_X1 U396 ( .A(n168), .ZN(n213) );
  XOR2_X1 U397 ( .A(n160), .B(n27), .Z(SUM[6]) );
  NAND2_X1 U398 ( .A1(n211), .A2(n159), .ZN(n27) );
  INV_X1 U399 ( .A(n158), .ZN(n211) );
  INV_X1 U400 ( .A(n138), .ZN(n136) );
  INV_X1 U401 ( .A(n169), .ZN(n167) );
  INV_X1 U402 ( .A(n377), .ZN(n208) );
  INV_X1 U403 ( .A(n362), .ZN(n210) );
  INV_X1 U404 ( .A(n371), .ZN(n212) );
  INV_X1 U405 ( .A(n386), .ZN(n214) );
  XOR2_X1 U406 ( .A(n165), .B(n28), .Z(SUM[5]) );
  NAND2_X1 U407 ( .A1(n212), .A2(n164), .ZN(n28) );
  AOI21_X1 U408 ( .B1(n170), .B2(n213), .A(n167), .ZN(n165) );
  XNOR2_X1 U409 ( .A(n170), .B(n29), .ZN(SUM[4]) );
  NAND2_X1 U410 ( .A1(n213), .A2(n169), .ZN(n29) );
  XNOR2_X1 U411 ( .A(n176), .B(n30), .ZN(SUM[3]) );
  NAND2_X1 U412 ( .A1(n214), .A2(n175), .ZN(n30) );
  OAI21_X1 U413 ( .B1(n179), .B2(n177), .A(n178), .ZN(n176) );
  XOR2_X1 U414 ( .A(n179), .B(n31), .Z(SUM[2]) );
  NAND2_X1 U415 ( .A1(n215), .A2(n178), .ZN(n31) );
  INV_X1 U416 ( .A(n177), .ZN(n215) );
  XOR2_X1 U417 ( .A(n32), .B(n184), .Z(SUM[1]) );
  NAND2_X1 U418 ( .A1(n216), .A2(n182), .ZN(n32) );
  INV_X1 U419 ( .A(n181), .ZN(n216) );
  AND2_X1 U420 ( .A1(n346), .A2(n184), .ZN(SUM[0]) );
  NAND2_X1 U421 ( .A1(n203), .A2(n112), .ZN(n19) );
  INV_X1 U422 ( .A(n111), .ZN(n203) );
  NAND2_X1 U423 ( .A1(n401), .A2(n109), .ZN(n18) );
  XNOR2_X1 U424 ( .A(n127), .B(n21), .ZN(SUM[12]) );
  NAND2_X1 U425 ( .A1(n398), .A2(n126), .ZN(n21) );
  XNOR2_X1 U426 ( .A(n139), .B(n23), .ZN(SUM[10]) );
  NAND2_X1 U427 ( .A1(n207), .A2(n138), .ZN(n23) );
  XNOR2_X1 U428 ( .A(n146), .B(n24), .ZN(SUM[9]) );
  NAND2_X1 U429 ( .A1(n208), .A2(n145), .ZN(n24) );
  OAI21_X1 U430 ( .B1(n149), .B2(n147), .A(n148), .ZN(n146) );
  XOR2_X1 U431 ( .A(n149), .B(n25), .Z(SUM[8]) );
  NAND2_X1 U432 ( .A1(n209), .A2(n148), .ZN(n25) );
  INV_X1 U433 ( .A(n147), .ZN(n209) );
  XNOR2_X1 U434 ( .A(n157), .B(n26), .ZN(SUM[7]) );
  NAND2_X1 U435 ( .A1(n210), .A2(n156), .ZN(n26) );
  OAI21_X1 U436 ( .B1(n160), .B2(n158), .A(n159), .ZN(n157) );
  NOR2_X1 U437 ( .A1(B[8]), .A2(A[8]), .ZN(n147) );
  NOR2_X1 U438 ( .A1(B[6]), .A2(A[6]), .ZN(n158) );
  NOR2_X1 U439 ( .A1(B[2]), .A2(A[2]), .ZN(n177) );
  NOR2_X1 U440 ( .A1(B[5]), .A2(A[5]), .ZN(n163) );
  OR2_X1 U441 ( .A1(B[12]), .A2(A[12]), .ZN(n398) );
  OR2_X1 U442 ( .A1(B[13]), .A2(A[13]), .ZN(n399) );
  NAND2_X1 U443 ( .A1(B[11]), .A2(A[11]), .ZN(n133) );
  NOR2_X1 U444 ( .A1(B[10]), .A2(A[10]), .ZN(n137) );
  NOR2_X1 U445 ( .A1(B[4]), .A2(A[4]), .ZN(n168) );
  NOR2_X1 U446 ( .A1(B[1]), .A2(A[1]), .ZN(n181) );
  NAND2_X1 U447 ( .A1(B[8]), .A2(A[8]), .ZN(n148) );
  NAND2_X1 U448 ( .A1(B[6]), .A2(A[6]), .ZN(n159) );
  OR2_X1 U449 ( .A1(B[19]), .A2(A[19]), .ZN(n400) );
  NAND2_X1 U450 ( .A1(B[0]), .A2(A[0]), .ZN(n184) );
  NAND2_X1 U451 ( .A1(B[10]), .A2(A[10]), .ZN(n138) );
  NAND2_X1 U452 ( .A1(B[4]), .A2(A[4]), .ZN(n169) );
  NAND2_X1 U453 ( .A1(B[9]), .A2(A[9]), .ZN(n145) );
  NAND2_X1 U454 ( .A1(B[3]), .A2(A[3]), .ZN(n175) );
  NAND2_X1 U455 ( .A1(B[1]), .A2(A[1]), .ZN(n182) );
  NAND2_X1 U456 ( .A1(B[5]), .A2(A[5]), .ZN(n164) );
  NAND2_X1 U457 ( .A1(B[7]), .A2(A[7]), .ZN(n156) );
  INV_X1 U458 ( .A(n45), .ZN(n43) );
  NOR2_X1 U459 ( .A1(B[20]), .A2(A[20]), .ZN(n87) );
  NOR2_X1 U460 ( .A1(B[18]), .A2(A[18]), .ZN(n95) );
  NOR2_X1 U461 ( .A1(B[14]), .A2(A[14]), .ZN(n111) );
  NOR2_X1 U462 ( .A1(B[16]), .A2(A[16]), .ZN(n103) );
  NOR2_X1 U463 ( .A1(B[30]), .A2(A[30]), .ZN(n47) );
  NOR2_X1 U464 ( .A1(B[28]), .A2(A[28]), .ZN(n55) );
  NOR2_X1 U465 ( .A1(B[26]), .A2(A[26]), .ZN(n63) );
  NOR2_X1 U466 ( .A1(B[24]), .A2(A[24]), .ZN(n71) );
  NOR2_X1 U467 ( .A1(B[22]), .A2(A[22]), .ZN(n79) );
  OR2_X1 U468 ( .A1(B[15]), .A2(A[15]), .ZN(n401) );
  OR2_X1 U469 ( .A1(B[17]), .A2(A[17]), .ZN(n402) );
  NAND2_X1 U470 ( .A1(B[21]), .A2(A[21]), .ZN(n85) );
  NAND2_X1 U471 ( .A1(B[12]), .A2(A[12]), .ZN(n126) );
  NAND2_X1 U472 ( .A1(B[19]), .A2(A[19]), .ZN(n93) );
  NAND2_X1 U473 ( .A1(B[13]), .A2(A[13]), .ZN(n121) );
  NAND2_X1 U474 ( .A1(B[15]), .A2(A[15]), .ZN(n109) );
  NAND2_X1 U475 ( .A1(B[17]), .A2(A[17]), .ZN(n101) );
  NAND2_X1 U476 ( .A1(B[23]), .A2(A[23]), .ZN(n77) );
  NAND2_X1 U477 ( .A1(B[25]), .A2(A[25]), .ZN(n69) );
  NAND2_X1 U478 ( .A1(B[27]), .A2(A[27]), .ZN(n61) );
  NAND2_X1 U479 ( .A1(B[29]), .A2(A[29]), .ZN(n53) );
  NAND2_X1 U480 ( .A1(B[31]), .A2(A[31]), .ZN(n45) );
  NAND2_X1 U481 ( .A1(B[20]), .A2(A[20]), .ZN(n88) );
  NAND2_X1 U482 ( .A1(B[18]), .A2(A[18]), .ZN(n96) );
  NAND2_X1 U483 ( .A1(B[14]), .A2(A[14]), .ZN(n112) );
  NAND2_X1 U484 ( .A1(B[16]), .A2(A[16]), .ZN(n104) );
  NAND2_X1 U485 ( .A1(B[30]), .A2(A[30]), .ZN(n48) );
  NAND2_X1 U486 ( .A1(B[28]), .A2(A[28]), .ZN(n56) );
  NAND2_X1 U487 ( .A1(B[26]), .A2(A[26]), .ZN(n64) );
  NAND2_X1 U488 ( .A1(B[24]), .A2(A[24]), .ZN(n72) );
  NAND2_X1 U489 ( .A1(B[22]), .A2(A[22]), .ZN(n80) );
  OR2_X1 U490 ( .A1(B[21]), .A2(A[21]), .ZN(n403) );
  OR2_X1 U491 ( .A1(B[23]), .A2(A[23]), .ZN(n404) );
  OR2_X1 U492 ( .A1(B[27]), .A2(A[27]), .ZN(n405) );
  OR2_X1 U493 ( .A1(B[25]), .A2(A[25]), .ZN(n406) );
  OR2_X1 U494 ( .A1(B[29]), .A2(A[29]), .ZN(n407) );
  OR2_X1 U495 ( .A1(B[31]), .A2(A[31]), .ZN(n408) );
  XNOR2_X1 U496 ( .A(n34), .B(n409), .ZN(SUM[39]) );
  XNOR2_X1 U497 ( .A(A[39]), .B(B[39]), .ZN(n409) );
  OAI21_X1 U498 ( .B1(n97), .B2(n95), .A(n96), .ZN(n94) );
  XOR2_X1 U499 ( .A(n393), .B(n15), .Z(SUM[18]) );
  XNOR2_X1 U500 ( .A(n360), .B(n8), .ZN(SUM[25]) );
  XNOR2_X1 U501 ( .A(n376), .B(n16), .ZN(SUM[17]) );
  XNOR2_X1 U502 ( .A(n370), .B(n6), .ZN(SUM[27]) );
  OAI21_X1 U503 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  AOI21_X1 U504 ( .B1(n54), .B2(n407), .A(n51), .ZN(n49) );
  XOR2_X1 U505 ( .A(n390), .B(n3), .Z(SUM[30]) );
  XOR2_X1 U506 ( .A(n388), .B(n17), .Z(SUM[16]) );
  OAI21_X1 U507 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  OAI21_X1 U508 ( .B1(n105), .B2(n103), .A(n104), .ZN(n102) );
  XNOR2_X1 U509 ( .A(n389), .B(n2), .ZN(SUM[31]) );
  XNOR2_X1 U510 ( .A(n392), .B(n10), .ZN(SUM[23]) );
  XNOR2_X1 U511 ( .A(n372), .B(n18), .ZN(SUM[15]) );
  INV_X1 U512 ( .A(n41), .ZN(n185) );
  AOI21_X1 U513 ( .B1(n46), .B2(n408), .A(n43), .ZN(n41) );
  AOI21_X1 U514 ( .B1(n78), .B2(n404), .A(n75), .ZN(n73) );
  XNOR2_X1 U515 ( .A(n391), .B(n12), .ZN(SUM[21]) );
  XOR2_X1 U516 ( .A(n368), .B(n19), .Z(SUM[14]) );
  XOR2_X1 U517 ( .A(n396), .B(n11), .Z(SUM[22]) );
  INV_X1 U518 ( .A(n150), .ZN(n149) );
  OAI21_X1 U519 ( .B1(n81), .B2(n79), .A(n80), .ZN(n78) );
  AOI21_X1 U520 ( .B1(n86), .B2(n403), .A(n83), .ZN(n81) );
  OAI21_X1 U521 ( .B1(n113), .B2(n111), .A(n112), .ZN(n110) );
  OAI21_X1 U522 ( .B1(n171), .B2(n151), .A(n152), .ZN(n150) );
  OAI21_X1 U523 ( .B1(n89), .B2(n87), .A(n88), .ZN(n86) );
  XOR2_X1 U524 ( .A(n366), .B(n7), .Z(SUM[26]) );
  XOR2_X1 U525 ( .A(n394), .B(n9), .Z(SUM[24]) );
  OAI21_X1 U526 ( .B1(n149), .B2(n128), .A(n369), .ZN(n127) );
  OAI21_X1 U527 ( .B1(n65), .B2(n63), .A(n64), .ZN(n62) );
  OAI21_X1 U528 ( .B1(n73), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U529 ( .B1(n129), .B2(n116), .A(n117), .ZN(n115) );
endmodule


module mac_6 ( clk, clear_acc, a, b, mac_out );
  input [19:0] a;
  input [19:0] b;
  output [39:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, n2, n3;
  wire   [39:0] mul;
  wire   [39:0] pipeline;
  wire   [39:0] sum;

  DFF_X1 \pipeline_reg[38]  ( .D(mul[38]), .CK(clk), .Q(pipeline[38]) );
  DFF_X1 \pipeline_reg[37]  ( .D(mul[37]), .CK(clk), .Q(pipeline[37]) );
  DFF_X1 \pipeline_reg[36]  ( .D(mul[36]), .CK(clk), .Q(pipeline[36]) );
  DFF_X1 \pipeline_reg[35]  ( .D(mul[35]), .CK(clk), .Q(pipeline[35]) );
  DFF_X1 \pipeline_reg[34]  ( .D(mul[34]), .CK(clk), .Q(pipeline[34]) );
  DFF_X1 \pipeline_reg[33]  ( .D(mul[33]), .CK(clk), .Q(pipeline[33]) );
  DFF_X1 \pipeline_reg[32]  ( .D(mul[32]), .CK(clk), .Q(pipeline[32]) );
  DFF_X1 \pipeline_reg[31]  ( .D(mul[31]), .CK(clk), .Q(pipeline[31]) );
  DFF_X1 \pipeline_reg[30]  ( .D(mul[30]), .CK(clk), .Q(pipeline[30]) );
  DFF_X1 \pipeline_reg[29]  ( .D(mul[29]), .CK(clk), .Q(pipeline[29]) );
  DFF_X1 \pipeline_reg[28]  ( .D(mul[28]), .CK(clk), .Q(pipeline[28]) );
  DFF_X1 \pipeline_reg[27]  ( .D(mul[27]), .CK(clk), .Q(pipeline[27]) );
  DFF_X1 \pipeline_reg[26]  ( .D(mul[26]), .CK(clk), .Q(pipeline[26]) );
  DFF_X1 \pipeline_reg[25]  ( .D(mul[25]), .CK(clk), .Q(pipeline[25]) );
  DFF_X1 \pipeline_reg[24]  ( .D(mul[24]), .CK(clk), .Q(pipeline[24]) );
  DFF_X1 \pipeline_reg[23]  ( .D(mul[23]), .CK(clk), .Q(pipeline[23]) );
  DFF_X1 \pipeline_reg[22]  ( .D(mul[22]), .CK(clk), .Q(pipeline[22]) );
  DFF_X1 \pipeline_reg[21]  ( .D(mul[21]), .CK(clk), .Q(pipeline[21]) );
  DFF_X1 \pipeline_reg[20]  ( .D(mul[20]), .CK(clk), .Q(pipeline[20]) );
  DFF_X1 \pipeline_reg[19]  ( .D(mul[19]), .CK(clk), .Q(pipeline[19]) );
  DFF_X1 \pipeline_reg[18]  ( .D(mul[18]), .CK(clk), .Q(pipeline[18]) );
  DFF_X1 \pipeline_reg[17]  ( .D(mul[17]), .CK(clk), .Q(pipeline[17]) );
  DFF_X1 \pipeline_reg[16]  ( .D(mul[16]), .CK(clk), .Q(pipeline[16]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \mac_out_reg[16]  ( .D(N19), .CK(clk), .Q(mac_out[16]) );
  DFF_X1 \mac_out_reg[17]  ( .D(N20), .CK(clk), .Q(mac_out[17]) );
  DFF_X1 \mac_out_reg[18]  ( .D(N21), .CK(clk), .Q(mac_out[18]) );
  DFF_X1 \mac_out_reg[19]  ( .D(N22), .CK(clk), .Q(mac_out[19]) );
  DFF_X1 \mac_out_reg[20]  ( .D(N23), .CK(clk), .Q(mac_out[20]) );
  DFF_X1 \mac_out_reg[21]  ( .D(N24), .CK(clk), .Q(mac_out[21]) );
  DFF_X1 \mac_out_reg[22]  ( .D(N25), .CK(clk), .Q(mac_out[22]) );
  DFF_X1 \mac_out_reg[23]  ( .D(N26), .CK(clk), .Q(mac_out[23]) );
  DFF_X1 \mac_out_reg[24]  ( .D(N27), .CK(clk), .Q(mac_out[24]) );
  DFF_X1 \mac_out_reg[25]  ( .D(N28), .CK(clk), .Q(mac_out[25]) );
  DFF_X1 \mac_out_reg[26]  ( .D(N29), .CK(clk), .Q(mac_out[26]) );
  DFF_X1 \mac_out_reg[27]  ( .D(N30), .CK(clk), .Q(mac_out[27]) );
  DFF_X1 \mac_out_reg[28]  ( .D(N31), .CK(clk), .Q(mac_out[28]) );
  DFF_X1 \mac_out_reg[29]  ( .D(N32), .CK(clk), .Q(mac_out[29]) );
  DFF_X1 \mac_out_reg[30]  ( .D(N33), .CK(clk), .Q(mac_out[30]) );
  DFF_X1 \mac_out_reg[31]  ( .D(N34), .CK(clk), .Q(mac_out[31]) );
  DFF_X1 \mac_out_reg[32]  ( .D(N35), .CK(clk), .Q(mac_out[32]) );
  DFF_X1 \mac_out_reg[33]  ( .D(N36), .CK(clk), .Q(mac_out[33]) );
  DFF_X1 \mac_out_reg[34]  ( .D(N37), .CK(clk), .Q(mac_out[34]) );
  DFF_X1 \mac_out_reg[35]  ( .D(N38), .CK(clk), .Q(mac_out[35]) );
  DFF_X1 \mac_out_reg[36]  ( .D(N39), .CK(clk), .Q(mac_out[36]) );
  DFF_X1 \mac_out_reg[37]  ( .D(N40), .CK(clk), .Q(mac_out[37]) );
  DFF_X1 \mac_out_reg[38]  ( .D(N41), .CK(clk), .Q(mac_out[38]) );
  DFF_X1 \mac_out_reg[39]  ( .D(N42), .CK(clk), .Q(mac_out[39]) );
  mac_6_DW_mult_tc_1 mult_355 ( .a(a), .b(b), .product(mul) );
  mac_6_DW01_add_1 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  DFF_X2 \pipeline_reg[39]  ( .D(mul[39]), .CK(clk), .Q(pipeline[39]) );
  BUF_X1 U3 ( .A(n3), .Z(n2) );
  INV_X1 U4 ( .A(clear_acc), .ZN(n3) );
  AND2_X1 U6 ( .A1(sum[39]), .A2(n2), .ZN(N42) );
  AND2_X1 U7 ( .A1(sum[38]), .A2(n2), .ZN(N41) );
  AND2_X1 U8 ( .A1(sum[37]), .A2(n2), .ZN(N40) );
  AND2_X1 U9 ( .A1(sum[36]), .A2(n2), .ZN(N39) );
  AND2_X1 U10 ( .A1(sum[35]), .A2(n2), .ZN(N38) );
  AND2_X1 U11 ( .A1(sum[34]), .A2(n2), .ZN(N37) );
  AND2_X1 U12 ( .A1(sum[33]), .A2(n2), .ZN(N36) );
  AND2_X1 U13 ( .A1(sum[32]), .A2(n2), .ZN(N35) );
  AND2_X1 U14 ( .A1(sum[31]), .A2(n2), .ZN(N34) );
  AND2_X1 U15 ( .A1(sum[30]), .A2(n2), .ZN(N33) );
  AND2_X1 U16 ( .A1(sum[29]), .A2(n2), .ZN(N32) );
  AND2_X1 U17 ( .A1(sum[28]), .A2(n3), .ZN(N31) );
  AND2_X1 U18 ( .A1(sum[27]), .A2(n3), .ZN(N30) );
  AND2_X1 U19 ( .A1(sum[26]), .A2(n3), .ZN(N29) );
  AND2_X1 U20 ( .A1(sum[25]), .A2(n3), .ZN(N28) );
  AND2_X1 U21 ( .A1(sum[24]), .A2(n3), .ZN(N27) );
  AND2_X1 U22 ( .A1(sum[23]), .A2(n3), .ZN(N26) );
  AND2_X1 U23 ( .A1(sum[22]), .A2(n3), .ZN(N25) );
  AND2_X1 U24 ( .A1(sum[21]), .A2(n3), .ZN(N24) );
  AND2_X1 U25 ( .A1(sum[20]), .A2(n3), .ZN(N23) );
  AND2_X1 U26 ( .A1(sum[19]), .A2(n3), .ZN(N22) );
  AND2_X1 U27 ( .A1(sum[18]), .A2(n3), .ZN(N21) );
  AND2_X1 U28 ( .A1(sum[17]), .A2(n3), .ZN(N20) );
  AND2_X1 U29 ( .A1(sum[16]), .A2(n3), .ZN(N19) );
  AND2_X1 U30 ( .A1(sum[15]), .A2(n3), .ZN(N18) );
  AND2_X1 U31 ( .A1(sum[14]), .A2(n3), .ZN(N17) );
  AND2_X1 U32 ( .A1(sum[13]), .A2(n3), .ZN(N16) );
  AND2_X1 U33 ( .A1(sum[12]), .A2(n3), .ZN(N15) );
  AND2_X1 U34 ( .A1(sum[11]), .A2(n3), .ZN(N14) );
  AND2_X1 U35 ( .A1(sum[10]), .A2(n3), .ZN(N13) );
  AND2_X1 U36 ( .A1(sum[9]), .A2(n3), .ZN(N12) );
  AND2_X1 U37 ( .A1(sum[8]), .A2(n3), .ZN(N11) );
  AND2_X1 U38 ( .A1(sum[7]), .A2(n3), .ZN(N10) );
  AND2_X1 U39 ( .A1(sum[6]), .A2(n3), .ZN(N9) );
  AND2_X1 U40 ( .A1(sum[5]), .A2(n3), .ZN(N8) );
  AND2_X1 U41 ( .A1(sum[4]), .A2(n3), .ZN(N7) );
  AND2_X1 U42 ( .A1(sum[3]), .A2(n3), .ZN(N6) );
  AND2_X1 U43 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U44 ( .A1(sum[1]), .A2(n3), .ZN(N4) );
  AND2_X1 U45 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
endmodule


module mac_5_DW_mult_tc_1 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n4, n6, n7, n9, n12, n13, n16, n19, n24, n25, n28, n31, n34, n36,
         n37, n40, n42, n43, n46, n48, n49, n52, n54, n55, n60, n61, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n97, n98, n99, n100, n101, n103, n105, n106, n107, n108,
         n109, n111, n113, n114, n115, n116, n117, n119, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n185, n186, n188, n193, n194, n195, n196, n198, n200, n201,
         n202, n203, n204, n205, n206, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n227,
         n228, n230, n232, n233, n234, n236, n238, n239, n240, n241, n242,
         n244, n246, n247, n248, n249, n250, n252, n254, n255, n256, n257,
         n258, n259, n260, n261, n263, n264, n266, n268, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n284, n285, n286,
         n287, n291, n293, n295, n296, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n643, n644, n646,
         n647, n649, n650, n652, n653, n655, n656, n658, n659, n661, n662,
         n664, n667, n668, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1115, n1117, n1119, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1233, n1234, n1235, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n37 = a[13];
  assign n43 = a[15];
  assign n49 = a[17];
  assign n55 = a[19];
  assign n61 = b[0];
  assign n668 = a[0];
  assign n1090 = b[19];
  assign n1091 = b[18];
  assign n1092 = b[17];
  assign n1093 = b[16];
  assign n1094 = b[15];
  assign n1095 = b[14];
  assign n1096 = b[13];
  assign n1097 = b[12];
  assign n1098 = b[11];
  assign n1099 = b[10];
  assign n1100 = b[9];
  assign n1101 = b[8];
  assign n1102 = b[7];
  assign n1103 = b[6];
  assign n1104 = b[5];
  assign n1105 = b[4];
  assign n1106 = b[3];
  assign n1107 = b[2];
  assign n1108 = b[1];

  FA_X1 U333 ( .A(n681), .B(n304), .CI(n700), .CO(n300), .S(n301) );
  FA_X1 U334 ( .A(n305), .B(n682), .CI(n308), .CO(n302), .S(n303) );
  FA_X1 U336 ( .A(n312), .B(n683), .CI(n309), .CO(n306), .S(n307) );
  FA_X1 U337 ( .A(n701), .B(n314), .CI(n720), .CO(n308), .S(n309) );
  FA_X1 U338 ( .A(n313), .B(n320), .CI(n318), .CO(n310), .S(n311) );
  FA_X1 U339 ( .A(n684), .B(n702), .CI(n315), .CO(n312), .S(n313) );
  FA_X1 U341 ( .A(n324), .B(n321), .CI(n319), .CO(n316), .S(n317) );
  FA_X1 U342 ( .A(n328), .B(n721), .CI(n326), .CO(n318), .S(n319) );
  FA_X1 U343 ( .A(n703), .B(n685), .CI(n740), .CO(n320), .S(n321) );
  FA_X1 U344 ( .A(n325), .B(n327), .CI(n332), .CO(n322), .S(n323) );
  FA_X1 U345 ( .A(n336), .B(n329), .CI(n334), .CO(n324), .S(n325) );
  FA_X1 U346 ( .A(n686), .B(n704), .CI(n722), .CO(n326), .S(n327) );
  FA_X1 U348 ( .A(n340), .B(n342), .CI(n333), .CO(n330), .S(n331) );
  FA_X1 U349 ( .A(n335), .B(n344), .CI(n337), .CO(n332), .S(n333) );
  FA_X1 U350 ( .A(n705), .B(n346), .CI(n723), .CO(n334), .S(n335) );
  FA_X1 U351 ( .A(n741), .B(n687), .CI(n760), .CO(n336), .S(n337) );
  FA_X1 U352 ( .A(n350), .B(n343), .CI(n341), .CO(n338), .S(n339) );
  FA_X1 U353 ( .A(n345), .B(n354), .CI(n352), .CO(n340), .S(n341) );
  FA_X1 U354 ( .A(n347), .B(n724), .CI(n356), .CO(n342), .S(n343) );
  FA_X1 U355 ( .A(n742), .B(n706), .CI(n688), .CO(n344), .S(n345) );
  FA_X1 U357 ( .A(n360), .B(n353), .CI(n351), .CO(n348), .S(n349) );
  FA_X1 U358 ( .A(n357), .B(n355), .CI(n362), .CO(n350), .S(n351) );
  FA_X1 U359 ( .A(n366), .B(n743), .CI(n364), .CO(n352), .S(n353) );
  FA_X1 U360 ( .A(n707), .B(n761), .CI(n725), .CO(n354), .S(n355) );
  FA_X1 U361 ( .A(n368), .B(n689), .CI(n780), .CO(n356), .S(n357) );
  FA_X1 U362 ( .A(n372), .B(n363), .CI(n361), .CO(n358), .S(n359) );
  FA_X1 U363 ( .A(n376), .B(n365), .CI(n374), .CO(n360), .S(n361) );
  FA_X1 U364 ( .A(n378), .B(n380), .CI(n367), .CO(n362), .S(n363) );
  FA_X1 U365 ( .A(n690), .B(n708), .CI(n369), .CO(n364), .S(n365) );
  FA_X1 U366 ( .A(n762), .B(n726), .CI(n744), .CO(n366), .S(n367) );
  FA_X1 U368 ( .A(n384), .B(n375), .CI(n373), .CO(n370), .S(n371) );
  FA_X1 U369 ( .A(n377), .B(n388), .CI(n386), .CO(n372), .S(n373) );
  FA_X1 U370 ( .A(n379), .B(n390), .CI(n381), .CO(n374), .S(n375) );
  FA_X1 U371 ( .A(n727), .B(n745), .CI(n392), .CO(n376), .S(n377) );
  FA_X1 U372 ( .A(n709), .B(n781), .CI(n763), .CO(n378), .S(n379) );
  FA_X1 U373 ( .A(n394), .B(n691), .CI(n800), .CO(n380), .S(n381) );
  FA_X1 U374 ( .A(n398), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U375 ( .A(n389), .B(n402), .CI(n400), .CO(n384), .S(n385) );
  FA_X1 U376 ( .A(n393), .B(n404), .CI(n391), .CO(n386), .S(n387) );
  FA_X1 U378 ( .A(n764), .B(n782), .CI(n746), .CO(n390), .S(n391) );
  FA_X1 U379 ( .A(n710), .B(n728), .CI(n692), .CO(n392), .S(n393) );
  FA_X1 U381 ( .A(n401), .B(n412), .CI(n399), .CO(n396), .S(n397) );
  FA_X1 U382 ( .A(n403), .B(n416), .CI(n414), .CO(n398), .S(n399) );
  FA_X1 U383 ( .A(n409), .B(n407), .CI(n418), .CO(n400), .S(n401) );
  FA_X1 U384 ( .A(n420), .B(n422), .CI(n405), .CO(n402), .S(n403) );
  FA_X1 U385 ( .A(n729), .B(n747), .CI(n765), .CO(n404), .S(n405) );
  FA_X1 U386 ( .A(n783), .B(n801), .CI(n711), .CO(n406), .S(n407) );
  FA_X1 U387 ( .A(n693), .B(n1362), .CI(n820), .CO(n408), .S(n409) );
  FA_X1 U391 ( .A(n436), .B(n438), .CI(n421), .CO(n416), .S(n417) );
  FA_X1 U392 ( .A(n748), .B(n425), .CI(n440), .CO(n418), .S(n419) );
  FA_X1 U393 ( .A(n694), .B(n766), .CI(n712), .CO(n420), .S(n421) );
  FA_X1 U394 ( .A(n802), .B(n730), .CI(n784), .CO(n422), .S(n423) );
  FA_X1 U398 ( .A(n450), .B(n441), .CI(n435), .CO(n430), .S(n431) );
  FA_X1 U399 ( .A(n437), .B(n452), .CI(n439), .CO(n432), .S(n433) );
  FA_X1 U401 ( .A(n731), .B(n785), .CI(n749), .CO(n436), .S(n437) );
  FA_X1 U402 ( .A(n458), .B(n803), .CI(n713), .CO(n438), .S(n439) );
  FA_X1 U406 ( .A(n468), .B(n453), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U407 ( .A(n455), .B(n470), .CI(n457), .CO(n448), .S(n449) );
  FA_X1 U408 ( .A(n472), .B(n476), .CI(n474), .CO(n450), .S(n451) );
  FA_X1 U409 ( .A(n768), .B(n786), .CI(n459), .CO(n452), .S(n453) );
  FA_X1 U411 ( .A(n696), .B(n822), .CI(n750), .CO(n456), .S(n457) );
  FA_X1 U413 ( .A(n465), .B(n480), .CI(n463), .CO(n460), .S(n461) );
  FA_X1 U414 ( .A(n467), .B(n484), .CI(n482), .CO(n462), .S(n463) );
  FA_X1 U416 ( .A(n473), .B(n488), .CI(n475), .CO(n466), .S(n467) );
  FA_X1 U417 ( .A(n492), .B(n477), .CI(n490), .CO(n468), .S(n469) );
  FA_X1 U418 ( .A(n805), .B(n823), .CI(n494), .CO(n470), .S(n471) );
  FA_X1 U419 ( .A(n841), .B(n733), .CI(n751), .CO(n472), .S(n473) );
  FA_X1 U420 ( .A(n860), .B(n697), .CI(n769), .CO(n474), .S(n475) );
  FA_X1 U423 ( .A(n498), .B(n483), .CI(n481), .CO(n478), .S(n479) );
  FA_X1 U424 ( .A(n485), .B(n487), .CI(n500), .CO(n480), .S(n481) );
  FA_X1 U426 ( .A(n489), .B(n506), .CI(n491), .CO(n484), .S(n485) );
  FA_X1 U427 ( .A(n510), .B(n495), .CI(n508), .CO(n486), .S(n487) );
  FA_X1 U428 ( .A(n770), .B(n842), .CI(n824), .CO(n488), .S(n489) );
  FA_X1 U429 ( .A(n861), .B(n806), .CI(n752), .CO(n490), .S(n491) );
  FA_X1 U430 ( .A(n734), .B(n670), .CI(n788), .CO(n492), .S(n493) );
  HA_X1 U431 ( .A(n698), .B(n716), .CO(n494), .S(n495) );
  FA_X1 U433 ( .A(n516), .B(n505), .CI(n503), .CO(n498), .S(n499) );
  FA_X1 U434 ( .A(n520), .B(n509), .CI(n518), .CO(n500), .S(n501) );
  FA_X1 U438 ( .A(n717), .B(n843), .CI(n753), .CO(n508), .S(n509) );
  FA_X1 U440 ( .A(n517), .B(n530), .CI(n515), .CO(n512), .S(n513) );
  FA_X1 U441 ( .A(n532), .B(n521), .CI(n519), .CO(n514), .S(n515) );
  FA_X1 U442 ( .A(n525), .B(n523), .CI(n534), .CO(n516), .S(n517) );
  FA_X1 U443 ( .A(n536), .B(n540), .CI(n538), .CO(n518), .S(n519) );
  FA_X1 U444 ( .A(n826), .B(n844), .CI(n527), .CO(n520), .S(n521) );
  FA_X1 U445 ( .A(n754), .B(n772), .CI(n808), .CO(n522), .S(n523) );
  FA_X1 U446 ( .A(n790), .B(n863), .CI(n671), .CO(n524), .S(n525) );
  HA_X1 U447 ( .A(n718), .B(n736), .CO(n526), .S(n527) );
  FA_X1 U448 ( .A(n544), .B(n533), .CI(n531), .CO(n528), .S(n529) );
  FA_X1 U449 ( .A(n535), .B(n548), .CI(n546), .CO(n530), .S(n531) );
  FA_X1 U451 ( .A(n552), .B(n554), .CI(n550), .CO(n534), .S(n535) );
  FA_X1 U452 ( .A(n827), .B(n791), .CI(n809), .CO(n536), .S(n537) );
  FA_X1 U453 ( .A(n845), .B(n773), .CI(n737), .CO(n538), .S(n539) );
  FA_X1 U457 ( .A(n562), .B(n564), .CI(n551), .CO(n546), .S(n547) );
  FA_X1 U458 ( .A(n555), .B(n846), .CI(n566), .CO(n548), .S(n549) );
  FA_X1 U459 ( .A(n865), .B(n792), .CI(n828), .CO(n550), .S(n551) );
  FA_X1 U460 ( .A(n774), .B(n672), .CI(n810), .CO(n552), .S(n553) );
  HA_X1 U461 ( .A(n738), .B(n756), .CO(n554), .S(n555) );
  FA_X1 U463 ( .A(n563), .B(n565), .CI(n572), .CO(n558), .S(n559) );
  FA_X1 U464 ( .A(n574), .B(n576), .CI(n567), .CO(n560), .S(n561) );
  FA_X1 U465 ( .A(n811), .B(n829), .CI(n578), .CO(n562), .S(n563) );
  FA_X1 U466 ( .A(n757), .B(n847), .CI(n793), .CO(n564), .S(n565) );
  FA_X1 U467 ( .A(n775), .B(n739), .CI(n866), .CO(n566), .S(n567) );
  FA_X1 U468 ( .A(n582), .B(n573), .CI(n571), .CO(n568), .S(n569) );
  FA_X1 U469 ( .A(n577), .B(n575), .CI(n584), .CO(n570), .S(n571) );
  FA_X1 U470 ( .A(n588), .B(n579), .CI(n586), .CO(n572), .S(n573) );
  FA_X1 U471 ( .A(n794), .B(n848), .CI(n830), .CO(n574), .S(n575) );
  FA_X1 U472 ( .A(n867), .B(n812), .CI(n673), .CO(n576), .S(n577) );
  HA_X1 U473 ( .A(n758), .B(n776), .CO(n578), .S(n579) );
  FA_X1 U474 ( .A(n585), .B(n592), .CI(n583), .CO(n580), .S(n581) );
  FA_X1 U475 ( .A(n587), .B(n589), .CI(n594), .CO(n582), .S(n583) );
  FA_X1 U476 ( .A(n598), .B(n831), .CI(n596), .CO(n584), .S(n585) );
  FA_X1 U477 ( .A(n777), .B(n849), .CI(n813), .CO(n586), .S(n587) );
  FA_X1 U478 ( .A(n795), .B(n759), .CI(n868), .CO(n588), .S(n589) );
  FA_X1 U479 ( .A(n602), .B(n595), .CI(n593), .CO(n590), .S(n591) );
  FA_X1 U480 ( .A(n604), .B(n606), .CI(n597), .CO(n592), .S(n593) );
  FA_X1 U481 ( .A(n814), .B(n850), .CI(n599), .CO(n594), .S(n595) );
  FA_X1 U482 ( .A(n674), .B(n832), .CI(n869), .CO(n596), .S(n597) );
  HA_X1 U483 ( .A(n778), .B(n796), .CO(n598), .S(n599) );
  FA_X1 U484 ( .A(n610), .B(n605), .CI(n603), .CO(n600), .S(n601) );
  FA_X1 U485 ( .A(n612), .B(n614), .CI(n607), .CO(n602), .S(n603) );
  FA_X1 U486 ( .A(n797), .B(n851), .CI(n833), .CO(n604), .S(n605) );
  FA_X1 U487 ( .A(n870), .B(n779), .CI(n815), .CO(n606), .S(n607) );
  FA_X1 U488 ( .A(n613), .B(n618), .CI(n611), .CO(n608), .S(n609) );
  FA_X1 U489 ( .A(n615), .B(n871), .CI(n620), .CO(n610), .S(n611) );
  FA_X1 U490 ( .A(n852), .B(n834), .CI(n675), .CO(n612), .S(n613) );
  HA_X1 U491 ( .A(n798), .B(n816), .CO(n614), .S(n615) );
  FA_X1 U492 ( .A(n621), .B(n624), .CI(n619), .CO(n616), .S(n617) );
  FA_X1 U493 ( .A(n817), .B(n853), .CI(n626), .CO(n618), .S(n619) );
  FA_X1 U494 ( .A(n835), .B(n799), .CI(n872), .CO(n620), .S(n621) );
  FA_X1 U495 ( .A(n630), .B(n627), .CI(n625), .CO(n622), .S(n623) );
  FA_X1 U496 ( .A(n854), .B(n873), .CI(n676), .CO(n624), .S(n625) );
  HA_X1 U497 ( .A(n818), .B(n836), .CO(n626), .S(n627) );
  FA_X1 U498 ( .A(n634), .B(n837), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U499 ( .A(n855), .B(n819), .CI(n874), .CO(n630), .S(n631) );
  FA_X1 U500 ( .A(n677), .B(n856), .CI(n635), .CO(n632), .S(n633) );
  HA_X1 U501 ( .A(n838), .B(n875), .CO(n634), .S(n635) );
  FA_X1 U502 ( .A(n876), .B(n839), .CI(n857), .CO(n636), .S(n637) );
  HA_X1 U503 ( .A(n858), .B(n877), .CO(n638), .S(n639) );
  BUF_X2 U1025 ( .A(n1102), .Z(n1556) );
  AND2_X1 U1026 ( .A1(n1330), .A2(n644), .ZN(n719) );
  BUF_X2 U1027 ( .A(n1450), .Z(n1514) );
  BUF_X2 U1028 ( .A(n52), .Z(n1412) );
  CLKBUF_X1 U1029 ( .A(n755), .Z(n1233) );
  BUF_X1 U1030 ( .A(n28), .Z(n1509) );
  BUF_X4 U1031 ( .A(n43), .Z(n1546) );
  OAI22_X1 U1032 ( .A1(n6), .A2(n1073), .B1(n1072), .B2(n4), .ZN(n1234) );
  BUF_X2 U1033 ( .A(n1093), .Z(n1564) );
  BUF_X2 U1034 ( .A(n1457), .Z(n1308) );
  BUF_X1 U1035 ( .A(n1101), .Z(n1557) );
  BUF_X2 U1036 ( .A(n40), .Z(n1510) );
  BUF_X2 U1037 ( .A(n1097), .Z(n1560) );
  BUF_X2 U1038 ( .A(n1095), .Z(n1562) );
  BUF_X2 U1039 ( .A(n55), .Z(n1548) );
  BUF_X2 U1040 ( .A(n1457), .Z(n1512) );
  BUF_X2 U1041 ( .A(n28), .Z(n1508) );
  BUF_X2 U1042 ( .A(n1092), .Z(n1565) );
  BUF_X1 U1043 ( .A(n49), .Z(n1547) );
  BUF_X1 U1044 ( .A(n1), .Z(n1540) );
  BUF_X2 U1045 ( .A(n16), .Z(n1507) );
  NAND3_X1 U1046 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n504) );
  BUF_X2 U1047 ( .A(n1091), .Z(n1566) );
  BUF_X2 U1048 ( .A(n1540), .Z(n1359) );
  OR2_X1 U1049 ( .A1(n513), .A2(n528), .ZN(n1497) );
  NOR2_X1 U1050 ( .A1(n497), .A2(n512), .ZN(n177) );
  NOR2_X1 U1051 ( .A1(n443), .A2(n460), .ZN(n161) );
  INV_X1 U1052 ( .A(n298), .ZN(n299) );
  INV_X1 U1053 ( .A(n1297), .ZN(n227) );
  BUF_X2 U1054 ( .A(n1107), .Z(n1552) );
  BUF_X1 U1055 ( .A(n1105), .Z(n1306) );
  OR2_X1 U1056 ( .A1(n679), .A2(n879), .ZN(n1235) );
  AND2_X1 U1057 ( .A1(n1235), .A2(n263), .ZN(product[1]) );
  CLKBUF_X1 U1058 ( .A(n840), .Z(n1237) );
  XNOR2_X1 U1059 ( .A(n499), .B(n1238), .ZN(n497) );
  XNOR2_X1 U1060 ( .A(n514), .B(n501), .ZN(n1238) );
  BUF_X2 U1061 ( .A(n25), .Z(n1327) );
  CLKBUF_X1 U1062 ( .A(n212), .Z(n1239) );
  BUF_X1 U1063 ( .A(n1561), .Z(n1336) );
  CLKBUF_X1 U1064 ( .A(n19), .Z(n1240) );
  CLKBUF_X1 U1065 ( .A(n1479), .Z(n1241) );
  BUF_X2 U1066 ( .A(n1479), .Z(n1242) );
  CLKBUF_X3 U1067 ( .A(n37), .Z(n1243) );
  CLKBUF_X1 U1068 ( .A(n37), .Z(n1545) );
  CLKBUF_X1 U1069 ( .A(a[2]), .Z(n1244) );
  CLKBUF_X1 U1070 ( .A(n539), .Z(n1245) );
  CLKBUF_X1 U1071 ( .A(n507), .Z(n1246) );
  INV_X1 U1072 ( .A(n668), .ZN(n1247) );
  INV_X2 U1073 ( .A(n668), .ZN(n4) );
  OR2_X1 U1074 ( .A1(n1462), .A2(n1360), .ZN(n1279) );
  OR2_X1 U1075 ( .A1(n1462), .A2(n1360), .ZN(n1463) );
  NOR2_X1 U1076 ( .A1(n371), .A2(n382), .ZN(n1248) );
  NOR2_X1 U1077 ( .A1(n371), .A2(n382), .ZN(n135) );
  XOR2_X1 U1078 ( .A(n804), .B(n732), .Z(n1249) );
  XOR2_X1 U1079 ( .A(n1249), .B(n714), .Z(n455) );
  NAND2_X1 U1080 ( .A1(n714), .A2(n804), .ZN(n1250) );
  NAND2_X1 U1081 ( .A1(n714), .A2(n732), .ZN(n1251) );
  NAND2_X1 U1082 ( .A1(n804), .A2(n732), .ZN(n1252) );
  NAND3_X1 U1083 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n454) );
  OR2_X2 U1084 ( .A1(n1504), .A2(n1505), .ZN(n755) );
  NAND2_X1 U1085 ( .A1(n1115), .A2(n28), .ZN(n1479) );
  CLKBUF_X1 U1086 ( .A(n48), .Z(n1253) );
  BUF_X1 U1087 ( .A(n1090), .Z(n1567) );
  BUF_X1 U1088 ( .A(n25), .Z(n1544) );
  CLKBUF_X1 U1089 ( .A(n1543), .Z(n1254) );
  XOR2_X1 U1090 ( .A(n526), .B(n807), .Z(n1255) );
  XOR2_X1 U1091 ( .A(n1255), .B(n524), .Z(n505) );
  NAND2_X1 U1092 ( .A1(n526), .A2(n807), .ZN(n1256) );
  NAND2_X1 U1093 ( .A1(n526), .A2(n524), .ZN(n1257) );
  NAND2_X1 U1094 ( .A1(n807), .A2(n524), .ZN(n1258) );
  XOR2_X1 U1095 ( .A(n493), .B(n502), .Z(n1259) );
  XOR2_X1 U1096 ( .A(n1259), .B(n504), .Z(n483) );
  NAND2_X1 U1097 ( .A1(n493), .A2(n502), .ZN(n1260) );
  NAND2_X1 U1098 ( .A1(n493), .A2(n504), .ZN(n1261) );
  NAND2_X1 U1099 ( .A1(n502), .A2(n504), .ZN(n1262) );
  NAND3_X1 U1100 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n482) );
  BUF_X2 U1101 ( .A(n54), .Z(n1320) );
  CLKBUF_X1 U1102 ( .A(n789), .Z(n1340) );
  CLKBUF_X1 U1103 ( .A(n148), .Z(n1263) );
  XNOR2_X1 U1104 ( .A(n1552), .B(n1548), .ZN(n1264) );
  XNOR2_X1 U1105 ( .A(n559), .B(n1265), .ZN(n557) );
  XNOR2_X1 U1106 ( .A(n570), .B(n561), .ZN(n1265) );
  NOR2_X1 U1107 ( .A1(n397), .A2(n410), .ZN(n1266) );
  XNOR2_X1 U1108 ( .A(n1556), .B(n1546), .ZN(n1267) );
  BUF_X2 U1109 ( .A(n1105), .Z(n1305) );
  NAND3_X1 U1110 ( .A1(n1379), .A2(n1380), .A3(n1381), .ZN(n1268) );
  CLKBUF_X3 U1111 ( .A(n31), .Z(n1455) );
  CLKBUF_X2 U1112 ( .A(n31), .Z(n1454) );
  NAND2_X1 U1113 ( .A1(n559), .A2(n570), .ZN(n1269) );
  NAND2_X1 U1114 ( .A1(n559), .A2(n561), .ZN(n1270) );
  NAND2_X1 U1115 ( .A1(n570), .A2(n561), .ZN(n1271) );
  NAND3_X1 U1116 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n556) );
  XOR2_X1 U1117 ( .A(n1542), .B(a[4]), .Z(n1272) );
  BUF_X2 U1118 ( .A(n13), .Z(n1542) );
  XNOR2_X1 U1119 ( .A(n408), .B(n1273), .ZN(n389) );
  XOR2_X1 U1120 ( .A(n406), .B(n394), .Z(n1273) );
  BUF_X2 U1121 ( .A(n1410), .Z(n1274) );
  INV_X1 U1122 ( .A(n647), .ZN(n1275) );
  BUF_X4 U1123 ( .A(n46), .Z(n1513) );
  BUF_X1 U1124 ( .A(n1557), .Z(n1352) );
  BUF_X2 U1125 ( .A(n1557), .Z(n1353) );
  INV_X1 U1126 ( .A(n1546), .ZN(n1276) );
  INV_X2 U1127 ( .A(n1276), .ZN(n1277) );
  CLKBUF_X1 U1128 ( .A(n194), .Z(n1278) );
  INV_X1 U1129 ( .A(n1366), .ZN(n185) );
  OR2_X2 U1130 ( .A1(n1462), .A2(n1360), .ZN(n1280) );
  OR2_X1 U1131 ( .A1(n1462), .A2(n1360), .ZN(n1464) );
  XNOR2_X1 U1132 ( .A(n1281), .B(n446), .ZN(n429) );
  XNOR2_X1 U1133 ( .A(n433), .B(n448), .ZN(n1281) );
  CLKBUF_X1 U1134 ( .A(n1466), .Z(n1282) );
  AND2_X1 U1135 ( .A1(n513), .A2(n528), .ZN(n1366) );
  NAND2_X1 U1136 ( .A1(n1486), .A2(n34), .ZN(n36) );
  OAI22_X1 U1137 ( .A1(n1481), .A2(n1029), .B1(n1028), .B2(n1507), .ZN(n821)
         );
  BUF_X2 U1138 ( .A(n1484), .Z(n1360) );
  NAND3_X1 U1139 ( .A1(n1375), .A2(n1374), .A3(n1373), .ZN(n1283) );
  BUF_X1 U1140 ( .A(n1106), .Z(n1553) );
  NOR2_X2 U1141 ( .A1(n581), .A2(n590), .ZN(n215) );
  XOR2_X1 U1142 ( .A(n469), .B(n471), .Z(n1284) );
  XOR2_X1 U1143 ( .A(n486), .B(n1284), .Z(n465) );
  NAND2_X1 U1144 ( .A1(n486), .A2(n469), .ZN(n1285) );
  NAND2_X1 U1145 ( .A1(n486), .A2(n471), .ZN(n1286) );
  NAND2_X1 U1146 ( .A1(n469), .A2(n471), .ZN(n1287) );
  NAND3_X1 U1147 ( .A1(n1285), .A2(n1286), .A3(n1287), .ZN(n464) );
  CLKBUF_X1 U1148 ( .A(n444), .Z(n1288) );
  XNOR2_X1 U1149 ( .A(n1306), .B(n1546), .ZN(n1289) );
  BUF_X2 U1150 ( .A(n1108), .Z(n1551) );
  CLKBUF_X2 U1151 ( .A(n1104), .Z(n1554) );
  CLKBUF_X1 U1152 ( .A(n1477), .Z(n1290) );
  CLKBUF_X3 U1153 ( .A(n49), .Z(n1410) );
  INV_X1 U1154 ( .A(n641), .ZN(n1407) );
  XOR2_X1 U1155 ( .A(n1237), .B(n695), .Z(n1291) );
  XOR2_X1 U1156 ( .A(n821), .B(n1291), .Z(n441) );
  NAND2_X1 U1157 ( .A1(n821), .A2(n840), .ZN(n1292) );
  NAND2_X1 U1158 ( .A1(n821), .A2(n695), .ZN(n1293) );
  NAND2_X1 U1159 ( .A1(n840), .A2(n695), .ZN(n1294) );
  NAND3_X1 U1160 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n440) );
  CLKBUF_X1 U1161 ( .A(n172), .Z(n1295) );
  CLKBUF_X1 U1162 ( .A(n1497), .Z(n1296) );
  AND2_X1 U1163 ( .A1(n601), .A2(n608), .ZN(n1297) );
  CLKBUF_X1 U1164 ( .A(n167), .Z(n1298) );
  OR2_X2 U1165 ( .A1(n529), .A2(n542), .ZN(n1299) );
  XOR2_X1 U1166 ( .A(n1567), .B(n1474), .Z(n1069) );
  BUF_X2 U1167 ( .A(n1482), .Z(n1318) );
  INV_X2 U1168 ( .A(n1474), .ZN(n1343) );
  CLKBUF_X1 U1169 ( .A(n1537), .Z(n1300) );
  NAND2_X1 U1170 ( .A1(n1395), .A2(n300), .ZN(n1301) );
  CLKBUF_X1 U1171 ( .A(n1538), .Z(n1302) );
  NAND3_X1 U1172 ( .A1(n1300), .A2(n1302), .A3(n1536), .ZN(n1303) );
  CLKBUF_X1 U1173 ( .A(n1392), .Z(n1304) );
  INV_X2 U1174 ( .A(n1140), .ZN(n1307) );
  BUF_X1 U1175 ( .A(n735), .Z(n1411) );
  INV_X1 U1176 ( .A(n1299), .ZN(n1309) );
  XNOR2_X1 U1177 ( .A(n1353), .B(n1327), .ZN(n1310) );
  CLKBUF_X1 U1178 ( .A(n1534), .Z(n1311) );
  CLKBUF_X1 U1179 ( .A(n1533), .Z(n1312) );
  BUF_X2 U1180 ( .A(n1557), .Z(n1354) );
  XNOR2_X1 U1181 ( .A(n1552), .B(n1454), .ZN(n1313) );
  BUF_X1 U1182 ( .A(n1461), .Z(n1314) );
  NAND2_X2 U1183 ( .A1(n1315), .A2(n1316), .ZN(n60) );
  XNOR2_X1 U1184 ( .A(n1547), .B(a[18]), .ZN(n1315) );
  XOR2_X1 U1185 ( .A(n55), .B(a[18]), .Z(n1316) );
  CLKBUF_X1 U1186 ( .A(n1100), .Z(n1356) );
  XOR2_X1 U1187 ( .A(n1542), .B(a[6]), .Z(n1317) );
  CLKBUF_X1 U1188 ( .A(n1100), .Z(n1357) );
  BUF_X2 U1189 ( .A(n1482), .Z(n1319) );
  NAND2_X1 U1190 ( .A1(n1117), .A2(n16), .ZN(n1482) );
  BUF_X2 U1191 ( .A(n54), .Z(n1401) );
  CLKBUF_X1 U1192 ( .A(n9), .Z(n1321) );
  BUF_X2 U1193 ( .A(n9), .Z(n1322) );
  INV_X1 U1194 ( .A(n1484), .ZN(n9) );
  OAI22_X1 U1195 ( .A1(n6), .A2(n1073), .B1(n1072), .B2(n4), .ZN(n1323) );
  INV_X1 U1196 ( .A(n1282), .ZN(n188) );
  AOI21_X1 U1197 ( .B1(n1502), .B2(n247), .A(n244), .ZN(n1324) );
  BUF_X1 U1198 ( .A(n6), .Z(n1325) );
  BUF_X2 U1199 ( .A(n1094), .Z(n1563) );
  BUF_X2 U1200 ( .A(n1103), .Z(n1555) );
  BUF_X1 U1201 ( .A(n40), .Z(n1358) );
  CLKBUF_X2 U1202 ( .A(n25), .Z(n1326) );
  XNOR2_X1 U1203 ( .A(n1328), .B(n454), .ZN(n435) );
  XNOR2_X1 U1204 ( .A(n456), .B(n767), .ZN(n1328) );
  XNOR2_X1 U1205 ( .A(n1305), .B(n1243), .ZN(n1329) );
  BUF_X2 U1206 ( .A(n61), .Z(n1330) );
  CLKBUF_X1 U1207 ( .A(n1510), .Z(n1331) );
  BUF_X1 U1208 ( .A(n6), .Z(n1332) );
  NAND2_X1 U1209 ( .A1(n1119), .A2(n4), .ZN(n6) );
  XNOR2_X1 U1210 ( .A(n1333), .B(n771), .ZN(n507) );
  XNOR2_X1 U1211 ( .A(n789), .B(n825), .ZN(n1333) );
  CLKBUF_X1 U1212 ( .A(n1562), .Z(n1334) );
  BUF_X1 U1213 ( .A(n1098), .Z(n1335) );
  BUF_X2 U1214 ( .A(n1561), .Z(n1337) );
  CLKBUF_X1 U1215 ( .A(n1561), .Z(n1338) );
  NOR2_X1 U1216 ( .A1(n557), .A2(n568), .ZN(n1339) );
  NAND2_X2 U1217 ( .A1(n1486), .A2(n34), .ZN(n1341) );
  AOI21_X1 U1218 ( .B1(n1459), .B2(n1427), .A(n134), .ZN(n1342) );
  INV_X1 U1219 ( .A(n1474), .ZN(n1344) );
  CLKBUF_X1 U1220 ( .A(n1565), .Z(n1345) );
  BUF_X2 U1221 ( .A(n1108), .Z(n1346) );
  NAND2_X1 U1222 ( .A1(n1119), .A2(n4), .ZN(n1461) );
  BUF_X1 U1223 ( .A(n1099), .Z(n1347) );
  BUF_X1 U1224 ( .A(n1099), .Z(n1348) );
  BUF_X1 U1225 ( .A(n1106), .Z(n1349) );
  BUF_X1 U1226 ( .A(n1106), .Z(n1350) );
  CLKBUF_X3 U1227 ( .A(n1090), .Z(n1351) );
  CLKBUF_X1 U1228 ( .A(n1564), .Z(n1355) );
  BUF_X4 U1229 ( .A(n13), .Z(n1361) );
  OAI22_X1 U1230 ( .A1(n1318), .A2(n1028), .B1(n1027), .B2(n1506), .ZN(n1362)
         );
  BUF_X1 U1231 ( .A(n825), .Z(n1363) );
  XNOR2_X1 U1232 ( .A(n1364), .B(n464), .ZN(n445) );
  XNOR2_X1 U1233 ( .A(n449), .B(n466), .ZN(n1364) );
  XNOR2_X1 U1234 ( .A(n1365), .B(n429), .ZN(n427) );
  XNOR2_X1 U1235 ( .A(n444), .B(n431), .ZN(n1365) );
  XNOR2_X1 U1236 ( .A(n1367), .B(n413), .ZN(n411) );
  XNOR2_X1 U1237 ( .A(n428), .B(n415), .ZN(n1367) );
  BUF_X2 U1238 ( .A(n52), .Z(n1413) );
  OR2_X1 U1239 ( .A1(n1368), .A2(n1369), .ZN(n24) );
  XNOR2_X1 U1240 ( .A(n1240), .B(a[6]), .ZN(n1368) );
  XOR2_X1 U1241 ( .A(n1542), .B(a[6]), .Z(n1369) );
  OR2_X2 U1242 ( .A1(n1368), .A2(n1369), .ZN(n1370) );
  OR2_X2 U1243 ( .A1(n1368), .A2(n1317), .ZN(n1371) );
  CLKBUF_X1 U1244 ( .A(n159), .Z(n1372) );
  NAND2_X1 U1245 ( .A1(n433), .A2(n448), .ZN(n1373) );
  NAND2_X1 U1246 ( .A1(n433), .A2(n446), .ZN(n1374) );
  NAND2_X1 U1247 ( .A1(n448), .A2(n446), .ZN(n1375) );
  NAND3_X1 U1248 ( .A1(n1375), .A2(n1374), .A3(n1373), .ZN(n428) );
  NAND2_X1 U1249 ( .A1(n1288), .A2(n431), .ZN(n1376) );
  NAND2_X1 U1250 ( .A1(n1288), .A2(n429), .ZN(n1377) );
  NAND2_X1 U1251 ( .A1(n431), .A2(n429), .ZN(n1378) );
  NAND3_X1 U1252 ( .A1(n1376), .A2(n1377), .A3(n1378), .ZN(n426) );
  NAND2_X1 U1253 ( .A1(n456), .A2(n767), .ZN(n1379) );
  NAND2_X1 U1254 ( .A1(n456), .A2(n454), .ZN(n1380) );
  NAND2_X1 U1255 ( .A1(n767), .A2(n454), .ZN(n1381) );
  NAND3_X1 U1256 ( .A1(n1379), .A2(n1380), .A3(n1381), .ZN(n434) );
  XOR2_X1 U1257 ( .A(n419), .B(n423), .Z(n1382) );
  XOR2_X1 U1258 ( .A(n1382), .B(n434), .Z(n415) );
  NAND2_X1 U1259 ( .A1(n423), .A2(n419), .ZN(n1383) );
  NAND2_X1 U1260 ( .A1(n423), .A2(n1268), .ZN(n1384) );
  NAND2_X1 U1261 ( .A1(n419), .A2(n434), .ZN(n1385) );
  NAND3_X1 U1262 ( .A1(n1383), .A2(n1384), .A3(n1385), .ZN(n414) );
  CLKBUF_X1 U1263 ( .A(n264), .Z(n1386) );
  XOR2_X1 U1264 ( .A(n1540), .B(n668), .Z(n1119) );
  CLKBUF_X1 U1265 ( .A(n1393), .Z(n1387) );
  CLKBUF_X1 U1266 ( .A(n1507), .Z(n1388) );
  NAND3_X1 U1267 ( .A1(n1393), .A2(n1392), .A3(n1394), .ZN(n1389) );
  NAND3_X1 U1268 ( .A1(n1304), .A2(n1387), .A3(n1394), .ZN(n1390) );
  XOR2_X1 U1269 ( .A(n307), .B(n310), .Z(n1391) );
  XOR2_X1 U1270 ( .A(n1386), .B(n1391), .Z(product[34]) );
  NAND2_X1 U1271 ( .A1(n264), .A2(n307), .ZN(n1392) );
  NAND2_X1 U1272 ( .A1(n264), .A2(n310), .ZN(n1393) );
  NAND2_X1 U1273 ( .A1(n307), .A2(n310), .ZN(n1394) );
  NAND3_X1 U1274 ( .A1(n1392), .A2(n1393), .A3(n1394), .ZN(n100) );
  NAND3_X1 U1275 ( .A1(n1537), .A2(n1538), .A3(n1536), .ZN(n1395) );
  NAND2_X1 U1276 ( .A1(n40), .A2(n1487), .ZN(n1396) );
  NAND2_X1 U1277 ( .A1(n1487), .A2(n1358), .ZN(n1397) );
  NAND2_X1 U1278 ( .A1(n1487), .A2(n1358), .ZN(n42) );
  NAND3_X1 U1279 ( .A1(n1301), .A2(n1440), .A3(n1441), .ZN(n1398) );
  NAND3_X1 U1280 ( .A1(n1440), .A2(n1301), .A3(n1441), .ZN(n1399) );
  CLKBUF_X1 U1281 ( .A(n114), .Z(n1400) );
  NAND2_X1 U1282 ( .A1(n1485), .A2(n52), .ZN(n54) );
  CLKBUF_X3 U1283 ( .A(n1446), .Z(n1402) );
  BUF_X1 U1284 ( .A(n1446), .Z(n1511) );
  NAND2_X1 U1285 ( .A1(n771), .A2(n1363), .ZN(n1403) );
  NAND2_X1 U1286 ( .A1(n771), .A2(n1340), .ZN(n1404) );
  NAND2_X1 U1287 ( .A1(n1363), .A2(n1340), .ZN(n1405) );
  NAND3_X1 U1288 ( .A1(n1403), .A2(n1404), .A3(n1405), .ZN(n506) );
  CLKBUF_X1 U1289 ( .A(n1253), .Z(n1406) );
  OR2_X1 U1290 ( .A1(n60), .A2(n898), .ZN(n1408) );
  OR2_X1 U1291 ( .A1(n897), .A2(n1514), .ZN(n1409) );
  NAND2_X1 U1292 ( .A1(n1408), .A2(n1409), .ZN(n697) );
  NAND2_X1 U1293 ( .A1(n408), .A2(n406), .ZN(n1414) );
  NAND2_X1 U1294 ( .A1(n408), .A2(n395), .ZN(n1415) );
  NAND2_X1 U1295 ( .A1(n406), .A2(n395), .ZN(n1416) );
  NAND3_X1 U1296 ( .A1(n1414), .A2(n1415), .A3(n1416), .ZN(n388) );
  INV_X1 U1297 ( .A(n139), .ZN(n1417) );
  CLKBUF_X1 U1298 ( .A(n165), .Z(n1418) );
  XNOR2_X1 U1299 ( .A(n1419), .B(n445), .ZN(n443) );
  XNOR2_X1 U1300 ( .A(n462), .B(n447), .ZN(n1419) );
  AND2_X1 U1301 ( .A1(n529), .A2(n542), .ZN(n1466) );
  XOR2_X1 U1302 ( .A(n417), .B(n432), .Z(n1420) );
  XOR2_X1 U1303 ( .A(n430), .B(n1420), .Z(n413) );
  NAND2_X1 U1304 ( .A1(n417), .A2(n432), .ZN(n1421) );
  NAND2_X1 U1305 ( .A1(n430), .A2(n417), .ZN(n1422) );
  NAND2_X1 U1306 ( .A1(n430), .A2(n432), .ZN(n1423) );
  NAND3_X1 U1307 ( .A1(n1421), .A2(n1422), .A3(n1423), .ZN(n412) );
  NAND2_X1 U1308 ( .A1(n1283), .A2(n415), .ZN(n1424) );
  NAND2_X1 U1309 ( .A1(n1283), .A2(n413), .ZN(n1425) );
  NAND2_X1 U1310 ( .A1(n415), .A2(n413), .ZN(n1426) );
  NAND3_X1 U1311 ( .A1(n1424), .A2(n1425), .A3(n1426), .ZN(n410) );
  CLKBUF_X1 U1312 ( .A(n133), .Z(n1427) );
  CLKBUF_X1 U1313 ( .A(n176), .Z(n1428) );
  NOR2_X1 U1314 ( .A1(n1266), .A2(n150), .ZN(n1429) );
  AND2_X1 U1315 ( .A1(n1429), .A2(n1430), .ZN(n126) );
  AND2_X1 U1316 ( .A1(n271), .A2(n133), .ZN(n1430) );
  CLKBUF_X1 U1317 ( .A(n1396), .Z(n1431) );
  NAND2_X1 U1318 ( .A1(n449), .A2(n466), .ZN(n1432) );
  NAND2_X1 U1319 ( .A1(n449), .A2(n464), .ZN(n1433) );
  NAND2_X1 U1320 ( .A1(n466), .A2(n464), .ZN(n1434) );
  NAND3_X1 U1321 ( .A1(n1432), .A2(n1433), .A3(n1434), .ZN(n444) );
  NAND2_X1 U1322 ( .A1(n462), .A2(n447), .ZN(n1435) );
  NAND2_X1 U1323 ( .A1(n462), .A2(n445), .ZN(n1436) );
  NAND2_X1 U1324 ( .A1(n447), .A2(n445), .ZN(n1437) );
  NAND3_X1 U1325 ( .A1(n1435), .A2(n1436), .A3(n1437), .ZN(n442) );
  XOR2_X1 U1326 ( .A(n300), .B(n299), .Z(n1438) );
  XOR2_X1 U1327 ( .A(n1303), .B(n1438), .Z(product[37]) );
  NAND2_X1 U1328 ( .A1(n1395), .A2(n300), .ZN(n1439) );
  NAND2_X1 U1329 ( .A1(n98), .A2(n299), .ZN(n1440) );
  NAND2_X1 U1330 ( .A1(n300), .A2(n299), .ZN(n1441) );
  NAND3_X1 U1331 ( .A1(n1440), .A2(n1439), .A3(n1441), .ZN(n97) );
  NAND3_X1 U1332 ( .A1(n1533), .A2(n1534), .A3(n1532), .ZN(n1442) );
  NAND3_X1 U1333 ( .A1(n1312), .A2(n1532), .A3(n1311), .ZN(n1443) );
  AOI21_X1 U1334 ( .B1(n1400), .B2(n1495), .A(n111), .ZN(n1444) );
  CLKBUF_X1 U1335 ( .A(n122), .Z(n1445) );
  XNOR2_X1 U1336 ( .A(n25), .B(a[10]), .ZN(n1446) );
  NAND2_X1 U1337 ( .A1(n499), .A2(n514), .ZN(n1447) );
  NAND2_X1 U1338 ( .A1(n499), .A2(n501), .ZN(n1448) );
  NAND2_X1 U1339 ( .A1(n514), .A2(n501), .ZN(n1449) );
  NAND3_X1 U1340 ( .A1(n1447), .A2(n1448), .A3(n1449), .ZN(n496) );
  XNOR2_X1 U1341 ( .A(n1547), .B(a[18]), .ZN(n1450) );
  CLKBUF_X1 U1342 ( .A(n60), .Z(n1451) );
  CLKBUF_X1 U1343 ( .A(n151), .Z(n1452) );
  CLKBUF_X1 U1344 ( .A(n1331), .Z(n1453) );
  AOI21_X1 U1345 ( .B1(n175), .B2(n1278), .A(n1428), .ZN(n1456) );
  XNOR2_X1 U1346 ( .A(n1542), .B(a[6]), .ZN(n1457) );
  XNOR2_X1 U1347 ( .A(n1458), .B(n862), .ZN(n511) );
  XNOR2_X1 U1348 ( .A(n735), .B(n699), .ZN(n1458) );
  CLKBUF_X1 U1349 ( .A(n146), .Z(n1459) );
  CLKBUF_X1 U1350 ( .A(n106), .Z(n1460) );
  OR2_X1 U1351 ( .A1(n1462), .A2(n1360), .ZN(n12) );
  XNOR2_X1 U1352 ( .A(n7), .B(n1244), .ZN(n1462) );
  XNOR2_X1 U1353 ( .A(n1465), .B(n511), .ZN(n503) );
  XNOR2_X1 U1354 ( .A(n522), .B(n1246), .ZN(n1465) );
  NAND2_X1 U1355 ( .A1(n1411), .A2(n699), .ZN(n1467) );
  NAND2_X1 U1356 ( .A1(n1411), .A2(n862), .ZN(n1468) );
  NAND2_X1 U1357 ( .A1(n699), .A2(n862), .ZN(n1469) );
  NAND3_X1 U1358 ( .A1(n1467), .A2(n1468), .A3(n1469), .ZN(n510) );
  NAND2_X1 U1359 ( .A1(n522), .A2(n507), .ZN(n1470) );
  NAND2_X1 U1360 ( .A1(n522), .A2(n511), .ZN(n1471) );
  NAND2_X1 U1361 ( .A1(n507), .A2(n511), .ZN(n1472) );
  NAND3_X1 U1362 ( .A1(n1470), .A2(n1471), .A3(n1472), .ZN(n502) );
  NOR2_X1 U1363 ( .A1(n478), .A2(n461), .ZN(n1473) );
  NOR2_X1 U1364 ( .A1(n461), .A2(n478), .ZN(n166) );
  INV_X1 U1365 ( .A(n1540), .ZN(n1474) );
  CLKBUF_X1 U1366 ( .A(n127), .Z(n1475) );
  AOI21_X1 U1367 ( .B1(n122), .B2(n1494), .A(n119), .ZN(n1476) );
  NOR2_X1 U1368 ( .A1(n427), .A2(n442), .ZN(n1477) );
  NAND2_X1 U1369 ( .A1(n1115), .A2(n28), .ZN(n1478) );
  CLKBUF_X1 U1370 ( .A(n153), .Z(n1480) );
  NAND2_X1 U1371 ( .A1(n1272), .A2(n16), .ZN(n1481) );
  AOI21_X1 U1372 ( .B1(n153), .B2(n126), .A(n127), .ZN(n1483) );
  XOR2_X1 U1373 ( .A(n1), .B(a[2]), .Z(n1484) );
  NOR2_X1 U1374 ( .A1(n359), .A2(n370), .ZN(n128) );
  OR2_X1 U1375 ( .A1(n339), .A2(n348), .ZN(n1494) );
  XOR2_X1 U1376 ( .A(n1547), .B(a[16]), .Z(n1485) );
  XOR2_X1 U1377 ( .A(n31), .B(a[10]), .Z(n1486) );
  XOR2_X1 U1378 ( .A(n37), .B(a[12]), .Z(n1487) );
  NAND2_X2 U1379 ( .A1(n46), .A2(n1488), .ZN(n48) );
  XOR2_X1 U1380 ( .A(n43), .B(a[14]), .Z(n1488) );
  OAI21_X1 U1381 ( .B1(n152), .B2(n143), .A(n144), .ZN(n142) );
  INV_X1 U1382 ( .A(n1459), .ZN(n144) );
  INV_X1 U1383 ( .A(n145), .ZN(n143) );
  INV_X1 U1384 ( .A(n1480), .ZN(n152) );
  NAND2_X1 U1385 ( .A1(n145), .A2(n1427), .ZN(n131) );
  XNOR2_X1 U1386 ( .A(n179), .B(n78), .ZN(product[18]) );
  NAND2_X1 U1387 ( .A1(n280), .A2(n178), .ZN(n78) );
  INV_X1 U1388 ( .A(n177), .ZN(n280) );
  INV_X1 U1389 ( .A(n171), .ZN(n279) );
  INV_X1 U1390 ( .A(n140), .ZN(n273) );
  XOR2_X1 U1391 ( .A(n168), .B(n76), .Z(product[20]) );
  NAND2_X1 U1392 ( .A1(n278), .A2(n1298), .ZN(n76) );
  AOI21_X1 U1393 ( .B1(n173), .B2(n279), .A(n170), .ZN(n168) );
  XOR2_X1 U1394 ( .A(n137), .B(n70), .Z(product[26]) );
  NAND2_X1 U1395 ( .A1(n272), .A2(n136), .ZN(n70) );
  AOI21_X1 U1396 ( .B1(n142), .B2(n273), .A(n139), .ZN(n137) );
  XOR2_X1 U1397 ( .A(n206), .B(n82), .Z(product[14]) );
  NAND2_X1 U1398 ( .A1(n284), .A2(n205), .ZN(n82) );
  AOI21_X1 U1399 ( .B1(n211), .B2(n285), .A(n208), .ZN(n206) );
  XOR2_X1 U1400 ( .A(n152), .B(n73), .Z(product[23]) );
  INV_X1 U1401 ( .A(n150), .ZN(n275) );
  XOR2_X1 U1402 ( .A(n163), .B(n75), .Z(product[21]) );
  NAND2_X1 U1403 ( .A1(n277), .A2(n162), .ZN(n75) );
  XOR2_X1 U1404 ( .A(n201), .B(n81), .Z(product[15]) );
  INV_X1 U1405 ( .A(n221), .ZN(n220) );
  INV_X1 U1406 ( .A(n234), .ZN(n233) );
  XNOR2_X1 U1407 ( .A(n160), .B(n74), .ZN(product[22]) );
  NAND2_X1 U1408 ( .A1(n276), .A2(n1372), .ZN(n74) );
  XNOR2_X1 U1409 ( .A(n173), .B(n77), .ZN(product[19]) );
  NAND2_X1 U1410 ( .A1(n279), .A2(n1295), .ZN(n77) );
  XNOR2_X1 U1411 ( .A(n130), .B(n69), .ZN(product[27]) );
  NAND2_X1 U1412 ( .A1(n271), .A2(n129), .ZN(n69) );
  INV_X1 U1413 ( .A(n128), .ZN(n271) );
  XNOR2_X1 U1414 ( .A(n149), .B(n72), .ZN(product[24]) );
  NAND2_X1 U1415 ( .A1(n274), .A2(n1263), .ZN(n72) );
  XNOR2_X1 U1416 ( .A(n142), .B(n71), .ZN(product[25]) );
  NAND2_X1 U1417 ( .A1(n273), .A2(n1417), .ZN(n71) );
  INV_X1 U1418 ( .A(n141), .ZN(n139) );
  INV_X1 U1419 ( .A(n1295), .ZN(n170) );
  INV_X1 U1420 ( .A(n121), .ZN(n119) );
  INV_X1 U1421 ( .A(n113), .ZN(n111) );
  NOR2_X1 U1422 ( .A1(n215), .A2(n218), .ZN(n213) );
  OAI21_X1 U1423 ( .B1(n215), .B2(n219), .A(n216), .ZN(n214) );
  AOI21_X1 U1424 ( .B1(n239), .B2(n1493), .A(n236), .ZN(n234) );
  INV_X1 U1425 ( .A(n238), .ZN(n236) );
  NOR2_X1 U1426 ( .A1(n427), .A2(n442), .ZN(n158) );
  NAND2_X1 U1427 ( .A1(n270), .A2(n124), .ZN(n68) );
  INV_X1 U1428 ( .A(n123), .ZN(n270) );
  NAND2_X1 U1429 ( .A1(n268), .A2(n116), .ZN(n66) );
  INV_X1 U1430 ( .A(n115), .ZN(n268) );
  NAND2_X1 U1431 ( .A1(n266), .A2(n108), .ZN(n64) );
  INV_X1 U1432 ( .A(n107), .ZN(n266) );
  INV_X1 U1433 ( .A(n209), .ZN(n285) );
  NAND2_X1 U1434 ( .A1(n443), .A2(n460), .ZN(n162) );
  OR2_X1 U1435 ( .A1(n543), .A2(n556), .ZN(n1489) );
  NAND2_X1 U1436 ( .A1(n1494), .A2(n121), .ZN(n67) );
  NAND2_X1 U1437 ( .A1(n1495), .A2(n113), .ZN(n65) );
  NAND2_X1 U1438 ( .A1(n1496), .A2(n105), .ZN(n63) );
  NOR2_X1 U1439 ( .A1(n411), .A2(n426), .ZN(n150) );
  XOR2_X1 U1440 ( .A(n220), .B(n85), .Z(product[11]) );
  NAND2_X1 U1441 ( .A1(n287), .A2(n219), .ZN(n85) );
  INV_X1 U1442 ( .A(n218), .ZN(n287) );
  XOR2_X1 U1443 ( .A(n228), .B(n86), .Z(product[10]) );
  AOI21_X1 U1444 ( .B1(n233), .B2(n1491), .A(n230), .ZN(n228) );
  XOR2_X1 U1445 ( .A(n193), .B(n80), .Z(product[16]) );
  NAND2_X1 U1446 ( .A1(n1299), .A2(n188), .ZN(n80) );
  NOR2_X1 U1447 ( .A1(n557), .A2(n568), .ZN(n204) );
  NOR2_X1 U1448 ( .A1(n479), .A2(n496), .ZN(n171) );
  XNOR2_X1 U1449 ( .A(n217), .B(n84), .ZN(product[12]) );
  NAND2_X1 U1450 ( .A1(n286), .A2(n216), .ZN(n84) );
  OAI21_X1 U1451 ( .B1(n220), .B2(n218), .A(n219), .ZN(n217) );
  INV_X1 U1452 ( .A(n215), .ZN(n286) );
  NOR2_X1 U1453 ( .A1(n383), .A2(n396), .ZN(n140) );
  XNOR2_X1 U1454 ( .A(n239), .B(n88), .ZN(product[8]) );
  NAND2_X1 U1455 ( .A1(n1493), .A2(n238), .ZN(n88) );
  NAND2_X1 U1456 ( .A1(n479), .A2(n496), .ZN(n172) );
  XNOR2_X1 U1457 ( .A(n211), .B(n83), .ZN(product[13]) );
  NAND2_X1 U1458 ( .A1(n285), .A2(n210), .ZN(n83) );
  XNOR2_X1 U1459 ( .A(n186), .B(n79), .ZN(product[17]) );
  OAI21_X1 U1460 ( .B1(n193), .B2(n1309), .A(n188), .ZN(n186) );
  XNOR2_X1 U1461 ( .A(n233), .B(n87), .ZN(product[9]) );
  NAND2_X1 U1462 ( .A1(n1491), .A2(n232), .ZN(n87) );
  NAND2_X1 U1463 ( .A1(n543), .A2(n556), .ZN(n200) );
  NAND2_X1 U1464 ( .A1(n359), .A2(n370), .ZN(n129) );
  NAND2_X1 U1465 ( .A1(n497), .A2(n512), .ZN(n178) );
  NAND2_X1 U1466 ( .A1(n557), .A2(n568), .ZN(n205) );
  INV_X1 U1467 ( .A(n210), .ZN(n208) );
  XNOR2_X1 U1468 ( .A(n1490), .B(n545), .ZN(n543) );
  XNOR2_X1 U1469 ( .A(n547), .B(n558), .ZN(n1490) );
  INV_X1 U1470 ( .A(n246), .ZN(n244) );
  NOR2_X1 U1471 ( .A1(n591), .A2(n600), .ZN(n218) );
  OAI21_X1 U1472 ( .B1(n256), .B2(n258), .A(n257), .ZN(n255) );
  AOI21_X1 U1473 ( .B1(n1501), .B2(n255), .A(n252), .ZN(n250) );
  INV_X1 U1474 ( .A(n254), .ZN(n252) );
  NAND2_X1 U1475 ( .A1(n581), .A2(n590), .ZN(n216) );
  NAND2_X1 U1476 ( .A1(n291), .A2(n241), .ZN(n89) );
  INV_X1 U1477 ( .A(n240), .ZN(n291) );
  OR2_X1 U1478 ( .A1(n609), .A2(n616), .ZN(n1491) );
  NAND2_X1 U1479 ( .A1(n591), .A2(n600), .ZN(n219) );
  NAND2_X1 U1480 ( .A1(n1502), .A2(n246), .ZN(n90) );
  XOR2_X1 U1481 ( .A(n93), .B(n258), .Z(product[3]) );
  NAND2_X1 U1482 ( .A1(n295), .A2(n257), .ZN(n93) );
  INV_X1 U1483 ( .A(n256), .ZN(n295) );
  XOR2_X1 U1484 ( .A(n91), .B(n250), .Z(product[5]) );
  NAND2_X1 U1485 ( .A1(n293), .A2(n249), .ZN(n91) );
  INV_X1 U1486 ( .A(n248), .ZN(n293) );
  OR2_X1 U1487 ( .A1(n601), .A2(n608), .ZN(n1492) );
  NOR2_X1 U1488 ( .A1(n569), .A2(n580), .ZN(n209) );
  NOR2_X1 U1489 ( .A1(n317), .A2(n322), .ZN(n107) );
  NOR2_X1 U1490 ( .A1(n331), .A2(n338), .ZN(n115) );
  NOR2_X1 U1491 ( .A1(n349), .A2(n358), .ZN(n123) );
  INV_X1 U1492 ( .A(n259), .ZN(n258) );
  OAI21_X1 U1493 ( .B1(n260), .B2(n263), .A(n261), .ZN(n259) );
  NAND2_X1 U1494 ( .A1(n569), .A2(n580), .ZN(n210) );
  OR2_X1 U1495 ( .A1(n617), .A2(n622), .ZN(n1493) );
  XNOR2_X1 U1496 ( .A(n92), .B(n255), .ZN(product[4]) );
  NAND2_X1 U1497 ( .A1(n1501), .A2(n254), .ZN(n92) );
  NAND2_X1 U1498 ( .A1(n339), .A2(n348), .ZN(n121) );
  NAND2_X1 U1499 ( .A1(n323), .A2(n330), .ZN(n113) );
  NAND2_X1 U1500 ( .A1(n617), .A2(n622), .ZN(n238) );
  NAND2_X1 U1501 ( .A1(n311), .A2(n316), .ZN(n105) );
  NAND2_X1 U1502 ( .A1(n609), .A2(n616), .ZN(n232) );
  NAND2_X1 U1503 ( .A1(n317), .A2(n322), .ZN(n108) );
  NAND2_X1 U1504 ( .A1(n331), .A2(n338), .ZN(n116) );
  NAND2_X1 U1505 ( .A1(n349), .A2(n358), .ZN(n124) );
  OR2_X1 U1506 ( .A1(n323), .A2(n330), .ZN(n1495) );
  OR2_X1 U1507 ( .A1(n311), .A2(n316), .ZN(n1496) );
  XOR2_X1 U1508 ( .A(n94), .B(n263), .Z(product[2]) );
  NAND2_X1 U1509 ( .A1(n296), .A2(n261), .ZN(n94) );
  INV_X1 U1510 ( .A(n260), .ZN(n296) );
  XNOR2_X1 U1511 ( .A(n1233), .B(n1498), .ZN(n541) );
  XNOR2_X1 U1512 ( .A(n1323), .B(n719), .ZN(n1498) );
  XNOR2_X1 U1513 ( .A(n1499), .B(n549), .ZN(n545) );
  XNOR2_X1 U1514 ( .A(n560), .B(n553), .ZN(n1499) );
  NOR2_X1 U1515 ( .A1(n639), .A2(n678), .ZN(n256) );
  NAND2_X1 U1516 ( .A1(n639), .A2(n678), .ZN(n257) );
  INV_X1 U1517 ( .A(n105), .ZN(n103) );
  NOR2_X1 U1518 ( .A1(n878), .A2(n859), .ZN(n260) );
  XNOR2_X1 U1519 ( .A(n1399), .B(n1500), .ZN(product[38]) );
  XNOR2_X1 U1520 ( .A(n680), .B(n298), .ZN(n1500) );
  NAND2_X1 U1521 ( .A1(n679), .A2(n879), .ZN(n263) );
  NAND2_X1 U1522 ( .A1(n878), .A2(n859), .ZN(n261) );
  OR2_X1 U1523 ( .A1(n637), .A2(n638), .ZN(n1501) );
  INV_X1 U1524 ( .A(n328), .ZN(n329) );
  INV_X1 U1525 ( .A(n394), .ZN(n395) );
  NOR2_X1 U1526 ( .A1(n633), .A2(n636), .ZN(n248) );
  NOR2_X1 U1527 ( .A1(n623), .A2(n628), .ZN(n240) );
  NAND2_X1 U1528 ( .A1(n629), .A2(n632), .ZN(n246) );
  NAND2_X1 U1529 ( .A1(n633), .A2(n636), .ZN(n249) );
  NAND2_X1 U1530 ( .A1(n623), .A2(n628), .ZN(n241) );
  NAND2_X1 U1531 ( .A1(n637), .A2(n638), .ZN(n254) );
  OR2_X1 U1532 ( .A1(n629), .A2(n632), .ZN(n1502) );
  AND3_X1 U1533 ( .A1(n1516), .A2(n1515), .A3(n1517), .ZN(product[39]) );
  OR2_X1 U1534 ( .A1(n1330), .A2(n1148), .ZN(n1068) );
  OAI22_X1 U1535 ( .A1(n1332), .A2(n1086), .B1(n1085), .B2(n1247), .ZN(n877)
         );
  OAI22_X1 U1536 ( .A1(n1332), .A2(n1088), .B1(n1087), .B2(n4), .ZN(n879) );
  OAI22_X1 U1537 ( .A1(n1332), .A2(n1149), .B1(n1089), .B2(n4), .ZN(n679) );
  OR2_X1 U1538 ( .A1(n1330), .A2(n1149), .ZN(n1089) );
  OAI22_X1 U1539 ( .A1(n1332), .A2(n1087), .B1(n1086), .B2(n1247), .ZN(n878)
         );
  AND2_X1 U1540 ( .A1(n1330), .A2(n656), .ZN(n799) );
  OAI22_X1 U1541 ( .A1(n1314), .A2(n1081), .B1(n1080), .B2(n1247), .ZN(n872)
         );
  OAI22_X1 U1542 ( .A1(n1461), .A2(n1074), .B1(n1073), .B2(n4), .ZN(n865) );
  OAI22_X1 U1543 ( .A1(n1314), .A2(n1076), .B1(n1075), .B2(n1247), .ZN(n867)
         );
  AND2_X1 U1544 ( .A1(n1330), .A2(n659), .ZN(n819) );
  OAI22_X1 U1545 ( .A1(n1325), .A2(n1083), .B1(n1082), .B2(n4), .ZN(n874) );
  OAI22_X1 U1546 ( .A1(n1069), .A2(n6), .B1(n1069), .B2(n4), .ZN(n667) );
  OR2_X1 U1547 ( .A1(n1330), .A2(n1147), .ZN(n1047) );
  AND2_X1 U1548 ( .A1(n1550), .A2(n662), .ZN(n839) );
  OAI22_X1 U1549 ( .A1(n1325), .A2(n1085), .B1(n1084), .B2(n4), .ZN(n876) );
  XNOR2_X1 U1550 ( .A(n1549), .B(n1410), .ZN(n920) );
  OAI22_X1 U1551 ( .A1(n1461), .A2(n1084), .B1(n1083), .B2(n4), .ZN(n875) );
  XNOR2_X1 U1552 ( .A(n1351), .B(n1274), .ZN(n901) );
  INV_X1 U1553 ( .A(n643), .ZN(n700) );
  INV_X1 U1554 ( .A(n304), .ZN(n305) );
  BUF_X2 U1555 ( .A(n16), .Z(n1506) );
  BUF_X1 U1556 ( .A(n1098), .Z(n1559) );
  BUF_X1 U1557 ( .A(n1096), .Z(n1561) );
  BUF_X1 U1558 ( .A(n1099), .Z(n1558) );
  XNOR2_X1 U1559 ( .A(n1334), .B(n1274), .ZN(n906) );
  XNOR2_X1 U1560 ( .A(n1338), .B(n1274), .ZN(n907) );
  XNOR2_X1 U1561 ( .A(n1306), .B(n1410), .ZN(n916) );
  XNOR2_X1 U1562 ( .A(n1553), .B(n1410), .ZN(n917) );
  XNOR2_X1 U1563 ( .A(n1560), .B(n1274), .ZN(n908) );
  XNOR2_X1 U1564 ( .A(n1552), .B(n1410), .ZN(n918) );
  XNOR2_X1 U1565 ( .A(n1554), .B(n1410), .ZN(n915) );
  XNOR2_X1 U1566 ( .A(n1357), .B(n1410), .ZN(n911) );
  XNOR2_X1 U1567 ( .A(n1353), .B(n1410), .ZN(n912) );
  XNOR2_X1 U1568 ( .A(n1556), .B(n1410), .ZN(n913) );
  XNOR2_X1 U1569 ( .A(n1346), .B(n1410), .ZN(n919) );
  XNOR2_X1 U1570 ( .A(n1555), .B(n1274), .ZN(n914) );
  XNOR2_X1 U1571 ( .A(n1348), .B(n1274), .ZN(n910) );
  XNOR2_X1 U1572 ( .A(n1559), .B(n1274), .ZN(n909) );
  XNOR2_X1 U1573 ( .A(n1563), .B(n1274), .ZN(n905) );
  XNOR2_X1 U1574 ( .A(n1566), .B(n1274), .ZN(n902) );
  XNOR2_X1 U1575 ( .A(n1355), .B(n1274), .ZN(n904) );
  XNOR2_X1 U1576 ( .A(n1345), .B(n1274), .ZN(n903) );
  XNOR2_X1 U1577 ( .A(n1335), .B(n1307), .ZN(n888) );
  XNOR2_X1 U1578 ( .A(n1558), .B(n1307), .ZN(n889) );
  XNOR2_X1 U1579 ( .A(n1556), .B(n1548), .ZN(n892) );
  XNOR2_X1 U1580 ( .A(n1555), .B(n1548), .ZN(n893) );
  XNOR2_X1 U1581 ( .A(n1554), .B(n1548), .ZN(n894) );
  XNOR2_X1 U1582 ( .A(n1553), .B(n1548), .ZN(n896) );
  XNOR2_X1 U1583 ( .A(n1105), .B(n1548), .ZN(n895) );
  XNOR2_X1 U1584 ( .A(n1354), .B(n1548), .ZN(n891) );
  XNOR2_X1 U1585 ( .A(n1551), .B(n1548), .ZN(n898) );
  XNOR2_X1 U1586 ( .A(n1552), .B(n1548), .ZN(n897) );
  XNOR2_X1 U1587 ( .A(n1356), .B(n1307), .ZN(n890) );
  XNOR2_X1 U1588 ( .A(n1560), .B(n1307), .ZN(n887) );
  XNOR2_X1 U1589 ( .A(n1337), .B(n1307), .ZN(n886) );
  XNOR2_X1 U1590 ( .A(n1334), .B(n1307), .ZN(n885) );
  XNOR2_X1 U1591 ( .A(n1563), .B(n1307), .ZN(n884) );
  XNOR2_X1 U1592 ( .A(n1355), .B(n1307), .ZN(n883) );
  XNOR2_X1 U1593 ( .A(n1345), .B(n1307), .ZN(n882) );
  XNOR2_X1 U1594 ( .A(n1566), .B(n1307), .ZN(n881) );
  AND2_X1 U1595 ( .A1(n1550), .A2(n1360), .ZN(n859) );
  INV_X1 U1596 ( .A(n314), .ZN(n315) );
  AND2_X1 U1597 ( .A1(n1330), .A2(n641), .ZN(n699) );
  OAI22_X1 U1598 ( .A1(n1325), .A2(n1071), .B1(n1070), .B2(n4), .ZN(n862) );
  OAI22_X1 U1599 ( .A1(n1461), .A2(n1072), .B1(n1071), .B2(n4), .ZN(n863) );
  INV_X1 U1600 ( .A(n649), .ZN(n740) );
  INV_X1 U1601 ( .A(n346), .ZN(n347) );
  AND2_X1 U1602 ( .A1(n1330), .A2(n650), .ZN(n759) );
  OAI22_X1 U1603 ( .A1(n1325), .A2(n1077), .B1(n1076), .B2(n4), .ZN(n868) );
  INV_X1 U1604 ( .A(n667), .ZN(n860) );
  INV_X1 U1605 ( .A(n652), .ZN(n760) );
  INV_X1 U1606 ( .A(n646), .ZN(n720) );
  OAI22_X1 U1607 ( .A1(n1332), .A2(n1080), .B1(n1079), .B2(n1247), .ZN(n871)
         );
  AND2_X1 U1608 ( .A1(n1550), .A2(n647), .ZN(n739) );
  OAI22_X1 U1609 ( .A1(n1332), .A2(n1075), .B1(n1074), .B2(n4), .ZN(n866) );
  AND2_X1 U1610 ( .A1(n1330), .A2(n653), .ZN(n779) );
  OAI22_X1 U1611 ( .A1(n1461), .A2(n1079), .B1(n1078), .B2(n4), .ZN(n870) );
  OAI22_X1 U1612 ( .A1(n1461), .A2(n1078), .B1(n1077), .B2(n4), .ZN(n869) );
  OAI22_X1 U1613 ( .A1(n1314), .A2(n1082), .B1(n1081), .B2(n1247), .ZN(n873)
         );
  INV_X1 U1614 ( .A(n458), .ZN(n459) );
  OAI22_X1 U1615 ( .A1(n1461), .A2(n1070), .B1(n1069), .B2(n4), .ZN(n861) );
  INV_X1 U1616 ( .A(n424), .ZN(n425) );
  INV_X1 U1617 ( .A(n368), .ZN(n369) );
  XNOR2_X1 U1618 ( .A(n1550), .B(n1548), .ZN(n899) );
  INV_X1 U1619 ( .A(n658), .ZN(n800) );
  INV_X1 U1620 ( .A(n661), .ZN(n820) );
  INV_X1 U1621 ( .A(n655), .ZN(n780) );
  INV_X1 U1622 ( .A(n664), .ZN(n840) );
  INV_X1 U1623 ( .A(n1410), .ZN(n1141) );
  INV_X1 U1624 ( .A(n1548), .ZN(n1140) );
  NOR2_X1 U1625 ( .A1(n42), .A2(n959), .ZN(n1504) );
  NOR2_X1 U1626 ( .A1(n958), .A2(n1358), .ZN(n1505) );
  OR2_X1 U1627 ( .A1(n1550), .A2(n1142), .ZN(n942) );
  OR2_X1 U1628 ( .A1(n1330), .A2(n1141), .ZN(n921) );
  OR2_X1 U1629 ( .A1(n1330), .A2(n1145), .ZN(n1005) );
  OR2_X1 U1630 ( .A1(n1330), .A2(n1140), .ZN(n900) );
  OR2_X1 U1631 ( .A1(n1330), .A2(n1143), .ZN(n963) );
  OR2_X1 U1632 ( .A1(n1330), .A2(n1144), .ZN(n984) );
  OR2_X1 U1633 ( .A1(n1330), .A2(n1146), .ZN(n1026) );
  XNOR2_X1 U1634 ( .A(n1351), .B(n1307), .ZN(n880) );
  BUF_X2 U1635 ( .A(n61), .Z(n1550) );
  BUF_X2 U1636 ( .A(n61), .Z(n1549) );
  AND2_X1 U1637 ( .A1(n1550), .A2(n668), .ZN(product[0]) );
  XNOR2_X1 U1638 ( .A(n7), .B(a[4]), .ZN(n16) );
  XNOR2_X1 U1639 ( .A(n43), .B(a[16]), .ZN(n52) );
  XNOR2_X1 U1640 ( .A(n19), .B(a[8]), .ZN(n28) );
  BUF_X4 U1641 ( .A(n7), .Z(n1541) );
  XNOR2_X1 U1642 ( .A(n31), .B(a[12]), .ZN(n40) );
  XNOR2_X1 U1643 ( .A(n25), .B(a[10]), .ZN(n34) );
  XNOR2_X1 U1644 ( .A(n37), .B(a[14]), .ZN(n46) );
  NAND2_X1 U1645 ( .A1(n97), .A2(n680), .ZN(n1515) );
  NAND2_X1 U1646 ( .A1(n1398), .A2(n298), .ZN(n1516) );
  NAND2_X1 U1647 ( .A1(n680), .A2(n298), .ZN(n1517) );
  NAND2_X1 U1648 ( .A1(n560), .A2(n553), .ZN(n1518) );
  NAND2_X1 U1649 ( .A1(n560), .A2(n549), .ZN(n1519) );
  NAND2_X1 U1650 ( .A1(n553), .A2(n549), .ZN(n1520) );
  NAND3_X1 U1651 ( .A1(n1518), .A2(n1519), .A3(n1520), .ZN(n544) );
  NAND2_X1 U1652 ( .A1(n547), .A2(n558), .ZN(n1521) );
  NAND2_X1 U1653 ( .A1(n547), .A2(n545), .ZN(n1522) );
  NAND2_X1 U1654 ( .A1(n558), .A2(n545), .ZN(n1523) );
  NAND3_X1 U1655 ( .A1(n1521), .A2(n1522), .A3(n1523), .ZN(n542) );
  INV_X1 U1656 ( .A(n640), .ZN(n680) );
  INV_X1 U1657 ( .A(n232), .ZN(n230) );
  XOR2_X1 U1658 ( .A(n1245), .B(n541), .Z(n1524) );
  XOR2_X1 U1659 ( .A(n537), .B(n1524), .Z(n533) );
  NAND2_X1 U1660 ( .A1(n537), .A2(n539), .ZN(n1525) );
  NAND2_X1 U1661 ( .A1(n537), .A2(n541), .ZN(n1526) );
  NAND2_X1 U1662 ( .A1(n539), .A2(n541), .ZN(n1527) );
  NAND3_X1 U1663 ( .A1(n1525), .A2(n1526), .A3(n1527), .ZN(n532) );
  INV_X1 U1664 ( .A(n161), .ZN(n277) );
  OAI21_X1 U1665 ( .B1(n163), .B2(n161), .A(n162), .ZN(n160) );
  XNOR2_X1 U1666 ( .A(n787), .B(n715), .ZN(n477) );
  OR2_X1 U1667 ( .A1(n787), .A2(n715), .ZN(n476) );
  NOR2_X1 U1668 ( .A1(n397), .A2(n410), .ZN(n147) );
  NAND2_X1 U1669 ( .A1(n383), .A2(n396), .ZN(n141) );
  XNOR2_X1 U1670 ( .A(n1554), .B(n1541), .ZN(n1062) );
  INV_X1 U1671 ( .A(n1541), .ZN(n1148) );
  XNOR2_X1 U1672 ( .A(n1354), .B(n1541), .ZN(n1059) );
  XNOR2_X1 U1673 ( .A(n1565), .B(n1541), .ZN(n1050) );
  XNOR2_X1 U1674 ( .A(n1563), .B(n1541), .ZN(n1052) );
  XNOR2_X1 U1675 ( .A(n1564), .B(n1541), .ZN(n1051) );
  XNOR2_X1 U1676 ( .A(n1566), .B(n1541), .ZN(n1049) );
  XNOR2_X1 U1677 ( .A(n1555), .B(n1541), .ZN(n1061) );
  XNOR2_X1 U1678 ( .A(n1556), .B(n1541), .ZN(n1060) );
  XNOR2_X1 U1679 ( .A(n1559), .B(n1541), .ZN(n1056) );
  XNOR2_X1 U1680 ( .A(n1560), .B(n1541), .ZN(n1055) );
  XNOR2_X1 U1681 ( .A(n1357), .B(n1541), .ZN(n1058) );
  XNOR2_X1 U1682 ( .A(n1550), .B(n1541), .ZN(n1067) );
  XNOR2_X1 U1683 ( .A(n1558), .B(n1541), .ZN(n1057) );
  XNOR2_X1 U1684 ( .A(n1350), .B(n1541), .ZN(n1064) );
  XNOR2_X1 U1685 ( .A(n1336), .B(n1541), .ZN(n1054) );
  XNOR2_X1 U1686 ( .A(n1305), .B(n1541), .ZN(n1063) );
  XNOR2_X1 U1687 ( .A(n1552), .B(n1541), .ZN(n1065) );
  XNOR2_X1 U1688 ( .A(n1562), .B(n1541), .ZN(n1053) );
  XNOR2_X1 U1689 ( .A(n1346), .B(n1541), .ZN(n1066) );
  XNOR2_X1 U1690 ( .A(n1567), .B(n7), .ZN(n1048) );
  NAND2_X1 U1691 ( .A1(n755), .A2(n1234), .ZN(n1528) );
  NAND2_X1 U1692 ( .A1(n755), .A2(n719), .ZN(n1529) );
  NAND2_X1 U1693 ( .A1(n1234), .A2(n719), .ZN(n1530) );
  NAND3_X1 U1694 ( .A1(n1528), .A2(n1529), .A3(n1530), .ZN(n540) );
  XNOR2_X1 U1695 ( .A(n1351), .B(n1326), .ZN(n985) );
  XNOR2_X1 U1696 ( .A(n1566), .B(n1327), .ZN(n986) );
  XNOR2_X1 U1697 ( .A(n1565), .B(n1327), .ZN(n987) );
  XNOR2_X1 U1698 ( .A(n1563), .B(n1326), .ZN(n989) );
  XNOR2_X1 U1699 ( .A(n1564), .B(n1326), .ZN(n988) );
  XNOR2_X1 U1700 ( .A(n1338), .B(n1327), .ZN(n991) );
  XNOR2_X1 U1701 ( .A(n1562), .B(n1327), .ZN(n990) );
  XNOR2_X1 U1702 ( .A(n1550), .B(n1327), .ZN(n1004) );
  INV_X1 U1703 ( .A(n1326), .ZN(n1145) );
  XNOR2_X1 U1704 ( .A(n1346), .B(n1326), .ZN(n1003) );
  XNOR2_X1 U1705 ( .A(n1100), .B(n1327), .ZN(n995) );
  XNOR2_X1 U1706 ( .A(n1554), .B(n1327), .ZN(n999) );
  XNOR2_X1 U1707 ( .A(n1558), .B(n1544), .ZN(n994) );
  XNOR2_X1 U1708 ( .A(n1335), .B(n1327), .ZN(n993) );
  XNOR2_X1 U1709 ( .A(n1560), .B(n1327), .ZN(n992) );
  XNOR2_X1 U1710 ( .A(n1555), .B(n1544), .ZN(n998) );
  XNOR2_X1 U1711 ( .A(n1305), .B(n1326), .ZN(n1000) );
  XNOR2_X1 U1712 ( .A(n1102), .B(n1544), .ZN(n997) );
  XNOR2_X1 U1713 ( .A(n1553), .B(n1326), .ZN(n1001) );
  XNOR2_X1 U1714 ( .A(n1552), .B(n1326), .ZN(n1002) );
  XNOR2_X1 U1715 ( .A(n1352), .B(n1544), .ZN(n996) );
  XOR2_X1 U1716 ( .A(n25), .B(a[8]), .Z(n1115) );
  OAI21_X1 U1717 ( .B1(n166), .B2(n172), .A(n167), .ZN(n165) );
  XNOR2_X1 U1718 ( .A(n1351), .B(n1243), .ZN(n943) );
  XNOR2_X1 U1719 ( .A(n1566), .B(n1545), .ZN(n944) );
  XNOR2_X1 U1720 ( .A(n1355), .B(n1243), .ZN(n946) );
  XNOR2_X1 U1721 ( .A(n1565), .B(n1243), .ZN(n945) );
  XNOR2_X1 U1722 ( .A(n1563), .B(n1243), .ZN(n947) );
  XNOR2_X1 U1723 ( .A(n1334), .B(n1243), .ZN(n948) );
  XNOR2_X1 U1724 ( .A(n1338), .B(n1243), .ZN(n949) );
  XNOR2_X1 U1725 ( .A(n1335), .B(n1243), .ZN(n951) );
  XNOR2_X1 U1726 ( .A(n1347), .B(n1243), .ZN(n952) );
  XNOR2_X1 U1727 ( .A(n1560), .B(n1243), .ZN(n950) );
  INV_X1 U1728 ( .A(n1545), .ZN(n1143) );
  XNOR2_X1 U1729 ( .A(n1554), .B(n1243), .ZN(n957) );
  XNOR2_X1 U1730 ( .A(n1555), .B(n1243), .ZN(n956) );
  XNOR2_X1 U1731 ( .A(n1556), .B(n1243), .ZN(n955) );
  XNOR2_X1 U1732 ( .A(n1552), .B(n1243), .ZN(n960) );
  XNOR2_X1 U1733 ( .A(n1352), .B(n1243), .ZN(n954) );
  XNOR2_X1 U1734 ( .A(n1100), .B(n1243), .ZN(n953) );
  XNOR2_X1 U1735 ( .A(n1350), .B(n1545), .ZN(n959) );
  XNOR2_X1 U1736 ( .A(n1549), .B(n1545), .ZN(n962) );
  XNOR2_X1 U1737 ( .A(n1305), .B(n1545), .ZN(n958) );
  XNOR2_X1 U1738 ( .A(n1551), .B(n1545), .ZN(n961) );
  NAND2_X1 U1739 ( .A1(n1492), .A2(n1491), .ZN(n222) );
  NAND2_X1 U1740 ( .A1(n1492), .A2(n227), .ZN(n86) );
  INV_X1 U1741 ( .A(n200), .ZN(n198) );
  AOI21_X1 U1742 ( .B1(n173), .B2(n164), .A(n1418), .ZN(n163) );
  NAND2_X1 U1743 ( .A1(n397), .A2(n410), .ZN(n148) );
  INV_X1 U1744 ( .A(n1239), .ZN(n211) );
  OAI21_X1 U1745 ( .B1(n152), .B2(n150), .A(n1452), .ZN(n149) );
  NAND2_X1 U1746 ( .A1(n275), .A2(n1452), .ZN(n73) );
  XOR2_X1 U1747 ( .A(n303), .B(n306), .Z(n1531) );
  XOR2_X1 U1748 ( .A(n1531), .B(n1390), .Z(product[35]) );
  NAND2_X1 U1749 ( .A1(n303), .A2(n306), .ZN(n1532) );
  NAND2_X1 U1750 ( .A1(n303), .A2(n100), .ZN(n1533) );
  NAND2_X1 U1751 ( .A1(n1389), .A2(n306), .ZN(n1534) );
  NAND3_X1 U1752 ( .A1(n1533), .A2(n1534), .A3(n1532), .ZN(n99) );
  XOR2_X1 U1753 ( .A(n302), .B(n301), .Z(n1535) );
  XOR2_X1 U1754 ( .A(n1535), .B(n1443), .Z(product[36]) );
  NAND2_X1 U1755 ( .A1(n302), .A2(n301), .ZN(n1536) );
  NAND2_X1 U1756 ( .A1(n302), .A2(n1442), .ZN(n1537) );
  NAND2_X1 U1757 ( .A1(n99), .A2(n301), .ZN(n1538) );
  NAND3_X1 U1758 ( .A1(n1537), .A2(n1538), .A3(n1536), .ZN(n98) );
  AOI21_X1 U1759 ( .B1(n1296), .B2(n1282), .A(n1366), .ZN(n1539) );
  AOI21_X1 U1760 ( .B1(n1497), .B2(n1466), .A(n1366), .ZN(n181) );
  AOI21_X1 U1761 ( .B1(n221), .B2(n213), .A(n214), .ZN(n212) );
  AOI21_X1 U1762 ( .B1(n1492), .B2(n230), .A(n1297), .ZN(n223) );
  AOI21_X1 U1763 ( .B1(n203), .B2(n1489), .A(n198), .ZN(n196) );
  NAND2_X1 U1764 ( .A1(n202), .A2(n1489), .ZN(n195) );
  NAND2_X1 U1765 ( .A1(n1489), .A2(n200), .ZN(n81) );
  NOR2_X1 U1766 ( .A1(n177), .A2(n180), .ZN(n175) );
  AOI21_X1 U1767 ( .B1(n146), .B2(n133), .A(n134), .ZN(n132) );
  NAND2_X1 U1768 ( .A1(n411), .A2(n426), .ZN(n151) );
  XNOR2_X1 U1769 ( .A(n1351), .B(n1543), .ZN(n1006) );
  INV_X1 U1770 ( .A(n1254), .ZN(n1146) );
  XNOR2_X1 U1771 ( .A(n1550), .B(n1254), .ZN(n1025) );
  XNOR2_X1 U1772 ( .A(n1566), .B(n1543), .ZN(n1007) );
  XNOR2_X1 U1773 ( .A(n1346), .B(n1254), .ZN(n1024) );
  XNOR2_X1 U1774 ( .A(n1565), .B(n1543), .ZN(n1008) );
  XNOR2_X1 U1775 ( .A(n1564), .B(n1543), .ZN(n1009) );
  XNOR2_X1 U1776 ( .A(n1559), .B(n1543), .ZN(n1014) );
  XNOR2_X1 U1777 ( .A(n1554), .B(n1543), .ZN(n1020) );
  XNOR2_X1 U1778 ( .A(n1337), .B(n1543), .ZN(n1012) );
  XNOR2_X1 U1779 ( .A(n1560), .B(n1543), .ZN(n1013) );
  XNOR2_X1 U1780 ( .A(n1552), .B(n1543), .ZN(n1023) );
  XNOR2_X1 U1781 ( .A(n1555), .B(n1543), .ZN(n1019) );
  XNOR2_X1 U1782 ( .A(n1556), .B(n1543), .ZN(n1018) );
  XNOR2_X1 U1783 ( .A(n1562), .B(n1543), .ZN(n1011) );
  XNOR2_X1 U1784 ( .A(n1563), .B(n1543), .ZN(n1010) );
  XNOR2_X1 U1785 ( .A(n1356), .B(n1543), .ZN(n1016) );
  XNOR2_X1 U1786 ( .A(n1354), .B(n1543), .ZN(n1017) );
  XNOR2_X1 U1787 ( .A(n1543), .B(n1347), .ZN(n1015) );
  XNOR2_X1 U1788 ( .A(n1350), .B(n1543), .ZN(n1022) );
  XNOR2_X1 U1789 ( .A(n1306), .B(n1543), .ZN(n1021) );
  INV_X1 U1790 ( .A(n1278), .ZN(n193) );
  AOI21_X1 U1791 ( .B1(n194), .B2(n175), .A(n176), .ZN(n174) );
  INV_X1 U1792 ( .A(n1361), .ZN(n1147) );
  XNOR2_X1 U1793 ( .A(n1563), .B(n1361), .ZN(n1031) );
  XNOR2_X1 U1794 ( .A(n1107), .B(n1361), .ZN(n1044) );
  XNOR2_X1 U1795 ( .A(n1555), .B(n1361), .ZN(n1040) );
  XNOR2_X1 U1796 ( .A(n1556), .B(n1361), .ZN(n1039) );
  XNOR2_X1 U1797 ( .A(n1550), .B(n1361), .ZN(n1046) );
  XNOR2_X1 U1798 ( .A(n1336), .B(n1361), .ZN(n1033) );
  XNOR2_X1 U1799 ( .A(n1354), .B(n1361), .ZN(n1038) );
  XNOR2_X1 U1800 ( .A(n1562), .B(n1361), .ZN(n1032) );
  XNOR2_X1 U1801 ( .A(n1346), .B(n1361), .ZN(n1045) );
  XNOR2_X1 U1802 ( .A(n1553), .B(n1361), .ZN(n1043) );
  XNOR2_X1 U1803 ( .A(n1356), .B(n1361), .ZN(n1037) );
  XNOR2_X1 U1804 ( .A(n1554), .B(n1361), .ZN(n1041) );
  XNOR2_X1 U1805 ( .A(n1306), .B(n1361), .ZN(n1042) );
  XNOR2_X1 U1806 ( .A(n1565), .B(n1361), .ZN(n1029) );
  XNOR2_X1 U1807 ( .A(n1564), .B(n1361), .ZN(n1030) );
  XNOR2_X1 U1808 ( .A(n1566), .B(n1361), .ZN(n1028) );
  XNOR2_X1 U1809 ( .A(n1351), .B(n1361), .ZN(n1027) );
  XNOR2_X1 U1810 ( .A(n1347), .B(n1361), .ZN(n1036) );
  XNOR2_X1 U1811 ( .A(n1559), .B(n1361), .ZN(n1035) );
  XNOR2_X1 U1812 ( .A(n1560), .B(n1361), .ZN(n1034) );
  XOR2_X1 U1813 ( .A(n1542), .B(a[4]), .Z(n1117) );
  NAND2_X1 U1814 ( .A1(n156), .A2(n164), .ZN(n154) );
  AOI21_X1 U1815 ( .B1(n165), .B2(n156), .A(n157), .ZN(n155) );
  XNOR2_X1 U1816 ( .A(n1277), .B(n1566), .ZN(n923) );
  XNOR2_X1 U1817 ( .A(n1351), .B(n1277), .ZN(n922) );
  XNOR2_X1 U1818 ( .A(n1345), .B(n1277), .ZN(n924) );
  XNOR2_X1 U1819 ( .A(n1563), .B(n1277), .ZN(n926) );
  XNOR2_X1 U1820 ( .A(n1355), .B(n1277), .ZN(n925) );
  XNOR2_X1 U1821 ( .A(n1334), .B(n1277), .ZN(n927) );
  XNOR2_X1 U1822 ( .A(n1337), .B(n1277), .ZN(n928) );
  XNOR2_X1 U1823 ( .A(n1560), .B(n1277), .ZN(n929) );
  XNOR2_X1 U1824 ( .A(n1335), .B(n1546), .ZN(n930) );
  XNOR2_X1 U1825 ( .A(n1357), .B(n1546), .ZN(n932) );
  XNOR2_X1 U1826 ( .A(n1558), .B(n1546), .ZN(n931) );
  XNOR2_X1 U1827 ( .A(n1354), .B(n1546), .ZN(n933) );
  XNOR2_X1 U1828 ( .A(n1555), .B(n1546), .ZN(n935) );
  XNOR2_X1 U1829 ( .A(n1550), .B(n1546), .ZN(n941) );
  XNOR2_X1 U1830 ( .A(n1556), .B(n1546), .ZN(n934) );
  INV_X1 U1831 ( .A(n1546), .ZN(n1142) );
  XNOR2_X1 U1832 ( .A(n1346), .B(n1546), .ZN(n940) );
  XNOR2_X1 U1833 ( .A(n1552), .B(n1546), .ZN(n939) );
  XNOR2_X1 U1834 ( .A(n1349), .B(n1546), .ZN(n938) );
  XNOR2_X1 U1835 ( .A(n1554), .B(n1546), .ZN(n936) );
  INV_X1 U1836 ( .A(n1343), .ZN(n1149) );
  XNOR2_X1 U1837 ( .A(n1346), .B(n1343), .ZN(n1087) );
  XNOR2_X1 U1838 ( .A(n1552), .B(n1359), .ZN(n1086) );
  XNOR2_X1 U1839 ( .A(n1348), .B(n1344), .ZN(n1078) );
  XNOR2_X1 U1840 ( .A(n1563), .B(n1344), .ZN(n1073) );
  XNOR2_X1 U1841 ( .A(n1305), .B(n1359), .ZN(n1084) );
  XNOR2_X1 U1842 ( .A(n1562), .B(n1344), .ZN(n1074) );
  XNOR2_X1 U1843 ( .A(n1566), .B(n1359), .ZN(n1070) );
  XNOR2_X1 U1844 ( .A(n1565), .B(n1359), .ZN(n1071) );
  XNOR2_X1 U1845 ( .A(n1556), .B(n1359), .ZN(n1081) );
  XNOR2_X1 U1846 ( .A(n1559), .B(n1343), .ZN(n1077) );
  XNOR2_X1 U1847 ( .A(n1353), .B(n1343), .ZN(n1080) );
  XNOR2_X1 U1848 ( .A(n1560), .B(n1359), .ZN(n1076) );
  XNOR2_X1 U1849 ( .A(n1338), .B(n1343), .ZN(n1075) );
  XNOR2_X1 U1850 ( .A(n1564), .B(n1359), .ZN(n1072) );
  XNOR2_X1 U1851 ( .A(n1555), .B(n1343), .ZN(n1082) );
  XNOR2_X1 U1852 ( .A(n1554), .B(n1343), .ZN(n1083) );
  XNOR2_X1 U1853 ( .A(n1357), .B(n1359), .ZN(n1079) );
  XNOR2_X1 U1854 ( .A(n1349), .B(n1359), .ZN(n1085) );
  XNOR2_X1 U1855 ( .A(n1550), .B(n1359), .ZN(n1088) );
  NAND2_X1 U1856 ( .A1(n371), .A2(n382), .ZN(n136) );
  NOR2_X1 U1857 ( .A1(n140), .A2(n1248), .ZN(n133) );
  INV_X1 U1858 ( .A(n1248), .ZN(n272) );
  OAI21_X1 U1859 ( .B1(n141), .B2(n135), .A(n136), .ZN(n134) );
  NAND2_X1 U1860 ( .A1(n1296), .A2(n185), .ZN(n79) );
  NAND2_X1 U1861 ( .A1(n1299), .A2(n1497), .ZN(n180) );
  XNOR2_X1 U1862 ( .A(n1351), .B(n1455), .ZN(n964) );
  XNOR2_X1 U1863 ( .A(n1566), .B(n1454), .ZN(n965) );
  XNOR2_X1 U1864 ( .A(n1565), .B(n1455), .ZN(n966) );
  XNOR2_X1 U1865 ( .A(n1564), .B(n1454), .ZN(n967) );
  XNOR2_X1 U1866 ( .A(n1335), .B(n1455), .ZN(n972) );
  XNOR2_X1 U1867 ( .A(n1560), .B(n1454), .ZN(n971) );
  INV_X1 U1868 ( .A(n1454), .ZN(n1144) );
  XNOR2_X1 U1869 ( .A(n1337), .B(n1454), .ZN(n970) );
  XNOR2_X1 U1870 ( .A(n1562), .B(n1455), .ZN(n969) );
  XNOR2_X1 U1871 ( .A(n1563), .B(n1455), .ZN(n968) );
  XNOR2_X1 U1872 ( .A(n1549), .B(n1455), .ZN(n983) );
  XNOR2_X1 U1873 ( .A(n1551), .B(n1455), .ZN(n982) );
  XNOR2_X1 U1874 ( .A(n1556), .B(n1455), .ZN(n976) );
  XNOR2_X1 U1875 ( .A(n1353), .B(n1454), .ZN(n975) );
  XNOR2_X1 U1876 ( .A(n1348), .B(n1455), .ZN(n973) );
  XNOR2_X1 U1877 ( .A(n1356), .B(n1454), .ZN(n974) );
  XNOR2_X1 U1878 ( .A(n1104), .B(n1454), .ZN(n978) );
  XNOR2_X1 U1879 ( .A(n1305), .B(n1454), .ZN(n979) );
  XNOR2_X1 U1880 ( .A(n1555), .B(n1455), .ZN(n977) );
  XNOR2_X1 U1881 ( .A(n1349), .B(n1455), .ZN(n980) );
  XNOR2_X1 U1882 ( .A(n1552), .B(n1454), .ZN(n981) );
  OAI21_X1 U1883 ( .B1(n152), .B2(n131), .A(n1342), .ZN(n130) );
  INV_X1 U1884 ( .A(n1266), .ZN(n274) );
  NOR2_X1 U1885 ( .A1(n150), .A2(n1266), .ZN(n145) );
  OAI21_X1 U1886 ( .B1(n195), .B2(n212), .A(n196), .ZN(n194) );
  OAI21_X1 U1887 ( .B1(n222), .B2(n234), .A(n223), .ZN(n221) );
  AOI21_X1 U1888 ( .B1(n211), .B2(n202), .A(n203), .ZN(n201) );
  INV_X1 U1889 ( .A(n1339), .ZN(n284) );
  NOR2_X1 U1890 ( .A1(n1339), .A2(n209), .ZN(n202) );
  OAI21_X1 U1891 ( .B1(n204), .B2(n210), .A(n205), .ZN(n203) );
  INV_X1 U1892 ( .A(n1290), .ZN(n276) );
  OAI22_X1 U1893 ( .A1(n880), .A2(n1451), .B1(n880), .B2(n1407), .ZN(n640) );
  OAI22_X1 U1894 ( .A1(n1451), .A2(n881), .B1(n880), .B2(n1407), .ZN(n298) );
  OAI22_X1 U1895 ( .A1(n1451), .A2(n882), .B1(n881), .B2(n1407), .ZN(n681) );
  OAI22_X1 U1896 ( .A1(n1451), .A2(n883), .B1(n882), .B2(n1407), .ZN(n682) );
  OAI22_X1 U1897 ( .A1(n1451), .A2(n884), .B1(n883), .B2(n1407), .ZN(n683) );
  NOR2_X1 U1898 ( .A1(n161), .A2(n1477), .ZN(n156) );
  OAI21_X1 U1899 ( .B1(n158), .B2(n162), .A(n159), .ZN(n157) );
  OAI22_X1 U1900 ( .A1(n1451), .A2(n886), .B1(n885), .B2(n1407), .ZN(n685) );
  OAI22_X1 U1901 ( .A1(n1451), .A2(n885), .B1(n884), .B2(n1407), .ZN(n684) );
  NAND2_X1 U1902 ( .A1(n427), .A2(n442), .ZN(n159) );
  OAI22_X1 U1903 ( .A1(n1451), .A2(n887), .B1(n886), .B2(n1407), .ZN(n686) );
  OAI22_X1 U1904 ( .A1(n1451), .A2(n888), .B1(n887), .B2(n1407), .ZN(n687) );
  OAI22_X1 U1905 ( .A1(n60), .A2(n889), .B1(n888), .B2(n1407), .ZN(n688) );
  OAI22_X1 U1906 ( .A1(n60), .A2(n890), .B1(n889), .B2(n1407), .ZN(n689) );
  OAI22_X1 U1907 ( .A1(n60), .A2(n891), .B1(n890), .B2(n1514), .ZN(n690) );
  OAI22_X1 U1908 ( .A1(n60), .A2(n892), .B1(n891), .B2(n1514), .ZN(n691) );
  OAI22_X1 U1909 ( .A1(n60), .A2(n894), .B1(n893), .B2(n1514), .ZN(n693) );
  OAI22_X1 U1910 ( .A1(n60), .A2(n893), .B1(n892), .B2(n1514), .ZN(n692) );
  OAI22_X1 U1911 ( .A1(n60), .A2(n895), .B1(n894), .B2(n1514), .ZN(n694) );
  OAI22_X1 U1912 ( .A1(n60), .A2(n899), .B1(n898), .B2(n1514), .ZN(n698) );
  OAI22_X1 U1913 ( .A1(n60), .A2(n896), .B1(n895), .B2(n1514), .ZN(n695) );
  OAI22_X1 U1914 ( .A1(n60), .A2(n1140), .B1(n900), .B2(n1514), .ZN(n670) );
  OAI22_X1 U1915 ( .A1(n60), .A2(n1264), .B1(n896), .B2(n1514), .ZN(n696) );
  INV_X1 U1916 ( .A(n1514), .ZN(n641) );
  INV_X1 U1917 ( .A(n1473), .ZN(n278) );
  OAI22_X1 U1918 ( .A1(n922), .A2(n1406), .B1(n922), .B2(n1275), .ZN(n646) );
  NOR2_X1 U1919 ( .A1(n1473), .A2(n171), .ZN(n164) );
  OAI22_X1 U1920 ( .A1(n1406), .A2(n924), .B1(n923), .B2(n1275), .ZN(n721) );
  OAI22_X1 U1921 ( .A1(n1406), .A2(n923), .B1(n922), .B2(n1275), .ZN(n314) );
  NAND2_X1 U1922 ( .A1(n461), .A2(n478), .ZN(n167) );
  OAI22_X1 U1923 ( .A1(n1406), .A2(n925), .B1(n924), .B2(n1275), .ZN(n722) );
  OAI22_X1 U1924 ( .A1(n1406), .A2(n927), .B1(n926), .B2(n1275), .ZN(n724) );
  OAI22_X1 U1925 ( .A1(n1406), .A2(n926), .B1(n925), .B2(n1275), .ZN(n723) );
  OAI22_X1 U1926 ( .A1(n1406), .A2(n928), .B1(n927), .B2(n1513), .ZN(n725) );
  OAI22_X1 U1927 ( .A1(n1253), .A2(n929), .B1(n928), .B2(n1513), .ZN(n726) );
  OAI22_X1 U1928 ( .A1(n1253), .A2(n930), .B1(n929), .B2(n1513), .ZN(n727) );
  OAI22_X1 U1929 ( .A1(n1253), .A2(n933), .B1(n932), .B2(n1513), .ZN(n730) );
  OAI22_X1 U1930 ( .A1(n48), .A2(n931), .B1(n930), .B2(n1513), .ZN(n728) );
  OAI22_X1 U1931 ( .A1(n48), .A2(n932), .B1(n931), .B2(n1513), .ZN(n729) );
  OAI22_X1 U1932 ( .A1(n48), .A2(n1142), .B1(n942), .B2(n1513), .ZN(n672) );
  OAI22_X1 U1933 ( .A1(n48), .A2(n1267), .B1(n933), .B2(n1513), .ZN(n731) );
  OAI22_X1 U1934 ( .A1(n48), .A2(n939), .B1(n938), .B2(n1513), .ZN(n736) );
  OAI22_X1 U1935 ( .A1(n48), .A2(n935), .B1(n934), .B2(n1513), .ZN(n732) );
  OAI22_X1 U1936 ( .A1(n48), .A2(n936), .B1(n935), .B2(n1513), .ZN(n733) );
  OAI22_X1 U1937 ( .A1(n48), .A2(n940), .B1(n939), .B2(n1513), .ZN(n737) );
  OAI22_X1 U1938 ( .A1(n48), .A2(n941), .B1(n940), .B2(n1513), .ZN(n738) );
  OAI22_X1 U1939 ( .A1(n48), .A2(n1289), .B1(n936), .B2(n1513), .ZN(n734) );
  OAI22_X1 U1940 ( .A1(n48), .A2(n938), .B1(n1289), .B2(n1513), .ZN(n735) );
  INV_X1 U1941 ( .A(n1513), .ZN(n647) );
  OAI21_X1 U1942 ( .B1(n193), .B2(n180), .A(n1539), .ZN(n179) );
  OAI21_X1 U1943 ( .B1(n181), .B2(n177), .A(n178), .ZN(n176) );
  OAI22_X1 U1944 ( .A1(n1318), .A2(n1039), .B1(n1038), .B2(n1506), .ZN(n831)
         );
  OAI22_X1 U1945 ( .A1(n1318), .A2(n1041), .B1(n1040), .B2(n1507), .ZN(n833)
         );
  OAI22_X1 U1946 ( .A1(n1318), .A2(n1045), .B1(n1044), .B2(n1388), .ZN(n837)
         );
  OAI22_X1 U1947 ( .A1(n1318), .A2(n1031), .B1(n1030), .B2(n1507), .ZN(n823)
         );
  OAI22_X1 U1948 ( .A1(n1318), .A2(n1147), .B1(n1047), .B2(n1506), .ZN(n677)
         );
  OAI22_X1 U1949 ( .A1(n1318), .A2(n1034), .B1(n1033), .B2(n1506), .ZN(n826)
         );
  OAI22_X1 U1950 ( .A1(n1319), .A2(n1032), .B1(n1031), .B2(n1506), .ZN(n824)
         );
  OAI22_X1 U1951 ( .A1(n1318), .A2(n1028), .B1(n1027), .B2(n1506), .ZN(n424)
         );
  OAI22_X1 U1952 ( .A1(n1318), .A2(n1044), .B1(n1043), .B2(n1506), .ZN(n836)
         );
  OAI22_X1 U1953 ( .A1(n1318), .A2(n1038), .B1(n1037), .B2(n1507), .ZN(n830)
         );
  OAI22_X1 U1954 ( .A1(n1027), .A2(n1319), .B1(n1027), .B2(n1506), .ZN(n661)
         );
  OAI22_X1 U1955 ( .A1(n1481), .A2(n1030), .B1(n1029), .B2(n1506), .ZN(n822)
         );
  OAI22_X1 U1956 ( .A1(n1319), .A2(n1040), .B1(n1039), .B2(n1507), .ZN(n832)
         );
  OAI22_X1 U1957 ( .A1(n1319), .A2(n1037), .B1(n1036), .B2(n1506), .ZN(n829)
         );
  OAI22_X1 U1958 ( .A1(n1318), .A2(n1046), .B1(n1045), .B2(n1507), .ZN(n838)
         );
  OAI22_X1 U1959 ( .A1(n1481), .A2(n1036), .B1(n1035), .B2(n1506), .ZN(n828)
         );
  OAI22_X1 U1960 ( .A1(n1319), .A2(n1043), .B1(n1042), .B2(n1507), .ZN(n835)
         );
  OAI22_X1 U1961 ( .A1(n1481), .A2(n1033), .B1(n1032), .B2(n1507), .ZN(n825)
         );
  OAI22_X1 U1962 ( .A1(n1319), .A2(n1042), .B1(n1041), .B2(n1507), .ZN(n834)
         );
  OAI22_X1 U1963 ( .A1(n1481), .A2(n1035), .B1(n1034), .B2(n1507), .ZN(n827)
         );
  INV_X1 U1964 ( .A(n1506), .ZN(n662) );
  OAI21_X1 U1965 ( .B1(n147), .B2(n151), .A(n148), .ZN(n146) );
  XNOR2_X1 U1966 ( .A(n90), .B(n247), .ZN(product[6]) );
  XOR2_X1 U1967 ( .A(n1324), .B(n89), .Z(product[7]) );
  OAI21_X1 U1968 ( .B1(n242), .B2(n240), .A(n241), .ZN(n239) );
  AOI21_X1 U1969 ( .B1(n1502), .B2(n247), .A(n244), .ZN(n242) );
  INV_X1 U1970 ( .A(n1456), .ZN(n173) );
  OAI22_X1 U1971 ( .A1(n901), .A2(n1401), .B1(n901), .B2(n1412), .ZN(n643) );
  OAI22_X1 U1972 ( .A1(n1320), .A2(n902), .B1(n901), .B2(n1413), .ZN(n304) );
  OAI22_X1 U1973 ( .A1(n1401), .A2(n903), .B1(n902), .B2(n1412), .ZN(n701) );
  OAI22_X1 U1974 ( .A1(n1401), .A2(n905), .B1(n904), .B2(n1412), .ZN(n703) );
  OAI22_X1 U1975 ( .A1(n1320), .A2(n904), .B1(n903), .B2(n1413), .ZN(n702) );
  OAI22_X1 U1976 ( .A1(n1320), .A2(n906), .B1(n905), .B2(n1413), .ZN(n704) );
  OAI22_X1 U1977 ( .A1(n1401), .A2(n907), .B1(n906), .B2(n1412), .ZN(n705) );
  OAI22_X1 U1978 ( .A1(n1320), .A2(n908), .B1(n907), .B2(n1413), .ZN(n706) );
  OAI22_X1 U1979 ( .A1(n1401), .A2(n909), .B1(n908), .B2(n1412), .ZN(n707) );
  OAI22_X1 U1980 ( .A1(n1320), .A2(n910), .B1(n909), .B2(n1413), .ZN(n708) );
  OAI22_X1 U1981 ( .A1(n1401), .A2(n911), .B1(n910), .B2(n1412), .ZN(n709) );
  OAI22_X1 U1982 ( .A1(n1320), .A2(n912), .B1(n911), .B2(n1413), .ZN(n710) );
  OAI22_X1 U1983 ( .A1(n1320), .A2(n913), .B1(n912), .B2(n1412), .ZN(n711) );
  OAI22_X1 U1984 ( .A1(n1401), .A2(n915), .B1(n914), .B2(n1412), .ZN(n713) );
  OAI22_X1 U1985 ( .A1(n1320), .A2(n914), .B1(n913), .B2(n1413), .ZN(n712) );
  OAI22_X1 U1986 ( .A1(n1320), .A2(n1141), .B1(n921), .B2(n1413), .ZN(n671) );
  OAI22_X1 U1987 ( .A1(n1401), .A2(n919), .B1(n918), .B2(n1412), .ZN(n717) );
  OAI22_X1 U1988 ( .A1(n1320), .A2(n918), .B1(n917), .B2(n1412), .ZN(n716) );
  OAI22_X1 U1989 ( .A1(n1401), .A2(n916), .B1(n915), .B2(n1412), .ZN(n714) );
  OAI22_X1 U1990 ( .A1(n1401), .A2(n917), .B1(n916), .B2(n1413), .ZN(n715) );
  OAI22_X1 U1991 ( .A1(n54), .A2(n920), .B1(n919), .B2(n1413), .ZN(n718) );
  INV_X1 U1992 ( .A(n1413), .ZN(n644) );
  OAI21_X1 U1993 ( .B1(n132), .B2(n128), .A(n129), .ZN(n127) );
  OAI22_X1 U1994 ( .A1(n1341), .A2(n965), .B1(n964), .B2(n1402), .ZN(n346) );
  OAI22_X1 U1995 ( .A1(n964), .A2(n1341), .B1(n964), .B2(n1402), .ZN(n652) );
  OAI22_X1 U1996 ( .A1(n1341), .A2(n966), .B1(n965), .B2(n1402), .ZN(n761) );
  OAI22_X1 U1997 ( .A1(n1341), .A2(n967), .B1(n966), .B2(n1402), .ZN(n762) );
  OAI22_X1 U1998 ( .A1(n1341), .A2(n968), .B1(n967), .B2(n1402), .ZN(n763) );
  OAI22_X1 U1999 ( .A1(n1341), .A2(n973), .B1(n972), .B2(n1402), .ZN(n768) );
  OAI22_X1 U2000 ( .A1(n1341), .A2(n972), .B1(n971), .B2(n1402), .ZN(n767) );
  OAI22_X1 U2001 ( .A1(n36), .A2(n975), .B1(n974), .B2(n1402), .ZN(n770) );
  OAI22_X1 U2002 ( .A1(n36), .A2(n969), .B1(n968), .B2(n1402), .ZN(n764) );
  OAI22_X1 U2003 ( .A1(n1341), .A2(n971), .B1(n970), .B2(n1402), .ZN(n766) );
  OAI22_X1 U2004 ( .A1(n1341), .A2(n977), .B1(n976), .B2(n1402), .ZN(n772) );
  OAI22_X1 U2005 ( .A1(n1341), .A2(n1144), .B1(n984), .B2(n1402), .ZN(n674) );
  OAI22_X1 U2006 ( .A1(n36), .A2(n970), .B1(n969), .B2(n1402), .ZN(n765) );
  OAI22_X1 U2007 ( .A1(n36), .A2(n983), .B1(n982), .B2(n1402), .ZN(n778) );
  OAI22_X1 U2008 ( .A1(n1341), .A2(n976), .B1(n975), .B2(n1402), .ZN(n771) );
  OAI22_X1 U2009 ( .A1(n1341), .A2(n982), .B1(n1313), .B2(n1402), .ZN(n777) );
  OAI22_X1 U2010 ( .A1(n36), .A2(n979), .B1(n978), .B2(n1511), .ZN(n774) );
  OAI22_X1 U2011 ( .A1(n1341), .A2(n974), .B1(n973), .B2(n1511), .ZN(n769) );
  OAI22_X1 U2012 ( .A1(n1341), .A2(n980), .B1(n979), .B2(n1402), .ZN(n775) );
  OAI22_X1 U2013 ( .A1(n36), .A2(n978), .B1(n977), .B2(n1511), .ZN(n773) );
  OAI22_X1 U2014 ( .A1(n36), .A2(n981), .B1(n980), .B2(n1511), .ZN(n776) );
  INV_X1 U2015 ( .A(n1511), .ZN(n653) );
  AOI21_X1 U2016 ( .B1(n1480), .B2(n126), .A(n1475), .ZN(n125) );
  OAI21_X1 U2017 ( .B1(n174), .B2(n154), .A(n155), .ZN(n153) );
  INV_X1 U2018 ( .A(n101), .ZN(n264) );
  OAI22_X1 U2019 ( .A1(n985), .A2(n1242), .B1(n985), .B2(n1508), .ZN(n655) );
  OAI22_X1 U2020 ( .A1(n1242), .A2(n986), .B1(n985), .B2(n1509), .ZN(n368) );
  OAI22_X1 U2021 ( .A1(n1242), .A2(n987), .B1(n986), .B2(n1508), .ZN(n781) );
  OAI22_X1 U2022 ( .A1(n1241), .A2(n989), .B1(n988), .B2(n1509), .ZN(n783) );
  OAI22_X1 U2023 ( .A1(n1241), .A2(n992), .B1(n991), .B2(n1508), .ZN(n786) );
  OAI22_X1 U2024 ( .A1(n1242), .A2(n990), .B1(n989), .B2(n1509), .ZN(n784) );
  OAI22_X1 U2025 ( .A1(n1241), .A2(n1003), .B1(n1002), .B2(n1509), .ZN(n797)
         );
  OAI22_X1 U2026 ( .A1(n1242), .A2(n988), .B1(n987), .B2(n1508), .ZN(n782) );
  OAI22_X1 U2027 ( .A1(n1242), .A2(n991), .B1(n990), .B2(n1509), .ZN(n785) );
  OAI22_X1 U2028 ( .A1(n1478), .A2(n1310), .B1(n995), .B2(n1508), .ZN(n790) );
  OAI22_X1 U2029 ( .A1(n1242), .A2(n999), .B1(n998), .B2(n1509), .ZN(n793) );
  OAI22_X1 U2030 ( .A1(n1478), .A2(n994), .B1(n993), .B2(n1508), .ZN(n788) );
  OAI22_X1 U2031 ( .A1(n1242), .A2(n993), .B1(n992), .B2(n1508), .ZN(n787) );
  OAI22_X1 U2032 ( .A1(n1242), .A2(n1000), .B1(n999), .B2(n1508), .ZN(n794) );
  OAI22_X1 U2033 ( .A1(n1478), .A2(n995), .B1(n994), .B2(n1509), .ZN(n789) );
  OAI22_X1 U2034 ( .A1(n1241), .A2(n1002), .B1(n1001), .B2(n1509), .ZN(n796)
         );
  OAI22_X1 U2035 ( .A1(n1242), .A2(n1004), .B1(n1003), .B2(n1509), .ZN(n798)
         );
  INV_X1 U2036 ( .A(n1508), .ZN(n656) );
  OAI22_X1 U2037 ( .A1(n1242), .A2(n1145), .B1(n1005), .B2(n1508), .ZN(n675)
         );
  OAI22_X1 U2038 ( .A1(n1478), .A2(n1001), .B1(n1000), .B2(n1509), .ZN(n795)
         );
  OAI22_X1 U2039 ( .A1(n1478), .A2(n998), .B1(n997), .B2(n1508), .ZN(n792) );
  OAI22_X1 U2040 ( .A1(n1478), .A2(n997), .B1(n996), .B2(n1508), .ZN(n791) );
  BUF_X4 U2041 ( .A(n19), .Z(n1543) );
  OAI22_X1 U2042 ( .A1(n943), .A2(n1431), .B1(n943), .B2(n1453), .ZN(n649) );
  OAI22_X1 U2043 ( .A1(n1431), .A2(n944), .B1(n943), .B2(n1453), .ZN(n328) );
  OAI22_X1 U2044 ( .A1(n1431), .A2(n945), .B1(n944), .B2(n1453), .ZN(n741) );
  OAI22_X1 U2045 ( .A1(n1431), .A2(n947), .B1(n946), .B2(n1453), .ZN(n743) );
  OAI22_X1 U2046 ( .A1(n1431), .A2(n946), .B1(n945), .B2(n1453), .ZN(n742) );
  OAI22_X1 U2047 ( .A1(n1431), .A2(n948), .B1(n947), .B2(n1331), .ZN(n744) );
  OAI22_X1 U2048 ( .A1(n1396), .A2(n949), .B1(n948), .B2(n1331), .ZN(n745) );
  OAI22_X1 U2049 ( .A1(n1397), .A2(n952), .B1(n951), .B2(n1331), .ZN(n748) );
  OAI22_X1 U2050 ( .A1(n1396), .A2(n950), .B1(n949), .B2(n1510), .ZN(n746) );
  OAI22_X1 U2051 ( .A1(n1396), .A2(n951), .B1(n950), .B2(n1510), .ZN(n747) );
  OAI22_X1 U2052 ( .A1(n1396), .A2(n953), .B1(n952), .B2(n1510), .ZN(n749) );
  OAI22_X1 U2053 ( .A1(n1396), .A2(n957), .B1(n956), .B2(n1331), .ZN(n753) );
  OAI22_X1 U2054 ( .A1(n1397), .A2(n956), .B1(n955), .B2(n1510), .ZN(n752) );
  OAI22_X1 U2055 ( .A1(n1397), .A2(n1329), .B1(n957), .B2(n1510), .ZN(n754) );
  OAI22_X1 U2056 ( .A1(n42), .A2(n955), .B1(n954), .B2(n1510), .ZN(n751) );
  OAI22_X1 U2057 ( .A1(n1397), .A2(n1143), .B1(n963), .B2(n1331), .ZN(n673) );
  OAI22_X1 U2058 ( .A1(n1396), .A2(n954), .B1(n953), .B2(n1510), .ZN(n750) );
  OAI22_X1 U2059 ( .A1(n1397), .A2(n960), .B1(n959), .B2(n1510), .ZN(n756) );
  OAI22_X1 U2060 ( .A1(n1397), .A2(n961), .B1(n960), .B2(n1510), .ZN(n757) );
  INV_X1 U2061 ( .A(n1510), .ZN(n650) );
  OAI22_X1 U2062 ( .A1(n42), .A2(n962), .B1(n1510), .B2(n961), .ZN(n758) );
  XNOR2_X1 U2063 ( .A(n1445), .B(n67), .ZN(product[29]) );
  XNOR2_X1 U2064 ( .A(n1400), .B(n65), .ZN(product[31]) );
  OAI22_X1 U2065 ( .A1(n1370), .A2(n1014), .B1(n1013), .B2(n1308), .ZN(n807)
         );
  OAI22_X1 U2066 ( .A1(n1370), .A2(n1007), .B1(n1006), .B2(n1308), .ZN(n394)
         );
  OAI22_X1 U2067 ( .A1(n1006), .A2(n1371), .B1(n1006), .B2(n1308), .ZN(n658)
         );
  OAI22_X1 U2068 ( .A1(n1371), .A2(n1012), .B1(n1011), .B2(n1308), .ZN(n805)
         );
  OAI22_X1 U2069 ( .A1(n1371), .A2(n1008), .B1(n1007), .B2(n1308), .ZN(n801)
         );
  OAI22_X1 U2070 ( .A1(n1371), .A2(n1021), .B1(n1020), .B2(n1512), .ZN(n814)
         );
  OAI22_X1 U2071 ( .A1(n1370), .A2(n1024), .B1(n1023), .B2(n1308), .ZN(n817)
         );
  OAI22_X1 U2072 ( .A1(n1371), .A2(n1009), .B1(n1008), .B2(n1512), .ZN(n802)
         );
  OAI22_X1 U2073 ( .A1(n1371), .A2(n1010), .B1(n1009), .B2(n1512), .ZN(n803)
         );
  OAI22_X1 U2074 ( .A1(n1370), .A2(n1015), .B1(n1014), .B2(n1308), .ZN(n808)
         );
  OAI22_X1 U2075 ( .A1(n24), .A2(n1013), .B1(n1012), .B2(n1308), .ZN(n806) );
  OAI22_X1 U2076 ( .A1(n1371), .A2(n1146), .B1(n1026), .B2(n1512), .ZN(n676)
         );
  OAI22_X1 U2077 ( .A1(n1371), .A2(n1011), .B1(n1010), .B2(n1512), .ZN(n804)
         );
  OAI22_X1 U2078 ( .A1(n1370), .A2(n1025), .B1(n1024), .B2(n1512), .ZN(n818)
         );
  OAI22_X1 U2079 ( .A1(n1371), .A2(n1019), .B1(n1018), .B2(n1512), .ZN(n812)
         );
  OAI22_X1 U2080 ( .A1(n1370), .A2(n1020), .B1(n1019), .B2(n1308), .ZN(n813)
         );
  OAI22_X1 U2081 ( .A1(n1371), .A2(n1018), .B1(n1017), .B2(n1512), .ZN(n811)
         );
  OAI22_X1 U2082 ( .A1(n1370), .A2(n1017), .B1(n1016), .B2(n1512), .ZN(n810)
         );
  OAI22_X1 U2083 ( .A1(n1370), .A2(n1023), .B1(n1022), .B2(n1308), .ZN(n816)
         );
  OAI22_X1 U2084 ( .A1(n1016), .A2(n24), .B1(n1015), .B2(n1308), .ZN(n809) );
  OAI22_X1 U2085 ( .A1(n1370), .A2(n1022), .B1(n1021), .B2(n1512), .ZN(n815)
         );
  INV_X1 U2086 ( .A(n1512), .ZN(n659) );
  OAI21_X1 U2087 ( .B1(n248), .B2(n250), .A(n249), .ZN(n247) );
  AOI21_X1 U2088 ( .B1(n114), .B2(n1495), .A(n111), .ZN(n109) );
  OAI21_X1 U2089 ( .B1(n1483), .B2(n123), .A(n124), .ZN(n122) );
  AOI21_X1 U2090 ( .B1(n1445), .B2(n1494), .A(n119), .ZN(n117) );
  XNOR2_X1 U2091 ( .A(n1460), .B(n63), .ZN(product[33]) );
  XOR2_X1 U2092 ( .A(n1444), .B(n64), .Z(product[32]) );
  XOR2_X1 U2093 ( .A(n117), .B(n66), .Z(product[30]) );
  XOR2_X1 U2094 ( .A(n125), .B(n68), .Z(product[28]) );
  AOI21_X1 U2095 ( .B1(n106), .B2(n1496), .A(n103), .ZN(n101) );
  OAI21_X1 U2096 ( .B1(n109), .B2(n107), .A(n108), .ZN(n106) );
  OAI21_X1 U2097 ( .B1(n1476), .B2(n115), .A(n116), .ZN(n114) );
  OAI22_X1 U2098 ( .A1(n1463), .A2(n1055), .B1(n1054), .B2(n1322), .ZN(n846)
         );
  OAI22_X1 U2099 ( .A1(n1463), .A2(n1051), .B1(n1050), .B2(n1322), .ZN(n842)
         );
  OAI22_X1 U2100 ( .A1(n1464), .A2(n1062), .B1(n1061), .B2(n1321), .ZN(n853)
         );
  OAI22_X1 U2101 ( .A1(n1463), .A2(n1059), .B1(n1058), .B2(n1321), .ZN(n850)
         );
  OAI22_X1 U2102 ( .A1(n1279), .A2(n1060), .B1(n1059), .B2(n1321), .ZN(n851)
         );
  OAI22_X1 U2103 ( .A1(n1280), .A2(n1053), .B1(n1052), .B2(n1322), .ZN(n844)
         );
  OAI22_X1 U2104 ( .A1(n1464), .A2(n1049), .B1(n1048), .B2(n1322), .ZN(n458)
         );
  OAI22_X1 U2105 ( .A1(n1463), .A2(n1052), .B1(n1051), .B2(n1321), .ZN(n843)
         );
  OAI22_X1 U2106 ( .A1(n1464), .A2(n1063), .B1(n1062), .B2(n1322), .ZN(n854)
         );
  OAI22_X1 U2107 ( .A1(n1279), .A2(n1050), .B1(n1049), .B2(n1322), .ZN(n841)
         );
  OAI22_X1 U2108 ( .A1(n1464), .A2(n1057), .B1(n1056), .B2(n1321), .ZN(n848)
         );
  OAI22_X1 U2109 ( .A1(n1279), .A2(n1065), .B1(n1064), .B2(n1322), .ZN(n856)
         );
  OAI22_X1 U2110 ( .A1(n1280), .A2(n1056), .B1(n1055), .B2(n1322), .ZN(n847)
         );
  OAI22_X1 U2111 ( .A1(n1464), .A2(n1058), .B1(n1057), .B2(n1322), .ZN(n849)
         );
  OAI22_X1 U2112 ( .A1(n1464), .A2(n1148), .B1(n1068), .B2(n1321), .ZN(n678)
         );
  OAI22_X1 U2113 ( .A1(n1280), .A2(n1054), .B1(n1053), .B2(n1322), .ZN(n845)
         );
  OAI22_X1 U2114 ( .A1(n1279), .A2(n1061), .B1(n1060), .B2(n1321), .ZN(n852)
         );
  OAI22_X1 U2115 ( .A1(n1048), .A2(n12), .B1(n1048), .B2(n9), .ZN(n664) );
  OAI22_X1 U2116 ( .A1(n1463), .A2(n1064), .B1(n1063), .B2(n1322), .ZN(n855)
         );
  OAI22_X1 U2117 ( .A1(n1279), .A2(n1067), .B1(n1066), .B2(n1322), .ZN(n858)
         );
  OAI22_X1 U2118 ( .A1(n1280), .A2(n1066), .B1(n1065), .B2(n1321), .ZN(n857)
         );
endmodule


module mac_5_DW01_add_1 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n34, n35, n36, n37, n38, n39, n40, n41, n43, n45, n46, n47,
         n48, n49, n51, n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65,
         n67, n69, n70, n71, n72, n73, n75, n77, n78, n79, n80, n81, n83, n85,
         n86, n87, n88, n89, n91, n93, n94, n95, n96, n97, n99, n101, n102,
         n103, n104, n105, n107, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n119, n121, n122, n124, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n184, n185, n187, n189, n191,
         n193, n195, n197, n199, n201, n203, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407;

  FA_X1 U3 ( .A(B[38]), .B(A[38]), .CI(n35), .CO(n34), .S(SUM[38]) );
  FA_X1 U6 ( .A(B[35]), .B(A[35]), .CI(n38), .CO(n37), .S(SUM[35]) );
  FA_X1 U7 ( .A(B[34]), .B(A[34]), .CI(n39), .CO(n38), .S(SUM[34]) );
  OR2_X1 U254 ( .A1(B[0]), .A2(A[0]), .ZN(n344) );
  XOR2_X1 U255 ( .A(B[36]), .B(A[36]), .Z(n345) );
  XOR2_X1 U256 ( .A(n37), .B(n345), .Z(SUM[36]) );
  NAND2_X1 U257 ( .A1(n37), .A2(B[36]), .ZN(n346) );
  NAND2_X1 U258 ( .A1(n37), .A2(A[36]), .ZN(n347) );
  NAND2_X1 U259 ( .A1(B[36]), .A2(A[36]), .ZN(n348) );
  NAND3_X1 U260 ( .A1(n346), .A2(n347), .A3(n348), .ZN(n36) );
  XOR2_X1 U261 ( .A(B[37]), .B(A[37]), .Z(n349) );
  XOR2_X1 U262 ( .A(n36), .B(n349), .Z(SUM[37]) );
  NAND2_X1 U263 ( .A1(n36), .A2(B[37]), .ZN(n350) );
  NAND2_X1 U264 ( .A1(n36), .A2(A[37]), .ZN(n351) );
  NAND2_X1 U265 ( .A1(B[37]), .A2(A[37]), .ZN(n352) );
  NAND3_X1 U266 ( .A1(n350), .A2(n351), .A3(n352), .ZN(n35) );
  NAND3_X1 U267 ( .A1(n381), .A2(n382), .A3(n383), .ZN(n353) );
  NAND3_X1 U268 ( .A1(n381), .A2(n382), .A3(n383), .ZN(n354) );
  XOR2_X1 U269 ( .A(B[33]), .B(A[33]), .Z(n355) );
  XOR2_X1 U270 ( .A(n354), .B(n355), .Z(SUM[33]) );
  NAND2_X1 U271 ( .A1(n353), .A2(B[33]), .ZN(n356) );
  NAND2_X1 U272 ( .A1(n40), .A2(A[33]), .ZN(n357) );
  NAND2_X1 U273 ( .A1(B[33]), .A2(A[33]), .ZN(n358) );
  NAND3_X1 U274 ( .A1(n356), .A2(n357), .A3(n358), .ZN(n39) );
  CLKBUF_X1 U275 ( .A(n110), .Z(n359) );
  CLKBUF_X1 U276 ( .A(n70), .Z(n360) );
  INV_X1 U277 ( .A(n136), .ZN(n361) );
  NOR2_X1 U278 ( .A1(B[9]), .A2(A[9]), .ZN(n362) );
  NOR2_X1 U279 ( .A1(B[9]), .A2(A[9]), .ZN(n144) );
  NOR2_X1 U280 ( .A1(B[3]), .A2(A[3]), .ZN(n363) );
  NOR2_X1 U281 ( .A1(B[3]), .A2(A[3]), .ZN(n174) );
  CLKBUF_X1 U282 ( .A(n130), .Z(n364) );
  NOR2_X1 U283 ( .A1(B[5]), .A2(A[5]), .ZN(n365) );
  AOI21_X1 U284 ( .B1(n172), .B2(n180), .A(n173), .ZN(n366) );
  NOR2_X1 U285 ( .A1(B[7]), .A2(A[7]), .ZN(n367) );
  CLKBUF_X1 U286 ( .A(n150), .Z(n368) );
  CLKBUF_X1 U287 ( .A(n143), .Z(n369) );
  NOR2_X1 U288 ( .A1(B[11]), .A2(A[11]), .ZN(n370) );
  NOR2_X1 U289 ( .A1(B[11]), .A2(A[11]), .ZN(n132) );
  CLKBUF_X1 U290 ( .A(n185), .Z(n371) );
  AOI21_X1 U291 ( .B1(n359), .B2(n401), .A(n107), .ZN(n372) );
  AOI21_X1 U292 ( .B1(n110), .B2(n401), .A(n107), .ZN(n105) );
  AOI21_X1 U293 ( .B1(n360), .B2(n403), .A(n67), .ZN(n373) );
  AOI21_X1 U294 ( .B1(n70), .B2(n403), .A(n67), .ZN(n65) );
  CLKBUF_X1 U295 ( .A(n131), .Z(n374) );
  AOI21_X1 U296 ( .B1(n364), .B2(n369), .A(n374), .ZN(n375) );
  CLKBUF_X1 U297 ( .A(n115), .Z(n376) );
  CLKBUF_X1 U298 ( .A(n62), .Z(n377) );
  CLKBUF_X1 U299 ( .A(n54), .Z(n378) );
  CLKBUF_X1 U300 ( .A(n78), .Z(n379) );
  XOR2_X1 U301 ( .A(B[32]), .B(A[32]), .Z(n380) );
  XOR2_X1 U302 ( .A(n371), .B(n380), .Z(SUM[32]) );
  NAND2_X1 U303 ( .A1(n185), .A2(B[32]), .ZN(n381) );
  NAND2_X1 U304 ( .A1(n185), .A2(A[32]), .ZN(n382) );
  NAND2_X1 U305 ( .A1(B[32]), .A2(A[32]), .ZN(n383) );
  NAND3_X1 U306 ( .A1(n381), .A2(n382), .A3(n383), .ZN(n40) );
  AOI21_X1 U307 ( .B1(n377), .B2(n404), .A(n59), .ZN(n384) );
  AOI21_X1 U308 ( .B1(n378), .B2(n405), .A(n51), .ZN(n385) );
  CLKBUF_X1 U309 ( .A(n102), .Z(n386) );
  CLKBUF_X1 U310 ( .A(n94), .Z(n387) );
  CLKBUF_X1 U311 ( .A(n46), .Z(n388) );
  CLKBUF_X1 U312 ( .A(n86), .Z(n389) );
  AOI21_X1 U313 ( .B1(n386), .B2(n399), .A(n99), .ZN(n390) );
  AOI21_X1 U314 ( .B1(n368), .B2(n114), .A(n376), .ZN(n391) );
  AOI21_X1 U315 ( .B1(n102), .B2(n399), .A(n99), .ZN(n97) );
  AOI21_X1 U316 ( .B1(n150), .B2(n114), .A(n115), .ZN(n113) );
  AOI21_X1 U317 ( .B1(n389), .B2(n400), .A(n83), .ZN(n392) );
  AOI21_X1 U318 ( .B1(n86), .B2(n400), .A(n83), .ZN(n81) );
  AOI21_X1 U319 ( .B1(n379), .B2(n402), .A(n75), .ZN(n393) );
  AOI21_X1 U320 ( .B1(n387), .B2(n398), .A(n91), .ZN(n394) );
  INV_X1 U321 ( .A(n368), .ZN(n149) );
  OAI21_X1 U322 ( .B1(n149), .B2(n128), .A(n375), .ZN(n127) );
  OAI21_X1 U323 ( .B1(n149), .B2(n140), .A(n141), .ZN(n139) );
  INV_X1 U324 ( .A(n369), .ZN(n141) );
  INV_X1 U325 ( .A(n142), .ZN(n140) );
  NAND2_X1 U326 ( .A1(n142), .A2(n130), .ZN(n128) );
  AOI21_X1 U327 ( .B1(n170), .B2(n161), .A(n162), .ZN(n160) );
  INV_X1 U328 ( .A(n366), .ZN(n170) );
  INV_X1 U329 ( .A(n180), .ZN(n179) );
  INV_X1 U330 ( .A(n85), .ZN(n83) );
  INV_X1 U331 ( .A(n77), .ZN(n75) );
  INV_X1 U332 ( .A(n61), .ZN(n59) );
  INV_X1 U333 ( .A(n53), .ZN(n51) );
  INV_X1 U334 ( .A(n109), .ZN(n107) );
  AOI21_X1 U335 ( .B1(n130), .B2(n143), .A(n131), .ZN(n129) );
  OAI21_X1 U336 ( .B1(n132), .B2(n138), .A(n133), .ZN(n131) );
  OAI21_X1 U337 ( .B1(n163), .B2(n169), .A(n164), .ZN(n162) );
  AOI21_X1 U338 ( .B1(n172), .B2(n180), .A(n173), .ZN(n171) );
  NOR2_X1 U339 ( .A1(n177), .A2(n363), .ZN(n172) );
  OAI21_X1 U340 ( .B1(n174), .B2(n178), .A(n175), .ZN(n173) );
  INV_X1 U341 ( .A(n69), .ZN(n67) );
  AOI21_X1 U342 ( .B1(n94), .B2(n398), .A(n91), .ZN(n89) );
  INV_X1 U343 ( .A(n93), .ZN(n91) );
  INV_X1 U344 ( .A(n101), .ZN(n99) );
  OAI21_X1 U345 ( .B1(n144), .B2(n148), .A(n145), .ZN(n143) );
  NOR2_X1 U346 ( .A1(n168), .A2(n365), .ZN(n161) );
  OAI21_X1 U347 ( .B1(n181), .B2(n184), .A(n182), .ZN(n180) );
  NOR2_X1 U348 ( .A1(n137), .A2(n370), .ZN(n130) );
  OAI21_X1 U349 ( .B1(n171), .B2(n151), .A(n152), .ZN(n150) );
  NAND2_X1 U350 ( .A1(n161), .A2(n153), .ZN(n151) );
  AOI21_X1 U351 ( .B1(n153), .B2(n162), .A(n154), .ZN(n152) );
  NOR2_X1 U352 ( .A1(n158), .A2(n367), .ZN(n153) );
  AOI21_X1 U353 ( .B1(n397), .B2(n124), .A(n119), .ZN(n117) );
  INV_X1 U354 ( .A(n121), .ZN(n119) );
  NAND2_X1 U355 ( .A1(n195), .A2(n80), .ZN(n11) );
  INV_X1 U356 ( .A(n79), .ZN(n195) );
  NAND2_X1 U357 ( .A1(n197), .A2(n88), .ZN(n13) );
  INV_X1 U358 ( .A(n87), .ZN(n197) );
  NAND2_X1 U359 ( .A1(n199), .A2(n96), .ZN(n15) );
  INV_X1 U360 ( .A(n95), .ZN(n199) );
  NAND2_X1 U361 ( .A1(n201), .A2(n104), .ZN(n17) );
  INV_X1 U362 ( .A(n103), .ZN(n201) );
  NOR2_X1 U363 ( .A1(n128), .A2(n116), .ZN(n114) );
  OAI21_X1 U364 ( .B1(n129), .B2(n116), .A(n117), .ZN(n115) );
  NAND2_X1 U365 ( .A1(n396), .A2(n397), .ZN(n116) );
  NOR2_X1 U366 ( .A1(n147), .A2(n362), .ZN(n142) );
  INV_X1 U367 ( .A(n126), .ZN(n124) );
  OAI21_X1 U368 ( .B1(n155), .B2(n159), .A(n156), .ZN(n154) );
  NAND2_X1 U369 ( .A1(n187), .A2(n48), .ZN(n3) );
  INV_X1 U370 ( .A(n47), .ZN(n187) );
  NAND2_X1 U371 ( .A1(n189), .A2(n56), .ZN(n5) );
  INV_X1 U372 ( .A(n55), .ZN(n189) );
  NAND2_X1 U373 ( .A1(n191), .A2(n64), .ZN(n7) );
  INV_X1 U374 ( .A(n63), .ZN(n191) );
  NAND2_X1 U375 ( .A1(n193), .A2(n72), .ZN(n9) );
  INV_X1 U376 ( .A(n71), .ZN(n193) );
  NAND2_X1 U377 ( .A1(n406), .A2(n45), .ZN(n2) );
  NAND2_X1 U378 ( .A1(n405), .A2(n53), .ZN(n4) );
  NAND2_X1 U379 ( .A1(n404), .A2(n61), .ZN(n6) );
  NAND2_X1 U380 ( .A1(n403), .A2(n69), .ZN(n8) );
  NAND2_X1 U381 ( .A1(n402), .A2(n77), .ZN(n10) );
  NAND2_X1 U382 ( .A1(n400), .A2(n85), .ZN(n12) );
  NAND2_X1 U383 ( .A1(n398), .A2(n93), .ZN(n14) );
  NAND2_X1 U384 ( .A1(n399), .A2(n101), .ZN(n16) );
  XOR2_X1 U385 ( .A(n122), .B(n20), .Z(SUM[13]) );
  NAND2_X1 U386 ( .A1(n397), .A2(n121), .ZN(n20) );
  AOI21_X1 U387 ( .B1(n127), .B2(n396), .A(n124), .ZN(n122) );
  XOR2_X1 U388 ( .A(n134), .B(n22), .Z(SUM[11]) );
  NAND2_X1 U389 ( .A1(n206), .A2(n133), .ZN(n22) );
  AOI21_X1 U390 ( .B1(n139), .B2(n207), .A(n136), .ZN(n134) );
  INV_X1 U391 ( .A(n137), .ZN(n207) );
  INV_X1 U392 ( .A(n168), .ZN(n213) );
  XOR2_X1 U393 ( .A(n160), .B(n27), .Z(SUM[6]) );
  NAND2_X1 U394 ( .A1(n211), .A2(n159), .ZN(n27) );
  INV_X1 U395 ( .A(n158), .ZN(n211) );
  INV_X1 U396 ( .A(n370), .ZN(n206) );
  INV_X1 U397 ( .A(n138), .ZN(n136) );
  INV_X1 U398 ( .A(n169), .ZN(n167) );
  INV_X1 U399 ( .A(n362), .ZN(n208) );
  INV_X1 U400 ( .A(n367), .ZN(n210) );
  INV_X1 U401 ( .A(n365), .ZN(n212) );
  INV_X1 U402 ( .A(n363), .ZN(n214) );
  XOR2_X1 U403 ( .A(n165), .B(n28), .Z(SUM[5]) );
  NAND2_X1 U404 ( .A1(n212), .A2(n164), .ZN(n28) );
  AOI21_X1 U405 ( .B1(n170), .B2(n213), .A(n167), .ZN(n165) );
  XNOR2_X1 U406 ( .A(n170), .B(n29), .ZN(SUM[4]) );
  NAND2_X1 U407 ( .A1(n213), .A2(n169), .ZN(n29) );
  XNOR2_X1 U408 ( .A(n176), .B(n30), .ZN(SUM[3]) );
  NAND2_X1 U409 ( .A1(n214), .A2(n175), .ZN(n30) );
  OAI21_X1 U410 ( .B1(n179), .B2(n177), .A(n178), .ZN(n176) );
  XOR2_X1 U411 ( .A(n179), .B(n31), .Z(SUM[2]) );
  NAND2_X1 U412 ( .A1(n215), .A2(n178), .ZN(n31) );
  INV_X1 U413 ( .A(n177), .ZN(n215) );
  XOR2_X1 U414 ( .A(n32), .B(n184), .Z(SUM[1]) );
  NAND2_X1 U415 ( .A1(n216), .A2(n182), .ZN(n32) );
  INV_X1 U416 ( .A(n181), .ZN(n216) );
  AND2_X1 U417 ( .A1(n344), .A2(n184), .ZN(SUM[0]) );
  NAND2_X1 U418 ( .A1(n203), .A2(n112), .ZN(n19) );
  INV_X1 U419 ( .A(n111), .ZN(n203) );
  NAND2_X1 U420 ( .A1(n401), .A2(n109), .ZN(n18) );
  XNOR2_X1 U421 ( .A(n127), .B(n21), .ZN(SUM[12]) );
  NAND2_X1 U422 ( .A1(n396), .A2(n126), .ZN(n21) );
  XNOR2_X1 U423 ( .A(n139), .B(n23), .ZN(SUM[10]) );
  NAND2_X1 U424 ( .A1(n207), .A2(n361), .ZN(n23) );
  XNOR2_X1 U425 ( .A(n146), .B(n24), .ZN(SUM[9]) );
  NAND2_X1 U426 ( .A1(n208), .A2(n145), .ZN(n24) );
  OAI21_X1 U427 ( .B1(n149), .B2(n147), .A(n148), .ZN(n146) );
  XOR2_X1 U428 ( .A(n149), .B(n25), .Z(SUM[8]) );
  NAND2_X1 U429 ( .A1(n209), .A2(n148), .ZN(n25) );
  INV_X1 U430 ( .A(n147), .ZN(n209) );
  XNOR2_X1 U431 ( .A(n157), .B(n26), .ZN(SUM[7]) );
  NAND2_X1 U432 ( .A1(n210), .A2(n156), .ZN(n26) );
  OAI21_X1 U433 ( .B1(n160), .B2(n158), .A(n159), .ZN(n157) );
  NOR2_X1 U434 ( .A1(B[6]), .A2(A[6]), .ZN(n158) );
  NOR2_X1 U435 ( .A1(B[2]), .A2(A[2]), .ZN(n177) );
  NOR2_X1 U436 ( .A1(B[8]), .A2(A[8]), .ZN(n147) );
  NOR2_X1 U437 ( .A1(B[5]), .A2(A[5]), .ZN(n163) );
  NOR2_X1 U438 ( .A1(B[7]), .A2(A[7]), .ZN(n155) );
  OR2_X1 U439 ( .A1(B[12]), .A2(A[12]), .ZN(n396) );
  OR2_X1 U440 ( .A1(B[13]), .A2(A[13]), .ZN(n397) );
  NAND2_X1 U441 ( .A1(B[11]), .A2(A[11]), .ZN(n133) );
  NOR2_X1 U442 ( .A1(B[10]), .A2(A[10]), .ZN(n137) );
  NOR2_X1 U443 ( .A1(B[4]), .A2(A[4]), .ZN(n168) );
  NOR2_X1 U444 ( .A1(B[1]), .A2(A[1]), .ZN(n181) );
  NAND2_X1 U445 ( .A1(B[8]), .A2(A[8]), .ZN(n148) );
  NAND2_X1 U446 ( .A1(B[2]), .A2(A[2]), .ZN(n178) );
  NAND2_X1 U447 ( .A1(B[6]), .A2(A[6]), .ZN(n159) );
  NAND2_X1 U448 ( .A1(B[0]), .A2(A[0]), .ZN(n184) );
  NAND2_X1 U449 ( .A1(B[10]), .A2(A[10]), .ZN(n138) );
  NAND2_X1 U450 ( .A1(B[4]), .A2(A[4]), .ZN(n169) );
  NAND2_X1 U451 ( .A1(B[9]), .A2(A[9]), .ZN(n145) );
  NAND2_X1 U452 ( .A1(B[3]), .A2(A[3]), .ZN(n175) );
  NAND2_X1 U453 ( .A1(B[1]), .A2(A[1]), .ZN(n182) );
  NAND2_X1 U454 ( .A1(B[5]), .A2(A[5]), .ZN(n164) );
  NAND2_X1 U455 ( .A1(B[7]), .A2(A[7]), .ZN(n156) );
  INV_X1 U456 ( .A(n45), .ZN(n43) );
  NOR2_X1 U457 ( .A1(B[20]), .A2(A[20]), .ZN(n87) );
  NOR2_X1 U458 ( .A1(B[18]), .A2(A[18]), .ZN(n95) );
  NOR2_X1 U459 ( .A1(B[14]), .A2(A[14]), .ZN(n111) );
  NOR2_X1 U460 ( .A1(B[16]), .A2(A[16]), .ZN(n103) );
  NOR2_X1 U461 ( .A1(B[30]), .A2(A[30]), .ZN(n47) );
  NOR2_X1 U462 ( .A1(B[28]), .A2(A[28]), .ZN(n55) );
  NOR2_X1 U463 ( .A1(B[26]), .A2(A[26]), .ZN(n63) );
  NOR2_X1 U464 ( .A1(B[24]), .A2(A[24]), .ZN(n71) );
  NOR2_X1 U465 ( .A1(B[22]), .A2(A[22]), .ZN(n79) );
  OR2_X1 U466 ( .A1(B[19]), .A2(A[19]), .ZN(n398) );
  OR2_X1 U467 ( .A1(B[17]), .A2(A[17]), .ZN(n399) );
  NAND2_X1 U468 ( .A1(B[21]), .A2(A[21]), .ZN(n85) );
  NAND2_X1 U469 ( .A1(B[12]), .A2(A[12]), .ZN(n126) );
  NAND2_X1 U470 ( .A1(B[19]), .A2(A[19]), .ZN(n93) );
  NAND2_X1 U471 ( .A1(B[13]), .A2(A[13]), .ZN(n121) );
  NAND2_X1 U472 ( .A1(B[15]), .A2(A[15]), .ZN(n109) );
  NAND2_X1 U473 ( .A1(B[17]), .A2(A[17]), .ZN(n101) );
  NAND2_X1 U474 ( .A1(B[23]), .A2(A[23]), .ZN(n77) );
  NAND2_X1 U475 ( .A1(B[25]), .A2(A[25]), .ZN(n69) );
  NAND2_X1 U476 ( .A1(B[27]), .A2(A[27]), .ZN(n61) );
  NAND2_X1 U477 ( .A1(B[29]), .A2(A[29]), .ZN(n53) );
  NAND2_X1 U478 ( .A1(B[31]), .A2(A[31]), .ZN(n45) );
  NAND2_X1 U479 ( .A1(B[20]), .A2(A[20]), .ZN(n88) );
  NAND2_X1 U480 ( .A1(B[18]), .A2(A[18]), .ZN(n96) );
  NAND2_X1 U481 ( .A1(B[14]), .A2(A[14]), .ZN(n112) );
  NAND2_X1 U482 ( .A1(B[16]), .A2(A[16]), .ZN(n104) );
  NAND2_X1 U483 ( .A1(B[30]), .A2(A[30]), .ZN(n48) );
  NAND2_X1 U484 ( .A1(B[28]), .A2(A[28]), .ZN(n56) );
  NAND2_X1 U485 ( .A1(B[26]), .A2(A[26]), .ZN(n64) );
  NAND2_X1 U486 ( .A1(B[24]), .A2(A[24]), .ZN(n72) );
  NAND2_X1 U487 ( .A1(B[22]), .A2(A[22]), .ZN(n80) );
  OR2_X1 U488 ( .A1(B[21]), .A2(A[21]), .ZN(n400) );
  OR2_X1 U489 ( .A1(B[15]), .A2(A[15]), .ZN(n401) );
  OR2_X1 U490 ( .A1(B[23]), .A2(A[23]), .ZN(n402) );
  OR2_X1 U491 ( .A1(B[25]), .A2(A[25]), .ZN(n403) );
  OR2_X1 U492 ( .A1(B[27]), .A2(A[27]), .ZN(n404) );
  OR2_X1 U493 ( .A1(B[29]), .A2(A[29]), .ZN(n405) );
  OR2_X1 U494 ( .A1(B[31]), .A2(A[31]), .ZN(n406) );
  XNOR2_X1 U495 ( .A(n34), .B(n407), .ZN(SUM[39]) );
  XNOR2_X1 U496 ( .A(A[39]), .B(B[39]), .ZN(n407) );
  XNOR2_X1 U497 ( .A(n389), .B(n12), .ZN(SUM[21]) );
  OAI21_X1 U498 ( .B1(n89), .B2(n87), .A(n88), .ZN(n86) );
  XOR2_X1 U499 ( .A(n394), .B(n13), .Z(SUM[20]) );
  XNOR2_X1 U500 ( .A(n387), .B(n14), .ZN(SUM[19]) );
  XNOR2_X1 U501 ( .A(n377), .B(n6), .ZN(SUM[27]) );
  AOI21_X1 U502 ( .B1(n62), .B2(n404), .A(n59), .ZN(n57) );
  XOR2_X1 U503 ( .A(n384), .B(n5), .Z(SUM[28]) );
  XOR2_X1 U504 ( .A(n373), .B(n7), .Z(SUM[26]) );
  XOR2_X1 U505 ( .A(n390), .B(n15), .Z(SUM[18]) );
  OAI21_X1 U506 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  OAI21_X1 U507 ( .B1(n65), .B2(n63), .A(n64), .ZN(n62) );
  OAI21_X1 U508 ( .B1(n97), .B2(n95), .A(n96), .ZN(n94) );
  XNOR2_X1 U509 ( .A(n378), .B(n4), .ZN(SUM[29]) );
  XNOR2_X1 U510 ( .A(n360), .B(n8), .ZN(SUM[25]) );
  XNOR2_X1 U511 ( .A(n386), .B(n16), .ZN(SUM[17]) );
  AOI21_X1 U512 ( .B1(n54), .B2(n405), .A(n51), .ZN(n49) );
  XOR2_X1 U513 ( .A(n393), .B(n9), .Z(SUM[24]) );
  XOR2_X1 U514 ( .A(n372), .B(n17), .Z(SUM[16]) );
  OAI21_X1 U515 ( .B1(n73), .B2(n71), .A(n72), .ZN(n70) );
  AOI21_X1 U516 ( .B1(n78), .B2(n402), .A(n75), .ZN(n73) );
  OAI21_X1 U517 ( .B1(n105), .B2(n103), .A(n104), .ZN(n102) );
  XNOR2_X1 U518 ( .A(n379), .B(n10), .ZN(SUM[23]) );
  XNOR2_X1 U519 ( .A(n359), .B(n18), .ZN(SUM[15]) );
  INV_X1 U520 ( .A(n41), .ZN(n185) );
  XNOR2_X1 U521 ( .A(n388), .B(n2), .ZN(SUM[31]) );
  XOR2_X1 U522 ( .A(n391), .B(n19), .Z(SUM[14]) );
  XOR2_X1 U523 ( .A(n392), .B(n11), .Z(SUM[22]) );
  XOR2_X1 U524 ( .A(n385), .B(n3), .Z(SUM[30]) );
  AOI21_X1 U525 ( .B1(n46), .B2(n406), .A(n43), .ZN(n41) );
  OAI21_X1 U526 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  OAI21_X1 U527 ( .B1(n81), .B2(n79), .A(n80), .ZN(n78) );
  OAI21_X1 U528 ( .B1(n113), .B2(n111), .A(n112), .ZN(n110) );
endmodule


module mac_5 ( clk, clear_acc, a, b, mac_out );
  input [19:0] a;
  input [19:0] b;
  output [39:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, n3, n4;
  wire   [39:0] mul;
  wire   [39:0] pipeline;
  wire   [39:0] sum;

  DFF_X1 \pipeline_reg[38]  ( .D(mul[38]), .CK(clk), .Q(pipeline[38]) );
  DFF_X1 \pipeline_reg[37]  ( .D(mul[37]), .CK(clk), .Q(pipeline[37]) );
  DFF_X1 \pipeline_reg[36]  ( .D(mul[36]), .CK(clk), .Q(pipeline[36]) );
  DFF_X1 \pipeline_reg[35]  ( .D(mul[35]), .CK(clk), .Q(pipeline[35]) );
  DFF_X1 \pipeline_reg[34]  ( .D(mul[34]), .CK(clk), .Q(pipeline[34]) );
  DFF_X1 \pipeline_reg[33]  ( .D(mul[33]), .CK(clk), .Q(pipeline[33]) );
  DFF_X1 \pipeline_reg[32]  ( .D(mul[32]), .CK(clk), .Q(pipeline[32]) );
  DFF_X1 \pipeline_reg[31]  ( .D(mul[31]), .CK(clk), .Q(pipeline[31]) );
  DFF_X1 \pipeline_reg[30]  ( .D(mul[30]), .CK(clk), .Q(pipeline[30]) );
  DFF_X1 \pipeline_reg[29]  ( .D(mul[29]), .CK(clk), .Q(pipeline[29]) );
  DFF_X1 \pipeline_reg[28]  ( .D(mul[28]), .CK(clk), .Q(pipeline[28]) );
  DFF_X1 \pipeline_reg[27]  ( .D(mul[27]), .CK(clk), .Q(pipeline[27]) );
  DFF_X1 \pipeline_reg[26]  ( .D(mul[26]), .CK(clk), .Q(pipeline[26]) );
  DFF_X1 \pipeline_reg[25]  ( .D(mul[25]), .CK(clk), .Q(pipeline[25]) );
  DFF_X1 \pipeline_reg[24]  ( .D(mul[24]), .CK(clk), .Q(pipeline[24]) );
  DFF_X1 \pipeline_reg[23]  ( .D(mul[23]), .CK(clk), .Q(pipeline[23]) );
  DFF_X1 \pipeline_reg[22]  ( .D(mul[22]), .CK(clk), .Q(pipeline[22]) );
  DFF_X1 \pipeline_reg[21]  ( .D(mul[21]), .CK(clk), .Q(pipeline[21]) );
  DFF_X1 \pipeline_reg[20]  ( .D(mul[20]), .CK(clk), .Q(pipeline[20]) );
  DFF_X1 \pipeline_reg[19]  ( .D(mul[19]), .CK(clk), .Q(pipeline[19]) );
  DFF_X1 \pipeline_reg[18]  ( .D(mul[18]), .CK(clk), .Q(pipeline[18]) );
  DFF_X1 \pipeline_reg[17]  ( .D(mul[17]), .CK(clk), .Q(pipeline[17]) );
  DFF_X1 \pipeline_reg[16]  ( .D(mul[16]), .CK(clk), .Q(pipeline[16]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \mac_out_reg[16]  ( .D(N19), .CK(clk), .Q(mac_out[16]) );
  DFF_X1 \mac_out_reg[17]  ( .D(N20), .CK(clk), .Q(mac_out[17]) );
  DFF_X1 \mac_out_reg[18]  ( .D(N21), .CK(clk), .Q(mac_out[18]) );
  DFF_X1 \mac_out_reg[19]  ( .D(N22), .CK(clk), .Q(mac_out[19]) );
  DFF_X1 \mac_out_reg[20]  ( .D(N23), .CK(clk), .Q(mac_out[20]) );
  DFF_X1 \mac_out_reg[21]  ( .D(N24), .CK(clk), .Q(mac_out[21]) );
  DFF_X1 \mac_out_reg[22]  ( .D(N25), .CK(clk), .Q(mac_out[22]) );
  DFF_X1 \mac_out_reg[23]  ( .D(N26), .CK(clk), .Q(mac_out[23]) );
  DFF_X1 \mac_out_reg[24]  ( .D(N27), .CK(clk), .Q(mac_out[24]) );
  DFF_X1 \mac_out_reg[25]  ( .D(N28), .CK(clk), .Q(mac_out[25]) );
  DFF_X1 \mac_out_reg[26]  ( .D(N29), .CK(clk), .Q(mac_out[26]) );
  DFF_X1 \mac_out_reg[27]  ( .D(N30), .CK(clk), .Q(mac_out[27]) );
  DFF_X1 \mac_out_reg[28]  ( .D(N31), .CK(clk), .Q(mac_out[28]) );
  DFF_X1 \mac_out_reg[29]  ( .D(N32), .CK(clk), .Q(mac_out[29]) );
  DFF_X1 \mac_out_reg[30]  ( .D(N33), .CK(clk), .Q(mac_out[30]) );
  DFF_X1 \mac_out_reg[31]  ( .D(N34), .CK(clk), .Q(mac_out[31]) );
  DFF_X1 \mac_out_reg[32]  ( .D(N35), .CK(clk), .Q(mac_out[32]) );
  DFF_X1 \mac_out_reg[33]  ( .D(N36), .CK(clk), .Q(mac_out[33]) );
  DFF_X1 \mac_out_reg[34]  ( .D(N37), .CK(clk), .Q(mac_out[34]) );
  DFF_X1 \mac_out_reg[35]  ( .D(N38), .CK(clk), .Q(mac_out[35]) );
  DFF_X1 \mac_out_reg[36]  ( .D(N39), .CK(clk), .Q(mac_out[36]) );
  DFF_X1 \mac_out_reg[37]  ( .D(N40), .CK(clk), .Q(mac_out[37]) );
  DFF_X1 \mac_out_reg[38]  ( .D(N41), .CK(clk), .Q(mac_out[38]) );
  DFF_X1 \mac_out_reg[39]  ( .D(N42), .CK(clk), .Q(mac_out[39]) );
  mac_5_DW_mult_tc_1 mult_355 ( .a(a), .b(b), .product(mul) );
  mac_5_DW01_add_1 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  DFF_X2 \pipeline_reg[39]  ( .D(mul[39]), .CK(clk), .Q(pipeline[39]) );
  SDFF_X1 \mac_out_reg[11]  ( .D(1'b0), .SI(n4), .SE(sum[11]), .CK(clk), .Q(
        mac_out[11]) );
  BUF_X1 U4 ( .A(n4), .Z(n3) );
  INV_X1 U6 ( .A(clear_acc), .ZN(n4) );
  AND2_X1 U7 ( .A1(sum[39]), .A2(n3), .ZN(N42) );
  AND2_X1 U8 ( .A1(sum[38]), .A2(n3), .ZN(N41) );
  AND2_X1 U9 ( .A1(sum[37]), .A2(n3), .ZN(N40) );
  AND2_X1 U10 ( .A1(sum[36]), .A2(n3), .ZN(N39) );
  AND2_X1 U11 ( .A1(sum[35]), .A2(n3), .ZN(N38) );
  AND2_X1 U12 ( .A1(sum[34]), .A2(n3), .ZN(N37) );
  AND2_X1 U13 ( .A1(sum[33]), .A2(n3), .ZN(N36) );
  AND2_X1 U14 ( .A1(sum[32]), .A2(n3), .ZN(N35) );
  AND2_X1 U15 ( .A1(sum[31]), .A2(n3), .ZN(N34) );
  AND2_X1 U16 ( .A1(sum[30]), .A2(n3), .ZN(N33) );
  AND2_X1 U17 ( .A1(sum[29]), .A2(n3), .ZN(N32) );
  AND2_X1 U18 ( .A1(sum[28]), .A2(n4), .ZN(N31) );
  AND2_X1 U19 ( .A1(sum[27]), .A2(n4), .ZN(N30) );
  AND2_X1 U20 ( .A1(sum[26]), .A2(n4), .ZN(N29) );
  AND2_X1 U21 ( .A1(sum[25]), .A2(n4), .ZN(N28) );
  AND2_X1 U22 ( .A1(sum[24]), .A2(n4), .ZN(N27) );
  AND2_X1 U23 ( .A1(sum[23]), .A2(n4), .ZN(N26) );
  AND2_X1 U24 ( .A1(sum[22]), .A2(n4), .ZN(N25) );
  AND2_X1 U25 ( .A1(sum[21]), .A2(n4), .ZN(N24) );
  AND2_X1 U26 ( .A1(sum[20]), .A2(n4), .ZN(N23) );
  AND2_X1 U27 ( .A1(sum[19]), .A2(n4), .ZN(N22) );
  AND2_X1 U28 ( .A1(sum[18]), .A2(n4), .ZN(N21) );
  AND2_X1 U29 ( .A1(sum[17]), .A2(n4), .ZN(N20) );
  AND2_X1 U30 ( .A1(sum[16]), .A2(n4), .ZN(N19) );
  AND2_X1 U31 ( .A1(sum[15]), .A2(n4), .ZN(N18) );
  AND2_X1 U32 ( .A1(sum[14]), .A2(n4), .ZN(N17) );
  AND2_X1 U33 ( .A1(sum[13]), .A2(n4), .ZN(N16) );
  AND2_X1 U34 ( .A1(sum[12]), .A2(n4), .ZN(N15) );
  AND2_X1 U35 ( .A1(sum[10]), .A2(n4), .ZN(N13) );
  AND2_X1 U36 ( .A1(sum[9]), .A2(n4), .ZN(N12) );
  AND2_X1 U37 ( .A1(sum[8]), .A2(n4), .ZN(N11) );
  AND2_X1 U38 ( .A1(sum[7]), .A2(n4), .ZN(N10) );
  AND2_X1 U39 ( .A1(sum[6]), .A2(n4), .ZN(N9) );
  AND2_X1 U40 ( .A1(sum[5]), .A2(n4), .ZN(N8) );
  AND2_X1 U41 ( .A1(sum[4]), .A2(n4), .ZN(N7) );
  AND2_X1 U42 ( .A1(sum[3]), .A2(n4), .ZN(N6) );
  AND2_X1 U43 ( .A1(sum[2]), .A2(n4), .ZN(N5) );
  AND2_X1 U44 ( .A1(sum[1]), .A2(n4), .ZN(N4) );
  AND2_X1 U45 ( .A1(sum[0]), .A2(n3), .ZN(N3) );
endmodule


module mac_4_DW_mult_tc_1 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n4, n6, n7, n9, n12, n13, n16, n18, n19, n22, n24, n25, n28, n30,
         n31, n34, n36, n37, n40, n42, n43, n46, n48, n49, n52, n54, n55, n58,
         n60, n61, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n97, n98, n99, n100, n101, n103, n105,
         n106, n107, n108, n109, n111, n113, n114, n115, n116, n117, n119,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n183, n185, n186, n187, n188, n190, n193,
         n194, n195, n196, n198, n200, n201, n202, n203, n204, n205, n206,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n225, n227, n228, n230, n232, n233,
         n234, n236, n238, n239, n240, n241, n242, n244, n246, n247, n248,
         n249, n250, n252, n254, n255, n256, n257, n258, n259, n260, n261,
         n263, n264, n266, n268, n270, n271, n272, n273, n274, n275, n277,
         n278, n279, n280, n284, n285, n286, n287, n291, n293, n295, n296,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n643, n644, n646, n647, n649, n650, n652, n653, n655,
         n656, n658, n659, n661, n662, n664, n665, n667, n668, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1119, n1141, n1142,
         n1144, n1145, n1146, n1147, n1148, n1149, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n37 = a[13];
  assign n43 = a[15];
  assign n49 = a[17];
  assign n55 = a[19];
  assign n61 = b[0];
  assign n668 = a[0];
  assign n1090 = b[19];
  assign n1091 = b[18];
  assign n1092 = b[17];
  assign n1093 = b[16];
  assign n1094 = b[15];
  assign n1095 = b[14];
  assign n1096 = b[13];
  assign n1097 = b[12];
  assign n1098 = b[11];
  assign n1099 = b[10];
  assign n1100 = b[9];
  assign n1101 = b[8];
  assign n1102 = b[7];
  assign n1103 = b[6];
  assign n1104 = b[5];
  assign n1105 = b[4];
  assign n1106 = b[3];
  assign n1107 = b[2];
  assign n1108 = b[1];

  FA_X1 U333 ( .A(n681), .B(n304), .CI(n700), .CO(n300), .S(n301) );
  FA_X1 U334 ( .A(n305), .B(n682), .CI(n308), .CO(n302), .S(n303) );
  FA_X1 U336 ( .A(n312), .B(n683), .CI(n309), .CO(n306), .S(n307) );
  FA_X1 U337 ( .A(n701), .B(n314), .CI(n720), .CO(n308), .S(n309) );
  FA_X1 U338 ( .A(n313), .B(n320), .CI(n318), .CO(n310), .S(n311) );
  FA_X1 U339 ( .A(n684), .B(n702), .CI(n315), .CO(n312), .S(n313) );
  FA_X1 U341 ( .A(n324), .B(n321), .CI(n319), .CO(n316), .S(n317) );
  FA_X1 U342 ( .A(n328), .B(n721), .CI(n326), .CO(n318), .S(n319) );
  FA_X1 U343 ( .A(n703), .B(n685), .CI(n740), .CO(n320), .S(n321) );
  FA_X1 U344 ( .A(n325), .B(n327), .CI(n332), .CO(n322), .S(n323) );
  FA_X1 U345 ( .A(n336), .B(n329), .CI(n334), .CO(n324), .S(n325) );
  FA_X1 U346 ( .A(n686), .B(n704), .CI(n722), .CO(n326), .S(n327) );
  FA_X1 U348 ( .A(n340), .B(n342), .CI(n333), .CO(n330), .S(n331) );
  FA_X1 U349 ( .A(n335), .B(n344), .CI(n337), .CO(n332), .S(n333) );
  FA_X1 U350 ( .A(n705), .B(n346), .CI(n723), .CO(n334), .S(n335) );
  FA_X1 U351 ( .A(n741), .B(n687), .CI(n760), .CO(n336), .S(n337) );
  FA_X1 U352 ( .A(n350), .B(n343), .CI(n341), .CO(n338), .S(n339) );
  FA_X1 U353 ( .A(n345), .B(n354), .CI(n352), .CO(n340), .S(n341) );
  FA_X1 U354 ( .A(n347), .B(n724), .CI(n356), .CO(n342), .S(n343) );
  FA_X1 U355 ( .A(n742), .B(n706), .CI(n688), .CO(n344), .S(n345) );
  FA_X1 U357 ( .A(n360), .B(n353), .CI(n351), .CO(n348), .S(n349) );
  FA_X1 U358 ( .A(n357), .B(n355), .CI(n362), .CO(n350), .S(n351) );
  FA_X1 U359 ( .A(n366), .B(n743), .CI(n364), .CO(n352), .S(n353) );
  FA_X1 U360 ( .A(n707), .B(n761), .CI(n725), .CO(n354), .S(n355) );
  FA_X1 U361 ( .A(n368), .B(n689), .CI(n780), .CO(n356), .S(n357) );
  FA_X1 U362 ( .A(n372), .B(n363), .CI(n361), .CO(n358), .S(n359) );
  FA_X1 U363 ( .A(n376), .B(n365), .CI(n374), .CO(n360), .S(n361) );
  FA_X1 U364 ( .A(n378), .B(n380), .CI(n367), .CO(n362), .S(n363) );
  FA_X1 U365 ( .A(n690), .B(n708), .CI(n369), .CO(n364), .S(n365) );
  FA_X1 U366 ( .A(n762), .B(n726), .CI(n744), .CO(n366), .S(n367) );
  FA_X1 U368 ( .A(n384), .B(n375), .CI(n373), .CO(n370), .S(n371) );
  FA_X1 U369 ( .A(n377), .B(n388), .CI(n386), .CO(n372), .S(n373) );
  FA_X1 U370 ( .A(n379), .B(n390), .CI(n381), .CO(n374), .S(n375) );
  FA_X1 U371 ( .A(n727), .B(n745), .CI(n392), .CO(n376), .S(n377) );
  FA_X1 U372 ( .A(n709), .B(n781), .CI(n763), .CO(n378), .S(n379) );
  FA_X1 U373 ( .A(n394), .B(n691), .CI(n800), .CO(n380), .S(n381) );
  FA_X1 U374 ( .A(n398), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U375 ( .A(n389), .B(n402), .CI(n400), .CO(n384), .S(n385) );
  FA_X1 U376 ( .A(n391), .B(n404), .CI(n393), .CO(n386), .S(n387) );
  FA_X1 U377 ( .A(n408), .B(n395), .CI(n406), .CO(n388), .S(n389) );
  FA_X1 U378 ( .A(n746), .B(n782), .CI(n764), .CO(n390), .S(n391) );
  FA_X1 U379 ( .A(n692), .B(n728), .CI(n710), .CO(n392), .S(n393) );
  FA_X1 U381 ( .A(n412), .B(n401), .CI(n399), .CO(n396), .S(n397) );
  FA_X1 U382 ( .A(n403), .B(n416), .CI(n414), .CO(n398), .S(n399) );
  FA_X1 U383 ( .A(n409), .B(n407), .CI(n418), .CO(n400), .S(n401) );
  FA_X1 U384 ( .A(n420), .B(n422), .CI(n405), .CO(n402), .S(n403) );
  FA_X1 U385 ( .A(n765), .B(n747), .CI(n729), .CO(n404), .S(n405) );
  FA_X1 U386 ( .A(n711), .B(n801), .CI(n783), .CO(n406), .S(n407) );
  FA_X1 U387 ( .A(n424), .B(n693), .CI(n820), .CO(n408), .S(n409) );
  FA_X1 U388 ( .A(n428), .B(n415), .CI(n413), .CO(n410), .S(n411) );
  FA_X1 U389 ( .A(n417), .B(n432), .CI(n430), .CO(n412), .S(n413) );
  FA_X1 U391 ( .A(n436), .B(n438), .CI(n421), .CO(n416), .S(n417) );
  FA_X1 U393 ( .A(n694), .B(n766), .CI(n712), .CO(n420), .S(n421) );
  FA_X1 U394 ( .A(n802), .B(n730), .CI(n784), .CO(n422), .S(n423) );
  FA_X1 U399 ( .A(n437), .B(n452), .CI(n439), .CO(n432), .S(n433) );
  FA_X1 U400 ( .A(n456), .B(n767), .CI(n454), .CO(n434), .S(n435) );
  FA_X1 U401 ( .A(n731), .B(n785), .CI(n749), .CO(n436), .S(n437) );
  FA_X1 U402 ( .A(n458), .B(n803), .CI(n713), .CO(n438), .S(n439) );
  FA_X1 U406 ( .A(n468), .B(n453), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U407 ( .A(n455), .B(n470), .CI(n457), .CO(n448), .S(n449) );
  FA_X1 U408 ( .A(n472), .B(n476), .CI(n474), .CO(n450), .S(n451) );
  FA_X1 U409 ( .A(n768), .B(n786), .CI(n459), .CO(n452), .S(n453) );
  FA_X1 U410 ( .A(n714), .B(n732), .CI(n804), .CO(n454), .S(n455) );
  FA_X1 U416 ( .A(n473), .B(n488), .CI(n475), .CO(n466), .S(n467) );
  FA_X1 U417 ( .A(n492), .B(n490), .CI(n477), .CO(n468), .S(n469) );
  FA_X1 U418 ( .A(n805), .B(n823), .CI(n494), .CO(n470), .S(n471) );
  FA_X1 U419 ( .A(n733), .B(n751), .CI(n841), .CO(n472), .S(n473) );
  FA_X1 U420 ( .A(n769), .B(n860), .CI(n697), .CO(n474), .S(n475) );
  FA_X1 U425 ( .A(n504), .B(n493), .CI(n502), .CO(n482), .S(n483) );
  FA_X1 U426 ( .A(n489), .B(n506), .CI(n491), .CO(n484), .S(n485) );
  FA_X1 U427 ( .A(n510), .B(n495), .CI(n508), .CO(n486), .S(n487) );
  FA_X1 U428 ( .A(n770), .B(n842), .CI(n824), .CO(n488), .S(n489) );
  FA_X1 U429 ( .A(n806), .B(n752), .CI(n861), .CO(n490), .S(n491) );
  FA_X1 U430 ( .A(n670), .B(n788), .CI(n734), .CO(n492), .S(n493) );
  HA_X1 U431 ( .A(n698), .B(n716), .CO(n494), .S(n495) );
  FA_X1 U433 ( .A(n516), .B(n505), .CI(n503), .CO(n498), .S(n499) );
  FA_X1 U436 ( .A(n526), .B(n807), .CI(n524), .CO(n504), .S(n505) );
  FA_X1 U437 ( .A(n771), .B(n789), .CI(n825), .CO(n506), .S(n507) );
  FA_X1 U438 ( .A(n717), .B(n843), .CI(n753), .CO(n508), .S(n509) );
  FA_X1 U443 ( .A(n536), .B(n540), .CI(n538), .CO(n518), .S(n519) );
  FA_X1 U444 ( .A(n826), .B(n844), .CI(n527), .CO(n520), .S(n521) );
  FA_X1 U445 ( .A(n754), .B(n772), .CI(n808), .CO(n522), .S(n523) );
  FA_X1 U446 ( .A(n863), .B(n671), .CI(n790), .CO(n524), .S(n525) );
  HA_X1 U447 ( .A(n736), .B(n718), .CO(n526), .S(n527) );
  FA_X1 U450 ( .A(n537), .B(n541), .CI(n539), .CO(n532), .S(n533) );
  FA_X1 U451 ( .A(n552), .B(n554), .CI(n550), .CO(n534), .S(n535) );
  FA_X1 U452 ( .A(n791), .B(n827), .CI(n809), .CO(n536), .S(n537) );
  FA_X1 U453 ( .A(n773), .B(n845), .CI(n737), .CO(n538), .S(n539) );
  FA_X1 U454 ( .A(n755), .B(n719), .CI(n864), .CO(n540), .S(n541) );
  FA_X1 U455 ( .A(n547), .B(n558), .CI(n545), .CO(n542), .S(n543) );
  FA_X1 U456 ( .A(n560), .B(n553), .CI(n549), .CO(n544), .S(n545) );
  FA_X1 U457 ( .A(n562), .B(n564), .CI(n551), .CO(n546), .S(n547) );
  FA_X1 U458 ( .A(n555), .B(n846), .CI(n566), .CO(n548), .S(n549) );
  FA_X1 U459 ( .A(n865), .B(n792), .CI(n828), .CO(n550), .S(n551) );
  FA_X1 U460 ( .A(n774), .B(n810), .CI(n672), .CO(n552), .S(n553) );
  HA_X1 U461 ( .A(n738), .B(n756), .CO(n554), .S(n555) );
  FA_X1 U462 ( .A(n561), .B(n570), .CI(n559), .CO(n556), .S(n557) );
  FA_X1 U463 ( .A(n563), .B(n565), .CI(n572), .CO(n558), .S(n559) );
  FA_X1 U465 ( .A(n811), .B(n829), .CI(n578), .CO(n562), .S(n563) );
  FA_X1 U466 ( .A(n757), .B(n847), .CI(n793), .CO(n564), .S(n565) );
  FA_X1 U468 ( .A(n582), .B(n573), .CI(n571), .CO(n568), .S(n569) );
  FA_X1 U469 ( .A(n577), .B(n575), .CI(n584), .CO(n570), .S(n571) );
  FA_X1 U470 ( .A(n588), .B(n579), .CI(n586), .CO(n572), .S(n573) );
  FA_X1 U471 ( .A(n794), .B(n830), .CI(n848), .CO(n574), .S(n575) );
  FA_X1 U472 ( .A(n867), .B(n812), .CI(n673), .CO(n576), .S(n577) );
  HA_X1 U473 ( .A(n776), .B(n758), .CO(n578), .S(n579) );
  FA_X1 U474 ( .A(n585), .B(n592), .CI(n583), .CO(n580), .S(n581) );
  FA_X1 U475 ( .A(n587), .B(n589), .CI(n594), .CO(n582), .S(n583) );
  FA_X1 U476 ( .A(n1238), .B(n831), .CI(n596), .CO(n584), .S(n585) );
  FA_X1 U477 ( .A(n777), .B(n813), .CI(n849), .CO(n586), .S(n587) );
  FA_X1 U478 ( .A(n868), .B(n759), .CI(n795), .CO(n588), .S(n589) );
  FA_X1 U479 ( .A(n602), .B(n595), .CI(n593), .CO(n590), .S(n591) );
  FA_X1 U480 ( .A(n604), .B(n606), .CI(n597), .CO(n592), .S(n593) );
  FA_X1 U481 ( .A(n814), .B(n850), .CI(n599), .CO(n594), .S(n595) );
  FA_X1 U482 ( .A(n674), .B(n832), .CI(n869), .CO(n596), .S(n597) );
  FA_X1 U486 ( .A(n797), .B(n851), .CI(n833), .CO(n604), .S(n605) );
  FA_X1 U488 ( .A(n613), .B(n618), .CI(n611), .CO(n608), .S(n609) );
  FA_X1 U489 ( .A(n615), .B(n871), .CI(n620), .CO(n610), .S(n611) );
  FA_X1 U490 ( .A(n852), .B(n834), .CI(n675), .CO(n612), .S(n613) );
  HA_X1 U491 ( .A(n798), .B(n816), .CO(n614), .S(n615) );
  FA_X1 U492 ( .A(n621), .B(n624), .CI(n619), .CO(n616), .S(n617) );
  FA_X1 U493 ( .A(n817), .B(n853), .CI(n626), .CO(n618), .S(n619) );
  FA_X1 U494 ( .A(n835), .B(n799), .CI(n872), .CO(n620), .S(n621) );
  FA_X1 U495 ( .A(n630), .B(n627), .CI(n625), .CO(n622), .S(n623) );
  FA_X1 U496 ( .A(n854), .B(n873), .CI(n676), .CO(n624), .S(n625) );
  HA_X1 U497 ( .A(n818), .B(n836), .CO(n626), .S(n627) );
  FA_X1 U498 ( .A(n634), .B(n837), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U499 ( .A(n874), .B(n819), .CI(n855), .CO(n630), .S(n631) );
  FA_X1 U500 ( .A(n677), .B(n856), .CI(n635), .CO(n632), .S(n633) );
  HA_X1 U501 ( .A(n838), .B(n875), .CO(n634), .S(n635) );
  FA_X1 U502 ( .A(n876), .B(n839), .CI(n857), .CO(n636), .S(n637) );
  HA_X1 U503 ( .A(n858), .B(n877), .CO(n638), .S(n639) );
  BUF_X2 U1025 ( .A(n13), .Z(n1349) );
  BUF_X2 U1026 ( .A(n16), .Z(n1507) );
  XNOR2_X1 U1027 ( .A(n1233), .B(n485), .ZN(n481) );
  BUF_X1 U1028 ( .A(n55), .Z(n1344) );
  BUF_X2 U1029 ( .A(n24), .Z(n1457) );
  CLKBUF_X3 U1030 ( .A(n55), .Z(n1369) );
  BUF_X1 U1031 ( .A(n16), .Z(n1346) );
  XNOR2_X1 U1032 ( .A(n500), .B(n487), .ZN(n1233) );
  CLKBUF_X1 U1033 ( .A(n501), .Z(n1234) );
  BUF_X2 U1034 ( .A(n1105), .Z(n1370) );
  INV_X1 U1035 ( .A(n220), .ZN(n1235) );
  NAND2_X1 U1036 ( .A1(n840), .A2(n821), .ZN(n1253) );
  BUF_X1 U1037 ( .A(n1554), .Z(n1374) );
  BUF_X2 U1038 ( .A(n1100), .Z(n1380) );
  BUF_X2 U1039 ( .A(n1460), .Z(n1390) );
  BUF_X2 U1040 ( .A(n1553), .Z(n1358) );
  BUF_X2 U1041 ( .A(n1554), .Z(n1375) );
  BUF_X2 U1042 ( .A(n19), .Z(n1275) );
  XOR2_X1 U1043 ( .A(n1252), .B(n1260), .Z(n441) );
  BUF_X2 U1044 ( .A(n1096), .Z(n1563) );
  BUF_X2 U1045 ( .A(n40), .Z(n1322) );
  BUF_X2 U1046 ( .A(n1094), .Z(n1564) );
  BUF_X2 U1047 ( .A(n1091), .Z(n1566) );
  BUF_X2 U1048 ( .A(n1360), .Z(n1509) );
  NAND2_X1 U1049 ( .A1(n434), .A2(n423), .ZN(n1296) );
  AOI21_X1 U1050 ( .B1(n1503), .B2(n247), .A(n244), .ZN(n242) );
  BUF_X4 U1051 ( .A(n1104), .Z(n1556) );
  CLKBUF_X1 U1052 ( .A(n126), .Z(n1236) );
  CLKBUF_X1 U1053 ( .A(n431), .Z(n1237) );
  AND2_X1 U1054 ( .A1(n796), .A2(n778), .ZN(n1238) );
  BUF_X2 U1055 ( .A(n37), .Z(n1278) );
  BUF_X2 U1056 ( .A(n1092), .Z(n1565) );
  BUF_X2 U1057 ( .A(n1097), .Z(n1562) );
  OR2_X1 U1058 ( .A1(n1334), .A2(n442), .ZN(n1239) );
  OR2_X1 U1059 ( .A1(n679), .A2(n879), .ZN(n1240) );
  AND2_X1 U1060 ( .A1(n1240), .A2(n263), .ZN(product[1]) );
  XNOR2_X1 U1061 ( .A(n463), .B(n1242), .ZN(n461) );
  XNOR2_X1 U1062 ( .A(n480), .B(n465), .ZN(n1242) );
  NAND2_X1 U1063 ( .A1(n58), .A2(n1477), .ZN(n1243) );
  NAND2_X1 U1064 ( .A1(n58), .A2(n1477), .ZN(n60) );
  OAI22_X1 U1065 ( .A1(n1283), .A2(n1075), .B1(n1074), .B2(n4), .ZN(n1244) );
  BUF_X1 U1066 ( .A(n46), .Z(n1245) );
  XNOR2_X1 U1067 ( .A(n19), .B(a[8]), .ZN(n1246) );
  BUF_X2 U1068 ( .A(n1561), .Z(n1362) );
  AOI21_X1 U1069 ( .B1(n1486), .B2(n190), .A(n183), .ZN(n1247) );
  XOR2_X1 U1070 ( .A(n435), .B(n441), .Z(n1248) );
  XOR2_X1 U1071 ( .A(n450), .B(n1248), .Z(n431) );
  NAND2_X1 U1072 ( .A1(n450), .A2(n435), .ZN(n1249) );
  NAND2_X1 U1073 ( .A1(n450), .A2(n441), .ZN(n1250) );
  NAND2_X1 U1074 ( .A1(n435), .A2(n441), .ZN(n1251) );
  NAND3_X1 U1075 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n430) );
  XOR2_X1 U1076 ( .A(n840), .B(n821), .Z(n1252) );
  NAND2_X1 U1077 ( .A1(n840), .A2(n695), .ZN(n1254) );
  NAND2_X1 U1078 ( .A1(n821), .A2(n695), .ZN(n1255) );
  NAND3_X1 U1079 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n440) );
  XOR2_X1 U1080 ( .A(n425), .B(n748), .Z(n1256) );
  XOR2_X1 U1081 ( .A(n1256), .B(n440), .Z(n419) );
  NAND2_X1 U1082 ( .A1(n425), .A2(n748), .ZN(n1257) );
  NAND2_X1 U1083 ( .A1(n425), .A2(n440), .ZN(n1258) );
  NAND2_X1 U1084 ( .A1(n748), .A2(n440), .ZN(n1259) );
  NAND3_X1 U1085 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n418) );
  CLKBUF_X1 U1086 ( .A(n695), .Z(n1260) );
  CLKBUF_X1 U1087 ( .A(n1506), .Z(n1261) );
  CLKBUF_X3 U1088 ( .A(n34), .Z(n1506) );
  XNOR2_X1 U1089 ( .A(n1324), .B(n1545), .ZN(n1262) );
  CLKBUF_X3 U1090 ( .A(n13), .Z(n1350) );
  BUF_X1 U1091 ( .A(n9), .Z(n1360) );
  XOR2_X1 U1092 ( .A(n486), .B(n471), .Z(n1263) );
  XOR2_X1 U1093 ( .A(n469), .B(n1263), .Z(n465) );
  NAND2_X1 U1094 ( .A1(n469), .A2(n486), .ZN(n1264) );
  NAND2_X1 U1095 ( .A1(n469), .A2(n471), .ZN(n1265) );
  NAND2_X1 U1096 ( .A1(n486), .A2(n471), .ZN(n1266) );
  NAND3_X1 U1097 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n464) );
  CLKBUF_X2 U1098 ( .A(n1), .Z(n1270) );
  BUF_X2 U1099 ( .A(n1090), .Z(n1324) );
  BUF_X1 U1100 ( .A(n48), .Z(n1473) );
  OAI22_X1 U1101 ( .A1(n1408), .A2(n1030), .B1(n1029), .B2(n1346), .ZN(n1267)
         );
  INV_X1 U1102 ( .A(n644), .ZN(n1268) );
  CLKBUF_X3 U1103 ( .A(n52), .Z(n1335) );
  XNOR2_X1 U1104 ( .A(n1370), .B(n1386), .ZN(n1269) );
  CLKBUF_X1 U1105 ( .A(n1), .Z(n1545) );
  CLKBUF_X1 U1106 ( .A(n1105), .Z(n1371) );
  XOR2_X1 U1107 ( .A(n576), .B(n574), .Z(n1271) );
  XOR2_X1 U1108 ( .A(n567), .B(n1271), .Z(n561) );
  NAND2_X1 U1109 ( .A1(n567), .A2(n576), .ZN(n1272) );
  NAND2_X1 U1110 ( .A1(n567), .A2(n574), .ZN(n1273) );
  NAND2_X1 U1111 ( .A1(n576), .A2(n574), .ZN(n1274) );
  NAND3_X1 U1112 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(n560) );
  CLKBUF_X3 U1113 ( .A(n25), .Z(n1331) );
  BUF_X2 U1114 ( .A(n52), .Z(n1504) );
  BUF_X2 U1115 ( .A(n1100), .Z(n1381) );
  BUF_X1 U1116 ( .A(n1246), .Z(n1453) );
  CLKBUF_X1 U1117 ( .A(n19), .Z(n1547) );
  OAI22_X1 U1118 ( .A1(n1243), .A2(n897), .B1(n896), .B2(n1390), .ZN(n1276) );
  XNOR2_X1 U1119 ( .A(n1559), .B(n1407), .ZN(n1277) );
  CLKBUF_X1 U1120 ( .A(n37), .Z(n1407) );
  BUF_X2 U1121 ( .A(n18), .Z(n1279) );
  CLKBUF_X1 U1122 ( .A(n1348), .Z(n1280) );
  BUF_X2 U1123 ( .A(n6), .Z(n1348) );
  BUF_X2 U1124 ( .A(n6), .Z(n1347) );
  XOR2_X1 U1125 ( .A(n796), .B(n778), .Z(n599) );
  AOI21_X1 U1126 ( .B1(n1235), .B2(n213), .A(n214), .ZN(n1281) );
  CLKBUF_X1 U1127 ( .A(n1566), .Z(n1282) );
  BUF_X1 U1128 ( .A(n42), .Z(n1429) );
  NAND2_X1 U1129 ( .A1(n1119), .A2(n1385), .ZN(n1283) );
  CLKBUF_X1 U1130 ( .A(n1), .Z(n1284) );
  NAND2_X2 U1131 ( .A1(n1480), .A2(n1360), .ZN(n1469) );
  XOR2_X1 U1132 ( .A(n523), .B(n525), .Z(n1285) );
  XOR2_X1 U1133 ( .A(n534), .B(n1285), .Z(n517) );
  NAND2_X1 U1134 ( .A1(n534), .A2(n523), .ZN(n1286) );
  NAND2_X1 U1135 ( .A1(n534), .A2(n525), .ZN(n1287) );
  NAND2_X1 U1136 ( .A1(n523), .A2(n525), .ZN(n1288) );
  NAND3_X1 U1137 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n516) );
  CLKBUF_X1 U1138 ( .A(n530), .Z(n1289) );
  CLKBUF_X1 U1139 ( .A(n134), .Z(n1290) );
  CLKBUF_X2 U1140 ( .A(n1245), .Z(n1291) );
  BUF_X2 U1141 ( .A(n1245), .Z(n1292) );
  CLKBUF_X1 U1142 ( .A(n46), .Z(n1508) );
  XOR2_X1 U1143 ( .A(n434), .B(n423), .Z(n1293) );
  XOR2_X1 U1144 ( .A(n419), .B(n1293), .Z(n415) );
  NAND2_X1 U1145 ( .A1(n419), .A2(n434), .ZN(n1294) );
  NAND2_X1 U1146 ( .A1(n419), .A2(n423), .ZN(n1295) );
  NAND3_X1 U1147 ( .A1(n1294), .A2(n1295), .A3(n1296), .ZN(n414) );
  NOR2_X2 U1148 ( .A1(n581), .A2(n590), .ZN(n215) );
  NOR2_X2 U1149 ( .A1(n371), .A2(n382), .ZN(n135) );
  XNOR2_X1 U1150 ( .A(n1556), .B(n1388), .ZN(n1297) );
  CLKBUF_X1 U1151 ( .A(n176), .Z(n1298) );
  XOR2_X1 U1152 ( .A(n750), .B(n1267), .Z(n1299) );
  XOR2_X1 U1153 ( .A(n1276), .B(n1299), .Z(n457) );
  NAND2_X1 U1154 ( .A1(n1276), .A2(n750), .ZN(n1300) );
  NAND2_X1 U1155 ( .A1(n696), .A2(n822), .ZN(n1301) );
  NAND2_X1 U1156 ( .A1(n750), .A2(n822), .ZN(n1302) );
  NAND3_X1 U1157 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n456) );
  XNOR2_X1 U1158 ( .A(n1303), .B(n481), .ZN(n479) );
  XNOR2_X1 U1159 ( .A(n498), .B(n483), .ZN(n1303) );
  NAND2_X1 U1160 ( .A1(n500), .A2(n487), .ZN(n1304) );
  NAND2_X1 U1161 ( .A1(n500), .A2(n485), .ZN(n1305) );
  NAND2_X1 U1162 ( .A1(n487), .A2(n485), .ZN(n1306) );
  NAND3_X1 U1163 ( .A1(n1304), .A2(n1305), .A3(n1306), .ZN(n480) );
  NAND2_X1 U1164 ( .A1(n498), .A2(n483), .ZN(n1307) );
  NAND2_X1 U1165 ( .A1(n498), .A2(n481), .ZN(n1308) );
  NAND2_X1 U1166 ( .A1(n483), .A2(n481), .ZN(n1309) );
  NAND3_X1 U1167 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n478) );
  XOR2_X1 U1168 ( .A(n518), .B(n509), .Z(n1310) );
  XOR2_X1 U1169 ( .A(n520), .B(n1310), .Z(n501) );
  NAND2_X1 U1170 ( .A1(n520), .A2(n518), .ZN(n1311) );
  NAND2_X1 U1171 ( .A1(n520), .A2(n509), .ZN(n1312) );
  NAND2_X1 U1172 ( .A1(n518), .A2(n509), .ZN(n1313) );
  NAND3_X1 U1173 ( .A1(n1311), .A2(n1312), .A3(n1313), .ZN(n500) );
  XOR2_X1 U1174 ( .A(n467), .B(n484), .Z(n1314) );
  XOR2_X1 U1175 ( .A(n1314), .B(n482), .Z(n463) );
  NAND2_X1 U1176 ( .A1(n467), .A2(n484), .ZN(n1315) );
  NAND2_X1 U1177 ( .A1(n467), .A2(n482), .ZN(n1316) );
  NAND2_X1 U1178 ( .A1(n484), .A2(n482), .ZN(n1317) );
  NAND3_X1 U1179 ( .A1(n1315), .A2(n1316), .A3(n1317), .ZN(n462) );
  NAND2_X1 U1180 ( .A1(n480), .A2(n465), .ZN(n1318) );
  NAND2_X1 U1181 ( .A1(n480), .A2(n463), .ZN(n1319) );
  NAND2_X1 U1182 ( .A1(n465), .A2(n463), .ZN(n1320) );
  NAND3_X1 U1183 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n460) );
  NOR2_X1 U1184 ( .A1(n557), .A2(n568), .ZN(n1321) );
  NOR2_X1 U1185 ( .A1(n557), .A2(n568), .ZN(n204) );
  CLKBUF_X1 U1186 ( .A(n40), .Z(n1323) );
  BUF_X1 U1187 ( .A(n42), .Z(n1431) );
  NAND2_X1 U1188 ( .A1(n1484), .A2(n28), .ZN(n30) );
  BUF_X2 U1189 ( .A(n9), .Z(n1510) );
  XNOR2_X1 U1190 ( .A(n1325), .B(n464), .ZN(n445) );
  XNOR2_X1 U1191 ( .A(n449), .B(n466), .ZN(n1325) );
  BUF_X2 U1192 ( .A(n1101), .Z(n1559) );
  NAND2_X1 U1193 ( .A1(n1524), .A2(n302), .ZN(n1326) );
  NAND2_X1 U1194 ( .A1(n1440), .A2(n300), .ZN(n1327) );
  XNOR2_X1 U1195 ( .A(n1565), .B(n1350), .ZN(n1328) );
  BUF_X2 U1196 ( .A(n18), .Z(n1408) );
  XOR2_X1 U1197 ( .A(n1549), .B(a[16]), .Z(n1329) );
  BUF_X2 U1198 ( .A(n49), .Z(n1549) );
  XNOR2_X1 U1199 ( .A(n1330), .B(n446), .ZN(n429) );
  XNOR2_X1 U1200 ( .A(n433), .B(n448), .ZN(n1330) );
  CLKBUF_X3 U1201 ( .A(n25), .Z(n1332) );
  BUF_X1 U1202 ( .A(n1553), .Z(n1356) );
  NAND3_X1 U1203 ( .A1(n1411), .A2(n1412), .A3(n1413), .ZN(n1333) );
  XNOR2_X1 U1204 ( .A(n1409), .B(n429), .ZN(n1334) );
  NAND2_X1 U1205 ( .A1(n1480), .A2(n1360), .ZN(n1336) );
  CLKBUF_X1 U1206 ( .A(n1528), .Z(n1337) );
  NAND3_X1 U1207 ( .A1(n1327), .A2(n1448), .A3(n1446), .ZN(n1338) );
  CLKBUF_X1 U1208 ( .A(n1434), .Z(n1339) );
  CLKBUF_X1 U1209 ( .A(n1326), .Z(n1340) );
  CLKBUF_X1 U1210 ( .A(n1532), .Z(n1341) );
  INV_X1 U1211 ( .A(n1278), .ZN(n1342) );
  INV_X2 U1212 ( .A(n1342), .ZN(n1343) );
  CLKBUF_X1 U1213 ( .A(n1431), .Z(n1345) );
  NAND2_X1 U1214 ( .A1(n1480), .A2(n9), .ZN(n12) );
  NAND2_X1 U1215 ( .A1(n1119), .A2(n1385), .ZN(n6) );
  OAI22_X1 U1216 ( .A1(n1473), .A2(n938), .B1(n937), .B2(n1292), .ZN(n1351) );
  BUF_X1 U1217 ( .A(n1095), .Z(n1352) );
  BUF_X1 U1218 ( .A(n1095), .Z(n1353) );
  BUF_X2 U1219 ( .A(n42), .Z(n1430) );
  BUF_X1 U1220 ( .A(n61), .Z(n1354) );
  BUF_X1 U1221 ( .A(n61), .Z(n1355) );
  BUF_X1 U1222 ( .A(n1553), .Z(n1357) );
  BUF_X1 U1223 ( .A(n1246), .Z(n1359) );
  BUF_X1 U1224 ( .A(n1108), .Z(n1361) );
  CLKBUF_X1 U1225 ( .A(n1108), .Z(n1552) );
  BUF_X2 U1226 ( .A(n1561), .Z(n1363) );
  CLKBUF_X1 U1227 ( .A(n1561), .Z(n1364) );
  CLKBUF_X1 U1228 ( .A(n1103), .Z(n1365) );
  CLKBUF_X1 U1229 ( .A(n1103), .Z(n1366) );
  CLKBUF_X1 U1230 ( .A(n1103), .Z(n1557) );
  BUF_X1 U1231 ( .A(n1102), .Z(n1367) );
  BUF_X1 U1232 ( .A(n1102), .Z(n1368) );
  BUF_X1 U1233 ( .A(n1099), .Z(n1372) );
  BUF_X1 U1234 ( .A(n1099), .Z(n1373) );
  XNOR2_X1 U1235 ( .A(n1393), .B(a[18]), .ZN(n1477) );
  NAND2_X1 U1236 ( .A1(n1329), .A2(n1504), .ZN(n1376) );
  NAND2_X1 U1237 ( .A1(n1482), .A2(n1504), .ZN(n1377) );
  NAND2_X1 U1238 ( .A1(n1329), .A2(n1504), .ZN(n1410) );
  CLKBUF_X1 U1239 ( .A(n150), .Z(n1378) );
  AOI21_X1 U1240 ( .B1(n1455), .B2(n133), .A(n1290), .ZN(n1379) );
  BUF_X1 U1241 ( .A(n1093), .Z(n1382) );
  BUF_X1 U1242 ( .A(n1093), .Z(n1383) );
  CLKBUF_X1 U1243 ( .A(n1324), .Z(n1384) );
  INV_X1 U1244 ( .A(n668), .ZN(n1385) );
  INV_X2 U1245 ( .A(n668), .ZN(n4) );
  BUF_X4 U1246 ( .A(n49), .Z(n1386) );
  CLKBUF_X3 U1247 ( .A(n43), .Z(n1387) );
  CLKBUF_X3 U1248 ( .A(n43), .Z(n1388) );
  CLKBUF_X1 U1249 ( .A(n1529), .Z(n1389) );
  CLKBUF_X1 U1250 ( .A(n148), .Z(n1391) );
  CLKBUF_X1 U1251 ( .A(n1243), .Z(n1392) );
  INV_X1 U1252 ( .A(n55), .ZN(n1393) );
  XNOR2_X1 U1253 ( .A(n1394), .B(n862), .ZN(n511) );
  XNOR2_X1 U1254 ( .A(n735), .B(n699), .ZN(n1394) );
  XNOR2_X1 U1255 ( .A(n1395), .B(n445), .ZN(n443) );
  XNOR2_X1 U1256 ( .A(n462), .B(n447), .ZN(n1395) );
  XOR2_X1 U1257 ( .A(n522), .B(n507), .Z(n1396) );
  XOR2_X1 U1258 ( .A(n1396), .B(n511), .Z(n503) );
  NAND2_X1 U1259 ( .A1(n1351), .A2(n699), .ZN(n1397) );
  NAND2_X1 U1260 ( .A1(n1351), .A2(n862), .ZN(n1398) );
  NAND2_X1 U1261 ( .A1(n699), .A2(n862), .ZN(n1399) );
  NAND3_X1 U1262 ( .A1(n1397), .A2(n1398), .A3(n1399), .ZN(n510) );
  NAND2_X1 U1263 ( .A1(n522), .A2(n507), .ZN(n1400) );
  NAND2_X1 U1264 ( .A1(n522), .A2(n511), .ZN(n1401) );
  NAND2_X1 U1265 ( .A1(n511), .A2(n507), .ZN(n1402) );
  NAND3_X1 U1266 ( .A1(n1400), .A2(n1401), .A3(n1402), .ZN(n502) );
  XOR2_X1 U1267 ( .A(n501), .B(n514), .Z(n1403) );
  XOR2_X1 U1268 ( .A(n499), .B(n1403), .Z(n497) );
  NAND2_X1 U1269 ( .A1(n499), .A2(n1234), .ZN(n1404) );
  NAND2_X1 U1270 ( .A1(n499), .A2(n514), .ZN(n1405) );
  NAND2_X1 U1271 ( .A1(n1234), .A2(n514), .ZN(n1406) );
  NAND3_X1 U1272 ( .A1(n1404), .A2(n1405), .A3(n1406), .ZN(n496) );
  XNOR2_X1 U1273 ( .A(n1409), .B(n429), .ZN(n427) );
  XNOR2_X1 U1274 ( .A(n444), .B(n431), .ZN(n1409) );
  BUF_X2 U1275 ( .A(n36), .Z(n1466) );
  NAND2_X1 U1276 ( .A1(n1484), .A2(n28), .ZN(n1435) );
  NAND2_X1 U1277 ( .A1(n1482), .A2(n1504), .ZN(n54) );
  NAND2_X1 U1278 ( .A1(n449), .A2(n466), .ZN(n1411) );
  NAND2_X1 U1279 ( .A1(n449), .A2(n464), .ZN(n1412) );
  NAND2_X1 U1280 ( .A1(n466), .A2(n464), .ZN(n1413) );
  NAND3_X1 U1281 ( .A1(n1411), .A2(n1412), .A3(n1413), .ZN(n444) );
  NAND2_X1 U1282 ( .A1(n462), .A2(n447), .ZN(n1414) );
  NAND2_X1 U1283 ( .A1(n462), .A2(n445), .ZN(n1415) );
  NAND2_X1 U1284 ( .A1(n447), .A2(n445), .ZN(n1416) );
  NAND3_X1 U1285 ( .A1(n1414), .A2(n1415), .A3(n1416), .ZN(n442) );
  INV_X1 U1286 ( .A(n277), .ZN(n1417) );
  NOR2_X1 U1287 ( .A1(n443), .A2(n460), .ZN(n161) );
  CLKBUF_X1 U1288 ( .A(n159), .Z(n1418) );
  XNOR2_X1 U1289 ( .A(n1419), .B(n1443), .ZN(product[38]) );
  XNOR2_X1 U1290 ( .A(n680), .B(n298), .ZN(n1419) );
  NOR2_X1 U1291 ( .A1(n497), .A2(n512), .ZN(n1420) );
  NOR2_X1 U1292 ( .A1(n497), .A2(n512), .ZN(n177) );
  AND3_X1 U1293 ( .A1(n1451), .A2(n1450), .A3(n1449), .ZN(product[39]) );
  BUF_X2 U1294 ( .A(n36), .Z(n1467) );
  NAND2_X1 U1295 ( .A1(n433), .A2(n448), .ZN(n1422) );
  NAND2_X1 U1296 ( .A1(n433), .A2(n446), .ZN(n1423) );
  NAND2_X1 U1297 ( .A1(n448), .A2(n446), .ZN(n1424) );
  NAND3_X1 U1298 ( .A1(n1422), .A2(n1423), .A3(n1424), .ZN(n428) );
  NAND2_X1 U1299 ( .A1(n1333), .A2(n1237), .ZN(n1425) );
  NAND2_X1 U1300 ( .A1(n429), .A2(n1333), .ZN(n1426) );
  NAND2_X1 U1301 ( .A1(n1237), .A2(n429), .ZN(n1427) );
  NAND3_X1 U1302 ( .A1(n1425), .A2(n1426), .A3(n1427), .ZN(n426) );
  CLKBUF_X1 U1303 ( .A(n194), .Z(n1428) );
  NAND2_X1 U1304 ( .A1(n40), .A2(n1481), .ZN(n42) );
  CLKBUF_X1 U1305 ( .A(n58), .Z(n1432) );
  CLKBUF_X1 U1306 ( .A(n264), .Z(n1433) );
  NAND3_X1 U1307 ( .A1(n1437), .A2(n1438), .A3(n1439), .ZN(n1434) );
  XOR2_X1 U1308 ( .A(n310), .B(n307), .Z(n1436) );
  XOR2_X1 U1309 ( .A(n1433), .B(n1436), .Z(product[34]) );
  NAND2_X1 U1310 ( .A1(n264), .A2(n310), .ZN(n1437) );
  NAND2_X1 U1311 ( .A1(n264), .A2(n307), .ZN(n1438) );
  NAND2_X1 U1312 ( .A1(n310), .A2(n307), .ZN(n1439) );
  NAND3_X1 U1313 ( .A1(n1438), .A2(n1437), .A3(n1439), .ZN(n100) );
  NAND3_X1 U1314 ( .A1(n1532), .A2(n1326), .A3(n1530), .ZN(n1440) );
  NAND3_X1 U1315 ( .A1(n1341), .A2(n1340), .A3(n1530), .ZN(n1441) );
  CLKBUF_X1 U1316 ( .A(n114), .Z(n1442) );
  NAND3_X1 U1317 ( .A1(n1327), .A2(n1446), .A3(n1448), .ZN(n1443) );
  AOI21_X1 U1318 ( .B1(n1442), .B2(n1491), .A(n111), .ZN(n1444) );
  NAND2_X1 U1319 ( .A1(n1479), .A2(n16), .ZN(n18) );
  XOR2_X1 U1320 ( .A(n300), .B(n299), .Z(n1445) );
  XOR2_X1 U1321 ( .A(n1445), .B(n1441), .Z(product[37]) );
  NAND2_X1 U1322 ( .A1(n300), .A2(n299), .ZN(n1446) );
  NAND2_X1 U1323 ( .A1(n1440), .A2(n300), .ZN(n1447) );
  NAND2_X1 U1324 ( .A1(n299), .A2(n98), .ZN(n1448) );
  NAND3_X1 U1325 ( .A1(n1448), .A2(n1447), .A3(n1446), .ZN(n97) );
  NAND2_X1 U1326 ( .A1(n680), .A2(n298), .ZN(n1449) );
  NAND2_X1 U1327 ( .A1(n97), .A2(n680), .ZN(n1450) );
  NAND2_X1 U1328 ( .A1(n1338), .A2(n298), .ZN(n1451) );
  CLKBUF_X1 U1329 ( .A(n1246), .Z(n1452) );
  CLKBUF_X1 U1330 ( .A(n151), .Z(n1454) );
  CLKBUF_X1 U1331 ( .A(n146), .Z(n1455) );
  BUF_X2 U1332 ( .A(n24), .Z(n1456) );
  NAND2_X1 U1333 ( .A1(n22), .A2(n1483), .ZN(n24) );
  BUF_X2 U1334 ( .A(n48), .Z(n1472) );
  CLKBUF_X1 U1335 ( .A(n127), .Z(n1458) );
  AOI21_X1 U1336 ( .B1(n1462), .B2(n1236), .A(n1458), .ZN(n1459) );
  XNOR2_X1 U1337 ( .A(n1549), .B(a[18]), .ZN(n1460) );
  CLKBUF_X1 U1338 ( .A(n1392), .Z(n1461) );
  CLKBUF_X1 U1339 ( .A(n153), .Z(n1462) );
  CLKBUF_X1 U1340 ( .A(n106), .Z(n1463) );
  AOI21_X1 U1341 ( .B1(n175), .B2(n1428), .A(n1298), .ZN(n1464) );
  NOR2_X1 U1342 ( .A1(n461), .A2(n478), .ZN(n1465) );
  NAND2_X1 U1343 ( .A1(n1478), .A2(n34), .ZN(n36) );
  NOR2_X1 U1344 ( .A1(n397), .A2(n410), .ZN(n1468) );
  CLKBUF_X1 U1345 ( .A(n122), .Z(n1470) );
  CLKBUF_X1 U1346 ( .A(n48), .Z(n1471) );
  NAND2_X1 U1347 ( .A1(n1476), .A2(n46), .ZN(n48) );
  AOI21_X1 U1348 ( .B1(n122), .B2(n1490), .A(n119), .ZN(n1474) );
  NOR2_X1 U1349 ( .A1(n442), .A2(n427), .ZN(n1475) );
  NOR2_X1 U1350 ( .A1(n359), .A2(n370), .ZN(n128) );
  OR2_X1 U1351 ( .A1(n339), .A2(n348), .ZN(n1490) );
  BUF_X4 U1352 ( .A(n22), .Z(n1505) );
  XOR2_X1 U1353 ( .A(n43), .B(a[14]), .Z(n1476) );
  XOR2_X1 U1354 ( .A(n31), .B(a[10]), .Z(n1478) );
  XOR2_X1 U1355 ( .A(n13), .B(a[4]), .Z(n1479) );
  XOR2_X1 U1356 ( .A(n7), .B(a[2]), .Z(n1480) );
  BUF_X1 U1357 ( .A(n61), .Z(n1550) );
  BUF_X1 U1358 ( .A(n61), .Z(n1551) );
  XOR2_X1 U1359 ( .A(n37), .B(a[12]), .Z(n1481) );
  XOR2_X1 U1360 ( .A(n1549), .B(a[16]), .Z(n1482) );
  XOR2_X1 U1361 ( .A(n19), .B(a[6]), .Z(n1483) );
  XOR2_X1 U1362 ( .A(n25), .B(a[8]), .Z(n1484) );
  OAI21_X1 U1363 ( .B1(n152), .B2(n143), .A(n144), .ZN(n142) );
  XNOR2_X1 U1364 ( .A(n130), .B(n69), .ZN(product[27]) );
  NAND2_X1 U1365 ( .A1(n271), .A2(n129), .ZN(n69) );
  INV_X1 U1366 ( .A(n128), .ZN(n271) );
  INV_X1 U1367 ( .A(n200), .ZN(n198) );
  AOI21_X1 U1368 ( .B1(n1486), .B2(n190), .A(n183), .ZN(n181) );
  INV_X1 U1369 ( .A(n185), .ZN(n183) );
  INV_X1 U1370 ( .A(n188), .ZN(n190) );
  INV_X1 U1371 ( .A(n140), .ZN(n273) );
  XOR2_X1 U1372 ( .A(n168), .B(n76), .Z(product[20]) );
  NAND2_X1 U1373 ( .A1(n278), .A2(n167), .ZN(n76) );
  AOI21_X1 U1374 ( .B1(n173), .B2(n279), .A(n170), .ZN(n168) );
  XOR2_X1 U1375 ( .A(n137), .B(n70), .Z(product[26]) );
  NAND2_X1 U1376 ( .A1(n272), .A2(n136), .ZN(n70) );
  AOI21_X1 U1377 ( .B1(n142), .B2(n273), .A(n139), .ZN(n137) );
  XOR2_X1 U1378 ( .A(n206), .B(n82), .Z(product[14]) );
  NAND2_X1 U1379 ( .A1(n284), .A2(n205), .ZN(n82) );
  AOI21_X1 U1380 ( .B1(n211), .B2(n285), .A(n208), .ZN(n206) );
  XOR2_X1 U1381 ( .A(n163), .B(n75), .Z(product[21]) );
  NAND2_X1 U1382 ( .A1(n277), .A2(n162), .ZN(n75) );
  INV_X1 U1383 ( .A(n161), .ZN(n277) );
  XOR2_X1 U1384 ( .A(n193), .B(n80), .Z(product[16]) );
  NAND2_X1 U1385 ( .A1(n1523), .A2(n188), .ZN(n80) );
  XOR2_X1 U1386 ( .A(n201), .B(n81), .Z(product[15]) );
  XOR2_X1 U1387 ( .A(n152), .B(n73), .Z(product[23]) );
  INV_X1 U1388 ( .A(n1378), .ZN(n275) );
  NAND2_X1 U1389 ( .A1(n1486), .A2(n1523), .ZN(n180) );
  XNOR2_X1 U1390 ( .A(n160), .B(n74), .ZN(product[22]) );
  NAND2_X1 U1391 ( .A1(n1239), .A2(n1418), .ZN(n74) );
  OAI21_X1 U1392 ( .B1(n163), .B2(n1417), .A(n162), .ZN(n160) );
  XNOR2_X1 U1393 ( .A(n149), .B(n72), .ZN(product[24]) );
  NAND2_X1 U1394 ( .A1(n274), .A2(n1391), .ZN(n72) );
  INV_X1 U1395 ( .A(n1468), .ZN(n274) );
  XNOR2_X1 U1396 ( .A(n142), .B(n71), .ZN(product[25]) );
  NAND2_X1 U1397 ( .A1(n273), .A2(n141), .ZN(n71) );
  XNOR2_X1 U1398 ( .A(n186), .B(n79), .ZN(product[17]) );
  INV_X1 U1399 ( .A(n1523), .ZN(n187) );
  INV_X1 U1400 ( .A(n141), .ZN(n139) );
  INV_X1 U1401 ( .A(n121), .ZN(n119) );
  INV_X1 U1402 ( .A(n113), .ZN(n111) );
  NOR2_X1 U1403 ( .A1(n1420), .A2(n180), .ZN(n175) );
  INV_X1 U1404 ( .A(n238), .ZN(n236) );
  INV_X1 U1405 ( .A(n227), .ZN(n225) );
  NOR2_X1 U1406 ( .A1(n397), .A2(n410), .ZN(n147) );
  NOR2_X1 U1407 ( .A1(n411), .A2(n426), .ZN(n150) );
  OR2_X1 U1408 ( .A1(n543), .A2(n556), .ZN(n1485) );
  NAND2_X1 U1409 ( .A1(n443), .A2(n460), .ZN(n162) );
  OR2_X1 U1410 ( .A1(n529), .A2(n542), .ZN(n1523) );
  NOR2_X1 U1411 ( .A1(n461), .A2(n478), .ZN(n166) );
  NOR2_X1 U1412 ( .A1(n1334), .A2(n442), .ZN(n158) );
  NAND2_X1 U1413 ( .A1(n268), .A2(n116), .ZN(n66) );
  INV_X1 U1414 ( .A(n115), .ZN(n268) );
  NAND2_X1 U1415 ( .A1(n266), .A2(n108), .ZN(n64) );
  INV_X1 U1416 ( .A(n107), .ZN(n266) );
  NAND2_X1 U1417 ( .A1(n270), .A2(n124), .ZN(n68) );
  INV_X1 U1418 ( .A(n123), .ZN(n270) );
  NAND2_X1 U1419 ( .A1(n529), .A2(n542), .ZN(n188) );
  INV_X1 U1420 ( .A(n209), .ZN(n285) );
  INV_X1 U1421 ( .A(n171), .ZN(n279) );
  NAND2_X1 U1422 ( .A1(n1490), .A2(n121), .ZN(n67) );
  NAND2_X1 U1423 ( .A1(n1491), .A2(n113), .ZN(n65) );
  NAND2_X1 U1424 ( .A1(n1493), .A2(n105), .ZN(n63) );
  NAND2_X1 U1425 ( .A1(n1492), .A2(n238), .ZN(n88) );
  XOR2_X1 U1426 ( .A(n228), .B(n86), .Z(product[10]) );
  AOI21_X1 U1427 ( .B1(n233), .B2(n1489), .A(n230), .ZN(n228) );
  XOR2_X1 U1428 ( .A(n220), .B(n85), .Z(product[11]) );
  NAND2_X1 U1429 ( .A1(n287), .A2(n219), .ZN(n85) );
  INV_X1 U1430 ( .A(n218), .ZN(n287) );
  OR2_X1 U1431 ( .A1(n513), .A2(n528), .ZN(n1486) );
  NAND2_X1 U1432 ( .A1(n557), .A2(n568), .ZN(n205) );
  XNOR2_X1 U1433 ( .A(n211), .B(n83), .ZN(product[13]) );
  NAND2_X1 U1434 ( .A1(n285), .A2(n210), .ZN(n83) );
  XNOR2_X1 U1435 ( .A(n173), .B(n77), .ZN(product[19]) );
  NAND2_X1 U1436 ( .A1(n279), .A2(n172), .ZN(n77) );
  XNOR2_X1 U1437 ( .A(n233), .B(n87), .ZN(product[9]) );
  NAND2_X1 U1438 ( .A1(n1489), .A2(n232), .ZN(n87) );
  XNOR2_X1 U1439 ( .A(n179), .B(n78), .ZN(product[18]) );
  NAND2_X1 U1440 ( .A1(n280), .A2(n178), .ZN(n78) );
  INV_X1 U1441 ( .A(n1420), .ZN(n280) );
  XNOR2_X1 U1442 ( .A(n217), .B(n84), .ZN(product[12]) );
  NAND2_X1 U1443 ( .A1(n286), .A2(n216), .ZN(n84) );
  OAI21_X1 U1444 ( .B1(n220), .B2(n218), .A(n219), .ZN(n217) );
  NAND2_X1 U1445 ( .A1(n359), .A2(n370), .ZN(n129) );
  INV_X1 U1446 ( .A(n232), .ZN(n230) );
  INV_X1 U1447 ( .A(n210), .ZN(n208) );
  INV_X1 U1448 ( .A(n172), .ZN(n170) );
  NAND2_X1 U1449 ( .A1(n543), .A2(n556), .ZN(n200) );
  INV_X1 U1450 ( .A(n246), .ZN(n244) );
  XNOR2_X1 U1451 ( .A(n1487), .B(n515), .ZN(n513) );
  XNOR2_X1 U1452 ( .A(n517), .B(n530), .ZN(n1487) );
  XNOR2_X1 U1453 ( .A(n531), .B(n1488), .ZN(n529) );
  XNOR2_X1 U1454 ( .A(n544), .B(n533), .ZN(n1488) );
  OAI21_X1 U1455 ( .B1(n256), .B2(n258), .A(n257), .ZN(n255) );
  NAND3_X1 U1456 ( .A1(n1542), .A2(n1543), .A3(n1544), .ZN(n512) );
  NOR2_X1 U1457 ( .A1(n591), .A2(n600), .ZN(n218) );
  AOI21_X1 U1458 ( .B1(n1502), .B2(n255), .A(n252), .ZN(n250) );
  INV_X1 U1459 ( .A(n254), .ZN(n252) );
  OAI21_X1 U1460 ( .B1(n242), .B2(n240), .A(n241), .ZN(n239) );
  OR2_X1 U1461 ( .A1(n609), .A2(n616), .ZN(n1489) );
  XOR2_X1 U1462 ( .A(n91), .B(n250), .Z(product[5]) );
  NAND2_X1 U1463 ( .A1(n293), .A2(n249), .ZN(n91) );
  INV_X1 U1464 ( .A(n248), .ZN(n293) );
  XOR2_X1 U1465 ( .A(n242), .B(n89), .Z(product[7]) );
  NAND2_X1 U1466 ( .A1(n291), .A2(n241), .ZN(n89) );
  INV_X1 U1467 ( .A(n240), .ZN(n291) );
  NOR2_X1 U1468 ( .A1(n479), .A2(n496), .ZN(n171) );
  NOR2_X1 U1469 ( .A1(n569), .A2(n580), .ZN(n209) );
  NOR2_X1 U1470 ( .A1(n349), .A2(n358), .ZN(n123) );
  NOR2_X1 U1471 ( .A1(n317), .A2(n322), .ZN(n107) );
  NOR2_X1 U1472 ( .A1(n331), .A2(n338), .ZN(n115) );
  XNOR2_X1 U1473 ( .A(n90), .B(n247), .ZN(product[6]) );
  NAND2_X1 U1474 ( .A1(n1503), .A2(n246), .ZN(n90) );
  NAND2_X1 U1475 ( .A1(n591), .A2(n600), .ZN(n219) );
  INV_X1 U1476 ( .A(n259), .ZN(n258) );
  OAI21_X1 U1477 ( .B1(n260), .B2(n263), .A(n261), .ZN(n259) );
  NAND2_X1 U1478 ( .A1(n479), .A2(n496), .ZN(n172) );
  NAND2_X1 U1479 ( .A1(n569), .A2(n580), .ZN(n210) );
  XNOR2_X1 U1480 ( .A(n92), .B(n255), .ZN(product[4]) );
  NAND2_X1 U1481 ( .A1(n1502), .A2(n254), .ZN(n92) );
  NAND2_X1 U1482 ( .A1(n339), .A2(n348), .ZN(n121) );
  NAND2_X1 U1483 ( .A1(n323), .A2(n330), .ZN(n113) );
  NAND2_X1 U1484 ( .A1(n609), .A2(n616), .ZN(n232) );
  NAND2_X1 U1485 ( .A1(n617), .A2(n622), .ZN(n238) );
  NAND2_X1 U1486 ( .A1(n311), .A2(n316), .ZN(n105) );
  NAND2_X1 U1487 ( .A1(n317), .A2(n322), .ZN(n108) );
  NAND2_X1 U1488 ( .A1(n349), .A2(n358), .ZN(n124) );
  NAND2_X1 U1489 ( .A1(n331), .A2(n338), .ZN(n116) );
  NAND2_X1 U1490 ( .A1(n497), .A2(n512), .ZN(n178) );
  OR2_X1 U1491 ( .A1(n323), .A2(n330), .ZN(n1491) );
  OR2_X1 U1492 ( .A1(n617), .A2(n622), .ZN(n1492) );
  OR2_X1 U1493 ( .A1(n311), .A2(n316), .ZN(n1493) );
  NAND2_X1 U1494 ( .A1(n581), .A2(n590), .ZN(n216) );
  XOR2_X1 U1495 ( .A(n93), .B(n258), .Z(product[3]) );
  NAND2_X1 U1496 ( .A1(n295), .A2(n257), .ZN(n93) );
  INV_X1 U1497 ( .A(n256), .ZN(n295) );
  OR2_X1 U1498 ( .A1(n601), .A2(n608), .ZN(n1494) );
  XOR2_X1 U1499 ( .A(n94), .B(n263), .Z(product[2]) );
  NAND2_X1 U1500 ( .A1(n296), .A2(n261), .ZN(n94) );
  INV_X1 U1501 ( .A(n260), .ZN(n296) );
  XNOR2_X1 U1502 ( .A(n1495), .B(n603), .ZN(n601) );
  XNOR2_X1 U1503 ( .A(n610), .B(n605), .ZN(n1495) );
  XNOR2_X1 U1504 ( .A(n1496), .B(n607), .ZN(n603) );
  XNOR2_X1 U1505 ( .A(n612), .B(n614), .ZN(n1496) );
  XNOR2_X1 U1506 ( .A(n1497), .B(n519), .ZN(n515) );
  XNOR2_X1 U1507 ( .A(n532), .B(n521), .ZN(n1497) );
  XNOR2_X1 U1508 ( .A(n1498), .B(n535), .ZN(n531) );
  XNOR2_X1 U1509 ( .A(n546), .B(n548), .ZN(n1498) );
  XNOR2_X1 U1510 ( .A(n815), .B(n1499), .ZN(n607) );
  XNOR2_X1 U1511 ( .A(n870), .B(n779), .ZN(n1499) );
  XNOR2_X1 U1512 ( .A(n775), .B(n1500), .ZN(n567) );
  XNOR2_X1 U1513 ( .A(n1244), .B(n739), .ZN(n1500) );
  NAND3_X1 U1514 ( .A1(n1517), .A2(n1518), .A3(n1519), .ZN(n600) );
  NAND2_X1 U1515 ( .A1(n639), .A2(n678), .ZN(n257) );
  INV_X1 U1516 ( .A(n105), .ZN(n103) );
  NOR2_X1 U1517 ( .A1(n639), .A2(n678), .ZN(n256) );
  NOR2_X1 U1518 ( .A1(n878), .A2(n859), .ZN(n260) );
  XNOR2_X1 U1519 ( .A(n1501), .B(n1525), .ZN(product[36]) );
  XNOR2_X1 U1520 ( .A(n302), .B(n301), .ZN(n1501) );
  NAND2_X1 U1521 ( .A1(n679), .A2(n879), .ZN(n263) );
  NAND2_X1 U1522 ( .A1(n878), .A2(n859), .ZN(n261) );
  NOR2_X1 U1523 ( .A1(n623), .A2(n628), .ZN(n240) );
  OR2_X1 U1524 ( .A1(n637), .A2(n638), .ZN(n1502) );
  INV_X1 U1525 ( .A(n328), .ZN(n329) );
  INV_X1 U1526 ( .A(n394), .ZN(n395) );
  NOR2_X1 U1527 ( .A1(n633), .A2(n636), .ZN(n248) );
  INV_X1 U1528 ( .A(n298), .ZN(n299) );
  NAND2_X1 U1529 ( .A1(n629), .A2(n632), .ZN(n246) );
  NAND2_X1 U1530 ( .A1(n623), .A2(n628), .ZN(n241) );
  OR2_X1 U1531 ( .A1(n629), .A2(n632), .ZN(n1503) );
  NAND2_X1 U1532 ( .A1(n633), .A2(n636), .ZN(n249) );
  OR2_X1 U1533 ( .A1(n1354), .A2(n1148), .ZN(n1068) );
  OAI22_X1 U1534 ( .A1(n1347), .A2(n1086), .B1(n1085), .B2(n4), .ZN(n877) );
  OAI22_X1 U1535 ( .A1(n1348), .A2(n1088), .B1(n1087), .B2(n4), .ZN(n879) );
  OAI22_X1 U1536 ( .A1(n1347), .A2(n1149), .B1(n1089), .B2(n4), .ZN(n679) );
  OR2_X1 U1537 ( .A1(n1355), .A2(n1149), .ZN(n1089) );
  OAI22_X1 U1538 ( .A1(n1347), .A2(n1087), .B1(n1086), .B2(n4), .ZN(n878) );
  OAI22_X1 U1539 ( .A1(n1280), .A2(n1082), .B1(n1081), .B2(n4), .ZN(n873) );
  OAI22_X1 U1540 ( .A1(n1347), .A2(n1078), .B1(n1077), .B2(n4), .ZN(n869) );
  INV_X1 U1541 ( .A(n661), .ZN(n820) );
  OAI22_X1 U1542 ( .A1(n1347), .A2(n1084), .B1(n1083), .B2(n4), .ZN(n875) );
  OAI22_X1 U1543 ( .A1(n1262), .A2(n1283), .B1(n1069), .B2(n4), .ZN(n667) );
  OR2_X1 U1544 ( .A1(n1355), .A2(n1147), .ZN(n1047) );
  XNOR2_X1 U1545 ( .A(n1354), .B(n1386), .ZN(n920) );
  AND2_X1 U1546 ( .A1(n1551), .A2(n662), .ZN(n839) );
  OAI22_X1 U1547 ( .A1(n1348), .A2(n1085), .B1(n1084), .B2(n4), .ZN(n876) );
  XNOR2_X1 U1548 ( .A(n1384), .B(n1386), .ZN(n901) );
  INV_X1 U1549 ( .A(n643), .ZN(n700) );
  INV_X1 U1550 ( .A(n304), .ZN(n305) );
  XNOR2_X1 U1551 ( .A(n1353), .B(n1386), .ZN(n906) );
  XNOR2_X1 U1552 ( .A(n1563), .B(n1386), .ZN(n907) );
  XNOR2_X1 U1553 ( .A(n1562), .B(n1386), .ZN(n908) );
  XNOR2_X1 U1554 ( .A(n1373), .B(n1386), .ZN(n910) );
  XNOR2_X1 U1555 ( .A(n1381), .B(n1386), .ZN(n911) );
  XNOR2_X1 U1556 ( .A(n1559), .B(n1386), .ZN(n912) );
  XNOR2_X1 U1557 ( .A(n1367), .B(n1386), .ZN(n913) );
  XNOR2_X1 U1558 ( .A(n1366), .B(n1386), .ZN(n914) );
  XNOR2_X1 U1559 ( .A(n1370), .B(n1386), .ZN(n916) );
  XNOR2_X1 U1560 ( .A(n1556), .B(n1386), .ZN(n915) );
  XNOR2_X1 U1561 ( .A(n1375), .B(n1386), .ZN(n917) );
  XNOR2_X1 U1562 ( .A(n1364), .B(n1386), .ZN(n909) );
  XNOR2_X1 U1563 ( .A(n1357), .B(n1386), .ZN(n918) );
  XNOR2_X1 U1564 ( .A(n1361), .B(n1386), .ZN(n919) );
  XNOR2_X1 U1565 ( .A(n1564), .B(n1386), .ZN(n905) );
  XNOR2_X1 U1566 ( .A(n1282), .B(n1386), .ZN(n902) );
  XNOR2_X1 U1567 ( .A(n1383), .B(n1386), .ZN(n904) );
  XNOR2_X1 U1568 ( .A(n1565), .B(n1386), .ZN(n903) );
  AND2_X1 U1569 ( .A1(n1551), .A2(n665), .ZN(n859) );
  BUF_X1 U1570 ( .A(n1098), .Z(n1561) );
  BUF_X1 U1571 ( .A(n1099), .Z(n1560) );
  BUF_X1 U1572 ( .A(n1102), .Z(n1558) );
  BUF_X1 U1573 ( .A(n1105), .Z(n1555) );
  BUF_X1 U1574 ( .A(n1106), .Z(n1554) );
  BUF_X1 U1575 ( .A(n1107), .Z(n1553) );
  INV_X1 U1576 ( .A(n655), .ZN(n780) );
  INV_X1 U1577 ( .A(n314), .ZN(n315) );
  AND2_X1 U1578 ( .A1(n1355), .A2(n641), .ZN(n699) );
  OAI22_X1 U1579 ( .A1(n1347), .A2(n1071), .B1(n1070), .B2(n4), .ZN(n862) );
  OAI22_X1 U1580 ( .A1(n1348), .A2(n1072), .B1(n1071), .B2(n4), .ZN(n863) );
  INV_X1 U1581 ( .A(n649), .ZN(n740) );
  INV_X1 U1582 ( .A(n346), .ZN(n347) );
  AND2_X1 U1583 ( .A1(n1355), .A2(n644), .ZN(n719) );
  OAI22_X1 U1584 ( .A1(n1347), .A2(n1073), .B1(n1072), .B2(n4), .ZN(n864) );
  OAI22_X1 U1585 ( .A1(n1077), .A2(n1348), .B1(n1076), .B2(n4), .ZN(n868) );
  AND2_X1 U1586 ( .A1(n1355), .A2(n650), .ZN(n759) );
  INV_X1 U1587 ( .A(n667), .ZN(n860) );
  INV_X1 U1588 ( .A(n652), .ZN(n760) );
  INV_X1 U1589 ( .A(n646), .ZN(n720) );
  INV_X1 U1590 ( .A(n424), .ZN(n425) );
  OAI22_X1 U1591 ( .A1(n1347), .A2(n1080), .B1(n1079), .B2(n4), .ZN(n871) );
  AND2_X1 U1592 ( .A1(n1355), .A2(n659), .ZN(n819) );
  OAI22_X1 U1593 ( .A1(n1348), .A2(n1083), .B1(n1082), .B2(n4), .ZN(n874) );
  OAI22_X1 U1594 ( .A1(n1347), .A2(n1076), .B1(n1075), .B2(n4), .ZN(n867) );
  INV_X1 U1595 ( .A(n458), .ZN(n459) );
  OAI22_X1 U1596 ( .A1(n1347), .A2(n1070), .B1(n1262), .B2(n4), .ZN(n861) );
  OAI22_X1 U1597 ( .A1(n1348), .A2(n1074), .B1(n1073), .B2(n4), .ZN(n865) );
  OAI22_X1 U1598 ( .A1(n1280), .A2(n1081), .B1(n1080), .B2(n4), .ZN(n872) );
  AND2_X1 U1599 ( .A1(n1355), .A2(n656), .ZN(n799) );
  INV_X1 U1600 ( .A(n640), .ZN(n680) );
  INV_X1 U1601 ( .A(n368), .ZN(n369) );
  INV_X1 U1602 ( .A(n658), .ZN(n800) );
  INV_X1 U1603 ( .A(n1386), .ZN(n1141) );
  OR2_X1 U1604 ( .A1(n1354), .A2(n1393), .ZN(n900) );
  OR2_X1 U1605 ( .A1(n1354), .A2(n1342), .ZN(n963) );
  OR2_X1 U1606 ( .A1(n1355), .A2(n1144), .ZN(n984) );
  OR2_X1 U1607 ( .A1(n1354), .A2(n1146), .ZN(n1026) );
  OR2_X1 U1608 ( .A1(n1551), .A2(n1142), .ZN(n942) );
  OR2_X1 U1609 ( .A1(n1551), .A2(n1141), .ZN(n921) );
  OR2_X1 U1610 ( .A1(n1354), .A2(n1145), .ZN(n1005) );
  AND2_X1 U1611 ( .A1(n1551), .A2(n668), .ZN(product[0]) );
  XNOR2_X1 U1612 ( .A(n43), .B(a[16]), .ZN(n52) );
  XNOR2_X1 U1613 ( .A(n13), .B(a[6]), .ZN(n22) );
  XNOR2_X1 U1614 ( .A(n25), .B(a[10]), .ZN(n34) );
  XNOR2_X1 U1615 ( .A(n7), .B(a[4]), .ZN(n16) );
  XNOR2_X1 U1616 ( .A(n19), .B(a[8]), .ZN(n28) );
  XNOR2_X1 U1617 ( .A(n31), .B(a[12]), .ZN(n40) );
  XNOR2_X1 U1618 ( .A(n1549), .B(a[18]), .ZN(n58) );
  XNOR2_X1 U1619 ( .A(n37), .B(a[14]), .ZN(n46) );
  XNOR2_X1 U1620 ( .A(n1), .B(a[2]), .ZN(n9) );
  XNOR2_X1 U1621 ( .A(n1282), .B(n1387), .ZN(n923) );
  XNOR2_X1 U1622 ( .A(n1384), .B(n1388), .ZN(n922) );
  XNOR2_X1 U1623 ( .A(n1565), .B(n1387), .ZN(n924) );
  XNOR2_X1 U1624 ( .A(n1564), .B(n1388), .ZN(n926) );
  XNOR2_X1 U1625 ( .A(n1382), .B(n1387), .ZN(n925) );
  XNOR2_X1 U1626 ( .A(n1352), .B(n1388), .ZN(n927) );
  XNOR2_X1 U1627 ( .A(n1563), .B(n1387), .ZN(n928) );
  XNOR2_X1 U1628 ( .A(n1562), .B(n1388), .ZN(n929) );
  XNOR2_X1 U1629 ( .A(n1362), .B(n1387), .ZN(n930) );
  XNOR2_X1 U1630 ( .A(n1380), .B(n1388), .ZN(n932) );
  XNOR2_X1 U1631 ( .A(n1372), .B(n1387), .ZN(n931) );
  XNOR2_X1 U1632 ( .A(n1559), .B(n1388), .ZN(n933) );
  XNOR2_X1 U1633 ( .A(n1557), .B(n1388), .ZN(n935) );
  XNOR2_X1 U1634 ( .A(n1368), .B(n1387), .ZN(n934) );
  XNOR2_X1 U1635 ( .A(n1358), .B(n1388), .ZN(n939) );
  XNOR2_X1 U1636 ( .A(n1550), .B(n1387), .ZN(n941) );
  XNOR2_X1 U1637 ( .A(n1361), .B(n1387), .ZN(n940) );
  XNOR2_X1 U1638 ( .A(n1375), .B(n1387), .ZN(n938) );
  XNOR2_X1 U1639 ( .A(n1555), .B(n1388), .ZN(n937) );
  XNOR2_X1 U1640 ( .A(n1556), .B(n1388), .ZN(n936) );
  INV_X1 U1641 ( .A(n1387), .ZN(n1142) );
  NAND2_X1 U1642 ( .A1(n815), .A2(n870), .ZN(n1511) );
  NAND2_X1 U1643 ( .A1(n815), .A2(n779), .ZN(n1512) );
  NAND2_X1 U1644 ( .A1(n870), .A2(n779), .ZN(n1513) );
  NAND3_X1 U1645 ( .A1(n1511), .A2(n1512), .A3(n1513), .ZN(n606) );
  NAND2_X1 U1646 ( .A1(n612), .A2(n614), .ZN(n1514) );
  NAND2_X1 U1647 ( .A1(n612), .A2(n607), .ZN(n1515) );
  NAND2_X1 U1648 ( .A1(n614), .A2(n607), .ZN(n1516) );
  NAND3_X1 U1649 ( .A1(n1514), .A2(n1515), .A3(n1516), .ZN(n602) );
  NAND2_X1 U1650 ( .A1(n610), .A2(n605), .ZN(n1517) );
  NAND2_X1 U1651 ( .A1(n610), .A2(n603), .ZN(n1518) );
  NAND2_X1 U1652 ( .A1(n605), .A2(n603), .ZN(n1519) );
  AND2_X1 U1653 ( .A1(n1355), .A2(n653), .ZN(n779) );
  OAI22_X1 U1654 ( .A1(n1280), .A2(n1079), .B1(n1078), .B2(n4), .ZN(n870) );
  XNOR2_X1 U1655 ( .A(n1384), .B(n1369), .ZN(n880) );
  XNOR2_X1 U1656 ( .A(n1282), .B(n1344), .ZN(n881) );
  XNOR2_X1 U1657 ( .A(n1565), .B(n1369), .ZN(n882) );
  XNOR2_X1 U1658 ( .A(n1382), .B(n1344), .ZN(n883) );
  XNOR2_X1 U1659 ( .A(n1352), .B(n1344), .ZN(n885) );
  XNOR2_X1 U1660 ( .A(n1564), .B(n1369), .ZN(n884) );
  XNOR2_X1 U1661 ( .A(n1563), .B(n1369), .ZN(n886) );
  XNOR2_X1 U1662 ( .A(n1562), .B(n1344), .ZN(n887) );
  XNOR2_X1 U1663 ( .A(n1362), .B(n1369), .ZN(n888) );
  XNOR2_X1 U1664 ( .A(n1372), .B(n1344), .ZN(n889) );
  XNOR2_X1 U1665 ( .A(n1380), .B(n1369), .ZN(n890) );
  XNOR2_X1 U1666 ( .A(n1559), .B(n1344), .ZN(n891) );
  XNOR2_X1 U1667 ( .A(n1367), .B(n1369), .ZN(n892) );
  XNOR2_X1 U1668 ( .A(n1556), .B(n55), .ZN(n894) );
  XNOR2_X1 U1669 ( .A(n1365), .B(n1369), .ZN(n893) );
  XNOR2_X1 U1670 ( .A(n1355), .B(n1369), .ZN(n899) );
  XNOR2_X1 U1671 ( .A(n1370), .B(n1369), .ZN(n895) );
  XNOR2_X1 U1672 ( .A(n1552), .B(n1369), .ZN(n898) );
  XNOR2_X1 U1673 ( .A(n1356), .B(n1369), .ZN(n897) );
  XNOR2_X1 U1674 ( .A(n1374), .B(n1369), .ZN(n896) );
  INV_X1 U1675 ( .A(n215), .ZN(n286) );
  NOR2_X1 U1676 ( .A1(n215), .A2(n218), .ZN(n213) );
  OAI21_X1 U1677 ( .B1(n215), .B2(n219), .A(n216), .ZN(n214) );
  NAND2_X1 U1678 ( .A1(n601), .A2(n608), .ZN(n227) );
  NAND2_X1 U1679 ( .A1(n866), .A2(n775), .ZN(n1520) );
  NAND2_X1 U1680 ( .A1(n775), .A2(n739), .ZN(n1521) );
  NAND2_X1 U1681 ( .A1(n866), .A2(n739), .ZN(n1522) );
  NAND3_X1 U1682 ( .A1(n1520), .A2(n1521), .A3(n1522), .ZN(n566) );
  AND2_X1 U1683 ( .A1(n1355), .A2(n647), .ZN(n739) );
  OAI22_X1 U1684 ( .A1(n1283), .A2(n1075), .B1(n1074), .B2(n4), .ZN(n866) );
  NOR2_X1 U1685 ( .A1(n383), .A2(n396), .ZN(n140) );
  NAND2_X1 U1686 ( .A1(n383), .A2(n396), .ZN(n141) );
  INV_X1 U1687 ( .A(n145), .ZN(n143) );
  NOR2_X1 U1688 ( .A1(n131), .A2(n128), .ZN(n126) );
  NAND3_X1 U1689 ( .A1(n1529), .A2(n1528), .A3(n1527), .ZN(n1524) );
  NAND3_X1 U1690 ( .A1(n1527), .A2(n1337), .A3(n1389), .ZN(n1525) );
  XOR2_X1 U1691 ( .A(n303), .B(n306), .Z(n1526) );
  XOR2_X1 U1692 ( .A(n1526), .B(n1339), .Z(product[35]) );
  NAND2_X1 U1693 ( .A1(n303), .A2(n306), .ZN(n1527) );
  NAND2_X1 U1694 ( .A1(n303), .A2(n100), .ZN(n1528) );
  NAND2_X1 U1695 ( .A1(n1434), .A2(n306), .ZN(n1529) );
  NAND3_X1 U1696 ( .A1(n1529), .A2(n1528), .A3(n1527), .ZN(n99) );
  NAND2_X1 U1697 ( .A1(n302), .A2(n301), .ZN(n1530) );
  NAND2_X1 U1698 ( .A1(n1524), .A2(n302), .ZN(n1531) );
  NAND2_X1 U1699 ( .A1(n301), .A2(n99), .ZN(n1532) );
  NAND3_X1 U1700 ( .A1(n1532), .A2(n1531), .A3(n1530), .ZN(n98) );
  NAND2_X1 U1701 ( .A1(n546), .A2(n548), .ZN(n1533) );
  NAND2_X1 U1702 ( .A1(n546), .A2(n535), .ZN(n1534) );
  NAND2_X1 U1703 ( .A1(n548), .A2(n535), .ZN(n1535) );
  NAND3_X1 U1704 ( .A1(n1533), .A2(n1534), .A3(n1535), .ZN(n530) );
  NAND2_X1 U1705 ( .A1(n544), .A2(n533), .ZN(n1536) );
  NAND2_X1 U1706 ( .A1(n531), .A2(n544), .ZN(n1537) );
  NAND2_X1 U1707 ( .A1(n531), .A2(n533), .ZN(n1538) );
  NAND3_X1 U1708 ( .A1(n1536), .A2(n1537), .A3(n1538), .ZN(n528) );
  NAND2_X1 U1709 ( .A1(n513), .A2(n528), .ZN(n185) );
  OAI21_X1 U1710 ( .B1(n166), .B2(n172), .A(n167), .ZN(n165) );
  XNOR2_X1 U1711 ( .A(n1384), .B(n1343), .ZN(n943) );
  XNOR2_X1 U1712 ( .A(n1282), .B(n1343), .ZN(n944) );
  XNOR2_X1 U1713 ( .A(n1383), .B(n1343), .ZN(n946) );
  XNOR2_X1 U1714 ( .A(n1565), .B(n1343), .ZN(n945) );
  XNOR2_X1 U1715 ( .A(n1564), .B(n1343), .ZN(n947) );
  XNOR2_X1 U1716 ( .A(n1353), .B(n1343), .ZN(n948) );
  XNOR2_X1 U1717 ( .A(n1563), .B(n1278), .ZN(n949) );
  XNOR2_X1 U1718 ( .A(n1362), .B(n1278), .ZN(n951) );
  XNOR2_X1 U1719 ( .A(n1373), .B(n1278), .ZN(n952) );
  XNOR2_X1 U1720 ( .A(n1562), .B(n1278), .ZN(n950) );
  XNOR2_X1 U1721 ( .A(n1366), .B(n1278), .ZN(n956) );
  XNOR2_X1 U1722 ( .A(n1368), .B(n1407), .ZN(n955) );
  XNOR2_X1 U1723 ( .A(n1556), .B(n1278), .ZN(n957) );
  XNOR2_X1 U1724 ( .A(n1100), .B(n1407), .ZN(n953) );
  XNOR2_X1 U1725 ( .A(n1559), .B(n1407), .ZN(n954) );
  XNOR2_X1 U1726 ( .A(n1357), .B(n1278), .ZN(n960) );
  XNOR2_X1 U1727 ( .A(n1374), .B(n1278), .ZN(n959) );
  XNOR2_X1 U1728 ( .A(n1555), .B(n1278), .ZN(n958) );
  XNOR2_X1 U1729 ( .A(n1550), .B(n1278), .ZN(n962) );
  XNOR2_X1 U1730 ( .A(n1552), .B(n1407), .ZN(n961) );
  OAI21_X1 U1731 ( .B1(n248), .B2(n250), .A(n249), .ZN(n247) );
  NAND2_X1 U1732 ( .A1(n1485), .A2(n200), .ZN(n81) );
  NAND2_X1 U1733 ( .A1(n202), .A2(n1485), .ZN(n195) );
  NAND2_X1 U1734 ( .A1(n532), .A2(n521), .ZN(n1539) );
  NAND2_X1 U1735 ( .A1(n532), .A2(n519), .ZN(n1540) );
  NAND2_X1 U1736 ( .A1(n521), .A2(n519), .ZN(n1541) );
  NAND3_X1 U1737 ( .A1(n1539), .A2(n1540), .A3(n1541), .ZN(n514) );
  NAND2_X1 U1738 ( .A1(n517), .A2(n1289), .ZN(n1542) );
  NAND2_X1 U1739 ( .A1(n517), .A2(n515), .ZN(n1543) );
  NAND2_X1 U1740 ( .A1(n1289), .A2(n515), .ZN(n1544) );
  XNOR2_X1 U1741 ( .A(n1556), .B(n1546), .ZN(n1062) );
  XNOR2_X1 U1742 ( .A(n1559), .B(n1546), .ZN(n1059) );
  INV_X1 U1743 ( .A(n1546), .ZN(n1148) );
  XNOR2_X1 U1744 ( .A(n1565), .B(n1546), .ZN(n1050) );
  XNOR2_X1 U1745 ( .A(n1566), .B(n1546), .ZN(n1049) );
  XNOR2_X1 U1746 ( .A(n1365), .B(n1546), .ZN(n1061) );
  XNOR2_X1 U1747 ( .A(n1558), .B(n1546), .ZN(n1060) );
  XNOR2_X1 U1748 ( .A(n1564), .B(n1546), .ZN(n1052) );
  XNOR2_X1 U1749 ( .A(n1382), .B(n1546), .ZN(n1051) );
  XNOR2_X1 U1750 ( .A(n1375), .B(n1546), .ZN(n1064) );
  XNOR2_X1 U1751 ( .A(n1370), .B(n1546), .ZN(n1063) );
  XNOR2_X1 U1752 ( .A(n1381), .B(n1546), .ZN(n1058) );
  XNOR2_X1 U1753 ( .A(n1562), .B(n1546), .ZN(n1055) );
  XNOR2_X1 U1754 ( .A(n1372), .B(n1546), .ZN(n1057) );
  XNOR2_X1 U1755 ( .A(n1364), .B(n1546), .ZN(n1056) );
  XNOR2_X1 U1756 ( .A(n1354), .B(n1546), .ZN(n1067) );
  XNOR2_X1 U1757 ( .A(n1090), .B(n7), .ZN(n1048) );
  XNOR2_X1 U1758 ( .A(n1563), .B(n1546), .ZN(n1054) );
  XNOR2_X1 U1759 ( .A(n1361), .B(n1546), .ZN(n1066) );
  XNOR2_X1 U1760 ( .A(n1352), .B(n1546), .ZN(n1053) );
  XNOR2_X1 U1761 ( .A(n1358), .B(n1546), .ZN(n1065) );
  BUF_X4 U1762 ( .A(n7), .Z(n1546) );
  INV_X1 U1763 ( .A(n1275), .ZN(n1146) );
  XNOR2_X1 U1764 ( .A(n1324), .B(n1275), .ZN(n1006) );
  XNOR2_X1 U1765 ( .A(n1383), .B(n1275), .ZN(n1009) );
  XNOR2_X1 U1766 ( .A(n1551), .B(n1275), .ZN(n1025) );
  XNOR2_X1 U1767 ( .A(n1565), .B(n1275), .ZN(n1008) );
  XNOR2_X1 U1768 ( .A(n1108), .B(n1275), .ZN(n1024) );
  XNOR2_X1 U1769 ( .A(n1566), .B(n1275), .ZN(n1007) );
  XNOR2_X1 U1770 ( .A(n1357), .B(n1275), .ZN(n1023) );
  XNOR2_X1 U1771 ( .A(n1364), .B(n1275), .ZN(n1014) );
  XNOR2_X1 U1772 ( .A(n1095), .B(n1547), .ZN(n1011) );
  XNOR2_X1 U1773 ( .A(n1556), .B(n1275), .ZN(n1020) );
  XNOR2_X1 U1774 ( .A(n1564), .B(n1547), .ZN(n1010) );
  XNOR2_X1 U1775 ( .A(n1562), .B(n1547), .ZN(n1013) );
  XNOR2_X1 U1776 ( .A(n1563), .B(n1547), .ZN(n1012) );
  XNOR2_X1 U1777 ( .A(n1558), .B(n1547), .ZN(n1018) );
  XNOR2_X1 U1778 ( .A(n1366), .B(n1547), .ZN(n1019) );
  XNOR2_X1 U1779 ( .A(n1375), .B(n1275), .ZN(n1022) );
  XNOR2_X1 U1780 ( .A(n1370), .B(n1275), .ZN(n1021) );
  XNOR2_X1 U1781 ( .A(n1373), .B(n1275), .ZN(n1015) );
  XNOR2_X1 U1782 ( .A(n1380), .B(n1547), .ZN(n1016) );
  XNOR2_X1 U1783 ( .A(n1559), .B(n19), .ZN(n1017) );
  XNOR2_X1 U1784 ( .A(n1384), .B(n1548), .ZN(n964) );
  XNOR2_X1 U1785 ( .A(n1566), .B(n1548), .ZN(n965) );
  XNOR2_X1 U1786 ( .A(n1565), .B(n1548), .ZN(n966) );
  XNOR2_X1 U1787 ( .A(n1382), .B(n1548), .ZN(n967) );
  XNOR2_X1 U1788 ( .A(n1362), .B(n1548), .ZN(n972) );
  XNOR2_X1 U1789 ( .A(n1564), .B(n1548), .ZN(n968) );
  XNOR2_X1 U1790 ( .A(n1562), .B(n1548), .ZN(n971) );
  XNOR2_X1 U1791 ( .A(n1563), .B(n1548), .ZN(n970) );
  XNOR2_X1 U1792 ( .A(n1353), .B(n1548), .ZN(n969) );
  INV_X1 U1793 ( .A(n1548), .ZN(n1144) );
  XNOR2_X1 U1794 ( .A(n1560), .B(n1548), .ZN(n973) );
  XNOR2_X1 U1795 ( .A(n1381), .B(n1548), .ZN(n974) );
  XNOR2_X1 U1796 ( .A(n1558), .B(n1548), .ZN(n976) );
  XNOR2_X1 U1797 ( .A(n1101), .B(n1548), .ZN(n975) );
  XNOR2_X1 U1798 ( .A(n1550), .B(n1548), .ZN(n983) );
  XNOR2_X1 U1799 ( .A(n1552), .B(n1548), .ZN(n982) );
  XNOR2_X1 U1800 ( .A(n1557), .B(n1548), .ZN(n977) );
  XNOR2_X1 U1801 ( .A(n1556), .B(n1548), .ZN(n978) );
  XNOR2_X1 U1802 ( .A(n1371), .B(n1548), .ZN(n979) );
  XNOR2_X1 U1803 ( .A(n1374), .B(n1548), .ZN(n980) );
  XNOR2_X1 U1804 ( .A(n1356), .B(n1548), .ZN(n981) );
  OAI21_X1 U1805 ( .B1(n151), .B2(n147), .A(n148), .ZN(n146) );
  OAI21_X1 U1806 ( .B1(n152), .B2(n1378), .A(n1454), .ZN(n149) );
  NAND2_X1 U1807 ( .A1(n275), .A2(n1454), .ZN(n73) );
  NAND2_X1 U1808 ( .A1(n411), .A2(n426), .ZN(n151) );
  AOI21_X1 U1809 ( .B1(n173), .B2(n164), .A(n165), .ZN(n163) );
  NAND2_X1 U1810 ( .A1(n461), .A2(n478), .ZN(n167) );
  NAND2_X1 U1811 ( .A1(n1494), .A2(n227), .ZN(n86) );
  INV_X1 U1812 ( .A(n221), .ZN(n220) );
  AOI21_X1 U1813 ( .B1(n221), .B2(n213), .A(n214), .ZN(n212) );
  NAND2_X1 U1814 ( .A1(n1494), .A2(n1489), .ZN(n222) );
  AOI21_X1 U1815 ( .B1(n1494), .B2(n230), .A(n225), .ZN(n223) );
  XNOR2_X1 U1816 ( .A(n1357), .B(n1349), .ZN(n1044) );
  INV_X1 U1817 ( .A(n1349), .ZN(n1147) );
  XNOR2_X1 U1818 ( .A(n1564), .B(n1349), .ZN(n1031) );
  XNOR2_X1 U1819 ( .A(n1365), .B(n1350), .ZN(n1040) );
  XNOR2_X1 U1820 ( .A(n1558), .B(n1349), .ZN(n1039) );
  XNOR2_X1 U1821 ( .A(n1559), .B(n1350), .ZN(n1038) );
  XNOR2_X1 U1822 ( .A(n1380), .B(n1349), .ZN(n1037) );
  XNOR2_X1 U1823 ( .A(n1551), .B(n1350), .ZN(n1046) );
  XNOR2_X1 U1824 ( .A(n1375), .B(n1350), .ZN(n1043) );
  XNOR2_X1 U1825 ( .A(n1361), .B(n1350), .ZN(n1045) );
  XNOR2_X1 U1826 ( .A(n1373), .B(n1349), .ZN(n1036) );
  XNOR2_X1 U1827 ( .A(n1324), .B(n1349), .ZN(n1027) );
  XNOR2_X1 U1828 ( .A(n1556), .B(n1350), .ZN(n1041) );
  XNOR2_X1 U1829 ( .A(n1371), .B(n1349), .ZN(n1042) );
  XNOR2_X1 U1830 ( .A(n1563), .B(n1350), .ZN(n1033) );
  XNOR2_X1 U1831 ( .A(n1565), .B(n1349), .ZN(n1029) );
  XNOR2_X1 U1832 ( .A(n1093), .B(n1350), .ZN(n1030) );
  XNOR2_X1 U1833 ( .A(n1353), .B(n1350), .ZN(n1032) );
  XNOR2_X1 U1834 ( .A(n1566), .B(n1349), .ZN(n1028) );
  XNOR2_X1 U1835 ( .A(n1363), .B(n1350), .ZN(n1035) );
  XNOR2_X1 U1836 ( .A(n1562), .B(n1349), .ZN(n1034) );
  AOI21_X1 U1837 ( .B1(n211), .B2(n202), .A(n203), .ZN(n201) );
  INV_X1 U1838 ( .A(n1321), .ZN(n284) );
  AOI21_X1 U1839 ( .B1(n203), .B2(n1485), .A(n198), .ZN(n196) );
  NOR2_X1 U1840 ( .A1(n1321), .A2(n209), .ZN(n202) );
  OAI21_X1 U1841 ( .B1(n204), .B2(n210), .A(n205), .ZN(n203) );
  INV_X1 U1842 ( .A(n135), .ZN(n272) );
  NOR2_X1 U1843 ( .A1(n140), .A2(n135), .ZN(n133) );
  OAI21_X1 U1844 ( .B1(n141), .B2(n135), .A(n136), .ZN(n134) );
  NAND2_X1 U1845 ( .A1(n371), .A2(n382), .ZN(n136) );
  XNOR2_X1 U1846 ( .A(n239), .B(n88), .ZN(product[8]) );
  INV_X1 U1847 ( .A(n234), .ZN(n233) );
  OAI21_X1 U1848 ( .B1(n222), .B2(n234), .A(n223), .ZN(n221) );
  AOI21_X1 U1849 ( .B1(n239), .B2(n1492), .A(n236), .ZN(n234) );
  NAND2_X1 U1850 ( .A1(n637), .A2(n638), .ZN(n254) );
  XNOR2_X1 U1851 ( .A(n1559), .B(n1270), .ZN(n1080) );
  XNOR2_X1 U1852 ( .A(n1367), .B(n1270), .ZN(n1081) );
  XNOR2_X1 U1853 ( .A(n1564), .B(n1270), .ZN(n1073) );
  XNOR2_X1 U1854 ( .A(n1565), .B(n1270), .ZN(n1071) );
  XNOR2_X1 U1855 ( .A(n1382), .B(n1284), .ZN(n1072) );
  XNOR2_X1 U1856 ( .A(n1566), .B(n1270), .ZN(n1070) );
  XNOR2_X1 U1857 ( .A(n1563), .B(n1270), .ZN(n1075) );
  XNOR2_X1 U1858 ( .A(n1562), .B(n1270), .ZN(n1076) );
  XNOR2_X1 U1859 ( .A(n1352), .B(n1545), .ZN(n1074) );
  XNOR2_X1 U1860 ( .A(n1363), .B(n1270), .ZN(n1077) );
  XNOR2_X1 U1861 ( .A(n1381), .B(n1284), .ZN(n1079) );
  XNOR2_X1 U1862 ( .A(n1366), .B(n1284), .ZN(n1082) );
  XNOR2_X1 U1863 ( .A(n1372), .B(n1270), .ZN(n1078) );
  XNOR2_X1 U1864 ( .A(n1556), .B(n1270), .ZN(n1083) );
  XNOR2_X1 U1865 ( .A(n1324), .B(n1545), .ZN(n1069) );
  XNOR2_X1 U1866 ( .A(n1354), .B(n1270), .ZN(n1088) );
  XNOR2_X1 U1867 ( .A(n1358), .B(n1284), .ZN(n1086) );
  XNOR2_X1 U1868 ( .A(n1375), .B(n1284), .ZN(n1085) );
  INV_X1 U1869 ( .A(n1284), .ZN(n1149) );
  XNOR2_X1 U1870 ( .A(n1108), .B(n1270), .ZN(n1087) );
  XNOR2_X1 U1871 ( .A(n1371), .B(n1270), .ZN(n1084) );
  XOR2_X1 U1872 ( .A(n1), .B(n668), .Z(n1119) );
  INV_X1 U1873 ( .A(n664), .ZN(n840) );
  NAND2_X1 U1874 ( .A1(n397), .A2(n410), .ZN(n148) );
  NAND2_X1 U1875 ( .A1(n145), .A2(n133), .ZN(n131) );
  INV_X1 U1876 ( .A(n1455), .ZN(n144) );
  AOI21_X1 U1877 ( .B1(n146), .B2(n133), .A(n134), .ZN(n132) );
  OAI21_X1 U1878 ( .B1(n193), .B2(n180), .A(n1247), .ZN(n179) );
  BUF_X4 U1879 ( .A(n31), .Z(n1548) );
  NAND2_X1 U1880 ( .A1(n1486), .A2(n185), .ZN(n79) );
  NAND2_X1 U1881 ( .A1(n156), .A2(n164), .ZN(n154) );
  AOI21_X1 U1882 ( .B1(n165), .B2(n156), .A(n157), .ZN(n155) );
  XNOR2_X1 U1883 ( .A(n787), .B(n715), .ZN(n477) );
  OR2_X1 U1884 ( .A1(n787), .A2(n715), .ZN(n476) );
  OAI21_X1 U1885 ( .B1(n193), .B2(n187), .A(n188), .ZN(n186) );
  NOR2_X1 U1886 ( .A1(n150), .A2(n1468), .ZN(n145) );
  NOR2_X1 U1887 ( .A1(n161), .A2(n1475), .ZN(n156) );
  OAI21_X1 U1888 ( .B1(n158), .B2(n162), .A(n159), .ZN(n157) );
  NAND2_X1 U1889 ( .A1(n427), .A2(n442), .ZN(n159) );
  OAI22_X1 U1890 ( .A1(n1466), .A2(n965), .B1(n964), .B2(n1506), .ZN(n346) );
  OAI22_X1 U1891 ( .A1(n964), .A2(n1467), .B1(n964), .B2(n1506), .ZN(n652) );
  OAI22_X1 U1892 ( .A1(n1467), .A2(n966), .B1(n965), .B2(n1506), .ZN(n761) );
  OAI22_X1 U1893 ( .A1(n1466), .A2(n967), .B1(n966), .B2(n1261), .ZN(n762) );
  XNOR2_X1 U1894 ( .A(n1384), .B(n1331), .ZN(n985) );
  OAI22_X1 U1895 ( .A1(n1467), .A2(n968), .B1(n967), .B2(n1261), .ZN(n763) );
  XNOR2_X1 U1896 ( .A(n1566), .B(n1332), .ZN(n986) );
  OAI22_X1 U1897 ( .A1(n1466), .A2(n972), .B1(n971), .B2(n1261), .ZN(n767) );
  OAI22_X1 U1898 ( .A1(n1467), .A2(n975), .B1(n974), .B2(n1506), .ZN(n770) );
  OAI22_X1 U1899 ( .A1(n1467), .A2(n973), .B1(n972), .B2(n1261), .ZN(n768) );
  OAI22_X1 U1900 ( .A1(n1466), .A2(n1144), .B1(n984), .B2(n1506), .ZN(n674) );
  OAI22_X1 U1901 ( .A1(n1467), .A2(n969), .B1(n968), .B2(n1506), .ZN(n764) );
  OAI22_X1 U1902 ( .A1(n1466), .A2(n983), .B1(n982), .B2(n1506), .ZN(n778) );
  OAI22_X1 U1903 ( .A1(n1467), .A2(n977), .B1(n976), .B2(n1506), .ZN(n772) );
  OAI22_X1 U1904 ( .A1(n1466), .A2(n971), .B1(n970), .B2(n1506), .ZN(n766) );
  OAI22_X1 U1905 ( .A1(n1466), .A2(n970), .B1(n969), .B2(n1506), .ZN(n765) );
  OAI22_X1 U1906 ( .A1(n1466), .A2(n978), .B1(n977), .B2(n1506), .ZN(n773) );
  OAI22_X1 U1907 ( .A1(n1466), .A2(n982), .B1(n981), .B2(n1506), .ZN(n777) );
  XNOR2_X1 U1908 ( .A(n1564), .B(n1332), .ZN(n989) );
  OAI22_X1 U1909 ( .A1(n1467), .A2(n979), .B1(n978), .B2(n1506), .ZN(n774) );
  OAI22_X1 U1910 ( .A1(n36), .A2(n976), .B1(n975), .B2(n1506), .ZN(n771) );
  OAI22_X1 U1911 ( .A1(n1467), .A2(n980), .B1(n979), .B2(n1506), .ZN(n775) );
  XNOR2_X1 U1912 ( .A(n1383), .B(n1332), .ZN(n988) );
  XNOR2_X1 U1913 ( .A(n1551), .B(n1332), .ZN(n1004) );
  XNOR2_X1 U1914 ( .A(n1565), .B(n1331), .ZN(n987) );
  XNOR2_X1 U1915 ( .A(n1556), .B(n1331), .ZN(n999) );
  XNOR2_X1 U1916 ( .A(n1358), .B(n1331), .ZN(n1002) );
  XNOR2_X1 U1917 ( .A(n1361), .B(n1331), .ZN(n1003) );
  OAI22_X1 U1918 ( .A1(n1467), .A2(n974), .B1(n973), .B2(n1506), .ZN(n769) );
  INV_X1 U1919 ( .A(n1261), .ZN(n653) );
  OAI22_X1 U1920 ( .A1(n1466), .A2(n981), .B1(n980), .B2(n1506), .ZN(n776) );
  XNOR2_X1 U1921 ( .A(n1563), .B(n1332), .ZN(n991) );
  XNOR2_X1 U1922 ( .A(n1380), .B(n1332), .ZN(n995) );
  INV_X1 U1923 ( .A(n1331), .ZN(n1145) );
  XNOR2_X1 U1924 ( .A(n1352), .B(n1332), .ZN(n990) );
  XNOR2_X1 U1925 ( .A(n1559), .B(n1332), .ZN(n996) );
  XNOR2_X1 U1926 ( .A(n1555), .B(n1331), .ZN(n1000) );
  XNOR2_X1 U1927 ( .A(n1375), .B(n1331), .ZN(n1001) );
  XNOR2_X1 U1928 ( .A(n1365), .B(n1332), .ZN(n998) );
  XNOR2_X1 U1929 ( .A(n1560), .B(n1331), .ZN(n994) );
  XNOR2_X1 U1930 ( .A(n1367), .B(n1332), .ZN(n997) );
  XNOR2_X1 U1931 ( .A(n1363), .B(n1332), .ZN(n993) );
  XNOR2_X1 U1932 ( .A(n1562), .B(n1331), .ZN(n992) );
  INV_X1 U1933 ( .A(n1428), .ZN(n193) );
  INV_X1 U1934 ( .A(n1281), .ZN(n211) );
  OAI21_X1 U1935 ( .B1(n195), .B2(n212), .A(n196), .ZN(n194) );
  OAI22_X1 U1936 ( .A1(n1336), .A2(n1053), .B1(n1052), .B2(n1509), .ZN(n844)
         );
  OAI22_X1 U1937 ( .A1(n1469), .A2(n1055), .B1(n1054), .B2(n1510), .ZN(n846)
         );
  OAI22_X1 U1938 ( .A1(n1469), .A2(n1051), .B1(n1050), .B2(n1509), .ZN(n842)
         );
  OAI22_X1 U1939 ( .A1(n1469), .A2(n1062), .B1(n1061), .B2(n1510), .ZN(n853)
         );
  OAI22_X1 U1940 ( .A1(n1336), .A2(n1059), .B1(n1058), .B2(n1509), .ZN(n850)
         );
  OAI22_X1 U1941 ( .A1(n1336), .A2(n1060), .B1(n1059), .B2(n1509), .ZN(n851)
         );
  OAI22_X1 U1942 ( .A1(n1336), .A2(n1063), .B1(n1062), .B2(n1509), .ZN(n854)
         );
  OAI22_X1 U1943 ( .A1(n12), .A2(n1054), .B1(n1053), .B2(n1510), .ZN(n845) );
  OAI22_X1 U1944 ( .A1(n12), .A2(n1049), .B1(n1048), .B2(n1509), .ZN(n458) );
  OAI22_X1 U1945 ( .A1(n1469), .A2(n1056), .B1(n1055), .B2(n1510), .ZN(n847)
         );
  OAI22_X1 U1946 ( .A1(n1336), .A2(n1052), .B1(n1051), .B2(n1509), .ZN(n843)
         );
  OAI22_X1 U1947 ( .A1(n1469), .A2(n1057), .B1(n1056), .B2(n1509), .ZN(n848)
         );
  OAI22_X1 U1948 ( .A1(n1050), .A2(n12), .B1(n1049), .B2(n1510), .ZN(n841) );
  OAI22_X1 U1949 ( .A1(n1469), .A2(n1065), .B1(n1064), .B2(n1510), .ZN(n856)
         );
  OAI22_X1 U1950 ( .A1(n1469), .A2(n1058), .B1(n1057), .B2(n1509), .ZN(n849)
         );
  OAI22_X1 U1951 ( .A1(n1469), .A2(n1148), .B1(n1068), .B2(n1510), .ZN(n678)
         );
  OAI22_X1 U1952 ( .A1(n1469), .A2(n1061), .B1(n1060), .B2(n1510), .ZN(n852)
         );
  OAI22_X1 U1953 ( .A1(n1048), .A2(n12), .B1(n1048), .B2(n1510), .ZN(n664) );
  OAI22_X1 U1954 ( .A1(n1336), .A2(n1064), .B1(n1063), .B2(n1509), .ZN(n855)
         );
  OAI22_X1 U1955 ( .A1(n1469), .A2(n1067), .B1(n1066), .B2(n1509), .ZN(n858)
         );
  OAI22_X1 U1956 ( .A1(n1336), .A2(n1066), .B1(n1065), .B2(n1510), .ZN(n857)
         );
  INV_X1 U1957 ( .A(n1510), .ZN(n665) );
  INV_X1 U1958 ( .A(n1464), .ZN(n173) );
  OAI22_X1 U1959 ( .A1(n985), .A2(n30), .B1(n985), .B2(n1453), .ZN(n655) );
  OAI22_X1 U1960 ( .A1(n1435), .A2(n986), .B1(n985), .B2(n1359), .ZN(n368) );
  OAI22_X1 U1961 ( .A1(n30), .A2(n987), .B1(n986), .B2(n1453), .ZN(n781) );
  OAI22_X1 U1962 ( .A1(n30), .A2(n989), .B1(n988), .B2(n1452), .ZN(n783) );
  OAI22_X1 U1963 ( .A1(n1435), .A2(n990), .B1(n989), .B2(n1453), .ZN(n784) );
  OAI22_X1 U1964 ( .A1(n1435), .A2(n992), .B1(n991), .B2(n1359), .ZN(n786) );
  OAI22_X1 U1965 ( .A1(n1435), .A2(n1003), .B1(n1002), .B2(n1452), .ZN(n797)
         );
  OAI22_X1 U1966 ( .A1(n30), .A2(n988), .B1(n987), .B2(n1359), .ZN(n782) );
  OAI22_X1 U1967 ( .A1(n1435), .A2(n996), .B1(n995), .B2(n1359), .ZN(n790) );
  OAI22_X1 U1968 ( .A1(n1435), .A2(n991), .B1(n990), .B2(n1452), .ZN(n785) );
  OAI22_X1 U1969 ( .A1(n1435), .A2(n999), .B1(n998), .B2(n1359), .ZN(n793) );
  OAI22_X1 U1970 ( .A1(n30), .A2(n995), .B1(n994), .B2(n1453), .ZN(n789) );
  OAI22_X1 U1971 ( .A1(n1435), .A2(n993), .B1(n992), .B2(n1453), .ZN(n787) );
  OAI22_X1 U1972 ( .A1(n30), .A2(n1000), .B1(n999), .B2(n1359), .ZN(n794) );
  OAI22_X1 U1973 ( .A1(n30), .A2(n994), .B1(n993), .B2(n1453), .ZN(n788) );
  OAI22_X1 U1974 ( .A1(n1435), .A2(n1004), .B1(n1003), .B2(n1246), .ZN(n798)
         );
  OAI22_X1 U1975 ( .A1(n1435), .A2(n998), .B1(n997), .B2(n1452), .ZN(n792) );
  OAI22_X1 U1976 ( .A1(n30), .A2(n1002), .B1(n1001), .B2(n1452), .ZN(n796) );
  OAI22_X1 U1977 ( .A1(n1435), .A2(n1145), .B1(n1005), .B2(n1359), .ZN(n675)
         );
  INV_X1 U1978 ( .A(n1452), .ZN(n656) );
  OAI22_X1 U1979 ( .A1(n1435), .A2(n1001), .B1(n1000), .B2(n1452), .ZN(n795)
         );
  OAI21_X1 U1980 ( .B1(n152), .B2(n131), .A(n1379), .ZN(n130) );
  OAI22_X1 U1981 ( .A1(n901), .A2(n1410), .B1(n901), .B2(n1268), .ZN(n643) );
  OAI22_X1 U1982 ( .A1(n1376), .A2(n902), .B1(n901), .B2(n1268), .ZN(n304) );
  OAI22_X1 U1983 ( .A1(n1377), .A2(n903), .B1(n902), .B2(n1268), .ZN(n701) );
  OAI21_X1 U1984 ( .B1(n132), .B2(n128), .A(n129), .ZN(n127) );
  OAI22_X1 U1985 ( .A1(n1376), .A2(n905), .B1(n904), .B2(n1268), .ZN(n703) );
  OAI22_X1 U1986 ( .A1(n1410), .A2(n904), .B1(n903), .B2(n1268), .ZN(n702) );
  OAI22_X1 U1987 ( .A1(n1377), .A2(n906), .B1(n905), .B2(n1268), .ZN(n704) );
  OAI22_X1 U1988 ( .A1(n1410), .A2(n907), .B1(n906), .B2(n1268), .ZN(n705) );
  OAI22_X1 U1989 ( .A1(n1376), .A2(n908), .B1(n907), .B2(n1335), .ZN(n706) );
  OAI22_X1 U1990 ( .A1(n1377), .A2(n909), .B1(n908), .B2(n1335), .ZN(n707) );
  OAI22_X1 U1991 ( .A1(n1410), .A2(n910), .B1(n909), .B2(n1335), .ZN(n708) );
  OAI22_X1 U1992 ( .A1(n1376), .A2(n911), .B1(n910), .B2(n1335), .ZN(n709) );
  OAI22_X1 U1993 ( .A1(n54), .A2(n1141), .B1(n921), .B2(n1335), .ZN(n671) );
  OAI22_X1 U1994 ( .A1(n1410), .A2(n915), .B1(n914), .B2(n1335), .ZN(n713) );
  OAI22_X1 U1995 ( .A1(n1377), .A2(n920), .B1(n919), .B2(n1335), .ZN(n718) );
  OAI22_X1 U1996 ( .A1(n1410), .A2(n912), .B1(n911), .B2(n1335), .ZN(n710) );
  OAI22_X1 U1997 ( .A1(n1377), .A2(n913), .B1(n912), .B2(n1335), .ZN(n711) );
  OAI22_X1 U1998 ( .A1(n1377), .A2(n914), .B1(n913), .B2(n1335), .ZN(n712) );
  OAI22_X1 U1999 ( .A1(n54), .A2(n918), .B1(n917), .B2(n1335), .ZN(n716) );
  OAI22_X1 U2000 ( .A1(n1376), .A2(n919), .B1(n918), .B2(n1335), .ZN(n717) );
  OAI22_X1 U2001 ( .A1(n1376), .A2(n917), .B1(n1269), .B2(n1335), .ZN(n715) );
  INV_X1 U2002 ( .A(n1504), .ZN(n644) );
  OAI22_X1 U2003 ( .A1(n54), .A2(n916), .B1(n915), .B2(n1335), .ZN(n714) );
  INV_X1 U2004 ( .A(n1465), .ZN(n278) );
  INV_X1 U2005 ( .A(n1462), .ZN(n152) );
  OAI22_X1 U2006 ( .A1(n922), .A2(n1471), .B1(n922), .B2(n1291), .ZN(n646) );
  NOR2_X1 U2007 ( .A1(n1465), .A2(n171), .ZN(n164) );
  OAI22_X1 U2008 ( .A1(n1472), .A2(n924), .B1(n923), .B2(n1292), .ZN(n721) );
  OAI22_X1 U2009 ( .A1(n1472), .A2(n923), .B1(n922), .B2(n1291), .ZN(n314) );
  OAI22_X1 U2010 ( .A1(n1471), .A2(n925), .B1(n924), .B2(n1292), .ZN(n722) );
  OAI22_X1 U2011 ( .A1(n1472), .A2(n927), .B1(n926), .B2(n1291), .ZN(n724) );
  OAI22_X1 U2012 ( .A1(n1472), .A2(n926), .B1(n925), .B2(n1292), .ZN(n723) );
  OAI22_X1 U2013 ( .A1(n1472), .A2(n928), .B1(n927), .B2(n1291), .ZN(n725) );
  OAI22_X1 U2014 ( .A1(n1471), .A2(n929), .B1(n928), .B2(n1292), .ZN(n726) );
  OAI22_X1 U2015 ( .A1(n1472), .A2(n930), .B1(n929), .B2(n1291), .ZN(n727) );
  OAI22_X1 U2016 ( .A1(n1471), .A2(n939), .B1(n938), .B2(n1291), .ZN(n736) );
  OAI22_X1 U2017 ( .A1(n1472), .A2(n931), .B1(n930), .B2(n1292), .ZN(n728) );
  OAI22_X1 U2018 ( .A1(n1472), .A2(n933), .B1(n932), .B2(n1292), .ZN(n730) );
  OAI22_X1 U2019 ( .A1(n1471), .A2(n1142), .B1(n942), .B2(n1291), .ZN(n672) );
  OAI22_X1 U2020 ( .A1(n1472), .A2(n940), .B1(n939), .B2(n1292), .ZN(n737) );
  OAI22_X1 U2021 ( .A1(n1471), .A2(n934), .B1(n933), .B2(n1291), .ZN(n731) );
  OAI22_X1 U2022 ( .A1(n1472), .A2(n932), .B1(n931), .B2(n1292), .ZN(n729) );
  OAI22_X1 U2023 ( .A1(n1473), .A2(n936), .B1(n935), .B2(n1508), .ZN(n733) );
  OAI22_X1 U2024 ( .A1(n1472), .A2(n937), .B1(n1297), .B2(n1292), .ZN(n734) );
  OAI22_X1 U2025 ( .A1(n1472), .A2(n941), .B1(n940), .B2(n1292), .ZN(n738) );
  OAI22_X1 U2026 ( .A1(n1473), .A2(n935), .B1(n934), .B2(n1508), .ZN(n732) );
  INV_X1 U2027 ( .A(n1508), .ZN(n647) );
  OAI22_X1 U2028 ( .A1(n1473), .A2(n938), .B1(n937), .B2(n1291), .ZN(n735) );
  OAI22_X1 U2029 ( .A1(n880), .A2(n1461), .B1(n880), .B2(n1432), .ZN(n640) );
  OAI22_X1 U2030 ( .A1(n1461), .A2(n881), .B1(n880), .B2(n1432), .ZN(n298) );
  OAI22_X1 U2031 ( .A1(n1461), .A2(n882), .B1(n881), .B2(n1432), .ZN(n681) );
  OAI22_X1 U2032 ( .A1(n1461), .A2(n883), .B1(n882), .B2(n1432), .ZN(n682) );
  OAI22_X1 U2033 ( .A1(n1461), .A2(n884), .B1(n883), .B2(n1432), .ZN(n683) );
  OAI22_X1 U2034 ( .A1(n1461), .A2(n886), .B1(n885), .B2(n1432), .ZN(n685) );
  OAI22_X1 U2035 ( .A1(n1461), .A2(n885), .B1(n884), .B2(n1432), .ZN(n684) );
  OAI22_X1 U2036 ( .A1(n1461), .A2(n887), .B1(n886), .B2(n1432), .ZN(n686) );
  OAI22_X1 U2037 ( .A1(n1461), .A2(n888), .B1(n887), .B2(n1432), .ZN(n687) );
  OAI22_X1 U2038 ( .A1(n1392), .A2(n889), .B1(n888), .B2(n1432), .ZN(n688) );
  OAI22_X1 U2039 ( .A1(n1392), .A2(n890), .B1(n889), .B2(n1432), .ZN(n689) );
  OAI22_X1 U2040 ( .A1(n1392), .A2(n891), .B1(n890), .B2(n1390), .ZN(n690) );
  OAI22_X1 U2041 ( .A1(n1243), .A2(n892), .B1(n891), .B2(n1390), .ZN(n691) );
  OAI22_X1 U2042 ( .A1(n1243), .A2(n894), .B1(n893), .B2(n1390), .ZN(n693) );
  OAI22_X1 U2043 ( .A1(n60), .A2(n893), .B1(n892), .B2(n58), .ZN(n692) );
  OAI22_X1 U2044 ( .A1(n1243), .A2(n899), .B1(n898), .B2(n1390), .ZN(n698) );
  OAI22_X1 U2045 ( .A1(n1243), .A2(n895), .B1(n894), .B2(n1390), .ZN(n694) );
  OAI22_X1 U2046 ( .A1(n60), .A2(n1393), .B1(n900), .B2(n1460), .ZN(n670) );
  OAI22_X1 U2047 ( .A1(n60), .A2(n898), .B1(n897), .B2(n1390), .ZN(n697) );
  OAI22_X1 U2048 ( .A1(n896), .A2(n60), .B1(n895), .B2(n1460), .ZN(n695) );
  OAI22_X1 U2049 ( .A1(n1243), .A2(n897), .B1(n1390), .B2(n896), .ZN(n696) );
  INV_X1 U2050 ( .A(n1460), .ZN(n641) );
  OAI21_X1 U2051 ( .B1(n174), .B2(n154), .A(n155), .ZN(n153) );
  AOI21_X1 U2052 ( .B1(n194), .B2(n175), .A(n176), .ZN(n174) );
  AOI21_X1 U2053 ( .B1(n153), .B2(n126), .A(n127), .ZN(n125) );
  OAI22_X1 U2054 ( .A1(n30), .A2(n997), .B1(n996), .B2(n1359), .ZN(n791) );
  OAI21_X1 U2055 ( .B1(n181), .B2(n177), .A(n178), .ZN(n176) );
  OAI22_X1 U2056 ( .A1(n943), .A2(n1345), .B1(n943), .B2(n1322), .ZN(n649) );
  OAI22_X1 U2057 ( .A1(n1431), .A2(n944), .B1(n943), .B2(n1323), .ZN(n328) );
  OAI22_X1 U2058 ( .A1(n1345), .A2(n945), .B1(n944), .B2(n1322), .ZN(n741) );
  OAI22_X1 U2059 ( .A1(n1430), .A2(n947), .B1(n946), .B2(n1323), .ZN(n743) );
  OAI22_X1 U2060 ( .A1(n1345), .A2(n946), .B1(n945), .B2(n1322), .ZN(n742) );
  OAI22_X1 U2061 ( .A1(n1430), .A2(n948), .B1(n947), .B2(n1323), .ZN(n744) );
  OAI22_X1 U2062 ( .A1(n1431), .A2(n949), .B1(n948), .B2(n1322), .ZN(n745) );
  OAI22_X1 U2063 ( .A1(n1430), .A2(n952), .B1(n951), .B2(n1323), .ZN(n748) );
  OAI22_X1 U2064 ( .A1(n1431), .A2(n957), .B1(n956), .B2(n1322), .ZN(n753) );
  OAI22_X1 U2065 ( .A1(n1430), .A2(n953), .B1(n952), .B2(n1323), .ZN(n749) );
  OAI22_X1 U2066 ( .A1(n1430), .A2(n956), .B1(n955), .B2(n1323), .ZN(n752) );
  OAI22_X1 U2067 ( .A1(n1430), .A2(n950), .B1(n949), .B2(n1322), .ZN(n746) );
  OAI22_X1 U2068 ( .A1(n1430), .A2(n951), .B1(n950), .B2(n1323), .ZN(n747) );
  OAI22_X1 U2069 ( .A1(n1430), .A2(n958), .B1(n957), .B2(n1323), .ZN(n754) );
  OAI22_X1 U2070 ( .A1(n1431), .A2(n1342), .B1(n963), .B2(n1322), .ZN(n673) );
  OAI22_X1 U2071 ( .A1(n1429), .A2(n955), .B1(n1323), .B2(n954), .ZN(n751) );
  OAI22_X1 U2072 ( .A1(n1431), .A2(n960), .B1(n959), .B2(n1322), .ZN(n756) );
  OAI22_X1 U2073 ( .A1(n1431), .A2(n961), .B1(n960), .B2(n1322), .ZN(n757) );
  OAI22_X1 U2074 ( .A1(n1277), .A2(n1429), .B1(n953), .B2(n1322), .ZN(n750) );
  INV_X1 U2075 ( .A(n1322), .ZN(n650) );
  OAI22_X1 U2076 ( .A1(n1430), .A2(n962), .B1(n961), .B2(n1322), .ZN(n758) );
  OAI22_X1 U2077 ( .A1(n959), .A2(n1430), .B1(n958), .B2(n1322), .ZN(n755) );
  XNOR2_X1 U2078 ( .A(n1470), .B(n67), .ZN(product[29]) );
  XOR2_X1 U2079 ( .A(n1444), .B(n64), .Z(product[32]) );
  XOR2_X1 U2080 ( .A(n1459), .B(n68), .Z(product[28]) );
  AOI21_X1 U2081 ( .B1(n114), .B2(n1491), .A(n111), .ZN(n109) );
  AOI21_X1 U2082 ( .B1(n1470), .B2(n1490), .A(n119), .ZN(n117) );
  OAI21_X1 U2083 ( .B1(n125), .B2(n123), .A(n124), .ZN(n122) );
  OAI22_X1 U2084 ( .A1(n1456), .A2(n1014), .B1(n1013), .B2(n1505), .ZN(n807)
         );
  OAI22_X1 U2085 ( .A1(n1457), .A2(n1007), .B1(n1006), .B2(n1505), .ZN(n394)
         );
  OAI22_X1 U2086 ( .A1(n1457), .A2(n1012), .B1(n1011), .B2(n1505), .ZN(n805)
         );
  OAI22_X1 U2087 ( .A1(n1006), .A2(n1457), .B1(n1006), .B2(n1505), .ZN(n658)
         );
  OAI22_X1 U2088 ( .A1(n1456), .A2(n1021), .B1(n1505), .B2(n1020), .ZN(n814)
         );
  OAI22_X1 U2089 ( .A1(n1456), .A2(n1024), .B1(n1023), .B2(n1505), .ZN(n817)
         );
  OAI22_X1 U2090 ( .A1(n1456), .A2(n1010), .B1(n1009), .B2(n1505), .ZN(n803)
         );
  OAI22_X1 U2091 ( .A1(n1456), .A2(n1008), .B1(n1007), .B2(n1505), .ZN(n801)
         );
  OAI22_X1 U2092 ( .A1(n1457), .A2(n1015), .B1(n1014), .B2(n1505), .ZN(n808)
         );
  OAI22_X1 U2093 ( .A1(n1456), .A2(n1009), .B1(n1008), .B2(n1505), .ZN(n802)
         );
  OAI22_X1 U2094 ( .A1(n1456), .A2(n1146), .B1(n1026), .B2(n1505), .ZN(n676)
         );
  OAI22_X1 U2095 ( .A1(n1457), .A2(n1013), .B1(n1012), .B2(n1505), .ZN(n806)
         );
  OAI22_X1 U2096 ( .A1(n1457), .A2(n1025), .B1(n1024), .B2(n1505), .ZN(n818)
         );
  OAI22_X1 U2097 ( .A1(n1456), .A2(n1019), .B1(n1018), .B2(n1505), .ZN(n812)
         );
  OAI22_X1 U2098 ( .A1(n1456), .A2(n1020), .B1(n1019), .B2(n1505), .ZN(n813)
         );
  OAI22_X1 U2099 ( .A1(n1457), .A2(n1018), .B1(n1017), .B2(n1505), .ZN(n811)
         );
  OAI22_X1 U2100 ( .A1(n1456), .A2(n1011), .B1(n1010), .B2(n1505), .ZN(n804)
         );
  OAI22_X1 U2101 ( .A1(n1457), .A2(n1017), .B1(n1016), .B2(n1505), .ZN(n810)
         );
  OAI22_X1 U2102 ( .A1(n1457), .A2(n1023), .B1(n1022), .B2(n1505), .ZN(n816)
         );
  OAI22_X1 U2103 ( .A1(n1456), .A2(n1016), .B1(n1015), .B2(n1505), .ZN(n809)
         );
  OAI22_X1 U2104 ( .A1(n1457), .A2(n1022), .B1(n1021), .B2(n1505), .ZN(n815)
         );
  INV_X1 U2105 ( .A(n1505), .ZN(n659) );
  XNOR2_X1 U2106 ( .A(n1442), .B(n65), .ZN(product[31]) );
  XNOR2_X1 U2107 ( .A(n1463), .B(n63), .ZN(product[33]) );
  XOR2_X1 U2108 ( .A(n117), .B(n66), .Z(product[30]) );
  INV_X1 U2109 ( .A(n101), .ZN(n264) );
  AOI21_X1 U2110 ( .B1(n106), .B2(n1493), .A(n103), .ZN(n101) );
  OAI21_X1 U2111 ( .B1(n1474), .B2(n115), .A(n116), .ZN(n114) );
  OAI22_X1 U2112 ( .A1(n1279), .A2(n1039), .B1(n1038), .B2(n1507), .ZN(n831)
         );
  OAI22_X1 U2113 ( .A1(n1279), .A2(n1031), .B1(n1030), .B2(n1507), .ZN(n823)
         );
  OAI22_X1 U2114 ( .A1(n1279), .A2(n1041), .B1(n1040), .B2(n1346), .ZN(n833)
         );
  OAI22_X1 U2115 ( .A1(n1279), .A2(n1032), .B1(n1031), .B2(n1346), .ZN(n824)
         );
  OAI22_X1 U2116 ( .A1(n1408), .A2(n1034), .B1(n1033), .B2(n1346), .ZN(n826)
         );
  OAI22_X1 U2117 ( .A1(n1408), .A2(n1045), .B1(n1044), .B2(n1346), .ZN(n837)
         );
  OAI22_X1 U2118 ( .A1(n1408), .A2(n1038), .B1(n1037), .B2(n1346), .ZN(n830)
         );
  OAI22_X1 U2119 ( .A1(n1408), .A2(n1044), .B1(n1043), .B2(n1346), .ZN(n836)
         );
  OAI22_X1 U2120 ( .A1(n1279), .A2(n1028), .B1(n1027), .B2(n1346), .ZN(n424)
         );
  OAI22_X1 U2121 ( .A1(n1408), .A2(n1040), .B1(n1039), .B2(n1507), .ZN(n832)
         );
  OAI22_X1 U2122 ( .A1(n1279), .A2(n1033), .B1(n1032), .B2(n1507), .ZN(n825)
         );
  OAI22_X1 U2123 ( .A1(n1408), .A2(n1037), .B1(n1036), .B2(n1507), .ZN(n829)
         );
  OAI22_X1 U2124 ( .A1(n1279), .A2(n1147), .B1(n1047), .B2(n1507), .ZN(n677)
         );
  OAI22_X1 U2125 ( .A1(n1027), .A2(n1279), .B1(n1027), .B2(n1507), .ZN(n661)
         );
  OAI22_X1 U2126 ( .A1(n1408), .A2(n1030), .B1(n1029), .B2(n1346), .ZN(n822)
         );
  OAI22_X1 U2127 ( .A1(n1328), .A2(n1408), .B1(n1028), .B2(n1507), .ZN(n821)
         );
  OAI22_X1 U2128 ( .A1(n1279), .A2(n1036), .B1(n1035), .B2(n1507), .ZN(n828)
         );
  OAI22_X1 U2129 ( .A1(n1408), .A2(n1043), .B1(n1042), .B2(n1346), .ZN(n835)
         );
  OAI22_X1 U2130 ( .A1(n1408), .A2(n1042), .B1(n1041), .B2(n1507), .ZN(n834)
         );
  OAI22_X1 U2131 ( .A1(n1279), .A2(n1035), .B1(n1034), .B2(n1346), .ZN(n827)
         );
  OAI22_X1 U2132 ( .A1(n1408), .A2(n1046), .B1(n1045), .B2(n1346), .ZN(n838)
         );
  INV_X1 U2133 ( .A(n1507), .ZN(n662) );
  OAI21_X1 U2134 ( .B1(n109), .B2(n107), .A(n108), .ZN(n106) );
endmodule


module mac_4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n34, n35, n36, n37, n38, n39, n40, n41, n43, n45, n46, n47,
         n48, n49, n51, n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65,
         n67, n69, n70, n71, n72, n73, n75, n77, n78, n79, n80, n81, n83, n85,
         n86, n87, n88, n89, n91, n93, n94, n95, n96, n97, n99, n101, n102,
         n103, n104, n105, n107, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n119, n121, n122, n124, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n184, n185, n187, n189, n191,
         n193, n195, n197, n199, n201, n203, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406;

  FA_X1 U3 ( .A(B[38]), .B(A[38]), .CI(n35), .CO(n34), .S(SUM[38]) );
  FA_X1 U4 ( .A(B[37]), .B(A[37]), .CI(n36), .CO(n35), .S(SUM[37]) );
  CLKBUF_X1 U254 ( .A(n131), .Z(n344) );
  CLKBUF_X1 U255 ( .A(n115), .Z(n345) );
  OR2_X1 U256 ( .A1(B[0]), .A2(A[0]), .ZN(n346) );
  CLKBUF_X1 U257 ( .A(n37), .Z(n347) );
  XOR2_X1 U258 ( .A(B[36]), .B(A[36]), .Z(n348) );
  XOR2_X1 U259 ( .A(n347), .B(n348), .Z(SUM[36]) );
  NAND2_X1 U260 ( .A1(n37), .A2(B[36]), .ZN(n349) );
  NAND2_X1 U261 ( .A1(n37), .A2(A[36]), .ZN(n350) );
  NAND2_X1 U262 ( .A1(B[36]), .A2(A[36]), .ZN(n351) );
  NAND3_X1 U263 ( .A1(n349), .A2(n350), .A3(n351), .ZN(n36) );
  CLKBUF_X1 U264 ( .A(n185), .Z(n352) );
  NAND3_X1 U265 ( .A1(n371), .A2(n372), .A3(n373), .ZN(n353) );
  NAND3_X1 U266 ( .A1(n371), .A2(n372), .A3(n373), .ZN(n354) );
  XOR2_X1 U267 ( .A(B[35]), .B(A[35]), .Z(n355) );
  XOR2_X1 U268 ( .A(n354), .B(n355), .Z(SUM[35]) );
  NAND2_X1 U269 ( .A1(n353), .A2(B[35]), .ZN(n356) );
  NAND2_X1 U270 ( .A1(n38), .A2(A[35]), .ZN(n357) );
  NAND2_X1 U271 ( .A1(B[35]), .A2(A[35]), .ZN(n358) );
  NAND3_X1 U272 ( .A1(n356), .A2(n357), .A3(n358), .ZN(n37) );
  NAND3_X1 U273 ( .A1(n378), .A2(n379), .A3(n380), .ZN(n359) );
  CLKBUF_X1 U274 ( .A(n94), .Z(n360) );
  NAND3_X1 U275 ( .A1(n386), .A2(n387), .A3(n388), .ZN(n361) );
  NAND3_X1 U276 ( .A1(n386), .A2(n387), .A3(n388), .ZN(n362) );
  AOI21_X1 U277 ( .B1(n150), .B2(n114), .A(n345), .ZN(n363) );
  AOI21_X1 U278 ( .B1(n150), .B2(n114), .A(n115), .ZN(n113) );
  AOI21_X1 U279 ( .B1(n360), .B2(n398), .A(n91), .ZN(n364) );
  AOI21_X1 U280 ( .B1(n94), .B2(n398), .A(n91), .ZN(n89) );
  NOR2_X1 U281 ( .A1(B[3]), .A2(A[3]), .ZN(n365) );
  AOI21_X1 U282 ( .B1(n130), .B2(n143), .A(n344), .ZN(n366) );
  CLKBUF_X1 U283 ( .A(n54), .Z(n367) );
  AOI21_X1 U284 ( .B1(n367), .B2(n404), .A(n51), .ZN(n368) );
  CLKBUF_X1 U285 ( .A(n102), .Z(n369) );
  XOR2_X1 U286 ( .A(B[34]), .B(A[34]), .Z(n370) );
  XOR2_X1 U287 ( .A(n359), .B(n370), .Z(SUM[34]) );
  NAND2_X1 U288 ( .A1(n359), .A2(B[34]), .ZN(n371) );
  NAND2_X1 U289 ( .A1(n39), .A2(A[34]), .ZN(n372) );
  NAND2_X1 U290 ( .A1(B[34]), .A2(A[34]), .ZN(n373) );
  NAND3_X1 U291 ( .A1(n371), .A2(n372), .A3(n373), .ZN(n38) );
  CLKBUF_X1 U292 ( .A(n46), .Z(n374) );
  AOI21_X1 U293 ( .B1(n369), .B2(n400), .A(n99), .ZN(n375) );
  CLKBUF_X1 U294 ( .A(n110), .Z(n376) );
  AOI21_X1 U295 ( .B1(n54), .B2(n404), .A(n51), .ZN(n49) );
  XOR2_X1 U296 ( .A(B[33]), .B(A[33]), .Z(n377) );
  XOR2_X1 U297 ( .A(n362), .B(n377), .Z(SUM[33]) );
  NAND2_X1 U298 ( .A1(n361), .A2(B[33]), .ZN(n378) );
  NAND2_X1 U299 ( .A1(n40), .A2(A[33]), .ZN(n379) );
  NAND2_X1 U300 ( .A1(B[33]), .A2(A[33]), .ZN(n380) );
  NAND3_X1 U301 ( .A1(n378), .A2(n379), .A3(n380), .ZN(n39) );
  CLKBUF_X1 U302 ( .A(n62), .Z(n381) );
  AOI21_X1 U303 ( .B1(n376), .B2(n399), .A(n107), .ZN(n382) );
  CLKBUF_X1 U304 ( .A(n70), .Z(n383) );
  CLKBUF_X1 U305 ( .A(n78), .Z(n384) );
  XOR2_X1 U306 ( .A(B[32]), .B(A[32]), .Z(n385) );
  XOR2_X1 U307 ( .A(n352), .B(n385), .Z(SUM[32]) );
  NAND2_X1 U308 ( .A1(n185), .A2(B[32]), .ZN(n386) );
  NAND2_X1 U309 ( .A1(n185), .A2(A[32]), .ZN(n387) );
  NAND2_X1 U310 ( .A1(B[32]), .A2(A[32]), .ZN(n388) );
  NAND3_X1 U311 ( .A1(n386), .A2(n387), .A3(n388), .ZN(n40) );
  AOI21_X1 U312 ( .B1(n384), .B2(n401), .A(n75), .ZN(n389) );
  AOI21_X1 U313 ( .B1(n383), .B2(n402), .A(n67), .ZN(n390) );
  CLKBUF_X1 U314 ( .A(n86), .Z(n391) );
  AOI21_X1 U315 ( .B1(n381), .B2(n403), .A(n59), .ZN(n392) );
  AOI21_X1 U316 ( .B1(n391), .B2(n397), .A(n83), .ZN(n393) );
  NOR2_X2 U317 ( .A1(B[9]), .A2(A[9]), .ZN(n144) );
  NOR2_X2 U318 ( .A1(B[11]), .A2(A[11]), .ZN(n132) );
  INV_X1 U319 ( .A(n150), .ZN(n149) );
  OAI21_X1 U320 ( .B1(n149), .B2(n140), .A(n141), .ZN(n139) );
  INV_X1 U321 ( .A(n143), .ZN(n141) );
  INV_X1 U322 ( .A(n142), .ZN(n140) );
  NAND2_X1 U323 ( .A1(n142), .A2(n130), .ZN(n128) );
  AOI21_X1 U324 ( .B1(n170), .B2(n161), .A(n162), .ZN(n160) );
  INV_X1 U325 ( .A(n171), .ZN(n170) );
  INV_X1 U326 ( .A(n180), .ZN(n179) );
  OAI21_X1 U327 ( .B1(n163), .B2(n169), .A(n164), .ZN(n162) );
  INV_X1 U328 ( .A(n69), .ZN(n67) );
  INV_X1 U329 ( .A(n61), .ZN(n59) );
  INV_X1 U330 ( .A(n53), .ZN(n51) );
  AOI21_X1 U331 ( .B1(n110), .B2(n399), .A(n107), .ZN(n105) );
  INV_X1 U332 ( .A(n109), .ZN(n107) );
  AOI21_X1 U333 ( .B1(n172), .B2(n180), .A(n173), .ZN(n171) );
  AOI21_X1 U334 ( .B1(n86), .B2(n397), .A(n83), .ZN(n81) );
  INV_X1 U335 ( .A(n85), .ZN(n83) );
  AOI21_X1 U336 ( .B1(n78), .B2(n401), .A(n75), .ZN(n73) );
  INV_X1 U337 ( .A(n77), .ZN(n75) );
  INV_X1 U338 ( .A(n93), .ZN(n91) );
  AOI21_X1 U339 ( .B1(n102), .B2(n400), .A(n99), .ZN(n97) );
  INV_X1 U340 ( .A(n101), .ZN(n99) );
  OAI21_X1 U341 ( .B1(n181), .B2(n184), .A(n182), .ZN(n180) );
  OAI21_X1 U342 ( .B1(n144), .B2(n148), .A(n145), .ZN(n143) );
  NOR2_X1 U343 ( .A1(n137), .A2(n132), .ZN(n130) );
  OAI21_X1 U344 ( .B1(n171), .B2(n151), .A(n152), .ZN(n150) );
  NAND2_X1 U345 ( .A1(n161), .A2(n153), .ZN(n151) );
  AOI21_X1 U346 ( .B1(n153), .B2(n162), .A(n154), .ZN(n152) );
  NAND2_X1 U347 ( .A1(n197), .A2(n88), .ZN(n13) );
  INV_X1 U348 ( .A(n87), .ZN(n197) );
  NAND2_X1 U349 ( .A1(n199), .A2(n96), .ZN(n15) );
  INV_X1 U350 ( .A(n95), .ZN(n199) );
  NOR2_X1 U351 ( .A1(n128), .A2(n116), .ZN(n114) );
  NAND2_X1 U352 ( .A1(n395), .A2(n396), .ZN(n116) );
  NOR2_X1 U353 ( .A1(n147), .A2(n144), .ZN(n142) );
  AOI21_X1 U354 ( .B1(n130), .B2(n143), .A(n131), .ZN(n129) );
  OAI21_X1 U355 ( .B1(n132), .B2(n138), .A(n133), .ZN(n131) );
  INV_X1 U356 ( .A(n126), .ZN(n124) );
  AOI21_X1 U357 ( .B1(n396), .B2(n124), .A(n119), .ZN(n117) );
  INV_X1 U358 ( .A(n121), .ZN(n119) );
  NAND2_X1 U359 ( .A1(n187), .A2(n48), .ZN(n3) );
  INV_X1 U360 ( .A(n47), .ZN(n187) );
  NAND2_X1 U361 ( .A1(n189), .A2(n56), .ZN(n5) );
  INV_X1 U362 ( .A(n55), .ZN(n189) );
  NAND2_X1 U363 ( .A1(n191), .A2(n64), .ZN(n7) );
  INV_X1 U364 ( .A(n63), .ZN(n191) );
  NAND2_X1 U365 ( .A1(n193), .A2(n72), .ZN(n9) );
  INV_X1 U366 ( .A(n71), .ZN(n193) );
  NAND2_X1 U367 ( .A1(n195), .A2(n80), .ZN(n11) );
  INV_X1 U368 ( .A(n79), .ZN(n195) );
  NAND2_X1 U369 ( .A1(n405), .A2(n45), .ZN(n2) );
  NAND2_X1 U370 ( .A1(n404), .A2(n53), .ZN(n4) );
  NAND2_X1 U371 ( .A1(n403), .A2(n61), .ZN(n6) );
  NAND2_X1 U372 ( .A1(n402), .A2(n69), .ZN(n8) );
  NAND2_X1 U373 ( .A1(n401), .A2(n77), .ZN(n10) );
  XNOR2_X1 U374 ( .A(n391), .B(n12), .ZN(SUM[21]) );
  NAND2_X1 U375 ( .A1(n397), .A2(n85), .ZN(n12) );
  NAND2_X1 U376 ( .A1(n398), .A2(n93), .ZN(n14) );
  NAND2_X1 U377 ( .A1(n400), .A2(n101), .ZN(n16) );
  XOR2_X1 U378 ( .A(n382), .B(n17), .Z(SUM[16]) );
  NAND2_X1 U379 ( .A1(n201), .A2(n104), .ZN(n17) );
  INV_X1 U380 ( .A(n103), .ZN(n201) );
  XOR2_X1 U381 ( .A(n122), .B(n20), .Z(SUM[13]) );
  NAND2_X1 U382 ( .A1(n396), .A2(n121), .ZN(n20) );
  AOI21_X1 U383 ( .B1(n127), .B2(n395), .A(n124), .ZN(n122) );
  XNOR2_X1 U384 ( .A(n127), .B(n21), .ZN(SUM[12]) );
  NAND2_X1 U385 ( .A1(n395), .A2(n126), .ZN(n21) );
  XOR2_X1 U386 ( .A(n134), .B(n22), .Z(SUM[11]) );
  NAND2_X1 U387 ( .A1(n206), .A2(n133), .ZN(n22) );
  AOI21_X1 U388 ( .B1(n139), .B2(n207), .A(n136), .ZN(n134) );
  NAND2_X1 U389 ( .A1(n203), .A2(n112), .ZN(n19) );
  INV_X1 U390 ( .A(n111), .ZN(n203) );
  XOR2_X1 U391 ( .A(n165), .B(n28), .Z(SUM[5]) );
  NAND2_X1 U392 ( .A1(n212), .A2(n164), .ZN(n28) );
  AOI21_X1 U393 ( .B1(n170), .B2(n213), .A(n167), .ZN(n165) );
  INV_X1 U394 ( .A(n137), .ZN(n207) );
  INV_X1 U395 ( .A(n168), .ZN(n213) );
  XNOR2_X1 U396 ( .A(n146), .B(n24), .ZN(SUM[9]) );
  NAND2_X1 U397 ( .A1(n208), .A2(n145), .ZN(n24) );
  OAI21_X1 U398 ( .B1(n149), .B2(n147), .A(n148), .ZN(n146) );
  INV_X1 U399 ( .A(n132), .ZN(n206) );
  INV_X1 U400 ( .A(n138), .ZN(n136) );
  INV_X1 U401 ( .A(n169), .ZN(n167) );
  INV_X1 U402 ( .A(n144), .ZN(n208) );
  XOR2_X1 U403 ( .A(n160), .B(n27), .Z(SUM[6]) );
  NAND2_X1 U404 ( .A1(n211), .A2(n159), .ZN(n27) );
  INV_X1 U405 ( .A(n158), .ZN(n211) );
  XNOR2_X1 U406 ( .A(n170), .B(n29), .ZN(SUM[4]) );
  NAND2_X1 U407 ( .A1(n213), .A2(n169), .ZN(n29) );
  XNOR2_X1 U408 ( .A(n176), .B(n30), .ZN(SUM[3]) );
  NAND2_X1 U409 ( .A1(n214), .A2(n175), .ZN(n30) );
  OAI21_X1 U410 ( .B1(n179), .B2(n177), .A(n178), .ZN(n176) );
  XOR2_X1 U411 ( .A(n179), .B(n31), .Z(SUM[2]) );
  NAND2_X1 U412 ( .A1(n215), .A2(n178), .ZN(n31) );
  INV_X1 U413 ( .A(n177), .ZN(n215) );
  XOR2_X1 U414 ( .A(n32), .B(n184), .Z(SUM[1]) );
  NAND2_X1 U415 ( .A1(n216), .A2(n182), .ZN(n32) );
  INV_X1 U416 ( .A(n181), .ZN(n216) );
  AND2_X1 U417 ( .A1(n346), .A2(n184), .ZN(SUM[0]) );
  NAND2_X1 U418 ( .A1(n399), .A2(n109), .ZN(n18) );
  XNOR2_X1 U419 ( .A(n139), .B(n23), .ZN(SUM[10]) );
  NAND2_X1 U420 ( .A1(n207), .A2(n138), .ZN(n23) );
  XOR2_X1 U421 ( .A(n149), .B(n25), .Z(SUM[8]) );
  NAND2_X1 U422 ( .A1(n209), .A2(n148), .ZN(n25) );
  INV_X1 U423 ( .A(n147), .ZN(n209) );
  XNOR2_X1 U424 ( .A(n157), .B(n26), .ZN(SUM[7]) );
  NAND2_X1 U425 ( .A1(n210), .A2(n156), .ZN(n26) );
  OAI21_X1 U426 ( .B1(n160), .B2(n158), .A(n159), .ZN(n157) );
  NOR2_X1 U427 ( .A1(B[8]), .A2(A[8]), .ZN(n147) );
  NAND2_X1 U428 ( .A1(B[0]), .A2(A[0]), .ZN(n184) );
  NOR2_X1 U429 ( .A1(B[5]), .A2(A[5]), .ZN(n163) );
  OR2_X1 U430 ( .A1(B[12]), .A2(A[12]), .ZN(n395) );
  OR2_X1 U431 ( .A1(B[13]), .A2(A[13]), .ZN(n396) );
  NOR2_X1 U432 ( .A1(B[6]), .A2(A[6]), .ZN(n158) );
  NOR2_X1 U433 ( .A1(B[2]), .A2(A[2]), .ZN(n177) );
  NOR2_X1 U434 ( .A1(B[7]), .A2(A[7]), .ZN(n155) );
  NOR2_X1 U435 ( .A1(B[3]), .A2(A[3]), .ZN(n174) );
  NAND2_X1 U436 ( .A1(B[11]), .A2(A[11]), .ZN(n133) );
  NOR2_X1 U437 ( .A1(B[10]), .A2(A[10]), .ZN(n137) );
  NOR2_X1 U438 ( .A1(B[1]), .A2(A[1]), .ZN(n181) );
  NAND2_X1 U439 ( .A1(B[8]), .A2(A[8]), .ZN(n148) );
  NAND2_X1 U440 ( .A1(B[10]), .A2(A[10]), .ZN(n138) );
  NAND2_X1 U441 ( .A1(B[2]), .A2(A[2]), .ZN(n178) );
  NAND2_X1 U442 ( .A1(B[6]), .A2(A[6]), .ZN(n159) );
  NAND2_X1 U443 ( .A1(B[4]), .A2(A[4]), .ZN(n169) );
  NAND2_X1 U444 ( .A1(B[1]), .A2(A[1]), .ZN(n182) );
  NAND2_X1 U445 ( .A1(B[9]), .A2(A[9]), .ZN(n145) );
  INV_X1 U446 ( .A(n45), .ZN(n43) );
  NOR2_X1 U447 ( .A1(B[4]), .A2(A[4]), .ZN(n168) );
  NOR2_X1 U448 ( .A1(B[20]), .A2(A[20]), .ZN(n87) );
  NOR2_X1 U449 ( .A1(B[18]), .A2(A[18]), .ZN(n95) );
  NOR2_X1 U450 ( .A1(B[14]), .A2(A[14]), .ZN(n111) );
  NOR2_X1 U451 ( .A1(B[16]), .A2(A[16]), .ZN(n103) );
  NOR2_X1 U452 ( .A1(B[30]), .A2(A[30]), .ZN(n47) );
  NOR2_X1 U453 ( .A1(B[28]), .A2(A[28]), .ZN(n55) );
  NOR2_X1 U454 ( .A1(B[26]), .A2(A[26]), .ZN(n63) );
  NOR2_X1 U455 ( .A1(B[24]), .A2(A[24]), .ZN(n71) );
  NOR2_X1 U456 ( .A1(B[22]), .A2(A[22]), .ZN(n79) );
  OR2_X1 U457 ( .A1(B[21]), .A2(A[21]), .ZN(n397) );
  OR2_X1 U458 ( .A1(B[19]), .A2(A[19]), .ZN(n398) );
  OR2_X1 U459 ( .A1(B[15]), .A2(A[15]), .ZN(n399) );
  OR2_X1 U460 ( .A1(B[17]), .A2(A[17]), .ZN(n400) );
  OR2_X1 U461 ( .A1(B[23]), .A2(A[23]), .ZN(n401) );
  NAND2_X1 U462 ( .A1(B[21]), .A2(A[21]), .ZN(n85) );
  NAND2_X1 U463 ( .A1(B[12]), .A2(A[12]), .ZN(n126) );
  NAND2_X1 U464 ( .A1(B[19]), .A2(A[19]), .ZN(n93) );
  NAND2_X1 U465 ( .A1(B[13]), .A2(A[13]), .ZN(n121) );
  NAND2_X1 U466 ( .A1(B[15]), .A2(A[15]), .ZN(n109) );
  NAND2_X1 U467 ( .A1(B[17]), .A2(A[17]), .ZN(n101) );
  NAND2_X1 U468 ( .A1(B[23]), .A2(A[23]), .ZN(n77) );
  NAND2_X1 U469 ( .A1(B[25]), .A2(A[25]), .ZN(n69) );
  NAND2_X1 U470 ( .A1(B[27]), .A2(A[27]), .ZN(n61) );
  NAND2_X1 U471 ( .A1(B[29]), .A2(A[29]), .ZN(n53) );
  NAND2_X1 U472 ( .A1(B[31]), .A2(A[31]), .ZN(n45) );
  NAND2_X1 U473 ( .A1(B[20]), .A2(A[20]), .ZN(n88) );
  NAND2_X1 U474 ( .A1(B[18]), .A2(A[18]), .ZN(n96) );
  NAND2_X1 U475 ( .A1(B[14]), .A2(A[14]), .ZN(n112) );
  NAND2_X1 U476 ( .A1(B[16]), .A2(A[16]), .ZN(n104) );
  NAND2_X1 U477 ( .A1(B[30]), .A2(A[30]), .ZN(n48) );
  NAND2_X1 U478 ( .A1(B[28]), .A2(A[28]), .ZN(n56) );
  NAND2_X1 U479 ( .A1(B[26]), .A2(A[26]), .ZN(n64) );
  NAND2_X1 U480 ( .A1(B[24]), .A2(A[24]), .ZN(n72) );
  NAND2_X1 U481 ( .A1(B[22]), .A2(A[22]), .ZN(n80) );
  OR2_X1 U482 ( .A1(B[25]), .A2(A[25]), .ZN(n402) );
  OR2_X1 U483 ( .A1(B[27]), .A2(A[27]), .ZN(n403) );
  OR2_X1 U484 ( .A1(B[29]), .A2(A[29]), .ZN(n404) );
  OR2_X1 U485 ( .A1(B[31]), .A2(A[31]), .ZN(n405) );
  XNOR2_X1 U486 ( .A(n34), .B(n406), .ZN(SUM[39]) );
  XNOR2_X1 U487 ( .A(A[39]), .B(B[39]), .ZN(n406) );
  OAI21_X1 U488 ( .B1(n89), .B2(n87), .A(n88), .ZN(n86) );
  XOR2_X1 U489 ( .A(n364), .B(n13), .Z(SUM[20]) );
  XNOR2_X1 U490 ( .A(n360), .B(n14), .ZN(SUM[19]) );
  OAI21_X1 U491 ( .B1(n97), .B2(n95), .A(n96), .ZN(n94) );
  XOR2_X1 U492 ( .A(n375), .B(n15), .Z(SUM[18]) );
  XNOR2_X1 U493 ( .A(n369), .B(n16), .ZN(SUM[17]) );
  OAI21_X1 U494 ( .B1(n105), .B2(n103), .A(n104), .ZN(n102) );
  XNOR2_X1 U495 ( .A(n384), .B(n10), .ZN(SUM[23]) );
  XNOR2_X1 U496 ( .A(n376), .B(n18), .ZN(SUM[15]) );
  INV_X1 U497 ( .A(n41), .ZN(n185) );
  XNOR2_X1 U498 ( .A(n374), .B(n2), .ZN(SUM[31]) );
  XOR2_X1 U499 ( .A(n393), .B(n11), .Z(SUM[22]) );
  XOR2_X1 U500 ( .A(n363), .B(n19), .Z(SUM[14]) );
  XOR2_X1 U501 ( .A(n368), .B(n3), .Z(SUM[30]) );
  AOI21_X1 U502 ( .B1(n46), .B2(n405), .A(n43), .ZN(n41) );
  OAI21_X1 U503 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  OAI21_X1 U504 ( .B1(n81), .B2(n79), .A(n80), .ZN(n78) );
  OAI21_X1 U505 ( .B1(n113), .B2(n111), .A(n112), .ZN(n110) );
  XNOR2_X1 U506 ( .A(n367), .B(n4), .ZN(SUM[29]) );
  INV_X1 U507 ( .A(n155), .ZN(n210) );
  NOR2_X1 U508 ( .A1(n158), .A2(n155), .ZN(n153) );
  OAI21_X1 U509 ( .B1(n155), .B2(n159), .A(n156), .ZN(n154) );
  NAND2_X1 U510 ( .A1(B[7]), .A2(A[7]), .ZN(n156) );
  XOR2_X1 U511 ( .A(n392), .B(n5), .Z(SUM[28]) );
  INV_X1 U512 ( .A(n163), .ZN(n212) );
  OAI21_X1 U513 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  AOI21_X1 U514 ( .B1(n62), .B2(n403), .A(n59), .ZN(n57) );
  NOR2_X1 U515 ( .A1(n168), .A2(n163), .ZN(n161) );
  NAND2_X1 U516 ( .A1(B[5]), .A2(A[5]), .ZN(n164) );
  XNOR2_X1 U517 ( .A(n381), .B(n6), .ZN(SUM[27]) );
  XNOR2_X1 U518 ( .A(n383), .B(n8), .ZN(SUM[25]) );
  INV_X1 U519 ( .A(n365), .ZN(n214) );
  AOI21_X1 U520 ( .B1(n70), .B2(n402), .A(n67), .ZN(n65) );
  NOR2_X1 U521 ( .A1(n177), .A2(n365), .ZN(n172) );
  OAI21_X1 U522 ( .B1(n174), .B2(n178), .A(n175), .ZN(n173) );
  NAND2_X1 U523 ( .A1(B[3]), .A2(A[3]), .ZN(n175) );
  XOR2_X1 U524 ( .A(n390), .B(n7), .Z(SUM[26]) );
  XOR2_X1 U525 ( .A(n389), .B(n9), .Z(SUM[24]) );
  OAI21_X1 U526 ( .B1(n149), .B2(n128), .A(n366), .ZN(n127) );
  OAI21_X1 U527 ( .B1(n65), .B2(n63), .A(n64), .ZN(n62) );
  OAI21_X1 U528 ( .B1(n73), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U529 ( .B1(n129), .B2(n116), .A(n117), .ZN(n115) );
endmodule


module mac_4 ( clk, clear_acc, a, b, mac_out );
  input [19:0] a;
  input [19:0] b;
  output [39:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, n2, n3;
  wire   [39:0] mul;
  wire   [39:0] pipeline;
  wire   [39:0] sum;

  DFF_X1 \pipeline_reg[38]  ( .D(mul[38]), .CK(clk), .Q(pipeline[38]) );
  DFF_X1 \pipeline_reg[37]  ( .D(mul[37]), .CK(clk), .Q(pipeline[37]) );
  DFF_X1 \pipeline_reg[36]  ( .D(mul[36]), .CK(clk), .Q(pipeline[36]) );
  DFF_X1 \pipeline_reg[35]  ( .D(mul[35]), .CK(clk), .Q(pipeline[35]) );
  DFF_X1 \pipeline_reg[34]  ( .D(mul[34]), .CK(clk), .Q(pipeline[34]) );
  DFF_X1 \pipeline_reg[33]  ( .D(mul[33]), .CK(clk), .Q(pipeline[33]) );
  DFF_X1 \pipeline_reg[32]  ( .D(mul[32]), .CK(clk), .Q(pipeline[32]) );
  DFF_X1 \pipeline_reg[31]  ( .D(mul[31]), .CK(clk), .Q(pipeline[31]) );
  DFF_X1 \pipeline_reg[30]  ( .D(mul[30]), .CK(clk), .Q(pipeline[30]) );
  DFF_X1 \pipeline_reg[29]  ( .D(mul[29]), .CK(clk), .Q(pipeline[29]) );
  DFF_X1 \pipeline_reg[28]  ( .D(mul[28]), .CK(clk), .Q(pipeline[28]) );
  DFF_X1 \pipeline_reg[27]  ( .D(mul[27]), .CK(clk), .Q(pipeline[27]) );
  DFF_X1 \pipeline_reg[26]  ( .D(mul[26]), .CK(clk), .Q(pipeline[26]) );
  DFF_X1 \pipeline_reg[25]  ( .D(mul[25]), .CK(clk), .Q(pipeline[25]) );
  DFF_X1 \pipeline_reg[24]  ( .D(mul[24]), .CK(clk), .Q(pipeline[24]) );
  DFF_X1 \pipeline_reg[23]  ( .D(mul[23]), .CK(clk), .Q(pipeline[23]) );
  DFF_X1 \pipeline_reg[22]  ( .D(mul[22]), .CK(clk), .Q(pipeline[22]) );
  DFF_X1 \pipeline_reg[21]  ( .D(mul[21]), .CK(clk), .Q(pipeline[21]) );
  DFF_X1 \pipeline_reg[20]  ( .D(mul[20]), .CK(clk), .Q(pipeline[20]) );
  DFF_X1 \pipeline_reg[19]  ( .D(mul[19]), .CK(clk), .Q(pipeline[19]) );
  DFF_X1 \pipeline_reg[18]  ( .D(mul[18]), .CK(clk), .Q(pipeline[18]) );
  DFF_X1 \pipeline_reg[17]  ( .D(mul[17]), .CK(clk), .Q(pipeline[17]) );
  DFF_X1 \pipeline_reg[16]  ( .D(mul[16]), .CK(clk), .Q(pipeline[16]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \mac_out_reg[16]  ( .D(N19), .CK(clk), .Q(mac_out[16]) );
  DFF_X1 \mac_out_reg[17]  ( .D(N20), .CK(clk), .Q(mac_out[17]) );
  DFF_X1 \mac_out_reg[18]  ( .D(N21), .CK(clk), .Q(mac_out[18]) );
  DFF_X1 \mac_out_reg[19]  ( .D(N22), .CK(clk), .Q(mac_out[19]) );
  DFF_X1 \mac_out_reg[20]  ( .D(N23), .CK(clk), .Q(mac_out[20]) );
  DFF_X1 \mac_out_reg[21]  ( .D(N24), .CK(clk), .Q(mac_out[21]) );
  DFF_X1 \mac_out_reg[22]  ( .D(N25), .CK(clk), .Q(mac_out[22]) );
  DFF_X1 \mac_out_reg[23]  ( .D(N26), .CK(clk), .Q(mac_out[23]) );
  DFF_X1 \mac_out_reg[24]  ( .D(N27), .CK(clk), .Q(mac_out[24]) );
  DFF_X1 \mac_out_reg[25]  ( .D(N28), .CK(clk), .Q(mac_out[25]) );
  DFF_X1 \mac_out_reg[26]  ( .D(N29), .CK(clk), .Q(mac_out[26]) );
  DFF_X1 \mac_out_reg[27]  ( .D(N30), .CK(clk), .Q(mac_out[27]) );
  DFF_X1 \mac_out_reg[28]  ( .D(N31), .CK(clk), .Q(mac_out[28]) );
  DFF_X1 \mac_out_reg[29]  ( .D(N32), .CK(clk), .Q(mac_out[29]) );
  DFF_X1 \mac_out_reg[30]  ( .D(N33), .CK(clk), .Q(mac_out[30]) );
  DFF_X1 \mac_out_reg[31]  ( .D(N34), .CK(clk), .Q(mac_out[31]) );
  DFF_X1 \mac_out_reg[32]  ( .D(N35), .CK(clk), .Q(mac_out[32]) );
  DFF_X1 \mac_out_reg[33]  ( .D(N36), .CK(clk), .Q(mac_out[33]) );
  DFF_X1 \mac_out_reg[34]  ( .D(N37), .CK(clk), .Q(mac_out[34]) );
  DFF_X1 \mac_out_reg[35]  ( .D(N38), .CK(clk), .Q(mac_out[35]) );
  DFF_X1 \mac_out_reg[36]  ( .D(N39), .CK(clk), .Q(mac_out[36]) );
  DFF_X1 \mac_out_reg[37]  ( .D(N40), .CK(clk), .Q(mac_out[37]) );
  DFF_X1 \mac_out_reg[38]  ( .D(N41), .CK(clk), .Q(mac_out[38]) );
  DFF_X1 \mac_out_reg[39]  ( .D(N42), .CK(clk), .Q(mac_out[39]) );
  mac_4_DW_mult_tc_1 mult_355 ( .a(a), .b(b), .product(mul) );
  mac_4_DW01_add_1 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  DFF_X2 \pipeline_reg[39]  ( .D(mul[39]), .CK(clk), .Q(pipeline[39]) );
  BUF_X1 U3 ( .A(n3), .Z(n2) );
  INV_X1 U4 ( .A(clear_acc), .ZN(n3) );
  AND2_X1 U6 ( .A1(sum[39]), .A2(n2), .ZN(N42) );
  AND2_X1 U7 ( .A1(sum[38]), .A2(n2), .ZN(N41) );
  AND2_X1 U8 ( .A1(sum[37]), .A2(n2), .ZN(N40) );
  AND2_X1 U9 ( .A1(sum[36]), .A2(n2), .ZN(N39) );
  AND2_X1 U10 ( .A1(sum[35]), .A2(n2), .ZN(N38) );
  AND2_X1 U11 ( .A1(sum[34]), .A2(n2), .ZN(N37) );
  AND2_X1 U12 ( .A1(sum[33]), .A2(n2), .ZN(N36) );
  AND2_X1 U13 ( .A1(sum[32]), .A2(n2), .ZN(N35) );
  AND2_X1 U14 ( .A1(sum[31]), .A2(n2), .ZN(N34) );
  AND2_X1 U15 ( .A1(sum[30]), .A2(n2), .ZN(N33) );
  AND2_X1 U16 ( .A1(sum[29]), .A2(n2), .ZN(N32) );
  AND2_X1 U17 ( .A1(sum[28]), .A2(n3), .ZN(N31) );
  AND2_X1 U18 ( .A1(sum[27]), .A2(n3), .ZN(N30) );
  AND2_X1 U19 ( .A1(sum[26]), .A2(n3), .ZN(N29) );
  AND2_X1 U20 ( .A1(sum[25]), .A2(n3), .ZN(N28) );
  AND2_X1 U21 ( .A1(sum[24]), .A2(n3), .ZN(N27) );
  AND2_X1 U22 ( .A1(sum[23]), .A2(n3), .ZN(N26) );
  AND2_X1 U23 ( .A1(sum[22]), .A2(n3), .ZN(N25) );
  AND2_X1 U24 ( .A1(sum[21]), .A2(n3), .ZN(N24) );
  AND2_X1 U25 ( .A1(sum[20]), .A2(n3), .ZN(N23) );
  AND2_X1 U26 ( .A1(sum[19]), .A2(n3), .ZN(N22) );
  AND2_X1 U27 ( .A1(sum[18]), .A2(n3), .ZN(N21) );
  AND2_X1 U28 ( .A1(sum[17]), .A2(n3), .ZN(N20) );
  AND2_X1 U29 ( .A1(sum[16]), .A2(n3), .ZN(N19) );
  AND2_X1 U30 ( .A1(sum[15]), .A2(n3), .ZN(N18) );
  AND2_X1 U31 ( .A1(sum[14]), .A2(n3), .ZN(N17) );
  AND2_X1 U32 ( .A1(sum[13]), .A2(n3), .ZN(N16) );
  AND2_X1 U33 ( .A1(sum[12]), .A2(n3), .ZN(N15) );
  AND2_X1 U34 ( .A1(sum[11]), .A2(n3), .ZN(N14) );
  AND2_X1 U35 ( .A1(sum[10]), .A2(n3), .ZN(N13) );
  AND2_X1 U36 ( .A1(sum[9]), .A2(n3), .ZN(N12) );
  AND2_X1 U37 ( .A1(sum[8]), .A2(n3), .ZN(N11) );
  AND2_X1 U38 ( .A1(sum[7]), .A2(n3), .ZN(N10) );
  AND2_X1 U39 ( .A1(sum[6]), .A2(n3), .ZN(N9) );
  AND2_X1 U40 ( .A1(sum[5]), .A2(n3), .ZN(N8) );
  AND2_X1 U41 ( .A1(sum[4]), .A2(n3), .ZN(N7) );
  AND2_X1 U42 ( .A1(sum[3]), .A2(n3), .ZN(N6) );
  AND2_X1 U43 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U44 ( .A1(sum[1]), .A2(n3), .ZN(N4) );
  AND2_X1 U45 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
endmodule


module mac_3_DW_mult_tc_1 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n4, n6, n7, n9, n12, n13, n16, n18, n19, n22, n24, n25, n28, n31,
         n34, n36, n37, n42, n43, n48, n49, n52, n54, n55, n60, n61, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n98, n99, n100, n101, n103, n105, n106, n107, n108, n109,
         n111, n113, n114, n115, n116, n117, n119, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n185, n186, n188, n193, n194, n195, n196, n200, n201, n202, n203,
         n204, n205, n206, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n225, n227, n228,
         n230, n232, n233, n234, n236, n238, n239, n240, n241, n242, n244,
         n246, n247, n248, n249, n250, n252, n254, n255, n256, n257, n258,
         n259, n260, n261, n263, n264, n266, n268, n270, n271, n273, n274,
         n275, n276, n277, n278, n279, n280, n284, n285, n286, n287, n291,
         n293, n295, n296, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n643, n644, n646, n649, n652, n653,
         n655, n656, n658, n659, n661, n662, n664, n665, n667, n668, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1115, n1119,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1233, n1234, n1235, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n37 = a[13];
  assign n43 = a[15];
  assign n49 = a[17];
  assign n55 = a[19];
  assign n61 = b[0];
  assign n668 = a[0];
  assign n1090 = b[19];
  assign n1091 = b[18];
  assign n1092 = b[17];
  assign n1093 = b[16];
  assign n1094 = b[15];
  assign n1095 = b[14];
  assign n1096 = b[13];
  assign n1097 = b[12];
  assign n1098 = b[11];
  assign n1099 = b[10];
  assign n1100 = b[9];
  assign n1101 = b[8];
  assign n1102 = b[7];
  assign n1103 = b[6];
  assign n1104 = b[5];
  assign n1105 = b[4];
  assign n1106 = b[3];
  assign n1107 = b[2];
  assign n1108 = b[1];

  FA_X1 U333 ( .A(n681), .B(n304), .CI(n700), .CO(n300), .S(n301) );
  FA_X1 U334 ( .A(n305), .B(n682), .CI(n308), .CO(n302), .S(n303) );
  FA_X1 U336 ( .A(n312), .B(n683), .CI(n309), .CO(n306), .S(n307) );
  FA_X1 U337 ( .A(n701), .B(n314), .CI(n720), .CO(n308), .S(n309) );
  FA_X1 U338 ( .A(n313), .B(n320), .CI(n318), .CO(n310), .S(n311) );
  FA_X1 U339 ( .A(n684), .B(n702), .CI(n315), .CO(n312), .S(n313) );
  FA_X1 U341 ( .A(n324), .B(n321), .CI(n319), .CO(n316), .S(n317) );
  FA_X1 U342 ( .A(n328), .B(n721), .CI(n326), .CO(n318), .S(n319) );
  FA_X1 U343 ( .A(n703), .B(n685), .CI(n740), .CO(n320), .S(n321) );
  FA_X1 U344 ( .A(n325), .B(n327), .CI(n332), .CO(n322), .S(n323) );
  FA_X1 U345 ( .A(n336), .B(n329), .CI(n334), .CO(n324), .S(n325) );
  FA_X1 U346 ( .A(n686), .B(n704), .CI(n722), .CO(n326), .S(n327) );
  FA_X1 U348 ( .A(n340), .B(n342), .CI(n333), .CO(n330), .S(n331) );
  FA_X1 U349 ( .A(n335), .B(n344), .CI(n337), .CO(n332), .S(n333) );
  FA_X1 U350 ( .A(n705), .B(n346), .CI(n723), .CO(n334), .S(n335) );
  FA_X1 U351 ( .A(n741), .B(n687), .CI(n760), .CO(n336), .S(n337) );
  FA_X1 U352 ( .A(n350), .B(n343), .CI(n341), .CO(n338), .S(n339) );
  FA_X1 U353 ( .A(n345), .B(n354), .CI(n352), .CO(n340), .S(n341) );
  FA_X1 U354 ( .A(n347), .B(n724), .CI(n356), .CO(n342), .S(n343) );
  FA_X1 U355 ( .A(n742), .B(n706), .CI(n688), .CO(n344), .S(n345) );
  FA_X1 U357 ( .A(n360), .B(n353), .CI(n351), .CO(n348), .S(n349) );
  FA_X1 U358 ( .A(n357), .B(n355), .CI(n362), .CO(n350), .S(n351) );
  FA_X1 U359 ( .A(n366), .B(n743), .CI(n364), .CO(n352), .S(n353) );
  FA_X1 U360 ( .A(n707), .B(n761), .CI(n725), .CO(n354), .S(n355) );
  FA_X1 U361 ( .A(n368), .B(n689), .CI(n780), .CO(n356), .S(n357) );
  FA_X1 U362 ( .A(n372), .B(n363), .CI(n361), .CO(n358), .S(n359) );
  FA_X1 U363 ( .A(n376), .B(n365), .CI(n374), .CO(n360), .S(n361) );
  FA_X1 U364 ( .A(n378), .B(n380), .CI(n367), .CO(n362), .S(n363) );
  FA_X1 U365 ( .A(n690), .B(n708), .CI(n369), .CO(n364), .S(n365) );
  FA_X1 U366 ( .A(n762), .B(n726), .CI(n744), .CO(n366), .S(n367) );
  FA_X1 U368 ( .A(n384), .B(n375), .CI(n373), .CO(n370), .S(n371) );
  FA_X1 U369 ( .A(n377), .B(n388), .CI(n386), .CO(n372), .S(n373) );
  FA_X1 U370 ( .A(n379), .B(n390), .CI(n381), .CO(n374), .S(n375) );
  FA_X1 U371 ( .A(n727), .B(n745), .CI(n392), .CO(n376), .S(n377) );
  FA_X1 U372 ( .A(n709), .B(n781), .CI(n763), .CO(n378), .S(n379) );
  FA_X1 U373 ( .A(n394), .B(n691), .CI(n800), .CO(n380), .S(n381) );
  FA_X1 U374 ( .A(n398), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U375 ( .A(n389), .B(n402), .CI(n400), .CO(n384), .S(n385) );
  FA_X1 U376 ( .A(n391), .B(n404), .CI(n393), .CO(n386), .S(n387) );
  FA_X1 U377 ( .A(n408), .B(n395), .CI(n406), .CO(n388), .S(n389) );
  FA_X1 U378 ( .A(n746), .B(n782), .CI(n764), .CO(n390), .S(n391) );
  FA_X1 U379 ( .A(n692), .B(n728), .CI(n710), .CO(n392), .S(n393) );
  FA_X1 U381 ( .A(n412), .B(n401), .CI(n399), .CO(n396), .S(n397) );
  FA_X1 U382 ( .A(n403), .B(n416), .CI(n414), .CO(n398), .S(n399) );
  FA_X1 U383 ( .A(n409), .B(n407), .CI(n418), .CO(n400), .S(n401) );
  FA_X1 U384 ( .A(n420), .B(n422), .CI(n405), .CO(n402), .S(n403) );
  FA_X1 U385 ( .A(n765), .B(n747), .CI(n729), .CO(n404), .S(n405) );
  FA_X1 U386 ( .A(n711), .B(n801), .CI(n783), .CO(n406), .S(n407) );
  FA_X1 U387 ( .A(n1274), .B(n693), .CI(n820), .CO(n408), .S(n409) );
  FA_X1 U388 ( .A(n428), .B(n415), .CI(n413), .CO(n410), .S(n411) );
  FA_X1 U391 ( .A(n438), .B(n436), .CI(n421), .CO(n416), .S(n417) );
  FA_X1 U393 ( .A(n694), .B(n766), .CI(n712), .CO(n420), .S(n421) );
  FA_X1 U394 ( .A(n802), .B(n730), .CI(n784), .CO(n422), .S(n423) );
  FA_X1 U399 ( .A(n437), .B(n452), .CI(n439), .CO(n432), .S(n433) );
  FA_X1 U400 ( .A(n456), .B(n767), .CI(n454), .CO(n434), .S(n435) );
  FA_X1 U401 ( .A(n731), .B(n785), .CI(n749), .CO(n436), .S(n437) );
  FA_X1 U402 ( .A(n713), .B(n803), .CI(n458), .CO(n438), .S(n439) );
  FA_X1 U403 ( .A(n821), .B(n695), .CI(n840), .CO(n440), .S(n441) );
  FA_X1 U406 ( .A(n468), .B(n453), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U407 ( .A(n455), .B(n470), .CI(n457), .CO(n448), .S(n449) );
  FA_X1 U408 ( .A(n476), .B(n474), .CI(n472), .CO(n450), .S(n451) );
  FA_X1 U409 ( .A(n768), .B(n786), .CI(n459), .CO(n452), .S(n453) );
  FA_X1 U410 ( .A(n732), .B(n714), .CI(n804), .CO(n454), .S(n455) );
  FA_X1 U411 ( .A(n822), .B(n696), .CI(n750), .CO(n456), .S(n457) );
  FA_X1 U413 ( .A(n480), .B(n465), .CI(n463), .CO(n460), .S(n461) );
  FA_X1 U414 ( .A(n467), .B(n484), .CI(n482), .CO(n462), .S(n463) );
  FA_X1 U416 ( .A(n473), .B(n488), .CI(n475), .CO(n466), .S(n467) );
  FA_X1 U417 ( .A(n492), .B(n477), .CI(n490), .CO(n468), .S(n469) );
  FA_X1 U418 ( .A(n805), .B(n823), .CI(n494), .CO(n470), .S(n471) );
  FA_X1 U419 ( .A(n751), .B(n733), .CI(n841), .CO(n472), .S(n473) );
  FA_X1 U420 ( .A(n860), .B(n697), .CI(n769), .CO(n474), .S(n475) );
  FA_X1 U426 ( .A(n489), .B(n506), .CI(n491), .CO(n484), .S(n485) );
  FA_X1 U427 ( .A(n510), .B(n495), .CI(n508), .CO(n486), .S(n487) );
  FA_X1 U428 ( .A(n770), .B(n842), .CI(n824), .CO(n488), .S(n489) );
  FA_X1 U429 ( .A(n861), .B(n806), .CI(n752), .CO(n490), .S(n491) );
  FA_X1 U430 ( .A(n788), .B(n670), .CI(n734), .CO(n492), .S(n493) );
  HA_X1 U431 ( .A(n698), .B(n716), .CO(n494), .S(n495) );
  FA_X1 U433 ( .A(n516), .B(n505), .CI(n503), .CO(n498), .S(n499) );
  FA_X1 U434 ( .A(n520), .B(n509), .CI(n518), .CO(n500), .S(n501) );
  FA_X1 U436 ( .A(n526), .B(n807), .CI(n524), .CO(n504), .S(n505) );
  FA_X1 U437 ( .A(n789), .B(n825), .CI(n771), .CO(n506), .S(n507) );
  FA_X1 U438 ( .A(n717), .B(n843), .CI(n753), .CO(n508), .S(n509) );
  FA_X1 U439 ( .A(n699), .B(n735), .CI(n862), .CO(n510), .S(n511) );
  FA_X1 U441 ( .A(n519), .B(n521), .CI(n532), .CO(n514), .S(n515) );
  FA_X1 U442 ( .A(n525), .B(n523), .CI(n534), .CO(n516), .S(n517) );
  FA_X1 U444 ( .A(n826), .B(n844), .CI(n527), .CO(n520), .S(n521) );
  FA_X1 U445 ( .A(n808), .B(n772), .CI(n754), .CO(n522), .S(n523) );
  FA_X1 U446 ( .A(n863), .B(n790), .CI(n671), .CO(n524), .S(n525) );
  HA_X1 U447 ( .A(n718), .B(n736), .CO(n526), .S(n527) );
  FA_X1 U448 ( .A(n533), .B(n544), .CI(n531), .CO(n528), .S(n529) );
  FA_X1 U449 ( .A(n546), .B(n548), .CI(n535), .CO(n530), .S(n531) );
  FA_X1 U450 ( .A(n537), .B(n541), .CI(n539), .CO(n532), .S(n533) );
  FA_X1 U452 ( .A(n791), .B(n827), .CI(n809), .CO(n536), .S(n537) );
  FA_X1 U453 ( .A(n737), .B(n845), .CI(n773), .CO(n538), .S(n539) );
  FA_X1 U458 ( .A(n555), .B(n846), .CI(n566), .CO(n548), .S(n549) );
  FA_X1 U459 ( .A(n865), .B(n792), .CI(n828), .CO(n550), .S(n551) );
  HA_X1 U461 ( .A(n738), .B(n756), .CO(n554), .S(n555) );
  FA_X1 U464 ( .A(n574), .B(n576), .CI(n567), .CO(n560), .S(n561) );
  FA_X1 U466 ( .A(n757), .B(n847), .CI(n793), .CO(n564), .S(n565) );
  FA_X1 U467 ( .A(n866), .B(n739), .CI(n775), .CO(n566), .S(n567) );
  FA_X1 U468 ( .A(n582), .B(n573), .CI(n571), .CO(n568), .S(n569) );
  FA_X1 U469 ( .A(n577), .B(n575), .CI(n584), .CO(n570), .S(n571) );
  FA_X1 U470 ( .A(n588), .B(n579), .CI(n586), .CO(n572), .S(n573) );
  FA_X1 U471 ( .A(n794), .B(n848), .CI(n830), .CO(n574), .S(n575) );
  FA_X1 U472 ( .A(n867), .B(n812), .CI(n673), .CO(n576), .S(n577) );
  HA_X1 U473 ( .A(n758), .B(n776), .CO(n578), .S(n579) );
  FA_X1 U474 ( .A(n585), .B(n592), .CI(n583), .CO(n580), .S(n581) );
  FA_X1 U475 ( .A(n587), .B(n589), .CI(n594), .CO(n582), .S(n583) );
  FA_X1 U476 ( .A(n598), .B(n831), .CI(n596), .CO(n584), .S(n585) );
  FA_X1 U477 ( .A(n777), .B(n849), .CI(n813), .CO(n586), .S(n587) );
  FA_X1 U478 ( .A(n795), .B(n759), .CI(n868), .CO(n588), .S(n589) );
  FA_X1 U479 ( .A(n602), .B(n595), .CI(n593), .CO(n590), .S(n591) );
  FA_X1 U480 ( .A(n604), .B(n606), .CI(n597), .CO(n592), .S(n593) );
  FA_X1 U481 ( .A(n814), .B(n850), .CI(n599), .CO(n594), .S(n595) );
  FA_X1 U482 ( .A(n832), .B(n674), .CI(n869), .CO(n596), .S(n597) );
  HA_X1 U483 ( .A(n778), .B(n796), .CO(n598), .S(n599) );
  FA_X1 U484 ( .A(n610), .B(n605), .CI(n603), .CO(n600), .S(n601) );
  FA_X1 U485 ( .A(n612), .B(n614), .CI(n607), .CO(n602), .S(n603) );
  FA_X1 U486 ( .A(n797), .B(n851), .CI(n833), .CO(n604), .S(n605) );
  FA_X1 U488 ( .A(n613), .B(n618), .CI(n611), .CO(n608), .S(n609) );
  FA_X1 U489 ( .A(n615), .B(n871), .CI(n620), .CO(n610), .S(n611) );
  FA_X1 U490 ( .A(n852), .B(n834), .CI(n675), .CO(n612), .S(n613) );
  HA_X1 U491 ( .A(n798), .B(n816), .CO(n614), .S(n615) );
  FA_X1 U492 ( .A(n621), .B(n624), .CI(n619), .CO(n616), .S(n617) );
  FA_X1 U493 ( .A(n817), .B(n853), .CI(n626), .CO(n618), .S(n619) );
  FA_X1 U494 ( .A(n835), .B(n799), .CI(n872), .CO(n620), .S(n621) );
  FA_X1 U495 ( .A(n630), .B(n627), .CI(n625), .CO(n622), .S(n623) );
  FA_X1 U496 ( .A(n854), .B(n873), .CI(n676), .CO(n624), .S(n625) );
  HA_X1 U497 ( .A(n818), .B(n836), .CO(n626), .S(n627) );
  FA_X1 U498 ( .A(n634), .B(n837), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U499 ( .A(n874), .B(n819), .CI(n855), .CO(n630), .S(n631) );
  FA_X1 U500 ( .A(n677), .B(n856), .CI(n635), .CO(n632), .S(n633) );
  HA_X1 U501 ( .A(n838), .B(n875), .CO(n634), .S(n635) );
  FA_X1 U502 ( .A(n876), .B(n839), .CI(n857), .CO(n636), .S(n637) );
  HA_X1 U503 ( .A(n858), .B(n877), .CO(n638), .S(n639) );
  CLKBUF_X3 U1025 ( .A(n37), .Z(n1365) );
  BUF_X2 U1026 ( .A(n1094), .Z(n1560) );
  BUF_X2 U1027 ( .A(n1312), .Z(n1241) );
  CLKBUF_X2 U1028 ( .A(n42), .Z(n1504) );
  BUF_X1 U1029 ( .A(n1100), .Z(n1337) );
  BUF_X1 U1030 ( .A(n1108), .Z(n1346) );
  CLKBUF_X3 U1031 ( .A(n1099), .Z(n1555) );
  BUF_X2 U1032 ( .A(n7), .Z(n1537) );
  BUF_X1 U1033 ( .A(n1097), .Z(n1557) );
  BUF_X1 U1034 ( .A(n28), .Z(n1514) );
  BUF_X1 U1035 ( .A(n28), .Z(n1312) );
  BUF_X2 U1036 ( .A(n1098), .Z(n1350) );
  BUF_X2 U1037 ( .A(n1103), .Z(n1551) );
  BUF_X2 U1038 ( .A(n49), .Z(n1544) );
  BUF_X2 U1039 ( .A(n1), .Z(n1447) );
  BUF_X1 U1040 ( .A(n6), .Z(n1272) );
  OR2_X1 U1041 ( .A1(n529), .A2(n542), .ZN(n1233) );
  OR2_X1 U1042 ( .A1(n371), .A2(n382), .ZN(n1234) );
  OR2_X1 U1043 ( .A1(n679), .A2(n879), .ZN(n1235) );
  AND2_X1 U1044 ( .A1(n1235), .A2(n263), .ZN(product[1]) );
  BUF_X4 U1045 ( .A(n19), .Z(n1539) );
  XNOR2_X1 U1046 ( .A(n1559), .B(n1316), .ZN(n1237) );
  NAND3_X1 U1047 ( .A1(n1386), .A2(n1387), .A3(n1388), .ZN(n1238) );
  NAND3_X1 U1048 ( .A1(n1386), .A2(n1387), .A3(n1388), .ZN(n1239) );
  XNOR2_X1 U1049 ( .A(n1559), .B(n1335), .ZN(n1240) );
  BUF_X2 U1050 ( .A(n1095), .Z(n1559) );
  CLKBUF_X3 U1051 ( .A(n1448), .Z(n1316) );
  XNOR2_X1 U1052 ( .A(n499), .B(n1242), .ZN(n497) );
  XNOR2_X1 U1053 ( .A(n514), .B(n501), .ZN(n1242) );
  BUF_X2 U1054 ( .A(n13), .Z(n1335) );
  XNOR2_X1 U1055 ( .A(n1243), .B(n1245), .ZN(n429) );
  XNOR2_X1 U1056 ( .A(n433), .B(n448), .ZN(n1243) );
  XNOR2_X1 U1057 ( .A(n1), .B(a[2]), .ZN(n1244) );
  INV_X1 U1058 ( .A(n1308), .ZN(n1533) );
  CLKBUF_X2 U1059 ( .A(n1308), .Z(n1507) );
  CLKBUF_X1 U1060 ( .A(n446), .Z(n1245) );
  BUF_X2 U1061 ( .A(n1101), .Z(n1553) );
  XNOR2_X1 U1062 ( .A(n1555), .B(n1543), .ZN(n1246) );
  CLKBUF_X1 U1063 ( .A(n1269), .Z(n1247) );
  BUF_X1 U1064 ( .A(n25), .Z(n1540) );
  CLKBUF_X3 U1065 ( .A(n25), .Z(n1334) );
  CLKBUF_X1 U1066 ( .A(n417), .Z(n1248) );
  CLKBUF_X2 U1067 ( .A(n34), .Z(n1513) );
  BUF_X1 U1068 ( .A(n9), .Z(n1324) );
  BUF_X2 U1069 ( .A(n6), .Z(n1508) );
  XOR2_X1 U1070 ( .A(n500), .B(n487), .Z(n1249) );
  XOR2_X1 U1071 ( .A(n1249), .B(n485), .Z(n481) );
  XOR2_X1 U1072 ( .A(n498), .B(n483), .Z(n1250) );
  XOR2_X1 U1073 ( .A(n1250), .B(n481), .Z(n479) );
  NAND2_X1 U1074 ( .A1(n500), .A2(n487), .ZN(n1251) );
  NAND2_X1 U1075 ( .A1(n500), .A2(n485), .ZN(n1252) );
  NAND2_X1 U1076 ( .A1(n487), .A2(n485), .ZN(n1253) );
  NAND3_X1 U1077 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n480) );
  NAND2_X1 U1078 ( .A1(n498), .A2(n483), .ZN(n1254) );
  NAND2_X1 U1079 ( .A1(n498), .A2(n481), .ZN(n1255) );
  NAND2_X1 U1080 ( .A1(n483), .A2(n481), .ZN(n1256) );
  NAND3_X1 U1081 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n478) );
  XNOR2_X1 U1082 ( .A(n1555), .B(n1317), .ZN(n1257) );
  BUF_X2 U1083 ( .A(n1100), .Z(n1554) );
  CLKBUF_X1 U1084 ( .A(n434), .Z(n1258) );
  INV_X1 U1085 ( .A(n1233), .ZN(n1259) );
  BUF_X2 U1086 ( .A(n18), .Z(n1260) );
  CLKBUF_X2 U1087 ( .A(n1312), .Z(n1515) );
  CLKBUF_X1 U1088 ( .A(n175), .Z(n1261) );
  XNOR2_X1 U1089 ( .A(n1564), .B(n1447), .ZN(n1262) );
  BUF_X2 U1090 ( .A(n1107), .Z(n1548) );
  XOR2_X1 U1091 ( .A(n486), .B(n471), .Z(n1263) );
  XOR2_X1 U1092 ( .A(n469), .B(n1263), .Z(n465) );
  NAND2_X1 U1093 ( .A1(n469), .A2(n486), .ZN(n1264) );
  NAND2_X1 U1094 ( .A1(n469), .A2(n471), .ZN(n1265) );
  NAND2_X1 U1095 ( .A1(n486), .A2(n471), .ZN(n1266) );
  NAND3_X1 U1096 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n464) );
  NOR2_X1 U1097 ( .A1(n371), .A2(n382), .ZN(n1267) );
  NOR2_X1 U1098 ( .A1(n371), .A2(n382), .ZN(n135) );
  CLKBUF_X1 U1099 ( .A(n1524), .Z(n1268) );
  AND2_X1 U1100 ( .A1(n529), .A2(n542), .ZN(n1524) );
  NAND2_X1 U1101 ( .A1(n1115), .A2(n1514), .ZN(n1269) );
  CLKBUF_X1 U1102 ( .A(n221), .Z(n1270) );
  BUF_X1 U1103 ( .A(n6), .Z(n1509) );
  CLKBUF_X1 U1104 ( .A(n1503), .Z(n1271) );
  CLKBUF_X3 U1105 ( .A(n13), .Z(n1538) );
  INV_X1 U1106 ( .A(n275), .ZN(n1273) );
  OAI22_X1 U1107 ( .A1(n1475), .A2(n1028), .B1(n1027), .B2(n1516), .ZN(n1274)
         );
  BUF_X2 U1108 ( .A(n18), .Z(n1475) );
  XNOR2_X1 U1109 ( .A(n1275), .B(n464), .ZN(n445) );
  XNOR2_X1 U1110 ( .A(n449), .B(n466), .ZN(n1275) );
  BUF_X2 U1111 ( .A(n12), .Z(n1309) );
  NOR2_X1 U1112 ( .A1(n443), .A2(n460), .ZN(n161) );
  NAND2_X2 U1113 ( .A1(n1336), .A2(n1324), .ZN(n1477) );
  CLKBUF_X1 U1114 ( .A(n1104), .Z(n1550) );
  CLKBUF_X1 U1115 ( .A(n1104), .Z(n1343) );
  INV_X1 U1116 ( .A(n193), .ZN(n1276) );
  NAND2_X1 U1117 ( .A1(n511), .A2(n522), .ZN(n1295) );
  CLKBUF_X1 U1118 ( .A(n1104), .Z(n1344) );
  CLKBUF_X1 U1119 ( .A(n176), .Z(n1277) );
  BUF_X2 U1120 ( .A(n1102), .Z(n1552) );
  AOI21_X1 U1121 ( .B1(n1270), .B2(n213), .A(n214), .ZN(n1278) );
  NOR2_X2 U1122 ( .A1(n581), .A2(n590), .ZN(n215) );
  CLKBUF_X3 U1123 ( .A(n61), .Z(n1546) );
  CLKBUF_X1 U1124 ( .A(n870), .Z(n1339) );
  INV_X1 U1125 ( .A(n170), .ZN(n1279) );
  XOR2_X1 U1126 ( .A(n719), .B(n864), .Z(n1280) );
  XOR2_X1 U1127 ( .A(n755), .B(n1280), .Z(n541) );
  NAND2_X1 U1128 ( .A1(n755), .A2(n719), .ZN(n1281) );
  NAND2_X1 U1129 ( .A1(n755), .A2(n864), .ZN(n1282) );
  NAND2_X1 U1130 ( .A1(n719), .A2(n864), .ZN(n1283) );
  NAND3_X1 U1131 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n540) );
  NAND3_X1 U1132 ( .A1(n1408), .A2(n1409), .A3(n1410), .ZN(n1284) );
  CLKBUF_X1 U1133 ( .A(n1493), .Z(n1285) );
  XOR2_X1 U1134 ( .A(n425), .B(n748), .Z(n1286) );
  XOR2_X1 U1135 ( .A(n1286), .B(n440), .Z(n419) );
  XOR2_X1 U1136 ( .A(n423), .B(n1258), .Z(n1287) );
  XOR2_X1 U1137 ( .A(n1287), .B(n419), .Z(n415) );
  NAND2_X1 U1138 ( .A1(n425), .A2(n748), .ZN(n1288) );
  NAND2_X1 U1139 ( .A1(n440), .A2(n425), .ZN(n1289) );
  NAND2_X1 U1140 ( .A1(n440), .A2(n748), .ZN(n1290) );
  NAND3_X1 U1141 ( .A1(n1288), .A2(n1289), .A3(n1290), .ZN(n418) );
  NAND2_X1 U1142 ( .A1(n423), .A2(n434), .ZN(n1291) );
  NAND2_X1 U1143 ( .A1(n423), .A2(n419), .ZN(n1292) );
  NAND2_X1 U1144 ( .A1(n434), .A2(n419), .ZN(n1293) );
  NAND3_X1 U1145 ( .A1(n1291), .A2(n1292), .A3(n1293), .ZN(n414) );
  XOR2_X1 U1146 ( .A(n511), .B(n522), .Z(n1294) );
  XOR2_X1 U1147 ( .A(n1294), .B(n507), .Z(n503) );
  NAND2_X1 U1148 ( .A1(n511), .A2(n507), .ZN(n1296) );
  NAND2_X1 U1149 ( .A1(n522), .A2(n507), .ZN(n1297) );
  NAND3_X1 U1150 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n502) );
  XOR2_X1 U1151 ( .A(n504), .B(n493), .Z(n1298) );
  XOR2_X1 U1152 ( .A(n1298), .B(n502), .Z(n483) );
  NAND2_X1 U1153 ( .A1(n504), .A2(n493), .ZN(n1299) );
  NAND2_X1 U1154 ( .A1(n504), .A2(n502), .ZN(n1300) );
  NAND2_X1 U1155 ( .A1(n493), .A2(n502), .ZN(n1301) );
  NAND3_X1 U1156 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n482) );
  CLKBUF_X3 U1157 ( .A(n36), .Z(n1480) );
  INV_X1 U1158 ( .A(n662), .ZN(n1302) );
  CLKBUF_X1 U1159 ( .A(n1369), .Z(n1303) );
  INV_X1 U1160 ( .A(n1142), .ZN(n1304) );
  XNOR2_X1 U1161 ( .A(n7), .B(a[4]), .ZN(n1305) );
  XNOR2_X1 U1162 ( .A(n1306), .B(n559), .ZN(n557) );
  XNOR2_X1 U1163 ( .A(n561), .B(n570), .ZN(n1306) );
  CLKBUF_X1 U1164 ( .A(n1564), .Z(n1307) );
  XNOR2_X1 U1165 ( .A(n31), .B(a[12]), .ZN(n1308) );
  NAND2_X1 U1166 ( .A1(n1489), .A2(n1244), .ZN(n12) );
  NOR2_X1 U1167 ( .A1(n411), .A2(n426), .ZN(n150) );
  XNOR2_X1 U1168 ( .A(n578), .B(n1310), .ZN(n563) );
  XNOR2_X1 U1169 ( .A(n829), .B(n811), .ZN(n1310) );
  XNOR2_X1 U1170 ( .A(n1453), .B(n1311), .ZN(product[38]) );
  AND3_X1 U1171 ( .A1(n1451), .A2(n1450), .A3(n1452), .ZN(n1311) );
  CLKBUF_X1 U1172 ( .A(n148), .Z(n1313) );
  CLKBUF_X1 U1173 ( .A(n1557), .Z(n1314) );
  BUF_X1 U1174 ( .A(n1244), .Z(n1505) );
  BUF_X1 U1175 ( .A(n9), .Z(n1506) );
  CLKBUF_X1 U1176 ( .A(n1448), .Z(n1315) );
  BUF_X1 U1177 ( .A(n1448), .Z(n1317) );
  CLKBUF_X1 U1178 ( .A(n1561), .Z(n1318) );
  BUF_X2 U1179 ( .A(n1093), .Z(n1561) );
  BUF_X2 U1180 ( .A(n37), .Z(n1542) );
  CLKBUF_X1 U1181 ( .A(n264), .Z(n1319) );
  CLKBUF_X1 U1182 ( .A(n100), .Z(n1320) );
  CLKBUF_X1 U1183 ( .A(n98), .Z(n1321) );
  INV_X1 U1184 ( .A(n1558), .ZN(n1322) );
  INV_X1 U1185 ( .A(n1322), .ZN(n1323) );
  BUF_X2 U1186 ( .A(n1096), .Z(n1558) );
  XNOR2_X1 U1187 ( .A(n1), .B(n1357), .ZN(n1119) );
  BUF_X1 U1188 ( .A(n1106), .Z(n1325) );
  BUF_X1 U1189 ( .A(n1106), .Z(n1326) );
  CLKBUF_X1 U1190 ( .A(n126), .Z(n1327) );
  XNOR2_X1 U1191 ( .A(n1328), .B(n552), .ZN(n535) );
  XNOR2_X1 U1192 ( .A(n554), .B(n550), .ZN(n1328) );
  BUF_X2 U1193 ( .A(n55), .Z(n1329) );
  CLKBUF_X2 U1194 ( .A(n55), .Z(n1330) );
  CLKBUF_X1 U1195 ( .A(n55), .Z(n1545) );
  CLKBUF_X1 U1196 ( .A(n1370), .Z(n1331) );
  XNOR2_X1 U1197 ( .A(n1564), .B(n1537), .ZN(n1332) );
  CLKBUF_X1 U1198 ( .A(n7), .Z(n1333) );
  BUF_X1 U1199 ( .A(n6), .Z(n1510) );
  CLKBUF_X1 U1200 ( .A(n1489), .Z(n1336) );
  CLKBUF_X1 U1201 ( .A(n1486), .Z(n1338) );
  INV_X1 U1202 ( .A(n1362), .ZN(n1486) );
  XNOR2_X1 U1203 ( .A(n1340), .B(n429), .ZN(n427) );
  XNOR2_X1 U1204 ( .A(n444), .B(n431), .ZN(n1340) );
  AOI21_X1 U1205 ( .B1(n1520), .B2(n1268), .A(n1528), .ZN(n1341) );
  CLKBUF_X1 U1206 ( .A(n1553), .Z(n1342) );
  BUF_X1 U1207 ( .A(n1107), .Z(n1345) );
  CLKBUF_X1 U1208 ( .A(n1108), .Z(n1347) );
  INV_X2 U1209 ( .A(n1141), .ZN(n1348) );
  CLKBUF_X1 U1210 ( .A(n1507), .Z(n1349) );
  CLKBUF_X1 U1211 ( .A(n1098), .Z(n1556) );
  CLKBUF_X1 U1212 ( .A(n1563), .Z(n1351) );
  BUF_X2 U1213 ( .A(n1091), .Z(n1563) );
  BUF_X2 U1214 ( .A(n1549), .Z(n1352) );
  CLKBUF_X1 U1215 ( .A(n1549), .Z(n1353) );
  BUF_X2 U1216 ( .A(n1562), .Z(n1354) );
  BUF_X1 U1217 ( .A(n1562), .Z(n1355) );
  BUF_X1 U1218 ( .A(n1106), .Z(n1356) );
  INV_X1 U1219 ( .A(n668), .ZN(n1357) );
  BUF_X2 U1220 ( .A(n1090), .Z(n1564) );
  NAND3_X1 U1221 ( .A1(n1370), .A2(n1369), .A3(n1368), .ZN(n1358) );
  NAND3_X1 U1222 ( .A1(n1368), .A2(n1303), .A3(n1331), .ZN(n1359) );
  NAND3_X1 U1223 ( .A1(n1373), .A2(n1374), .A3(n1372), .ZN(n1360) );
  AOI21_X1 U1224 ( .B1(n1261), .B2(n1276), .A(n1277), .ZN(n1361) );
  XOR2_X1 U1225 ( .A(n49), .B(a[18]), .Z(n1362) );
  NOR2_X1 U1226 ( .A1(n427), .A2(n442), .ZN(n1493) );
  NAND3_X1 U1227 ( .A1(n1394), .A2(n1395), .A3(n1396), .ZN(n1363) );
  CLKBUF_X1 U1228 ( .A(n134), .Z(n1364) );
  XNOR2_X1 U1229 ( .A(n1366), .B(n445), .ZN(n443) );
  XNOR2_X1 U1230 ( .A(n462), .B(n447), .ZN(n1366) );
  XOR2_X1 U1231 ( .A(n303), .B(n306), .Z(n1367) );
  XOR2_X1 U1232 ( .A(n1367), .B(n1320), .Z(product[35]) );
  NAND2_X1 U1233 ( .A1(n303), .A2(n306), .ZN(n1368) );
  NAND2_X1 U1234 ( .A1(n303), .A2(n1363), .ZN(n1369) );
  NAND2_X1 U1235 ( .A1(n100), .A2(n306), .ZN(n1370) );
  NAND3_X1 U1236 ( .A1(n1370), .A2(n1369), .A3(n1368), .ZN(n99) );
  XOR2_X1 U1237 ( .A(n302), .B(n301), .Z(n1371) );
  XOR2_X1 U1238 ( .A(n1371), .B(n1359), .Z(product[36]) );
  NAND2_X1 U1239 ( .A1(n302), .A2(n301), .ZN(n1372) );
  NAND2_X1 U1240 ( .A1(n1358), .A2(n302), .ZN(n1373) );
  NAND2_X1 U1241 ( .A1(n99), .A2(n301), .ZN(n1374) );
  NAND3_X1 U1242 ( .A1(n1374), .A2(n1373), .A3(n1372), .ZN(n98) );
  INV_X1 U1243 ( .A(n1428), .ZN(n1375) );
  BUF_X2 U1244 ( .A(n42), .Z(n1503) );
  AND3_X1 U1245 ( .A1(n1456), .A2(n1455), .A3(n1454), .ZN(product[39]) );
  NAND3_X1 U1246 ( .A1(n1451), .A2(n1452), .A3(n1450), .ZN(n1377) );
  CLKBUF_X1 U1247 ( .A(n114), .Z(n1378) );
  NAND2_X1 U1248 ( .A1(n433), .A2(n448), .ZN(n1379) );
  NAND2_X1 U1249 ( .A1(n446), .A2(n433), .ZN(n1380) );
  NAND2_X1 U1250 ( .A1(n446), .A2(n448), .ZN(n1381) );
  NAND3_X1 U1251 ( .A1(n1379), .A2(n1380), .A3(n1381), .ZN(n428) );
  NAND2_X1 U1252 ( .A1(n1284), .A2(n431), .ZN(n1382) );
  NAND2_X1 U1253 ( .A1(n1284), .A2(n429), .ZN(n1383) );
  NAND2_X1 U1254 ( .A1(n431), .A2(n429), .ZN(n1384) );
  NAND3_X1 U1255 ( .A1(n1382), .A2(n1383), .A3(n1384), .ZN(n426) );
  OR2_X2 U1256 ( .A1(n1439), .A2(n1440), .ZN(n60) );
  XOR2_X1 U1257 ( .A(n450), .B(n441), .Z(n1385) );
  XOR2_X1 U1258 ( .A(n1385), .B(n435), .Z(n431) );
  NAND2_X1 U1259 ( .A1(n450), .A2(n441), .ZN(n1386) );
  NAND2_X1 U1260 ( .A1(n450), .A2(n435), .ZN(n1387) );
  NAND2_X1 U1261 ( .A1(n441), .A2(n435), .ZN(n1388) );
  NAND3_X1 U1262 ( .A1(n1386), .A2(n1387), .A3(n1388), .ZN(n430) );
  XOR2_X1 U1263 ( .A(n417), .B(n432), .Z(n1389) );
  XOR2_X1 U1264 ( .A(n1389), .B(n1239), .Z(n413) );
  NAND2_X1 U1265 ( .A1(n1248), .A2(n432), .ZN(n1390) );
  NAND2_X1 U1266 ( .A1(n417), .A2(n1238), .ZN(n1391) );
  NAND2_X1 U1267 ( .A1(n432), .A2(n430), .ZN(n1392) );
  NAND3_X1 U1268 ( .A1(n1390), .A2(n1391), .A3(n1392), .ZN(n412) );
  XOR2_X1 U1269 ( .A(n307), .B(n310), .Z(n1393) );
  XOR2_X1 U1270 ( .A(n1319), .B(n1393), .Z(product[34]) );
  NAND2_X1 U1271 ( .A1(n264), .A2(n307), .ZN(n1394) );
  NAND2_X1 U1272 ( .A1(n264), .A2(n310), .ZN(n1395) );
  NAND2_X1 U1273 ( .A1(n307), .A2(n310), .ZN(n1396) );
  NAND3_X1 U1274 ( .A1(n1395), .A2(n1394), .A3(n1396), .ZN(n100) );
  XOR2_X1 U1275 ( .A(n672), .B(n774), .Z(n1397) );
  XOR2_X1 U1276 ( .A(n1397), .B(n810), .Z(n553) );
  NAND2_X1 U1277 ( .A1(n774), .A2(n672), .ZN(n1398) );
  NAND2_X1 U1278 ( .A1(n774), .A2(n810), .ZN(n1399) );
  NAND2_X1 U1279 ( .A1(n672), .A2(n810), .ZN(n1400) );
  NAND3_X1 U1280 ( .A1(n1398), .A2(n1399), .A3(n1400), .ZN(n552) );
  NAND2_X1 U1281 ( .A1(n554), .A2(n550), .ZN(n1401) );
  NAND2_X1 U1282 ( .A1(n554), .A2(n552), .ZN(n1402) );
  NAND2_X1 U1283 ( .A1(n550), .A2(n552), .ZN(n1403) );
  NAND3_X1 U1284 ( .A1(n1401), .A2(n1402), .A3(n1403), .ZN(n534) );
  NAND2_X1 U1285 ( .A1(n499), .A2(n514), .ZN(n1404) );
  NAND2_X1 U1286 ( .A1(n499), .A2(n501), .ZN(n1405) );
  NAND2_X1 U1287 ( .A1(n514), .A2(n501), .ZN(n1406) );
  NAND3_X1 U1288 ( .A1(n1404), .A2(n1405), .A3(n1406), .ZN(n496) );
  XNOR2_X1 U1289 ( .A(n540), .B(n1407), .ZN(n519) );
  XNOR2_X1 U1290 ( .A(n536), .B(n538), .ZN(n1407) );
  NAND2_X1 U1291 ( .A1(n449), .A2(n466), .ZN(n1408) );
  NAND2_X1 U1292 ( .A1(n449), .A2(n464), .ZN(n1409) );
  NAND2_X1 U1293 ( .A1(n466), .A2(n464), .ZN(n1410) );
  NAND3_X1 U1294 ( .A1(n1410), .A2(n1409), .A3(n1408), .ZN(n444) );
  NAND2_X1 U1295 ( .A1(n462), .A2(n447), .ZN(n1411) );
  NAND2_X1 U1296 ( .A1(n462), .A2(n445), .ZN(n1412) );
  NAND2_X1 U1297 ( .A1(n447), .A2(n445), .ZN(n1413) );
  NAND3_X1 U1298 ( .A1(n1411), .A2(n1412), .A3(n1413), .ZN(n442) );
  OR2_X1 U1299 ( .A1(n54), .A2(n919), .ZN(n1414) );
  OR2_X1 U1300 ( .A1(n918), .A2(n1511), .ZN(n1415) );
  NAND2_X1 U1301 ( .A1(n1414), .A2(n1415), .ZN(n717) );
  CLKBUF_X3 U1302 ( .A(n52), .Z(n1511) );
  CLKBUF_X1 U1303 ( .A(n127), .Z(n1416) );
  NAND2_X1 U1304 ( .A1(n1115), .A2(n1514), .ZN(n1417) );
  NAND2_X1 U1305 ( .A1(n1115), .A2(n1514), .ZN(n1484) );
  CLKBUF_X1 U1306 ( .A(n165), .Z(n1418) );
  XOR2_X1 U1307 ( .A(n560), .B(n553), .Z(n1419) );
  XOR2_X1 U1308 ( .A(n1419), .B(n549), .Z(n545) );
  XOR2_X1 U1309 ( .A(n547), .B(n558), .Z(n1420) );
  XOR2_X1 U1310 ( .A(n1420), .B(n545), .Z(n543) );
  NAND2_X1 U1311 ( .A1(n1427), .A2(n553), .ZN(n1421) );
  NAND2_X1 U1312 ( .A1(n1427), .A2(n549), .ZN(n1422) );
  NAND2_X1 U1313 ( .A1(n553), .A2(n549), .ZN(n1423) );
  NAND3_X1 U1314 ( .A1(n1421), .A2(n1422), .A3(n1423), .ZN(n544) );
  NAND2_X1 U1315 ( .A1(n547), .A2(n558), .ZN(n1424) );
  NAND2_X1 U1316 ( .A1(n547), .A2(n545), .ZN(n1425) );
  NAND2_X1 U1317 ( .A1(n558), .A2(n545), .ZN(n1426) );
  NAND3_X1 U1318 ( .A1(n1424), .A2(n1425), .A3(n1426), .ZN(n542) );
  CLKBUF_X1 U1319 ( .A(n560), .Z(n1427) );
  XOR2_X1 U1320 ( .A(n1542), .B(a[14]), .Z(n1428) );
  XOR2_X1 U1321 ( .A(n563), .B(n565), .Z(n1429) );
  XOR2_X1 U1322 ( .A(n1429), .B(n572), .Z(n559) );
  NAND2_X1 U1323 ( .A1(n563), .A2(n565), .ZN(n1430) );
  NAND2_X1 U1324 ( .A1(n563), .A2(n572), .ZN(n1431) );
  NAND2_X1 U1325 ( .A1(n565), .A2(n572), .ZN(n1432) );
  NAND3_X1 U1326 ( .A1(n1430), .A2(n1431), .A3(n1432), .ZN(n558) );
  NAND2_X1 U1327 ( .A1(n561), .A2(n570), .ZN(n1433) );
  NAND2_X1 U1328 ( .A1(n561), .A2(n559), .ZN(n1434) );
  NAND2_X1 U1329 ( .A1(n570), .A2(n559), .ZN(n1435) );
  NAND3_X1 U1330 ( .A1(n1433), .A2(n1434), .A3(n1435), .ZN(n556) );
  NAND2_X1 U1331 ( .A1(n578), .A2(n829), .ZN(n1436) );
  NAND2_X1 U1332 ( .A1(n578), .A2(n811), .ZN(n1437) );
  NAND2_X1 U1333 ( .A1(n829), .A2(n811), .ZN(n1438) );
  NAND3_X1 U1334 ( .A1(n1436), .A2(n1437), .A3(n1438), .ZN(n562) );
  CLKBUF_X3 U1335 ( .A(n34), .Z(n1512) );
  BUF_X1 U1336 ( .A(n36), .Z(n1479) );
  XNOR2_X1 U1337 ( .A(n55), .B(a[18]), .ZN(n1439) );
  XOR2_X1 U1338 ( .A(n49), .B(a[18]), .Z(n1440) );
  OR2_X2 U1339 ( .A1(n1439), .A2(n1440), .ZN(n1441) );
  OR2_X2 U1340 ( .A1(n1439), .A2(n1440), .ZN(n1442) );
  XNOR2_X1 U1341 ( .A(n1443), .B(n515), .ZN(n513) );
  XNOR2_X1 U1342 ( .A(n517), .B(n530), .ZN(n1443) );
  AOI21_X1 U1343 ( .B1(n1445), .B2(n133), .A(n1364), .ZN(n1444) );
  CLKBUF_X1 U1344 ( .A(n146), .Z(n1445) );
  CLKBUF_X1 U1345 ( .A(n106), .Z(n1446) );
  BUF_X1 U1346 ( .A(n1), .Z(n1448) );
  XOR2_X1 U1347 ( .A(n300), .B(n299), .Z(n1449) );
  XOR2_X1 U1348 ( .A(n1449), .B(n1321), .Z(product[37]) );
  NAND2_X1 U1349 ( .A1(n300), .A2(n299), .ZN(n1450) );
  NAND2_X1 U1350 ( .A1(n98), .A2(n300), .ZN(n1451) );
  NAND2_X1 U1351 ( .A1(n299), .A2(n1360), .ZN(n1452) );
  XOR2_X1 U1352 ( .A(n680), .B(n298), .Z(n1453) );
  NAND2_X1 U1353 ( .A1(n680), .A2(n298), .ZN(n1454) );
  NAND2_X1 U1354 ( .A1(n1377), .A2(n680), .ZN(n1455) );
  NAND2_X1 U1355 ( .A1(n1377), .A2(n298), .ZN(n1456) );
  NAND2_X1 U1356 ( .A1(n515), .A2(n517), .ZN(n1457) );
  NAND2_X1 U1357 ( .A1(n515), .A2(n530), .ZN(n1458) );
  NAND2_X1 U1358 ( .A1(n517), .A2(n530), .ZN(n1459) );
  NAND3_X1 U1359 ( .A1(n1457), .A2(n1458), .A3(n1459), .ZN(n512) );
  NAND2_X1 U1360 ( .A1(n540), .A2(n536), .ZN(n1460) );
  NAND2_X1 U1361 ( .A1(n540), .A2(n538), .ZN(n1461) );
  NAND2_X1 U1362 ( .A1(n536), .A2(n538), .ZN(n1462) );
  NAND3_X1 U1363 ( .A1(n1460), .A2(n1461), .A3(n1462), .ZN(n518) );
  CLKBUF_X1 U1364 ( .A(n1511), .Z(n1463) );
  CLKBUF_X1 U1365 ( .A(n151), .Z(n1464) );
  INV_X1 U1366 ( .A(n54), .ZN(n1465) );
  INV_X1 U1367 ( .A(n1465), .ZN(n1466) );
  OR2_X2 U1368 ( .A1(n513), .A2(n528), .ZN(n1520) );
  OR2_X1 U1369 ( .A1(n1467), .A2(n1468), .ZN(n48) );
  XNOR2_X1 U1370 ( .A(n43), .B(a[14]), .ZN(n1467) );
  XOR2_X1 U1371 ( .A(n1542), .B(a[14]), .Z(n1468) );
  OR2_X2 U1372 ( .A1(n1467), .A2(n1468), .ZN(n1469) );
  OR2_X2 U1373 ( .A1(n1467), .A2(n1428), .ZN(n1470) );
  BUF_X1 U1374 ( .A(n18), .Z(n1474) );
  AOI21_X1 U1375 ( .B1(n114), .B2(n1498), .A(n111), .ZN(n1471) );
  BUF_X4 U1376 ( .A(n24), .Z(n1472) );
  NAND2_X1 U1377 ( .A1(n1492), .A2(n22), .ZN(n24) );
  CLKBUF_X1 U1378 ( .A(n122), .Z(n1473) );
  NAND2_X1 U1379 ( .A1(n1487), .A2(n16), .ZN(n18) );
  AOI21_X1 U1380 ( .B1(n122), .B2(n1497), .A(n119), .ZN(n1476) );
  NOR2_X1 U1381 ( .A1(n497), .A2(n512), .ZN(n1478) );
  BUF_X2 U1382 ( .A(n36), .Z(n1481) );
  NAND2_X1 U1383 ( .A1(n1488), .A2(n34), .ZN(n36) );
  CLKBUF_X1 U1384 ( .A(n153), .Z(n1482) );
  NAND2_X1 U1385 ( .A1(n1115), .A2(n1514), .ZN(n1483) );
  INV_X2 U1386 ( .A(n668), .ZN(n4) );
  AOI21_X1 U1387 ( .B1(n153), .B2(n126), .A(n127), .ZN(n1485) );
  NOR2_X1 U1388 ( .A1(n497), .A2(n512), .ZN(n177) );
  NOR2_X1 U1389 ( .A1(n359), .A2(n370), .ZN(n128) );
  OR2_X1 U1390 ( .A1(n323), .A2(n330), .ZN(n1498) );
  XOR2_X1 U1391 ( .A(n13), .B(a[4]), .Z(n1487) );
  XOR2_X1 U1392 ( .A(n31), .B(a[10]), .Z(n1488) );
  XOR2_X1 U1393 ( .A(n7), .B(a[2]), .Z(n1489) );
  NAND2_X2 U1394 ( .A1(n1490), .A2(n52), .ZN(n54) );
  XOR2_X1 U1395 ( .A(n49), .B(a[16]), .Z(n1490) );
  NAND2_X1 U1396 ( .A1(n1491), .A2(n1308), .ZN(n42) );
  XOR2_X1 U1397 ( .A(n1542), .B(a[12]), .Z(n1491) );
  XOR2_X1 U1398 ( .A(n19), .B(a[6]), .Z(n1492) );
  OAI21_X1 U1399 ( .B1(n152), .B2(n143), .A(n144), .ZN(n142) );
  NAND2_X1 U1400 ( .A1(n270), .A2(n124), .ZN(n68) );
  INV_X1 U1401 ( .A(n123), .ZN(n270) );
  INV_X1 U1402 ( .A(n140), .ZN(n273) );
  INV_X1 U1403 ( .A(n171), .ZN(n279) );
  XOR2_X1 U1404 ( .A(n168), .B(n76), .Z(product[20]) );
  AOI21_X1 U1405 ( .B1(n173), .B2(n279), .A(n170), .ZN(n168) );
  XOR2_X1 U1406 ( .A(n137), .B(n70), .Z(product[26]) );
  NAND2_X1 U1407 ( .A1(n1234), .A2(n136), .ZN(n70) );
  AOI21_X1 U1408 ( .B1(n142), .B2(n273), .A(n139), .ZN(n137) );
  XOR2_X1 U1409 ( .A(n206), .B(n82), .Z(product[14]) );
  NAND2_X1 U1410 ( .A1(n284), .A2(n205), .ZN(n82) );
  AOI21_X1 U1411 ( .B1(n211), .B2(n285), .A(n208), .ZN(n206) );
  XOR2_X1 U1412 ( .A(n152), .B(n73), .Z(product[23]) );
  NAND2_X1 U1413 ( .A1(n275), .A2(n1464), .ZN(n73) );
  XOR2_X1 U1414 ( .A(n193), .B(n80), .Z(product[16]) );
  NAND2_X1 U1415 ( .A1(n1233), .A2(n188), .ZN(n80) );
  XOR2_X1 U1416 ( .A(n163), .B(n75), .Z(product[21]) );
  INV_X1 U1417 ( .A(n234), .ZN(n233) );
  XNOR2_X1 U1418 ( .A(n160), .B(n74), .ZN(product[22]) );
  NAND2_X1 U1419 ( .A1(n276), .A2(n159), .ZN(n74) );
  XNOR2_X1 U1420 ( .A(n173), .B(n77), .ZN(product[19]) );
  NAND2_X1 U1421 ( .A1(n279), .A2(n1279), .ZN(n77) );
  XNOR2_X1 U1422 ( .A(n149), .B(n72), .ZN(product[24]) );
  NAND2_X1 U1423 ( .A1(n274), .A2(n1313), .ZN(n72) );
  XNOR2_X1 U1424 ( .A(n130), .B(n69), .ZN(product[27]) );
  NAND2_X1 U1425 ( .A1(n271), .A2(n129), .ZN(n69) );
  INV_X1 U1426 ( .A(n128), .ZN(n271) );
  XNOR2_X1 U1427 ( .A(n142), .B(n71), .ZN(product[25]) );
  NAND2_X1 U1428 ( .A1(n273), .A2(n141), .ZN(n71) );
  XNOR2_X1 U1429 ( .A(n179), .B(n78), .ZN(product[18]) );
  NAND2_X1 U1430 ( .A1(n280), .A2(n178), .ZN(n78) );
  INV_X1 U1431 ( .A(n1478), .ZN(n280) );
  INV_X1 U1432 ( .A(n172), .ZN(n170) );
  INV_X1 U1433 ( .A(n141), .ZN(n139) );
  INV_X1 U1434 ( .A(n113), .ZN(n111) );
  NAND2_X1 U1435 ( .A1(n1495), .A2(n1494), .ZN(n222) );
  AOI21_X1 U1436 ( .B1(n1495), .B2(n230), .A(n225), .ZN(n223) );
  INV_X1 U1437 ( .A(n227), .ZN(n225) );
  AOI21_X1 U1438 ( .B1(n239), .B2(n1496), .A(n236), .ZN(n234) );
  INV_X1 U1439 ( .A(n238), .ZN(n236) );
  AOI21_X1 U1440 ( .B1(n1473), .B2(n1497), .A(n119), .ZN(n117) );
  INV_X1 U1441 ( .A(n121), .ZN(n119) );
  NOR2_X1 U1442 ( .A1(n383), .A2(n396), .ZN(n140) );
  NAND2_X1 U1443 ( .A1(n268), .A2(n116), .ZN(n66) );
  INV_X1 U1444 ( .A(n115), .ZN(n268) );
  NAND2_X1 U1445 ( .A1(n266), .A2(n108), .ZN(n64) );
  INV_X1 U1446 ( .A(n107), .ZN(n266) );
  NAND2_X1 U1447 ( .A1(n383), .A2(n396), .ZN(n141) );
  INV_X1 U1448 ( .A(n232), .ZN(n230) );
  INV_X1 U1449 ( .A(n209), .ZN(n285) );
  NAND2_X1 U1450 ( .A1(n411), .A2(n426), .ZN(n151) );
  NAND2_X1 U1451 ( .A1(n1497), .A2(n121), .ZN(n67) );
  NAND2_X1 U1452 ( .A1(n1499), .A2(n105), .ZN(n63) );
  NAND2_X1 U1453 ( .A1(n1498), .A2(n113), .ZN(n65) );
  XOR2_X1 U1454 ( .A(n228), .B(n86), .Z(product[10]) );
  NAND2_X1 U1455 ( .A1(n1495), .A2(n227), .ZN(n86) );
  AOI21_X1 U1456 ( .B1(n233), .B2(n1494), .A(n230), .ZN(n228) );
  XOR2_X1 U1457 ( .A(n201), .B(n81), .Z(product[15]) );
  AOI21_X1 U1458 ( .B1(n211), .B2(n202), .A(n1522), .ZN(n201) );
  INV_X1 U1459 ( .A(n1526), .ZN(n200) );
  XOR2_X1 U1460 ( .A(n220), .B(n85), .Z(product[11]) );
  NAND2_X1 U1461 ( .A1(n287), .A2(n219), .ZN(n85) );
  INV_X1 U1462 ( .A(n218), .ZN(n287) );
  NOR2_X1 U1463 ( .A1(n349), .A2(n358), .ZN(n123) );
  XNOR2_X1 U1464 ( .A(n211), .B(n83), .ZN(product[13]) );
  NAND2_X1 U1465 ( .A1(n285), .A2(n210), .ZN(n83) );
  NOR2_X1 U1466 ( .A1(n479), .A2(n496), .ZN(n171) );
  XNOR2_X1 U1467 ( .A(n239), .B(n88), .ZN(product[8]) );
  NAND2_X1 U1468 ( .A1(n1496), .A2(n238), .ZN(n88) );
  XNOR2_X1 U1469 ( .A(n186), .B(n79), .ZN(product[17]) );
  INV_X1 U1470 ( .A(n1528), .ZN(n185) );
  XNOR2_X1 U1471 ( .A(n233), .B(n87), .ZN(product[9]) );
  NAND2_X1 U1472 ( .A1(n1494), .A2(n232), .ZN(n87) );
  XNOR2_X1 U1473 ( .A(n217), .B(n84), .ZN(product[12]) );
  NAND2_X1 U1474 ( .A1(n286), .A2(n216), .ZN(n84) );
  OAI21_X1 U1475 ( .B1(n220), .B2(n218), .A(n219), .ZN(n217) );
  NAND2_X1 U1476 ( .A1(n557), .A2(n568), .ZN(n205) );
  NAND2_X1 U1477 ( .A1(n497), .A2(n512), .ZN(n178) );
  NAND2_X1 U1478 ( .A1(n349), .A2(n358), .ZN(n124) );
  NAND2_X1 U1479 ( .A1(n359), .A2(n370), .ZN(n129) );
  NAND2_X1 U1480 ( .A1(n427), .A2(n442), .ZN(n159) );
  INV_X1 U1481 ( .A(n210), .ZN(n208) );
  INV_X1 U1482 ( .A(n1268), .ZN(n188) );
  AOI21_X1 U1483 ( .B1(n1501), .B2(n255), .A(n252), .ZN(n250) );
  INV_X1 U1484 ( .A(n254), .ZN(n252) );
  OR2_X1 U1485 ( .A1(n609), .A2(n616), .ZN(n1494) );
  OAI21_X1 U1486 ( .B1(n256), .B2(n258), .A(n257), .ZN(n255) );
  OR2_X1 U1487 ( .A1(n601), .A2(n608), .ZN(n1495) );
  AOI21_X1 U1488 ( .B1(n1502), .B2(n247), .A(n244), .ZN(n242) );
  INV_X1 U1489 ( .A(n246), .ZN(n244) );
  NOR2_X1 U1490 ( .A1(n591), .A2(n600), .ZN(n218) );
  OAI21_X1 U1491 ( .B1(n248), .B2(n250), .A(n249), .ZN(n247) );
  NAND2_X1 U1492 ( .A1(n291), .A2(n241), .ZN(n89) );
  INV_X1 U1493 ( .A(n240), .ZN(n291) );
  XOR2_X1 U1494 ( .A(n91), .B(n250), .Z(product[5]) );
  NAND2_X1 U1495 ( .A1(n293), .A2(n249), .ZN(n91) );
  INV_X1 U1496 ( .A(n248), .ZN(n293) );
  NAND2_X1 U1497 ( .A1(n591), .A2(n600), .ZN(n219) );
  NOR2_X1 U1498 ( .A1(n569), .A2(n580), .ZN(n209) );
  NOR2_X1 U1499 ( .A1(n331), .A2(n338), .ZN(n115) );
  NOR2_X1 U1500 ( .A1(n317), .A2(n322), .ZN(n107) );
  NAND2_X1 U1501 ( .A1(n569), .A2(n580), .ZN(n210) );
  INV_X1 U1502 ( .A(n259), .ZN(n258) );
  OAI21_X1 U1503 ( .B1(n260), .B2(n263), .A(n261), .ZN(n259) );
  OR2_X1 U1504 ( .A1(n617), .A2(n622), .ZN(n1496) );
  XNOR2_X1 U1505 ( .A(n92), .B(n255), .ZN(product[4]) );
  NAND2_X1 U1506 ( .A1(n1501), .A2(n254), .ZN(n92) );
  OR2_X1 U1507 ( .A1(n339), .A2(n348), .ZN(n1497) );
  XNOR2_X1 U1508 ( .A(n90), .B(n247), .ZN(product[6]) );
  NAND2_X1 U1509 ( .A1(n1502), .A2(n246), .ZN(n90) );
  NAND2_X1 U1510 ( .A1(n323), .A2(n330), .ZN(n113) );
  NAND2_X1 U1511 ( .A1(n617), .A2(n622), .ZN(n238) );
  NAND2_X1 U1512 ( .A1(n311), .A2(n316), .ZN(n105) );
  NAND2_X1 U1513 ( .A1(n339), .A2(n348), .ZN(n121) );
  NAND2_X1 U1514 ( .A1(n331), .A2(n338), .ZN(n116) );
  NAND2_X1 U1515 ( .A1(n317), .A2(n322), .ZN(n108) );
  NAND2_X1 U1516 ( .A1(n601), .A2(n608), .ZN(n227) );
  OR2_X1 U1517 ( .A1(n311), .A2(n316), .ZN(n1499) );
  NAND2_X1 U1518 ( .A1(n581), .A2(n590), .ZN(n216) );
  XOR2_X1 U1519 ( .A(n93), .B(n258), .Z(product[3]) );
  NAND2_X1 U1520 ( .A1(n295), .A2(n257), .ZN(n93) );
  INV_X1 U1521 ( .A(n256), .ZN(n295) );
  OR2_X1 U1522 ( .A1(n543), .A2(n556), .ZN(n1523) );
  XOR2_X1 U1523 ( .A(n94), .B(n263), .Z(product[2]) );
  NAND2_X1 U1524 ( .A1(n296), .A2(n261), .ZN(n94) );
  INV_X1 U1525 ( .A(n260), .ZN(n296) );
  NOR2_X1 U1526 ( .A1(n633), .A2(n636), .ZN(n248) );
  XNOR2_X1 U1527 ( .A(n1500), .B(n815), .ZN(n607) );
  XNOR2_X1 U1528 ( .A(n870), .B(n779), .ZN(n1500) );
  NAND2_X1 U1529 ( .A1(n639), .A2(n678), .ZN(n257) );
  NOR2_X1 U1530 ( .A1(n639), .A2(n678), .ZN(n256) );
  NOR2_X1 U1531 ( .A1(n878), .A2(n859), .ZN(n260) );
  NAND2_X1 U1532 ( .A1(n679), .A2(n879), .ZN(n263) );
  NAND2_X1 U1533 ( .A1(n878), .A2(n859), .ZN(n261) );
  OR2_X1 U1534 ( .A1(n637), .A2(n638), .ZN(n1501) );
  INV_X1 U1535 ( .A(n394), .ZN(n395) );
  INV_X1 U1536 ( .A(n328), .ZN(n329) );
  INV_X1 U1537 ( .A(n424), .ZN(n425) );
  NOR2_X1 U1538 ( .A1(n623), .A2(n628), .ZN(n240) );
  INV_X1 U1539 ( .A(n105), .ZN(n103) );
  INV_X1 U1540 ( .A(n298), .ZN(n299) );
  NAND2_X1 U1541 ( .A1(n629), .A2(n632), .ZN(n246) );
  OR2_X1 U1542 ( .A1(n629), .A2(n632), .ZN(n1502) );
  NAND2_X1 U1543 ( .A1(n623), .A2(n628), .ZN(n241) );
  OAI22_X1 U1544 ( .A1(n1508), .A2(n1086), .B1(n1085), .B2(n4), .ZN(n877) );
  OAI22_X1 U1545 ( .A1(n1272), .A2(n1088), .B1(n1087), .B2(n4), .ZN(n879) );
  OAI22_X1 U1546 ( .A1(n1510), .A2(n1149), .B1(n1089), .B2(n4), .ZN(n679) );
  OR2_X1 U1547 ( .A1(n1547), .A2(n1149), .ZN(n1089) );
  OAI22_X1 U1548 ( .A1(n1272), .A2(n1087), .B1(n1086), .B2(n4), .ZN(n878) );
  INV_X1 U1549 ( .A(n314), .ZN(n315) );
  INV_X1 U1550 ( .A(n667), .ZN(n860) );
  OAI22_X1 U1551 ( .A1(n1237), .A2(n1508), .B1(n1073), .B2(n4), .ZN(n865) );
  INV_X1 U1552 ( .A(n458), .ZN(n459) );
  OAI22_X1 U1553 ( .A1(n1510), .A2(n1257), .B1(n1077), .B2(n4), .ZN(n869) );
  OAI22_X1 U1554 ( .A1(n1262), .A2(n1509), .B1(n1069), .B2(n4), .ZN(n667) );
  OAI22_X1 U1555 ( .A1(n1510), .A2(n1076), .B1(n1075), .B2(n4), .ZN(n867) );
  AND2_X1 U1556 ( .A1(n1547), .A2(n662), .ZN(n839) );
  OAI22_X1 U1557 ( .A1(n1272), .A2(n1085), .B1(n1084), .B2(n4), .ZN(n876) );
  OAI22_X1 U1558 ( .A1(n1508), .A2(n1084), .B1(n1083), .B2(n4), .ZN(n875) );
  XNOR2_X1 U1559 ( .A(n1552), .B(n1329), .ZN(n892) );
  XNOR2_X1 U1560 ( .A(n1342), .B(n1330), .ZN(n891) );
  XNOR2_X1 U1561 ( .A(n1551), .B(n1329), .ZN(n893) );
  XNOR2_X1 U1562 ( .A(n1343), .B(n1329), .ZN(n894) );
  XNOR2_X1 U1563 ( .A(n1352), .B(n1545), .ZN(n895) );
  XNOR2_X1 U1564 ( .A(n1325), .B(n1545), .ZN(n896) );
  XNOR2_X1 U1565 ( .A(n1555), .B(n1330), .ZN(n889) );
  XNOR2_X1 U1566 ( .A(n1350), .B(n1329), .ZN(n888) );
  XNOR2_X1 U1567 ( .A(n1554), .B(n1329), .ZN(n890) );
  XNOR2_X1 U1568 ( .A(n1548), .B(n1545), .ZN(n897) );
  XNOR2_X1 U1569 ( .A(n1108), .B(n1330), .ZN(n898) );
  XNOR2_X1 U1570 ( .A(n1314), .B(n1330), .ZN(n887) );
  XNOR2_X1 U1571 ( .A(n1323), .B(n1329), .ZN(n886) );
  XNOR2_X1 U1572 ( .A(n1559), .B(n1330), .ZN(n885) );
  XNOR2_X1 U1573 ( .A(n1560), .B(n1329), .ZN(n884) );
  XNOR2_X1 U1574 ( .A(n1318), .B(n1330), .ZN(n883) );
  XNOR2_X1 U1575 ( .A(n1354), .B(n1329), .ZN(n882) );
  XNOR2_X1 U1576 ( .A(n1351), .B(n1330), .ZN(n881) );
  AND2_X1 U1577 ( .A1(n1547), .A2(n665), .ZN(n859) );
  OR2_X1 U1578 ( .A1(n1547), .A2(n1147), .ZN(n1047) );
  BUF_X1 U1579 ( .A(n1105), .Z(n1549) );
  BUF_X1 U1580 ( .A(n1092), .Z(n1562) );
  INV_X1 U1581 ( .A(n661), .ZN(n820) );
  INV_X1 U1582 ( .A(n655), .ZN(n780) );
  INV_X1 U1583 ( .A(n304), .ZN(n305) );
  AND2_X1 U1584 ( .A1(n1547), .A2(n1440), .ZN(n699) );
  OAI22_X1 U1585 ( .A1(n1508), .A2(n1071), .B1(n1070), .B2(n4), .ZN(n862) );
  OAI22_X1 U1586 ( .A1(n1272), .A2(n1072), .B1(n1071), .B2(n4), .ZN(n863) );
  INV_X1 U1587 ( .A(n649), .ZN(n740) );
  INV_X1 U1588 ( .A(n643), .ZN(n700) );
  INV_X1 U1589 ( .A(n346), .ZN(n347) );
  OAI22_X1 U1590 ( .A1(n1272), .A2(n1077), .B1(n1076), .B2(n4), .ZN(n868) );
  INV_X1 U1591 ( .A(n652), .ZN(n760) );
  INV_X1 U1592 ( .A(n646), .ZN(n720) );
  OAI22_X1 U1593 ( .A1(n1510), .A2(n1080), .B1(n1079), .B2(n4), .ZN(n871) );
  AND2_X1 U1594 ( .A1(n1547), .A2(n1428), .ZN(n739) );
  OAI22_X1 U1595 ( .A1(n1510), .A2(n1075), .B1(n1074), .B2(n4), .ZN(n866) );
  OAI22_X1 U1596 ( .A1(n1272), .A2(n1082), .B1(n1081), .B2(n4), .ZN(n873) );
  OAI22_X1 U1597 ( .A1(n1272), .A2(n1083), .B1(n1082), .B2(n4), .ZN(n874) );
  AND2_X1 U1598 ( .A1(n1547), .A2(n659), .ZN(n819) );
  OAI22_X1 U1599 ( .A1(n1508), .A2(n1073), .B1(n1072), .B2(n4), .ZN(n864) );
  AND2_X1 U1600 ( .A1(n1547), .A2(n644), .ZN(n719) );
  INV_X1 U1601 ( .A(n664), .ZN(n840) );
  OAI22_X1 U1602 ( .A1(n1508), .A2(n1070), .B1(n1262), .B2(n4), .ZN(n861) );
  AND2_X1 U1603 ( .A1(n1547), .A2(n656), .ZN(n799) );
  OAI22_X1 U1604 ( .A1(n1510), .A2(n1081), .B1(n1080), .B2(n4), .ZN(n872) );
  INV_X1 U1605 ( .A(n640), .ZN(n680) );
  INV_X1 U1606 ( .A(n368), .ZN(n369) );
  XNOR2_X1 U1607 ( .A(n1546), .B(n1330), .ZN(n899) );
  INV_X1 U1608 ( .A(n658), .ZN(n800) );
  INV_X1 U1609 ( .A(n55), .ZN(n1140) );
  OR2_X1 U1610 ( .A1(n1546), .A2(n1142), .ZN(n942) );
  OR2_X1 U1611 ( .A1(n1546), .A2(n1141), .ZN(n921) );
  OR2_X1 U1612 ( .A1(n1547), .A2(n1144), .ZN(n984) );
  OR2_X1 U1613 ( .A1(n1547), .A2(n1140), .ZN(n900) );
  OR2_X1 U1614 ( .A1(n1547), .A2(n1146), .ZN(n1026) );
  XNOR2_X1 U1615 ( .A(n1307), .B(n1329), .ZN(n880) );
  BUF_X2 U1616 ( .A(n61), .Z(n1547) );
  AND2_X1 U1617 ( .A1(n1547), .A2(n668), .ZN(product[0]) );
  XNOR2_X1 U1618 ( .A(n1), .B(a[2]), .ZN(n9) );
  NAND2_X1 U1619 ( .A1(n1119), .A2(n1357), .ZN(n6) );
  XNOR2_X1 U1620 ( .A(n43), .B(a[16]), .ZN(n52) );
  XNOR2_X1 U1621 ( .A(n25), .B(a[10]), .ZN(n34) );
  XNOR2_X1 U1622 ( .A(n19), .B(a[8]), .ZN(n28) );
  BUF_X4 U1623 ( .A(n1305), .Z(n1516) );
  XNOR2_X1 U1624 ( .A(n7), .B(a[4]), .ZN(n16) );
  BUF_X4 U1625 ( .A(n22), .Z(n1517) );
  XNOR2_X1 U1626 ( .A(n13), .B(a[6]), .ZN(n22) );
  XNOR2_X1 U1627 ( .A(n1542), .B(a[14]), .ZN(n1518) );
  XNOR2_X1 U1628 ( .A(n1542), .B(a[14]), .ZN(n1519) );
  OR2_X1 U1629 ( .A1(n1547), .A2(n1143), .ZN(n963) );
  CLKBUF_X1 U1630 ( .A(n167), .Z(n1521) );
  OAI21_X1 U1631 ( .B1(n204), .B2(n210), .A(n205), .ZN(n1522) );
  NAND2_X1 U1632 ( .A1(n609), .A2(n616), .ZN(n232) );
  NOR2_X1 U1633 ( .A1(n461), .A2(n478), .ZN(n1525) );
  OAI21_X1 U1634 ( .B1(n215), .B2(n219), .A(n216), .ZN(n214) );
  NOR2_X1 U1635 ( .A1(n215), .A2(n218), .ZN(n213) );
  INV_X1 U1636 ( .A(n215), .ZN(n286) );
  AOI21_X1 U1637 ( .B1(n173), .B2(n164), .A(n1418), .ZN(n163) );
  AND2_X1 U1638 ( .A1(n543), .A2(n556), .ZN(n1526) );
  OR2_X1 U1639 ( .A1(n1546), .A2(n1145), .ZN(n1005) );
  NAND2_X1 U1640 ( .A1(n479), .A2(n496), .ZN(n172) );
  AND2_X1 U1641 ( .A1(n1547), .A2(n1533), .ZN(n759) );
  NAND2_X1 U1642 ( .A1(n278), .A2(n1521), .ZN(n76) );
  NOR2_X1 U1643 ( .A1(n410), .A2(n397), .ZN(n1527) );
  NOR2_X1 U1644 ( .A1(n397), .A2(n410), .ZN(n147) );
  XNOR2_X1 U1645 ( .A(n1307), .B(n1348), .ZN(n901) );
  XNOR2_X1 U1646 ( .A(n1351), .B(n1348), .ZN(n902) );
  XNOR2_X1 U1647 ( .A(n1318), .B(n1348), .ZN(n904) );
  XNOR2_X1 U1648 ( .A(n1355), .B(n1348), .ZN(n903) );
  XNOR2_X1 U1649 ( .A(n1560), .B(n1348), .ZN(n905) );
  XNOR2_X1 U1650 ( .A(n1559), .B(n1348), .ZN(n906) );
  XNOR2_X1 U1651 ( .A(n1323), .B(n1348), .ZN(n907) );
  XNOR2_X1 U1652 ( .A(n1314), .B(n1348), .ZN(n908) );
  XNOR2_X1 U1653 ( .A(n1350), .B(n1348), .ZN(n909) );
  XNOR2_X1 U1654 ( .A(n1555), .B(n1348), .ZN(n910) );
  XNOR2_X1 U1655 ( .A(n1554), .B(n1544), .ZN(n911) );
  XNOR2_X1 U1656 ( .A(n1552), .B(n1544), .ZN(n913) );
  XNOR2_X1 U1657 ( .A(n1553), .B(n1544), .ZN(n912) );
  XNOR2_X1 U1658 ( .A(n1551), .B(n1544), .ZN(n914) );
  XNOR2_X1 U1659 ( .A(n1326), .B(n1544), .ZN(n917) );
  XNOR2_X1 U1660 ( .A(n1548), .B(n1544), .ZN(n918) );
  XNOR2_X1 U1661 ( .A(n1353), .B(n1544), .ZN(n916) );
  XNOR2_X1 U1662 ( .A(n1546), .B(n1348), .ZN(n920) );
  XNOR2_X1 U1663 ( .A(n1344), .B(n1544), .ZN(n915) );
  INV_X1 U1664 ( .A(n49), .ZN(n1141) );
  XNOR2_X1 U1665 ( .A(n1346), .B(n1544), .ZN(n919) );
  NOR2_X1 U1666 ( .A1(n461), .A2(n478), .ZN(n166) );
  AND2_X1 U1667 ( .A1(n513), .A2(n528), .ZN(n1528) );
  OR2_X1 U1668 ( .A1(n1547), .A2(n1148), .ZN(n1068) );
  XOR2_X1 U1669 ( .A(n551), .B(n564), .Z(n1529) );
  XOR2_X1 U1670 ( .A(n562), .B(n1529), .Z(n547) );
  NAND2_X1 U1671 ( .A1(n562), .A2(n551), .ZN(n1530) );
  NAND2_X1 U1672 ( .A1(n562), .A2(n564), .ZN(n1531) );
  NAND2_X1 U1673 ( .A1(n551), .A2(n564), .ZN(n1532) );
  NAND3_X1 U1674 ( .A1(n1530), .A2(n1531), .A3(n1532), .ZN(n546) );
  NOR2_X1 U1675 ( .A1(n131), .A2(n128), .ZN(n126) );
  NAND2_X1 U1676 ( .A1(n277), .A2(n162), .ZN(n75) );
  XNOR2_X1 U1677 ( .A(n1351), .B(n1304), .ZN(n923) );
  XNOR2_X1 U1678 ( .A(n1564), .B(n1304), .ZN(n922) );
  XNOR2_X1 U1679 ( .A(n1354), .B(n1304), .ZN(n924) );
  XNOR2_X1 U1680 ( .A(n1560), .B(n1304), .ZN(n926) );
  XNOR2_X1 U1681 ( .A(n1318), .B(n1304), .ZN(n925) );
  XNOR2_X1 U1682 ( .A(n1559), .B(n1304), .ZN(n927) );
  XNOR2_X1 U1683 ( .A(n1323), .B(n1543), .ZN(n928) );
  XNOR2_X1 U1684 ( .A(n1314), .B(n1543), .ZN(n929) );
  XNOR2_X1 U1685 ( .A(n787), .B(n715), .ZN(n477) );
  OR2_X1 U1686 ( .A1(n787), .A2(n715), .ZN(n476) );
  XNOR2_X1 U1687 ( .A(n1350), .B(n1543), .ZN(n930) );
  XNOR2_X1 U1688 ( .A(n1337), .B(n1543), .ZN(n932) );
  XNOR2_X1 U1689 ( .A(n1555), .B(n1543), .ZN(n931) );
  XNOR2_X1 U1690 ( .A(n1553), .B(n1543), .ZN(n933) );
  XNOR2_X1 U1691 ( .A(n1551), .B(n1543), .ZN(n935) );
  XNOR2_X1 U1692 ( .A(n1552), .B(n1543), .ZN(n934) );
  XNOR2_X1 U1693 ( .A(n1546), .B(n1543), .ZN(n941) );
  XNOR2_X1 U1694 ( .A(n1550), .B(n1543), .ZN(n936) );
  XNOR2_X1 U1695 ( .A(n1347), .B(n1543), .ZN(n940) );
  XNOR2_X1 U1696 ( .A(n1548), .B(n1543), .ZN(n939) );
  XNOR2_X1 U1697 ( .A(n1326), .B(n1543), .ZN(n938) );
  INV_X1 U1698 ( .A(n1543), .ZN(n1142) );
  XNOR2_X1 U1699 ( .A(n1352), .B(n1543), .ZN(n937) );
  BUF_X4 U1700 ( .A(n43), .Z(n1543) );
  INV_X1 U1701 ( .A(n1445), .ZN(n144) );
  NOR2_X1 U1702 ( .A1(n1478), .A2(n180), .ZN(n175) );
  XNOR2_X1 U1703 ( .A(n1564), .B(n1539), .ZN(n1006) );
  INV_X1 U1704 ( .A(n1539), .ZN(n1146) );
  XNOR2_X1 U1705 ( .A(n1355), .B(n1539), .ZN(n1008) );
  XNOR2_X1 U1706 ( .A(n1563), .B(n1539), .ZN(n1007) );
  XNOR2_X1 U1707 ( .A(n1546), .B(n1539), .ZN(n1025) );
  XNOR2_X1 U1708 ( .A(n1346), .B(n1539), .ZN(n1024) );
  XNOR2_X1 U1709 ( .A(n1561), .B(n1539), .ZN(n1009) );
  XNOR2_X1 U1710 ( .A(n1350), .B(n1539), .ZN(n1014) );
  XNOR2_X1 U1711 ( .A(n1557), .B(n1539), .ZN(n1013) );
  XNOR2_X1 U1712 ( .A(n1558), .B(n1539), .ZN(n1012) );
  XNOR2_X1 U1713 ( .A(n1352), .B(n1539), .ZN(n1021) );
  XNOR2_X1 U1714 ( .A(n1344), .B(n1539), .ZN(n1020) );
  XNOR2_X1 U1715 ( .A(n1345), .B(n1539), .ZN(n1023) );
  XNOR2_X1 U1716 ( .A(n1356), .B(n1539), .ZN(n1022) );
  XNOR2_X1 U1717 ( .A(n1559), .B(n1539), .ZN(n1011) );
  XNOR2_X1 U1718 ( .A(n1552), .B(n1539), .ZN(n1018) );
  XNOR2_X1 U1719 ( .A(n1551), .B(n1539), .ZN(n1019) );
  XNOR2_X1 U1720 ( .A(n1560), .B(n1539), .ZN(n1010) );
  XNOR2_X1 U1721 ( .A(n1555), .B(n1539), .ZN(n1015) );
  XNOR2_X1 U1722 ( .A(n1553), .B(n19), .ZN(n1017) );
  XNOR2_X1 U1723 ( .A(n1337), .B(n1539), .ZN(n1016) );
  XNOR2_X1 U1724 ( .A(n1564), .B(n1365), .ZN(n943) );
  XNOR2_X1 U1725 ( .A(n1351), .B(n1365), .ZN(n944) );
  XNOR2_X1 U1726 ( .A(n1318), .B(n1365), .ZN(n946) );
  XNOR2_X1 U1727 ( .A(n1355), .B(n1365), .ZN(n945) );
  XNOR2_X1 U1728 ( .A(n1560), .B(n1365), .ZN(n947) );
  XNOR2_X1 U1729 ( .A(n1559), .B(n1365), .ZN(n948) );
  XNOR2_X1 U1730 ( .A(n1350), .B(n1365), .ZN(n951) );
  XNOR2_X1 U1731 ( .A(n1557), .B(n1365), .ZN(n950) );
  XNOR2_X1 U1732 ( .A(n1558), .B(n1365), .ZN(n949) );
  XNOR2_X1 U1733 ( .A(n1555), .B(n1365), .ZN(n952) );
  XNOR2_X1 U1734 ( .A(n1551), .B(n1365), .ZN(n956) );
  INV_X1 U1735 ( .A(n1365), .ZN(n1143) );
  XNOR2_X1 U1736 ( .A(n1552), .B(n1365), .ZN(n955) );
  XNOR2_X1 U1737 ( .A(n1344), .B(n1365), .ZN(n957) );
  XNOR2_X1 U1738 ( .A(n1345), .B(n1365), .ZN(n960) );
  XNOR2_X1 U1739 ( .A(n1337), .B(n1365), .ZN(n953) );
  XNOR2_X1 U1740 ( .A(n1553), .B(n1365), .ZN(n954) );
  XNOR2_X1 U1741 ( .A(n1546), .B(n1365), .ZN(n962) );
  XNOR2_X1 U1742 ( .A(n1325), .B(n1365), .ZN(n959) );
  XNOR2_X1 U1743 ( .A(n1347), .B(n1365), .ZN(n961) );
  XNOR2_X1 U1744 ( .A(n1352), .B(n1365), .ZN(n958) );
  INV_X1 U1745 ( .A(n1285), .ZN(n276) );
  NAND2_X1 U1746 ( .A1(n156), .A2(n164), .ZN(n154) );
  INV_X1 U1747 ( .A(n145), .ZN(n143) );
  NAND2_X1 U1748 ( .A1(n815), .A2(n1339), .ZN(n1534) );
  NAND2_X1 U1749 ( .A1(n815), .A2(n779), .ZN(n1535) );
  NAND2_X1 U1750 ( .A1(n870), .A2(n779), .ZN(n1536) );
  NAND3_X1 U1751 ( .A1(n1534), .A2(n1535), .A3(n1536), .ZN(n606) );
  AND2_X1 U1752 ( .A1(n1547), .A2(n653), .ZN(n779) );
  OAI22_X1 U1753 ( .A1(n1272), .A2(n1079), .B1(n1078), .B2(n4), .ZN(n870) );
  NAND2_X1 U1754 ( .A1(n461), .A2(n478), .ZN(n167) );
  XNOR2_X1 U1755 ( .A(n1550), .B(n1333), .ZN(n1062) );
  INV_X1 U1756 ( .A(n1333), .ZN(n1148) );
  XNOR2_X1 U1757 ( .A(n1553), .B(n1333), .ZN(n1059) );
  XNOR2_X1 U1758 ( .A(n1560), .B(n1537), .ZN(n1052) );
  XNOR2_X1 U1759 ( .A(n1561), .B(n1537), .ZN(n1051) );
  XNOR2_X1 U1760 ( .A(n1356), .B(n1333), .ZN(n1064) );
  XNOR2_X1 U1761 ( .A(n1353), .B(n1333), .ZN(n1063) );
  XNOR2_X1 U1762 ( .A(n1354), .B(n1537), .ZN(n1050) );
  XNOR2_X1 U1763 ( .A(n1350), .B(n1537), .ZN(n1056) );
  XNOR2_X1 U1764 ( .A(n1557), .B(n1333), .ZN(n1055) );
  XNOR2_X1 U1765 ( .A(n1554), .B(n1537), .ZN(n1058) );
  XNOR2_X1 U1766 ( .A(n1563), .B(n1537), .ZN(n1049) );
  XNOR2_X1 U1767 ( .A(n1551), .B(n1537), .ZN(n1061) );
  XNOR2_X1 U1768 ( .A(n1552), .B(n1537), .ZN(n1060) );
  XNOR2_X1 U1769 ( .A(n1555), .B(n1537), .ZN(n1057) );
  XNOR2_X1 U1770 ( .A(n1345), .B(n1333), .ZN(n1065) );
  XNOR2_X1 U1771 ( .A(n1546), .B(n1333), .ZN(n1067) );
  XNOR2_X1 U1772 ( .A(n1558), .B(n1537), .ZN(n1054) );
  XNOR2_X1 U1773 ( .A(n1346), .B(n1333), .ZN(n1066) );
  XNOR2_X1 U1774 ( .A(n1559), .B(n1537), .ZN(n1053) );
  XNOR2_X1 U1775 ( .A(n1564), .B(n1537), .ZN(n1048) );
  XNOR2_X1 U1776 ( .A(n1564), .B(n1541), .ZN(n964) );
  XNOR2_X1 U1777 ( .A(n1351), .B(n1541), .ZN(n965) );
  XNOR2_X1 U1778 ( .A(n1354), .B(n1541), .ZN(n966) );
  XNOR2_X1 U1779 ( .A(n1318), .B(n1541), .ZN(n967) );
  XNOR2_X1 U1780 ( .A(n1560), .B(n1541), .ZN(n968) );
  XNOR2_X1 U1781 ( .A(n1350), .B(n1541), .ZN(n972) );
  XNOR2_X1 U1782 ( .A(n1559), .B(n1541), .ZN(n969) );
  XNOR2_X1 U1783 ( .A(n1558), .B(n1541), .ZN(n970) );
  XNOR2_X1 U1784 ( .A(n1557), .B(n1541), .ZN(n971) );
  INV_X1 U1785 ( .A(n1541), .ZN(n1144) );
  XNOR2_X1 U1786 ( .A(n1551), .B(n1541), .ZN(n977) );
  XNOR2_X1 U1787 ( .A(n1546), .B(n1541), .ZN(n983) );
  XNOR2_X1 U1788 ( .A(n1552), .B(n1541), .ZN(n976) );
  XNOR2_X1 U1789 ( .A(n1555), .B(n1541), .ZN(n973) );
  XNOR2_X1 U1790 ( .A(n1337), .B(n1541), .ZN(n974) );
  XNOR2_X1 U1791 ( .A(n1346), .B(n1541), .ZN(n982) );
  XNOR2_X1 U1792 ( .A(n1553), .B(n1541), .ZN(n975) );
  XNOR2_X1 U1793 ( .A(n1550), .B(n1541), .ZN(n978) );
  XNOR2_X1 U1794 ( .A(n1353), .B(n1541), .ZN(n979) );
  XNOR2_X1 U1795 ( .A(n1356), .B(n1541), .ZN(n980) );
  XNOR2_X1 U1796 ( .A(n1345), .B(n1541), .ZN(n981) );
  INV_X1 U1797 ( .A(n1538), .ZN(n1147) );
  XNOR2_X1 U1798 ( .A(n1345), .B(n1538), .ZN(n1044) );
  XNOR2_X1 U1799 ( .A(n1560), .B(n1538), .ZN(n1031) );
  XNOR2_X1 U1800 ( .A(n1546), .B(n1538), .ZN(n1046) );
  XNOR2_X1 U1801 ( .A(n1564), .B(n1335), .ZN(n1027) );
  XNOR2_X1 U1802 ( .A(n1553), .B(n1538), .ZN(n1038) );
  XNOR2_X1 U1803 ( .A(n1346), .B(n1538), .ZN(n1045) );
  XNOR2_X1 U1804 ( .A(n1551), .B(n1538), .ZN(n1040) );
  XNOR2_X1 U1805 ( .A(n1552), .B(n1538), .ZN(n1039) );
  XNOR2_X1 U1806 ( .A(n1563), .B(n1335), .ZN(n1028) );
  XNOR2_X1 U1807 ( .A(n1554), .B(n1538), .ZN(n1037) );
  XNOR2_X1 U1808 ( .A(n1561), .B(n1335), .ZN(n1030) );
  XNOR2_X1 U1809 ( .A(n1092), .B(n1335), .ZN(n1029) );
  XNOR2_X1 U1810 ( .A(n1325), .B(n1538), .ZN(n1043) );
  XNOR2_X1 U1811 ( .A(n1352), .B(n1538), .ZN(n1042) );
  XNOR2_X1 U1812 ( .A(n1343), .B(n1538), .ZN(n1041) );
  XNOR2_X1 U1813 ( .A(n1558), .B(n1335), .ZN(n1033) );
  XNOR2_X1 U1814 ( .A(n1555), .B(n1538), .ZN(n1036) );
  XNOR2_X1 U1815 ( .A(n1559), .B(n1335), .ZN(n1032) );
  XNOR2_X1 U1816 ( .A(n1556), .B(n1538), .ZN(n1035) );
  XNOR2_X1 U1817 ( .A(n1557), .B(n1538), .ZN(n1034) );
  NAND2_X1 U1818 ( .A1(n1523), .A2(n200), .ZN(n81) );
  NAND2_X1 U1819 ( .A1(n202), .A2(n1523), .ZN(n195) );
  XNOR2_X1 U1820 ( .A(n1564), .B(n1334), .ZN(n985) );
  XNOR2_X1 U1821 ( .A(n1563), .B(n1334), .ZN(n986) );
  XNOR2_X1 U1822 ( .A(n1560), .B(n1334), .ZN(n989) );
  XNOR2_X1 U1823 ( .A(n1561), .B(n1334), .ZN(n988) );
  XNOR2_X1 U1824 ( .A(n1355), .B(n1334), .ZN(n987) );
  XNOR2_X1 U1825 ( .A(n1558), .B(n1334), .ZN(n991) );
  XNOR2_X1 U1826 ( .A(n1559), .B(n1334), .ZN(n990) );
  XNOR2_X1 U1827 ( .A(n1546), .B(n1334), .ZN(n1004) );
  INV_X1 U1828 ( .A(n1334), .ZN(n1145) );
  XNOR2_X1 U1829 ( .A(n1347), .B(n1334), .ZN(n1003) );
  XNOR2_X1 U1830 ( .A(n1554), .B(n1540), .ZN(n995) );
  XNOR2_X1 U1831 ( .A(n1557), .B(n1334), .ZN(n992) );
  XNOR2_X1 U1832 ( .A(n1540), .B(n1556), .ZN(n993) );
  XNOR2_X1 U1833 ( .A(n1099), .B(n25), .ZN(n994) );
  XNOR2_X1 U1834 ( .A(n1343), .B(n1334), .ZN(n999) );
  XNOR2_X1 U1835 ( .A(n1352), .B(n1334), .ZN(n1000) );
  XNOR2_X1 U1836 ( .A(n1551), .B(n1540), .ZN(n998) );
  XNOR2_X1 U1837 ( .A(n1325), .B(n1540), .ZN(n1001) );
  XNOR2_X1 U1838 ( .A(n1548), .B(n1540), .ZN(n1002) );
  XNOR2_X1 U1839 ( .A(n1552), .B(n1540), .ZN(n997) );
  XNOR2_X1 U1840 ( .A(n1553), .B(n1334), .ZN(n996) );
  XOR2_X1 U1841 ( .A(n25), .B(a[8]), .Z(n1115) );
  INV_X1 U1842 ( .A(n204), .ZN(n284) );
  NOR2_X1 U1843 ( .A1(n204), .A2(n209), .ZN(n202) );
  OAI21_X1 U1844 ( .B1(n204), .B2(n210), .A(n205), .ZN(n203) );
  NOR2_X2 U1845 ( .A1(n557), .A2(n568), .ZN(n204) );
  XOR2_X1 U1846 ( .A(n242), .B(n89), .Z(product[7]) );
  OAI21_X1 U1847 ( .B1(n242), .B2(n240), .A(n241), .ZN(n239) );
  NAND2_X1 U1848 ( .A1(n633), .A2(n636), .ZN(n249) );
  NOR2_X1 U1849 ( .A1(n140), .A2(n1267), .ZN(n133) );
  OAI21_X1 U1850 ( .B1(n141), .B2(n135), .A(n136), .ZN(n134) );
  NAND2_X1 U1851 ( .A1(n371), .A2(n382), .ZN(n136) );
  INV_X1 U1852 ( .A(n1278), .ZN(n211) );
  INV_X1 U1853 ( .A(n1270), .ZN(n220) );
  AOI21_X1 U1854 ( .B1(n221), .B2(n213), .A(n214), .ZN(n212) );
  AOI21_X1 U1855 ( .B1(n203), .B2(n1523), .A(n1526), .ZN(n196) );
  XNOR2_X1 U1856 ( .A(n1553), .B(n1447), .ZN(n1080) );
  XNOR2_X1 U1857 ( .A(n1552), .B(n1316), .ZN(n1081) );
  XNOR2_X1 U1858 ( .A(n1561), .B(n1447), .ZN(n1072) );
  XNOR2_X1 U1859 ( .A(n1560), .B(n1447), .ZN(n1073) );
  XNOR2_X1 U1860 ( .A(n1562), .B(n1315), .ZN(n1071) );
  XNOR2_X1 U1861 ( .A(n1563), .B(n1447), .ZN(n1070) );
  XNOR2_X1 U1862 ( .A(n1558), .B(n1316), .ZN(n1075) );
  XNOR2_X1 U1863 ( .A(n1337), .B(n1447), .ZN(n1079) );
  XNOR2_X1 U1864 ( .A(n1559), .B(n1316), .ZN(n1074) );
  XNOR2_X1 U1865 ( .A(n1555), .B(n1317), .ZN(n1078) );
  XNOR2_X1 U1866 ( .A(n1557), .B(n1317), .ZN(n1076) );
  XNOR2_X1 U1867 ( .A(n1556), .B(n1447), .ZN(n1077) );
  XNOR2_X1 U1868 ( .A(n1551), .B(n1317), .ZN(n1082) );
  XNOR2_X1 U1869 ( .A(n1550), .B(n1447), .ZN(n1083) );
  XNOR2_X1 U1870 ( .A(n1353), .B(n1316), .ZN(n1084) );
  XNOR2_X1 U1871 ( .A(n1326), .B(n1447), .ZN(n1085) );
  XNOR2_X1 U1872 ( .A(n1564), .B(n1447), .ZN(n1069) );
  XNOR2_X1 U1873 ( .A(n1546), .B(n1447), .ZN(n1088) );
  XNOR2_X1 U1874 ( .A(n1345), .B(n1317), .ZN(n1086) );
  INV_X1 U1875 ( .A(n1447), .ZN(n1149) );
  XNOR2_X1 U1876 ( .A(n1347), .B(n1316), .ZN(n1087) );
  AOI21_X1 U1877 ( .B1(n146), .B2(n133), .A(n134), .ZN(n132) );
  NAND2_X1 U1878 ( .A1(n145), .A2(n133), .ZN(n131) );
  NAND2_X1 U1879 ( .A1(n1233), .A2(n1520), .ZN(n180) );
  NAND2_X1 U1880 ( .A1(n1520), .A2(n185), .ZN(n79) );
  AOI21_X1 U1881 ( .B1(n1520), .B2(n1524), .A(n1528), .ZN(n181) );
  INV_X1 U1882 ( .A(n1527), .ZN(n274) );
  OAI21_X1 U1883 ( .B1(n147), .B2(n151), .A(n148), .ZN(n146) );
  NAND2_X1 U1884 ( .A1(n397), .A2(n410), .ZN(n148) );
  OAI21_X1 U1885 ( .B1(n193), .B2(n1259), .A(n188), .ZN(n186) );
  AOI21_X1 U1886 ( .B1(n165), .B2(n156), .A(n157), .ZN(n155) );
  OAI21_X1 U1887 ( .B1(n166), .B2(n172), .A(n167), .ZN(n165) );
  OAI21_X1 U1888 ( .B1(n158), .B2(n162), .A(n159), .ZN(n157) );
  NAND2_X1 U1889 ( .A1(n443), .A2(n460), .ZN(n162) );
  NOR2_X1 U1890 ( .A1(n427), .A2(n442), .ZN(n158) );
  OAI21_X1 U1891 ( .B1(n152), .B2(n1273), .A(n1464), .ZN(n149) );
  INV_X1 U1892 ( .A(n150), .ZN(n275) );
  NOR2_X1 U1893 ( .A1(n150), .A2(n1527), .ZN(n145) );
  INV_X1 U1894 ( .A(n161), .ZN(n277) );
  OAI21_X1 U1895 ( .B1(n163), .B2(n161), .A(n162), .ZN(n160) );
  NOR2_X1 U1896 ( .A1(n161), .A2(n1493), .ZN(n156) );
  OAI21_X1 U1897 ( .B1(n193), .B2(n180), .A(n1341), .ZN(n179) );
  OAI21_X1 U1898 ( .B1(n181), .B2(n177), .A(n178), .ZN(n176) );
  OAI22_X1 U1899 ( .A1(n1472), .A2(n1024), .B1(n1023), .B2(n1517), .ZN(n817)
         );
  OAI22_X1 U1900 ( .A1(n1472), .A2(n1014), .B1(n1013), .B2(n1517), .ZN(n807)
         );
  OAI22_X1 U1901 ( .A1(n1472), .A2(n1146), .B1(n1026), .B2(n1517), .ZN(n676)
         );
  OAI22_X1 U1902 ( .A1(n1472), .A2(n1007), .B1(n1006), .B2(n1517), .ZN(n394)
         );
  OAI22_X1 U1903 ( .A1(n1472), .A2(n1021), .B1(n1020), .B2(n1517), .ZN(n814)
         );
  OAI22_X1 U1904 ( .A1(n1006), .A2(n1472), .B1(n1006), .B2(n1517), .ZN(n658)
         );
  OAI22_X1 U1905 ( .A1(n1472), .A2(n1025), .B1(n1024), .B2(n1517), .ZN(n818)
         );
  OAI22_X1 U1906 ( .A1(n1472), .A2(n1012), .B1(n1011), .B2(n1517), .ZN(n805)
         );
  OAI22_X1 U1907 ( .A1(n1472), .A2(n1008), .B1(n1007), .B2(n1517), .ZN(n801)
         );
  OAI22_X1 U1908 ( .A1(n1472), .A2(n1009), .B1(n1008), .B2(n1517), .ZN(n802)
         );
  OAI22_X1 U1909 ( .A1(n1015), .A2(n1472), .B1(n1014), .B2(n1517), .ZN(n808)
         );
  OAI22_X1 U1910 ( .A1(n1472), .A2(n1023), .B1(n1022), .B2(n1517), .ZN(n816)
         );
  OAI22_X1 U1911 ( .A1(n1472), .A2(n1010), .B1(n1009), .B2(n1517), .ZN(n803)
         );
  OAI22_X1 U1912 ( .A1(n1472), .A2(n1020), .B1(n1019), .B2(n1517), .ZN(n813)
         );
  OAI22_X1 U1913 ( .A1(n1472), .A2(n1019), .B1(n1018), .B2(n1517), .ZN(n812)
         );
  OAI22_X1 U1914 ( .A1(n1472), .A2(n1013), .B1(n1012), .B2(n1517), .ZN(n806)
         );
  OAI22_X1 U1915 ( .A1(n1472), .A2(n1018), .B1(n1017), .B2(n1517), .ZN(n811)
         );
  OAI22_X1 U1916 ( .A1(n1472), .A2(n1022), .B1(n1021), .B2(n1517), .ZN(n815)
         );
  OAI22_X1 U1917 ( .A1(n1472), .A2(n1011), .B1(n1010), .B2(n1517), .ZN(n804)
         );
  OAI22_X1 U1918 ( .A1(n1472), .A2(n1017), .B1(n1016), .B2(n1517), .ZN(n810)
         );
  INV_X1 U1919 ( .A(n1517), .ZN(n659) );
  OAI22_X1 U1920 ( .A1(n1472), .A2(n1016), .B1(n1015), .B2(n1517), .ZN(n809)
         );
  NAND2_X1 U1921 ( .A1(n637), .A2(n638), .ZN(n254) );
  OAI21_X1 U1922 ( .B1(n222), .B2(n234), .A(n223), .ZN(n221) );
  OAI21_X1 U1923 ( .B1(n195), .B2(n212), .A(n196), .ZN(n194) );
  OAI21_X1 U1924 ( .B1(n152), .B2(n131), .A(n1444), .ZN(n130) );
  OAI22_X1 U1925 ( .A1(n901), .A2(n1466), .B1(n901), .B2(n1463), .ZN(n643) );
  OAI22_X1 U1926 ( .A1(n1466), .A2(n902), .B1(n901), .B2(n1463), .ZN(n304) );
  OAI22_X1 U1927 ( .A1(n1466), .A2(n903), .B1(n902), .B2(n1463), .ZN(n701) );
  OAI21_X1 U1928 ( .B1(n132), .B2(n128), .A(n129), .ZN(n127) );
  OAI22_X1 U1929 ( .A1(n1466), .A2(n905), .B1(n904), .B2(n1463), .ZN(n703) );
  OAI22_X1 U1930 ( .A1(n1466), .A2(n904), .B1(n903), .B2(n1463), .ZN(n702) );
  OAI22_X1 U1931 ( .A1(n1466), .A2(n906), .B1(n905), .B2(n1463), .ZN(n704) );
  OAI22_X1 U1932 ( .A1(n1466), .A2(n907), .B1(n906), .B2(n1463), .ZN(n705) );
  OAI22_X1 U1933 ( .A1(n1466), .A2(n908), .B1(n907), .B2(n1463), .ZN(n706) );
  OAI22_X1 U1934 ( .A1(n54), .A2(n909), .B1(n908), .B2(n1511), .ZN(n707) );
  OAI22_X1 U1935 ( .A1(n54), .A2(n910), .B1(n909), .B2(n1511), .ZN(n708) );
  OAI22_X1 U1936 ( .A1(n54), .A2(n911), .B1(n910), .B2(n1511), .ZN(n709) );
  OAI22_X1 U1937 ( .A1(n54), .A2(n1141), .B1(n921), .B2(n1511), .ZN(n671) );
  OAI22_X1 U1938 ( .A1(n54), .A2(n915), .B1(n914), .B2(n1511), .ZN(n713) );
  OAI22_X1 U1939 ( .A1(n54), .A2(n912), .B1(n911), .B2(n1511), .ZN(n710) );
  OAI22_X1 U1940 ( .A1(n54), .A2(n913), .B1(n912), .B2(n1511), .ZN(n711) );
  OAI22_X1 U1941 ( .A1(n54), .A2(n914), .B1(n913), .B2(n1511), .ZN(n712) );
  OAI22_X1 U1942 ( .A1(n54), .A2(n918), .B1(n917), .B2(n1511), .ZN(n716) );
  OAI22_X1 U1943 ( .A1(n54), .A2(n920), .B1(n919), .B2(n1511), .ZN(n718) );
  OAI22_X1 U1944 ( .A1(n54), .A2(n917), .B1(n916), .B2(n1511), .ZN(n715) );
  OAI22_X1 U1945 ( .A1(n54), .A2(n916), .B1(n915), .B2(n1511), .ZN(n714) );
  INV_X1 U1946 ( .A(n1511), .ZN(n644) );
  INV_X1 U1947 ( .A(n1525), .ZN(n278) );
  OAI22_X1 U1948 ( .A1(n922), .A2(n1469), .B1(n922), .B2(n1375), .ZN(n646) );
  NOR2_X1 U1949 ( .A1(n1525), .A2(n171), .ZN(n164) );
  OAI22_X1 U1950 ( .A1(n1469), .A2(n924), .B1(n923), .B2(n1375), .ZN(n721) );
  OAI22_X1 U1951 ( .A1(n1469), .A2(n923), .B1(n922), .B2(n1375), .ZN(n314) );
  OAI22_X1 U1952 ( .A1(n1469), .A2(n925), .B1(n924), .B2(n1519), .ZN(n722) );
  OAI22_X1 U1953 ( .A1(n1469), .A2(n927), .B1(n926), .B2(n1375), .ZN(n724) );
  OAI22_X1 U1954 ( .A1(n1469), .A2(n926), .B1(n925), .B2(n1519), .ZN(n723) );
  OAI22_X1 U1955 ( .A1(n1469), .A2(n928), .B1(n927), .B2(n1375), .ZN(n725) );
  OAI22_X1 U1956 ( .A1(n1469), .A2(n929), .B1(n928), .B2(n1519), .ZN(n726) );
  OAI22_X1 U1957 ( .A1(n1469), .A2(n930), .B1(n929), .B2(n1375), .ZN(n727) );
  OAI22_X1 U1958 ( .A1(n1470), .A2(n1246), .B1(n930), .B2(n1375), .ZN(n728) );
  OAI22_X1 U1959 ( .A1(n1469), .A2(n933), .B1(n932), .B2(n1519), .ZN(n730) );
  OAI22_X1 U1960 ( .A1(n1470), .A2(n934), .B1(n933), .B2(n1519), .ZN(n731) );
  OAI22_X1 U1961 ( .A1(n48), .A2(n1142), .B1(n942), .B2(n1518), .ZN(n672) );
  OAI22_X1 U1962 ( .A1(n1469), .A2(n941), .B1(n940), .B2(n1519), .ZN(n738) );
  OAI22_X1 U1963 ( .A1(n1470), .A2(n932), .B1(n931), .B2(n1518), .ZN(n729) );
  OAI22_X1 U1964 ( .A1(n1470), .A2(n936), .B1(n935), .B2(n1518), .ZN(n733) );
  OAI22_X1 U1965 ( .A1(n1470), .A2(n939), .B1(n938), .B2(n1518), .ZN(n736) );
  OAI22_X1 U1966 ( .A1(n48), .A2(n937), .B1(n936), .B2(n1518), .ZN(n734) );
  OAI22_X1 U1967 ( .A1(n1470), .A2(n940), .B1(n939), .B2(n1518), .ZN(n737) );
  OAI22_X1 U1968 ( .A1(n935), .A2(n1470), .B1(n934), .B2(n1518), .ZN(n732) );
  OAI22_X1 U1969 ( .A1(n48), .A2(n938), .B1(n937), .B2(n1519), .ZN(n735) );
  OAI22_X1 U1970 ( .A1(n880), .A2(n1441), .B1(n880), .B2(n1338), .ZN(n640) );
  OAI22_X1 U1971 ( .A1(n1442), .A2(n881), .B1(n880), .B2(n1338), .ZN(n298) );
  OAI22_X1 U1972 ( .A1(n1441), .A2(n882), .B1(n881), .B2(n1338), .ZN(n681) );
  OAI22_X1 U1973 ( .A1(n1442), .A2(n883), .B1(n882), .B2(n1338), .ZN(n682) );
  OAI22_X1 U1974 ( .A1(n1441), .A2(n884), .B1(n883), .B2(n1338), .ZN(n683) );
  OAI22_X1 U1975 ( .A1(n1441), .A2(n886), .B1(n885), .B2(n1338), .ZN(n685) );
  OAI22_X1 U1976 ( .A1(n1442), .A2(n885), .B1(n884), .B2(n1338), .ZN(n684) );
  OAI22_X1 U1977 ( .A1(n1442), .A2(n887), .B1(n886), .B2(n1338), .ZN(n686) );
  OAI22_X1 U1978 ( .A1(n1441), .A2(n888), .B1(n887), .B2(n1338), .ZN(n687) );
  OAI22_X1 U1979 ( .A1(n1442), .A2(n889), .B1(n888), .B2(n1338), .ZN(n688) );
  OAI22_X1 U1980 ( .A1(n1441), .A2(n890), .B1(n889), .B2(n1338), .ZN(n689) );
  OAI22_X1 U1981 ( .A1(n1442), .A2(n891), .B1(n890), .B2(n1486), .ZN(n690) );
  OAI22_X1 U1982 ( .A1(n1441), .A2(n892), .B1(n891), .B2(n1486), .ZN(n691) );
  OAI22_X1 U1983 ( .A1(n1441), .A2(n894), .B1(n893), .B2(n1486), .ZN(n693) );
  OAI22_X1 U1984 ( .A1(n1442), .A2(n893), .B1(n892), .B2(n1486), .ZN(n692) );
  OAI22_X1 U1985 ( .A1(n1441), .A2(n899), .B1(n898), .B2(n1486), .ZN(n698) );
  OAI22_X1 U1986 ( .A1(n1442), .A2(n895), .B1(n894), .B2(n1486), .ZN(n694) );
  OAI22_X1 U1987 ( .A1(n60), .A2(n1140), .B1(n900), .B2(n1486), .ZN(n670) );
  OAI22_X1 U1988 ( .A1(n60), .A2(n898), .B1(n897), .B2(n1486), .ZN(n697) );
  OAI22_X1 U1989 ( .A1(n60), .A2(n896), .B1(n895), .B2(n1486), .ZN(n695) );
  OAI22_X1 U1990 ( .A1(n60), .A2(n897), .B1(n896), .B2(n1486), .ZN(n696) );
  INV_X1 U1991 ( .A(n194), .ZN(n193) );
  INV_X1 U1992 ( .A(n1482), .ZN(n152) );
  AOI21_X1 U1993 ( .B1(n1482), .B2(n1327), .A(n1416), .ZN(n125) );
  AOI21_X1 U1994 ( .B1(n194), .B2(n175), .A(n176), .ZN(n174) );
  OAI22_X1 U1995 ( .A1(n1481), .A2(n965), .B1(n964), .B2(n1512), .ZN(n346) );
  OAI22_X1 U1996 ( .A1(n964), .A2(n1480), .B1(n964), .B2(n1513), .ZN(n652) );
  OAI22_X1 U1997 ( .A1(n1480), .A2(n966), .B1(n965), .B2(n1512), .ZN(n761) );
  OAI22_X1 U1998 ( .A1(n1481), .A2(n967), .B1(n966), .B2(n1513), .ZN(n762) );
  OAI22_X1 U1999 ( .A1(n1481), .A2(n968), .B1(n967), .B2(n1512), .ZN(n763) );
  OAI22_X1 U2000 ( .A1(n1481), .A2(n973), .B1(n972), .B2(n1513), .ZN(n768) );
  OAI22_X1 U2001 ( .A1(n1480), .A2(n972), .B1(n971), .B2(n1513), .ZN(n767) );
  OAI22_X1 U2002 ( .A1(n1481), .A2(n975), .B1(n974), .B2(n1512), .ZN(n770) );
  OAI22_X1 U2003 ( .A1(n1481), .A2(n969), .B1(n968), .B2(n1512), .ZN(n764) );
  OAI22_X1 U2004 ( .A1(n1479), .A2(n971), .B1(n970), .B2(n1512), .ZN(n766) );
  OAI22_X1 U2005 ( .A1(n1481), .A2(n970), .B1(n969), .B2(n1513), .ZN(n765) );
  OAI22_X1 U2006 ( .A1(n1480), .A2(n977), .B1(n976), .B2(n1512), .ZN(n772) );
  OAI22_X1 U2007 ( .A1(n1480), .A2(n1144), .B1(n984), .B2(n1513), .ZN(n674) );
  OAI22_X1 U2008 ( .A1(n1480), .A2(n983), .B1(n982), .B2(n1512), .ZN(n778) );
  OAI22_X1 U2009 ( .A1(n1480), .A2(n982), .B1(n981), .B2(n1513), .ZN(n777) );
  OAI22_X1 U2010 ( .A1(n1481), .A2(n974), .B1(n973), .B2(n1512), .ZN(n769) );
  OAI22_X1 U2011 ( .A1(n1479), .A2(n976), .B1(n975), .B2(n1512), .ZN(n771) );
  OAI22_X1 U2012 ( .A1(n979), .A2(n1481), .B1(n978), .B2(n1513), .ZN(n774) );
  OAI22_X1 U2013 ( .A1(n1480), .A2(n978), .B1(n977), .B2(n1512), .ZN(n773) );
  OAI22_X1 U2014 ( .A1(n1481), .A2(n980), .B1(n979), .B2(n1512), .ZN(n775) );
  OAI22_X1 U2015 ( .A1(n1481), .A2(n981), .B1(n980), .B2(n1513), .ZN(n776) );
  INV_X1 U2016 ( .A(n1513), .ZN(n653) );
  INV_X1 U2017 ( .A(n1361), .ZN(n173) );
  OAI21_X1 U2018 ( .B1(n174), .B2(n154), .A(n155), .ZN(n153) );
  OAI22_X1 U2019 ( .A1(n985), .A2(n1483), .B1(n985), .B2(n1515), .ZN(n655) );
  OAI22_X1 U2020 ( .A1(n1484), .A2(n986), .B1(n985), .B2(n1241), .ZN(n368) );
  OAI22_X1 U2021 ( .A1(n1247), .A2(n987), .B1(n986), .B2(n1515), .ZN(n781) );
  OAI22_X1 U2022 ( .A1(n1269), .A2(n989), .B1(n988), .B2(n1241), .ZN(n783) );
  OAI22_X1 U2023 ( .A1(n1484), .A2(n992), .B1(n991), .B2(n1515), .ZN(n786) );
  OAI22_X1 U2024 ( .A1(n1483), .A2(n990), .B1(n989), .B2(n1241), .ZN(n784) );
  OAI22_X1 U2025 ( .A1(n1483), .A2(n1003), .B1(n1002), .B2(n1241), .ZN(n797)
         );
  OAI22_X1 U2026 ( .A1(n1269), .A2(n988), .B1(n987), .B2(n1515), .ZN(n782) );
  OAI22_X1 U2027 ( .A1(n1417), .A2(n991), .B1(n990), .B2(n1515), .ZN(n785) );
  OAI22_X1 U2028 ( .A1(n1483), .A2(n996), .B1(n995), .B2(n1515), .ZN(n790) );
  OAI22_X1 U2029 ( .A1(n1484), .A2(n993), .B1(n992), .B2(n1241), .ZN(n787) );
  OAI22_X1 U2030 ( .A1(n1484), .A2(n994), .B1(n993), .B2(n1241), .ZN(n788) );
  OAI22_X1 U2031 ( .A1(n1247), .A2(n999), .B1(n998), .B2(n1241), .ZN(n793) );
  OAI22_X1 U2032 ( .A1(n1417), .A2(n995), .B1(n994), .B2(n1514), .ZN(n789) );
  OAI22_X1 U2033 ( .A1(n1483), .A2(n1000), .B1(n999), .B2(n1515), .ZN(n794) );
  OAI22_X1 U2034 ( .A1(n1484), .A2(n1004), .B1(n1003), .B2(n1515), .ZN(n798)
         );
  OAI22_X1 U2035 ( .A1(n1483), .A2(n1002), .B1(n1001), .B2(n1241), .ZN(n796)
         );
  OAI22_X1 U2036 ( .A1(n1247), .A2(n1145), .B1(n1005), .B2(n1241), .ZN(n675)
         );
  OAI22_X1 U2037 ( .A1(n1269), .A2(n998), .B1(n997), .B2(n1241), .ZN(n792) );
  INV_X1 U2038 ( .A(n1241), .ZN(n656) );
  OAI22_X1 U2039 ( .A1(n1484), .A2(n1001), .B1(n1000), .B2(n1241), .ZN(n795)
         );
  OAI22_X1 U2040 ( .A1(n1483), .A2(n997), .B1(n996), .B2(n1515), .ZN(n791) );
  INV_X1 U2041 ( .A(n101), .ZN(n264) );
  OAI22_X1 U2042 ( .A1(n943), .A2(n1271), .B1(n943), .B2(n1349), .ZN(n649) );
  OAI22_X1 U2043 ( .A1(n1503), .A2(n944), .B1(n943), .B2(n1349), .ZN(n328) );
  OAI22_X1 U2044 ( .A1(n1271), .A2(n945), .B1(n944), .B2(n1349), .ZN(n741) );
  OAI22_X1 U2045 ( .A1(n1503), .A2(n947), .B1(n946), .B2(n1349), .ZN(n743) );
  OAI22_X1 U2046 ( .A1(n1271), .A2(n946), .B1(n945), .B2(n1349), .ZN(n742) );
  OAI22_X1 U2047 ( .A1(n1503), .A2(n948), .B1(n947), .B2(n1349), .ZN(n744) );
  OAI22_X1 U2048 ( .A1(n1503), .A2(n949), .B1(n948), .B2(n1507), .ZN(n745) );
  OAI22_X1 U2049 ( .A1(n1503), .A2(n952), .B1(n951), .B2(n1507), .ZN(n748) );
  OAI22_X1 U2050 ( .A1(n1503), .A2(n957), .B1(n956), .B2(n1507), .ZN(n753) );
  OAI22_X1 U2051 ( .A1(n951), .A2(n1504), .B1(n950), .B2(n1507), .ZN(n747) );
  OAI22_X1 U2052 ( .A1(n1504), .A2(n950), .B1(n949), .B2(n1507), .ZN(n746) );
  OAI22_X1 U2053 ( .A1(n1504), .A2(n953), .B1(n952), .B2(n1507), .ZN(n749) );
  OAI22_X1 U2054 ( .A1(n1503), .A2(n956), .B1(n955), .B2(n1507), .ZN(n752) );
  OAI22_X1 U2055 ( .A1(n1503), .A2(n958), .B1(n957), .B2(n1507), .ZN(n754) );
  OAI22_X1 U2056 ( .A1(n1504), .A2(n955), .B1(n954), .B2(n1507), .ZN(n751) );
  OAI22_X1 U2057 ( .A1(n1503), .A2(n1143), .B1(n963), .B2(n1507), .ZN(n673) );
  OAI22_X1 U2058 ( .A1(n1504), .A2(n954), .B1(n953), .B2(n1507), .ZN(n750) );
  OAI22_X1 U2059 ( .A1(n1503), .A2(n961), .B1(n960), .B2(n1507), .ZN(n757) );
  OAI22_X1 U2060 ( .A1(n1503), .A2(n960), .B1(n959), .B2(n1507), .ZN(n756) );
  OAI22_X1 U2061 ( .A1(n1504), .A2(n962), .B1(n961), .B2(n1507), .ZN(n758) );
  OAI22_X1 U2062 ( .A1(n1503), .A2(n959), .B1(n958), .B2(n1507), .ZN(n755) );
  BUF_X4 U2063 ( .A(n31), .Z(n1541) );
  OAI21_X1 U2064 ( .B1(n1485), .B2(n123), .A(n124), .ZN(n122) );
  XNOR2_X1 U2065 ( .A(n1473), .B(n67), .ZN(product[29]) );
  XNOR2_X1 U2066 ( .A(n1378), .B(n65), .ZN(product[31]) );
  AOI21_X1 U2067 ( .B1(n1378), .B2(n1498), .A(n111), .ZN(n109) );
  OAI22_X1 U2068 ( .A1(n1475), .A2(n1039), .B1(n1038), .B2(n1302), .ZN(n831)
         );
  OAI22_X1 U2069 ( .A1(n1475), .A2(n1031), .B1(n1030), .B2(n1516), .ZN(n823)
         );
  OAI22_X1 U2070 ( .A1(n1475), .A2(n1240), .B1(n1031), .B2(n1516), .ZN(n824)
         );
  OAI22_X1 U2071 ( .A1(n1260), .A2(n1041), .B1(n1040), .B2(n1516), .ZN(n833)
         );
  OAI22_X1 U2072 ( .A1(n1475), .A2(n1034), .B1(n1033), .B2(n1516), .ZN(n826)
         );
  OAI22_X1 U2073 ( .A1(n1475), .A2(n1045), .B1(n1044), .B2(n1302), .ZN(n837)
         );
  OAI22_X1 U2074 ( .A1(n1475), .A2(n1028), .B1(n1027), .B2(n1516), .ZN(n424)
         );
  OAI22_X1 U2075 ( .A1(n1027), .A2(n1475), .B1(n1027), .B2(n1516), .ZN(n661)
         );
  OAI22_X1 U2076 ( .A1(n1260), .A2(n1038), .B1(n1037), .B2(n1516), .ZN(n830)
         );
  OAI22_X1 U2077 ( .A1(n1260), .A2(n1044), .B1(n1043), .B2(n1516), .ZN(n836)
         );
  OAI22_X1 U2078 ( .A1(n1474), .A2(n1030), .B1(n1029), .B2(n1516), .ZN(n822)
         );
  OAI22_X1 U2079 ( .A1(n1029), .A2(n1474), .B1(n1516), .B2(n1028), .ZN(n821)
         );
  OAI22_X1 U2080 ( .A1(n1474), .A2(n1033), .B1(n1032), .B2(n1516), .ZN(n825)
         );
  OAI22_X1 U2081 ( .A1(n1260), .A2(n1040), .B1(n1039), .B2(n1516), .ZN(n832)
         );
  OAI22_X1 U2082 ( .A1(n1475), .A2(n1037), .B1(n1036), .B2(n1516), .ZN(n829)
         );
  OAI22_X1 U2083 ( .A1(n1260), .A2(n1147), .B1(n1047), .B2(n1516), .ZN(n677)
         );
  OAI22_X1 U2084 ( .A1(n1475), .A2(n1036), .B1(n1035), .B2(n1516), .ZN(n828)
         );
  OAI22_X1 U2085 ( .A1(n1260), .A2(n1043), .B1(n1042), .B2(n1516), .ZN(n835)
         );
  OAI22_X1 U2086 ( .A1(n1260), .A2(n1042), .B1(n1041), .B2(n1516), .ZN(n834)
         );
  OAI22_X1 U2087 ( .A1(n1260), .A2(n1035), .B1(n1034), .B2(n1516), .ZN(n827)
         );
  OAI22_X1 U2088 ( .A1(n1260), .A2(n1046), .B1(n1045), .B2(n1516), .ZN(n838)
         );
  INV_X1 U2089 ( .A(n1516), .ZN(n662) );
  XNOR2_X1 U2090 ( .A(n1446), .B(n63), .ZN(product[33]) );
  XOR2_X1 U2091 ( .A(n109), .B(n64), .Z(product[32]) );
  XOR2_X1 U2092 ( .A(n117), .B(n66), .Z(product[30]) );
  XOR2_X1 U2093 ( .A(n125), .B(n68), .Z(product[28]) );
  AOI21_X1 U2094 ( .B1(n106), .B2(n1499), .A(n103), .ZN(n101) );
  OAI21_X1 U2095 ( .B1(n1471), .B2(n107), .A(n108), .ZN(n106) );
  OAI21_X1 U2096 ( .B1(n1476), .B2(n115), .A(n116), .ZN(n114) );
  OAI22_X1 U2097 ( .A1(n1309), .A2(n1055), .B1(n1054), .B2(n1505), .ZN(n846)
         );
  OAI22_X1 U2098 ( .A1(n1309), .A2(n1051), .B1(n1050), .B2(n1505), .ZN(n842)
         );
  OAI22_X1 U2099 ( .A1(n1477), .A2(n1062), .B1(n1061), .B2(n1506), .ZN(n853)
         );
  OAI22_X1 U2100 ( .A1(n1309), .A2(n1059), .B1(n1058), .B2(n1506), .ZN(n850)
         );
  OAI22_X1 U2101 ( .A1(n1477), .A2(n1060), .B1(n1059), .B2(n1505), .ZN(n851)
         );
  OAI22_X1 U2102 ( .A1(n1477), .A2(n1053), .B1(n1052), .B2(n1505), .ZN(n844)
         );
  OAI22_X1 U2103 ( .A1(n1309), .A2(n1049), .B1(n1332), .B2(n1505), .ZN(n458)
         );
  OAI22_X1 U2104 ( .A1(n1477), .A2(n1052), .B1(n1051), .B2(n1506), .ZN(n843)
         );
  OAI22_X1 U2105 ( .A1(n1477), .A2(n1063), .B1(n1062), .B2(n1506), .ZN(n854)
         );
  OAI22_X1 U2106 ( .A1(n1477), .A2(n1050), .B1(n1049), .B2(n1506), .ZN(n841)
         );
  OAI22_X1 U2107 ( .A1(n1477), .A2(n1057), .B1(n1056), .B2(n1505), .ZN(n848)
         );
  OAI22_X1 U2108 ( .A1(n1309), .A2(n1065), .B1(n1064), .B2(n1505), .ZN(n856)
         );
  OAI22_X1 U2109 ( .A1(n1477), .A2(n1056), .B1(n1055), .B2(n1506), .ZN(n847)
         );
  OAI22_X1 U2110 ( .A1(n1309), .A2(n1058), .B1(n1057), .B2(n1505), .ZN(n849)
         );
  OAI22_X1 U2111 ( .A1(n1309), .A2(n1148), .B1(n1068), .B2(n1505), .ZN(n678)
         );
  OAI22_X1 U2112 ( .A1(n1309), .A2(n1054), .B1(n1053), .B2(n1506), .ZN(n845)
         );
  OAI22_X1 U2113 ( .A1(n1477), .A2(n1061), .B1(n1060), .B2(n1505), .ZN(n852)
         );
  OAI22_X1 U2114 ( .A1(n1332), .A2(n12), .B1(n1048), .B2(n1506), .ZN(n664) );
  OAI22_X1 U2115 ( .A1(n1309), .A2(n1064), .B1(n1063), .B2(n1505), .ZN(n855)
         );
  OAI22_X1 U2116 ( .A1(n1309), .A2(n1067), .B1(n1066), .B2(n1505), .ZN(n858)
         );
  OAI22_X1 U2117 ( .A1(n1477), .A2(n1066), .B1(n1065), .B2(n1506), .ZN(n857)
         );
  INV_X1 U2118 ( .A(n1506), .ZN(n665) );
endmodule


module mac_3_DW01_add_1 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n34, n35, n36, n37, n38, n39, n40, n41, n43, n45, n46, n47,
         n48, n49, n51, n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65,
         n67, n69, n70, n71, n72, n73, n75, n77, n78, n79, n80, n81, n83, n85,
         n86, n87, n88, n89, n91, n93, n94, n95, n96, n97, n99, n101, n102,
         n103, n104, n105, n107, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n119, n121, n122, n124, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n184, n185, n187, n189, n191,
         n193, n195, n197, n199, n201, n203, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405;

  FA_X1 U8 ( .A(B[33]), .B(A[33]), .CI(n40), .CO(n39), .S(SUM[33]) );
  FA_X1 U9 ( .A(B[32]), .B(A[32]), .CI(n185), .CO(n40), .S(SUM[32]) );
  CLKBUF_X1 U254 ( .A(n37), .Z(n344) );
  NAND3_X1 U255 ( .A1(n388), .A2(n387), .A3(n386), .ZN(n345) );
  CLKBUF_X1 U256 ( .A(n46), .Z(n346) );
  OR2_X1 U257 ( .A1(B[0]), .A2(A[0]), .ZN(n347) );
  CLKBUF_X1 U258 ( .A(n363), .Z(n348) );
  CLKBUF_X1 U259 ( .A(n86), .Z(n349) );
  XOR2_X1 U260 ( .A(B[35]), .B(A[35]), .Z(n350) );
  XOR2_X1 U261 ( .A(n38), .B(n350), .Z(SUM[35]) );
  NAND2_X1 U262 ( .A1(n38), .A2(B[35]), .ZN(n351) );
  NAND2_X1 U263 ( .A1(n38), .A2(A[35]), .ZN(n352) );
  NAND2_X1 U264 ( .A1(B[35]), .A2(A[35]), .ZN(n353) );
  NAND3_X1 U265 ( .A1(n351), .A2(n352), .A3(n353), .ZN(n37) );
  CLKBUF_X1 U266 ( .A(n62), .Z(n354) );
  CLKBUF_X1 U267 ( .A(n110), .Z(n355) );
  CLKBUF_X1 U268 ( .A(n150), .Z(n356) );
  AOI21_X1 U269 ( .B1(n355), .B2(n396), .A(n107), .ZN(n357) );
  AOI21_X1 U270 ( .B1(n110), .B2(n396), .A(n107), .ZN(n105) );
  AOI21_X1 U271 ( .B1(n349), .B2(n397), .A(n83), .ZN(n358) );
  AOI21_X1 U272 ( .B1(n86), .B2(n397), .A(n83), .ZN(n81) );
  AOI21_X1 U273 ( .B1(n354), .B2(n402), .A(n59), .ZN(n359) );
  AOI21_X1 U274 ( .B1(n62), .B2(n402), .A(n59), .ZN(n57) );
  AOI21_X1 U275 ( .B1(n130), .B2(n143), .A(n131), .ZN(n360) );
  AOI21_X1 U276 ( .B1(n356), .B2(n114), .A(n115), .ZN(n361) );
  AOI21_X1 U277 ( .B1(n150), .B2(n114), .A(n115), .ZN(n113) );
  CLKBUF_X1 U278 ( .A(n94), .Z(n362) );
  NAND3_X1 U279 ( .A1(n376), .A2(n377), .A3(n378), .ZN(n363) );
  CLKBUF_X1 U280 ( .A(n70), .Z(n364) );
  AOI21_X1 U281 ( .B1(n362), .B2(n400), .A(n91), .ZN(n365) );
  CLKBUF_X1 U282 ( .A(n102), .Z(n366) );
  XOR2_X1 U283 ( .A(B[34]), .B(A[34]), .Z(n367) );
  XOR2_X1 U284 ( .A(n39), .B(n367), .Z(SUM[34]) );
  NAND2_X1 U285 ( .A1(n39), .A2(B[34]), .ZN(n368) );
  NAND2_X1 U286 ( .A1(n39), .A2(A[34]), .ZN(n369) );
  NAND2_X1 U287 ( .A1(B[34]), .A2(A[34]), .ZN(n370) );
  NAND3_X1 U288 ( .A1(n368), .A2(n369), .A3(n370), .ZN(n38) );
  AOI21_X1 U289 ( .B1(n366), .B2(n398), .A(n99), .ZN(n371) );
  NOR2_X2 U290 ( .A1(B[5]), .A2(A[5]), .ZN(n163) );
  NOR2_X2 U291 ( .A1(B[7]), .A2(A[7]), .ZN(n155) );
  NOR2_X1 U292 ( .A1(B[3]), .A2(A[3]), .ZN(n372) );
  NOR2_X1 U293 ( .A1(B[3]), .A2(A[3]), .ZN(n174) );
  NOR2_X1 U294 ( .A1(B[9]), .A2(A[9]), .ZN(n373) );
  NOR2_X1 U295 ( .A1(B[9]), .A2(A[9]), .ZN(n144) );
  NOR2_X1 U296 ( .A1(B[11]), .A2(A[11]), .ZN(n374) );
  NOR2_X1 U297 ( .A1(B[11]), .A2(A[11]), .ZN(n132) );
  XOR2_X1 U298 ( .A(B[36]), .B(A[36]), .Z(n375) );
  XOR2_X1 U299 ( .A(n344), .B(n375), .Z(SUM[36]) );
  NAND2_X1 U300 ( .A1(n37), .A2(B[36]), .ZN(n376) );
  NAND2_X1 U301 ( .A1(n37), .A2(A[36]), .ZN(n377) );
  NAND2_X1 U302 ( .A1(B[36]), .A2(A[36]), .ZN(n378) );
  NAND3_X1 U303 ( .A1(n376), .A2(n377), .A3(n378), .ZN(n36) );
  CLKBUF_X1 U304 ( .A(n54), .Z(n379) );
  CLKBUF_X1 U305 ( .A(n78), .Z(n380) );
  AOI21_X1 U306 ( .B1(n364), .B2(n401), .A(n67), .ZN(n381) );
  AOI21_X1 U307 ( .B1(n70), .B2(n401), .A(n67), .ZN(n65) );
  NAND3_X1 U308 ( .A1(n387), .A2(n386), .A3(n388), .ZN(n382) );
  AOI21_X1 U309 ( .B1(n379), .B2(n403), .A(n51), .ZN(n383) );
  AOI21_X1 U310 ( .B1(n380), .B2(n399), .A(n75), .ZN(n384) );
  XOR2_X1 U311 ( .A(B[37]), .B(A[37]), .Z(n385) );
  XOR2_X1 U312 ( .A(n385), .B(n348), .Z(SUM[37]) );
  NAND2_X1 U313 ( .A1(B[37]), .A2(A[37]), .ZN(n386) );
  NAND2_X1 U314 ( .A1(B[37]), .A2(n36), .ZN(n387) );
  NAND2_X1 U315 ( .A1(A[37]), .A2(n363), .ZN(n388) );
  NAND3_X1 U316 ( .A1(n388), .A2(n387), .A3(n386), .ZN(n35) );
  XOR2_X1 U317 ( .A(B[38]), .B(A[38]), .Z(n389) );
  XOR2_X1 U318 ( .A(n389), .B(n382), .Z(SUM[38]) );
  NAND2_X1 U319 ( .A1(B[38]), .A2(A[38]), .ZN(n390) );
  NAND2_X1 U320 ( .A1(n345), .A2(B[38]), .ZN(n391) );
  NAND2_X1 U321 ( .A1(n35), .A2(A[38]), .ZN(n392) );
  NAND3_X1 U322 ( .A1(n390), .A2(n391), .A3(n392), .ZN(n34) );
  OR2_X1 U323 ( .A1(B[13]), .A2(A[13]), .ZN(n395) );
  OR2_X1 U324 ( .A1(B[12]), .A2(A[12]), .ZN(n394) );
  OR2_X1 U325 ( .A1(B[15]), .A2(A[15]), .ZN(n396) );
  INV_X1 U326 ( .A(n356), .ZN(n149) );
  OAI21_X1 U327 ( .B1(n149), .B2(n128), .A(n360), .ZN(n127) );
  OAI21_X1 U328 ( .B1(n149), .B2(n140), .A(n141), .ZN(n139) );
  INV_X1 U329 ( .A(n143), .ZN(n141) );
  INV_X1 U330 ( .A(n142), .ZN(n140) );
  NAND2_X1 U331 ( .A1(n142), .A2(n130), .ZN(n128) );
  AOI21_X1 U332 ( .B1(n170), .B2(n161), .A(n162), .ZN(n160) );
  INV_X1 U333 ( .A(n171), .ZN(n170) );
  INV_X1 U334 ( .A(n180), .ZN(n179) );
  INV_X1 U335 ( .A(n61), .ZN(n59) );
  INV_X1 U336 ( .A(n93), .ZN(n91) );
  INV_X1 U337 ( .A(n53), .ZN(n51) );
  AOI21_X1 U338 ( .B1(n130), .B2(n143), .A(n131), .ZN(n129) );
  INV_X1 U339 ( .A(n109), .ZN(n107) );
  AOI21_X1 U340 ( .B1(n102), .B2(n398), .A(n99), .ZN(n97) );
  INV_X1 U341 ( .A(n101), .ZN(n99) );
  NOR2_X1 U342 ( .A1(n128), .A2(n116), .ZN(n114) );
  OAI21_X1 U343 ( .B1(n129), .B2(n116), .A(n117), .ZN(n115) );
  NAND2_X1 U344 ( .A1(n394), .A2(n395), .ZN(n116) );
  OAI21_X1 U345 ( .B1(n163), .B2(n169), .A(n164), .ZN(n162) );
  AOI21_X1 U346 ( .B1(n172), .B2(n180), .A(n173), .ZN(n171) );
  NOR2_X1 U347 ( .A1(n177), .A2(n372), .ZN(n172) );
  OAI21_X1 U348 ( .B1(n174), .B2(n178), .A(n175), .ZN(n173) );
  OAI21_X1 U349 ( .B1(n113), .B2(n111), .A(n112), .ZN(n110) );
  INV_X1 U350 ( .A(n85), .ZN(n83) );
  AOI21_X1 U351 ( .B1(n78), .B2(n399), .A(n75), .ZN(n73) );
  INV_X1 U352 ( .A(n77), .ZN(n75) );
  INV_X1 U353 ( .A(n69), .ZN(n67) );
  NOR2_X1 U354 ( .A1(n168), .A2(n163), .ZN(n161) );
  OAI21_X1 U355 ( .B1(n181), .B2(n184), .A(n182), .ZN(n180) );
  AOI21_X1 U356 ( .B1(n395), .B2(n124), .A(n119), .ZN(n117) );
  INV_X1 U357 ( .A(n121), .ZN(n119) );
  NAND2_X1 U358 ( .A1(n195), .A2(n80), .ZN(n11) );
  INV_X1 U359 ( .A(n79), .ZN(n195) );
  NAND2_X1 U360 ( .A1(n197), .A2(n88), .ZN(n13) );
  INV_X1 U361 ( .A(n87), .ZN(n197) );
  OAI21_X1 U362 ( .B1(n171), .B2(n151), .A(n152), .ZN(n150) );
  NAND2_X1 U363 ( .A1(n161), .A2(n153), .ZN(n151) );
  AOI21_X1 U364 ( .B1(n153), .B2(n162), .A(n154), .ZN(n152) );
  NOR2_X1 U365 ( .A1(n158), .A2(n155), .ZN(n153) );
  INV_X1 U366 ( .A(n126), .ZN(n124) );
  OAI21_X1 U367 ( .B1(n155), .B2(n159), .A(n156), .ZN(n154) );
  XOR2_X1 U368 ( .A(n371), .B(n15), .Z(SUM[18]) );
  NAND2_X1 U369 ( .A1(n199), .A2(n96), .ZN(n15) );
  INV_X1 U370 ( .A(n95), .ZN(n199) );
  XOR2_X1 U371 ( .A(n357), .B(n17), .Z(SUM[16]) );
  NAND2_X1 U372 ( .A1(n201), .A2(n104), .ZN(n17) );
  INV_X1 U373 ( .A(n103), .ZN(n201) );
  NAND2_X1 U374 ( .A1(n187), .A2(n48), .ZN(n3) );
  INV_X1 U375 ( .A(n47), .ZN(n187) );
  NAND2_X1 U376 ( .A1(n189), .A2(n56), .ZN(n5) );
  INV_X1 U377 ( .A(n55), .ZN(n189) );
  NAND2_X1 U378 ( .A1(n191), .A2(n64), .ZN(n7) );
  INV_X1 U379 ( .A(n63), .ZN(n191) );
  NAND2_X1 U380 ( .A1(n193), .A2(n72), .ZN(n9) );
  INV_X1 U381 ( .A(n71), .ZN(n193) );
  NAND2_X1 U382 ( .A1(n404), .A2(n45), .ZN(n2) );
  XNOR2_X1 U383 ( .A(n379), .B(n4), .ZN(SUM[29]) );
  NAND2_X1 U384 ( .A1(n403), .A2(n53), .ZN(n4) );
  NAND2_X1 U385 ( .A1(n402), .A2(n61), .ZN(n6) );
  XNOR2_X1 U386 ( .A(n364), .B(n8), .ZN(SUM[25]) );
  NAND2_X1 U387 ( .A1(n401), .A2(n69), .ZN(n8) );
  NAND2_X1 U388 ( .A1(n399), .A2(n77), .ZN(n10) );
  NAND2_X1 U389 ( .A1(n397), .A2(n85), .ZN(n12) );
  NAND2_X1 U390 ( .A1(n400), .A2(n93), .ZN(n14) );
  NAND2_X1 U391 ( .A1(n398), .A2(n101), .ZN(n16) );
  XOR2_X1 U392 ( .A(n122), .B(n20), .Z(SUM[13]) );
  NAND2_X1 U393 ( .A1(n395), .A2(n121), .ZN(n20) );
  AOI21_X1 U394 ( .B1(n127), .B2(n394), .A(n124), .ZN(n122) );
  XOR2_X1 U395 ( .A(n134), .B(n22), .Z(SUM[11]) );
  NAND2_X1 U396 ( .A1(n206), .A2(n133), .ZN(n22) );
  AOI21_X1 U397 ( .B1(n139), .B2(n207), .A(n136), .ZN(n134) );
  INV_X1 U398 ( .A(n168), .ZN(n213) );
  INV_X1 U399 ( .A(n137), .ZN(n207) );
  XOR2_X1 U400 ( .A(n160), .B(n27), .Z(SUM[6]) );
  NAND2_X1 U401 ( .A1(n211), .A2(n159), .ZN(n27) );
  INV_X1 U402 ( .A(n158), .ZN(n211) );
  INV_X1 U403 ( .A(n169), .ZN(n167) );
  INV_X1 U404 ( .A(n138), .ZN(n136) );
  INV_X1 U405 ( .A(n155), .ZN(n210) );
  INV_X1 U406 ( .A(n163), .ZN(n212) );
  INV_X1 U407 ( .A(n372), .ZN(n214) );
  XOR2_X1 U408 ( .A(n165), .B(n28), .Z(SUM[5]) );
  NAND2_X1 U409 ( .A1(n212), .A2(n164), .ZN(n28) );
  AOI21_X1 U410 ( .B1(n170), .B2(n213), .A(n167), .ZN(n165) );
  XNOR2_X1 U411 ( .A(n170), .B(n29), .ZN(SUM[4]) );
  NAND2_X1 U412 ( .A1(n213), .A2(n169), .ZN(n29) );
  XNOR2_X1 U413 ( .A(n176), .B(n30), .ZN(SUM[3]) );
  NAND2_X1 U414 ( .A1(n214), .A2(n175), .ZN(n30) );
  OAI21_X1 U415 ( .B1(n179), .B2(n177), .A(n178), .ZN(n176) );
  XOR2_X1 U416 ( .A(n179), .B(n31), .Z(SUM[2]) );
  NAND2_X1 U417 ( .A1(n215), .A2(n178), .ZN(n31) );
  INV_X1 U418 ( .A(n177), .ZN(n215) );
  XOR2_X1 U419 ( .A(n32), .B(n184), .Z(SUM[1]) );
  NAND2_X1 U420 ( .A1(n216), .A2(n182), .ZN(n32) );
  INV_X1 U421 ( .A(n181), .ZN(n216) );
  AND2_X1 U422 ( .A1(n347), .A2(n184), .ZN(SUM[0]) );
  NAND2_X1 U423 ( .A1(n203), .A2(n112), .ZN(n19) );
  INV_X1 U424 ( .A(n111), .ZN(n203) );
  NAND2_X1 U425 ( .A1(n396), .A2(n109), .ZN(n18) );
  XNOR2_X1 U426 ( .A(n127), .B(n21), .ZN(SUM[12]) );
  NAND2_X1 U427 ( .A1(n394), .A2(n126), .ZN(n21) );
  XNOR2_X1 U428 ( .A(n139), .B(n23), .ZN(SUM[10]) );
  NAND2_X1 U429 ( .A1(n207), .A2(n138), .ZN(n23) );
  XNOR2_X1 U430 ( .A(n146), .B(n24), .ZN(SUM[9]) );
  NAND2_X1 U431 ( .A1(n208), .A2(n145), .ZN(n24) );
  OAI21_X1 U432 ( .B1(n149), .B2(n147), .A(n148), .ZN(n146) );
  XOR2_X1 U433 ( .A(n149), .B(n25), .Z(SUM[8]) );
  NAND2_X1 U434 ( .A1(n209), .A2(n148), .ZN(n25) );
  INV_X1 U435 ( .A(n147), .ZN(n209) );
  XNOR2_X1 U436 ( .A(n157), .B(n26), .ZN(SUM[7]) );
  NAND2_X1 U437 ( .A1(n210), .A2(n156), .ZN(n26) );
  OAI21_X1 U438 ( .B1(n160), .B2(n158), .A(n159), .ZN(n157) );
  NOR2_X1 U439 ( .A1(B[6]), .A2(A[6]), .ZN(n158) );
  NOR2_X1 U440 ( .A1(B[2]), .A2(A[2]), .ZN(n177) );
  NOR2_X1 U441 ( .A1(B[8]), .A2(A[8]), .ZN(n147) );
  NOR2_X1 U442 ( .A1(B[4]), .A2(A[4]), .ZN(n168) );
  NOR2_X1 U443 ( .A1(B[1]), .A2(A[1]), .ZN(n181) );
  NAND2_X1 U444 ( .A1(B[6]), .A2(A[6]), .ZN(n159) );
  NAND2_X1 U445 ( .A1(B[2]), .A2(A[2]), .ZN(n178) );
  NAND2_X1 U446 ( .A1(B[0]), .A2(A[0]), .ZN(n184) );
  NAND2_X1 U447 ( .A1(B[4]), .A2(A[4]), .ZN(n169) );
  NOR2_X1 U448 ( .A1(B[14]), .A2(A[14]), .ZN(n111) );
  NAND2_X1 U449 ( .A1(B[8]), .A2(A[8]), .ZN(n148) );
  NAND2_X1 U450 ( .A1(B[5]), .A2(A[5]), .ZN(n164) );
  NAND2_X1 U451 ( .A1(B[7]), .A2(A[7]), .ZN(n156) );
  NAND2_X1 U452 ( .A1(B[3]), .A2(A[3]), .ZN(n175) );
  NAND2_X1 U453 ( .A1(B[1]), .A2(A[1]), .ZN(n182) );
  NAND2_X1 U454 ( .A1(B[11]), .A2(A[11]), .ZN(n133) );
  NAND2_X1 U455 ( .A1(B[10]), .A2(A[10]), .ZN(n138) );
  INV_X1 U456 ( .A(n41), .ZN(n185) );
  INV_X1 U457 ( .A(n45), .ZN(n43) );
  NOR2_X1 U458 ( .A1(B[10]), .A2(A[10]), .ZN(n137) );
  NOR2_X1 U459 ( .A1(B[20]), .A2(A[20]), .ZN(n87) );
  NOR2_X1 U460 ( .A1(B[18]), .A2(A[18]), .ZN(n95) );
  NOR2_X1 U461 ( .A1(B[16]), .A2(A[16]), .ZN(n103) );
  NOR2_X1 U462 ( .A1(B[30]), .A2(A[30]), .ZN(n47) );
  NOR2_X1 U463 ( .A1(B[28]), .A2(A[28]), .ZN(n55) );
  NOR2_X1 U464 ( .A1(B[26]), .A2(A[26]), .ZN(n63) );
  NOR2_X1 U465 ( .A1(B[24]), .A2(A[24]), .ZN(n71) );
  NOR2_X1 U466 ( .A1(B[22]), .A2(A[22]), .ZN(n79) );
  OR2_X1 U467 ( .A1(B[21]), .A2(A[21]), .ZN(n397) );
  OR2_X1 U468 ( .A1(B[17]), .A2(A[17]), .ZN(n398) );
  OR2_X1 U469 ( .A1(B[23]), .A2(A[23]), .ZN(n399) );
  NAND2_X1 U470 ( .A1(B[19]), .A2(A[19]), .ZN(n93) );
  NAND2_X1 U471 ( .A1(B[15]), .A2(A[15]), .ZN(n109) );
  NAND2_X1 U472 ( .A1(B[12]), .A2(A[12]), .ZN(n126) );
  NAND2_X1 U473 ( .A1(B[13]), .A2(A[13]), .ZN(n121) );
  NAND2_X1 U474 ( .A1(B[21]), .A2(A[21]), .ZN(n85) );
  NAND2_X1 U475 ( .A1(B[17]), .A2(A[17]), .ZN(n101) );
  NAND2_X1 U476 ( .A1(B[23]), .A2(A[23]), .ZN(n77) );
  NAND2_X1 U477 ( .A1(B[25]), .A2(A[25]), .ZN(n69) );
  NAND2_X1 U478 ( .A1(B[27]), .A2(A[27]), .ZN(n61) );
  NAND2_X1 U479 ( .A1(B[29]), .A2(A[29]), .ZN(n53) );
  NAND2_X1 U480 ( .A1(B[31]), .A2(A[31]), .ZN(n45) );
  NAND2_X1 U481 ( .A1(B[14]), .A2(A[14]), .ZN(n112) );
  NAND2_X1 U482 ( .A1(B[20]), .A2(A[20]), .ZN(n88) );
  NAND2_X1 U483 ( .A1(B[18]), .A2(A[18]), .ZN(n96) );
  NAND2_X1 U484 ( .A1(B[16]), .A2(A[16]), .ZN(n104) );
  NAND2_X1 U485 ( .A1(B[30]), .A2(A[30]), .ZN(n48) );
  NAND2_X1 U486 ( .A1(B[28]), .A2(A[28]), .ZN(n56) );
  NAND2_X1 U487 ( .A1(B[26]), .A2(A[26]), .ZN(n64) );
  NAND2_X1 U488 ( .A1(B[24]), .A2(A[24]), .ZN(n72) );
  NAND2_X1 U489 ( .A1(B[22]), .A2(A[22]), .ZN(n80) );
  OR2_X1 U490 ( .A1(B[19]), .A2(A[19]), .ZN(n400) );
  OR2_X1 U491 ( .A1(B[25]), .A2(A[25]), .ZN(n401) );
  OR2_X1 U492 ( .A1(B[27]), .A2(A[27]), .ZN(n402) );
  OR2_X1 U493 ( .A1(B[29]), .A2(A[29]), .ZN(n403) );
  OR2_X1 U494 ( .A1(B[31]), .A2(A[31]), .ZN(n404) );
  XNOR2_X1 U495 ( .A(n34), .B(n405), .ZN(SUM[39]) );
  XNOR2_X1 U496 ( .A(A[39]), .B(B[39]), .ZN(n405) );
  OAI21_X1 U497 ( .B1(n73), .B2(n71), .A(n72), .ZN(n70) );
  XOR2_X1 U498 ( .A(n384), .B(n9), .Z(SUM[24]) );
  XNOR2_X1 U499 ( .A(n366), .B(n16), .ZN(SUM[17]) );
  XNOR2_X1 U500 ( .A(n362), .B(n14), .ZN(SUM[19]) );
  AOI21_X1 U501 ( .B1(n94), .B2(n400), .A(n91), .ZN(n89) );
  OAI21_X1 U502 ( .B1(n144), .B2(n148), .A(n145), .ZN(n143) );
  NOR2_X1 U503 ( .A1(n147), .A2(n373), .ZN(n142) );
  INV_X1 U504 ( .A(n373), .ZN(n208) );
  OAI21_X1 U505 ( .B1(n132), .B2(n138), .A(n133), .ZN(n131) );
  NOR2_X1 U506 ( .A1(n137), .A2(n374), .ZN(n130) );
  INV_X1 U507 ( .A(n374), .ZN(n206) );
  XNOR2_X1 U508 ( .A(n380), .B(n10), .ZN(SUM[23]) );
  NAND2_X1 U509 ( .A1(B[9]), .A2(A[9]), .ZN(n145) );
  XNOR2_X1 U510 ( .A(n349), .B(n12), .ZN(SUM[21]) );
  XOR2_X1 U511 ( .A(n359), .B(n5), .Z(SUM[28]) );
  XNOR2_X1 U512 ( .A(n354), .B(n6), .ZN(SUM[27]) );
  XNOR2_X1 U513 ( .A(n355), .B(n18), .ZN(SUM[15]) );
  XOR2_X1 U514 ( .A(n381), .B(n7), .Z(SUM[26]) );
  XOR2_X1 U515 ( .A(n365), .B(n13), .Z(SUM[20]) );
  OAI21_X1 U516 ( .B1(n65), .B2(n63), .A(n64), .ZN(n62) );
  OAI21_X1 U517 ( .B1(n89), .B2(n87), .A(n88), .ZN(n86) );
  OAI21_X1 U518 ( .B1(n97), .B2(n95), .A(n96), .ZN(n94) );
  OAI21_X1 U519 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  OAI21_X1 U520 ( .B1(n105), .B2(n103), .A(n104), .ZN(n102) );
  AOI21_X1 U521 ( .B1(n54), .B2(n403), .A(n51), .ZN(n49) );
  XNOR2_X1 U522 ( .A(n346), .B(n2), .ZN(SUM[31]) );
  XOR2_X1 U523 ( .A(n361), .B(n19), .Z(SUM[14]) );
  XOR2_X1 U524 ( .A(n358), .B(n11), .Z(SUM[22]) );
  XOR2_X1 U525 ( .A(n383), .B(n3), .Z(SUM[30]) );
  AOI21_X1 U526 ( .B1(n46), .B2(n404), .A(n43), .ZN(n41) );
  OAI21_X1 U527 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  OAI21_X1 U528 ( .B1(n81), .B2(n79), .A(n80), .ZN(n78) );
endmodule


module mac_3 ( clk, clear_acc, a, b, mac_out );
  input [19:0] a;
  input [19:0] b;
  output [39:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, n2, n3;
  wire   [39:0] mul;
  wire   [39:0] pipeline;
  wire   [39:0] sum;

  DFF_X1 \pipeline_reg[37]  ( .D(mul[37]), .CK(clk), .Q(pipeline[37]) );
  DFF_X1 \pipeline_reg[36]  ( .D(mul[36]), .CK(clk), .Q(pipeline[36]) );
  DFF_X1 \pipeline_reg[35]  ( .D(mul[35]), .CK(clk), .Q(pipeline[35]) );
  DFF_X1 \pipeline_reg[34]  ( .D(mul[34]), .CK(clk), .Q(pipeline[34]) );
  DFF_X1 \pipeline_reg[33]  ( .D(mul[33]), .CK(clk), .Q(pipeline[33]) );
  DFF_X1 \pipeline_reg[32]  ( .D(mul[32]), .CK(clk), .Q(pipeline[32]) );
  DFF_X1 \pipeline_reg[31]  ( .D(mul[31]), .CK(clk), .Q(pipeline[31]) );
  DFF_X1 \pipeline_reg[30]  ( .D(mul[30]), .CK(clk), .Q(pipeline[30]) );
  DFF_X1 \pipeline_reg[29]  ( .D(mul[29]), .CK(clk), .Q(pipeline[29]) );
  DFF_X1 \pipeline_reg[28]  ( .D(mul[28]), .CK(clk), .Q(pipeline[28]) );
  DFF_X1 \pipeline_reg[27]  ( .D(mul[27]), .CK(clk), .Q(pipeline[27]) );
  DFF_X1 \pipeline_reg[26]  ( .D(mul[26]), .CK(clk), .Q(pipeline[26]) );
  DFF_X1 \pipeline_reg[25]  ( .D(mul[25]), .CK(clk), .Q(pipeline[25]) );
  DFF_X1 \pipeline_reg[24]  ( .D(mul[24]), .CK(clk), .Q(pipeline[24]) );
  DFF_X1 \pipeline_reg[23]  ( .D(mul[23]), .CK(clk), .Q(pipeline[23]) );
  DFF_X1 \pipeline_reg[22]  ( .D(mul[22]), .CK(clk), .Q(pipeline[22]) );
  DFF_X1 \pipeline_reg[21]  ( .D(mul[21]), .CK(clk), .Q(pipeline[21]) );
  DFF_X1 \pipeline_reg[20]  ( .D(mul[20]), .CK(clk), .Q(pipeline[20]) );
  DFF_X1 \pipeline_reg[19]  ( .D(mul[19]), .CK(clk), .Q(pipeline[19]) );
  DFF_X1 \pipeline_reg[18]  ( .D(mul[18]), .CK(clk), .Q(pipeline[18]) );
  DFF_X1 \pipeline_reg[17]  ( .D(mul[17]), .CK(clk), .Q(pipeline[17]) );
  DFF_X1 \pipeline_reg[16]  ( .D(mul[16]), .CK(clk), .Q(pipeline[16]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \mac_out_reg[16]  ( .D(N19), .CK(clk), .Q(mac_out[16]) );
  DFF_X1 \mac_out_reg[17]  ( .D(N20), .CK(clk), .Q(mac_out[17]) );
  DFF_X1 \mac_out_reg[18]  ( .D(N21), .CK(clk), .Q(mac_out[18]) );
  DFF_X1 \mac_out_reg[19]  ( .D(N22), .CK(clk), .Q(mac_out[19]) );
  DFF_X1 \mac_out_reg[20]  ( .D(N23), .CK(clk), .Q(mac_out[20]) );
  DFF_X1 \mac_out_reg[21]  ( .D(N24), .CK(clk), .Q(mac_out[21]) );
  DFF_X1 \mac_out_reg[22]  ( .D(N25), .CK(clk), .Q(mac_out[22]) );
  DFF_X1 \mac_out_reg[23]  ( .D(N26), .CK(clk), .Q(mac_out[23]) );
  DFF_X1 \mac_out_reg[24]  ( .D(N27), .CK(clk), .Q(mac_out[24]) );
  DFF_X1 \mac_out_reg[25]  ( .D(N28), .CK(clk), .Q(mac_out[25]) );
  DFF_X1 \mac_out_reg[26]  ( .D(N29), .CK(clk), .Q(mac_out[26]) );
  DFF_X1 \mac_out_reg[27]  ( .D(N30), .CK(clk), .Q(mac_out[27]) );
  DFF_X1 \mac_out_reg[28]  ( .D(N31), .CK(clk), .Q(mac_out[28]) );
  DFF_X1 \mac_out_reg[29]  ( .D(N32), .CK(clk), .Q(mac_out[29]) );
  DFF_X1 \mac_out_reg[30]  ( .D(N33), .CK(clk), .Q(mac_out[30]) );
  DFF_X1 \mac_out_reg[31]  ( .D(N34), .CK(clk), .Q(mac_out[31]) );
  DFF_X1 \mac_out_reg[32]  ( .D(N35), .CK(clk), .Q(mac_out[32]) );
  DFF_X1 \mac_out_reg[33]  ( .D(N36), .CK(clk), .Q(mac_out[33]) );
  DFF_X1 \mac_out_reg[34]  ( .D(N37), .CK(clk), .Q(mac_out[34]) );
  DFF_X1 \mac_out_reg[35]  ( .D(N38), .CK(clk), .Q(mac_out[35]) );
  DFF_X1 \mac_out_reg[36]  ( .D(N39), .CK(clk), .Q(mac_out[36]) );
  DFF_X1 \mac_out_reg[37]  ( .D(N40), .CK(clk), .Q(mac_out[37]) );
  DFF_X1 \mac_out_reg[38]  ( .D(N41), .CK(clk), .Q(mac_out[38]) );
  DFF_X1 \mac_out_reg[39]  ( .D(N42), .CK(clk), .Q(mac_out[39]) );
  mac_3_DW_mult_tc_1 mult_355 ( .a(a), .b(b), .product(mul) );
  mac_3_DW01_add_1 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  DFF_X1 \pipeline_reg[38]  ( .D(mul[38]), .CK(clk), .Q(pipeline[38]) );
  DFF_X2 \pipeline_reg[39]  ( .D(mul[39]), .CK(clk), .Q(pipeline[39]) );
  BUF_X1 U3 ( .A(n3), .Z(n2) );
  INV_X1 U4 ( .A(clear_acc), .ZN(n3) );
  AND2_X1 U6 ( .A1(sum[39]), .A2(n2), .ZN(N42) );
  AND2_X1 U7 ( .A1(sum[38]), .A2(n2), .ZN(N41) );
  AND2_X1 U8 ( .A1(sum[37]), .A2(n2), .ZN(N40) );
  AND2_X1 U9 ( .A1(sum[36]), .A2(n2), .ZN(N39) );
  AND2_X1 U10 ( .A1(sum[35]), .A2(n2), .ZN(N38) );
  AND2_X1 U11 ( .A1(sum[34]), .A2(n2), .ZN(N37) );
  AND2_X1 U12 ( .A1(sum[33]), .A2(n2), .ZN(N36) );
  AND2_X1 U13 ( .A1(sum[32]), .A2(n2), .ZN(N35) );
  AND2_X1 U14 ( .A1(sum[31]), .A2(n2), .ZN(N34) );
  AND2_X1 U15 ( .A1(sum[30]), .A2(n2), .ZN(N33) );
  AND2_X1 U16 ( .A1(sum[29]), .A2(n2), .ZN(N32) );
  AND2_X1 U17 ( .A1(sum[28]), .A2(n3), .ZN(N31) );
  AND2_X1 U18 ( .A1(sum[27]), .A2(n3), .ZN(N30) );
  AND2_X1 U19 ( .A1(sum[26]), .A2(n3), .ZN(N29) );
  AND2_X1 U20 ( .A1(sum[25]), .A2(n3), .ZN(N28) );
  AND2_X1 U21 ( .A1(sum[24]), .A2(n3), .ZN(N27) );
  AND2_X1 U22 ( .A1(sum[23]), .A2(n3), .ZN(N26) );
  AND2_X1 U23 ( .A1(sum[22]), .A2(n3), .ZN(N25) );
  AND2_X1 U24 ( .A1(sum[21]), .A2(n3), .ZN(N24) );
  AND2_X1 U25 ( .A1(sum[20]), .A2(n3), .ZN(N23) );
  AND2_X1 U26 ( .A1(sum[19]), .A2(n3), .ZN(N22) );
  AND2_X1 U27 ( .A1(sum[18]), .A2(n3), .ZN(N21) );
  AND2_X1 U28 ( .A1(sum[17]), .A2(n3), .ZN(N20) );
  AND2_X1 U29 ( .A1(sum[16]), .A2(n3), .ZN(N19) );
  AND2_X1 U30 ( .A1(sum[15]), .A2(n3), .ZN(N18) );
  AND2_X1 U31 ( .A1(sum[14]), .A2(n3), .ZN(N17) );
  AND2_X1 U32 ( .A1(sum[13]), .A2(n3), .ZN(N16) );
  AND2_X1 U33 ( .A1(sum[12]), .A2(n3), .ZN(N15) );
  AND2_X1 U34 ( .A1(sum[11]), .A2(n3), .ZN(N14) );
  AND2_X1 U35 ( .A1(sum[10]), .A2(n3), .ZN(N13) );
  AND2_X1 U36 ( .A1(sum[9]), .A2(n3), .ZN(N12) );
  AND2_X1 U37 ( .A1(sum[8]), .A2(n3), .ZN(N11) );
  AND2_X1 U38 ( .A1(sum[7]), .A2(n3), .ZN(N10) );
  AND2_X1 U39 ( .A1(sum[6]), .A2(n3), .ZN(N9) );
  AND2_X1 U40 ( .A1(sum[5]), .A2(n3), .ZN(N8) );
  AND2_X1 U41 ( .A1(sum[4]), .A2(n3), .ZN(N7) );
  AND2_X1 U42 ( .A1(sum[3]), .A2(n3), .ZN(N6) );
  AND2_X1 U43 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U44 ( .A1(sum[1]), .A2(n3), .ZN(N4) );
  AND2_X1 U45 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
endmodule


module mac_2_DW_mult_tc_1 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n4, n6, n7, n9, n12, n13, n16, n18, n19, n24, n25, n28, n31, n34,
         n37, n42, n43, n46, n49, n52, n54, n55, n58, n60, n61, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n97, n98, n99, n100, n101, n103, n105, n106, n107, n108, n109,
         n111, n113, n114, n115, n116, n117, n119, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n141, n142, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n185,
         n186, n187, n188, n193, n194, n195, n196, n198, n200, n201, n202,
         n203, n204, n205, n206, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n225, n227,
         n228, n230, n232, n233, n234, n236, n238, n239, n240, n241, n242,
         n244, n246, n247, n248, n249, n250, n252, n254, n255, n256, n257,
         n258, n259, n260, n261, n263, n264, n266, n268, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n284, n285, n286,
         n287, n291, n293, n295, n296, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n643, n644, n646,
         n647, n649, n652, n653, n655, n656, n658, n659, n661, n662, n664,
         n665, n667, n668, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1115, n1116, n1119, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1233, n1234, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n37 = a[13];
  assign n43 = a[15];
  assign n49 = a[17];
  assign n55 = a[19];
  assign n61 = b[0];
  assign n668 = a[0];
  assign n1090 = b[19];
  assign n1091 = b[18];
  assign n1092 = b[17];
  assign n1093 = b[16];
  assign n1094 = b[15];
  assign n1095 = b[14];
  assign n1096 = b[13];
  assign n1097 = b[12];
  assign n1098 = b[11];
  assign n1099 = b[10];
  assign n1100 = b[9];
  assign n1101 = b[8];
  assign n1102 = b[7];
  assign n1103 = b[6];
  assign n1104 = b[5];
  assign n1105 = b[4];
  assign n1106 = b[3];
  assign n1107 = b[2];
  assign n1108 = b[1];

  FA_X1 U333 ( .A(n681), .B(n304), .CI(n700), .CO(n300), .S(n301) );
  FA_X1 U334 ( .A(n305), .B(n682), .CI(n308), .CO(n302), .S(n303) );
  FA_X1 U336 ( .A(n312), .B(n683), .CI(n309), .CO(n306), .S(n307) );
  FA_X1 U337 ( .A(n701), .B(n314), .CI(n720), .CO(n308), .S(n309) );
  FA_X1 U338 ( .A(n313), .B(n320), .CI(n318), .CO(n310), .S(n311) );
  FA_X1 U339 ( .A(n684), .B(n702), .CI(n315), .CO(n312), .S(n313) );
  FA_X1 U341 ( .A(n324), .B(n321), .CI(n319), .CO(n316), .S(n317) );
  FA_X1 U342 ( .A(n328), .B(n721), .CI(n326), .CO(n318), .S(n319) );
  FA_X1 U343 ( .A(n703), .B(n685), .CI(n740), .CO(n320), .S(n321) );
  FA_X1 U344 ( .A(n325), .B(n327), .CI(n332), .CO(n322), .S(n323) );
  FA_X1 U345 ( .A(n336), .B(n329), .CI(n334), .CO(n324), .S(n325) );
  FA_X1 U346 ( .A(n686), .B(n704), .CI(n722), .CO(n326), .S(n327) );
  FA_X1 U348 ( .A(n340), .B(n342), .CI(n333), .CO(n330), .S(n331) );
  FA_X1 U349 ( .A(n335), .B(n344), .CI(n337), .CO(n332), .S(n333) );
  FA_X1 U350 ( .A(n705), .B(n346), .CI(n723), .CO(n334), .S(n335) );
  FA_X1 U351 ( .A(n741), .B(n687), .CI(n760), .CO(n336), .S(n337) );
  FA_X1 U352 ( .A(n350), .B(n343), .CI(n341), .CO(n338), .S(n339) );
  FA_X1 U353 ( .A(n345), .B(n354), .CI(n352), .CO(n340), .S(n341) );
  FA_X1 U354 ( .A(n347), .B(n724), .CI(n356), .CO(n342), .S(n343) );
  FA_X1 U355 ( .A(n742), .B(n706), .CI(n688), .CO(n344), .S(n345) );
  FA_X1 U357 ( .A(n360), .B(n353), .CI(n351), .CO(n348), .S(n349) );
  FA_X1 U358 ( .A(n357), .B(n355), .CI(n362), .CO(n350), .S(n351) );
  FA_X1 U359 ( .A(n366), .B(n743), .CI(n364), .CO(n352), .S(n353) );
  FA_X1 U360 ( .A(n707), .B(n761), .CI(n725), .CO(n354), .S(n355) );
  FA_X1 U361 ( .A(n368), .B(n689), .CI(n780), .CO(n356), .S(n357) );
  FA_X1 U362 ( .A(n372), .B(n363), .CI(n361), .CO(n358), .S(n359) );
  FA_X1 U363 ( .A(n376), .B(n365), .CI(n374), .CO(n360), .S(n361) );
  FA_X1 U364 ( .A(n378), .B(n380), .CI(n367), .CO(n362), .S(n363) );
  FA_X1 U365 ( .A(n690), .B(n708), .CI(n369), .CO(n364), .S(n365) );
  FA_X1 U366 ( .A(n762), .B(n726), .CI(n744), .CO(n366), .S(n367) );
  FA_X1 U368 ( .A(n384), .B(n375), .CI(n373), .CO(n370), .S(n371) );
  FA_X1 U369 ( .A(n377), .B(n388), .CI(n386), .CO(n372), .S(n373) );
  FA_X1 U370 ( .A(n379), .B(n390), .CI(n381), .CO(n374), .S(n375) );
  FA_X1 U371 ( .A(n727), .B(n745), .CI(n392), .CO(n376), .S(n377) );
  FA_X1 U372 ( .A(n709), .B(n781), .CI(n763), .CO(n378), .S(n379) );
  FA_X1 U373 ( .A(n394), .B(n691), .CI(n800), .CO(n380), .S(n381) );
  FA_X1 U374 ( .A(n398), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U375 ( .A(n389), .B(n402), .CI(n400), .CO(n384), .S(n385) );
  FA_X1 U376 ( .A(n393), .B(n404), .CI(n391), .CO(n386), .S(n387) );
  FA_X1 U377 ( .A(n408), .B(n395), .CI(n406), .CO(n388), .S(n389) );
  FA_X1 U378 ( .A(n746), .B(n782), .CI(n764), .CO(n390), .S(n391) );
  FA_X1 U379 ( .A(n710), .B(n728), .CI(n692), .CO(n392), .S(n393) );
  FA_X1 U381 ( .A(n412), .B(n401), .CI(n399), .CO(n396), .S(n397) );
  FA_X1 U382 ( .A(n403), .B(n416), .CI(n414), .CO(n398), .S(n399) );
  FA_X1 U383 ( .A(n409), .B(n407), .CI(n418), .CO(n400), .S(n401) );
  FA_X1 U384 ( .A(n420), .B(n422), .CI(n405), .CO(n402), .S(n403) );
  FA_X1 U385 ( .A(n729), .B(n747), .CI(n765), .CO(n404), .S(n405) );
  FA_X1 U386 ( .A(n711), .B(n783), .CI(n801), .CO(n406), .S(n407) );
  FA_X1 U387 ( .A(n424), .B(n693), .CI(n820), .CO(n408), .S(n409) );
  FA_X1 U388 ( .A(n428), .B(n415), .CI(n413), .CO(n410), .S(n411) );
  FA_X1 U389 ( .A(n417), .B(n432), .CI(n430), .CO(n412), .S(n413) );
  FA_X1 U391 ( .A(n436), .B(n438), .CI(n421), .CO(n416), .S(n417) );
  FA_X1 U392 ( .A(n425), .B(n748), .CI(n440), .CO(n418), .S(n419) );
  FA_X1 U393 ( .A(n694), .B(n712), .CI(n766), .CO(n420), .S(n421) );
  FA_X1 U394 ( .A(n802), .B(n730), .CI(n784), .CO(n422), .S(n423) );
  FA_X1 U397 ( .A(n433), .B(n448), .CI(n446), .CO(n428), .S(n429) );
  FA_X1 U399 ( .A(n437), .B(n452), .CI(n439), .CO(n432), .S(n433) );
  FA_X1 U400 ( .A(n456), .B(n767), .CI(n454), .CO(n434), .S(n435) );
  FA_X1 U401 ( .A(n731), .B(n785), .CI(n749), .CO(n436), .S(n437) );
  FA_X1 U402 ( .A(n458), .B(n803), .CI(n713), .CO(n438), .S(n439) );
  FA_X1 U403 ( .A(n840), .B(n695), .CI(n821), .CO(n440), .S(n441) );
  FA_X1 U404 ( .A(n462), .B(n447), .CI(n445), .CO(n442), .S(n443) );
  FA_X1 U405 ( .A(n449), .B(n466), .CI(n464), .CO(n444), .S(n445) );
  FA_X1 U407 ( .A(n455), .B(n470), .CI(n457), .CO(n448), .S(n449) );
  FA_X1 U408 ( .A(n472), .B(n476), .CI(n474), .CO(n450), .S(n451) );
  FA_X1 U409 ( .A(n768), .B(n786), .CI(n459), .CO(n452), .S(n453) );
  FA_X1 U410 ( .A(n714), .B(n732), .CI(n804), .CO(n454), .S(n455) );
  FA_X1 U414 ( .A(n467), .B(n484), .CI(n482), .CO(n462), .S(n463) );
  FA_X1 U416 ( .A(n473), .B(n488), .CI(n475), .CO(n466), .S(n467) );
  FA_X1 U417 ( .A(n490), .B(n477), .CI(n492), .CO(n468), .S(n469) );
  FA_X1 U418 ( .A(n805), .B(n823), .CI(n494), .CO(n470), .S(n471) );
  FA_X1 U419 ( .A(n733), .B(n841), .CI(n751), .CO(n472), .S(n473) );
  FA_X1 U420 ( .A(n697), .B(n860), .CI(n769), .CO(n474), .S(n475) );
  FA_X1 U423 ( .A(n498), .B(n483), .CI(n481), .CO(n478), .S(n479) );
  FA_X1 U424 ( .A(n500), .B(n487), .CI(n485), .CO(n480), .S(n481) );
  FA_X1 U426 ( .A(n489), .B(n506), .CI(n491), .CO(n484), .S(n485) );
  FA_X1 U428 ( .A(n770), .B(n842), .CI(n824), .CO(n488), .S(n489) );
  FA_X1 U430 ( .A(n734), .B(n670), .CI(n788), .CO(n492), .S(n493) );
  HA_X1 U431 ( .A(n698), .B(n716), .CO(n494), .S(n495) );
  FA_X1 U433 ( .A(n516), .B(n505), .CI(n503), .CO(n498), .S(n499) );
  FA_X1 U434 ( .A(n520), .B(n509), .CI(n518), .CO(n500), .S(n501) );
  FA_X1 U436 ( .A(n526), .B(n807), .CI(n524), .CO(n504), .S(n505) );
  FA_X1 U437 ( .A(n771), .B(n789), .CI(n825), .CO(n506), .S(n507) );
  FA_X1 U438 ( .A(n753), .B(n717), .CI(n843), .CO(n508), .S(n509) );
  FA_X1 U442 ( .A(n525), .B(n523), .CI(n534), .CO(n516), .S(n517) );
  FA_X1 U444 ( .A(n826), .B(n844), .CI(n527), .CO(n520), .S(n521) );
  FA_X1 U445 ( .A(n754), .B(n772), .CI(n808), .CO(n522), .S(n523) );
  FA_X1 U446 ( .A(n863), .B(n790), .CI(n671), .CO(n524), .S(n525) );
  HA_X1 U447 ( .A(n736), .B(n718), .CO(n526), .S(n527) );
  FA_X1 U448 ( .A(n544), .B(n533), .CI(n531), .CO(n528), .S(n529) );
  FA_X1 U449 ( .A(n546), .B(n548), .CI(n535), .CO(n530), .S(n531) );
  FA_X1 U450 ( .A(n537), .B(n541), .CI(n539), .CO(n532), .S(n533) );
  FA_X1 U453 ( .A(n737), .B(n845), .CI(n773), .CO(n538), .S(n539) );
  FA_X1 U454 ( .A(n755), .B(n719), .CI(n864), .CO(n540), .S(n541) );
  FA_X1 U458 ( .A(n566), .B(n846), .CI(n555), .CO(n548), .S(n549) );
  FA_X1 U459 ( .A(n865), .B(n792), .CI(n828), .CO(n550), .S(n551) );
  FA_X1 U460 ( .A(n774), .B(n810), .CI(n672), .CO(n552), .S(n553) );
  HA_X1 U461 ( .A(n738), .B(n756), .CO(n554), .S(n555) );
  FA_X1 U462 ( .A(n561), .B(n570), .CI(n559), .CO(n556), .S(n557) );
  FA_X1 U463 ( .A(n563), .B(n565), .CI(n572), .CO(n558), .S(n559) );
  FA_X1 U464 ( .A(n574), .B(n576), .CI(n567), .CO(n560), .S(n561) );
  FA_X1 U466 ( .A(n757), .B(n847), .CI(n793), .CO(n564), .S(n565) );
  FA_X1 U467 ( .A(n866), .B(n739), .CI(n775), .CO(n566), .S(n567) );
  FA_X1 U468 ( .A(n582), .B(n573), .CI(n571), .CO(n568), .S(n569) );
  FA_X1 U469 ( .A(n577), .B(n575), .CI(n584), .CO(n570), .S(n571) );
  FA_X1 U471 ( .A(n794), .B(n848), .CI(n830), .CO(n574), .S(n575) );
  FA_X1 U472 ( .A(n867), .B(n812), .CI(n673), .CO(n576), .S(n577) );
  HA_X1 U473 ( .A(n776), .B(n758), .CO(n578), .S(n579) );
  FA_X1 U474 ( .A(n585), .B(n592), .CI(n583), .CO(n580), .S(n581) );
  FA_X1 U475 ( .A(n587), .B(n589), .CI(n594), .CO(n582), .S(n583) );
  FA_X1 U476 ( .A(n598), .B(n831), .CI(n596), .CO(n584), .S(n585) );
  FA_X1 U478 ( .A(n795), .B(n759), .CI(n868), .CO(n588), .S(n589) );
  FA_X1 U479 ( .A(n602), .B(n595), .CI(n593), .CO(n590), .S(n591) );
  FA_X1 U480 ( .A(n604), .B(n606), .CI(n597), .CO(n592), .S(n593) );
  FA_X1 U481 ( .A(n814), .B(n850), .CI(n599), .CO(n594), .S(n595) );
  FA_X1 U482 ( .A(n869), .B(n832), .CI(n674), .CO(n596), .S(n597) );
  HA_X1 U483 ( .A(n778), .B(n796), .CO(n598), .S(n599) );
  FA_X1 U485 ( .A(n612), .B(n614), .CI(n607), .CO(n602), .S(n603) );
  FA_X1 U486 ( .A(n797), .B(n851), .CI(n833), .CO(n604), .S(n605) );
  FA_X1 U488 ( .A(n613), .B(n618), .CI(n611), .CO(n608), .S(n609) );
  FA_X1 U489 ( .A(n615), .B(n871), .CI(n620), .CO(n610), .S(n611) );
  FA_X1 U490 ( .A(n852), .B(n834), .CI(n675), .CO(n612), .S(n613) );
  HA_X1 U491 ( .A(n798), .B(n816), .CO(n614), .S(n615) );
  FA_X1 U492 ( .A(n621), .B(n624), .CI(n619), .CO(n616), .S(n617) );
  FA_X1 U493 ( .A(n817), .B(n853), .CI(n626), .CO(n618), .S(n619) );
  FA_X1 U494 ( .A(n835), .B(n799), .CI(n872), .CO(n620), .S(n621) );
  FA_X1 U495 ( .A(n630), .B(n627), .CI(n625), .CO(n622), .S(n623) );
  FA_X1 U496 ( .A(n854), .B(n873), .CI(n676), .CO(n624), .S(n625) );
  HA_X1 U497 ( .A(n818), .B(n836), .CO(n626), .S(n627) );
  FA_X1 U498 ( .A(n634), .B(n837), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U499 ( .A(n874), .B(n819), .CI(n855), .CO(n630), .S(n631) );
  FA_X1 U500 ( .A(n677), .B(n856), .CI(n635), .CO(n632), .S(n633) );
  HA_X1 U501 ( .A(n838), .B(n875), .CO(n634), .S(n635) );
  FA_X1 U502 ( .A(n876), .B(n839), .CI(n857), .CO(n636), .S(n637) );
  HA_X1 U503 ( .A(n858), .B(n877), .CO(n638), .S(n639) );
  AND2_X2 U1025 ( .A1(n46), .A2(n1514), .ZN(n1529) );
  CLKBUF_X1 U1026 ( .A(n450), .Z(n1233) );
  BUF_X4 U1027 ( .A(n1329), .Z(n1539) );
  BUF_X2 U1028 ( .A(n1095), .Z(n1584) );
  BUF_X2 U1029 ( .A(n1), .Z(n1470) );
  OR2_X1 U1030 ( .A1(n529), .A2(n542), .ZN(n1312) );
  BUF_X1 U1031 ( .A(n1096), .Z(n1333) );
  BUF_X1 U1032 ( .A(n1096), .Z(n1583) );
  NOR2_X1 U1033 ( .A1(n497), .A2(n512), .ZN(n1234) );
  NOR2_X1 U1034 ( .A1(n497), .A2(n512), .ZN(n177) );
  CLKBUF_X3 U1035 ( .A(n13), .Z(n1252) );
  BUF_X2 U1036 ( .A(n1099), .Z(n1285) );
  BUF_X2 U1037 ( .A(n1099), .Z(n1580) );
  NOR2_X2 U1038 ( .A1(n557), .A2(n568), .ZN(n204) );
  NAND3_X1 U1039 ( .A1(n1289), .A2(n1290), .A3(n1291), .ZN(n536) );
  BUF_X1 U1040 ( .A(n25), .Z(n1564) );
  BUF_X1 U1041 ( .A(n1578), .Z(n1379) );
  AND2_X1 U1042 ( .A1(n1115), .A2(n28), .ZN(n1530) );
  BUF_X2 U1043 ( .A(n31), .Z(n1400) );
  BUF_X1 U1044 ( .A(n1541), .Z(n1495) );
  BUF_X1 U1045 ( .A(n37), .Z(n1566) );
  BUF_X2 U1046 ( .A(n1575), .Z(n1366) );
  BUF_X1 U1047 ( .A(n1106), .Z(n1363) );
  BUF_X2 U1048 ( .A(n1541), .Z(n1496) );
  BUF_X2 U1049 ( .A(n1313), .Z(n1542) );
  BUF_X2 U1050 ( .A(n1329), .Z(n1540) );
  NAND3_X1 U1051 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n486) );
  BUF_X2 U1052 ( .A(n1092), .Z(n1587) );
  NAND3_X1 U1053 ( .A1(n1454), .A2(n1455), .A3(n1456), .ZN(n514) );
  BUF_X2 U1054 ( .A(n1), .Z(n1471) );
  BUF_X2 U1055 ( .A(n6), .Z(n1536) );
  INV_X1 U1056 ( .A(n1312), .ZN(n187) );
  AND2_X1 U1057 ( .A1(n1510), .A2(n263), .ZN(product[1]) );
  BUF_X2 U1058 ( .A(n1104), .Z(n1576) );
  OAI22_X1 U1059 ( .A1(n1486), .A2(n956), .B1(n1324), .B2(n1545), .ZN(n1236)
         );
  XNOR2_X1 U1060 ( .A(n1322), .B(n1271), .ZN(n1237) );
  CLKBUF_X3 U1061 ( .A(n25), .Z(n1271) );
  BUF_X1 U1062 ( .A(n953), .Z(n1238) );
  BUF_X2 U1063 ( .A(n52), .Z(n1498) );
  BUF_X1 U1064 ( .A(n1353), .Z(n1506) );
  NAND2_X1 U1065 ( .A1(n1315), .A2(n1518), .ZN(n1239) );
  NAND2_X1 U1066 ( .A1(n1315), .A2(n1518), .ZN(n1383) );
  CLKBUF_X3 U1067 ( .A(n28), .Z(n1314) );
  BUF_X2 U1068 ( .A(n1100), .Z(n1579) );
  INV_X2 U1069 ( .A(n1142), .ZN(n1323) );
  CLKBUF_X1 U1070 ( .A(n1502), .Z(n1240) );
  INV_X1 U1071 ( .A(n1368), .ZN(n1241) );
  BUF_X2 U1072 ( .A(n1270), .Z(n1532) );
  CLKBUF_X1 U1073 ( .A(n465), .Z(n1242) );
  BUF_X2 U1074 ( .A(n18), .Z(n1262) );
  BUF_X1 U1075 ( .A(n1586), .Z(n1337) );
  OR2_X2 U1076 ( .A1(n1484), .A2(n1399), .ZN(n42) );
  AND2_X1 U1077 ( .A1(n1513), .A2(n34), .ZN(n1243) );
  AND2_X1 U1078 ( .A1(n34), .A2(n1513), .ZN(n1244) );
  AND2_X1 U1079 ( .A1(n1513), .A2(n34), .ZN(n1531) );
  XOR2_X1 U1080 ( .A(n468), .B(n453), .Z(n1245) );
  XOR2_X1 U1081 ( .A(n451), .B(n1245), .Z(n447) );
  NAND2_X1 U1082 ( .A1(n451), .A2(n468), .ZN(n1246) );
  NAND2_X1 U1083 ( .A1(n451), .A2(n453), .ZN(n1247) );
  NAND2_X1 U1084 ( .A1(n468), .A2(n453), .ZN(n1248) );
  NAND3_X1 U1085 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n446) );
  CLKBUF_X2 U1086 ( .A(n7), .Z(n1358) );
  XNOR2_X1 U1087 ( .A(n1377), .B(n1509), .ZN(n1249) );
  CLKBUF_X1 U1088 ( .A(n140), .Z(n1250) );
  OR2_X1 U1089 ( .A1(n150), .A2(n1546), .ZN(n1251) );
  XOR2_X1 U1090 ( .A(n510), .B(n495), .Z(n1253) );
  XOR2_X1 U1091 ( .A(n1253), .B(n508), .Z(n487) );
  NAND2_X1 U1092 ( .A1(n510), .A2(n495), .ZN(n1254) );
  NAND2_X1 U1093 ( .A1(n510), .A2(n508), .ZN(n1255) );
  NAND2_X1 U1094 ( .A1(n495), .A2(n508), .ZN(n1256) );
  XOR2_X1 U1095 ( .A(n471), .B(n469), .Z(n1257) );
  XOR2_X1 U1096 ( .A(n1257), .B(n486), .Z(n465) );
  NAND2_X1 U1097 ( .A1(n471), .A2(n469), .ZN(n1258) );
  NAND2_X1 U1098 ( .A1(n471), .A2(n486), .ZN(n1259) );
  NAND2_X1 U1099 ( .A1(n469), .A2(n486), .ZN(n1260) );
  NAND3_X1 U1100 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n464) );
  BUF_X2 U1101 ( .A(n18), .Z(n1261) );
  CLKBUF_X1 U1102 ( .A(n18), .Z(n1367) );
  BUF_X1 U1103 ( .A(n1578), .Z(n1380) );
  BUF_X2 U1104 ( .A(n1353), .Z(n1505) );
  BUF_X2 U1105 ( .A(n1558), .Z(n1263) );
  CLKBUF_X1 U1106 ( .A(n1485), .Z(n1264) );
  BUF_X2 U1107 ( .A(n1573), .Z(n1265) );
  BUF_X1 U1108 ( .A(n1573), .Z(n1266) );
  BUF_X2 U1109 ( .A(n1107), .Z(n1573) );
  NOR2_X1 U1110 ( .A1(n171), .A2(n1507), .ZN(n1267) );
  NAND2_X1 U1111 ( .A1(n1398), .A2(n302), .ZN(n1268) );
  NAND2_X1 U1112 ( .A1(n98), .A2(n300), .ZN(n1269) );
  XNOR2_X1 U1113 ( .A(a[2]), .B(n1), .ZN(n1270) );
  CLKBUF_X3 U1114 ( .A(n25), .Z(n1385) );
  CLKBUF_X3 U1115 ( .A(n1108), .Z(n1572) );
  CLKBUF_X1 U1116 ( .A(n1101), .Z(n1370) );
  XNOR2_X1 U1117 ( .A(n1272), .B(n536), .ZN(n519) );
  XNOR2_X1 U1118 ( .A(n540), .B(n538), .ZN(n1272) );
  XNOR2_X1 U1119 ( .A(n499), .B(n1273), .ZN(n497) );
  XNOR2_X1 U1120 ( .A(n514), .B(n501), .ZN(n1273) );
  XNOR2_X1 U1121 ( .A(n1354), .B(n1274), .ZN(n457) );
  XNOR2_X1 U1122 ( .A(n822), .B(n696), .ZN(n1274) );
  XNOR2_X1 U1123 ( .A(n1233), .B(n1275), .ZN(n431) );
  XNOR2_X1 U1124 ( .A(n435), .B(n441), .ZN(n1275) );
  OR2_X1 U1125 ( .A1(n513), .A2(n528), .ZN(n1547) );
  BUF_X2 U1126 ( .A(n61), .Z(n1570) );
  BUF_X2 U1127 ( .A(n31), .Z(n1565) );
  BUF_X1 U1128 ( .A(n16), .Z(n1541) );
  XNOR2_X1 U1129 ( .A(n603), .B(n1276), .ZN(n601) );
  XNOR2_X1 U1130 ( .A(n610), .B(n605), .ZN(n1276) );
  XOR2_X1 U1131 ( .A(n522), .B(n511), .Z(n1277) );
  XOR2_X1 U1132 ( .A(n1277), .B(n507), .Z(n503) );
  NAND2_X1 U1133 ( .A1(n511), .A2(n522), .ZN(n1278) );
  NAND2_X1 U1134 ( .A1(n511), .A2(n507), .ZN(n1279) );
  NAND2_X1 U1135 ( .A1(n522), .A2(n507), .ZN(n1280) );
  NAND3_X1 U1136 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n502) );
  XOR2_X1 U1137 ( .A(n504), .B(n493), .Z(n1281) );
  XOR2_X1 U1138 ( .A(n1281), .B(n502), .Z(n483) );
  NAND2_X1 U1139 ( .A1(n504), .A2(n493), .ZN(n1282) );
  NAND2_X1 U1140 ( .A1(n504), .A2(n502), .ZN(n1283) );
  NAND2_X1 U1141 ( .A1(n493), .A2(n502), .ZN(n1284) );
  NAND3_X1 U1142 ( .A1(n1282), .A2(n1283), .A3(n1284), .ZN(n482) );
  CLKBUF_X1 U1143 ( .A(n141), .Z(n1286) );
  BUF_X2 U1144 ( .A(n1585), .Z(n1378) );
  INV_X1 U1145 ( .A(n1530), .ZN(n1492) );
  INV_X1 U1146 ( .A(n1140), .ZN(n1287) );
  CLKBUF_X3 U1147 ( .A(n55), .Z(n1569) );
  XOR2_X1 U1148 ( .A(n791), .B(n827), .Z(n1288) );
  XOR2_X1 U1149 ( .A(n1288), .B(n809), .Z(n537) );
  NAND2_X1 U1150 ( .A1(n791), .A2(n827), .ZN(n1289) );
  NAND2_X1 U1151 ( .A1(n791), .A2(n809), .ZN(n1290) );
  NAND2_X1 U1152 ( .A1(n827), .A2(n809), .ZN(n1291) );
  NAND2_X1 U1153 ( .A1(n540), .A2(n538), .ZN(n1292) );
  NAND2_X1 U1154 ( .A1(n540), .A2(n536), .ZN(n1293) );
  NAND2_X1 U1155 ( .A1(n538), .A2(n536), .ZN(n1294) );
  NAND3_X1 U1156 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n518) );
  CLKBUF_X1 U1157 ( .A(n19), .Z(n1538) );
  NAND2_X1 U1158 ( .A1(n435), .A2(n450), .ZN(n1295) );
  NAND2_X1 U1159 ( .A1(n450), .A2(n441), .ZN(n1296) );
  NAND2_X1 U1160 ( .A1(n435), .A2(n441), .ZN(n1297) );
  NAND3_X1 U1161 ( .A1(n1297), .A2(n1295), .A3(n1296), .ZN(n430) );
  XOR2_X1 U1162 ( .A(n1), .B(n668), .Z(n1119) );
  NAND2_X1 U1163 ( .A1(n603), .A2(n610), .ZN(n1298) );
  NAND2_X1 U1164 ( .A1(n603), .A2(n605), .ZN(n1299) );
  NAND2_X1 U1165 ( .A1(n610), .A2(n605), .ZN(n1300) );
  NAND3_X1 U1166 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n600) );
  OR2_X2 U1167 ( .A1(n1399), .A2(n1484), .ZN(n1486) );
  XOR2_X1 U1168 ( .A(n419), .B(n423), .Z(n1301) );
  XOR2_X1 U1169 ( .A(n434), .B(n1301), .Z(n415) );
  NAND2_X1 U1170 ( .A1(n434), .A2(n419), .ZN(n1302) );
  NAND2_X1 U1171 ( .A1(n434), .A2(n423), .ZN(n1303) );
  NAND2_X1 U1172 ( .A1(n419), .A2(n423), .ZN(n1304) );
  NAND3_X1 U1173 ( .A1(n1302), .A2(n1304), .A3(n1303), .ZN(n414) );
  XNOR2_X1 U1174 ( .A(n735), .B(n1305), .ZN(n511) );
  XNOR2_X1 U1175 ( .A(n862), .B(n699), .ZN(n1305) );
  CLKBUF_X1 U1176 ( .A(n134), .Z(n1306) );
  CLKBUF_X1 U1177 ( .A(n150), .Z(n1307) );
  NOR2_X1 U1178 ( .A1(n426), .A2(n411), .ZN(n150) );
  CLKBUF_X1 U1179 ( .A(n1373), .Z(n1308) );
  NAND3_X1 U1180 ( .A1(n1407), .A2(n1408), .A3(n1409), .ZN(n1309) );
  NAND3_X1 U1181 ( .A1(n1407), .A2(n1408), .A3(n1409), .ZN(n1310) );
  CLKBUF_X1 U1182 ( .A(n1463), .Z(n1311) );
  XNOR2_X1 U1183 ( .A(n1564), .B(a[10]), .ZN(n1313) );
  CLKBUF_X1 U1184 ( .A(n28), .Z(n1537) );
  XOR2_X1 U1185 ( .A(n1538), .B(a[6]), .Z(n1315) );
  CLKBUF_X1 U1186 ( .A(n171), .Z(n1316) );
  XNOR2_X1 U1187 ( .A(n1576), .B(n1567), .ZN(n1317) );
  XNOR2_X1 U1188 ( .A(n1318), .B(n549), .ZN(n545) );
  XNOR2_X1 U1189 ( .A(n560), .B(n553), .ZN(n1318) );
  BUF_X1 U1190 ( .A(n1103), .Z(n1319) );
  CLKBUF_X1 U1191 ( .A(n165), .Z(n1320) );
  CLKBUF_X1 U1192 ( .A(n176), .Z(n1321) );
  BUF_X1 U1193 ( .A(n24), .Z(n1348) );
  BUF_X2 U1194 ( .A(n1578), .Z(n1322) );
  BUF_X2 U1195 ( .A(n1106), .Z(n1574) );
  BUF_X1 U1196 ( .A(n1589), .Z(n1376) );
  XNOR2_X1 U1197 ( .A(n1380), .B(n1387), .ZN(n1324) );
  XNOR2_X1 U1198 ( .A(n1265), .B(n1489), .ZN(n1325) );
  CLKBUF_X1 U1199 ( .A(n1355), .Z(n1326) );
  CLKBUF_X1 U1200 ( .A(n1467), .Z(n1327) );
  XNOR2_X1 U1201 ( .A(n463), .B(n1328), .ZN(n461) );
  XNOR2_X1 U1202 ( .A(n480), .B(n465), .ZN(n1328) );
  XNOR2_X1 U1203 ( .A(n1566), .B(a[14]), .ZN(n1329) );
  INV_X1 U1204 ( .A(n1244), .ZN(n1330) );
  INV_X1 U1205 ( .A(n1243), .ZN(n1331) );
  NOR2_X1 U1206 ( .A1(n581), .A2(n590), .ZN(n1332) );
  CLKBUF_X1 U1207 ( .A(n1462), .Z(n1389) );
  NAND3_X1 U1208 ( .A1(n1463), .A2(n1462), .A3(n1461), .ZN(n1334) );
  CLKBUF_X1 U1209 ( .A(n1268), .Z(n1335) );
  NAND3_X1 U1210 ( .A1(n1327), .A2(n1335), .A3(n1465), .ZN(n1336) );
  BUF_X1 U1211 ( .A(n1586), .Z(n1338) );
  BUF_X2 U1212 ( .A(n1586), .Z(n1339) );
  XNOR2_X1 U1213 ( .A(n1355), .B(n1470), .ZN(n1340) );
  CLKBUF_X1 U1214 ( .A(n1396), .Z(n1341) );
  CLKBUF_X1 U1215 ( .A(n1518), .Z(n1342) );
  BUF_X2 U1216 ( .A(n1518), .Z(n1343) );
  CLKBUF_X1 U1217 ( .A(n1518), .Z(n1344) );
  XNOR2_X1 U1218 ( .A(n13), .B(a[6]), .ZN(n1518) );
  BUF_X1 U1219 ( .A(n1097), .Z(n1345) );
  XNOR2_X2 U1220 ( .A(n1565), .B(a[12]), .ZN(n1545) );
  NAND3_X1 U1221 ( .A1(n1395), .A2(n1396), .A3(n1397), .ZN(n1346) );
  NAND3_X1 U1222 ( .A1(n1395), .A2(n1341), .A3(n1397), .ZN(n1347) );
  BUF_X2 U1223 ( .A(n24), .Z(n1349) );
  NAND2_X1 U1224 ( .A1(n1116), .A2(n1518), .ZN(n24) );
  BUF_X2 U1225 ( .A(n9), .Z(n1533) );
  NAND2_X1 U1226 ( .A1(n1516), .A2(n1270), .ZN(n1501) );
  NAND2_X1 U1227 ( .A1(n1516), .A2(n1270), .ZN(n1502) );
  BUF_X1 U1228 ( .A(n1376), .Z(n1350) );
  CLKBUF_X1 U1229 ( .A(n1573), .Z(n1351) );
  CLKBUF_X1 U1230 ( .A(n1573), .Z(n1352) );
  XNOR2_X1 U1231 ( .A(n1568), .B(a[18]), .ZN(n1353) );
  BUF_X2 U1232 ( .A(n49), .Z(n1568) );
  OAI22_X1 U1233 ( .A1(n1486), .A2(n954), .B1(n953), .B2(n1545), .ZN(n1354) );
  BUF_X2 U1234 ( .A(n1589), .Z(n1355) );
  CLKBUF_X1 U1235 ( .A(n61), .Z(n1356) );
  XNOR2_X1 U1236 ( .A(n1376), .B(n1470), .ZN(n1357) );
  CLKBUF_X2 U1237 ( .A(n7), .Z(n1359) );
  XNOR2_X1 U1238 ( .A(n552), .B(n1360), .ZN(n535) );
  XNOR2_X1 U1239 ( .A(n550), .B(n554), .ZN(n1360) );
  OAI22_X1 U1240 ( .A1(n1239), .A2(n1013), .B1(n1012), .B2(n1343), .ZN(n1361)
         );
  BUF_X1 U1241 ( .A(n1098), .Z(n1362) );
  CLKBUF_X1 U1242 ( .A(n54), .Z(n1364) );
  CLKBUF_X1 U1243 ( .A(n1575), .Z(n1365) );
  INV_X1 U1244 ( .A(n668), .ZN(n1368) );
  INV_X2 U1245 ( .A(n1241), .ZN(n4) );
  BUF_X1 U1246 ( .A(n1101), .Z(n1369) );
  CLKBUF_X1 U1247 ( .A(n1509), .Z(n1384) );
  BUF_X4 U1248 ( .A(n19), .Z(n1509) );
  CLKBUF_X1 U1249 ( .A(n1587), .Z(n1371) );
  AOI21_X1 U1250 ( .B1(n1547), .B2(n1548), .A(n1557), .ZN(n1372) );
  CLKBUF_X1 U1251 ( .A(n13), .Z(n1373) );
  INV_X1 U1252 ( .A(n1588), .ZN(n1374) );
  INV_X1 U1253 ( .A(n1374), .ZN(n1375) );
  BUF_X2 U1254 ( .A(n1091), .Z(n1588) );
  BUF_X2 U1255 ( .A(n1585), .Z(n1377) );
  CLKBUF_X1 U1256 ( .A(n1584), .Z(n1381) );
  BUF_X1 U1257 ( .A(n1103), .Z(n1382) );
  XNOR2_X1 U1258 ( .A(n1386), .B(n532), .ZN(n515) );
  XNOR2_X1 U1259 ( .A(n519), .B(n521), .ZN(n1386) );
  BUF_X4 U1260 ( .A(n37), .Z(n1387) );
  INV_X1 U1261 ( .A(n1529), .ZN(n1388) );
  CLKBUF_X1 U1262 ( .A(n264), .Z(n1390) );
  NAND2_X1 U1263 ( .A1(n499), .A2(n514), .ZN(n1391) );
  NAND2_X1 U1264 ( .A1(n499), .A2(n501), .ZN(n1392) );
  NAND2_X1 U1265 ( .A1(n514), .A2(n501), .ZN(n1393) );
  NAND3_X1 U1266 ( .A1(n1391), .A2(n1392), .A3(n1393), .ZN(n496) );
  XOR2_X1 U1267 ( .A(n310), .B(n307), .Z(n1394) );
  XOR2_X1 U1268 ( .A(n1390), .B(n1394), .Z(product[34]) );
  NAND2_X1 U1269 ( .A1(n264), .A2(n310), .ZN(n1395) );
  NAND2_X1 U1270 ( .A1(n264), .A2(n307), .ZN(n1396) );
  NAND2_X1 U1271 ( .A1(n310), .A2(n307), .ZN(n1397) );
  NAND3_X1 U1272 ( .A1(n1395), .A2(n1396), .A3(n1397), .ZN(n100) );
  NAND3_X1 U1273 ( .A1(n1463), .A2(n1462), .A3(n1461), .ZN(n1398) );
  XOR2_X1 U1274 ( .A(n1565), .B(a[12]), .Z(n1399) );
  NAND3_X1 U1275 ( .A1(n1467), .A2(n1466), .A3(n1465), .ZN(n1401) );
  XNOR2_X1 U1276 ( .A(n1469), .B(n1402), .ZN(product[38]) );
  NAND3_X1 U1277 ( .A1(n1269), .A2(n1477), .A3(n1479), .ZN(n1402) );
  AND3_X1 U1278 ( .A1(n1482), .A2(n1481), .A3(n1480), .ZN(product[39]) );
  INV_X1 U1279 ( .A(n1544), .ZN(n1404) );
  INV_X1 U1280 ( .A(n1404), .ZN(n1405) );
  XOR2_X1 U1281 ( .A(n811), .B(n829), .Z(n1406) );
  XOR2_X1 U1282 ( .A(n578), .B(n1406), .Z(n563) );
  NAND2_X1 U1283 ( .A1(n578), .A2(n811), .ZN(n1407) );
  NAND2_X1 U1284 ( .A1(n578), .A2(n829), .ZN(n1408) );
  NAND2_X1 U1285 ( .A1(n811), .A2(n829), .ZN(n1409) );
  NAND3_X1 U1286 ( .A1(n1407), .A2(n1408), .A3(n1409), .ZN(n562) );
  XOR2_X1 U1287 ( .A(n547), .B(n558), .Z(n1410) );
  XOR2_X1 U1288 ( .A(n1410), .B(n545), .Z(n543) );
  NAND2_X1 U1289 ( .A1(n560), .A2(n553), .ZN(n1411) );
  NAND2_X1 U1290 ( .A1(n560), .A2(n549), .ZN(n1412) );
  NAND2_X1 U1291 ( .A1(n553), .A2(n549), .ZN(n1413) );
  NAND3_X1 U1292 ( .A1(n1411), .A2(n1412), .A3(n1413), .ZN(n544) );
  NAND2_X1 U1293 ( .A1(n547), .A2(n558), .ZN(n1414) );
  NAND2_X1 U1294 ( .A1(n547), .A2(n545), .ZN(n1415) );
  NAND2_X1 U1295 ( .A1(n558), .A2(n545), .ZN(n1416) );
  NAND3_X1 U1296 ( .A1(n1414), .A2(n1415), .A3(n1416), .ZN(n542) );
  NOR2_X2 U1297 ( .A1(n371), .A2(n382), .ZN(n135) );
  CLKBUF_X1 U1298 ( .A(n172), .Z(n1417) );
  XOR2_X1 U1299 ( .A(n861), .B(n752), .Z(n1418) );
  XOR2_X1 U1300 ( .A(n1422), .B(n1418), .Z(n491) );
  NAND2_X1 U1301 ( .A1(n1361), .A2(n752), .ZN(n1419) );
  NAND2_X1 U1302 ( .A1(n861), .A2(n806), .ZN(n1420) );
  NAND2_X1 U1303 ( .A1(n1236), .A2(n861), .ZN(n1421) );
  NAND3_X1 U1304 ( .A1(n1419), .A2(n1421), .A3(n1420), .ZN(n490) );
  CLKBUF_X1 U1305 ( .A(n1361), .Z(n1422) );
  XOR2_X1 U1306 ( .A(n588), .B(n579), .Z(n1423) );
  XOR2_X1 U1307 ( .A(n586), .B(n1423), .Z(n573) );
  NAND2_X1 U1308 ( .A1(n586), .A2(n588), .ZN(n1424) );
  NAND2_X1 U1309 ( .A1(n586), .A2(n579), .ZN(n1425) );
  NAND2_X1 U1310 ( .A1(n588), .A2(n579), .ZN(n1426) );
  NAND3_X1 U1311 ( .A1(n1424), .A2(n1425), .A3(n1426), .ZN(n572) );
  XOR2_X1 U1312 ( .A(n813), .B(n849), .Z(n1427) );
  XOR2_X1 U1313 ( .A(n777), .B(n1427), .Z(n587) );
  NAND2_X1 U1314 ( .A1(n777), .A2(n813), .ZN(n1428) );
  NAND2_X1 U1315 ( .A1(n777), .A2(n849), .ZN(n1429) );
  NAND2_X1 U1316 ( .A1(n813), .A2(n849), .ZN(n1430) );
  NAND3_X1 U1317 ( .A1(n1428), .A2(n1429), .A3(n1430), .ZN(n586) );
  NAND2_X1 U1318 ( .A1(n1354), .A2(n822), .ZN(n1431) );
  NAND2_X1 U1319 ( .A1(n750), .A2(n696), .ZN(n1432) );
  NAND2_X1 U1320 ( .A1(n822), .A2(n696), .ZN(n1433) );
  NAND3_X1 U1321 ( .A1(n1431), .A2(n1432), .A3(n1433), .ZN(n456) );
  INV_X1 U1322 ( .A(n1529), .ZN(n1558) );
  CLKBUF_X1 U1323 ( .A(n161), .Z(n1434) );
  INV_X1 U1324 ( .A(n1530), .ZN(n1435) );
  CLKBUF_X1 U1325 ( .A(n60), .Z(n1436) );
  XNOR2_X1 U1326 ( .A(n429), .B(n1437), .ZN(n427) );
  XNOR2_X1 U1327 ( .A(n444), .B(n431), .ZN(n1437) );
  NAND2_X1 U1328 ( .A1(n429), .A2(n444), .ZN(n1438) );
  NAND2_X1 U1329 ( .A1(n429), .A2(n431), .ZN(n1439) );
  NAND2_X1 U1330 ( .A1(n444), .A2(n431), .ZN(n1440) );
  NAND3_X1 U1331 ( .A1(n1438), .A2(n1439), .A3(n1440), .ZN(n426) );
  CLKBUF_X1 U1332 ( .A(n194), .Z(n1441) );
  NAND2_X1 U1333 ( .A1(n735), .A2(n699), .ZN(n1442) );
  NAND2_X1 U1334 ( .A1(n735), .A2(n862), .ZN(n1443) );
  NAND2_X1 U1335 ( .A1(n699), .A2(n862), .ZN(n1444) );
  NAND3_X1 U1336 ( .A1(n1442), .A2(n1443), .A3(n1444), .ZN(n510) );
  NAND2_X1 U1337 ( .A1(n463), .A2(n480), .ZN(n1445) );
  NAND2_X1 U1338 ( .A1(n463), .A2(n1242), .ZN(n1446) );
  NAND2_X1 U1339 ( .A1(n480), .A2(n1242), .ZN(n1447) );
  NAND3_X1 U1340 ( .A1(n1445), .A2(n1446), .A3(n1447), .ZN(n460) );
  OR2_X1 U1341 ( .A1(n1388), .A2(n938), .ZN(n1448) );
  OR2_X1 U1342 ( .A1(n937), .A2(n1540), .ZN(n1449) );
  NAND2_X1 U1343 ( .A1(n1448), .A2(n1449), .ZN(n735) );
  NAND2_X1 U1344 ( .A1(n552), .A2(n554), .ZN(n1450) );
  NAND2_X1 U1345 ( .A1(n552), .A2(n550), .ZN(n1451) );
  NAND2_X1 U1346 ( .A1(n554), .A2(n550), .ZN(n1452) );
  NAND3_X1 U1347 ( .A1(n1450), .A2(n1451), .A3(n1452), .ZN(n534) );
  XNOR2_X1 U1348 ( .A(n1453), .B(n515), .ZN(n513) );
  XNOR2_X1 U1349 ( .A(n517), .B(n530), .ZN(n1453) );
  NOR2_X1 U1350 ( .A1(n443), .A2(n460), .ZN(n161) );
  NAND2_X1 U1351 ( .A1(n519), .A2(n521), .ZN(n1454) );
  NAND2_X1 U1352 ( .A1(n519), .A2(n532), .ZN(n1455) );
  NAND2_X1 U1353 ( .A1(n521), .A2(n532), .ZN(n1456) );
  NAND2_X1 U1354 ( .A1(n517), .A2(n530), .ZN(n1457) );
  NAND2_X1 U1355 ( .A1(n517), .A2(n515), .ZN(n1458) );
  NAND2_X1 U1356 ( .A1(n530), .A2(n515), .ZN(n1459) );
  NAND3_X1 U1357 ( .A1(n1457), .A2(n1458), .A3(n1459), .ZN(n512) );
  BUF_X2 U1358 ( .A(n1313), .Z(n1543) );
  XOR2_X1 U1359 ( .A(n303), .B(n306), .Z(n1460) );
  XOR2_X1 U1360 ( .A(n1460), .B(n1347), .Z(product[35]) );
  NAND2_X1 U1361 ( .A1(n303), .A2(n306), .ZN(n1461) );
  NAND2_X1 U1362 ( .A1(n100), .A2(n303), .ZN(n1462) );
  NAND2_X1 U1363 ( .A1(n306), .A2(n1346), .ZN(n1463) );
  NAND3_X1 U1364 ( .A1(n1311), .A2(n1389), .A3(n1461), .ZN(n99) );
  XOR2_X1 U1365 ( .A(n302), .B(n301), .Z(n1464) );
  XOR2_X1 U1366 ( .A(n1464), .B(n99), .Z(product[36]) );
  NAND2_X1 U1367 ( .A1(n302), .A2(n301), .ZN(n1465) );
  NAND2_X1 U1368 ( .A1(n1398), .A2(n302), .ZN(n1466) );
  NAND2_X1 U1369 ( .A1(n301), .A2(n1334), .ZN(n1467) );
  NAND3_X1 U1370 ( .A1(n1467), .A2(n1268), .A3(n1465), .ZN(n98) );
  CLKBUF_X1 U1371 ( .A(n162), .Z(n1468) );
  XNOR2_X1 U1372 ( .A(n680), .B(n298), .ZN(n1469) );
  INV_X1 U1373 ( .A(n1530), .ZN(n1563) );
  CLKBUF_X1 U1374 ( .A(n127), .Z(n1472) );
  NAND3_X1 U1375 ( .A1(n1269), .A2(n1479), .A3(n1477), .ZN(n1473) );
  CLKBUF_X1 U1376 ( .A(n106), .Z(n1474) );
  CLKBUF_X1 U1377 ( .A(n114), .Z(n1475) );
  XOR2_X1 U1378 ( .A(n300), .B(n299), .Z(n1476) );
  XOR2_X1 U1379 ( .A(n1476), .B(n1336), .Z(product[37]) );
  NAND2_X1 U1380 ( .A1(n300), .A2(n299), .ZN(n1477) );
  NAND2_X1 U1381 ( .A1(n98), .A2(n300), .ZN(n1478) );
  NAND2_X1 U1382 ( .A1(n299), .A2(n1401), .ZN(n1479) );
  NAND3_X1 U1383 ( .A1(n1479), .A2(n1478), .A3(n1477), .ZN(n97) );
  NAND2_X1 U1384 ( .A1(n680), .A2(n298), .ZN(n1480) );
  NAND2_X1 U1385 ( .A1(n97), .A2(n680), .ZN(n1481) );
  NAND2_X1 U1386 ( .A1(n1473), .A2(n298), .ZN(n1482) );
  INV_X1 U1387 ( .A(n1531), .ZN(n1551) );
  INV_X1 U1388 ( .A(n1529), .ZN(n1559) );
  CLKBUF_X1 U1389 ( .A(n151), .Z(n1483) );
  XNOR2_X1 U1390 ( .A(n1566), .B(a[12]), .ZN(n1484) );
  OR2_X2 U1391 ( .A1(n1484), .A2(n1399), .ZN(n1485) );
  CLKBUF_X1 U1392 ( .A(n146), .Z(n1487) );
  AOI21_X1 U1393 ( .B1(n1487), .B2(n133), .A(n1306), .ZN(n1488) );
  BUF_X4 U1394 ( .A(n49), .Z(n1489) );
  CLKBUF_X1 U1395 ( .A(n1436), .Z(n1490) );
  AOI21_X1 U1396 ( .B1(n175), .B2(n1441), .A(n1321), .ZN(n1491) );
  NAND2_X1 U1397 ( .A1(n16), .A2(n1515), .ZN(n18) );
  AOI21_X1 U1398 ( .B1(n114), .B2(n1525), .A(n111), .ZN(n1493) );
  CLKBUF_X1 U1399 ( .A(n1541), .Z(n1494) );
  CLKBUF_X1 U1400 ( .A(n122), .Z(n1497) );
  CLKBUF_X2 U1401 ( .A(n52), .Z(n1499) );
  AOI21_X1 U1402 ( .B1(n122), .B2(n1524), .A(n119), .ZN(n1500) );
  NAND2_X1 U1403 ( .A1(n1516), .A2(n1270), .ZN(n12) );
  BUF_X1 U1404 ( .A(n58), .Z(n1504) );
  NOR2_X1 U1405 ( .A1(n427), .A2(n442), .ZN(n1503) );
  NOR2_X1 U1406 ( .A1(n461), .A2(n478), .ZN(n1507) );
  BUF_X4 U1407 ( .A(n43), .Z(n1567) );
  CLKBUF_X1 U1408 ( .A(n153), .Z(n1508) );
  OR2_X1 U1409 ( .A1(n679), .A2(n879), .ZN(n1510) );
  NAND2_X2 U1410 ( .A1(n58), .A2(n1511), .ZN(n60) );
  XOR2_X1 U1411 ( .A(n55), .B(a[18]), .Z(n1511) );
  NAND2_X2 U1412 ( .A1(n1512), .A2(n52), .ZN(n54) );
  XOR2_X1 U1413 ( .A(n1568), .B(a[16]), .Z(n1512) );
  XOR2_X1 U1414 ( .A(n1565), .B(a[10]), .Z(n1513) );
  XOR2_X1 U1415 ( .A(n43), .B(a[14]), .Z(n1514) );
  BUF_X1 U1416 ( .A(n61), .Z(n1571) );
  XNOR2_X1 U1417 ( .A(n19), .B(a[8]), .ZN(n28) );
  XOR2_X1 U1418 ( .A(n13), .B(a[4]), .Z(n1515) );
  XOR2_X1 U1419 ( .A(a[2]), .B(n7), .Z(n1516) );
  AOI21_X1 U1420 ( .B1(n153), .B2(n126), .A(n127), .ZN(n1517) );
  OAI21_X1 U1421 ( .B1(n152), .B2(n1251), .A(n144), .ZN(n142) );
  INV_X1 U1422 ( .A(n1487), .ZN(n144) );
  AOI21_X1 U1423 ( .B1(n146), .B2(n133), .A(n134), .ZN(n132) );
  NAND2_X1 U1424 ( .A1(n268), .A2(n116), .ZN(n66) );
  INV_X1 U1425 ( .A(n115), .ZN(n268) );
  INV_X1 U1426 ( .A(n1316), .ZN(n279) );
  XOR2_X1 U1427 ( .A(n137), .B(n70), .Z(product[26]) );
  NAND2_X1 U1428 ( .A1(n272), .A2(n136), .ZN(n70) );
  AOI21_X1 U1429 ( .B1(n142), .B2(n273), .A(n139), .ZN(n137) );
  INV_X1 U1430 ( .A(n135), .ZN(n272) );
  XOR2_X1 U1431 ( .A(n206), .B(n82), .Z(product[14]) );
  NAND2_X1 U1432 ( .A1(n284), .A2(n205), .ZN(n82) );
  AOI21_X1 U1433 ( .B1(n211), .B2(n285), .A(n208), .ZN(n206) );
  XOR2_X1 U1434 ( .A(n168), .B(n76), .Z(product[20]) );
  NAND2_X1 U1435 ( .A1(n278), .A2(n167), .ZN(n76) );
  AOI21_X1 U1436 ( .B1(n173), .B2(n279), .A(n170), .ZN(n168) );
  XOR2_X1 U1437 ( .A(n163), .B(n75), .Z(product[21]) );
  NAND2_X1 U1438 ( .A1(n277), .A2(n1468), .ZN(n75) );
  XOR2_X1 U1439 ( .A(n193), .B(n80), .Z(product[16]) );
  NAND2_X1 U1440 ( .A1(n1312), .A2(n188), .ZN(n80) );
  XOR2_X1 U1441 ( .A(n152), .B(n73), .Z(product[23]) );
  INV_X1 U1442 ( .A(n221), .ZN(n220) );
  XNOR2_X1 U1443 ( .A(n160), .B(n74), .ZN(product[22]) );
  NAND2_X1 U1444 ( .A1(n276), .A2(n159), .ZN(n74) );
  XNOR2_X1 U1445 ( .A(n173), .B(n77), .ZN(product[19]) );
  NAND2_X1 U1446 ( .A1(n279), .A2(n1417), .ZN(n77) );
  XNOR2_X1 U1447 ( .A(n149), .B(n72), .ZN(product[24]) );
  NAND2_X1 U1448 ( .A1(n274), .A2(n148), .ZN(n72) );
  XNOR2_X1 U1449 ( .A(n130), .B(n69), .ZN(product[27]) );
  NAND2_X1 U1450 ( .A1(n271), .A2(n129), .ZN(n69) );
  INV_X1 U1451 ( .A(n128), .ZN(n271) );
  XNOR2_X1 U1452 ( .A(n142), .B(n71), .ZN(product[25]) );
  XNOR2_X1 U1453 ( .A(n179), .B(n78), .ZN(product[18]) );
  NAND2_X1 U1454 ( .A1(n280), .A2(n178), .ZN(n78) );
  INV_X1 U1455 ( .A(n1250), .ZN(n273) );
  INV_X1 U1456 ( .A(n1417), .ZN(n170) );
  NAND2_X1 U1457 ( .A1(n1520), .A2(n1519), .ZN(n222) );
  AOI21_X1 U1458 ( .B1(n1520), .B2(n230), .A(n225), .ZN(n223) );
  INV_X1 U1459 ( .A(n121), .ZN(n119) );
  INV_X1 U1460 ( .A(n113), .ZN(n111) );
  INV_X1 U1461 ( .A(n200), .ZN(n198) );
  AOI21_X1 U1462 ( .B1(n221), .B2(n213), .A(n214), .ZN(n212) );
  NOR2_X1 U1463 ( .A1(n461), .A2(n478), .ZN(n166) );
  NOR2_X1 U1464 ( .A1(n427), .A2(n442), .ZN(n158) );
  NAND2_X1 U1465 ( .A1(n266), .A2(n108), .ZN(n64) );
  INV_X1 U1466 ( .A(n107), .ZN(n266) );
  NAND2_X1 U1467 ( .A1(n270), .A2(n124), .ZN(n68) );
  INV_X1 U1468 ( .A(n123), .ZN(n270) );
  INV_X1 U1469 ( .A(n232), .ZN(n230) );
  NAND2_X1 U1470 ( .A1(n443), .A2(n460), .ZN(n162) );
  NOR2_X1 U1471 ( .A1(n359), .A2(n370), .ZN(n128) );
  INV_X1 U1472 ( .A(n209), .ZN(n285) );
  NAND2_X1 U1473 ( .A1(n1525), .A2(n113), .ZN(n65) );
  NAND2_X1 U1474 ( .A1(n1523), .A2(n105), .ZN(n63) );
  NAND2_X1 U1475 ( .A1(n1524), .A2(n121), .ZN(n67) );
  XOR2_X1 U1476 ( .A(n220), .B(n85), .Z(product[11]) );
  NAND2_X1 U1477 ( .A1(n287), .A2(n219), .ZN(n85) );
  INV_X1 U1478 ( .A(n218), .ZN(n287) );
  XOR2_X1 U1479 ( .A(n228), .B(n86), .Z(product[10]) );
  NAND2_X1 U1480 ( .A1(n1520), .A2(n227), .ZN(n86) );
  AOI21_X1 U1481 ( .B1(n233), .B2(n1519), .A(n230), .ZN(n228) );
  XOR2_X1 U1482 ( .A(n201), .B(n81), .Z(product[15]) );
  AOI21_X1 U1483 ( .B1(n211), .B2(n202), .A(n203), .ZN(n201) );
  NOR2_X1 U1484 ( .A1(n479), .A2(n496), .ZN(n171) );
  NAND2_X1 U1485 ( .A1(n557), .A2(n568), .ZN(n205) );
  NAND2_X1 U1486 ( .A1(n371), .A2(n382), .ZN(n136) );
  NOR2_X1 U1487 ( .A1(n331), .A2(n338), .ZN(n115) );
  XNOR2_X1 U1488 ( .A(n239), .B(n88), .ZN(product[8]) );
  NAND2_X1 U1489 ( .A1(n1522), .A2(n238), .ZN(n88) );
  NAND2_X1 U1490 ( .A1(n479), .A2(n496), .ZN(n172) );
  XNOR2_X1 U1491 ( .A(n211), .B(n83), .ZN(product[13]) );
  NAND2_X1 U1492 ( .A1(n285), .A2(n210), .ZN(n83) );
  XNOR2_X1 U1493 ( .A(n186), .B(n79), .ZN(product[17]) );
  INV_X1 U1494 ( .A(n1557), .ZN(n185) );
  XNOR2_X1 U1495 ( .A(n233), .B(n87), .ZN(product[9]) );
  NAND2_X1 U1496 ( .A1(n1519), .A2(n232), .ZN(n87) );
  XNOR2_X1 U1497 ( .A(n217), .B(n84), .ZN(product[12]) );
  NAND2_X1 U1498 ( .A1(n286), .A2(n216), .ZN(n84) );
  OAI21_X1 U1499 ( .B1(n220), .B2(n218), .A(n219), .ZN(n217) );
  NAND2_X1 U1500 ( .A1(n497), .A2(n512), .ZN(n178) );
  NAND2_X1 U1501 ( .A1(n359), .A2(n370), .ZN(n129) );
  NAND2_X1 U1502 ( .A1(n331), .A2(n338), .ZN(n116) );
  INV_X1 U1503 ( .A(n210), .ZN(n208) );
  INV_X1 U1504 ( .A(n227), .ZN(n225) );
  INV_X1 U1505 ( .A(n1548), .ZN(n188) );
  INV_X1 U1506 ( .A(n238), .ZN(n236) );
  INV_X1 U1507 ( .A(n246), .ZN(n244) );
  OR2_X1 U1508 ( .A1(n609), .A2(n616), .ZN(n1519) );
  OR2_X1 U1509 ( .A1(n601), .A2(n608), .ZN(n1520) );
  OAI21_X1 U1510 ( .B1(n256), .B2(n258), .A(n257), .ZN(n255) );
  NOR2_X1 U1511 ( .A1(n591), .A2(n600), .ZN(n218) );
  AOI21_X1 U1512 ( .B1(n1527), .B2(n255), .A(n252), .ZN(n250) );
  INV_X1 U1513 ( .A(n254), .ZN(n252) );
  NAND2_X1 U1514 ( .A1(n291), .A2(n241), .ZN(n89) );
  INV_X1 U1515 ( .A(n240), .ZN(n291) );
  OR2_X1 U1516 ( .A1(n543), .A2(n556), .ZN(n1521) );
  NAND2_X1 U1517 ( .A1(n1528), .A2(n246), .ZN(n90) );
  XOR2_X1 U1518 ( .A(n91), .B(n250), .Z(product[5]) );
  NAND2_X1 U1519 ( .A1(n293), .A2(n249), .ZN(n91) );
  NAND2_X1 U1520 ( .A1(n591), .A2(n600), .ZN(n219) );
  NOR2_X1 U1521 ( .A1(n569), .A2(n580), .ZN(n209) );
  NOR2_X1 U1522 ( .A1(n317), .A2(n322), .ZN(n107) );
  NOR2_X1 U1523 ( .A1(n349), .A2(n358), .ZN(n123) );
  INV_X1 U1524 ( .A(n259), .ZN(n258) );
  OAI21_X1 U1525 ( .B1(n260), .B2(n263), .A(n261), .ZN(n259) );
  NAND2_X1 U1526 ( .A1(n569), .A2(n580), .ZN(n210) );
  OR2_X1 U1527 ( .A1(n617), .A2(n622), .ZN(n1522) );
  XNOR2_X1 U1528 ( .A(n92), .B(n255), .ZN(product[4]) );
  NAND2_X1 U1529 ( .A1(n1527), .A2(n254), .ZN(n92) );
  OR2_X1 U1530 ( .A1(n311), .A2(n316), .ZN(n1523) );
  NAND2_X1 U1531 ( .A1(n617), .A2(n622), .ZN(n238) );
  NAND2_X1 U1532 ( .A1(n311), .A2(n316), .ZN(n105) );
  NAND2_X1 U1533 ( .A1(n339), .A2(n348), .ZN(n121) );
  NAND2_X1 U1534 ( .A1(n323), .A2(n330), .ZN(n113) );
  NAND2_X1 U1535 ( .A1(n317), .A2(n322), .ZN(n108) );
  NAND2_X1 U1536 ( .A1(n349), .A2(n358), .ZN(n124) );
  NAND2_X1 U1537 ( .A1(n601), .A2(n608), .ZN(n227) );
  OR2_X1 U1538 ( .A1(n339), .A2(n348), .ZN(n1524) );
  OR2_X1 U1539 ( .A1(n323), .A2(n330), .ZN(n1525) );
  NAND2_X1 U1540 ( .A1(n581), .A2(n590), .ZN(n216) );
  XOR2_X1 U1541 ( .A(n93), .B(n258), .Z(product[3]) );
  NAND2_X1 U1542 ( .A1(n295), .A2(n257), .ZN(n93) );
  INV_X1 U1543 ( .A(n256), .ZN(n295) );
  NAND2_X1 U1544 ( .A1(n543), .A2(n556), .ZN(n200) );
  XOR2_X1 U1545 ( .A(n94), .B(n263), .Z(product[2]) );
  NAND2_X1 U1546 ( .A1(n296), .A2(n261), .ZN(n94) );
  INV_X1 U1547 ( .A(n260), .ZN(n296) );
  NOR2_X1 U1548 ( .A1(n639), .A2(n678), .ZN(n256) );
  XNOR2_X1 U1549 ( .A(n815), .B(n1526), .ZN(n607) );
  XNOR2_X1 U1550 ( .A(n870), .B(n779), .ZN(n1526) );
  NOR2_X1 U1551 ( .A1(n878), .A2(n859), .ZN(n260) );
  NAND2_X1 U1552 ( .A1(n679), .A2(n879), .ZN(n263) );
  NAND2_X1 U1553 ( .A1(n878), .A2(n859), .ZN(n261) );
  OR2_X1 U1554 ( .A1(n637), .A2(n638), .ZN(n1527) );
  INV_X1 U1555 ( .A(n394), .ZN(n395) );
  INV_X1 U1556 ( .A(n328), .ZN(n329) );
  INV_X1 U1557 ( .A(n346), .ZN(n347) );
  NOR2_X1 U1558 ( .A1(n623), .A2(n628), .ZN(n240) );
  INV_X1 U1559 ( .A(n105), .ZN(n103) );
  INV_X1 U1560 ( .A(n298), .ZN(n299) );
  NAND2_X1 U1561 ( .A1(n629), .A2(n632), .ZN(n246) );
  NAND2_X1 U1562 ( .A1(n623), .A2(n628), .ZN(n241) );
  OR2_X1 U1563 ( .A1(n629), .A2(n632), .ZN(n1528) );
  NAND2_X1 U1564 ( .A1(n633), .A2(n636), .ZN(n249) );
  OAI22_X1 U1565 ( .A1(n1535), .A2(n1088), .B1(n1087), .B2(n4), .ZN(n879) );
  OAI22_X1 U1566 ( .A1(n1536), .A2(n1149), .B1(n1089), .B2(n4), .ZN(n679) );
  OR2_X1 U1567 ( .A1(n1571), .A2(n1149), .ZN(n1089) );
  OAI22_X1 U1568 ( .A1(n1535), .A2(n1087), .B1(n1086), .B2(n4), .ZN(n878) );
  OR2_X1 U1569 ( .A1(n61), .A2(n1148), .ZN(n1068) );
  OAI22_X1 U1570 ( .A1(n1534), .A2(n1070), .B1(n1340), .B2(n4), .ZN(n861) );
  AND2_X1 U1571 ( .A1(n1571), .A2(n1404), .ZN(n759) );
  OAI22_X1 U1572 ( .A1(n1536), .A2(n1077), .B1(n1076), .B2(n4), .ZN(n868) );
  INV_X1 U1573 ( .A(n667), .ZN(n860) );
  OAI22_X1 U1574 ( .A1(n1536), .A2(n1082), .B1(n1081), .B2(n4), .ZN(n873) );
  OAI22_X1 U1575 ( .A1(n1069), .A2(n1534), .B1(n1357), .B2(n4), .ZN(n667) );
  BUF_X1 U1576 ( .A(n6), .Z(n1535) );
  AND2_X1 U1577 ( .A1(n1356), .A2(n662), .ZN(n839) );
  OAI22_X1 U1578 ( .A1(n1535), .A2(n1085), .B1(n1084), .B2(n4), .ZN(n876) );
  OAI22_X1 U1579 ( .A1(n1536), .A2(n1084), .B1(n1083), .B2(n4), .ZN(n875) );
  OR2_X1 U1580 ( .A1(n1571), .A2(n1147), .ZN(n1047) );
  XNOR2_X1 U1581 ( .A(n1285), .B(n1569), .ZN(n889) );
  XNOR2_X1 U1582 ( .A(n1581), .B(n1569), .ZN(n888) );
  XNOR2_X1 U1583 ( .A(n1345), .B(n1287), .ZN(n887) );
  XNOR2_X1 U1584 ( .A(n1574), .B(n1569), .ZN(n896) );
  XNOR2_X1 U1585 ( .A(n1573), .B(n1569), .ZN(n897) );
  XNOR2_X1 U1586 ( .A(n1572), .B(n1569), .ZN(n898) );
  XNOR2_X1 U1587 ( .A(n1365), .B(n1569), .ZN(n895) );
  XNOR2_X1 U1588 ( .A(n1576), .B(n1569), .ZN(n894) );
  XNOR2_X1 U1589 ( .A(n1319), .B(n1569), .ZN(n893) );
  XNOR2_X1 U1590 ( .A(n1322), .B(n1569), .ZN(n892) );
  XNOR2_X1 U1591 ( .A(n1369), .B(n1569), .ZN(n891) );
  XNOR2_X1 U1592 ( .A(n1579), .B(n1569), .ZN(n890) );
  XNOR2_X1 U1593 ( .A(n1583), .B(n1287), .ZN(n886) );
  XNOR2_X1 U1594 ( .A(n1381), .B(n1287), .ZN(n885) );
  XNOR2_X1 U1595 ( .A(n1377), .B(n1287), .ZN(n884) );
  XNOR2_X1 U1596 ( .A(n1338), .B(n1287), .ZN(n883) );
  XNOR2_X1 U1597 ( .A(n1371), .B(n1287), .ZN(n882) );
  XNOR2_X1 U1598 ( .A(n1375), .B(n1287), .ZN(n881) );
  AND2_X1 U1599 ( .A1(n1356), .A2(n665), .ZN(n859) );
  BUF_X1 U1600 ( .A(n1090), .Z(n1589) );
  BUF_X1 U1601 ( .A(n1094), .Z(n1585) );
  BUF_X1 U1602 ( .A(n1105), .Z(n1575) );
  BUF_X1 U1603 ( .A(n1103), .Z(n1577) );
  BUF_X1 U1604 ( .A(n1097), .Z(n1582) );
  BUF_X1 U1605 ( .A(n1102), .Z(n1578) );
  BUF_X1 U1606 ( .A(n1098), .Z(n1581) );
  BUF_X1 U1607 ( .A(n1093), .Z(n1586) );
  INV_X1 U1608 ( .A(n655), .ZN(n780) );
  INV_X1 U1609 ( .A(n314), .ZN(n315) );
  INV_X1 U1610 ( .A(n304), .ZN(n305) );
  AND2_X1 U1611 ( .A1(n1356), .A2(n641), .ZN(n699) );
  OAI22_X1 U1612 ( .A1(n1534), .A2(n1071), .B1(n1070), .B2(n4), .ZN(n862) );
  OAI22_X1 U1613 ( .A1(n1536), .A2(n1072), .B1(n1071), .B2(n4), .ZN(n863) );
  OAI22_X1 U1614 ( .A1(n1535), .A2(n1076), .B1(n1075), .B2(n4), .ZN(n867) );
  INV_X1 U1615 ( .A(n649), .ZN(n740) );
  INV_X1 U1616 ( .A(n643), .ZN(n700) );
  INV_X1 U1617 ( .A(n458), .ZN(n459) );
  INV_X1 U1618 ( .A(n658), .ZN(n800) );
  INV_X1 U1619 ( .A(n652), .ZN(n760) );
  INV_X1 U1620 ( .A(n646), .ZN(n720) );
  OAI22_X1 U1621 ( .A1(n1535), .A2(n1080), .B1(n1079), .B2(n4), .ZN(n871) );
  INV_X1 U1622 ( .A(n424), .ZN(n425) );
  AND2_X1 U1623 ( .A1(n1571), .A2(n647), .ZN(n739) );
  OAI22_X1 U1624 ( .A1(n1535), .A2(n1075), .B1(n1074), .B2(n4), .ZN(n866) );
  AND2_X1 U1625 ( .A1(n1571), .A2(n659), .ZN(n819) );
  OAI22_X1 U1626 ( .A1(n1536), .A2(n1083), .B1(n1082), .B2(n4), .ZN(n874) );
  OAI22_X1 U1627 ( .A1(n1536), .A2(n1073), .B1(n1072), .B2(n4), .ZN(n864) );
  AND2_X1 U1628 ( .A1(n1571), .A2(n644), .ZN(n719) );
  OAI22_X1 U1629 ( .A1(n1536), .A2(n1074), .B1(n1073), .B2(n4), .ZN(n865) );
  AND2_X1 U1630 ( .A1(n1571), .A2(n656), .ZN(n799) );
  OAI22_X1 U1631 ( .A1(n1536), .A2(n1081), .B1(n1080), .B2(n4), .ZN(n872) );
  OAI22_X1 U1632 ( .A1(n1536), .A2(n1078), .B1(n1077), .B2(n4), .ZN(n869) );
  INV_X1 U1633 ( .A(n640), .ZN(n680) );
  INV_X1 U1634 ( .A(n368), .ZN(n369) );
  XNOR2_X1 U1635 ( .A(n1570), .B(n1569), .ZN(n899) );
  INV_X1 U1636 ( .A(n1569), .ZN(n1140) );
  INV_X1 U1637 ( .A(n661), .ZN(n820) );
  OR2_X1 U1638 ( .A1(n1356), .A2(n1143), .ZN(n963) );
  OR2_X1 U1639 ( .A1(n1570), .A2(n1140), .ZN(n900) );
  OR2_X1 U1640 ( .A1(n1356), .A2(n1146), .ZN(n1026) );
  OR2_X1 U1641 ( .A1(n1571), .A2(n1142), .ZN(n942) );
  OR2_X1 U1642 ( .A1(n1570), .A2(n1145), .ZN(n1005) );
  OR2_X1 U1643 ( .A1(n1571), .A2(n1141), .ZN(n921) );
  XNOR2_X1 U1644 ( .A(n1350), .B(n1287), .ZN(n880) );
  AND2_X1 U1645 ( .A1(n1571), .A2(n1241), .ZN(product[0]) );
  XNOR2_X1 U1646 ( .A(n1), .B(a[2]), .ZN(n9) );
  BUF_X1 U1647 ( .A(n6), .Z(n1534) );
  NAND2_X1 U1648 ( .A1(n1119), .A2(n1368), .ZN(n6) );
  AOI21_X1 U1649 ( .B1(n1528), .B2(n247), .A(n244), .ZN(n242) );
  XNOR2_X1 U1650 ( .A(n90), .B(n247), .ZN(product[6]) );
  XNOR2_X1 U1651 ( .A(n43), .B(a[16]), .ZN(n52) );
  XNOR2_X1 U1652 ( .A(n1566), .B(a[14]), .ZN(n46) );
  XNOR2_X1 U1653 ( .A(n1568), .B(a[18]), .ZN(n58) );
  XNOR2_X1 U1654 ( .A(n7), .B(a[4]), .ZN(n16) );
  XNOR2_X1 U1655 ( .A(n1564), .B(a[10]), .ZN(n34) );
  XNOR2_X1 U1656 ( .A(n1565), .B(a[12]), .ZN(n1544) );
  NOR2_X1 U1657 ( .A1(n397), .A2(n410), .ZN(n1546) );
  NOR2_X1 U1658 ( .A1(n397), .A2(n410), .ZN(n147) );
  NAND2_X1 U1659 ( .A1(n609), .A2(n616), .ZN(n232) );
  OAI21_X1 U1660 ( .B1(n248), .B2(n250), .A(n249), .ZN(n247) );
  INV_X1 U1661 ( .A(n248), .ZN(n293) );
  NOR2_X1 U1662 ( .A1(n633), .A2(n636), .ZN(n248) );
  NAND2_X1 U1663 ( .A1(n427), .A2(n442), .ZN(n159) );
  OAI21_X1 U1664 ( .B1(n163), .B2(n1434), .A(n1468), .ZN(n160) );
  INV_X1 U1665 ( .A(n1434), .ZN(n277) );
  XNOR2_X1 U1666 ( .A(n1375), .B(n1323), .ZN(n923) );
  XNOR2_X1 U1667 ( .A(n1350), .B(n1323), .ZN(n922) );
  XNOR2_X1 U1668 ( .A(n1371), .B(n1323), .ZN(n924) );
  XNOR2_X1 U1669 ( .A(n1377), .B(n1323), .ZN(n926) );
  XNOR2_X1 U1670 ( .A(n1338), .B(n1323), .ZN(n925) );
  XNOR2_X1 U1671 ( .A(n1381), .B(n1323), .ZN(n927) );
  XNOR2_X1 U1672 ( .A(n1333), .B(n1323), .ZN(n928) );
  XNOR2_X1 U1673 ( .A(n1345), .B(n1567), .ZN(n929) );
  XNOR2_X1 U1674 ( .A(n1362), .B(n1567), .ZN(n930) );
  XNOR2_X1 U1675 ( .A(n1579), .B(n1567), .ZN(n932) );
  XNOR2_X1 U1676 ( .A(n1580), .B(n1567), .ZN(n931) );
  XNOR2_X1 U1677 ( .A(n1370), .B(n1567), .ZN(n933) );
  XNOR2_X1 U1678 ( .A(n1382), .B(n1567), .ZN(n935) );
  XNOR2_X1 U1679 ( .A(n1380), .B(n1567), .ZN(n934) );
  XNOR2_X1 U1680 ( .A(n1571), .B(n1567), .ZN(n941) );
  XNOR2_X1 U1681 ( .A(n1352), .B(n1567), .ZN(n939) );
  XNOR2_X1 U1682 ( .A(n1572), .B(n1567), .ZN(n940) );
  XNOR2_X1 U1683 ( .A(n1574), .B(n1567), .ZN(n938) );
  XNOR2_X1 U1684 ( .A(n1576), .B(n1567), .ZN(n936) );
  XNOR2_X1 U1685 ( .A(n1366), .B(n1567), .ZN(n937) );
  INV_X1 U1686 ( .A(n1567), .ZN(n1142) );
  OAI21_X1 U1687 ( .B1(n215), .B2(n219), .A(n216), .ZN(n214) );
  NOR2_X1 U1688 ( .A1(n1332), .A2(n218), .ZN(n213) );
  INV_X1 U1689 ( .A(n1332), .ZN(n286) );
  NOR2_X1 U1690 ( .A1(n581), .A2(n590), .ZN(n215) );
  INV_X1 U1691 ( .A(n1234), .ZN(n280) );
  NOR2_X1 U1692 ( .A1(n1234), .A2(n180), .ZN(n175) );
  AOI21_X1 U1693 ( .B1(n173), .B2(n1267), .A(n1320), .ZN(n163) );
  AND2_X1 U1694 ( .A1(n529), .A2(n542), .ZN(n1548) );
  XNOR2_X1 U1695 ( .A(n1326), .B(n1489), .ZN(n901) );
  XNOR2_X1 U1696 ( .A(n1375), .B(n1489), .ZN(n902) );
  NOR2_X1 U1697 ( .A1(n131), .A2(n128), .ZN(n126) );
  XNOR2_X1 U1698 ( .A(n1339), .B(n1489), .ZN(n904) );
  XNOR2_X1 U1699 ( .A(n1371), .B(n1489), .ZN(n903) );
  XNOR2_X1 U1700 ( .A(n1378), .B(n1489), .ZN(n905) );
  XNOR2_X1 U1701 ( .A(n1381), .B(n1489), .ZN(n906) );
  XNOR2_X1 U1702 ( .A(n1583), .B(n1489), .ZN(n907) );
  XNOR2_X1 U1703 ( .A(n1582), .B(n1489), .ZN(n908) );
  XNOR2_X1 U1704 ( .A(n1362), .B(n1489), .ZN(n909) );
  XNOR2_X1 U1705 ( .A(n1580), .B(n1489), .ZN(n910) );
  XNOR2_X1 U1706 ( .A(n1579), .B(n1489), .ZN(n911) );
  XNOR2_X1 U1707 ( .A(n1370), .B(n1489), .ZN(n912) );
  XNOR2_X1 U1708 ( .A(n1577), .B(n1489), .ZN(n914) );
  XNOR2_X1 U1709 ( .A(n1322), .B(n1489), .ZN(n913) );
  XNOR2_X1 U1710 ( .A(n1266), .B(n1489), .ZN(n918) );
  XNOR2_X1 U1711 ( .A(n1363), .B(n1489), .ZN(n917) );
  XNOR2_X1 U1712 ( .A(n1570), .B(n1489), .ZN(n920) );
  XNOR2_X1 U1713 ( .A(n1365), .B(n1489), .ZN(n916) );
  XNOR2_X1 U1714 ( .A(n1576), .B(n1489), .ZN(n915) );
  XNOR2_X1 U1715 ( .A(n1572), .B(n1489), .ZN(n919) );
  INV_X1 U1716 ( .A(n1489), .ZN(n1141) );
  NAND2_X1 U1717 ( .A1(n156), .A2(n164), .ZN(n154) );
  XNOR2_X1 U1718 ( .A(n1326), .B(n1387), .ZN(n943) );
  XNOR2_X1 U1719 ( .A(n1375), .B(n1387), .ZN(n944) );
  XNOR2_X1 U1720 ( .A(n1339), .B(n1387), .ZN(n946) );
  XNOR2_X1 U1721 ( .A(n1371), .B(n1387), .ZN(n945) );
  XNOR2_X1 U1722 ( .A(n1378), .B(n1387), .ZN(n947) );
  XNOR2_X1 U1723 ( .A(n1381), .B(n1387), .ZN(n948) );
  XNOR2_X1 U1724 ( .A(n1362), .B(n1387), .ZN(n951) );
  XNOR2_X1 U1725 ( .A(n1345), .B(n1387), .ZN(n950) );
  XNOR2_X1 U1726 ( .A(n1333), .B(n1387), .ZN(n949) );
  XNOR2_X1 U1727 ( .A(n1285), .B(n1387), .ZN(n952) );
  XNOR2_X1 U1728 ( .A(n1382), .B(n1387), .ZN(n956) );
  INV_X1 U1729 ( .A(n1387), .ZN(n1143) );
  XNOR2_X1 U1730 ( .A(n1576), .B(n1387), .ZN(n957) );
  XNOR2_X1 U1731 ( .A(n1265), .B(n1387), .ZN(n960) );
  XNOR2_X1 U1732 ( .A(n1369), .B(n1387), .ZN(n954) );
  XNOR2_X1 U1733 ( .A(n1579), .B(n1387), .ZN(n953) );
  XNOR2_X1 U1734 ( .A(n1570), .B(n1387), .ZN(n962) );
  XNOR2_X1 U1735 ( .A(n1363), .B(n1387), .ZN(n959) );
  XNOR2_X1 U1736 ( .A(n1365), .B(n1387), .ZN(n958) );
  XNOR2_X1 U1737 ( .A(n1572), .B(n1387), .ZN(n961) );
  INV_X1 U1738 ( .A(n1243), .ZN(n1549) );
  INV_X1 U1739 ( .A(n1244), .ZN(n1550) );
  NAND2_X1 U1740 ( .A1(n275), .A2(n1483), .ZN(n73) );
  XOR2_X1 U1741 ( .A(n1310), .B(n564), .Z(n1552) );
  XOR2_X1 U1742 ( .A(n551), .B(n1552), .Z(n547) );
  NAND2_X1 U1743 ( .A1(n551), .A2(n1309), .ZN(n1553) );
  NAND2_X1 U1744 ( .A1(n551), .A2(n564), .ZN(n1554) );
  NAND2_X1 U1745 ( .A1(n562), .A2(n564), .ZN(n1555) );
  NAND3_X1 U1746 ( .A1(n1553), .A2(n1554), .A3(n1555), .ZN(n546) );
  AOI21_X1 U1747 ( .B1(n239), .B2(n1522), .A(n236), .ZN(n1556) );
  AND2_X1 U1748 ( .A1(n513), .A2(n528), .ZN(n1557) );
  OR2_X1 U1749 ( .A1(n1571), .A2(n1144), .ZN(n984) );
  XNOR2_X1 U1750 ( .A(n1350), .B(n1384), .ZN(n1006) );
  INV_X1 U1751 ( .A(n1509), .ZN(n1146) );
  XNOR2_X1 U1752 ( .A(n1588), .B(n1509), .ZN(n1007) );
  XNOR2_X1 U1753 ( .A(n1587), .B(n1509), .ZN(n1008) );
  XNOR2_X1 U1754 ( .A(n1339), .B(n1509), .ZN(n1009) );
  XNOR2_X1 U1755 ( .A(n1570), .B(n1384), .ZN(n1025) );
  XNOR2_X1 U1756 ( .A(n1572), .B(n1384), .ZN(n1024) );
  XNOR2_X1 U1757 ( .A(n1581), .B(n1509), .ZN(n1014) );
  XNOR2_X1 U1758 ( .A(n1584), .B(n1509), .ZN(n1011) );
  XNOR2_X1 U1759 ( .A(n1576), .B(n1509), .ZN(n1020) );
  XNOR2_X1 U1760 ( .A(n1366), .B(n1384), .ZN(n1021) );
  XNOR2_X1 U1761 ( .A(n1582), .B(n1509), .ZN(n1013) );
  XNOR2_X1 U1762 ( .A(n1583), .B(n1509), .ZN(n1012) );
  XNOR2_X1 U1763 ( .A(n1377), .B(n1509), .ZN(n1010) );
  XNOR2_X1 U1764 ( .A(n1319), .B(n1509), .ZN(n1019) );
  XNOR2_X1 U1765 ( .A(n1352), .B(n1509), .ZN(n1023) );
  XNOR2_X1 U1766 ( .A(n1363), .B(n1509), .ZN(n1022) );
  XNOR2_X1 U1767 ( .A(n1322), .B(n1509), .ZN(n1018) );
  XNOR2_X1 U1768 ( .A(n1580), .B(n1509), .ZN(n1015) );
  XNOR2_X1 U1769 ( .A(n1369), .B(n1509), .ZN(n1017) );
  XNOR2_X1 U1770 ( .A(n1579), .B(n1509), .ZN(n1016) );
  XOR2_X1 U1771 ( .A(n1538), .B(a[6]), .Z(n1116) );
  NAND2_X1 U1772 ( .A1(n411), .A2(n426), .ZN(n151) );
  NAND2_X1 U1773 ( .A1(n815), .A2(n870), .ZN(n1560) );
  NAND2_X1 U1774 ( .A1(n815), .A2(n779), .ZN(n1561) );
  NAND2_X1 U1775 ( .A1(n870), .A2(n779), .ZN(n1562) );
  NAND3_X1 U1776 ( .A1(n1560), .A2(n1561), .A3(n1562), .ZN(n606) );
  AND2_X1 U1777 ( .A1(n1356), .A2(n653), .ZN(n779) );
  OAI22_X1 U1778 ( .A1(n1536), .A2(n1079), .B1(n1078), .B2(n4), .ZN(n870) );
  INV_X1 U1779 ( .A(n1471), .ZN(n1149) );
  XNOR2_X1 U1780 ( .A(n1265), .B(n1471), .ZN(n1086) );
  XNOR2_X1 U1781 ( .A(n1574), .B(n1471), .ZN(n1085) );
  XNOR2_X1 U1782 ( .A(n1366), .B(n1470), .ZN(n1084) );
  XNOR2_X1 U1783 ( .A(n1584), .B(n1471), .ZN(n1074) );
  XNOR2_X1 U1784 ( .A(n1094), .B(n1470), .ZN(n1073) );
  XNOR2_X1 U1785 ( .A(n1577), .B(n1470), .ZN(n1082) );
  XNOR2_X1 U1786 ( .A(n1587), .B(n1471), .ZN(n1071) );
  XNOR2_X1 U1787 ( .A(n1345), .B(n1471), .ZN(n1076) );
  XNOR2_X1 U1788 ( .A(n1581), .B(n1470), .ZN(n1077) );
  XNOR2_X1 U1789 ( .A(n1369), .B(n1471), .ZN(n1080) );
  XNOR2_X1 U1790 ( .A(n1379), .B(n1471), .ZN(n1081) );
  XNOR2_X1 U1791 ( .A(n1333), .B(n1471), .ZN(n1075) );
  XNOR2_X1 U1792 ( .A(n1588), .B(n1470), .ZN(n1070) );
  XNOR2_X1 U1793 ( .A(n1576), .B(n1471), .ZN(n1083) );
  XNOR2_X1 U1794 ( .A(n1579), .B(n1470), .ZN(n1079) );
  XNOR2_X1 U1795 ( .A(n1339), .B(n1471), .ZN(n1072) );
  XNOR2_X1 U1796 ( .A(n1285), .B(n1471), .ZN(n1078) );
  XNOR2_X1 U1797 ( .A(n1571), .B(n1470), .ZN(n1088) );
  XNOR2_X1 U1798 ( .A(n1572), .B(n1471), .ZN(n1087) );
  XNOR2_X1 U1799 ( .A(n1355), .B(n1470), .ZN(n1069) );
  NAND2_X1 U1800 ( .A1(n639), .A2(n678), .ZN(n257) );
  OAI22_X1 U1801 ( .A1(n1535), .A2(n1086), .B1(n1085), .B2(n4), .ZN(n877) );
  INV_X1 U1802 ( .A(n1546), .ZN(n274) );
  OAI21_X1 U1803 ( .B1(n151), .B2(n147), .A(n148), .ZN(n146) );
  NAND2_X1 U1804 ( .A1(n397), .A2(n410), .ZN(n148) );
  INV_X1 U1805 ( .A(n204), .ZN(n284) );
  NOR2_X1 U1806 ( .A1(n204), .A2(n209), .ZN(n202) );
  OAI21_X1 U1807 ( .B1(n204), .B2(n210), .A(n205), .ZN(n203) );
  XNOR2_X1 U1808 ( .A(n1326), .B(n1385), .ZN(n985) );
  XNOR2_X1 U1809 ( .A(n1375), .B(n1385), .ZN(n986) );
  XNOR2_X1 U1810 ( .A(n1338), .B(n1385), .ZN(n988) );
  XNOR2_X1 U1811 ( .A(n1587), .B(n1385), .ZN(n987) );
  XNOR2_X1 U1812 ( .A(n1377), .B(n1385), .ZN(n989) );
  XNOR2_X1 U1813 ( .A(n1583), .B(n1385), .ZN(n991) );
  XNOR2_X1 U1814 ( .A(n1584), .B(n1385), .ZN(n990) );
  XNOR2_X1 U1815 ( .A(n1356), .B(n1271), .ZN(n1004) );
  XNOR2_X1 U1816 ( .A(n1576), .B(n1385), .ZN(n999) );
  XNOR2_X1 U1817 ( .A(n1579), .B(n1385), .ZN(n995) );
  XNOR2_X1 U1818 ( .A(n1345), .B(n1271), .ZN(n992) );
  INV_X1 U1819 ( .A(n1271), .ZN(n1145) );
  XNOR2_X1 U1820 ( .A(n1572), .B(n1271), .ZN(n1003) );
  XNOR2_X1 U1821 ( .A(n1362), .B(n1271), .ZN(n993) );
  XNOR2_X1 U1822 ( .A(n1580), .B(n1385), .ZN(n994) );
  XNOR2_X1 U1823 ( .A(n1266), .B(n1271), .ZN(n1002) );
  XNOR2_X1 U1824 ( .A(n1319), .B(n1271), .ZN(n998) );
  XNOR2_X1 U1825 ( .A(n1322), .B(n1271), .ZN(n997) );
  XNOR2_X1 U1826 ( .A(n1366), .B(n1271), .ZN(n1000) );
  XNOR2_X1 U1827 ( .A(n1574), .B(n1385), .ZN(n1001) );
  XNOR2_X1 U1828 ( .A(n1369), .B(n1271), .ZN(n996) );
  XOR2_X1 U1829 ( .A(n25), .B(a[8]), .Z(n1115) );
  XNOR2_X1 U1830 ( .A(n1350), .B(n1400), .ZN(n964) );
  XNOR2_X1 U1831 ( .A(n1375), .B(n1400), .ZN(n965) );
  XNOR2_X1 U1832 ( .A(n1371), .B(n1400), .ZN(n966) );
  XNOR2_X1 U1833 ( .A(n1338), .B(n1400), .ZN(n967) );
  XNOR2_X1 U1834 ( .A(n1098), .B(n1400), .ZN(n972) );
  XNOR2_X1 U1835 ( .A(n1377), .B(n1400), .ZN(n968) );
  XNOR2_X1 U1836 ( .A(n1584), .B(n1400), .ZN(n969) );
  XNOR2_X1 U1837 ( .A(n1333), .B(n1400), .ZN(n970) );
  XNOR2_X1 U1838 ( .A(n1582), .B(n1400), .ZN(n971) );
  XNOR2_X1 U1839 ( .A(n1379), .B(n1400), .ZN(n976) );
  INV_X1 U1840 ( .A(n1400), .ZN(n1144) );
  XNOR2_X1 U1841 ( .A(n1369), .B(n1400), .ZN(n975) );
  XNOR2_X1 U1842 ( .A(n1570), .B(n1400), .ZN(n983) );
  XNOR2_X1 U1843 ( .A(n1577), .B(n1400), .ZN(n977) );
  XNOR2_X1 U1844 ( .A(n1285), .B(n1400), .ZN(n973) );
  XNOR2_X1 U1845 ( .A(n1579), .B(n1400), .ZN(n974) );
  XNOR2_X1 U1846 ( .A(n1572), .B(n1400), .ZN(n982) );
  XNOR2_X1 U1847 ( .A(n1576), .B(n1400), .ZN(n978) );
  XNOR2_X1 U1848 ( .A(n1366), .B(n1400), .ZN(n979) );
  XNOR2_X1 U1849 ( .A(n1363), .B(n1400), .ZN(n980) );
  XNOR2_X1 U1850 ( .A(n1351), .B(n1400), .ZN(n981) );
  INV_X1 U1851 ( .A(n1503), .ZN(n276) );
  OAI21_X1 U1852 ( .B1(n162), .B2(n158), .A(n159), .ZN(n157) );
  INV_X1 U1853 ( .A(n1286), .ZN(n139) );
  OAI21_X1 U1854 ( .B1(n141), .B2(n135), .A(n136), .ZN(n134) );
  NAND2_X1 U1855 ( .A1(n273), .A2(n1286), .ZN(n71) );
  NAND2_X1 U1856 ( .A1(n383), .A2(n396), .ZN(n141) );
  XNOR2_X1 U1857 ( .A(n1351), .B(n1308), .ZN(n1044) );
  XNOR2_X1 U1858 ( .A(n1378), .B(n1252), .ZN(n1031) );
  INV_X1 U1859 ( .A(n1308), .ZN(n1147) );
  XNOR2_X1 U1860 ( .A(n1370), .B(n1308), .ZN(n1038) );
  XNOR2_X1 U1861 ( .A(n1579), .B(n1252), .ZN(n1037) );
  XNOR2_X1 U1862 ( .A(n1356), .B(n1252), .ZN(n1046) );
  XNOR2_X1 U1863 ( .A(n1583), .B(n1373), .ZN(n1033) );
  XNOR2_X1 U1864 ( .A(n1363), .B(n1373), .ZN(n1043) );
  XNOR2_X1 U1865 ( .A(n1285), .B(n1252), .ZN(n1036) );
  XNOR2_X1 U1866 ( .A(n1355), .B(n1252), .ZN(n1027) );
  XNOR2_X1 U1867 ( .A(n1337), .B(n1373), .ZN(n1030) );
  XNOR2_X1 U1868 ( .A(n1366), .B(n1252), .ZN(n1042) );
  XNOR2_X1 U1869 ( .A(n1576), .B(n1373), .ZN(n1041) );
  XNOR2_X1 U1870 ( .A(n1587), .B(n1252), .ZN(n1029) );
  XNOR2_X1 U1871 ( .A(n1584), .B(n1373), .ZN(n1032) );
  XNOR2_X1 U1872 ( .A(n1572), .B(n1252), .ZN(n1045) );
  XNOR2_X1 U1873 ( .A(n1577), .B(n1252), .ZN(n1040) );
  XNOR2_X1 U1874 ( .A(n1379), .B(n1252), .ZN(n1039) );
  XNOR2_X1 U1875 ( .A(n1588), .B(n1252), .ZN(n1028) );
  XNOR2_X1 U1876 ( .A(n1581), .B(n1252), .ZN(n1035) );
  XNOR2_X1 U1877 ( .A(n1582), .B(n1252), .ZN(n1034) );
  XNOR2_X1 U1878 ( .A(n1576), .B(n1359), .ZN(n1062) );
  XNOR2_X1 U1879 ( .A(n1370), .B(n1358), .ZN(n1059) );
  INV_X1 U1880 ( .A(n1358), .ZN(n1148) );
  XNOR2_X1 U1881 ( .A(n1582), .B(n1358), .ZN(n1055) );
  XNOR2_X1 U1882 ( .A(n1581), .B(n1359), .ZN(n1056) );
  XNOR2_X1 U1883 ( .A(n1363), .B(n1358), .ZN(n1064) );
  XNOR2_X1 U1884 ( .A(n1379), .B(n1358), .ZN(n1060) );
  XNOR2_X1 U1885 ( .A(n1319), .B(n1359), .ZN(n1061) );
  XNOR2_X1 U1886 ( .A(n1366), .B(n1359), .ZN(n1063) );
  XNOR2_X1 U1887 ( .A(n1337), .B(n1358), .ZN(n1051) );
  XNOR2_X1 U1888 ( .A(n1378), .B(n1358), .ZN(n1052) );
  XNOR2_X1 U1889 ( .A(n1333), .B(n1359), .ZN(n1054) );
  XNOR2_X1 U1890 ( .A(n1580), .B(n1358), .ZN(n1057) );
  XNOR2_X1 U1891 ( .A(n1579), .B(n1359), .ZN(n1058) );
  XNOR2_X1 U1892 ( .A(n1571), .B(n1359), .ZN(n1067) );
  XNOR2_X1 U1893 ( .A(n1584), .B(n1358), .ZN(n1053) );
  XNOR2_X1 U1894 ( .A(n1266), .B(n1359), .ZN(n1065) );
  XNOR2_X1 U1895 ( .A(n1572), .B(n1358), .ZN(n1066) );
  XNOR2_X1 U1896 ( .A(n1587), .B(n1359), .ZN(n1050) );
  XNOR2_X1 U1897 ( .A(n1588), .B(n1358), .ZN(n1049) );
  XNOR2_X1 U1898 ( .A(n1090), .B(n7), .ZN(n1048) );
  OR2_X1 U1899 ( .A1(n787), .A2(n715), .ZN(n476) );
  NAND2_X1 U1900 ( .A1(n637), .A2(n638), .ZN(n254) );
  NAND2_X1 U1901 ( .A1(n145), .A2(n133), .ZN(n131) );
  INV_X1 U1902 ( .A(n212), .ZN(n211) );
  OAI21_X1 U1903 ( .B1(n152), .B2(n131), .A(n1488), .ZN(n130) );
  AOI21_X1 U1904 ( .B1(n203), .B2(n1521), .A(n198), .ZN(n196) );
  NAND2_X1 U1905 ( .A1(n202), .A2(n1521), .ZN(n195) );
  NAND2_X1 U1906 ( .A1(n1521), .A2(n200), .ZN(n81) );
  AOI21_X1 U1907 ( .B1(n239), .B2(n1522), .A(n236), .ZN(n234) );
  NOR2_X1 U1908 ( .A1(n140), .A2(n135), .ZN(n133) );
  NOR2_X1 U1909 ( .A1(n383), .A2(n396), .ZN(n140) );
  INV_X1 U1910 ( .A(n664), .ZN(n840) );
  NAND2_X1 U1911 ( .A1(n1547), .A2(n1312), .ZN(n180) );
  NAND2_X1 U1912 ( .A1(n1547), .A2(n185), .ZN(n79) );
  AOI21_X1 U1913 ( .B1(n1547), .B2(n1548), .A(n1557), .ZN(n181) );
  OAI21_X1 U1914 ( .B1(n193), .B2(n187), .A(n188), .ZN(n186) );
  NOR2_X1 U1915 ( .A1(n161), .A2(n1503), .ZN(n156) );
  XNOR2_X1 U1916 ( .A(n787), .B(n715), .ZN(n477) );
  INV_X1 U1917 ( .A(n1441), .ZN(n193) );
  INV_X1 U1918 ( .A(n1542), .ZN(n653) );
  INV_X1 U1919 ( .A(n1507), .ZN(n278) );
  OAI22_X1 U1920 ( .A1(n922), .A2(n1263), .B1(n922), .B2(n1539), .ZN(n646) );
  NOR2_X1 U1921 ( .A1(n171), .A2(n1507), .ZN(n164) );
  OAI21_X1 U1922 ( .B1(n166), .B2(n172), .A(n167), .ZN(n165) );
  OAI22_X1 U1923 ( .A1(n1263), .A2(n924), .B1(n923), .B2(n1539), .ZN(n721) );
  OAI22_X1 U1924 ( .A1(n1388), .A2(n923), .B1(n922), .B2(n1539), .ZN(n314) );
  NAND2_X1 U1925 ( .A1(n461), .A2(n478), .ZN(n167) );
  OAI22_X1 U1926 ( .A1(n1263), .A2(n925), .B1(n924), .B2(n1539), .ZN(n722) );
  OAI22_X1 U1927 ( .A1(n1388), .A2(n927), .B1(n926), .B2(n1539), .ZN(n724) );
  OAI22_X1 U1928 ( .A1(n1388), .A2(n926), .B1(n925), .B2(n1539), .ZN(n723) );
  OAI22_X1 U1929 ( .A1(n1263), .A2(n928), .B1(n927), .B2(n1539), .ZN(n725) );
  OAI22_X1 U1930 ( .A1(n1263), .A2(n929), .B1(n928), .B2(n1539), .ZN(n726) );
  OAI22_X1 U1931 ( .A1(n1388), .A2(n930), .B1(n929), .B2(n1539), .ZN(n727) );
  OAI22_X1 U1932 ( .A1(n1388), .A2(n933), .B1(n932), .B2(n1539), .ZN(n730) );
  OAI22_X1 U1933 ( .A1(n1558), .A2(n931), .B1(n930), .B2(n1539), .ZN(n728) );
  OAI22_X1 U1934 ( .A1(n1559), .A2(n932), .B1(n931), .B2(n1539), .ZN(n729) );
  OAI22_X1 U1935 ( .A1(n1559), .A2(n935), .B1(n934), .B2(n1540), .ZN(n732) );
  OAI22_X1 U1936 ( .A1(n1388), .A2(n934), .B1(n933), .B2(n1539), .ZN(n731) );
  OAI22_X1 U1937 ( .A1(n1558), .A2(n939), .B1(n938), .B2(n1539), .ZN(n736) );
  OAI22_X1 U1938 ( .A1(n1559), .A2(n936), .B1(n935), .B2(n1540), .ZN(n733) );
  OAI22_X1 U1939 ( .A1(n1559), .A2(n940), .B1(n939), .B2(n1540), .ZN(n737) );
  OAI22_X1 U1940 ( .A1(n1388), .A2(n941), .B1(n940), .B2(n1539), .ZN(n738) );
  OAI22_X1 U1941 ( .A1(n1263), .A2(n1142), .B1(n942), .B2(n1539), .ZN(n672) );
  OAI22_X1 U1942 ( .A1(n1558), .A2(n937), .B1(n1540), .B2(n1317), .ZN(n734) );
  INV_X1 U1943 ( .A(n1540), .ZN(n647) );
  OAI21_X1 U1944 ( .B1(n152), .B2(n1307), .A(n1483), .ZN(n149) );
  INV_X1 U1945 ( .A(n1307), .ZN(n275) );
  OAI22_X1 U1946 ( .A1(n880), .A2(n1490), .B1(n880), .B2(n1505), .ZN(n640) );
  OAI22_X1 U1947 ( .A1(n1490), .A2(n881), .B1(n880), .B2(n1506), .ZN(n298) );
  OAI22_X1 U1948 ( .A1(n1490), .A2(n882), .B1(n881), .B2(n1505), .ZN(n681) );
  OAI22_X1 U1949 ( .A1(n1490), .A2(n883), .B1(n882), .B2(n1506), .ZN(n682) );
  OAI22_X1 U1950 ( .A1(n1490), .A2(n884), .B1(n883), .B2(n1505), .ZN(n683) );
  NOR2_X1 U1951 ( .A1(n150), .A2(n1546), .ZN(n145) );
  OAI22_X1 U1952 ( .A1(n1436), .A2(n886), .B1(n885), .B2(n1505), .ZN(n685) );
  OAI22_X1 U1953 ( .A1(n1436), .A2(n885), .B1(n884), .B2(n1506), .ZN(n684) );
  OAI22_X1 U1954 ( .A1(n1436), .A2(n887), .B1(n886), .B2(n1506), .ZN(n686) );
  OAI22_X1 U1955 ( .A1(n1436), .A2(n888), .B1(n887), .B2(n1505), .ZN(n687) );
  OAI22_X1 U1956 ( .A1(n1436), .A2(n889), .B1(n888), .B2(n1506), .ZN(n688) );
  OAI22_X1 U1957 ( .A1(n1436), .A2(n890), .B1(n889), .B2(n1505), .ZN(n689) );
  OAI22_X1 U1958 ( .A1(n60), .A2(n891), .B1(n890), .B2(n1506), .ZN(n690) );
  OAI22_X1 U1959 ( .A1(n60), .A2(n892), .B1(n891), .B2(n1505), .ZN(n691) );
  OAI22_X1 U1960 ( .A1(n60), .A2(n894), .B1(n893), .B2(n1506), .ZN(n693) );
  OAI22_X1 U1961 ( .A1(n60), .A2(n893), .B1(n892), .B2(n1506), .ZN(n692) );
  OAI22_X1 U1962 ( .A1(n60), .A2(n899), .B1(n898), .B2(n1505), .ZN(n698) );
  OAI22_X1 U1963 ( .A1(n60), .A2(n895), .B1(n894), .B2(n1505), .ZN(n694) );
  OAI22_X1 U1964 ( .A1(n60), .A2(n1140), .B1(n900), .B2(n1505), .ZN(n670) );
  OAI22_X1 U1965 ( .A1(n896), .A2(n60), .B1(n895), .B2(n1505), .ZN(n695) );
  OAI22_X1 U1966 ( .A1(n60), .A2(n898), .B1(n897), .B2(n1504), .ZN(n697) );
  INV_X1 U1967 ( .A(n1504), .ZN(n641) );
  OAI22_X1 U1968 ( .A1(n60), .A2(n897), .B1(n896), .B2(n1504), .ZN(n696) );
  OAI21_X1 U1969 ( .B1(n195), .B2(n212), .A(n196), .ZN(n194) );
  XOR2_X1 U1970 ( .A(n242), .B(n89), .Z(product[7]) );
  INV_X1 U1971 ( .A(n1556), .ZN(n233) );
  OAI21_X1 U1972 ( .B1(n222), .B2(n234), .A(n223), .ZN(n221) );
  OAI21_X1 U1973 ( .B1(n242), .B2(n240), .A(n241), .ZN(n239) );
  OAI22_X1 U1974 ( .A1(n1501), .A2(n1053), .B1(n1052), .B2(n1533), .ZN(n844)
         );
  OAI22_X1 U1975 ( .A1(n1501), .A2(n1055), .B1(n1054), .B2(n1532), .ZN(n846)
         );
  OAI22_X1 U1976 ( .A1(n1501), .A2(n1051), .B1(n1050), .B2(n1533), .ZN(n842)
         );
  OAI22_X1 U1977 ( .A1(n1240), .A2(n1062), .B1(n1061), .B2(n1532), .ZN(n853)
         );
  OAI22_X1 U1978 ( .A1(n1240), .A2(n1059), .B1(n1058), .B2(n1533), .ZN(n850)
         );
  OAI22_X1 U1979 ( .A1(n1240), .A2(n1060), .B1(n1059), .B2(n1533), .ZN(n851)
         );
  OAI22_X1 U1980 ( .A1(n1052), .A2(n1502), .B1(n1051), .B2(n1532), .ZN(n843)
         );
  OAI22_X1 U1981 ( .A1(n1502), .A2(n1063), .B1(n1062), .B2(n1532), .ZN(n854)
         );
  OAI22_X1 U1982 ( .A1(n1501), .A2(n1054), .B1(n1053), .B2(n1532), .ZN(n845)
         );
  OAI22_X1 U1983 ( .A1(n1501), .A2(n1049), .B1(n1048), .B2(n1533), .ZN(n458)
         );
  OAI22_X1 U1984 ( .A1(n1501), .A2(n1056), .B1(n1055), .B2(n1532), .ZN(n847)
         );
  OAI22_X1 U1985 ( .A1(n1502), .A2(n1057), .B1(n1056), .B2(n1532), .ZN(n848)
         );
  OAI22_X1 U1986 ( .A1(n1501), .A2(n1065), .B1(n1064), .B2(n1532), .ZN(n856)
         );
  OAI22_X1 U1987 ( .A1(n1502), .A2(n1050), .B1(n1049), .B2(n1532), .ZN(n841)
         );
  OAI22_X1 U1988 ( .A1(n1502), .A2(n1058), .B1(n1057), .B2(n1532), .ZN(n849)
         );
  OAI22_X1 U1989 ( .A1(n1501), .A2(n1148), .B1(n1068), .B2(n1533), .ZN(n678)
         );
  OAI22_X1 U1990 ( .A1(n1240), .A2(n1061), .B1(n1060), .B2(n1532), .ZN(n852)
         );
  OAI22_X1 U1991 ( .A1(n12), .A2(n1048), .B1(n1048), .B2(n1533), .ZN(n664) );
  OAI22_X1 U1992 ( .A1(n1502), .A2(n1064), .B1(n1063), .B2(n1533), .ZN(n855)
         );
  OAI22_X1 U1993 ( .A1(n1501), .A2(n1067), .B1(n1066), .B2(n1533), .ZN(n858)
         );
  OAI22_X1 U1994 ( .A1(n1502), .A2(n1066), .B1(n1065), .B2(n1533), .ZN(n857)
         );
  INV_X1 U1995 ( .A(n1533), .ZN(n665) );
  OAI22_X1 U1996 ( .A1(n901), .A2(n1364), .B1(n901), .B2(n1498), .ZN(n643) );
  OAI22_X1 U1997 ( .A1(n1364), .A2(n902), .B1(n901), .B2(n1499), .ZN(n304) );
  OAI22_X1 U1998 ( .A1(n1364), .A2(n903), .B1(n902), .B2(n1498), .ZN(n701) );
  OAI22_X1 U1999 ( .A1(n1364), .A2(n904), .B1(n903), .B2(n1499), .ZN(n702) );
  OAI22_X1 U2000 ( .A1(n1364), .A2(n905), .B1(n904), .B2(n1498), .ZN(n703) );
  OAI22_X1 U2001 ( .A1(n1364), .A2(n906), .B1(n905), .B2(n1499), .ZN(n704) );
  OAI22_X1 U2002 ( .A1(n1364), .A2(n907), .B1(n906), .B2(n1498), .ZN(n705) );
  OAI22_X1 U2003 ( .A1(n1364), .A2(n908), .B1(n907), .B2(n1499), .ZN(n706) );
  OAI22_X1 U2004 ( .A1(n1364), .A2(n909), .B1(n908), .B2(n1498), .ZN(n707) );
  OAI22_X1 U2005 ( .A1(n1364), .A2(n910), .B1(n909), .B2(n1499), .ZN(n708) );
  OAI22_X1 U2006 ( .A1(n54), .A2(n911), .B1(n910), .B2(n1498), .ZN(n709) );
  OAI22_X1 U2007 ( .A1(n54), .A2(n912), .B1(n911), .B2(n1499), .ZN(n710) );
  OAI22_X1 U2008 ( .A1(n54), .A2(n913), .B1(n912), .B2(n1499), .ZN(n711) );
  OAI22_X1 U2009 ( .A1(n54), .A2(n915), .B1(n914), .B2(n1499), .ZN(n713) );
  OAI22_X1 U2010 ( .A1(n54), .A2(n1141), .B1(n921), .B2(n1498), .ZN(n671) );
  OAI22_X1 U2011 ( .A1(n54), .A2(n914), .B1(n913), .B2(n1498), .ZN(n712) );
  OAI22_X1 U2012 ( .A1(n54), .A2(n920), .B1(n919), .B2(n1499), .ZN(n718) );
  OAI22_X1 U2013 ( .A1(n54), .A2(n918), .B1(n917), .B2(n1499), .ZN(n716) );
  OAI22_X1 U2014 ( .A1(n54), .A2(n919), .B1(n1325), .B2(n1498), .ZN(n717) );
  OAI22_X1 U2015 ( .A1(n54), .A2(n917), .B1(n916), .B2(n1499), .ZN(n715) );
  OAI22_X1 U2016 ( .A1(n54), .A2(n916), .B1(n915), .B2(n1498), .ZN(n714) );
  INV_X1 U2017 ( .A(n1498), .ZN(n644) );
  INV_X1 U2018 ( .A(n1491), .ZN(n173) );
  INV_X1 U2019 ( .A(n1508), .ZN(n152) );
  OAI22_X1 U2020 ( .A1(n985), .A2(n1435), .B1(n985), .B2(n1314), .ZN(n655) );
  OAI22_X1 U2021 ( .A1(n1435), .A2(n986), .B1(n985), .B2(n1314), .ZN(n368) );
  OAI22_X1 U2022 ( .A1(n1435), .A2(n987), .B1(n986), .B2(n1537), .ZN(n781) );
  OAI22_X1 U2023 ( .A1(n1563), .A2(n989), .B1(n988), .B2(n1314), .ZN(n783) );
  OAI22_X1 U2024 ( .A1(n1435), .A2(n992), .B1(n991), .B2(n1314), .ZN(n786) );
  OAI22_X1 U2025 ( .A1(n1435), .A2(n990), .B1(n989), .B2(n1314), .ZN(n784) );
  OAI22_X1 U2026 ( .A1(n1435), .A2(n988), .B1(n987), .B2(n1537), .ZN(n782) );
  OAI22_X1 U2027 ( .A1(n1435), .A2(n1003), .B1(n1002), .B2(n1314), .ZN(n797)
         );
  OAI22_X1 U2028 ( .A1(n1492), .A2(n991), .B1(n990), .B2(n1314), .ZN(n785) );
  OAI22_X1 U2029 ( .A1(n1492), .A2(n996), .B1(n995), .B2(n1314), .ZN(n790) );
  OAI22_X1 U2030 ( .A1(n1435), .A2(n999), .B1(n998), .B2(n1314), .ZN(n793) );
  OAI22_X1 U2031 ( .A1(n1563), .A2(n993), .B1(n992), .B2(n1537), .ZN(n787) );
  OAI22_X1 U2032 ( .A1(n1563), .A2(n995), .B1(n994), .B2(n1537), .ZN(n789) );
  OAI22_X1 U2033 ( .A1(n994), .A2(n1563), .B1(n993), .B2(n1537), .ZN(n788) );
  OAI22_X1 U2034 ( .A1(n1237), .A2(n1563), .B1(n996), .B2(n1537), .ZN(n791) );
  OAI22_X1 U2035 ( .A1(n1492), .A2(n1000), .B1(n999), .B2(n1314), .ZN(n794) );
  OAI22_X1 U2036 ( .A1(n1492), .A2(n998), .B1(n997), .B2(n1314), .ZN(n792) );
  OAI22_X1 U2037 ( .A1(n1563), .A2(n1004), .B1(n1003), .B2(n1537), .ZN(n798)
         );
  OAI22_X1 U2038 ( .A1(n1492), .A2(n1002), .B1(n1001), .B2(n1314), .ZN(n796)
         );
  OAI22_X1 U2039 ( .A1(n1435), .A2(n1145), .B1(n1005), .B2(n1314), .ZN(n675)
         );
  INV_X1 U2040 ( .A(n1314), .ZN(n656) );
  OAI22_X1 U2041 ( .A1(n1492), .A2(n1001), .B1(n1000), .B2(n1537), .ZN(n795)
         );
  AOI21_X1 U2042 ( .B1(n1508), .B2(n126), .A(n1472), .ZN(n125) );
  OAI21_X1 U2043 ( .B1(n132), .B2(n128), .A(n129), .ZN(n127) );
  OAI21_X1 U2044 ( .B1(n174), .B2(n154), .A(n155), .ZN(n153) );
  AOI21_X1 U2045 ( .B1(n194), .B2(n175), .A(n176), .ZN(n174) );
  AOI21_X1 U2046 ( .B1(n156), .B2(n165), .A(n157), .ZN(n155) );
  OAI22_X1 U2047 ( .A1(n1330), .A2(n965), .B1(n964), .B2(n1543), .ZN(n346) );
  OAI22_X1 U2048 ( .A1(n964), .A2(n1551), .B1(n964), .B2(n1543), .ZN(n652) );
  OAI22_X1 U2049 ( .A1(n1330), .A2(n966), .B1(n965), .B2(n1543), .ZN(n761) );
  OAI22_X1 U2050 ( .A1(n1551), .A2(n967), .B1(n966), .B2(n1543), .ZN(n762) );
  OAI22_X1 U2051 ( .A1(n1551), .A2(n968), .B1(n967), .B2(n1543), .ZN(n763) );
  OAI22_X1 U2052 ( .A1(n1330), .A2(n973), .B1(n972), .B2(n1543), .ZN(n768) );
  OAI22_X1 U2053 ( .A1(n1550), .A2(n972), .B1(n971), .B2(n1543), .ZN(n767) );
  OAI22_X1 U2054 ( .A1(n1551), .A2(n975), .B1(n974), .B2(n1543), .ZN(n770) );
  OAI22_X1 U2055 ( .A1(n1550), .A2(n969), .B1(n968), .B2(n1542), .ZN(n764) );
  OAI22_X1 U2056 ( .A1(n1330), .A2(n971), .B1(n970), .B2(n1543), .ZN(n766) );
  OAI22_X1 U2057 ( .A1(n1551), .A2(n978), .B1(n977), .B2(n1542), .ZN(n773) );
  OAI22_X1 U2058 ( .A1(n1330), .A2(n977), .B1(n976), .B2(n1542), .ZN(n772) );
  OAI22_X1 U2059 ( .A1(n1331), .A2(n970), .B1(n969), .B2(n1543), .ZN(n765) );
  OAI22_X1 U2060 ( .A1(n1331), .A2(n1144), .B1(n984), .B2(n1543), .ZN(n674) );
  OAI22_X1 U2061 ( .A1(n1330), .A2(n979), .B1(n978), .B2(n1542), .ZN(n774) );
  OAI22_X1 U2062 ( .A1(n1549), .A2(n976), .B1(n975), .B2(n1542), .ZN(n771) );
  OAI22_X1 U2063 ( .A1(n1550), .A2(n983), .B1(n982), .B2(n1543), .ZN(n778) );
  OAI22_X1 U2064 ( .A1(n1550), .A2(n974), .B1(n973), .B2(n1542), .ZN(n769) );
  OAI22_X1 U2065 ( .A1(n1551), .A2(n982), .B1(n1542), .B2(n981), .ZN(n777) );
  OAI22_X1 U2066 ( .A1(n1331), .A2(n980), .B1(n979), .B2(n1542), .ZN(n775) );
  OAI22_X1 U2067 ( .A1(n1331), .A2(n981), .B1(n980), .B2(n1542), .ZN(n776) );
  OAI21_X1 U2068 ( .B1(n193), .B2(n180), .A(n1372), .ZN(n179) );
  OAI21_X1 U2069 ( .B1(n181), .B2(n177), .A(n178), .ZN(n176) );
  OAI22_X1 U2070 ( .A1(n943), .A2(n42), .B1(n943), .B2(n1544), .ZN(n649) );
  OAI22_X1 U2071 ( .A1(n1264), .A2(n944), .B1(n943), .B2(n1405), .ZN(n328) );
  OAI22_X1 U2072 ( .A1(n1264), .A2(n945), .B1(n944), .B2(n1545), .ZN(n741) );
  OAI22_X1 U2073 ( .A1(n42), .A2(n947), .B1(n946), .B2(n1405), .ZN(n743) );
  OAI22_X1 U2074 ( .A1(n1264), .A2(n946), .B1(n945), .B2(n1544), .ZN(n742) );
  OAI22_X1 U2075 ( .A1(n42), .A2(n948), .B1(n947), .B2(n1405), .ZN(n744) );
  OAI22_X1 U2076 ( .A1(n1264), .A2(n949), .B1(n948), .B2(n1544), .ZN(n745) );
  OAI22_X1 U2077 ( .A1(n1485), .A2(n957), .B1(n956), .B2(n1544), .ZN(n753) );
  OAI22_X1 U2078 ( .A1(n1485), .A2(n952), .B1(n951), .B2(n1405), .ZN(n748) );
  OAI22_X1 U2079 ( .A1(n42), .A2(n1238), .B1(n952), .B2(n1405), .ZN(n749) );
  OAI22_X1 U2080 ( .A1(n1486), .A2(n956), .B1(n1324), .B2(n1545), .ZN(n752) );
  OAI22_X1 U2081 ( .A1(n42), .A2(n951), .B1(n950), .B2(n1545), .ZN(n747) );
  OAI22_X1 U2082 ( .A1(n1485), .A2(n950), .B1(n949), .B2(n1545), .ZN(n746) );
  OAI22_X1 U2083 ( .A1(n1485), .A2(n958), .B1(n957), .B2(n1405), .ZN(n754) );
  OAI22_X1 U2084 ( .A1(n1485), .A2(n1143), .B1(n963), .B2(n1405), .ZN(n673) );
  OAI22_X1 U2085 ( .A1(n1324), .A2(n1486), .B1(n954), .B2(n1545), .ZN(n751) );
  OAI22_X1 U2086 ( .A1(n1485), .A2(n961), .B1(n960), .B2(n1545), .ZN(n757) );
  OAI22_X1 U2087 ( .A1(n42), .A2(n960), .B1(n959), .B2(n1545), .ZN(n756) );
  OAI22_X1 U2088 ( .A1(n1486), .A2(n954), .B1(n953), .B2(n1545), .ZN(n750) );
  OAI22_X1 U2089 ( .A1(n1485), .A2(n962), .B1(n961), .B2(n1545), .ZN(n758) );
  OAI22_X1 U2090 ( .A1(n1486), .A2(n959), .B1(n958), .B2(n1545), .ZN(n755) );
  XNOR2_X1 U2091 ( .A(n1475), .B(n65), .ZN(product[31]) );
  XNOR2_X1 U2092 ( .A(n1497), .B(n67), .ZN(product[29]) );
  INV_X1 U2093 ( .A(n101), .ZN(n264) );
  AOI21_X1 U2094 ( .B1(n1475), .B2(n1525), .A(n111), .ZN(n109) );
  AOI21_X1 U2095 ( .B1(n1497), .B2(n1524), .A(n119), .ZN(n117) );
  OAI22_X1 U2096 ( .A1(n1349), .A2(n1014), .B1(n1013), .B2(n1344), .ZN(n807)
         );
  OAI22_X1 U2097 ( .A1(n1349), .A2(n1007), .B1(n1006), .B2(n1344), .ZN(n394)
         );
  OAI22_X1 U2098 ( .A1(n1349), .A2(n1012), .B1(n1011), .B2(n1344), .ZN(n805)
         );
  OAI22_X1 U2099 ( .A1(n1006), .A2(n1349), .B1(n1006), .B2(n1343), .ZN(n658)
         );
  OAI22_X1 U2100 ( .A1(n1349), .A2(n1024), .B1(n1023), .B2(n1343), .ZN(n817)
         );
  OAI22_X1 U2101 ( .A1(n1239), .A2(n1021), .B1(n1020), .B2(n1343), .ZN(n814)
         );
  OAI22_X1 U2102 ( .A1(n1348), .A2(n1008), .B1(n1007), .B2(n1344), .ZN(n801)
         );
  OAI22_X1 U2103 ( .A1(n1349), .A2(n1249), .B1(n1009), .B2(n1343), .ZN(n803)
         );
  OAI22_X1 U2104 ( .A1(n1349), .A2(n1009), .B1(n1008), .B2(n1344), .ZN(n802)
         );
  OAI22_X1 U2105 ( .A1(n1239), .A2(n1146), .B1(n1026), .B2(n1344), .ZN(n676)
         );
  OAI22_X1 U2106 ( .A1(n1349), .A2(n1015), .B1(n1014), .B2(n1343), .ZN(n808)
         );
  OAI22_X1 U2107 ( .A1(n1383), .A2(n1013), .B1(n1012), .B2(n1342), .ZN(n806)
         );
  OAI22_X1 U2108 ( .A1(n1349), .A2(n1025), .B1(n1024), .B2(n1344), .ZN(n818)
         );
  OAI22_X1 U2109 ( .A1(n1349), .A2(n1019), .B1(n1018), .B2(n1344), .ZN(n812)
         );
  OAI22_X1 U2110 ( .A1(n1348), .A2(n1020), .B1(n1019), .B2(n1343), .ZN(n813)
         );
  OAI22_X1 U2111 ( .A1(n1383), .A2(n1018), .B1(n1017), .B2(n1343), .ZN(n811)
         );
  OAI22_X1 U2112 ( .A1(n1349), .A2(n1023), .B1(n1022), .B2(n1343), .ZN(n816)
         );
  OAI22_X1 U2113 ( .A1(n1383), .A2(n1011), .B1(n1010), .B2(n1342), .ZN(n804)
         );
  OAI22_X1 U2114 ( .A1(n1239), .A2(n1017), .B1(n1016), .B2(n1343), .ZN(n810)
         );
  OAI22_X1 U2115 ( .A1(n1239), .A2(n1016), .B1(n1015), .B2(n1343), .ZN(n809)
         );
  OAI22_X1 U2116 ( .A1(n1383), .A2(n1022), .B1(n1021), .B2(n1343), .ZN(n815)
         );
  INV_X1 U2117 ( .A(n1342), .ZN(n659) );
  XNOR2_X1 U2118 ( .A(n1474), .B(n63), .ZN(product[33]) );
  XOR2_X1 U2119 ( .A(n109), .B(n64), .Z(product[32]) );
  XOR2_X1 U2120 ( .A(n117), .B(n66), .Z(product[30]) );
  XOR2_X1 U2121 ( .A(n125), .B(n68), .Z(product[28]) );
  AOI21_X1 U2122 ( .B1(n106), .B2(n1523), .A(n103), .ZN(n101) );
  OAI21_X1 U2123 ( .B1(n1500), .B2(n115), .A(n116), .ZN(n114) );
  OAI21_X1 U2124 ( .B1(n1517), .B2(n123), .A(n124), .ZN(n122) );
  OAI22_X1 U2125 ( .A1(n1261), .A2(n1039), .B1(n1038), .B2(n1496), .ZN(n831)
         );
  OAI22_X1 U2126 ( .A1(n1261), .A2(n1031), .B1(n1030), .B2(n1496), .ZN(n823)
         );
  OAI22_X1 U2127 ( .A1(n1262), .A2(n1041), .B1(n1040), .B2(n1496), .ZN(n833)
         );
  OAI22_X1 U2128 ( .A1(n1261), .A2(n1032), .B1(n1031), .B2(n1494), .ZN(n824)
         );
  OAI22_X1 U2129 ( .A1(n1261), .A2(n1034), .B1(n1033), .B2(n1496), .ZN(n826)
         );
  OAI22_X1 U2130 ( .A1(n1261), .A2(n1045), .B1(n1044), .B2(n1494), .ZN(n837)
         );
  OAI22_X1 U2131 ( .A1(n1262), .A2(n1038), .B1(n1037), .B2(n1496), .ZN(n830)
         );
  OAI22_X1 U2132 ( .A1(n1261), .A2(n1044), .B1(n1043), .B2(n1494), .ZN(n836)
         );
  OAI22_X1 U2133 ( .A1(n1262), .A2(n1040), .B1(n1039), .B2(n1496), .ZN(n832)
         );
  OAI22_X1 U2134 ( .A1(n1261), .A2(n1028), .B1(n1027), .B2(n1495), .ZN(n424)
         );
  OAI22_X1 U2135 ( .A1(n1261), .A2(n1037), .B1(n1496), .B2(n1036), .ZN(n829)
         );
  OAI22_X1 U2136 ( .A1(n1367), .A2(n1030), .B1(n1029), .B2(n1495), .ZN(n822)
         );
  OAI22_X1 U2137 ( .A1(n1261), .A2(n1033), .B1(n1032), .B2(n1496), .ZN(n825)
         );
  OAI22_X1 U2138 ( .A1(n1262), .A2(n1147), .B1(n1047), .B2(n1494), .ZN(n677)
         );
  OAI22_X1 U2139 ( .A1(n1027), .A2(n1261), .B1(n1027), .B2(n1495), .ZN(n661)
         );
  OAI22_X1 U2140 ( .A1(n1262), .A2(n1043), .B1(n1042), .B2(n1494), .ZN(n835)
         );
  OAI22_X1 U2141 ( .A1(n1367), .A2(n1029), .B1(n1028), .B2(n1495), .ZN(n821)
         );
  OAI22_X1 U2142 ( .A1(n1262), .A2(n1036), .B1(n1035), .B2(n1495), .ZN(n828)
         );
  OAI22_X1 U2143 ( .A1(n1262), .A2(n1042), .B1(n1041), .B2(n1496), .ZN(n834)
         );
  OAI22_X1 U2144 ( .A1(n1262), .A2(n1035), .B1(n1034), .B2(n1496), .ZN(n827)
         );
  OAI22_X1 U2145 ( .A1(n1262), .A2(n1046), .B1(n1045), .B2(n1494), .ZN(n838)
         );
  INV_X1 U2146 ( .A(n1496), .ZN(n662) );
  OAI21_X1 U2147 ( .B1(n1493), .B2(n107), .A(n108), .ZN(n106) );
endmodule


module mac_2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n34, n35, n36, n37, n38, n39, n40, n41, n43, n45, n46, n47,
         n48, n49, n51, n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65,
         n67, n69, n70, n71, n72, n73, n75, n77, n78, n79, n80, n81, n83, n85,
         n86, n87, n88, n89, n91, n93, n94, n95, n96, n97, n99, n101, n102,
         n103, n104, n105, n107, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n119, n121, n122, n124, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n184, n185, n187, n189, n191,
         n193, n195, n197, n199, n201, n203, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409;

  FA_X1 U7 ( .A(B[34]), .B(A[34]), .CI(n39), .CO(n38), .S(SUM[34]) );
  FA_X1 U8 ( .A(B[33]), .B(A[33]), .CI(n40), .CO(n39), .S(SUM[33]) );
  FA_X1 U9 ( .A(B[32]), .B(A[32]), .CI(n185), .CO(n40), .S(SUM[32]) );
  OR2_X1 U254 ( .A1(B[12]), .A2(A[12]), .ZN(n398) );
  NAND2_X1 U255 ( .A1(B[8]), .A2(A[8]), .ZN(n148) );
  OR2_X1 U256 ( .A1(B[0]), .A2(A[0]), .ZN(n344) );
  NAND3_X1 U257 ( .A1(n349), .A2(n350), .A3(n351), .ZN(n345) );
  NAND3_X1 U258 ( .A1(n349), .A2(n350), .A3(n351), .ZN(n346) );
  NAND3_X1 U259 ( .A1(n355), .A2(n356), .A3(n357), .ZN(n347) );
  XOR2_X1 U260 ( .A(B[35]), .B(A[35]), .Z(n348) );
  XOR2_X1 U261 ( .A(n38), .B(n348), .Z(SUM[35]) );
  NAND2_X1 U262 ( .A1(n38), .A2(B[35]), .ZN(n349) );
  NAND2_X1 U263 ( .A1(n38), .A2(A[35]), .ZN(n350) );
  NAND2_X1 U264 ( .A1(B[35]), .A2(A[35]), .ZN(n351) );
  NAND3_X1 U265 ( .A1(n349), .A2(n350), .A3(n351), .ZN(n37) );
  AOI21_X1 U266 ( .B1(n172), .B2(n180), .A(n173), .ZN(n352) );
  NOR2_X1 U267 ( .A1(B[9]), .A2(A[9]), .ZN(n353) );
  NOR2_X1 U268 ( .A1(B[9]), .A2(A[9]), .ZN(n144) );
  XOR2_X1 U269 ( .A(B[36]), .B(A[36]), .Z(n354) );
  XOR2_X1 U270 ( .A(n346), .B(n354), .Z(SUM[36]) );
  NAND2_X1 U271 ( .A1(n345), .A2(B[36]), .ZN(n355) );
  NAND2_X1 U272 ( .A1(n37), .A2(A[36]), .ZN(n356) );
  NAND2_X1 U273 ( .A1(B[36]), .A2(A[36]), .ZN(n357) );
  NAND3_X1 U274 ( .A1(n355), .A2(n356), .A3(n357), .ZN(n36) );
  CLKBUF_X1 U275 ( .A(n78), .Z(n358) );
  CLKBUF_X1 U276 ( .A(n62), .Z(n359) );
  CLKBUF_X1 U277 ( .A(n130), .Z(n360) );
  NOR2_X1 U278 ( .A1(B[5]), .A2(A[5]), .ZN(n361) );
  NOR2_X1 U279 ( .A1(B[7]), .A2(A[7]), .ZN(n362) );
  CLKBUF_X1 U280 ( .A(n143), .Z(n363) );
  NOR2_X1 U281 ( .A1(B[11]), .A2(A[11]), .ZN(n364) );
  NOR2_X1 U282 ( .A1(B[11]), .A2(A[11]), .ZN(n132) );
  CLKBUF_X1 U283 ( .A(n36), .Z(n365) );
  AOI21_X1 U284 ( .B1(n358), .B2(n404), .A(n75), .ZN(n366) );
  AOI21_X1 U285 ( .B1(n78), .B2(n404), .A(n75), .ZN(n73) );
  AOI21_X1 U286 ( .B1(n359), .B2(n406), .A(n59), .ZN(n367) );
  AOI21_X1 U287 ( .B1(n62), .B2(n406), .A(n59), .ZN(n57) );
  NOR2_X1 U288 ( .A1(B[3]), .A2(A[3]), .ZN(n368) );
  CLKBUF_X1 U289 ( .A(n131), .Z(n369) );
  CLKBUF_X1 U290 ( .A(n115), .Z(n370) );
  CLKBUF_X1 U291 ( .A(n150), .Z(n371) );
  AOI21_X1 U292 ( .B1(n360), .B2(n363), .A(n369), .ZN(n372) );
  CLKBUF_X1 U293 ( .A(n110), .Z(n373) );
  CLKBUF_X1 U294 ( .A(n86), .Z(n374) );
  BUF_X1 U295 ( .A(n383), .Z(n375) );
  AOI21_X1 U296 ( .B1(n371), .B2(n114), .A(n370), .ZN(n376) );
  AOI21_X1 U297 ( .B1(n150), .B2(n114), .A(n115), .ZN(n113) );
  NAND3_X1 U298 ( .A1(n382), .A2(n375), .A3(n384), .ZN(n377) );
  CLKBUF_X1 U299 ( .A(n54), .Z(n378) );
  CLKBUF_X1 U300 ( .A(n94), .Z(n379) );
  CLKBUF_X1 U301 ( .A(n70), .Z(n380) );
  XOR2_X1 U302 ( .A(B[37]), .B(A[37]), .Z(n381) );
  XOR2_X1 U303 ( .A(n381), .B(n365), .Z(SUM[37]) );
  NAND2_X1 U304 ( .A1(B[37]), .A2(A[37]), .ZN(n382) );
  NAND2_X1 U305 ( .A1(n36), .A2(B[37]), .ZN(n383) );
  NAND2_X1 U306 ( .A1(n347), .A2(A[37]), .ZN(n384) );
  NAND3_X1 U307 ( .A1(n384), .A2(n383), .A3(n382), .ZN(n35) );
  XOR2_X1 U308 ( .A(B[38]), .B(A[38]), .Z(n385) );
  XOR2_X1 U309 ( .A(n385), .B(n377), .Z(SUM[38]) );
  NAND2_X1 U310 ( .A1(B[38]), .A2(A[38]), .ZN(n386) );
  NAND2_X1 U311 ( .A1(n35), .A2(B[38]), .ZN(n387) );
  NAND2_X1 U312 ( .A1(n35), .A2(A[38]), .ZN(n388) );
  NAND3_X1 U313 ( .A1(n386), .A2(n387), .A3(n388), .ZN(n34) );
  AOI21_X1 U314 ( .B1(n374), .B2(n402), .A(n83), .ZN(n389) );
  AOI21_X1 U315 ( .B1(n86), .B2(n402), .A(n83), .ZN(n81) );
  AOI21_X1 U316 ( .B1(n393), .B2(n400), .A(n99), .ZN(n390) );
  CLKBUF_X1 U317 ( .A(n46), .Z(n391) );
  AOI21_X1 U318 ( .B1(n378), .B2(n407), .A(n51), .ZN(n392) );
  CLKBUF_X1 U319 ( .A(n102), .Z(n393) );
  AOI21_X1 U320 ( .B1(n102), .B2(n400), .A(n99), .ZN(n97) );
  AOI21_X1 U321 ( .B1(n380), .B2(n405), .A(n67), .ZN(n394) );
  AOI21_X1 U322 ( .B1(n373), .B2(n401), .A(n107), .ZN(n395) );
  AOI21_X1 U323 ( .B1(n379), .B2(n403), .A(n91), .ZN(n396) );
  NOR2_X1 U324 ( .A1(B[7]), .A2(A[7]), .ZN(n155) );
  NOR2_X1 U325 ( .A1(B[5]), .A2(A[5]), .ZN(n163) );
  NOR2_X1 U326 ( .A1(B[8]), .A2(A[8]), .ZN(n147) );
  NOR2_X1 U327 ( .A1(B[6]), .A2(A[6]), .ZN(n158) );
  NOR2_X1 U328 ( .A1(B[10]), .A2(A[10]), .ZN(n137) );
  NAND2_X1 U329 ( .A1(B[10]), .A2(A[10]), .ZN(n138) );
  OR2_X1 U330 ( .A1(B[17]), .A2(A[17]), .ZN(n400) );
  OAI21_X1 U331 ( .B1(n149), .B2(n140), .A(n141), .ZN(n139) );
  INV_X1 U332 ( .A(n363), .ZN(n141) );
  INV_X1 U333 ( .A(n142), .ZN(n140) );
  NAND2_X1 U334 ( .A1(n142), .A2(n130), .ZN(n128) );
  AOI21_X1 U335 ( .B1(n170), .B2(n161), .A(n162), .ZN(n160) );
  INV_X1 U336 ( .A(n352), .ZN(n170) );
  INV_X1 U337 ( .A(n180), .ZN(n179) );
  INV_X1 U338 ( .A(n101), .ZN(n99) );
  INV_X1 U339 ( .A(n85), .ZN(n83) );
  INV_X1 U340 ( .A(n77), .ZN(n75) );
  INV_X1 U341 ( .A(n69), .ZN(n67) );
  INV_X1 U342 ( .A(n61), .ZN(n59) );
  INV_X1 U343 ( .A(n53), .ZN(n51) );
  NAND2_X1 U344 ( .A1(n161), .A2(n153), .ZN(n151) );
  AOI21_X1 U345 ( .B1(n153), .B2(n162), .A(n154), .ZN(n152) );
  NOR2_X1 U346 ( .A1(n158), .A2(n362), .ZN(n153) );
  OAI21_X1 U347 ( .B1(n163), .B2(n169), .A(n164), .ZN(n162) );
  AOI21_X1 U348 ( .B1(n110), .B2(n401), .A(n107), .ZN(n105) );
  INV_X1 U349 ( .A(n109), .ZN(n107) );
  OAI21_X1 U350 ( .B1(n97), .B2(n95), .A(n96), .ZN(n94) );
  OAI21_X1 U351 ( .B1(n144), .B2(n148), .A(n145), .ZN(n143) );
  NOR2_X1 U352 ( .A1(n168), .A2(n361), .ZN(n161) );
  OAI21_X1 U353 ( .B1(n181), .B2(n184), .A(n182), .ZN(n180) );
  NOR2_X1 U354 ( .A1(n137), .A2(n364), .ZN(n130) );
  AOI21_X1 U355 ( .B1(n94), .B2(n403), .A(n91), .ZN(n89) );
  INV_X1 U356 ( .A(n93), .ZN(n91) );
  AOI21_X1 U357 ( .B1(n172), .B2(n180), .A(n173), .ZN(n171) );
  NOR2_X1 U358 ( .A1(n177), .A2(n368), .ZN(n172) );
  OAI21_X1 U359 ( .B1(n174), .B2(n178), .A(n175), .ZN(n173) );
  NOR2_X1 U360 ( .A1(n128), .A2(n116), .ZN(n114) );
  NAND2_X1 U361 ( .A1(n398), .A2(n399), .ZN(n116) );
  NAND2_X1 U362 ( .A1(n195), .A2(n80), .ZN(n11) );
  INV_X1 U363 ( .A(n79), .ZN(n195) );
  NOR2_X1 U364 ( .A1(n147), .A2(n353), .ZN(n142) );
  AOI21_X1 U365 ( .B1(n130), .B2(n143), .A(n131), .ZN(n129) );
  OAI21_X1 U366 ( .B1(n132), .B2(n138), .A(n133), .ZN(n131) );
  INV_X1 U367 ( .A(n126), .ZN(n124) );
  OAI21_X1 U368 ( .B1(n155), .B2(n159), .A(n156), .ZN(n154) );
  XOR2_X1 U369 ( .A(n396), .B(n13), .Z(SUM[20]) );
  NAND2_X1 U370 ( .A1(n197), .A2(n88), .ZN(n13) );
  INV_X1 U371 ( .A(n87), .ZN(n197) );
  XOR2_X1 U372 ( .A(n390), .B(n15), .Z(SUM[18]) );
  NAND2_X1 U373 ( .A1(n199), .A2(n96), .ZN(n15) );
  INV_X1 U374 ( .A(n95), .ZN(n199) );
  AOI21_X1 U375 ( .B1(n399), .B2(n124), .A(n119), .ZN(n117) );
  INV_X1 U376 ( .A(n121), .ZN(n119) );
  NAND2_X1 U377 ( .A1(n187), .A2(n48), .ZN(n3) );
  INV_X1 U378 ( .A(n47), .ZN(n187) );
  NAND2_X1 U379 ( .A1(n189), .A2(n56), .ZN(n5) );
  INV_X1 U380 ( .A(n55), .ZN(n189) );
  NAND2_X1 U381 ( .A1(n191), .A2(n64), .ZN(n7) );
  INV_X1 U382 ( .A(n63), .ZN(n191) );
  NAND2_X1 U383 ( .A1(n193), .A2(n72), .ZN(n9) );
  INV_X1 U384 ( .A(n71), .ZN(n193) );
  NAND2_X1 U385 ( .A1(n408), .A2(n45), .ZN(n2) );
  NAND2_X1 U386 ( .A1(n407), .A2(n53), .ZN(n4) );
  NAND2_X1 U387 ( .A1(n406), .A2(n61), .ZN(n6) );
  NAND2_X1 U388 ( .A1(n405), .A2(n69), .ZN(n8) );
  NAND2_X1 U389 ( .A1(n404), .A2(n77), .ZN(n10) );
  NAND2_X1 U390 ( .A1(n402), .A2(n85), .ZN(n12) );
  XNOR2_X1 U391 ( .A(n379), .B(n14), .ZN(SUM[19]) );
  NAND2_X1 U392 ( .A1(n403), .A2(n93), .ZN(n14) );
  NAND2_X1 U393 ( .A1(n400), .A2(n101), .ZN(n16) );
  XOR2_X1 U394 ( .A(n122), .B(n20), .Z(SUM[13]) );
  NAND2_X1 U395 ( .A1(n399), .A2(n121), .ZN(n20) );
  AOI21_X1 U396 ( .B1(n127), .B2(n398), .A(n124), .ZN(n122) );
  XOR2_X1 U397 ( .A(n134), .B(n22), .Z(SUM[11]) );
  NAND2_X1 U398 ( .A1(n206), .A2(n133), .ZN(n22) );
  AOI21_X1 U399 ( .B1(n139), .B2(n207), .A(n136), .ZN(n134) );
  NAND2_X1 U400 ( .A1(n201), .A2(n104), .ZN(n17) );
  INV_X1 U401 ( .A(n103), .ZN(n201) );
  INV_X1 U402 ( .A(n137), .ZN(n207) );
  INV_X1 U403 ( .A(n168), .ZN(n213) );
  XOR2_X1 U404 ( .A(n160), .B(n27), .Z(SUM[6]) );
  NAND2_X1 U405 ( .A1(n211), .A2(n159), .ZN(n27) );
  INV_X1 U406 ( .A(n158), .ZN(n211) );
  INV_X1 U407 ( .A(n364), .ZN(n206) );
  INV_X1 U408 ( .A(n138), .ZN(n136) );
  INV_X1 U409 ( .A(n169), .ZN(n167) );
  INV_X1 U410 ( .A(n353), .ZN(n208) );
  INV_X1 U411 ( .A(n362), .ZN(n210) );
  INV_X1 U412 ( .A(n361), .ZN(n212) );
  INV_X1 U413 ( .A(n368), .ZN(n214) );
  XOR2_X1 U414 ( .A(n165), .B(n28), .Z(SUM[5]) );
  NAND2_X1 U415 ( .A1(n212), .A2(n164), .ZN(n28) );
  AOI21_X1 U416 ( .B1(n170), .B2(n213), .A(n167), .ZN(n165) );
  XNOR2_X1 U417 ( .A(n170), .B(n29), .ZN(SUM[4]) );
  NAND2_X1 U418 ( .A1(n213), .A2(n169), .ZN(n29) );
  XNOR2_X1 U419 ( .A(n176), .B(n30), .ZN(SUM[3]) );
  NAND2_X1 U420 ( .A1(n214), .A2(n175), .ZN(n30) );
  OAI21_X1 U421 ( .B1(n179), .B2(n177), .A(n178), .ZN(n176) );
  XOR2_X1 U422 ( .A(n179), .B(n31), .Z(SUM[2]) );
  NAND2_X1 U423 ( .A1(n215), .A2(n178), .ZN(n31) );
  INV_X1 U424 ( .A(n177), .ZN(n215) );
  XOR2_X1 U425 ( .A(n32), .B(n184), .Z(SUM[1]) );
  NAND2_X1 U426 ( .A1(n216), .A2(n182), .ZN(n32) );
  INV_X1 U427 ( .A(n181), .ZN(n216) );
  AND2_X1 U428 ( .A1(n344), .A2(n184), .ZN(SUM[0]) );
  NAND2_X1 U429 ( .A1(n203), .A2(n112), .ZN(n19) );
  INV_X1 U430 ( .A(n111), .ZN(n203) );
  NAND2_X1 U431 ( .A1(n401), .A2(n109), .ZN(n18) );
  XNOR2_X1 U432 ( .A(n127), .B(n21), .ZN(SUM[12]) );
  NAND2_X1 U433 ( .A1(n398), .A2(n126), .ZN(n21) );
  XNOR2_X1 U434 ( .A(n139), .B(n23), .ZN(SUM[10]) );
  NAND2_X1 U435 ( .A1(n207), .A2(n138), .ZN(n23) );
  XNOR2_X1 U436 ( .A(n146), .B(n24), .ZN(SUM[9]) );
  NAND2_X1 U437 ( .A1(n208), .A2(n145), .ZN(n24) );
  OAI21_X1 U438 ( .B1(n149), .B2(n147), .A(n148), .ZN(n146) );
  XOR2_X1 U439 ( .A(n149), .B(n25), .Z(SUM[8]) );
  NAND2_X1 U440 ( .A1(n209), .A2(n148), .ZN(n25) );
  INV_X1 U441 ( .A(n147), .ZN(n209) );
  XNOR2_X1 U442 ( .A(n157), .B(n26), .ZN(SUM[7]) );
  NAND2_X1 U443 ( .A1(n210), .A2(n156), .ZN(n26) );
  OAI21_X1 U444 ( .B1(n160), .B2(n158), .A(n159), .ZN(n157) );
  NOR2_X1 U445 ( .A1(B[2]), .A2(A[2]), .ZN(n177) );
  NOR2_X1 U446 ( .A1(B[3]), .A2(A[3]), .ZN(n174) );
  OR2_X2 U447 ( .A1(B[13]), .A2(A[13]), .ZN(n399) );
  NAND2_X1 U448 ( .A1(B[11]), .A2(A[11]), .ZN(n133) );
  NOR2_X1 U449 ( .A1(B[4]), .A2(A[4]), .ZN(n168) );
  NOR2_X1 U450 ( .A1(B[18]), .A2(A[18]), .ZN(n95) );
  NOR2_X1 U451 ( .A1(B[1]), .A2(A[1]), .ZN(n181) );
  NAND2_X1 U452 ( .A1(B[6]), .A2(A[6]), .ZN(n159) );
  NAND2_X1 U453 ( .A1(B[2]), .A2(A[2]), .ZN(n178) );
  NAND2_X1 U454 ( .A1(B[0]), .A2(A[0]), .ZN(n184) );
  NAND2_X1 U455 ( .A1(B[4]), .A2(A[4]), .ZN(n169) );
  NAND2_X1 U456 ( .A1(B[9]), .A2(A[9]), .ZN(n145) );
  NAND2_X1 U457 ( .A1(B[5]), .A2(A[5]), .ZN(n164) );
  NAND2_X1 U458 ( .A1(B[7]), .A2(A[7]), .ZN(n156) );
  NAND2_X1 U459 ( .A1(B[3]), .A2(A[3]), .ZN(n175) );
  NAND2_X1 U460 ( .A1(B[1]), .A2(A[1]), .ZN(n182) );
  NAND2_X1 U461 ( .A1(B[18]), .A2(A[18]), .ZN(n96) );
  INV_X1 U462 ( .A(n45), .ZN(n43) );
  NOR2_X1 U463 ( .A1(B[14]), .A2(A[14]), .ZN(n111) );
  NOR2_X1 U464 ( .A1(B[20]), .A2(A[20]), .ZN(n87) );
  NOR2_X1 U465 ( .A1(B[16]), .A2(A[16]), .ZN(n103) );
  NOR2_X1 U466 ( .A1(B[30]), .A2(A[30]), .ZN(n47) );
  NOR2_X1 U467 ( .A1(B[28]), .A2(A[28]), .ZN(n55) );
  NOR2_X1 U468 ( .A1(B[26]), .A2(A[26]), .ZN(n63) );
  NOR2_X1 U469 ( .A1(B[24]), .A2(A[24]), .ZN(n71) );
  NOR2_X1 U470 ( .A1(B[22]), .A2(A[22]), .ZN(n79) );
  OR2_X1 U471 ( .A1(B[15]), .A2(A[15]), .ZN(n401) );
  NAND2_X1 U472 ( .A1(B[21]), .A2(A[21]), .ZN(n85) );
  NAND2_X1 U473 ( .A1(B[12]), .A2(A[12]), .ZN(n126) );
  NAND2_X1 U474 ( .A1(B[13]), .A2(A[13]), .ZN(n121) );
  NAND2_X1 U475 ( .A1(B[19]), .A2(A[19]), .ZN(n93) );
  NAND2_X1 U476 ( .A1(B[17]), .A2(A[17]), .ZN(n101) );
  NAND2_X1 U477 ( .A1(B[15]), .A2(A[15]), .ZN(n109) );
  NAND2_X1 U478 ( .A1(B[23]), .A2(A[23]), .ZN(n77) );
  NAND2_X1 U479 ( .A1(B[25]), .A2(A[25]), .ZN(n69) );
  NAND2_X1 U480 ( .A1(B[27]), .A2(A[27]), .ZN(n61) );
  NAND2_X1 U481 ( .A1(B[29]), .A2(A[29]), .ZN(n53) );
  NAND2_X1 U482 ( .A1(B[31]), .A2(A[31]), .ZN(n45) );
  NAND2_X1 U483 ( .A1(B[14]), .A2(A[14]), .ZN(n112) );
  NAND2_X1 U484 ( .A1(B[20]), .A2(A[20]), .ZN(n88) );
  NAND2_X1 U485 ( .A1(B[16]), .A2(A[16]), .ZN(n104) );
  NAND2_X1 U486 ( .A1(B[30]), .A2(A[30]), .ZN(n48) );
  NAND2_X1 U487 ( .A1(B[28]), .A2(A[28]), .ZN(n56) );
  NAND2_X1 U488 ( .A1(B[26]), .A2(A[26]), .ZN(n64) );
  NAND2_X1 U489 ( .A1(B[24]), .A2(A[24]), .ZN(n72) );
  NAND2_X1 U490 ( .A1(B[22]), .A2(A[22]), .ZN(n80) );
  OR2_X1 U491 ( .A1(B[21]), .A2(A[21]), .ZN(n402) );
  OR2_X1 U492 ( .A1(B[19]), .A2(A[19]), .ZN(n403) );
  OR2_X1 U493 ( .A1(B[23]), .A2(A[23]), .ZN(n404) );
  OR2_X1 U494 ( .A1(B[25]), .A2(A[25]), .ZN(n405) );
  OR2_X1 U495 ( .A1(B[27]), .A2(A[27]), .ZN(n406) );
  OR2_X1 U496 ( .A1(B[29]), .A2(A[29]), .ZN(n407) );
  OR2_X1 U497 ( .A1(B[31]), .A2(A[31]), .ZN(n408) );
  XNOR2_X1 U498 ( .A(n34), .B(n409), .ZN(SUM[39]) );
  XNOR2_X1 U499 ( .A(A[39]), .B(B[39]), .ZN(n409) );
  XNOR2_X1 U500 ( .A(n393), .B(n16), .ZN(SUM[17]) );
  OAI21_X1 U501 ( .B1(n105), .B2(n103), .A(n104), .ZN(n102) );
  XOR2_X1 U502 ( .A(n395), .B(n17), .Z(SUM[16]) );
  XNOR2_X1 U503 ( .A(n380), .B(n8), .ZN(SUM[25]) );
  AOI21_X1 U504 ( .B1(n70), .B2(n405), .A(n67), .ZN(n65) );
  XNOR2_X1 U505 ( .A(n359), .B(n6), .ZN(SUM[27]) );
  XNOR2_X1 U506 ( .A(n373), .B(n18), .ZN(SUM[15]) );
  XNOR2_X1 U507 ( .A(n378), .B(n4), .ZN(SUM[29]) );
  AOI21_X1 U508 ( .B1(n54), .B2(n407), .A(n51), .ZN(n49) );
  XNOR2_X1 U509 ( .A(n391), .B(n2), .ZN(SUM[31]) );
  XNOR2_X1 U510 ( .A(n358), .B(n10), .ZN(SUM[23]) );
  XOR2_X1 U511 ( .A(n392), .B(n3), .Z(SUM[30]) );
  XOR2_X1 U512 ( .A(n367), .B(n5), .Z(SUM[28]) );
  AOI21_X1 U513 ( .B1(n46), .B2(n408), .A(n43), .ZN(n41) );
  OAI21_X1 U514 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  OAI21_X1 U515 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  XNOR2_X1 U516 ( .A(n374), .B(n12), .ZN(SUM[21]) );
  XOR2_X1 U517 ( .A(n376), .B(n19), .Z(SUM[14]) );
  XOR2_X1 U518 ( .A(n389), .B(n11), .Z(SUM[22]) );
  INV_X1 U519 ( .A(n371), .ZN(n149) );
  INV_X1 U520 ( .A(n41), .ZN(n185) );
  OAI21_X1 U521 ( .B1(n81), .B2(n79), .A(n80), .ZN(n78) );
  OAI21_X1 U522 ( .B1(n113), .B2(n111), .A(n112), .ZN(n110) );
  OAI21_X1 U523 ( .B1(n171), .B2(n151), .A(n152), .ZN(n150) );
  OAI21_X1 U524 ( .B1(n89), .B2(n87), .A(n88), .ZN(n86) );
  XOR2_X1 U525 ( .A(n394), .B(n7), .Z(SUM[26]) );
  XOR2_X1 U526 ( .A(n366), .B(n9), .Z(SUM[24]) );
  OAI21_X1 U527 ( .B1(n149), .B2(n128), .A(n372), .ZN(n127) );
  OAI21_X1 U528 ( .B1(n65), .B2(n63), .A(n64), .ZN(n62) );
  OAI21_X1 U529 ( .B1(n73), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U530 ( .B1(n129), .B2(n116), .A(n117), .ZN(n115) );
endmodule


module mac_2 ( clk, clear_acc, a, b, mac_out );
  input [19:0] a;
  input [19:0] b;
  output [39:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, n2, n3;
  wire   [39:0] mul;
  wire   [39:0] pipeline;
  wire   [39:0] sum;

  DFF_X1 \pipeline_reg[37]  ( .D(mul[37]), .CK(clk), .Q(pipeline[37]) );
  DFF_X1 \pipeline_reg[36]  ( .D(mul[36]), .CK(clk), .Q(pipeline[36]) );
  DFF_X1 \pipeline_reg[35]  ( .D(mul[35]), .CK(clk), .Q(pipeline[35]) );
  DFF_X1 \pipeline_reg[34]  ( .D(mul[34]), .CK(clk), .Q(pipeline[34]) );
  DFF_X1 \pipeline_reg[33]  ( .D(mul[33]), .CK(clk), .Q(pipeline[33]) );
  DFF_X1 \pipeline_reg[32]  ( .D(mul[32]), .CK(clk), .Q(pipeline[32]) );
  DFF_X1 \pipeline_reg[31]  ( .D(mul[31]), .CK(clk), .Q(pipeline[31]) );
  DFF_X1 \pipeline_reg[30]  ( .D(mul[30]), .CK(clk), .Q(pipeline[30]) );
  DFF_X1 \pipeline_reg[29]  ( .D(mul[29]), .CK(clk), .Q(pipeline[29]) );
  DFF_X1 \pipeline_reg[28]  ( .D(mul[28]), .CK(clk), .Q(pipeline[28]) );
  DFF_X1 \pipeline_reg[27]  ( .D(mul[27]), .CK(clk), .Q(pipeline[27]) );
  DFF_X1 \pipeline_reg[26]  ( .D(mul[26]), .CK(clk), .Q(pipeline[26]) );
  DFF_X1 \pipeline_reg[25]  ( .D(mul[25]), .CK(clk), .Q(pipeline[25]) );
  DFF_X1 \pipeline_reg[24]  ( .D(mul[24]), .CK(clk), .Q(pipeline[24]) );
  DFF_X1 \pipeline_reg[23]  ( .D(mul[23]), .CK(clk), .Q(pipeline[23]) );
  DFF_X1 \pipeline_reg[22]  ( .D(mul[22]), .CK(clk), .Q(pipeline[22]) );
  DFF_X1 \pipeline_reg[21]  ( .D(mul[21]), .CK(clk), .Q(pipeline[21]) );
  DFF_X1 \pipeline_reg[20]  ( .D(mul[20]), .CK(clk), .Q(pipeline[20]) );
  DFF_X1 \pipeline_reg[19]  ( .D(mul[19]), .CK(clk), .Q(pipeline[19]) );
  DFF_X1 \pipeline_reg[18]  ( .D(mul[18]), .CK(clk), .Q(pipeline[18]) );
  DFF_X1 \pipeline_reg[17]  ( .D(mul[17]), .CK(clk), .Q(pipeline[17]) );
  DFF_X1 \pipeline_reg[16]  ( .D(mul[16]), .CK(clk), .Q(pipeline[16]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \mac_out_reg[16]  ( .D(N19), .CK(clk), .Q(mac_out[16]) );
  DFF_X1 \mac_out_reg[17]  ( .D(N20), .CK(clk), .Q(mac_out[17]) );
  DFF_X1 \mac_out_reg[18]  ( .D(N21), .CK(clk), .Q(mac_out[18]) );
  DFF_X1 \mac_out_reg[19]  ( .D(N22), .CK(clk), .Q(mac_out[19]) );
  DFF_X1 \mac_out_reg[20]  ( .D(N23), .CK(clk), .Q(mac_out[20]) );
  DFF_X1 \mac_out_reg[21]  ( .D(N24), .CK(clk), .Q(mac_out[21]) );
  DFF_X1 \mac_out_reg[22]  ( .D(N25), .CK(clk), .Q(mac_out[22]) );
  DFF_X1 \mac_out_reg[23]  ( .D(N26), .CK(clk), .Q(mac_out[23]) );
  DFF_X1 \mac_out_reg[24]  ( .D(N27), .CK(clk), .Q(mac_out[24]) );
  DFF_X1 \mac_out_reg[25]  ( .D(N28), .CK(clk), .Q(mac_out[25]) );
  DFF_X1 \mac_out_reg[26]  ( .D(N29), .CK(clk), .Q(mac_out[26]) );
  DFF_X1 \mac_out_reg[27]  ( .D(N30), .CK(clk), .Q(mac_out[27]) );
  DFF_X1 \mac_out_reg[28]  ( .D(N31), .CK(clk), .Q(mac_out[28]) );
  DFF_X1 \mac_out_reg[29]  ( .D(N32), .CK(clk), .Q(mac_out[29]) );
  DFF_X1 \mac_out_reg[30]  ( .D(N33), .CK(clk), .Q(mac_out[30]) );
  DFF_X1 \mac_out_reg[31]  ( .D(N34), .CK(clk), .Q(mac_out[31]) );
  DFF_X1 \mac_out_reg[32]  ( .D(N35), .CK(clk), .Q(mac_out[32]) );
  DFF_X1 \mac_out_reg[33]  ( .D(N36), .CK(clk), .Q(mac_out[33]) );
  DFF_X1 \mac_out_reg[34]  ( .D(N37), .CK(clk), .Q(mac_out[34]) );
  DFF_X1 \mac_out_reg[35]  ( .D(N38), .CK(clk), .Q(mac_out[35]) );
  DFF_X1 \mac_out_reg[36]  ( .D(N39), .CK(clk), .Q(mac_out[36]) );
  DFF_X1 \mac_out_reg[37]  ( .D(N40), .CK(clk), .Q(mac_out[37]) );
  DFF_X1 \mac_out_reg[38]  ( .D(N41), .CK(clk), .Q(mac_out[38]) );
  DFF_X1 \mac_out_reg[39]  ( .D(N42), .CK(clk), .Q(mac_out[39]) );
  mac_2_DW_mult_tc_1 mult_355 ( .a(a), .b(b), .product(mul) );
  mac_2_DW01_add_1 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  DFF_X2 \pipeline_reg[39]  ( .D(mul[39]), .CK(clk), .Q(pipeline[39]) );
  DFF_X1 \pipeline_reg[38]  ( .D(mul[38]), .CK(clk), .Q(pipeline[38]) );
  BUF_X1 U3 ( .A(n3), .Z(n2) );
  INV_X1 U4 ( .A(clear_acc), .ZN(n3) );
  AND2_X1 U6 ( .A1(sum[39]), .A2(n2), .ZN(N42) );
  AND2_X1 U7 ( .A1(sum[38]), .A2(n2), .ZN(N41) );
  AND2_X1 U8 ( .A1(sum[37]), .A2(n2), .ZN(N40) );
  AND2_X1 U9 ( .A1(sum[36]), .A2(n2), .ZN(N39) );
  AND2_X1 U10 ( .A1(sum[35]), .A2(n2), .ZN(N38) );
  AND2_X1 U11 ( .A1(sum[34]), .A2(n2), .ZN(N37) );
  AND2_X1 U12 ( .A1(sum[33]), .A2(n2), .ZN(N36) );
  AND2_X1 U13 ( .A1(sum[32]), .A2(n2), .ZN(N35) );
  AND2_X1 U14 ( .A1(sum[31]), .A2(n2), .ZN(N34) );
  AND2_X1 U15 ( .A1(sum[30]), .A2(n2), .ZN(N33) );
  AND2_X1 U16 ( .A1(sum[29]), .A2(n2), .ZN(N32) );
  AND2_X1 U17 ( .A1(sum[28]), .A2(n3), .ZN(N31) );
  AND2_X1 U18 ( .A1(sum[27]), .A2(n3), .ZN(N30) );
  AND2_X1 U19 ( .A1(sum[26]), .A2(n3), .ZN(N29) );
  AND2_X1 U20 ( .A1(sum[25]), .A2(n3), .ZN(N28) );
  AND2_X1 U21 ( .A1(sum[24]), .A2(n3), .ZN(N27) );
  AND2_X1 U22 ( .A1(sum[23]), .A2(n3), .ZN(N26) );
  AND2_X1 U23 ( .A1(sum[22]), .A2(n3), .ZN(N25) );
  AND2_X1 U24 ( .A1(sum[21]), .A2(n3), .ZN(N24) );
  AND2_X1 U25 ( .A1(sum[20]), .A2(n3), .ZN(N23) );
  AND2_X1 U26 ( .A1(sum[19]), .A2(n3), .ZN(N22) );
  AND2_X1 U27 ( .A1(sum[18]), .A2(n3), .ZN(N21) );
  AND2_X1 U28 ( .A1(sum[17]), .A2(n3), .ZN(N20) );
  AND2_X1 U29 ( .A1(sum[16]), .A2(n3), .ZN(N19) );
  AND2_X1 U30 ( .A1(sum[15]), .A2(n3), .ZN(N18) );
  AND2_X1 U31 ( .A1(sum[14]), .A2(n3), .ZN(N17) );
  AND2_X1 U32 ( .A1(sum[13]), .A2(n3), .ZN(N16) );
  AND2_X1 U33 ( .A1(sum[12]), .A2(n3), .ZN(N15) );
  AND2_X1 U34 ( .A1(sum[11]), .A2(n3), .ZN(N14) );
  AND2_X1 U35 ( .A1(sum[10]), .A2(n3), .ZN(N13) );
  AND2_X1 U36 ( .A1(sum[9]), .A2(n3), .ZN(N12) );
  AND2_X1 U37 ( .A1(sum[8]), .A2(n3), .ZN(N11) );
  AND2_X1 U38 ( .A1(sum[7]), .A2(n3), .ZN(N10) );
  AND2_X1 U39 ( .A1(sum[6]), .A2(n3), .ZN(N9) );
  AND2_X1 U40 ( .A1(sum[5]), .A2(n3), .ZN(N8) );
  AND2_X1 U41 ( .A1(sum[4]), .A2(n3), .ZN(N7) );
  AND2_X1 U42 ( .A1(sum[3]), .A2(n3), .ZN(N6) );
  AND2_X1 U43 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U44 ( .A1(sum[1]), .A2(n3), .ZN(N4) );
  AND2_X1 U45 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
endmodule


module mac_1_DW_mult_tc_1 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n4, n6, n7, n9, n12, n13, n16, n19, n22, n25, n28, n31, n34, n37,
         n40, n42, n43, n46, n49, n52, n55, n58, n60, n61, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n97, n98, n99, n100, n101, n103, n105, n106, n107, n108, n109, n111,
         n113, n114, n115, n116, n117, n119, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n185,
         n186, n187, n188, n190, n193, n194, n195, n196, n198, n200, n201,
         n202, n203, n204, n205, n206, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n225,
         n227, n228, n230, n232, n233, n234, n236, n238, n239, n240, n241,
         n242, n244, n246, n247, n248, n249, n250, n252, n254, n255, n256,
         n257, n258, n259, n260, n261, n263, n264, n266, n268, n270, n271,
         n272, n273, n274, n275, n276, n278, n279, n280, n285, n286, n287,
         n291, n293, n295, n296, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n643, n644, n646, n649,
         n650, n652, n653, n655, n656, n658, n659, n661, n662, n664, n665,
         n667, n668, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1110, n1111, n1119, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1233, n1234, n1235, n1236, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n37 = a[13];
  assign n43 = a[15];
  assign n49 = a[17];
  assign n55 = a[19];
  assign n61 = b[0];
  assign n668 = a[0];
  assign n1090 = b[19];
  assign n1091 = b[18];
  assign n1092 = b[17];
  assign n1093 = b[16];
  assign n1094 = b[15];
  assign n1095 = b[14];
  assign n1096 = b[13];
  assign n1097 = b[12];
  assign n1098 = b[11];
  assign n1099 = b[10];
  assign n1100 = b[9];
  assign n1101 = b[8];
  assign n1102 = b[7];
  assign n1103 = b[6];
  assign n1104 = b[5];
  assign n1105 = b[4];
  assign n1106 = b[3];
  assign n1107 = b[2];
  assign n1108 = b[1];

  FA_X1 U333 ( .A(n681), .B(n304), .CI(n700), .CO(n300), .S(n301) );
  FA_X1 U334 ( .A(n305), .B(n682), .CI(n308), .CO(n302), .S(n303) );
  FA_X1 U336 ( .A(n312), .B(n683), .CI(n309), .CO(n306), .S(n307) );
  FA_X1 U337 ( .A(n701), .B(n314), .CI(n720), .CO(n308), .S(n309) );
  FA_X1 U338 ( .A(n313), .B(n320), .CI(n318), .CO(n310), .S(n311) );
  FA_X1 U339 ( .A(n684), .B(n702), .CI(n315), .CO(n312), .S(n313) );
  FA_X1 U341 ( .A(n324), .B(n321), .CI(n319), .CO(n316), .S(n317) );
  FA_X1 U342 ( .A(n328), .B(n721), .CI(n326), .CO(n318), .S(n319) );
  FA_X1 U343 ( .A(n703), .B(n685), .CI(n740), .CO(n320), .S(n321) );
  FA_X1 U344 ( .A(n325), .B(n327), .CI(n332), .CO(n322), .S(n323) );
  FA_X1 U345 ( .A(n336), .B(n329), .CI(n334), .CO(n324), .S(n325) );
  FA_X1 U346 ( .A(n686), .B(n704), .CI(n722), .CO(n326), .S(n327) );
  FA_X1 U348 ( .A(n340), .B(n342), .CI(n333), .CO(n330), .S(n331) );
  FA_X1 U349 ( .A(n335), .B(n344), .CI(n337), .CO(n332), .S(n333) );
  FA_X1 U350 ( .A(n705), .B(n346), .CI(n723), .CO(n334), .S(n335) );
  FA_X1 U351 ( .A(n741), .B(n687), .CI(n760), .CO(n336), .S(n337) );
  FA_X1 U352 ( .A(n350), .B(n343), .CI(n341), .CO(n338), .S(n339) );
  FA_X1 U353 ( .A(n345), .B(n354), .CI(n352), .CO(n340), .S(n341) );
  FA_X1 U354 ( .A(n347), .B(n724), .CI(n356), .CO(n342), .S(n343) );
  FA_X1 U355 ( .A(n742), .B(n706), .CI(n688), .CO(n344), .S(n345) );
  FA_X1 U357 ( .A(n360), .B(n353), .CI(n351), .CO(n348), .S(n349) );
  FA_X1 U358 ( .A(n357), .B(n355), .CI(n362), .CO(n350), .S(n351) );
  FA_X1 U359 ( .A(n366), .B(n743), .CI(n364), .CO(n352), .S(n353) );
  FA_X1 U360 ( .A(n707), .B(n761), .CI(n725), .CO(n354), .S(n355) );
  FA_X1 U361 ( .A(n368), .B(n689), .CI(n780), .CO(n356), .S(n357) );
  FA_X1 U362 ( .A(n372), .B(n363), .CI(n361), .CO(n358), .S(n359) );
  FA_X1 U363 ( .A(n376), .B(n365), .CI(n374), .CO(n360), .S(n361) );
  FA_X1 U364 ( .A(n378), .B(n380), .CI(n367), .CO(n362), .S(n363) );
  FA_X1 U365 ( .A(n690), .B(n708), .CI(n369), .CO(n364), .S(n365) );
  FA_X1 U366 ( .A(n762), .B(n726), .CI(n744), .CO(n366), .S(n367) );
  FA_X1 U368 ( .A(n384), .B(n375), .CI(n373), .CO(n370), .S(n371) );
  FA_X1 U369 ( .A(n377), .B(n388), .CI(n386), .CO(n372), .S(n373) );
  FA_X1 U370 ( .A(n379), .B(n390), .CI(n381), .CO(n374), .S(n375) );
  FA_X1 U371 ( .A(n727), .B(n745), .CI(n392), .CO(n376), .S(n377) );
  FA_X1 U372 ( .A(n709), .B(n781), .CI(n763), .CO(n378), .S(n379) );
  FA_X1 U373 ( .A(n394), .B(n691), .CI(n800), .CO(n380), .S(n381) );
  FA_X1 U374 ( .A(n398), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U375 ( .A(n389), .B(n402), .CI(n400), .CO(n384), .S(n385) );
  FA_X1 U376 ( .A(n391), .B(n404), .CI(n393), .CO(n386), .S(n387) );
  FA_X1 U378 ( .A(n746), .B(n782), .CI(n764), .CO(n390), .S(n391) );
  FA_X1 U379 ( .A(n692), .B(n728), .CI(n710), .CO(n392), .S(n393) );
  FA_X1 U382 ( .A(n403), .B(n416), .CI(n414), .CO(n398), .S(n399) );
  FA_X1 U383 ( .A(n409), .B(n407), .CI(n418), .CO(n400), .S(n401) );
  FA_X1 U384 ( .A(n420), .B(n422), .CI(n405), .CO(n402), .S(n403) );
  FA_X1 U385 ( .A(n729), .B(n765), .CI(n747), .CO(n404), .S(n405) );
  FA_X1 U386 ( .A(n711), .B(n801), .CI(n783), .CO(n406), .S(n407) );
  FA_X1 U387 ( .A(n424), .B(n693), .CI(n820), .CO(n408), .S(n409) );
  FA_X1 U388 ( .A(n428), .B(n415), .CI(n413), .CO(n410), .S(n411) );
  FA_X1 U391 ( .A(n436), .B(n438), .CI(n421), .CO(n416), .S(n417) );
  FA_X1 U393 ( .A(n766), .B(n712), .CI(n694), .CO(n420), .S(n421) );
  FA_X1 U394 ( .A(n802), .B(n730), .CI(n784), .CO(n422), .S(n423) );
  FA_X1 U397 ( .A(n433), .B(n448), .CI(n446), .CO(n428), .S(n429) );
  FA_X1 U398 ( .A(n450), .B(n441), .CI(n435), .CO(n430), .S(n431) );
  FA_X1 U399 ( .A(n437), .B(n452), .CI(n439), .CO(n432), .S(n433) );
  FA_X1 U400 ( .A(n454), .B(n767), .CI(n456), .CO(n434), .S(n435) );
  FA_X1 U401 ( .A(n731), .B(n785), .CI(n749), .CO(n436), .S(n437) );
  FA_X1 U402 ( .A(n458), .B(n803), .CI(n713), .CO(n438), .S(n439) );
  FA_X1 U404 ( .A(n462), .B(n447), .CI(n445), .CO(n442), .S(n443) );
  FA_X1 U405 ( .A(n449), .B(n466), .CI(n464), .CO(n444), .S(n445) );
  FA_X1 U406 ( .A(n468), .B(n453), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U407 ( .A(n455), .B(n470), .CI(n457), .CO(n448), .S(n449) );
  FA_X1 U408 ( .A(n474), .B(n476), .CI(n472), .CO(n450), .S(n451) );
  FA_X1 U409 ( .A(n768), .B(n786), .CI(n459), .CO(n452), .S(n453) );
  FA_X1 U410 ( .A(n732), .B(n804), .CI(n714), .CO(n454), .S(n455) );
  FA_X1 U411 ( .A(n696), .B(n750), .CI(n822), .CO(n456), .S(n457) );
  FA_X1 U416 ( .A(n473), .B(n488), .CI(n475), .CO(n466), .S(n467) );
  FA_X1 U417 ( .A(n477), .B(n490), .CI(n492), .CO(n468), .S(n469) );
  FA_X1 U418 ( .A(n805), .B(n823), .CI(n494), .CO(n470), .S(n471) );
  FA_X1 U419 ( .A(n841), .B(n751), .CI(n733), .CO(n472), .S(n473) );
  FA_X1 U423 ( .A(n498), .B(n483), .CI(n481), .CO(n478), .S(n479) );
  FA_X1 U424 ( .A(n500), .B(n487), .CI(n485), .CO(n480), .S(n481) );
  FA_X1 U425 ( .A(n504), .B(n493), .CI(n502), .CO(n482), .S(n483) );
  FA_X1 U426 ( .A(n491), .B(n506), .CI(n489), .CO(n484), .S(n485) );
  FA_X1 U428 ( .A(n770), .B(n824), .CI(n842), .CO(n488), .S(n489) );
  FA_X1 U429 ( .A(n861), .B(n806), .CI(n752), .CO(n490), .S(n491) );
  FA_X1 U430 ( .A(n788), .B(n670), .CI(n734), .CO(n492), .S(n493) );
  HA_X1 U431 ( .A(n716), .B(n698), .CO(n494), .S(n495) );
  FA_X1 U432 ( .A(n514), .B(n501), .CI(n499), .CO(n496), .S(n497) );
  FA_X1 U434 ( .A(n520), .B(n509), .CI(n518), .CO(n500), .S(n501) );
  FA_X1 U435 ( .A(n511), .B(n522), .CI(n507), .CO(n502), .S(n503) );
  FA_X1 U436 ( .A(n526), .B(n807), .CI(n524), .CO(n504), .S(n505) );
  FA_X1 U437 ( .A(n789), .B(n825), .CI(n771), .CO(n506), .S(n507) );
  FA_X1 U438 ( .A(n717), .B(n753), .CI(n843), .CO(n508), .S(n509) );
  FA_X1 U439 ( .A(n862), .B(n699), .CI(n735), .CO(n510), .S(n511) );
  FA_X1 U440 ( .A(n517), .B(n530), .CI(n515), .CO(n512), .S(n513) );
  FA_X1 U441 ( .A(n532), .B(n521), .CI(n519), .CO(n514), .S(n515) );
  FA_X1 U443 ( .A(n540), .B(n538), .CI(n536), .CO(n518), .S(n519) );
  FA_X1 U444 ( .A(n826), .B(n844), .CI(n527), .CO(n520), .S(n521) );
  FA_X1 U445 ( .A(n754), .B(n772), .CI(n808), .CO(n522), .S(n523) );
  FA_X1 U446 ( .A(n863), .B(n790), .CI(n671), .CO(n524), .S(n525) );
  HA_X1 U447 ( .A(n736), .B(n718), .CO(n526), .S(n527) );
  FA_X1 U451 ( .A(n552), .B(n554), .CI(n550), .CO(n534), .S(n535) );
  FA_X1 U453 ( .A(n773), .B(n737), .CI(n845), .CO(n538), .S(n539) );
  FA_X1 U457 ( .A(n562), .B(n564), .CI(n551), .CO(n546), .S(n547) );
  FA_X1 U458 ( .A(n555), .B(n846), .CI(n566), .CO(n548), .S(n549) );
  FA_X1 U459 ( .A(n865), .B(n792), .CI(n828), .CO(n550), .S(n551) );
  FA_X1 U460 ( .A(n774), .B(n672), .CI(n810), .CO(n552), .S(n553) );
  HA_X1 U461 ( .A(n738), .B(n756), .CO(n554), .S(n555) );
  FA_X1 U462 ( .A(n561), .B(n570), .CI(n559), .CO(n556), .S(n557) );
  FA_X1 U463 ( .A(n563), .B(n565), .CI(n572), .CO(n558), .S(n559) );
  FA_X1 U466 ( .A(n757), .B(n847), .CI(n793), .CO(n564), .S(n565) );
  FA_X1 U467 ( .A(n866), .B(n739), .CI(n775), .CO(n566), .S(n567) );
  FA_X1 U468 ( .A(n582), .B(n573), .CI(n571), .CO(n568), .S(n569) );
  FA_X1 U469 ( .A(n577), .B(n575), .CI(n584), .CO(n570), .S(n571) );
  FA_X1 U470 ( .A(n588), .B(n579), .CI(n586), .CO(n572), .S(n573) );
  FA_X1 U471 ( .A(n794), .B(n848), .CI(n830), .CO(n574), .S(n575) );
  FA_X1 U472 ( .A(n867), .B(n812), .CI(n673), .CO(n576), .S(n577) );
  HA_X1 U473 ( .A(n758), .B(n776), .CO(n578), .S(n579) );
  FA_X1 U474 ( .A(n585), .B(n592), .CI(n583), .CO(n580), .S(n581) );
  FA_X1 U475 ( .A(n587), .B(n589), .CI(n594), .CO(n582), .S(n583) );
  FA_X1 U476 ( .A(n598), .B(n831), .CI(n596), .CO(n584), .S(n585) );
  FA_X1 U477 ( .A(n777), .B(n849), .CI(n813), .CO(n586), .S(n587) );
  FA_X1 U478 ( .A(n868), .B(n759), .CI(n795), .CO(n588), .S(n589) );
  FA_X1 U479 ( .A(n602), .B(n595), .CI(n593), .CO(n590), .S(n591) );
  FA_X1 U480 ( .A(n604), .B(n606), .CI(n597), .CO(n592), .S(n593) );
  FA_X1 U481 ( .A(n814), .B(n850), .CI(n599), .CO(n594), .S(n595) );
  FA_X1 U482 ( .A(n869), .B(n832), .CI(n674), .CO(n596), .S(n597) );
  HA_X1 U483 ( .A(n796), .B(n778), .CO(n598), .S(n599) );
  FA_X1 U484 ( .A(n610), .B(n605), .CI(n603), .CO(n600), .S(n601) );
  FA_X1 U485 ( .A(n612), .B(n614), .CI(n607), .CO(n602), .S(n603) );
  FA_X1 U486 ( .A(n797), .B(n851), .CI(n833), .CO(n604), .S(n605) );
  FA_X1 U487 ( .A(n815), .B(n779), .CI(n870), .CO(n606), .S(n607) );
  FA_X1 U488 ( .A(n613), .B(n618), .CI(n611), .CO(n608), .S(n609) );
  FA_X1 U489 ( .A(n615), .B(n871), .CI(n620), .CO(n610), .S(n611) );
  FA_X1 U490 ( .A(n852), .B(n834), .CI(n675), .CO(n612), .S(n613) );
  HA_X1 U491 ( .A(n798), .B(n816), .CO(n614), .S(n615) );
  FA_X1 U492 ( .A(n621), .B(n624), .CI(n619), .CO(n616), .S(n617) );
  FA_X1 U493 ( .A(n817), .B(n853), .CI(n626), .CO(n618), .S(n619) );
  FA_X1 U494 ( .A(n835), .B(n799), .CI(n872), .CO(n620), .S(n621) );
  FA_X1 U495 ( .A(n630), .B(n627), .CI(n625), .CO(n622), .S(n623) );
  FA_X1 U496 ( .A(n854), .B(n873), .CI(n676), .CO(n624), .S(n625) );
  HA_X1 U497 ( .A(n818), .B(n836), .CO(n626), .S(n627) );
  FA_X1 U498 ( .A(n634), .B(n837), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U499 ( .A(n874), .B(n819), .CI(n855), .CO(n630), .S(n631) );
  FA_X1 U500 ( .A(n677), .B(n856), .CI(n635), .CO(n632), .S(n633) );
  HA_X1 U501 ( .A(n838), .B(n875), .CO(n634), .S(n635) );
  FA_X1 U502 ( .A(n876), .B(n839), .CI(n857), .CO(n636), .S(n637) );
  HA_X1 U503 ( .A(n858), .B(n877), .CO(n638), .S(n639) );
  BUF_X2 U1025 ( .A(n6), .Z(n1506) );
  AND2_X1 U1026 ( .A1(n40), .A2(n1483), .ZN(n1499) );
  BUF_X1 U1027 ( .A(n1564), .Z(n1253) );
  BUF_X1 U1028 ( .A(n1102), .Z(n1264) );
  XNOR2_X1 U1029 ( .A(n1565), .B(n1539), .ZN(n1233) );
  BUF_X2 U1030 ( .A(n1245), .Z(n1503) );
  AND2_X1 U1031 ( .A1(n513), .A2(n528), .ZN(n1408) );
  BUF_X1 U1032 ( .A(n1098), .Z(n1557) );
  BUF_X1 U1033 ( .A(n1099), .Z(n1371) );
  BUF_X1 U1034 ( .A(n1098), .Z(n1316) );
  BUF_X2 U1035 ( .A(n43), .Z(n1545) );
  BUF_X1 U1036 ( .A(n1099), .Z(n1373) );
  BUF_X2 U1037 ( .A(n7), .Z(n1539) );
  BUF_X2 U1038 ( .A(n1096), .Z(n1559) );
  BUF_X2 U1039 ( .A(n19), .Z(n1541) );
  BUF_X2 U1040 ( .A(n1515), .Z(n1309) );
  BUF_X2 U1041 ( .A(n1097), .Z(n1558) );
  NAND3_X1 U1042 ( .A1(n1287), .A2(n1288), .A3(n1289), .ZN(n486) );
  BUF_X2 U1043 ( .A(n1093), .Z(n1562) );
  BUF_X2 U1044 ( .A(n55), .Z(n1366) );
  INV_X1 U1045 ( .A(n1408), .ZN(n185) );
  AND2_X1 U1046 ( .A1(n1478), .A2(n9), .ZN(n1234) );
  BUF_X1 U1047 ( .A(n1104), .Z(n1552) );
  BUF_X1 U1048 ( .A(n1098), .Z(n1315) );
  OR2_X1 U1049 ( .A1(n557), .A2(n568), .ZN(n1235) );
  OR2_X1 U1050 ( .A1(n679), .A2(n879), .ZN(n1236) );
  AND2_X1 U1051 ( .A1(n1236), .A2(n263), .ZN(product[1]) );
  CLKBUF_X2 U1052 ( .A(n25), .Z(n1542) );
  CLKBUF_X2 U1053 ( .A(n25), .Z(n1362) );
  CLKBUF_X1 U1054 ( .A(n164), .Z(n1238) );
  BUF_X2 U1055 ( .A(n1514), .Z(n1467) );
  BUF_X2 U1056 ( .A(n1540), .Z(n1239) );
  CLKBUF_X2 U1057 ( .A(n1540), .Z(n1240) );
  CLKBUF_X3 U1058 ( .A(n1540), .Z(n1241) );
  BUF_X1 U1059 ( .A(n13), .Z(n1540) );
  NAND2_X1 U1060 ( .A1(n1245), .A2(n1377), .ZN(n1242) );
  NAND2_X1 U1061 ( .A1(n1245), .A2(n1377), .ZN(n12) );
  CLKBUF_X2 U1062 ( .A(n16), .Z(n1517) );
  BUF_X1 U1063 ( .A(n16), .Z(n1518) );
  INV_X1 U1064 ( .A(n220), .ZN(n1243) );
  INV_X1 U1065 ( .A(n1499), .ZN(n1244) );
  INV_X1 U1066 ( .A(n1499), .ZN(n42) );
  CLKBUF_X2 U1067 ( .A(n40), .Z(n1297) );
  BUF_X2 U1068 ( .A(n1514), .Z(n1466) );
  XNOR2_X1 U1069 ( .A(n1), .B(a[2]), .ZN(n1245) );
  CLKBUF_X1 U1070 ( .A(n668), .Z(n1246) );
  CLKBUF_X3 U1071 ( .A(n9), .Z(n1504) );
  XOR2_X1 U1072 ( .A(n537), .B(n539), .Z(n1247) );
  XOR2_X1 U1073 ( .A(n541), .B(n1247), .Z(n533) );
  NAND2_X1 U1074 ( .A1(n541), .A2(n537), .ZN(n1248) );
  NAND2_X1 U1075 ( .A1(n541), .A2(n539), .ZN(n1249) );
  NAND2_X1 U1076 ( .A1(n539), .A2(n537), .ZN(n1250) );
  NAND3_X1 U1077 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n532) );
  INV_X1 U1078 ( .A(n659), .ZN(n1251) );
  CLKBUF_X3 U1079 ( .A(n22), .Z(n1512) );
  CLKBUF_X3 U1080 ( .A(n7), .Z(n1321) );
  CLKBUF_X1 U1081 ( .A(n52), .Z(n1511) );
  CLKBUF_X2 U1082 ( .A(n19), .Z(n1332) );
  INV_X1 U1083 ( .A(n46), .ZN(n1252) );
  CLKBUF_X3 U1084 ( .A(n46), .Z(n1513) );
  CLKBUF_X1 U1085 ( .A(n1104), .Z(n1365) );
  BUF_X2 U1086 ( .A(n1091), .Z(n1564) );
  XNOR2_X1 U1087 ( .A(n1254), .B(n430), .ZN(n413) );
  XNOR2_X1 U1088 ( .A(n432), .B(n417), .ZN(n1254) );
  CLKBUF_X1 U1089 ( .A(n141), .Z(n1255) );
  XOR2_X1 U1090 ( .A(n419), .B(n423), .Z(n1256) );
  XOR2_X1 U1091 ( .A(n434), .B(n1256), .Z(n415) );
  NAND2_X1 U1092 ( .A1(n434), .A2(n419), .ZN(n1257) );
  NAND2_X1 U1093 ( .A1(n434), .A2(n423), .ZN(n1258) );
  NAND2_X1 U1094 ( .A1(n419), .A2(n423), .ZN(n1259) );
  NAND3_X1 U1095 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n414) );
  CLKBUF_X3 U1096 ( .A(n37), .Z(n1325) );
  BUF_X1 U1097 ( .A(n1496), .Z(n1456) );
  CLKBUF_X3 U1098 ( .A(n31), .Z(n1260) );
  CLKBUF_X1 U1099 ( .A(n31), .Z(n1543) );
  OR2_X1 U1100 ( .A1(n1497), .A2(n1498), .ZN(n1327) );
  CLKBUF_X1 U1101 ( .A(n482), .Z(n1261) );
  BUF_X2 U1102 ( .A(n1103), .Z(n1553) );
  CLKBUF_X1 U1103 ( .A(n1521), .Z(n1262) );
  OR2_X1 U1104 ( .A1(n513), .A2(n528), .ZN(n1521) );
  NAND2_X1 U1105 ( .A1(n1433), .A2(n301), .ZN(n1263) );
  BUF_X2 U1106 ( .A(n1108), .Z(n1548) );
  BUF_X1 U1107 ( .A(n1105), .Z(n1265) );
  BUF_X2 U1108 ( .A(n1107), .Z(n1549) );
  OR2_X2 U1109 ( .A1(n1497), .A2(n1252), .ZN(n1266) );
  CLKBUF_X1 U1110 ( .A(n1108), .Z(n1351) );
  XOR2_X1 U1111 ( .A(n811), .B(n829), .Z(n1267) );
  XOR2_X1 U1112 ( .A(n578), .B(n1267), .Z(n563) );
  NAND2_X1 U1113 ( .A1(n578), .A2(n811), .ZN(n1268) );
  NAND2_X1 U1114 ( .A1(n578), .A2(n829), .ZN(n1269) );
  NAND2_X1 U1115 ( .A1(n811), .A2(n829), .ZN(n1270) );
  NAND3_X1 U1116 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n562) );
  BUF_X2 U1117 ( .A(n1100), .Z(n1556) );
  XOR2_X1 U1118 ( .A(n560), .B(n553), .Z(n1271) );
  XOR2_X1 U1119 ( .A(n1271), .B(n549), .Z(n545) );
  XOR2_X1 U1120 ( .A(n547), .B(n558), .Z(n1272) );
  XOR2_X1 U1121 ( .A(n1272), .B(n545), .Z(n543) );
  NAND2_X1 U1122 ( .A1(n560), .A2(n553), .ZN(n1273) );
  NAND2_X1 U1123 ( .A1(n560), .A2(n549), .ZN(n1274) );
  NAND2_X1 U1124 ( .A1(n553), .A2(n549), .ZN(n1275) );
  NAND3_X1 U1125 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n544) );
  NAND2_X1 U1126 ( .A1(n547), .A2(n558), .ZN(n1276) );
  NAND2_X1 U1127 ( .A1(n547), .A2(n545), .ZN(n1277) );
  NAND2_X1 U1128 ( .A1(n558), .A2(n545), .ZN(n1278) );
  NAND3_X1 U1129 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n542) );
  XOR2_X1 U1130 ( .A(n567), .B(n576), .Z(n1279) );
  XOR2_X1 U1131 ( .A(n574), .B(n1279), .Z(n561) );
  NAND2_X1 U1132 ( .A1(n574), .A2(n567), .ZN(n1280) );
  NAND2_X1 U1133 ( .A1(n574), .A2(n576), .ZN(n1281) );
  NAND2_X1 U1134 ( .A1(n567), .A2(n576), .ZN(n1282) );
  NAND3_X1 U1135 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n560) );
  XNOR2_X1 U1136 ( .A(n769), .B(n1283), .ZN(n475) );
  XNOR2_X1 U1137 ( .A(n860), .B(n697), .ZN(n1283) );
  XNOR2_X1 U1138 ( .A(n1284), .B(n1261), .ZN(n463) );
  XNOR2_X1 U1139 ( .A(n467), .B(n484), .ZN(n1284) );
  CLKBUF_X1 U1140 ( .A(n172), .Z(n1285) );
  XOR2_X1 U1141 ( .A(n510), .B(n495), .Z(n1286) );
  XOR2_X1 U1142 ( .A(n1286), .B(n508), .Z(n487) );
  NAND2_X1 U1143 ( .A1(n510), .A2(n495), .ZN(n1287) );
  NAND2_X1 U1144 ( .A1(n510), .A2(n508), .ZN(n1288) );
  NAND2_X1 U1145 ( .A1(n495), .A2(n508), .ZN(n1289) );
  XOR2_X1 U1146 ( .A(n469), .B(n471), .Z(n1290) );
  XOR2_X1 U1147 ( .A(n1290), .B(n486), .Z(n465) );
  NAND2_X1 U1148 ( .A1(n471), .A2(n469), .ZN(n1291) );
  NAND2_X1 U1149 ( .A1(n471), .A2(n486), .ZN(n1292) );
  NAND2_X1 U1150 ( .A1(n469), .A2(n486), .ZN(n1293) );
  NAND3_X1 U1151 ( .A1(n1291), .A2(n1292), .A3(n1293), .ZN(n464) );
  CLKBUF_X1 U1152 ( .A(n1364), .Z(n1294) );
  BUF_X2 U1153 ( .A(n1364), .Z(n1295) );
  XNOR2_X1 U1154 ( .A(n1546), .B(a[18]), .ZN(n1364) );
  BUF_X2 U1155 ( .A(n49), .Z(n1546) );
  NOR2_X1 U1156 ( .A1(n557), .A2(n568), .ZN(n1296) );
  NOR2_X1 U1157 ( .A1(n557), .A2(n568), .ZN(n204) );
  CLKBUF_X1 U1158 ( .A(n40), .Z(n1508) );
  BUF_X2 U1159 ( .A(n1106), .Z(n1356) );
  BUF_X2 U1160 ( .A(n1365), .Z(n1304) );
  XNOR2_X1 U1161 ( .A(n1298), .B(n516), .ZN(n499) );
  XNOR2_X1 U1162 ( .A(n503), .B(n505), .ZN(n1298) );
  XNOR2_X1 U1163 ( .A(n1558), .B(n1332), .ZN(n1299) );
  NAND2_X1 U1164 ( .A1(n769), .A2(n860), .ZN(n1300) );
  NAND2_X1 U1165 ( .A1(n769), .A2(n697), .ZN(n1301) );
  NAND2_X1 U1166 ( .A1(n860), .A2(n697), .ZN(n1302) );
  NAND3_X1 U1167 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n474) );
  CLKBUF_X1 U1168 ( .A(n1457), .Z(n1303) );
  CLKBUF_X3 U1169 ( .A(n1496), .Z(n1457) );
  BUF_X1 U1170 ( .A(n1502), .Z(n1474) );
  BUF_X1 U1171 ( .A(n1365), .Z(n1305) );
  AND2_X2 U1172 ( .A1(n1482), .A2(n34), .ZN(n1501) );
  OR2_X1 U1173 ( .A1(n1497), .A2(n1498), .ZN(n1375) );
  CLKBUF_X1 U1174 ( .A(n1512), .Z(n1306) );
  INV_X1 U1175 ( .A(n394), .ZN(n395) );
  XNOR2_X1 U1176 ( .A(n1565), .B(n1538), .ZN(n1307) );
  CLKBUF_X1 U1177 ( .A(n1515), .Z(n1308) );
  BUF_X1 U1178 ( .A(n1502), .Z(n1310) );
  BUF_X1 U1179 ( .A(n1502), .Z(n1311) );
  BUF_X1 U1180 ( .A(n1100), .Z(n1318) );
  XNOR2_X1 U1181 ( .A(n1564), .B(n1342), .ZN(n1312) );
  CLKBUF_X1 U1182 ( .A(n150), .Z(n1313) );
  OAI22_X1 U1183 ( .A1(n1536), .A2(n1028), .B1(n1027), .B2(n1518), .ZN(n1314)
         );
  XNOR2_X1 U1184 ( .A(n1559), .B(n1541), .ZN(n1317) );
  XNOR2_X1 U1185 ( .A(n1319), .B(n827), .ZN(n537) );
  XNOR2_X1 U1186 ( .A(n809), .B(n791), .ZN(n1319) );
  BUF_X1 U1187 ( .A(n1472), .Z(n1320) );
  NAND2_X1 U1188 ( .A1(n1111), .A2(n1509), .ZN(n1472) );
  INV_X1 U1189 ( .A(n193), .ZN(n1322) );
  XNOR2_X1 U1190 ( .A(n1316), .B(n1362), .ZN(n1323) );
  CLKBUF_X1 U1191 ( .A(n1513), .Z(n1324) );
  CLKBUF_X1 U1192 ( .A(n37), .Z(n1544) );
  OR2_X2 U1193 ( .A1(n1497), .A2(n1252), .ZN(n1326) );
  XNOR2_X1 U1194 ( .A(n755), .B(n1328), .ZN(n541) );
  XNOR2_X1 U1195 ( .A(n864), .B(n719), .ZN(n1328) );
  INV_X1 U1196 ( .A(n1144), .ZN(n1329) );
  XNOR2_X1 U1197 ( .A(n399), .B(n1330), .ZN(n397) );
  XNOR2_X1 U1198 ( .A(n412), .B(n401), .ZN(n1330) );
  XNOR2_X1 U1199 ( .A(n1331), .B(n463), .ZN(n461) );
  XNOR2_X1 U1200 ( .A(n480), .B(n465), .ZN(n1331) );
  OAI22_X1 U1201 ( .A1(n1475), .A2(n997), .B1(n996), .B2(n1467), .ZN(n1333) );
  CLKBUF_X1 U1202 ( .A(n1102), .Z(n1554) );
  CLKBUF_X1 U1203 ( .A(n1102), .Z(n1363) );
  CLKBUF_X1 U1204 ( .A(n1560), .Z(n1334) );
  BUF_X2 U1205 ( .A(n1095), .Z(n1560) );
  CLKBUF_X1 U1206 ( .A(n1442), .Z(n1335) );
  CLKBUF_X1 U1207 ( .A(n1263), .Z(n1336) );
  NAND3_X1 U1208 ( .A1(n1336), .A2(n1335), .A3(n1443), .ZN(n1337) );
  CLKBUF_X1 U1209 ( .A(n443), .Z(n1338) );
  BUF_X2 U1210 ( .A(n61), .Z(n1339) );
  BUF_X1 U1211 ( .A(n61), .Z(n1340) );
  CLKBUF_X1 U1212 ( .A(n61), .Z(n1547) );
  CLKBUF_X2 U1213 ( .A(n1), .Z(n1341) );
  CLKBUF_X3 U1214 ( .A(n1), .Z(n1342) );
  CLKBUF_X1 U1215 ( .A(n1), .Z(n1538) );
  OR2_X1 U1216 ( .A1(n1338), .A2(n460), .ZN(n1343) );
  CLKBUF_X1 U1217 ( .A(n162), .Z(n1344) );
  CLKBUF_X1 U1218 ( .A(n1433), .Z(n1345) );
  NAND3_X1 U1219 ( .A1(n1431), .A2(n1430), .A3(n1432), .ZN(n1346) );
  CLKBUF_X1 U1220 ( .A(n1558), .Z(n1347) );
  BUF_X1 U1221 ( .A(n1107), .Z(n1348) );
  CLKBUF_X1 U1222 ( .A(n1559), .Z(n1349) );
  XNOR2_X1 U1223 ( .A(n1371), .B(n1542), .ZN(n1350) );
  INV_X2 U1224 ( .A(n1142), .ZN(n1352) );
  OR2_X2 U1225 ( .A1(n1497), .A2(n1498), .ZN(n1374) );
  OAI22_X1 U1226 ( .A1(n1507), .A2(n1073), .B1(n1072), .B2(n4), .ZN(n1353) );
  BUF_X1 U1227 ( .A(n1103), .Z(n1354) );
  XNOR2_X1 U1228 ( .A(n429), .B(n1355), .ZN(n427) );
  XNOR2_X1 U1229 ( .A(n444), .B(n431), .ZN(n1355) );
  CLKBUF_X3 U1230 ( .A(n52), .Z(n1510) );
  INV_X1 U1231 ( .A(n1343), .ZN(n1357) );
  CLKBUF_X1 U1232 ( .A(n1565), .Z(n1358) );
  BUF_X2 U1233 ( .A(n1090), .Z(n1565) );
  BUF_X2 U1234 ( .A(n1101), .Z(n1359) );
  CLKBUF_X1 U1235 ( .A(n1101), .Z(n1555) );
  CLKBUF_X1 U1236 ( .A(n1563), .Z(n1360) );
  BUF_X2 U1237 ( .A(n1092), .Z(n1563) );
  CLKBUF_X1 U1238 ( .A(n1562), .Z(n1361) );
  CLKBUF_X3 U1239 ( .A(n1094), .Z(n1561) );
  CLKBUF_X3 U1240 ( .A(n55), .Z(n1367) );
  BUF_X1 U1241 ( .A(n1105), .Z(n1368) );
  BUF_X1 U1242 ( .A(n1105), .Z(n1369) );
  INV_X1 U1243 ( .A(n1246), .ZN(n1370) );
  BUF_X1 U1244 ( .A(n1099), .Z(n1372) );
  CLKBUF_X1 U1245 ( .A(n1346), .Z(n1376) );
  XOR2_X1 U1246 ( .A(n7), .B(a[2]), .Z(n1377) );
  NOR2_X2 U1247 ( .A1(n581), .A2(n590), .ZN(n215) );
  NAND2_X1 U1248 ( .A1(n827), .A2(n1333), .ZN(n1378) );
  NAND2_X1 U1249 ( .A1(n827), .A2(n809), .ZN(n1379) );
  NAND2_X1 U1250 ( .A1(n1333), .A2(n809), .ZN(n1380) );
  NAND3_X1 U1251 ( .A1(n1378), .A2(n1379), .A3(n1380), .ZN(n536) );
  CLKBUF_X1 U1252 ( .A(n151), .Z(n1381) );
  OAI22_X1 U1253 ( .A1(n1405), .A2(n1049), .B1(n1233), .B2(n1503), .ZN(n1382)
         );
  OAI22_X1 U1254 ( .A1(n1405), .A2(n1049), .B1(n1048), .B2(n1503), .ZN(n458)
         );
  INV_X2 U1255 ( .A(n1500), .ZN(n1535) );
  XOR2_X1 U1256 ( .A(n406), .B(n395), .Z(n1383) );
  XOR2_X1 U1257 ( .A(n408), .B(n1383), .Z(n389) );
  NAND2_X1 U1258 ( .A1(n408), .A2(n406), .ZN(n1384) );
  NAND2_X1 U1259 ( .A1(n408), .A2(n395), .ZN(n1385) );
  NAND2_X1 U1260 ( .A1(n406), .A2(n395), .ZN(n1386) );
  NAND3_X1 U1261 ( .A1(n1384), .A2(n1385), .A3(n1386), .ZN(n388) );
  CLKBUF_X1 U1262 ( .A(n140), .Z(n1387) );
  NOR2_X1 U1263 ( .A1(n371), .A2(n382), .ZN(n1388) );
  NOR2_X1 U1264 ( .A1(n371), .A2(n382), .ZN(n135) );
  XOR2_X1 U1265 ( .A(n525), .B(n523), .Z(n1389) );
  XOR2_X1 U1266 ( .A(n1389), .B(n534), .Z(n517) );
  NAND2_X1 U1267 ( .A1(n525), .A2(n523), .ZN(n1390) );
  NAND2_X1 U1268 ( .A1(n525), .A2(n534), .ZN(n1391) );
  NAND2_X1 U1269 ( .A1(n523), .A2(n534), .ZN(n1392) );
  NAND3_X1 U1270 ( .A1(n1390), .A2(n1391), .A3(n1392), .ZN(n516) );
  NAND2_X1 U1271 ( .A1(n505), .A2(n503), .ZN(n1393) );
  NAND2_X1 U1272 ( .A1(n505), .A2(n516), .ZN(n1394) );
  NAND2_X1 U1273 ( .A1(n503), .A2(n516), .ZN(n1395) );
  NAND3_X1 U1274 ( .A1(n1393), .A2(n1394), .A3(n1395), .ZN(n498) );
  CLKBUF_X1 U1275 ( .A(n264), .Z(n1396) );
  CLKBUF_X1 U1276 ( .A(n176), .Z(n1397) );
  NAND3_X1 U1277 ( .A1(n1441), .A2(n1442), .A3(n1443), .ZN(n1398) );
  AOI21_X1 U1278 ( .B1(n175), .B2(n1322), .A(n1397), .ZN(n1399) );
  CLKBUF_X1 U1279 ( .A(n106), .Z(n1400) );
  NAND2_X1 U1280 ( .A1(n429), .A2(n444), .ZN(n1401) );
  NAND2_X1 U1281 ( .A1(n429), .A2(n431), .ZN(n1402) );
  NAND2_X1 U1282 ( .A1(n444), .A2(n431), .ZN(n1403) );
  NAND3_X1 U1283 ( .A1(n1401), .A2(n1402), .A3(n1403), .ZN(n426) );
  INV_X1 U1284 ( .A(n1234), .ZN(n1404) );
  INV_X1 U1285 ( .A(n1234), .ZN(n1405) );
  NAND3_X1 U1286 ( .A1(n1409), .A2(n1410), .A3(n1411), .ZN(n1406) );
  XNOR2_X1 U1287 ( .A(n1407), .B(n440), .ZN(n419) );
  XNOR2_X1 U1288 ( .A(n425), .B(n748), .ZN(n1407) );
  NAND2_X1 U1289 ( .A1(n430), .A2(n432), .ZN(n1409) );
  NAND2_X1 U1290 ( .A1(n430), .A2(n417), .ZN(n1410) );
  NAND2_X1 U1291 ( .A1(n432), .A2(n417), .ZN(n1411) );
  NAND3_X1 U1292 ( .A1(n1409), .A2(n1410), .A3(n1411), .ZN(n412) );
  NOR2_X1 U1293 ( .A1(n427), .A2(n442), .ZN(n1412) );
  NOR2_X1 U1294 ( .A1(n427), .A2(n442), .ZN(n158) );
  XOR2_X1 U1295 ( .A(n821), .B(n695), .Z(n1413) );
  XOR2_X1 U1296 ( .A(n1413), .B(n840), .Z(n441) );
  NAND2_X1 U1297 ( .A1(n821), .A2(n695), .ZN(n1414) );
  NAND2_X1 U1298 ( .A1(n821), .A2(n840), .ZN(n1415) );
  NAND2_X1 U1299 ( .A1(n695), .A2(n840), .ZN(n1416) );
  NAND3_X1 U1300 ( .A1(n1414), .A2(n1415), .A3(n1416), .ZN(n440) );
  NAND2_X1 U1301 ( .A1(n425), .A2(n748), .ZN(n1417) );
  NAND2_X1 U1302 ( .A1(n425), .A2(n440), .ZN(n1418) );
  NAND2_X1 U1303 ( .A1(n748), .A2(n440), .ZN(n1419) );
  NAND3_X1 U1304 ( .A1(n1417), .A2(n1418), .A3(n1419), .ZN(n418) );
  NAND2_X1 U1305 ( .A1(n467), .A2(n484), .ZN(n1420) );
  NAND2_X1 U1306 ( .A1(n467), .A2(n482), .ZN(n1421) );
  NAND2_X1 U1307 ( .A1(n484), .A2(n482), .ZN(n1422) );
  NAND3_X1 U1308 ( .A1(n1420), .A2(n1421), .A3(n1422), .ZN(n462) );
  NAND2_X1 U1309 ( .A1(n480), .A2(n465), .ZN(n1423) );
  NAND2_X1 U1310 ( .A1(n480), .A2(n463), .ZN(n1424) );
  NAND2_X1 U1311 ( .A1(n465), .A2(n463), .ZN(n1425) );
  NAND3_X1 U1312 ( .A1(n1423), .A2(n1424), .A3(n1425), .ZN(n460) );
  NAND2_X1 U1313 ( .A1(n399), .A2(n1406), .ZN(n1426) );
  NAND2_X1 U1314 ( .A1(n399), .A2(n401), .ZN(n1427) );
  NAND2_X1 U1315 ( .A1(n1406), .A2(n401), .ZN(n1428) );
  NAND3_X1 U1316 ( .A1(n1426), .A2(n1427), .A3(n1428), .ZN(n396) );
  XOR2_X1 U1317 ( .A(n310), .B(n307), .Z(n1429) );
  XOR2_X1 U1318 ( .A(n1396), .B(n1429), .Z(product[34]) );
  NAND2_X1 U1319 ( .A1(n264), .A2(n310), .ZN(n1430) );
  NAND2_X1 U1320 ( .A1(n264), .A2(n307), .ZN(n1431) );
  NAND2_X1 U1321 ( .A1(n310), .A2(n307), .ZN(n1432) );
  NAND3_X1 U1322 ( .A1(n1430), .A2(n1431), .A3(n1432), .ZN(n100) );
  NAND3_X1 U1323 ( .A1(n1436), .A2(n1435), .A3(n1437), .ZN(n1433) );
  INV_X1 U1324 ( .A(n1500), .ZN(n1537) );
  XOR2_X1 U1325 ( .A(n306), .B(n303), .Z(n1434) );
  XOR2_X1 U1326 ( .A(n1376), .B(n1434), .Z(product[35]) );
  NAND2_X1 U1327 ( .A1(n100), .A2(n306), .ZN(n1435) );
  NAND2_X1 U1328 ( .A1(n1346), .A2(n303), .ZN(n1436) );
  NAND2_X1 U1329 ( .A1(n306), .A2(n303), .ZN(n1437) );
  NAND3_X1 U1330 ( .A1(n1436), .A2(n1435), .A3(n1437), .ZN(n99) );
  CLKBUF_X1 U1331 ( .A(n127), .Z(n1438) );
  AND3_X1 U1332 ( .A1(n1453), .A2(n1452), .A3(n1451), .ZN(product[39]) );
  XOR2_X1 U1333 ( .A(n301), .B(n302), .Z(n1440) );
  XOR2_X1 U1334 ( .A(n1345), .B(n1440), .Z(product[36]) );
  NAND2_X1 U1335 ( .A1(n1433), .A2(n301), .ZN(n1441) );
  NAND2_X1 U1336 ( .A1(n99), .A2(n302), .ZN(n1442) );
  NAND2_X1 U1337 ( .A1(n301), .A2(n302), .ZN(n1443) );
  NAND3_X1 U1338 ( .A1(n1263), .A2(n1442), .A3(n1443), .ZN(n98) );
  NAND3_X1 U1339 ( .A1(n1448), .A2(n1449), .A3(n1447), .ZN(n1444) );
  CLKBUF_X1 U1340 ( .A(n114), .Z(n1445) );
  XOR2_X1 U1341 ( .A(n300), .B(n299), .Z(n1446) );
  XOR2_X1 U1342 ( .A(n1446), .B(n1337), .Z(product[37]) );
  NAND2_X1 U1343 ( .A1(n300), .A2(n299), .ZN(n1447) );
  NAND2_X1 U1344 ( .A1(n98), .A2(n300), .ZN(n1448) );
  NAND2_X1 U1345 ( .A1(n299), .A2(n1398), .ZN(n1449) );
  NAND3_X1 U1346 ( .A1(n1448), .A2(n1449), .A3(n1447), .ZN(n97) );
  XOR2_X1 U1347 ( .A(n680), .B(n298), .Z(n1450) );
  XOR2_X1 U1348 ( .A(n1444), .B(n1450), .Z(product[38]) );
  NAND2_X1 U1349 ( .A1(n680), .A2(n298), .ZN(n1451) );
  NAND2_X1 U1350 ( .A1(n97), .A2(n680), .ZN(n1452) );
  NAND2_X1 U1351 ( .A1(n97), .A2(n298), .ZN(n1453) );
  INV_X1 U1352 ( .A(n650), .ZN(n1454) );
  CLKBUF_X1 U1353 ( .A(n146), .Z(n1455) );
  NAND2_X1 U1354 ( .A1(n1479), .A2(n22), .ZN(n1496) );
  BUF_X4 U1355 ( .A(n49), .Z(n1458) );
  INV_X1 U1356 ( .A(n60), .ZN(n1459) );
  INV_X1 U1357 ( .A(n1459), .ZN(n1460) );
  AND2_X2 U1358 ( .A1(n1481), .A2(n16), .ZN(n1500) );
  AOI21_X1 U1359 ( .B1(n1262), .B2(n190), .A(n1408), .ZN(n1461) );
  AOI21_X1 U1360 ( .B1(n1455), .B2(n133), .A(n134), .ZN(n1462) );
  AOI21_X1 U1361 ( .B1(n114), .B2(n1492), .A(n111), .ZN(n1463) );
  CLKBUF_X1 U1362 ( .A(n153), .Z(n1464) );
  INV_X1 U1363 ( .A(n1499), .ZN(n1469) );
  CLKBUF_X1 U1364 ( .A(n122), .Z(n1465) );
  BUF_X1 U1365 ( .A(n28), .Z(n1514) );
  NAND2_X1 U1366 ( .A1(n1509), .A2(n1111), .ZN(n1471) );
  AOI21_X1 U1367 ( .B1(n122), .B2(n1491), .A(n119), .ZN(n1468) );
  NOR2_X1 U1368 ( .A1(n397), .A2(n410), .ZN(n1470) );
  AOI21_X1 U1369 ( .B1(n153), .B2(n126), .A(n127), .ZN(n1473) );
  BUF_X1 U1370 ( .A(n1502), .Z(n1475) );
  NAND2_X1 U1371 ( .A1(n1480), .A2(n28), .ZN(n1502) );
  NOR2_X1 U1372 ( .A1(n497), .A2(n512), .ZN(n1476) );
  INV_X1 U1373 ( .A(n1501), .ZN(n1477) );
  XOR2_X1 U1374 ( .A(n7), .B(a[2]), .Z(n1478) );
  XOR2_X1 U1375 ( .A(n19), .B(a[6]), .Z(n1479) );
  XOR2_X1 U1376 ( .A(n25), .B(a[8]), .Z(n1480) );
  XOR2_X1 U1377 ( .A(n13), .B(a[4]), .Z(n1481) );
  XOR2_X1 U1378 ( .A(n31), .B(a[10]), .Z(n1482) );
  XOR2_X1 U1379 ( .A(n37), .B(a[12]), .Z(n1483) );
  NOR2_X1 U1380 ( .A1(n461), .A2(n478), .ZN(n1484) );
  AOI21_X1 U1381 ( .B1(n173), .B2(n1238), .A(n165), .ZN(n163) );
  OAI21_X1 U1382 ( .B1(n152), .B2(n143), .A(n144), .ZN(n142) );
  INV_X1 U1383 ( .A(n145), .ZN(n143) );
  INV_X1 U1384 ( .A(n209), .ZN(n285) );
  INV_X1 U1385 ( .A(n171), .ZN(n279) );
  INV_X1 U1386 ( .A(n1387), .ZN(n273) );
  INV_X1 U1387 ( .A(n1520), .ZN(n211) );
  XOR2_X1 U1388 ( .A(n137), .B(n70), .Z(product[26]) );
  NAND2_X1 U1389 ( .A1(n272), .A2(n136), .ZN(n70) );
  AOI21_X1 U1390 ( .B1(n142), .B2(n273), .A(n139), .ZN(n137) );
  XOR2_X1 U1391 ( .A(n206), .B(n82), .Z(product[14]) );
  NAND2_X1 U1392 ( .A1(n1235), .A2(n205), .ZN(n82) );
  AOI21_X1 U1393 ( .B1(n211), .B2(n285), .A(n208), .ZN(n206) );
  XOR2_X1 U1394 ( .A(n168), .B(n76), .Z(product[20]) );
  NAND2_X1 U1395 ( .A1(n278), .A2(n167), .ZN(n76) );
  AOI21_X1 U1396 ( .B1(n173), .B2(n279), .A(n170), .ZN(n168) );
  XOR2_X1 U1397 ( .A(n163), .B(n75), .Z(product[21]) );
  NAND2_X1 U1398 ( .A1(n1343), .A2(n1344), .ZN(n75) );
  XOR2_X1 U1399 ( .A(n201), .B(n81), .Z(product[15]) );
  NAND2_X1 U1400 ( .A1(n1485), .A2(n200), .ZN(n81) );
  XOR2_X1 U1401 ( .A(n193), .B(n80), .Z(product[16]) );
  XOR2_X1 U1402 ( .A(n152), .B(n73), .Z(product[23]) );
  XNOR2_X1 U1403 ( .A(n173), .B(n77), .ZN(product[19]) );
  NAND2_X1 U1404 ( .A1(n279), .A2(n1285), .ZN(n77) );
  XNOR2_X1 U1405 ( .A(n149), .B(n72), .ZN(product[24]) );
  INV_X1 U1406 ( .A(n1470), .ZN(n274) );
  XNOR2_X1 U1407 ( .A(n130), .B(n69), .ZN(product[27]) );
  NAND2_X1 U1408 ( .A1(n271), .A2(n129), .ZN(n69) );
  INV_X1 U1409 ( .A(n128), .ZN(n271) );
  XNOR2_X1 U1410 ( .A(n142), .B(n71), .ZN(product[25]) );
  NAND2_X1 U1411 ( .A1(n273), .A2(n1255), .ZN(n71) );
  XNOR2_X1 U1412 ( .A(n211), .B(n83), .ZN(product[13]) );
  NAND2_X1 U1413 ( .A1(n285), .A2(n210), .ZN(n83) );
  XNOR2_X1 U1414 ( .A(n160), .B(n74), .ZN(product[22]) );
  NAND2_X1 U1415 ( .A1(n276), .A2(n159), .ZN(n74) );
  OAI21_X1 U1416 ( .B1(n163), .B2(n1357), .A(n1344), .ZN(n160) );
  INV_X1 U1417 ( .A(n210), .ZN(n208) );
  INV_X1 U1418 ( .A(n1285), .ZN(n170) );
  INV_X1 U1419 ( .A(n1255), .ZN(n139) );
  INV_X1 U1420 ( .A(n200), .ZN(n198) );
  AOI21_X1 U1421 ( .B1(n1488), .B2(n230), .A(n225), .ZN(n223) );
  INV_X1 U1422 ( .A(n227), .ZN(n225) );
  INV_X1 U1423 ( .A(n121), .ZN(n119) );
  INV_X1 U1424 ( .A(n113), .ZN(n111) );
  INV_X1 U1425 ( .A(n238), .ZN(n236) );
  NOR2_X1 U1426 ( .A1(n397), .A2(n410), .ZN(n147) );
  NAND2_X1 U1427 ( .A1(n443), .A2(n460), .ZN(n162) );
  NOR2_X1 U1428 ( .A1(n443), .A2(n460), .ZN(n161) );
  NOR2_X1 U1429 ( .A1(n461), .A2(n478), .ZN(n166) );
  OR2_X1 U1430 ( .A1(n529), .A2(n542), .ZN(n1528) );
  NAND2_X1 U1431 ( .A1(n268), .A2(n116), .ZN(n66) );
  INV_X1 U1432 ( .A(n115), .ZN(n268) );
  NAND2_X1 U1433 ( .A1(n266), .A2(n108), .ZN(n64) );
  INV_X1 U1434 ( .A(n107), .ZN(n266) );
  NAND2_X1 U1435 ( .A1(n291), .A2(n241), .ZN(n89) );
  INV_X1 U1436 ( .A(n240), .ZN(n291) );
  NAND2_X1 U1437 ( .A1(n270), .A2(n124), .ZN(n68) );
  INV_X1 U1438 ( .A(n123), .ZN(n270) );
  NOR2_X1 U1439 ( .A1(n359), .A2(n370), .ZN(n128) );
  NAND2_X1 U1440 ( .A1(n1492), .A2(n113), .ZN(n65) );
  NAND2_X1 U1441 ( .A1(n1490), .A2(n105), .ZN(n63) );
  NAND2_X1 U1442 ( .A1(n1491), .A2(n121), .ZN(n67) );
  NAND2_X1 U1443 ( .A1(n1489), .A2(n238), .ZN(n88) );
  XOR2_X1 U1444 ( .A(n228), .B(n86), .Z(product[10]) );
  AOI21_X1 U1445 ( .B1(n233), .B2(n1487), .A(n230), .ZN(n228) );
  AOI21_X1 U1446 ( .B1(n1521), .B2(n190), .A(n1408), .ZN(n181) );
  XOR2_X1 U1447 ( .A(n220), .B(n85), .Z(product[11]) );
  NAND2_X1 U1448 ( .A1(n287), .A2(n219), .ZN(n85) );
  INV_X1 U1449 ( .A(n218), .ZN(n287) );
  NOR2_X1 U1450 ( .A1(n383), .A2(n396), .ZN(n140) );
  NOR2_X1 U1451 ( .A1(n479), .A2(n496), .ZN(n171) );
  NOR2_X1 U1452 ( .A1(n569), .A2(n580), .ZN(n209) );
  NOR2_X1 U1453 ( .A1(n411), .A2(n426), .ZN(n150) );
  NAND2_X1 U1454 ( .A1(n383), .A2(n396), .ZN(n141) );
  NAND2_X1 U1455 ( .A1(n479), .A2(n496), .ZN(n172) );
  NAND2_X1 U1456 ( .A1(n569), .A2(n580), .ZN(n210) );
  INV_X1 U1457 ( .A(n232), .ZN(n230) );
  OR2_X1 U1458 ( .A1(n543), .A2(n556), .ZN(n1485) );
  XNOR2_X1 U1459 ( .A(n233), .B(n87), .ZN(product[9]) );
  NAND2_X1 U1460 ( .A1(n1487), .A2(n232), .ZN(n87) );
  XNOR2_X1 U1461 ( .A(n186), .B(n79), .ZN(product[17]) );
  INV_X1 U1462 ( .A(n1528), .ZN(n187) );
  XNOR2_X1 U1463 ( .A(n179), .B(n78), .ZN(product[18]) );
  NAND2_X1 U1464 ( .A1(n280), .A2(n178), .ZN(n78) );
  XNOR2_X1 U1465 ( .A(n217), .B(n84), .ZN(product[12]) );
  NAND2_X1 U1466 ( .A1(n286), .A2(n216), .ZN(n84) );
  OAI21_X1 U1467 ( .B1(n220), .B2(n218), .A(n219), .ZN(n217) );
  NAND2_X1 U1468 ( .A1(n359), .A2(n370), .ZN(n129) );
  NAND2_X1 U1469 ( .A1(n543), .A2(n556), .ZN(n200) );
  NAND2_X1 U1470 ( .A1(n557), .A2(n568), .ZN(n205) );
  NAND2_X1 U1471 ( .A1(n1521), .A2(n1528), .ZN(n180) );
  XNOR2_X1 U1472 ( .A(n1486), .B(n531), .ZN(n529) );
  XNOR2_X1 U1473 ( .A(n544), .B(n533), .ZN(n1486) );
  OAI21_X1 U1474 ( .B1(n256), .B2(n258), .A(n257), .ZN(n255) );
  AOI21_X1 U1475 ( .B1(n1495), .B2(n247), .A(n244), .ZN(n242) );
  INV_X1 U1476 ( .A(n246), .ZN(n244) );
  NOR2_X1 U1477 ( .A1(n591), .A2(n600), .ZN(n218) );
  NOR2_X1 U1478 ( .A1(n497), .A2(n512), .ZN(n177) );
  AOI21_X1 U1479 ( .B1(n1494), .B2(n255), .A(n252), .ZN(n250) );
  INV_X1 U1480 ( .A(n254), .ZN(n252) );
  OR2_X1 U1481 ( .A1(n609), .A2(n616), .ZN(n1487) );
  OR2_X1 U1482 ( .A1(n601), .A2(n608), .ZN(n1488) );
  NAND2_X1 U1483 ( .A1(n1495), .A2(n246), .ZN(n90) );
  NAND2_X1 U1484 ( .A1(n591), .A2(n600), .ZN(n219) );
  NOR2_X1 U1485 ( .A1(n317), .A2(n322), .ZN(n107) );
  NOR2_X1 U1486 ( .A1(n623), .A2(n628), .ZN(n240) );
  NOR2_X1 U1487 ( .A1(n349), .A2(n358), .ZN(n123) );
  NOR2_X1 U1488 ( .A1(n331), .A2(n338), .ZN(n115) );
  INV_X1 U1489 ( .A(n259), .ZN(n258) );
  OAI21_X1 U1490 ( .B1(n260), .B2(n263), .A(n261), .ZN(n259) );
  XNOR2_X1 U1491 ( .A(n92), .B(n255), .ZN(product[4]) );
  NAND2_X1 U1492 ( .A1(n1494), .A2(n254), .ZN(n92) );
  NAND2_X1 U1493 ( .A1(n609), .A2(n616), .ZN(n232) );
  NAND2_X1 U1494 ( .A1(n617), .A2(n622), .ZN(n238) );
  NAND2_X1 U1495 ( .A1(n311), .A2(n316), .ZN(n105) );
  NAND2_X1 U1496 ( .A1(n339), .A2(n348), .ZN(n121) );
  NAND2_X1 U1497 ( .A1(n323), .A2(n330), .ZN(n113) );
  NAND2_X1 U1498 ( .A1(n317), .A2(n322), .ZN(n108) );
  NAND2_X1 U1499 ( .A1(n623), .A2(n628), .ZN(n241) );
  NAND2_X1 U1500 ( .A1(n349), .A2(n358), .ZN(n124) );
  NAND2_X1 U1501 ( .A1(n331), .A2(n338), .ZN(n116) );
  NAND2_X1 U1502 ( .A1(n497), .A2(n512), .ZN(n178) );
  NAND2_X1 U1503 ( .A1(n581), .A2(n590), .ZN(n216) );
  OR2_X1 U1504 ( .A1(n617), .A2(n622), .ZN(n1489) );
  OR2_X1 U1505 ( .A1(n311), .A2(n316), .ZN(n1490) );
  OR2_X1 U1506 ( .A1(n339), .A2(n348), .ZN(n1491) );
  OR2_X1 U1507 ( .A1(n323), .A2(n330), .ZN(n1492) );
  NAND2_X1 U1508 ( .A1(n601), .A2(n608), .ZN(n227) );
  XOR2_X1 U1509 ( .A(n93), .B(n258), .Z(product[3]) );
  NAND2_X1 U1510 ( .A1(n295), .A2(n257), .ZN(n93) );
  INV_X1 U1511 ( .A(n256), .ZN(n295) );
  XOR2_X1 U1512 ( .A(n94), .B(n263), .Z(product[2]) );
  NAND2_X1 U1513 ( .A1(n296), .A2(n261), .ZN(n94) );
  INV_X1 U1514 ( .A(n260), .ZN(n296) );
  XOR2_X1 U1515 ( .A(n91), .B(n250), .Z(product[5]) );
  NAND2_X1 U1516 ( .A1(n293), .A2(n249), .ZN(n91) );
  INV_X1 U1517 ( .A(n248), .ZN(n293) );
  XNOR2_X1 U1518 ( .A(n1493), .B(n535), .ZN(n531) );
  XNOR2_X1 U1519 ( .A(n546), .B(n548), .ZN(n1493) );
  NAND2_X1 U1520 ( .A1(n639), .A2(n678), .ZN(n257) );
  NOR2_X1 U1521 ( .A1(n639), .A2(n678), .ZN(n256) );
  NOR2_X1 U1522 ( .A1(n878), .A2(n859), .ZN(n260) );
  NAND2_X1 U1523 ( .A1(n679), .A2(n879), .ZN(n263) );
  NAND2_X1 U1524 ( .A1(n878), .A2(n859), .ZN(n261) );
  OR2_X1 U1525 ( .A1(n637), .A2(n638), .ZN(n1494) );
  INV_X1 U1526 ( .A(n328), .ZN(n329) );
  NOR2_X1 U1527 ( .A1(n633), .A2(n636), .ZN(n248) );
  INV_X1 U1528 ( .A(n105), .ZN(n103) );
  INV_X1 U1529 ( .A(n298), .ZN(n299) );
  NAND2_X1 U1530 ( .A1(n629), .A2(n632), .ZN(n246) );
  OR2_X1 U1531 ( .A1(n629), .A2(n632), .ZN(n1495) );
  NAND2_X1 U1532 ( .A1(n633), .A2(n636), .ZN(n249) );
  NAND2_X1 U1533 ( .A1(n637), .A2(n638), .ZN(n254) );
  OR2_X1 U1534 ( .A1(n1340), .A2(n1148), .ZN(n1068) );
  OAI22_X1 U1535 ( .A1(n1507), .A2(n1086), .B1(n1085), .B2(n4), .ZN(n877) );
  OAI22_X1 U1536 ( .A1(n1507), .A2(n1088), .B1(n1087), .B2(n4), .ZN(n879) );
  OAI22_X1 U1537 ( .A1(n1507), .A2(n1149), .B1(n1089), .B2(n4), .ZN(n679) );
  OR2_X1 U1538 ( .A1(n1340), .A2(n1149), .ZN(n1089) );
  OAI22_X1 U1539 ( .A1(n1507), .A2(n1087), .B1(n1086), .B2(n4), .ZN(n878) );
  INV_X1 U1540 ( .A(n1382), .ZN(n459) );
  OAI22_X1 U1541 ( .A1(n1505), .A2(n1076), .B1(n1075), .B2(n4), .ZN(n867) );
  OAI22_X1 U1542 ( .A1(n1506), .A2(n1312), .B1(n1069), .B2(n4), .ZN(n861) );
  OAI22_X1 U1543 ( .A1(n1507), .A2(n1074), .B1(n1073), .B2(n4), .ZN(n865) );
  OAI22_X1 U1544 ( .A1(n1507), .A2(n1072), .B1(n1071), .B2(n4), .ZN(n863) );
  OAI22_X1 U1545 ( .A1(n1505), .A2(n1084), .B1(n1083), .B2(n4), .ZN(n875) );
  OR2_X1 U1546 ( .A1(n1340), .A2(n1147), .ZN(n1047) );
  AND2_X1 U1547 ( .A1(n1339), .A2(n662), .ZN(n839) );
  OAI22_X1 U1548 ( .A1(n1507), .A2(n1085), .B1(n1084), .B2(n4), .ZN(n876) );
  BUF_X1 U1549 ( .A(n34), .Z(n1516) );
  BUF_X1 U1550 ( .A(n34), .Z(n1515) );
  AND2_X1 U1551 ( .A1(n1339), .A2(n665), .ZN(n859) );
  BUF_X1 U1552 ( .A(n1105), .Z(n1551) );
  BUF_X1 U1553 ( .A(n1106), .Z(n1550) );
  INV_X1 U1554 ( .A(n655), .ZN(n780) );
  INV_X1 U1555 ( .A(n304), .ZN(n305) );
  AND2_X1 U1556 ( .A1(n1339), .A2(n641), .ZN(n699) );
  OAI22_X1 U1557 ( .A1(n1506), .A2(n1071), .B1(n1070), .B2(n4), .ZN(n862) );
  INV_X1 U1558 ( .A(n649), .ZN(n740) );
  INV_X1 U1559 ( .A(n643), .ZN(n700) );
  INV_X1 U1560 ( .A(n346), .ZN(n347) );
  OAI22_X1 U1561 ( .A1(n1506), .A2(n1077), .B1(n1076), .B2(n4), .ZN(n868) );
  AND2_X1 U1562 ( .A1(n1340), .A2(n650), .ZN(n759) );
  INV_X1 U1563 ( .A(n667), .ZN(n860) );
  INV_X1 U1564 ( .A(n652), .ZN(n760) );
  INV_X1 U1565 ( .A(n646), .ZN(n720) );
  OAI22_X1 U1566 ( .A1(n1507), .A2(n1080), .B1(n1079), .B2(n4), .ZN(n871) );
  AND2_X1 U1567 ( .A1(n1340), .A2(n653), .ZN(n779) );
  OAI22_X1 U1568 ( .A1(n1507), .A2(n1079), .B1(n1078), .B2(n4), .ZN(n870) );
  AND2_X1 U1569 ( .A1(n1339), .A2(n1252), .ZN(n739) );
  OAI22_X1 U1570 ( .A1(n1507), .A2(n1075), .B1(n1074), .B2(n4), .ZN(n866) );
  OAI22_X1 U1571 ( .A1(n1505), .A2(n1082), .B1(n1081), .B2(n4), .ZN(n873) );
  AND2_X1 U1572 ( .A1(n1339), .A2(n659), .ZN(n819) );
  OAI22_X1 U1573 ( .A1(n1505), .A2(n1083), .B1(n1082), .B2(n4), .ZN(n874) );
  OAI22_X1 U1574 ( .A1(n1505), .A2(n1081), .B1(n1080), .B2(n4), .ZN(n872) );
  AND2_X1 U1575 ( .A1(n1340), .A2(n656), .ZN(n799) );
  OAI22_X1 U1576 ( .A1(n1505), .A2(n1078), .B1(n1077), .B2(n4), .ZN(n869) );
  INV_X1 U1577 ( .A(n640), .ZN(n680) );
  INV_X1 U1578 ( .A(n368), .ZN(n369) );
  INV_X1 U1579 ( .A(n314), .ZN(n315) );
  OAI22_X1 U1580 ( .A1(n1307), .A2(n1506), .B1(n1307), .B2(n4), .ZN(n667) );
  INV_X1 U1581 ( .A(n661), .ZN(n820) );
  INV_X1 U1582 ( .A(n658), .ZN(n800) );
  OR2_X1 U1583 ( .A1(n1547), .A2(n1140), .ZN(n900) );
  OR2_X1 U1584 ( .A1(n1339), .A2(n1143), .ZN(n963) );
  OR2_X1 U1585 ( .A1(n1339), .A2(n1144), .ZN(n984) );
  OR2_X1 U1586 ( .A1(n1340), .A2(n1146), .ZN(n1026) );
  OR2_X1 U1587 ( .A1(n1340), .A2(n1142), .ZN(n942) );
  OR2_X1 U1588 ( .A1(n1339), .A2(n1141), .ZN(n921) );
  OR2_X1 U1589 ( .A1(n1340), .A2(n1145), .ZN(n1005) );
  INV_X2 U1590 ( .A(n668), .ZN(n4) );
  XNOR2_X1 U1591 ( .A(n43), .B(a[14]), .ZN(n1497) );
  INV_X1 U1592 ( .A(n46), .ZN(n1498) );
  AND2_X1 U1593 ( .A1(n1340), .A2(n1246), .ZN(product[0]) );
  XNOR2_X1 U1594 ( .A(n1), .B(a[2]), .ZN(n9) );
  CLKBUF_X1 U1595 ( .A(n6), .Z(n1505) );
  BUF_X2 U1596 ( .A(n6), .Z(n1507) );
  NAND2_X1 U1597 ( .A1(n1119), .A2(n1370), .ZN(n6) );
  XNOR2_X1 U1598 ( .A(n31), .B(a[12]), .ZN(n40) );
  CLKBUF_X1 U1599 ( .A(n52), .Z(n1509) );
  XNOR2_X1 U1600 ( .A(n43), .B(a[16]), .ZN(n52) );
  XNOR2_X1 U1601 ( .A(n13), .B(a[6]), .ZN(n22) );
  XNOR2_X1 U1602 ( .A(a[14]), .B(n37), .ZN(n46) );
  XNOR2_X1 U1603 ( .A(n19), .B(a[8]), .ZN(n28) );
  XNOR2_X1 U1604 ( .A(n25), .B(a[10]), .ZN(n34) );
  XNOR2_X1 U1605 ( .A(n7), .B(a[4]), .ZN(n16) );
  XNOR2_X1 U1606 ( .A(n1546), .B(a[18]), .ZN(n1519) );
  XNOR2_X1 U1607 ( .A(n1546), .B(a[18]), .ZN(n58) );
  AOI21_X1 U1608 ( .B1(n1243), .B2(n213), .A(n214), .ZN(n1520) );
  AOI21_X1 U1609 ( .B1(n221), .B2(n213), .A(n214), .ZN(n212) );
  INV_X1 U1610 ( .A(n215), .ZN(n286) );
  NOR2_X1 U1611 ( .A1(n215), .A2(n218), .ZN(n213) );
  OAI21_X1 U1612 ( .B1(n215), .B2(n219), .A(n216), .ZN(n214) );
  AOI21_X1 U1613 ( .B1(n211), .B2(n202), .A(n203), .ZN(n201) );
  NAND2_X1 U1614 ( .A1(n202), .A2(n1485), .ZN(n195) );
  NOR2_X1 U1615 ( .A1(n1296), .A2(n209), .ZN(n202) );
  INV_X1 U1616 ( .A(n1476), .ZN(n280) );
  NOR2_X1 U1617 ( .A1(n1476), .A2(n180), .ZN(n175) );
  NAND2_X1 U1618 ( .A1(n274), .A2(n148), .ZN(n72) );
  NAND2_X1 U1619 ( .A1(n397), .A2(n410), .ZN(n148) );
  INV_X1 U1620 ( .A(n1314), .ZN(n425) );
  NAND2_X1 U1621 ( .A1(n1528), .A2(n188), .ZN(n80) );
  INV_X1 U1622 ( .A(n188), .ZN(n190) );
  NAND2_X1 U1623 ( .A1(n529), .A2(n542), .ZN(n188) );
  XNOR2_X1 U1624 ( .A(n1358), .B(n1325), .ZN(n943) );
  XNOR2_X1 U1625 ( .A(n1253), .B(n1325), .ZN(n944) );
  XNOR2_X1 U1626 ( .A(n1361), .B(n1325), .ZN(n946) );
  XNOR2_X1 U1627 ( .A(n1360), .B(n1325), .ZN(n945) );
  XNOR2_X1 U1628 ( .A(n1561), .B(n1325), .ZN(n947) );
  XNOR2_X1 U1629 ( .A(n1334), .B(n1325), .ZN(n948) );
  XNOR2_X1 U1630 ( .A(n1559), .B(n1325), .ZN(n949) );
  XNOR2_X1 U1631 ( .A(n1316), .B(n1325), .ZN(n951) );
  XNOR2_X1 U1632 ( .A(n1558), .B(n1325), .ZN(n950) );
  XNOR2_X1 U1633 ( .A(n1373), .B(n1325), .ZN(n952) );
  XNOR2_X1 U1634 ( .A(n1553), .B(n1544), .ZN(n956) );
  XNOR2_X1 U1635 ( .A(n1264), .B(n1544), .ZN(n955) );
  XNOR2_X1 U1636 ( .A(n1552), .B(n1325), .ZN(n957) );
  XNOR2_X1 U1637 ( .A(n1368), .B(n1544), .ZN(n958) );
  XNOR2_X1 U1638 ( .A(n1555), .B(n1325), .ZN(n954) );
  XNOR2_X1 U1639 ( .A(n1556), .B(n1325), .ZN(n953) );
  INV_X1 U1640 ( .A(n1325), .ZN(n1143) );
  XNOR2_X1 U1641 ( .A(n1348), .B(n1544), .ZN(n960) );
  XNOR2_X1 U1642 ( .A(n1356), .B(n1544), .ZN(n959) );
  XNOR2_X1 U1643 ( .A(n1547), .B(n1544), .ZN(n962) );
  XNOR2_X1 U1644 ( .A(n1548), .B(n1544), .ZN(n961) );
  OAI21_X1 U1645 ( .B1(n204), .B2(n210), .A(n205), .ZN(n203) );
  OR2_X1 U1646 ( .A1(n787), .A2(n715), .ZN(n476) );
  XNOR2_X1 U1647 ( .A(n715), .B(n787), .ZN(n477) );
  NAND2_X1 U1648 ( .A1(n461), .A2(n478), .ZN(n167) );
  INV_X1 U1649 ( .A(n221), .ZN(n220) );
  NAND2_X1 U1650 ( .A1(n546), .A2(n548), .ZN(n1522) );
  NAND2_X1 U1651 ( .A1(n546), .A2(n535), .ZN(n1523) );
  NAND2_X1 U1652 ( .A1(n548), .A2(n535), .ZN(n1524) );
  NAND3_X1 U1653 ( .A1(n1522), .A2(n1523), .A3(n1524), .ZN(n530) );
  NAND2_X1 U1654 ( .A1(n544), .A2(n533), .ZN(n1525) );
  NAND2_X1 U1655 ( .A1(n544), .A2(n531), .ZN(n1526) );
  NAND2_X1 U1656 ( .A1(n533), .A2(n531), .ZN(n1527) );
  NAND3_X1 U1657 ( .A1(n1525), .A2(n1526), .A3(n1527), .ZN(n528) );
  XNOR2_X1 U1658 ( .A(n1358), .B(n1458), .ZN(n901) );
  XNOR2_X1 U1659 ( .A(n1253), .B(n1458), .ZN(n902) );
  XNOR2_X1 U1660 ( .A(n1361), .B(n1458), .ZN(n904) );
  XNOR2_X1 U1661 ( .A(n1360), .B(n1458), .ZN(n903) );
  XNOR2_X1 U1662 ( .A(n1561), .B(n1458), .ZN(n905) );
  XNOR2_X1 U1663 ( .A(n1334), .B(n1458), .ZN(n906) );
  XNOR2_X1 U1664 ( .A(n1349), .B(n1458), .ZN(n907) );
  XNOR2_X1 U1665 ( .A(n1347), .B(n1458), .ZN(n908) );
  XNOR2_X1 U1666 ( .A(n1316), .B(n1458), .ZN(n909) );
  XNOR2_X1 U1667 ( .A(n1373), .B(n1458), .ZN(n910) );
  XNOR2_X1 U1668 ( .A(n1556), .B(n1458), .ZN(n911) );
  XNOR2_X1 U1669 ( .A(n1354), .B(n1458), .ZN(n914) );
  XNOR2_X1 U1670 ( .A(n1363), .B(n1458), .ZN(n913) );
  XNOR2_X1 U1671 ( .A(n1359), .B(n1458), .ZN(n912) );
  XNOR2_X1 U1672 ( .A(n1549), .B(n1458), .ZN(n918) );
  XNOR2_X1 U1673 ( .A(n1552), .B(n1458), .ZN(n915) );
  INV_X1 U1674 ( .A(n1458), .ZN(n1141) );
  XNOR2_X1 U1675 ( .A(n1339), .B(n1458), .ZN(n920) );
  XNOR2_X1 U1676 ( .A(n1548), .B(n1458), .ZN(n919) );
  XNOR2_X1 U1677 ( .A(n1550), .B(n1458), .ZN(n917) );
  XNOR2_X1 U1678 ( .A(n1265), .B(n1458), .ZN(n916) );
  XOR2_X1 U1679 ( .A(n1546), .B(a[16]), .Z(n1111) );
  NAND2_X1 U1680 ( .A1(n1262), .A2(n185), .ZN(n79) );
  NAND2_X1 U1681 ( .A1(n275), .A2(n1381), .ZN(n73) );
  XNOR2_X1 U1682 ( .A(n1358), .B(n1366), .ZN(n880) );
  XNOR2_X1 U1683 ( .A(n1253), .B(n1367), .ZN(n881) );
  XNOR2_X1 U1684 ( .A(n1360), .B(n1366), .ZN(n882) );
  XNOR2_X1 U1685 ( .A(n1361), .B(n1367), .ZN(n883) );
  XNOR2_X1 U1686 ( .A(n1334), .B(n1367), .ZN(n885) );
  XNOR2_X1 U1687 ( .A(n1561), .B(n1366), .ZN(n884) );
  XNOR2_X1 U1688 ( .A(n1349), .B(n1366), .ZN(n886) );
  XNOR2_X1 U1689 ( .A(n1347), .B(n1367), .ZN(n887) );
  XNOR2_X1 U1690 ( .A(n1315), .B(n1366), .ZN(n888) );
  XNOR2_X1 U1691 ( .A(n1372), .B(n1367), .ZN(n889) );
  XNOR2_X1 U1692 ( .A(n1318), .B(n1366), .ZN(n890) );
  XNOR2_X1 U1693 ( .A(n1359), .B(n1367), .ZN(n891) );
  XNOR2_X1 U1694 ( .A(n1102), .B(n1366), .ZN(n892) );
  XNOR2_X1 U1695 ( .A(n1553), .B(n1367), .ZN(n893) );
  XNOR2_X1 U1696 ( .A(n1305), .B(n1367), .ZN(n894) );
  XNOR2_X1 U1697 ( .A(n1547), .B(n1366), .ZN(n899) );
  XNOR2_X1 U1698 ( .A(n1368), .B(n1366), .ZN(n895) );
  XNOR2_X1 U1699 ( .A(n1548), .B(n1366), .ZN(n898) );
  INV_X1 U1700 ( .A(n1367), .ZN(n1140) );
  XNOR2_X1 U1701 ( .A(n1549), .B(n1366), .ZN(n897) );
  XNOR2_X1 U1702 ( .A(n1550), .B(n1367), .ZN(n896) );
  XOR2_X1 U1703 ( .A(n55), .B(a[18]), .Z(n1110) );
  NAND2_X1 U1704 ( .A1(n755), .A2(n1353), .ZN(n1529) );
  NAND2_X1 U1705 ( .A1(n755), .A2(n719), .ZN(n1530) );
  NAND2_X1 U1706 ( .A1(n1353), .A2(n719), .ZN(n1531) );
  NAND3_X1 U1707 ( .A1(n1529), .A2(n1530), .A3(n1531), .ZN(n540) );
  AND2_X1 U1708 ( .A1(n1339), .A2(n644), .ZN(n719) );
  OAI22_X1 U1709 ( .A1(n1507), .A2(n1073), .B1(n1072), .B2(n4), .ZN(n864) );
  XNOR2_X1 U1710 ( .A(n1555), .B(n1362), .ZN(n996) );
  XNOR2_X1 U1711 ( .A(n1369), .B(n1542), .ZN(n1000) );
  XNOR2_X1 U1712 ( .A(n1348), .B(n1542), .ZN(n1002) );
  XNOR2_X1 U1713 ( .A(n1558), .B(n1362), .ZN(n992) );
  XNOR2_X1 U1714 ( .A(n1371), .B(n1542), .ZN(n994) );
  XNOR2_X1 U1715 ( .A(n1318), .B(n1542), .ZN(n995) );
  INV_X1 U1716 ( .A(n1362), .ZN(n1145) );
  XNOR2_X1 U1717 ( .A(n1560), .B(n1362), .ZN(n990) );
  XNOR2_X1 U1718 ( .A(n1562), .B(n1362), .ZN(n988) );
  XNOR2_X1 U1719 ( .A(n1563), .B(n1362), .ZN(n987) );
  XNOR2_X1 U1720 ( .A(n1358), .B(n1362), .ZN(n985) );
  XNOR2_X1 U1721 ( .A(n1253), .B(n1542), .ZN(n986) );
  XNOR2_X1 U1722 ( .A(n1561), .B(n1542), .ZN(n989) );
  XNOR2_X1 U1723 ( .A(n1559), .B(n1542), .ZN(n991) );
  XNOR2_X1 U1724 ( .A(n1340), .B(n1362), .ZN(n1004) );
  XNOR2_X1 U1725 ( .A(n1351), .B(n1542), .ZN(n1003) );
  XNOR2_X1 U1726 ( .A(n1557), .B(n1362), .ZN(n993) );
  XNOR2_X1 U1727 ( .A(n1304), .B(n1362), .ZN(n999) );
  XNOR2_X1 U1728 ( .A(n1553), .B(n1542), .ZN(n998) );
  XNOR2_X1 U1729 ( .A(n1550), .B(n1362), .ZN(n1001) );
  XNOR2_X1 U1730 ( .A(n1264), .B(n1542), .ZN(n997) );
  XNOR2_X1 U1731 ( .A(n1253), .B(n1352), .ZN(n923) );
  XNOR2_X1 U1732 ( .A(n1358), .B(n1352), .ZN(n922) );
  XNOR2_X1 U1733 ( .A(n1360), .B(n1352), .ZN(n924) );
  XNOR2_X1 U1734 ( .A(n1561), .B(n1352), .ZN(n926) );
  XNOR2_X1 U1735 ( .A(n1361), .B(n1352), .ZN(n925) );
  XNOR2_X1 U1736 ( .A(n1334), .B(n1352), .ZN(n927) );
  XNOR2_X1 U1737 ( .A(n1349), .B(n1352), .ZN(n928) );
  XNOR2_X1 U1738 ( .A(n1347), .B(n1352), .ZN(n929) );
  XNOR2_X1 U1739 ( .A(n1315), .B(n1545), .ZN(n930) );
  XNOR2_X1 U1740 ( .A(n1318), .B(n1545), .ZN(n932) );
  XNOR2_X1 U1741 ( .A(n1372), .B(n1545), .ZN(n931) );
  XNOR2_X1 U1742 ( .A(n1359), .B(n1545), .ZN(n933) );
  XNOR2_X1 U1743 ( .A(n1553), .B(n1545), .ZN(n935) );
  XNOR2_X1 U1744 ( .A(n1554), .B(n1545), .ZN(n934) );
  XNOR2_X1 U1745 ( .A(n1547), .B(n1545), .ZN(n941) );
  XNOR2_X1 U1746 ( .A(n1552), .B(n1545), .ZN(n936) );
  INV_X1 U1747 ( .A(n1545), .ZN(n1142) );
  XNOR2_X1 U1748 ( .A(n1551), .B(n43), .ZN(n937) );
  XNOR2_X1 U1749 ( .A(n1550), .B(n1545), .ZN(n938) );
  XNOR2_X1 U1750 ( .A(n1548), .B(n1545), .ZN(n940) );
  XNOR2_X1 U1751 ( .A(n1549), .B(n1545), .ZN(n939) );
  INV_X1 U1752 ( .A(n1501), .ZN(n1532) );
  INV_X1 U1753 ( .A(n1501), .ZN(n1533) );
  INV_X1 U1754 ( .A(n1501), .ZN(n1534) );
  INV_X1 U1755 ( .A(n1500), .ZN(n1536) );
  NAND2_X1 U1756 ( .A1(n156), .A2(n164), .ZN(n154) );
  XNOR2_X1 U1757 ( .A(n1565), .B(n1332), .ZN(n1006) );
  INV_X1 U1758 ( .A(n1541), .ZN(n1146) );
  XNOR2_X1 U1759 ( .A(n1562), .B(n1332), .ZN(n1009) );
  XNOR2_X1 U1760 ( .A(n1563), .B(n1541), .ZN(n1008) );
  XNOR2_X1 U1761 ( .A(n1564), .B(n1332), .ZN(n1007) );
  XNOR2_X1 U1762 ( .A(n1340), .B(n1541), .ZN(n1025) );
  XNOR2_X1 U1763 ( .A(n1351), .B(n1332), .ZN(n1024) );
  XNOR2_X1 U1764 ( .A(n1316), .B(n1541), .ZN(n1014) );
  XNOR2_X1 U1765 ( .A(n1560), .B(n1541), .ZN(n1011) );
  XNOR2_X1 U1766 ( .A(n1561), .B(n1332), .ZN(n1010) );
  XNOR2_X1 U1767 ( .A(n1348), .B(n1332), .ZN(n1023) );
  XNOR2_X1 U1768 ( .A(n1558), .B(n1332), .ZN(n1013) );
  XNOR2_X1 U1769 ( .A(n1559), .B(n1541), .ZN(n1012) );
  XNOR2_X1 U1770 ( .A(n1305), .B(n1541), .ZN(n1020) );
  XNOR2_X1 U1771 ( .A(n1363), .B(n1332), .ZN(n1018) );
  XNOR2_X1 U1772 ( .A(n1354), .B(n1541), .ZN(n1019) );
  XNOR2_X1 U1773 ( .A(n1356), .B(n1332), .ZN(n1022) );
  XNOR2_X1 U1774 ( .A(n1359), .B(n1541), .ZN(n1017) );
  XNOR2_X1 U1775 ( .A(n1369), .B(n1541), .ZN(n1021) );
  XNOR2_X1 U1776 ( .A(n1556), .B(n1332), .ZN(n1016) );
  XNOR2_X1 U1777 ( .A(n1371), .B(n1541), .ZN(n1015) );
  XNOR2_X1 U1778 ( .A(n1359), .B(n1341), .ZN(n1080) );
  XNOR2_X1 U1779 ( .A(n1554), .B(n1342), .ZN(n1081) );
  XNOR2_X1 U1780 ( .A(n1563), .B(n1538), .ZN(n1071) );
  XNOR2_X1 U1781 ( .A(n1564), .B(n1342), .ZN(n1070) );
  XNOR2_X1 U1782 ( .A(n1354), .B(n1341), .ZN(n1082) );
  XNOR2_X1 U1783 ( .A(n1550), .B(n1341), .ZN(n1085) );
  XNOR2_X1 U1784 ( .A(n1559), .B(n1342), .ZN(n1075) );
  XNOR2_X1 U1785 ( .A(n1304), .B(n1342), .ZN(n1083) );
  XNOR2_X1 U1786 ( .A(n1318), .B(n1342), .ZN(n1079) );
  XNOR2_X1 U1787 ( .A(n1348), .B(n1341), .ZN(n1086) );
  XNOR2_X1 U1788 ( .A(n1368), .B(n1342), .ZN(n1084) );
  XNOR2_X1 U1789 ( .A(n1558), .B(n1341), .ZN(n1076) );
  XNOR2_X1 U1790 ( .A(n1372), .B(n1341), .ZN(n1078) );
  XNOR2_X1 U1791 ( .A(n1557), .B(n1342), .ZN(n1077) );
  XNOR2_X1 U1792 ( .A(n1340), .B(n1342), .ZN(n1088) );
  XNOR2_X1 U1793 ( .A(n1560), .B(n1341), .ZN(n1074) );
  XNOR2_X1 U1794 ( .A(n1351), .B(n1341), .ZN(n1087) );
  XNOR2_X1 U1795 ( .A(n1561), .B(n1538), .ZN(n1073) );
  XNOR2_X1 U1796 ( .A(n1562), .B(n1538), .ZN(n1072) );
  INV_X1 U1797 ( .A(n1342), .ZN(n1149) );
  XNOR2_X1 U1798 ( .A(n1565), .B(n1538), .ZN(n1069) );
  XOR2_X1 U1799 ( .A(n1), .B(n668), .Z(n1119) );
  INV_X1 U1800 ( .A(n1240), .ZN(n1147) );
  XNOR2_X1 U1801 ( .A(n1561), .B(n1240), .ZN(n1031) );
  XNOR2_X1 U1802 ( .A(n1348), .B(n1241), .ZN(n1044) );
  XNOR2_X1 U1803 ( .A(n1340), .B(n1241), .ZN(n1046) );
  XNOR2_X1 U1804 ( .A(n1351), .B(n1241), .ZN(n1045) );
  XNOR2_X1 U1805 ( .A(n1562), .B(n1240), .ZN(n1030) );
  XNOR2_X1 U1806 ( .A(n1563), .B(n1241), .ZN(n1029) );
  XNOR2_X1 U1807 ( .A(n1359), .B(n1240), .ZN(n1038) );
  XNOR2_X1 U1808 ( .A(n1564), .B(n1239), .ZN(n1028) );
  XNOR2_X1 U1809 ( .A(n1559), .B(n1239), .ZN(n1033) );
  XNOR2_X1 U1810 ( .A(n1305), .B(n1240), .ZN(n1041) );
  XNOR2_X1 U1811 ( .A(n1356), .B(n1240), .ZN(n1043) );
  XNOR2_X1 U1812 ( .A(n1265), .B(n1241), .ZN(n1042) );
  XNOR2_X1 U1813 ( .A(n1556), .B(n1241), .ZN(n1037) );
  XNOR2_X1 U1814 ( .A(n1354), .B(n1241), .ZN(n1040) );
  XNOR2_X1 U1815 ( .A(n1554), .B(n1240), .ZN(n1039) );
  XNOR2_X1 U1816 ( .A(n1239), .B(n1560), .ZN(n1032) );
  XNOR2_X1 U1817 ( .A(n1565), .B(n1239), .ZN(n1027) );
  XNOR2_X1 U1818 ( .A(n1372), .B(n1239), .ZN(n1036) );
  XNOR2_X1 U1819 ( .A(n1316), .B(n1239), .ZN(n1035) );
  XNOR2_X1 U1820 ( .A(n1558), .B(n1239), .ZN(n1034) );
  XNOR2_X1 U1821 ( .A(n1304), .B(n1321), .ZN(n1062) );
  INV_X1 U1822 ( .A(n1321), .ZN(n1148) );
  XNOR2_X1 U1823 ( .A(n1359), .B(n1321), .ZN(n1059) );
  XNOR2_X1 U1824 ( .A(n1563), .B(n1321), .ZN(n1050) );
  XNOR2_X1 U1825 ( .A(n1564), .B(n1539), .ZN(n1049) );
  XNOR2_X1 U1826 ( .A(n1340), .B(n1321), .ZN(n1067) );
  XNOR2_X1 U1827 ( .A(n1561), .B(n1539), .ZN(n1052) );
  XNOR2_X1 U1828 ( .A(n1562), .B(n1321), .ZN(n1051) );
  XNOR2_X1 U1829 ( .A(n1356), .B(n1321), .ZN(n1064) );
  XNOR2_X1 U1830 ( .A(n1354), .B(n1321), .ZN(n1061) );
  XNOR2_X1 U1831 ( .A(n1264), .B(n1321), .ZN(n1060) );
  XNOR2_X1 U1832 ( .A(n1369), .B(n1321), .ZN(n1063) );
  XNOR2_X1 U1833 ( .A(n1351), .B(n1321), .ZN(n1066) );
  XNOR2_X1 U1834 ( .A(n1315), .B(n1539), .ZN(n1056) );
  XNOR2_X1 U1835 ( .A(n1558), .B(n1321), .ZN(n1055) );
  XNOR2_X1 U1836 ( .A(n1565), .B(n1539), .ZN(n1048) );
  XNOR2_X1 U1837 ( .A(n1348), .B(n1321), .ZN(n1065) );
  XNOR2_X1 U1838 ( .A(n1318), .B(n1539), .ZN(n1058) );
  XNOR2_X1 U1839 ( .A(n1373), .B(n1539), .ZN(n1057) );
  XNOR2_X1 U1840 ( .A(n1559), .B(n1539), .ZN(n1054) );
  XNOR2_X1 U1841 ( .A(n1560), .B(n1539), .ZN(n1053) );
  XNOR2_X1 U1842 ( .A(n1358), .B(n1329), .ZN(n964) );
  XNOR2_X1 U1843 ( .A(n1253), .B(n1329), .ZN(n965) );
  XNOR2_X1 U1844 ( .A(n1360), .B(n1329), .ZN(n966) );
  XNOR2_X1 U1845 ( .A(n1562), .B(n1329), .ZN(n967) );
  XNOR2_X1 U1846 ( .A(n1315), .B(n1260), .ZN(n972) );
  XNOR2_X1 U1847 ( .A(n1561), .B(n1260), .ZN(n968) );
  XNOR2_X1 U1848 ( .A(n1558), .B(n1543), .ZN(n971) );
  XNOR2_X1 U1849 ( .A(n1560), .B(n1260), .ZN(n969) );
  XNOR2_X1 U1850 ( .A(n1559), .B(n1543), .ZN(n970) );
  XNOR2_X1 U1851 ( .A(n1373), .B(n1260), .ZN(n973) );
  XNOR2_X1 U1852 ( .A(n1556), .B(n1260), .ZN(n974) );
  INV_X1 U1853 ( .A(n1260), .ZN(n1144) );
  XNOR2_X1 U1854 ( .A(n1363), .B(n1260), .ZN(n976) );
  XNOR2_X1 U1855 ( .A(n1359), .B(n1260), .ZN(n975) );
  XNOR2_X1 U1856 ( .A(n1339), .B(n1260), .ZN(n983) );
  XNOR2_X1 U1857 ( .A(n1351), .B(n1260), .ZN(n982) );
  XNOR2_X1 U1858 ( .A(n1552), .B(n1543), .ZN(n978) );
  XNOR2_X1 U1859 ( .A(n1103), .B(n1543), .ZN(n977) );
  XNOR2_X1 U1860 ( .A(n1551), .B(n1260), .ZN(n979) );
  XNOR2_X1 U1861 ( .A(n1356), .B(n1260), .ZN(n980) );
  XNOR2_X1 U1862 ( .A(n1549), .B(n1543), .ZN(n981) );
  INV_X1 U1863 ( .A(n234), .ZN(n233) );
  OAI21_X1 U1864 ( .B1(n222), .B2(n234), .A(n223), .ZN(n221) );
  AOI21_X1 U1865 ( .B1(n239), .B2(n1489), .A(n236), .ZN(n234) );
  XNOR2_X1 U1866 ( .A(n239), .B(n88), .ZN(product[8]) );
  OAI21_X1 U1867 ( .B1(n193), .B2(n187), .A(n188), .ZN(n186) );
  INV_X1 U1868 ( .A(n1517), .ZN(n662) );
  INV_X1 U1869 ( .A(n664), .ZN(n840) );
  NOR2_X1 U1870 ( .A1(n131), .A2(n128), .ZN(n126) );
  NAND2_X1 U1871 ( .A1(n1488), .A2(n1487), .ZN(n222) );
  NAND2_X1 U1872 ( .A1(n1488), .A2(n227), .ZN(n86) );
  XOR2_X1 U1873 ( .A(n242), .B(n89), .Z(product[7]) );
  INV_X1 U1874 ( .A(n194), .ZN(n193) );
  OAI21_X1 U1875 ( .B1(n242), .B2(n240), .A(n241), .ZN(n239) );
  NAND2_X1 U1876 ( .A1(n145), .A2(n133), .ZN(n131) );
  INV_X1 U1877 ( .A(n1388), .ZN(n272) );
  OAI21_X1 U1878 ( .B1(n141), .B2(n135), .A(n136), .ZN(n134) );
  NOR2_X1 U1879 ( .A1(n140), .A2(n1388), .ZN(n133) );
  NAND2_X1 U1880 ( .A1(n371), .A2(n382), .ZN(n136) );
  INV_X1 U1881 ( .A(n1412), .ZN(n276) );
  NOR2_X1 U1882 ( .A1(n161), .A2(n1412), .ZN(n156) );
  OAI21_X1 U1883 ( .B1(n158), .B2(n162), .A(n159), .ZN(n157) );
  NAND2_X1 U1884 ( .A1(n427), .A2(n442), .ZN(n159) );
  INV_X1 U1885 ( .A(n1455), .ZN(n144) );
  AOI21_X1 U1886 ( .B1(n133), .B2(n146), .A(n134), .ZN(n132) );
  OAI21_X1 U1887 ( .B1(n151), .B2(n147), .A(n148), .ZN(n146) );
  NAND2_X1 U1888 ( .A1(n411), .A2(n426), .ZN(n151) );
  AOI21_X1 U1889 ( .B1(n203), .B2(n1485), .A(n198), .ZN(n196) );
  OAI21_X1 U1890 ( .B1(n195), .B2(n212), .A(n196), .ZN(n194) );
  INV_X1 U1891 ( .A(n1484), .ZN(n278) );
  OAI22_X1 U1892 ( .A1(n922), .A2(n1266), .B1(n922), .B2(n1324), .ZN(n646) );
  NOR2_X1 U1893 ( .A1(n1484), .A2(n171), .ZN(n164) );
  OAI21_X1 U1894 ( .B1(n166), .B2(n172), .A(n167), .ZN(n165) );
  OAI22_X1 U1895 ( .A1(n1326), .A2(n924), .B1(n923), .B2(n1324), .ZN(n721) );
  OAI22_X1 U1896 ( .A1(n1327), .A2(n923), .B1(n922), .B2(n1324), .ZN(n314) );
  OAI22_X1 U1897 ( .A1(n1374), .A2(n925), .B1(n924), .B2(n1324), .ZN(n722) );
  OAI22_X1 U1898 ( .A1(n1326), .A2(n927), .B1(n926), .B2(n1324), .ZN(n724) );
  OAI22_X1 U1899 ( .A1(n1327), .A2(n926), .B1(n925), .B2(n1324), .ZN(n723) );
  OAI22_X1 U1900 ( .A1(n1374), .A2(n928), .B1(n927), .B2(n1324), .ZN(n725) );
  OAI22_X1 U1901 ( .A1(n1266), .A2(n929), .B1(n928), .B2(n1513), .ZN(n726) );
  OAI22_X1 U1902 ( .A1(n1326), .A2(n930), .B1(n929), .B2(n1513), .ZN(n727) );
  OAI22_X1 U1903 ( .A1(n1327), .A2(n933), .B1(n932), .B2(n1513), .ZN(n730) );
  OAI22_X1 U1904 ( .A1(n1374), .A2(n931), .B1(n930), .B2(n1513), .ZN(n728) );
  OAI22_X1 U1905 ( .A1(n1266), .A2(n932), .B1(n931), .B2(n1513), .ZN(n729) );
  OAI22_X1 U1906 ( .A1(n1326), .A2(n934), .B1(n933), .B2(n1513), .ZN(n731) );
  OAI22_X1 U1907 ( .A1(n1266), .A2(n939), .B1(n938), .B2(n1513), .ZN(n736) );
  OAI22_X1 U1908 ( .A1(n1326), .A2(n936), .B1(n935), .B2(n1513), .ZN(n733) );
  OAI22_X1 U1909 ( .A1(n1375), .A2(n940), .B1(n1513), .B2(n939), .ZN(n737) );
  OAI22_X1 U1910 ( .A1(n1326), .A2(n935), .B1(n934), .B2(n1513), .ZN(n732) );
  OAI22_X1 U1911 ( .A1(n1374), .A2(n1142), .B1(n942), .B2(n1513), .ZN(n672) );
  OAI22_X1 U1912 ( .A1(n1327), .A2(n937), .B1(n936), .B2(n1513), .ZN(n734) );
  OAI22_X1 U1913 ( .A1(n1327), .A2(n941), .B1(n940), .B2(n1513), .ZN(n738) );
  OAI22_X1 U1914 ( .A1(n1374), .A2(n938), .B1(n937), .B2(n1513), .ZN(n735) );
  XNOR2_X1 U1915 ( .A(n90), .B(n247), .ZN(product[6]) );
  OAI22_X1 U1916 ( .A1(n1535), .A2(n1034), .B1(n1033), .B2(n1517), .ZN(n826)
         );
  OAI22_X1 U1917 ( .A1(n1536), .A2(n1039), .B1(n1038), .B2(n1518), .ZN(n831)
         );
  OAI22_X1 U1918 ( .A1(n1536), .A2(n1031), .B1(n1030), .B2(n1518), .ZN(n823)
         );
  OAI22_X1 U1919 ( .A1(n1536), .A2(n1032), .B1(n1031), .B2(n1518), .ZN(n824)
         );
  OAI22_X1 U1920 ( .A1(n1536), .A2(n1041), .B1(n1040), .B2(n1518), .ZN(n833)
         );
  OAI22_X1 U1921 ( .A1(n1536), .A2(n1045), .B1(n1044), .B2(n1517), .ZN(n837)
         );
  OAI22_X1 U1922 ( .A1(n1536), .A2(n1028), .B1(n1027), .B2(n1518), .ZN(n424)
         );
  OAI22_X1 U1923 ( .A1(n1535), .A2(n1037), .B1(n1036), .B2(n1517), .ZN(n829)
         );
  OAI22_X1 U1924 ( .A1(n1535), .A2(n1044), .B1(n1043), .B2(n1517), .ZN(n836)
         );
  OAI22_X1 U1925 ( .A1(n1536), .A2(n1038), .B1(n1037), .B2(n1517), .ZN(n830)
         );
  OAI22_X1 U1926 ( .A1(n1537), .A2(n1035), .B1(n1034), .B2(n1518), .ZN(n827)
         );
  OAI22_X1 U1927 ( .A1(n1027), .A2(n1535), .B1(n1027), .B2(n1517), .ZN(n661)
         );
  OAI22_X1 U1928 ( .A1(n1535), .A2(n1030), .B1(n1029), .B2(n1517), .ZN(n822)
         );
  OAI22_X1 U1929 ( .A1(n1537), .A2(n1036), .B1(n1035), .B2(n1518), .ZN(n828)
         );
  OAI22_X1 U1930 ( .A1(n1535), .A2(n1147), .B1(n1047), .B2(n1517), .ZN(n677)
         );
  OAI22_X1 U1931 ( .A1(n1537), .A2(n1033), .B1(n1032), .B2(n1518), .ZN(n825)
         );
  OAI22_X1 U1932 ( .A1(n1535), .A2(n1029), .B1(n1028), .B2(n1517), .ZN(n821)
         );
  OAI22_X1 U1933 ( .A1(n1535), .A2(n1040), .B1(n1039), .B2(n1517), .ZN(n832)
         );
  OAI22_X1 U1934 ( .A1(n1535), .A2(n1043), .B1(n1042), .B2(n1518), .ZN(n835)
         );
  OAI22_X1 U1935 ( .A1(n1535), .A2(n1042), .B1(n1041), .B2(n1517), .ZN(n834)
         );
  OAI22_X1 U1936 ( .A1(n1536), .A2(n1046), .B1(n1045), .B2(n1518), .ZN(n838)
         );
  OAI21_X1 U1937 ( .B1(n152), .B2(n1313), .A(n1381), .ZN(n149) );
  INV_X1 U1938 ( .A(n1313), .ZN(n275) );
  OAI22_X1 U1939 ( .A1(n901), .A2(n1320), .B1(n901), .B2(n1510), .ZN(n643) );
  OAI22_X1 U1940 ( .A1(n1320), .A2(n902), .B1(n901), .B2(n1511), .ZN(n304) );
  OAI22_X1 U1941 ( .A1(n1320), .A2(n903), .B1(n902), .B2(n1510), .ZN(n701) );
  NOR2_X1 U1942 ( .A1(n150), .A2(n1470), .ZN(n145) );
  OAI22_X1 U1943 ( .A1(n1320), .A2(n905), .B1(n904), .B2(n1511), .ZN(n703) );
  OAI22_X1 U1944 ( .A1(n1320), .A2(n904), .B1(n903), .B2(n1510), .ZN(n702) );
  OAI22_X1 U1945 ( .A1(n1320), .A2(n906), .B1(n905), .B2(n1511), .ZN(n704) );
  OAI22_X1 U1946 ( .A1(n1320), .A2(n907), .B1(n906), .B2(n1510), .ZN(n705) );
  OAI22_X1 U1947 ( .A1(n1320), .A2(n908), .B1(n907), .B2(n1511), .ZN(n706) );
  OAI22_X1 U1948 ( .A1(n1320), .A2(n909), .B1(n908), .B2(n1510), .ZN(n707) );
  OAI22_X1 U1949 ( .A1(n1320), .A2(n910), .B1(n909), .B2(n1511), .ZN(n708) );
  OAI22_X1 U1950 ( .A1(n1472), .A2(n911), .B1(n910), .B2(n1510), .ZN(n709) );
  OAI22_X1 U1951 ( .A1(n1472), .A2(n912), .B1(n911), .B2(n1511), .ZN(n710) );
  OAI22_X1 U1952 ( .A1(n1472), .A2(n913), .B1(n912), .B2(n1510), .ZN(n711) );
  OAI22_X1 U1953 ( .A1(n1472), .A2(n915), .B1(n914), .B2(n1510), .ZN(n713) );
  OAI22_X1 U1954 ( .A1(n1472), .A2(n1141), .B1(n921), .B2(n1511), .ZN(n671) );
  OAI22_X1 U1955 ( .A1(n1471), .A2(n914), .B1(n913), .B2(n1511), .ZN(n712) );
  OAI22_X1 U1956 ( .A1(n1471), .A2(n919), .B1(n918), .B2(n1510), .ZN(n717) );
  OAI22_X1 U1957 ( .A1(n1471), .A2(n920), .B1(n919), .B2(n1510), .ZN(n718) );
  OAI22_X1 U1958 ( .A1(n1471), .A2(n918), .B1(n917), .B2(n1511), .ZN(n716) );
  INV_X1 U1959 ( .A(n1510), .ZN(n644) );
  OAI22_X1 U1960 ( .A1(n1471), .A2(n917), .B1(n916), .B2(n1511), .ZN(n715) );
  OAI22_X1 U1961 ( .A1(n1472), .A2(n916), .B1(n915), .B2(n1510), .ZN(n714) );
  INV_X1 U1962 ( .A(n1464), .ZN(n152) );
  AOI21_X1 U1963 ( .B1(n1464), .B2(n126), .A(n1438), .ZN(n125) );
  OAI22_X1 U1964 ( .A1(n985), .A2(n1475), .B1(n985), .B2(n1466), .ZN(n655) );
  OAI22_X1 U1965 ( .A1(n1310), .A2(n986), .B1(n985), .B2(n1467), .ZN(n368) );
  OAI22_X1 U1966 ( .A1(n1311), .A2(n987), .B1(n986), .B2(n1466), .ZN(n781) );
  OAI22_X1 U1967 ( .A1(n1310), .A2(n992), .B1(n991), .B2(n1467), .ZN(n786) );
  OAI22_X1 U1968 ( .A1(n1311), .A2(n989), .B1(n988), .B2(n1467), .ZN(n783) );
  OAI22_X1 U1969 ( .A1(n1475), .A2(n990), .B1(n989), .B2(n1467), .ZN(n784) );
  OAI22_X1 U1970 ( .A1(n1310), .A2(n1003), .B1(n1002), .B2(n1467), .ZN(n797)
         );
  OAI22_X1 U1971 ( .A1(n1310), .A2(n988), .B1(n987), .B2(n1467), .ZN(n782) );
  OAI22_X1 U1972 ( .A1(n1475), .A2(n991), .B1(n990), .B2(n1466), .ZN(n785) );
  OAI22_X1 U1973 ( .A1(n1310), .A2(n996), .B1(n995), .B2(n1467), .ZN(n790) );
  OAI22_X1 U1974 ( .A1(n1310), .A2(n999), .B1(n998), .B2(n1466), .ZN(n793) );
  OAI22_X1 U1975 ( .A1(n994), .A2(n1474), .B1(n993), .B2(n1514), .ZN(n788) );
  OAI22_X1 U1976 ( .A1(n1311), .A2(n1323), .B1(n992), .B2(n1466), .ZN(n787) );
  OAI22_X1 U1977 ( .A1(n1474), .A2(n995), .B1(n1350), .B2(n1467), .ZN(n789) );
  OAI22_X1 U1978 ( .A1(n1310), .A2(n1000), .B1(n999), .B2(n1466), .ZN(n794) );
  OAI22_X1 U1979 ( .A1(n997), .A2(n1311), .B1(n996), .B2(n1467), .ZN(n791) );
  OAI22_X1 U1980 ( .A1(n1310), .A2(n1002), .B1(n1001), .B2(n1467), .ZN(n796)
         );
  OAI22_X1 U1981 ( .A1(n1475), .A2(n998), .B1(n997), .B2(n1466), .ZN(n792) );
  OAI22_X1 U1982 ( .A1(n1311), .A2(n1004), .B1(n1003), .B2(n1466), .ZN(n798)
         );
  INV_X1 U1983 ( .A(n1466), .ZN(n656) );
  OAI22_X1 U1984 ( .A1(n1475), .A2(n1145), .B1(n1005), .B2(n1466), .ZN(n675)
         );
  OAI22_X1 U1985 ( .A1(n1311), .A2(n1001), .B1(n1000), .B2(n1466), .ZN(n795)
         );
  OAI21_X1 U1986 ( .B1(n152), .B2(n131), .A(n1462), .ZN(n130) );
  OAI22_X1 U1987 ( .A1(n880), .A2(n1460), .B1(n880), .B2(n1294), .ZN(n640) );
  OAI22_X1 U1988 ( .A1(n1460), .A2(n881), .B1(n880), .B2(n1519), .ZN(n298) );
  OAI22_X1 U1989 ( .A1(n1460), .A2(n882), .B1(n881), .B2(n1295), .ZN(n681) );
  OAI22_X1 U1990 ( .A1(n1460), .A2(n883), .B1(n882), .B2(n1519), .ZN(n682) );
  OAI22_X1 U1991 ( .A1(n1460), .A2(n884), .B1(n883), .B2(n1295), .ZN(n683) );
  OAI21_X1 U1992 ( .B1(n132), .B2(n128), .A(n129), .ZN(n127) );
  OAI22_X1 U1993 ( .A1(n1460), .A2(n886), .B1(n885), .B2(n1519), .ZN(n685) );
  OAI22_X1 U1994 ( .A1(n1460), .A2(n885), .B1(n884), .B2(n1295), .ZN(n684) );
  OAI22_X1 U1995 ( .A1(n1460), .A2(n887), .B1(n886), .B2(n1519), .ZN(n686) );
  OAI22_X1 U1996 ( .A1(n1460), .A2(n888), .B1(n887), .B2(n1295), .ZN(n687) );
  OAI22_X1 U1997 ( .A1(n1460), .A2(n889), .B1(n888), .B2(n1519), .ZN(n688) );
  OAI22_X1 U1998 ( .A1(n1460), .A2(n890), .B1(n889), .B2(n1295), .ZN(n689) );
  OAI22_X1 U1999 ( .A1(n60), .A2(n891), .B1(n890), .B2(n1295), .ZN(n690) );
  OAI22_X1 U2000 ( .A1(n60), .A2(n892), .B1(n891), .B2(n1519), .ZN(n691) );
  OAI22_X1 U2001 ( .A1(n60), .A2(n894), .B1(n893), .B2(n1295), .ZN(n693) );
  OAI22_X1 U2002 ( .A1(n60), .A2(n899), .B1(n898), .B2(n1295), .ZN(n698) );
  OAI22_X1 U2003 ( .A1(n60), .A2(n893), .B1(n892), .B2(n1519), .ZN(n692) );
  OAI22_X1 U2004 ( .A1(n60), .A2(n895), .B1(n894), .B2(n1519), .ZN(n694) );
  OAI22_X1 U2005 ( .A1(n60), .A2(n1140), .B1(n900), .B2(n1295), .ZN(n670) );
  INV_X1 U2006 ( .A(n1294), .ZN(n641) );
  OAI22_X1 U2007 ( .A1(n60), .A2(n898), .B1(n897), .B2(n1295), .ZN(n697) );
  OAI22_X1 U2008 ( .A1(n60), .A2(n896), .B1(n895), .B2(n1519), .ZN(n695) );
  OAI22_X1 U2009 ( .A1(n60), .A2(n897), .B1(n896), .B2(n1294), .ZN(n696) );
  NAND2_X2 U2010 ( .A1(n1110), .A2(n58), .ZN(n60) );
  AOI21_X1 U2011 ( .B1(n194), .B2(n175), .A(n176), .ZN(n174) );
  AOI21_X1 U2012 ( .B1(n165), .B2(n156), .A(n157), .ZN(n155) );
  INV_X1 U2013 ( .A(n1399), .ZN(n173) );
  OAI21_X1 U2014 ( .B1(n174), .B2(n154), .A(n155), .ZN(n153) );
  OAI22_X1 U2015 ( .A1(n1533), .A2(n965), .B1(n964), .B2(n1309), .ZN(n346) );
  OAI22_X1 U2016 ( .A1(n964), .A2(n1477), .B1(n964), .B2(n1516), .ZN(n652) );
  OAI22_X1 U2017 ( .A1(n1532), .A2(n966), .B1(n965), .B2(n1309), .ZN(n761) );
  OAI22_X1 U2018 ( .A1(n1477), .A2(n967), .B1(n966), .B2(n1516), .ZN(n762) );
  OAI22_X1 U2019 ( .A1(n1533), .A2(n968), .B1(n967), .B2(n1309), .ZN(n763) );
  OAI22_X1 U2020 ( .A1(n1532), .A2(n972), .B1(n971), .B2(n1516), .ZN(n767) );
  OAI22_X1 U2021 ( .A1(n1477), .A2(n973), .B1(n972), .B2(n1309), .ZN(n768) );
  OAI22_X1 U2022 ( .A1(n1533), .A2(n975), .B1(n974), .B2(n1309), .ZN(n770) );
  OAI22_X1 U2023 ( .A1(n1532), .A2(n969), .B1(n968), .B2(n1516), .ZN(n764) );
  OAI22_X1 U2024 ( .A1(n1532), .A2(n971), .B1(n970), .B2(n1309), .ZN(n766) );
  OAI22_X1 U2025 ( .A1(n1533), .A2(n970), .B1(n969), .B2(n1309), .ZN(n765) );
  OAI22_X1 U2026 ( .A1(n1534), .A2(n978), .B1(n977), .B2(n1308), .ZN(n773) );
  OAI22_X1 U2027 ( .A1(n1532), .A2(n977), .B1(n976), .B2(n1516), .ZN(n772) );
  OAI22_X1 U2028 ( .A1(n1477), .A2(n1144), .B1(n984), .B2(n1516), .ZN(n674) );
  OAI22_X1 U2029 ( .A1(n1477), .A2(n979), .B1(n978), .B2(n1309), .ZN(n774) );
  OAI22_X1 U2030 ( .A1(n1477), .A2(n976), .B1(n975), .B2(n1516), .ZN(n771) );
  OAI22_X1 U2031 ( .A1(n1532), .A2(n974), .B1(n973), .B2(n1516), .ZN(n769) );
  OAI22_X1 U2032 ( .A1(n1533), .A2(n983), .B1(n982), .B2(n1516), .ZN(n778) );
  OAI22_X1 U2033 ( .A1(n1533), .A2(n982), .B1(n981), .B2(n1309), .ZN(n777) );
  OAI22_X1 U2034 ( .A1(n1534), .A2(n980), .B1(n979), .B2(n1516), .ZN(n775) );
  INV_X1 U2035 ( .A(n1516), .ZN(n653) );
  OAI22_X1 U2036 ( .A1(n1534), .A2(n981), .B1(n980), .B2(n1308), .ZN(n776) );
  OAI21_X1 U2037 ( .B1(n193), .B2(n180), .A(n1461), .ZN(n179) );
  INV_X1 U2038 ( .A(n101), .ZN(n264) );
  OAI21_X1 U2039 ( .B1(n181), .B2(n177), .A(n178), .ZN(n176) );
  XNOR2_X1 U2040 ( .A(n1465), .B(n67), .ZN(product[29]) );
  OAI22_X1 U2041 ( .A1(n943), .A2(n1469), .B1(n943), .B2(n1454), .ZN(n649) );
  OAI22_X1 U2042 ( .A1(n42), .A2(n944), .B1(n943), .B2(n1454), .ZN(n328) );
  OAI22_X1 U2043 ( .A1(n1469), .A2(n945), .B1(n944), .B2(n1454), .ZN(n741) );
  OAI22_X1 U2044 ( .A1(n42), .A2(n947), .B1(n946), .B2(n1454), .ZN(n743) );
  OAI22_X1 U2045 ( .A1(n1244), .A2(n946), .B1(n945), .B2(n1454), .ZN(n742) );
  OAI22_X1 U2046 ( .A1(n1244), .A2(n948), .B1(n947), .B2(n1454), .ZN(n744) );
  OAI22_X1 U2047 ( .A1(n1244), .A2(n949), .B1(n948), .B2(n1297), .ZN(n745) );
  OAI22_X1 U2048 ( .A1(n1244), .A2(n952), .B1(n951), .B2(n1297), .ZN(n748) );
  OAI22_X1 U2049 ( .A1(n1244), .A2(n957), .B1(n956), .B2(n1297), .ZN(n753) );
  OAI22_X1 U2050 ( .A1(n1244), .A2(n951), .B1(n950), .B2(n1297), .ZN(n747) );
  OAI22_X1 U2051 ( .A1(n1469), .A2(n950), .B1(n949), .B2(n1297), .ZN(n746) );
  OAI22_X1 U2052 ( .A1(n42), .A2(n953), .B1(n952), .B2(n1297), .ZN(n749) );
  OAI22_X1 U2053 ( .A1(n42), .A2(n956), .B1(n955), .B2(n1508), .ZN(n752) );
  OAI22_X1 U2054 ( .A1(n1244), .A2(n958), .B1(n957), .B2(n1297), .ZN(n754) );
  OAI22_X1 U2055 ( .A1(n42), .A2(n955), .B1(n954), .B2(n1297), .ZN(n751) );
  OAI22_X1 U2056 ( .A1(n1469), .A2(n1143), .B1(n963), .B2(n1297), .ZN(n673) );
  OAI22_X1 U2057 ( .A1(n1469), .A2(n954), .B1(n953), .B2(n1297), .ZN(n750) );
  OAI22_X1 U2058 ( .A1(n1469), .A2(n961), .B1(n960), .B2(n1297), .ZN(n757) );
  OAI22_X1 U2059 ( .A1(n1244), .A2(n960), .B1(n959), .B2(n1297), .ZN(n756) );
  INV_X1 U2060 ( .A(n1508), .ZN(n650) );
  OAI22_X1 U2061 ( .A1(n1469), .A2(n962), .B1(n961), .B2(n1508), .ZN(n758) );
  OAI22_X1 U2062 ( .A1(n42), .A2(n959), .B1(n958), .B2(n1297), .ZN(n755) );
  XNOR2_X1 U2063 ( .A(n1445), .B(n65), .ZN(product[31]) );
  OAI22_X1 U2064 ( .A1(n1457), .A2(n1007), .B1(n1006), .B2(n1512), .ZN(n394)
         );
  OAI22_X1 U2065 ( .A1(n1303), .A2(n1014), .B1(n1299), .B2(n1306), .ZN(n807)
         );
  OAI22_X1 U2066 ( .A1(n1006), .A2(n1303), .B1(n1006), .B2(n1306), .ZN(n658)
         );
  OAI22_X1 U2067 ( .A1(n1457), .A2(n1317), .B1(n1011), .B2(n1251), .ZN(n805)
         );
  OAI22_X1 U2068 ( .A1(n1457), .A2(n1008), .B1(n1007), .B2(n1512), .ZN(n801)
         );
  OAI22_X1 U2069 ( .A1(n1457), .A2(n1009), .B1(n1008), .B2(n1251), .ZN(n802)
         );
  OAI22_X1 U2070 ( .A1(n1303), .A2(n1024), .B1(n1023), .B2(n1306), .ZN(n817)
         );
  OAI22_X1 U2071 ( .A1(n1457), .A2(n1021), .B1(n1020), .B2(n1306), .ZN(n814)
         );
  OAI22_X1 U2072 ( .A1(n1457), .A2(n1010), .B1(n1009), .B2(n1512), .ZN(n803)
         );
  OAI22_X1 U2073 ( .A1(n1457), .A2(n1015), .B1(n1014), .B2(n1512), .ZN(n808)
         );
  OAI22_X1 U2074 ( .A1(n1457), .A2(n1146), .B1(n1026), .B2(n1306), .ZN(n676)
         );
  OAI22_X1 U2075 ( .A1(n1013), .A2(n1456), .B1(n1012), .B2(n1512), .ZN(n806)
         );
  OAI22_X1 U2076 ( .A1(n1457), .A2(n1025), .B1(n1024), .B2(n1306), .ZN(n818)
         );
  OAI22_X1 U2077 ( .A1(n1456), .A2(n1011), .B1(n1010), .B2(n1512), .ZN(n804)
         );
  OAI22_X1 U2078 ( .A1(n1457), .A2(n1019), .B1(n1018), .B2(n1512), .ZN(n812)
         );
  OAI22_X1 U2079 ( .A1(n1457), .A2(n1020), .B1(n1019), .B2(n1512), .ZN(n813)
         );
  OAI22_X1 U2080 ( .A1(n1457), .A2(n1018), .B1(n1017), .B2(n1512), .ZN(n811)
         );
  OAI22_X1 U2081 ( .A1(n1457), .A2(n1023), .B1(n1022), .B2(n1251), .ZN(n816)
         );
  OAI22_X1 U2082 ( .A1(n1457), .A2(n1017), .B1(n1016), .B2(n1512), .ZN(n810)
         );
  OAI22_X1 U2083 ( .A1(n1456), .A2(n1016), .B1(n1015), .B2(n1512), .ZN(n809)
         );
  OAI22_X1 U2084 ( .A1(n1456), .A2(n1022), .B1(n1021), .B2(n1512), .ZN(n815)
         );
  INV_X1 U2085 ( .A(n1512), .ZN(n659) );
  OAI21_X1 U2086 ( .B1(n248), .B2(n250), .A(n249), .ZN(n247) );
  AOI21_X1 U2087 ( .B1(n1445), .B2(n1492), .A(n111), .ZN(n109) );
  OAI21_X1 U2088 ( .B1(n1473), .B2(n123), .A(n124), .ZN(n122) );
  AOI21_X1 U2089 ( .B1(n1465), .B2(n1491), .A(n119), .ZN(n117) );
  XNOR2_X1 U2090 ( .A(n1400), .B(n63), .ZN(product[33]) );
  XOR2_X1 U2091 ( .A(n109), .B(n64), .Z(product[32]) );
  XOR2_X1 U2092 ( .A(n117), .B(n66), .Z(product[30]) );
  XOR2_X1 U2093 ( .A(n125), .B(n68), .Z(product[28]) );
  AOI21_X1 U2094 ( .B1(n106), .B2(n1490), .A(n103), .ZN(n101) );
  OAI21_X1 U2095 ( .B1(n1463), .B2(n107), .A(n108), .ZN(n106) );
  OAI21_X1 U2096 ( .B1(n1468), .B2(n115), .A(n116), .ZN(n114) );
  OAI22_X1 U2097 ( .A1(n1405), .A2(n1055), .B1(n1054), .B2(n1503), .ZN(n846)
         );
  OAI22_X1 U2098 ( .A1(n1405), .A2(n1051), .B1(n1050), .B2(n1504), .ZN(n842)
         );
  OAI22_X1 U2099 ( .A1(n1404), .A2(n1062), .B1(n1061), .B2(n1503), .ZN(n853)
         );
  OAI22_X1 U2100 ( .A1(n1242), .A2(n1059), .B1(n1058), .B2(n1504), .ZN(n850)
         );
  OAI22_X1 U2101 ( .A1(n1242), .A2(n1060), .B1(n1059), .B2(n1504), .ZN(n851)
         );
  OAI22_X1 U2102 ( .A1(n1242), .A2(n1053), .B1(n1052), .B2(n1504), .ZN(n844)
         );
  OAI22_X1 U2103 ( .A1(n1242), .A2(n1052), .B1(n1051), .B2(n1504), .ZN(n843)
         );
  OAI22_X1 U2104 ( .A1(n1405), .A2(n1063), .B1(n1062), .B2(n1504), .ZN(n854)
         );
  OAI22_X1 U2105 ( .A1(n1404), .A2(n1050), .B1(n1049), .B2(n1504), .ZN(n841)
         );
  OAI22_X1 U2106 ( .A1(n1242), .A2(n1057), .B1(n1056), .B2(n1504), .ZN(n848)
         );
  OAI22_X1 U2107 ( .A1(n1242), .A2(n1065), .B1(n1064), .B2(n1503), .ZN(n856)
         );
  OAI22_X1 U2108 ( .A1(n1405), .A2(n1056), .B1(n1055), .B2(n1503), .ZN(n847)
         );
  OAI22_X1 U2109 ( .A1(n1404), .A2(n1058), .B1(n1057), .B2(n1504), .ZN(n849)
         );
  OAI22_X1 U2110 ( .A1(n1242), .A2(n1148), .B1(n1068), .B2(n1503), .ZN(n678)
         );
  OAI22_X1 U2111 ( .A1(n12), .A2(n1054), .B1(n1053), .B2(n1504), .ZN(n845) );
  OAI22_X1 U2112 ( .A1(n1242), .A2(n1061), .B1(n1060), .B2(n1503), .ZN(n852)
         );
  OAI22_X1 U2113 ( .A1(n1233), .A2(n12), .B1(n1048), .B2(n1503), .ZN(n664) );
  OAI22_X1 U2114 ( .A1(n1242), .A2(n1064), .B1(n1063), .B2(n1504), .ZN(n855)
         );
  OAI22_X1 U2115 ( .A1(n1405), .A2(n1067), .B1(n1066), .B2(n1504), .ZN(n858)
         );
  OAI22_X1 U2116 ( .A1(n1404), .A2(n1066), .B1(n1065), .B2(n1503), .ZN(n857)
         );
  INV_X1 U2117 ( .A(n1503), .ZN(n665) );
endmodule


module mac_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n34, n35, n36, n37, n38, n39, n40, n41, n43, n45, n46, n47,
         n48, n49, n51, n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65,
         n67, n69, n70, n71, n72, n73, n75, n77, n78, n79, n80, n81, n83, n85,
         n86, n87, n88, n89, n91, n93, n94, n95, n96, n97, n99, n101, n102,
         n103, n104, n105, n107, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n119, n121, n122, n124, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n184, n185, n187, n189, n191,
         n193, n195, n197, n199, n201, n203, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405;

  FA_X1 U3 ( .A(B[38]), .B(A[38]), .CI(n35), .CO(n34), .S(SUM[38]) );
  FA_X1 U7 ( .A(B[34]), .B(A[34]), .CI(n39), .CO(n38), .S(SUM[34]) );
  NAND2_X1 U254 ( .A1(B[8]), .A2(A[8]), .ZN(n148) );
  OR2_X1 U255 ( .A1(B[0]), .A2(A[0]), .ZN(n344) );
  XOR2_X1 U256 ( .A(B[35]), .B(A[35]), .Z(n345) );
  XOR2_X1 U257 ( .A(n38), .B(n345), .Z(SUM[35]) );
  NAND2_X1 U258 ( .A1(n38), .A2(B[35]), .ZN(n346) );
  NAND2_X1 U259 ( .A1(n38), .A2(A[35]), .ZN(n347) );
  NAND2_X1 U260 ( .A1(B[35]), .A2(A[35]), .ZN(n348) );
  NAND3_X1 U261 ( .A1(n346), .A2(n347), .A3(n348), .ZN(n37) );
  CLKBUF_X1 U262 ( .A(n36), .Z(n349) );
  XOR2_X1 U263 ( .A(B[36]), .B(A[36]), .Z(n350) );
  XOR2_X1 U264 ( .A(n37), .B(n350), .Z(SUM[36]) );
  NAND2_X1 U265 ( .A1(n37), .A2(B[36]), .ZN(n351) );
  NAND2_X1 U266 ( .A1(n37), .A2(A[36]), .ZN(n352) );
  NAND2_X1 U267 ( .A1(B[36]), .A2(A[36]), .ZN(n353) );
  NAND3_X1 U268 ( .A1(n351), .A2(n352), .A3(n353), .ZN(n36) );
  XOR2_X1 U269 ( .A(B[37]), .B(A[37]), .Z(n354) );
  XOR2_X1 U270 ( .A(n349), .B(n354), .Z(SUM[37]) );
  NAND2_X1 U271 ( .A1(n36), .A2(B[37]), .ZN(n355) );
  NAND2_X1 U272 ( .A1(n36), .A2(A[37]), .ZN(n356) );
  NAND2_X1 U273 ( .A1(B[37]), .A2(A[37]), .ZN(n357) );
  NAND3_X1 U274 ( .A1(n355), .A2(n356), .A3(n357), .ZN(n35) );
  CLKBUF_X1 U275 ( .A(n185), .Z(n358) );
  CLKBUF_X1 U276 ( .A(n94), .Z(n359) );
  NOR2_X1 U277 ( .A1(B[7]), .A2(A[7]), .ZN(n360) );
  CLKBUF_X1 U278 ( .A(n143), .Z(n361) );
  NOR2_X1 U279 ( .A1(B[11]), .A2(A[11]), .ZN(n362) );
  NOR2_X1 U280 ( .A1(B[11]), .A2(A[11]), .ZN(n132) );
  NAND3_X1 U281 ( .A1(n383), .A2(n384), .A3(n385), .ZN(n363) );
  NAND3_X1 U282 ( .A1(n383), .A2(n384), .A3(n385), .ZN(n364) );
  AOI21_X1 U283 ( .B1(n359), .B2(n396), .A(n91), .ZN(n365) );
  AOI21_X1 U284 ( .B1(n94), .B2(n396), .A(n91), .ZN(n89) );
  NOR2_X1 U285 ( .A1(B[3]), .A2(A[3]), .ZN(n366) );
  CLKBUF_X1 U286 ( .A(n150), .Z(n367) );
  AOI21_X1 U287 ( .B1(n130), .B2(n361), .A(n131), .ZN(n368) );
  CLKBUF_X1 U288 ( .A(n102), .Z(n369) );
  AOI21_X1 U289 ( .B1(n369), .B2(n398), .A(n99), .ZN(n370) );
  CLKBUF_X1 U290 ( .A(n110), .Z(n371) );
  CLKBUF_X1 U291 ( .A(n62), .Z(n372) );
  CLKBUF_X1 U292 ( .A(n70), .Z(n373) );
  XOR2_X1 U293 ( .A(B[33]), .B(A[33]), .Z(n374) );
  XOR2_X1 U294 ( .A(n364), .B(n374), .Z(SUM[33]) );
  NAND2_X1 U295 ( .A1(n363), .A2(B[33]), .ZN(n375) );
  NAND2_X1 U296 ( .A1(n40), .A2(A[33]), .ZN(n376) );
  NAND2_X1 U297 ( .A1(B[33]), .A2(A[33]), .ZN(n377) );
  NAND3_X1 U298 ( .A1(n375), .A2(n376), .A3(n377), .ZN(n39) );
  AOI21_X1 U299 ( .B1(n373), .B2(n401), .A(n67), .ZN(n378) );
  AOI21_X1 U300 ( .B1(n372), .B2(n402), .A(n59), .ZN(n379) );
  AOI21_X1 U301 ( .B1(n371), .B2(n397), .A(n107), .ZN(n380) );
  CLKBUF_X1 U302 ( .A(n78), .Z(n381) );
  XOR2_X1 U303 ( .A(B[32]), .B(A[32]), .Z(n382) );
  XOR2_X1 U304 ( .A(n358), .B(n382), .Z(SUM[32]) );
  NAND2_X1 U305 ( .A1(n185), .A2(B[32]), .ZN(n383) );
  NAND2_X1 U306 ( .A1(n185), .A2(A[32]), .ZN(n384) );
  NAND2_X1 U307 ( .A1(B[32]), .A2(A[32]), .ZN(n385) );
  NAND3_X1 U308 ( .A1(n383), .A2(n384), .A3(n385), .ZN(n40) );
  AOI21_X1 U309 ( .B1(n381), .B2(n399), .A(n75), .ZN(n386) );
  CLKBUF_X1 U310 ( .A(n54), .Z(n387) );
  CLKBUF_X1 U311 ( .A(n86), .Z(n388) );
  CLKBUF_X1 U312 ( .A(n46), .Z(n389) );
  AOI21_X1 U313 ( .B1(n387), .B2(n403), .A(n51), .ZN(n390) );
  AOI21_X1 U314 ( .B1(n388), .B2(n400), .A(n83), .ZN(n391) );
  AOI21_X1 U315 ( .B1(n367), .B2(n114), .A(n115), .ZN(n392) );
  AOI21_X1 U316 ( .B1(n150), .B2(n114), .A(n115), .ZN(n113) );
  NOR2_X1 U317 ( .A1(B[7]), .A2(A[7]), .ZN(n155) );
  NOR2_X1 U318 ( .A1(B[5]), .A2(A[5]), .ZN(n163) );
  NOR2_X1 U319 ( .A1(B[6]), .A2(A[6]), .ZN(n158) );
  NOR2_X1 U320 ( .A1(B[10]), .A2(A[10]), .ZN(n137) );
  OR2_X1 U321 ( .A1(B[13]), .A2(A[13]), .ZN(n395) );
  OR2_X1 U322 ( .A1(B[12]), .A2(A[12]), .ZN(n394) );
  INV_X1 U323 ( .A(n367), .ZN(n149) );
  OAI21_X1 U324 ( .B1(n149), .B2(n128), .A(n368), .ZN(n127) );
  OAI21_X1 U325 ( .B1(n149), .B2(n140), .A(n141), .ZN(n139) );
  INV_X1 U326 ( .A(n361), .ZN(n141) );
  INV_X1 U327 ( .A(n142), .ZN(n140) );
  NAND2_X1 U328 ( .A1(n142), .A2(n130), .ZN(n128) );
  AOI21_X1 U329 ( .B1(n170), .B2(n161), .A(n162), .ZN(n160) );
  INV_X1 U330 ( .A(n171), .ZN(n170) );
  INV_X1 U331 ( .A(n180), .ZN(n179) );
  INV_X1 U332 ( .A(n85), .ZN(n83) );
  INV_X1 U333 ( .A(n61), .ZN(n59) );
  INV_X1 U334 ( .A(n53), .ZN(n51) );
  AOI21_X1 U335 ( .B1(n143), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U336 ( .B1(n132), .B2(n138), .A(n133), .ZN(n131) );
  AOI21_X1 U337 ( .B1(n78), .B2(n399), .A(n75), .ZN(n73) );
  INV_X1 U338 ( .A(n77), .ZN(n75) );
  AOI21_X1 U339 ( .B1(n110), .B2(n397), .A(n107), .ZN(n105) );
  INV_X1 U340 ( .A(n109), .ZN(n107) );
  AOI21_X1 U341 ( .B1(n102), .B2(n398), .A(n99), .ZN(n97) );
  INV_X1 U342 ( .A(n101), .ZN(n99) );
  OAI21_X1 U343 ( .B1(n163), .B2(n169), .A(n164), .ZN(n162) );
  AOI21_X1 U344 ( .B1(n172), .B2(n180), .A(n173), .ZN(n171) );
  NOR2_X1 U345 ( .A1(n177), .A2(n366), .ZN(n172) );
  OAI21_X1 U346 ( .B1(n174), .B2(n178), .A(n175), .ZN(n173) );
  AOI21_X1 U347 ( .B1(n70), .B2(n401), .A(n67), .ZN(n65) );
  INV_X1 U348 ( .A(n69), .ZN(n67) );
  INV_X1 U349 ( .A(n93), .ZN(n91) );
  OAI21_X1 U350 ( .B1(n144), .B2(n148), .A(n145), .ZN(n143) );
  NOR2_X1 U351 ( .A1(n168), .A2(n163), .ZN(n161) );
  OAI21_X1 U352 ( .B1(n181), .B2(n184), .A(n182), .ZN(n180) );
  NOR2_X1 U353 ( .A1(n137), .A2(n362), .ZN(n130) );
  OAI21_X1 U354 ( .B1(n171), .B2(n151), .A(n152), .ZN(n150) );
  NAND2_X1 U355 ( .A1(n161), .A2(n153), .ZN(n151) );
  AOI21_X1 U356 ( .B1(n153), .B2(n162), .A(n154), .ZN(n152) );
  NOR2_X1 U357 ( .A1(n158), .A2(n360), .ZN(n153) );
  AOI21_X1 U358 ( .B1(n395), .B2(n124), .A(n119), .ZN(n117) );
  INV_X1 U359 ( .A(n121), .ZN(n119) );
  NAND2_X1 U360 ( .A1(n195), .A2(n80), .ZN(n11) );
  INV_X1 U361 ( .A(n79), .ZN(n195) );
  NAND2_X1 U362 ( .A1(n197), .A2(n88), .ZN(n13) );
  INV_X1 U363 ( .A(n87), .ZN(n197) );
  NOR2_X1 U364 ( .A1(n128), .A2(n116), .ZN(n114) );
  OAI21_X1 U365 ( .B1(n129), .B2(n116), .A(n117), .ZN(n115) );
  NAND2_X1 U366 ( .A1(n394), .A2(n395), .ZN(n116) );
  NOR2_X1 U367 ( .A1(n147), .A2(n144), .ZN(n142) );
  INV_X1 U368 ( .A(n126), .ZN(n124) );
  OAI21_X1 U369 ( .B1(n155), .B2(n159), .A(n156), .ZN(n154) );
  NAND2_X1 U370 ( .A1(n187), .A2(n48), .ZN(n3) );
  INV_X1 U371 ( .A(n47), .ZN(n187) );
  NAND2_X1 U372 ( .A1(n189), .A2(n56), .ZN(n5) );
  INV_X1 U373 ( .A(n55), .ZN(n189) );
  NAND2_X1 U374 ( .A1(n191), .A2(n64), .ZN(n7) );
  INV_X1 U375 ( .A(n63), .ZN(n191) );
  NAND2_X1 U376 ( .A1(n404), .A2(n45), .ZN(n2) );
  NAND2_X1 U377 ( .A1(n403), .A2(n53), .ZN(n4) );
  NAND2_X1 U378 ( .A1(n402), .A2(n61), .ZN(n6) );
  NAND2_X1 U379 ( .A1(n401), .A2(n69), .ZN(n8) );
  XOR2_X1 U380 ( .A(n386), .B(n9), .Z(SUM[24]) );
  NAND2_X1 U381 ( .A1(n193), .A2(n72), .ZN(n9) );
  INV_X1 U382 ( .A(n71), .ZN(n193) );
  NAND2_X1 U383 ( .A1(n399), .A2(n77), .ZN(n10) );
  NAND2_X1 U384 ( .A1(n400), .A2(n85), .ZN(n12) );
  NAND2_X1 U385 ( .A1(n396), .A2(n93), .ZN(n14) );
  XOR2_X1 U386 ( .A(n370), .B(n15), .Z(SUM[18]) );
  NAND2_X1 U387 ( .A1(n199), .A2(n96), .ZN(n15) );
  INV_X1 U388 ( .A(n95), .ZN(n199) );
  NAND2_X1 U389 ( .A1(n398), .A2(n101), .ZN(n16) );
  XOR2_X1 U390 ( .A(n380), .B(n17), .Z(SUM[16]) );
  NAND2_X1 U391 ( .A1(n201), .A2(n104), .ZN(n17) );
  INV_X1 U392 ( .A(n103), .ZN(n201) );
  XOR2_X1 U393 ( .A(n122), .B(n20), .Z(SUM[13]) );
  NAND2_X1 U394 ( .A1(n395), .A2(n121), .ZN(n20) );
  AOI21_X1 U395 ( .B1(n127), .B2(n394), .A(n124), .ZN(n122) );
  XOR2_X1 U396 ( .A(n134), .B(n22), .Z(SUM[11]) );
  NAND2_X1 U397 ( .A1(n206), .A2(n133), .ZN(n22) );
  AOI21_X1 U398 ( .B1(n139), .B2(n207), .A(n136), .ZN(n134) );
  INV_X1 U399 ( .A(n137), .ZN(n207) );
  INV_X1 U400 ( .A(n168), .ZN(n213) );
  XOR2_X1 U401 ( .A(n160), .B(n27), .Z(SUM[6]) );
  NAND2_X1 U402 ( .A1(n211), .A2(n159), .ZN(n27) );
  INV_X1 U403 ( .A(n158), .ZN(n211) );
  INV_X1 U404 ( .A(n362), .ZN(n206) );
  INV_X1 U405 ( .A(n138), .ZN(n136) );
  INV_X1 U406 ( .A(n169), .ZN(n167) );
  INV_X1 U407 ( .A(n144), .ZN(n208) );
  INV_X1 U408 ( .A(n360), .ZN(n210) );
  INV_X1 U409 ( .A(n163), .ZN(n212) );
  INV_X1 U410 ( .A(n366), .ZN(n214) );
  XOR2_X1 U411 ( .A(n165), .B(n28), .Z(SUM[5]) );
  NAND2_X1 U412 ( .A1(n212), .A2(n164), .ZN(n28) );
  AOI21_X1 U413 ( .B1(n170), .B2(n213), .A(n167), .ZN(n165) );
  XNOR2_X1 U414 ( .A(n170), .B(n29), .ZN(SUM[4]) );
  NAND2_X1 U415 ( .A1(n213), .A2(n169), .ZN(n29) );
  XNOR2_X1 U416 ( .A(n176), .B(n30), .ZN(SUM[3]) );
  NAND2_X1 U417 ( .A1(n214), .A2(n175), .ZN(n30) );
  OAI21_X1 U418 ( .B1(n179), .B2(n177), .A(n178), .ZN(n176) );
  XOR2_X1 U419 ( .A(n179), .B(n31), .Z(SUM[2]) );
  NAND2_X1 U420 ( .A1(n215), .A2(n178), .ZN(n31) );
  INV_X1 U421 ( .A(n177), .ZN(n215) );
  XOR2_X1 U422 ( .A(n32), .B(n184), .Z(SUM[1]) );
  NAND2_X1 U423 ( .A1(n216), .A2(n182), .ZN(n32) );
  INV_X1 U424 ( .A(n181), .ZN(n216) );
  AND2_X1 U425 ( .A1(n344), .A2(n184), .ZN(SUM[0]) );
  NAND2_X1 U426 ( .A1(n203), .A2(n112), .ZN(n19) );
  INV_X1 U427 ( .A(n111), .ZN(n203) );
  NAND2_X1 U428 ( .A1(n397), .A2(n109), .ZN(n18) );
  XNOR2_X1 U429 ( .A(n127), .B(n21), .ZN(SUM[12]) );
  NAND2_X1 U430 ( .A1(n394), .A2(n126), .ZN(n21) );
  XNOR2_X1 U431 ( .A(n139), .B(n23), .ZN(SUM[10]) );
  NAND2_X1 U432 ( .A1(n207), .A2(n138), .ZN(n23) );
  XNOR2_X1 U433 ( .A(n146), .B(n24), .ZN(SUM[9]) );
  NAND2_X1 U434 ( .A1(n208), .A2(n145), .ZN(n24) );
  OAI21_X1 U435 ( .B1(n149), .B2(n147), .A(n148), .ZN(n146) );
  XOR2_X1 U436 ( .A(n149), .B(n25), .Z(SUM[8]) );
  NAND2_X1 U437 ( .A1(n209), .A2(n148), .ZN(n25) );
  INV_X1 U438 ( .A(n147), .ZN(n209) );
  XNOR2_X1 U439 ( .A(n157), .B(n26), .ZN(SUM[7]) );
  NAND2_X1 U440 ( .A1(n210), .A2(n156), .ZN(n26) );
  OAI21_X1 U441 ( .B1(n160), .B2(n158), .A(n159), .ZN(n157) );
  NOR2_X1 U442 ( .A1(B[2]), .A2(A[2]), .ZN(n177) );
  NOR2_X1 U443 ( .A1(B[8]), .A2(A[8]), .ZN(n147) );
  NOR2_X2 U444 ( .A1(B[9]), .A2(A[9]), .ZN(n144) );
  NOR2_X1 U445 ( .A1(B[3]), .A2(A[3]), .ZN(n174) );
  NAND2_X1 U446 ( .A1(B[11]), .A2(A[11]), .ZN(n133) );
  NOR2_X1 U447 ( .A1(B[4]), .A2(A[4]), .ZN(n168) );
  NOR2_X1 U448 ( .A1(B[1]), .A2(A[1]), .ZN(n181) );
  NAND2_X1 U449 ( .A1(B[6]), .A2(A[6]), .ZN(n159) );
  NAND2_X1 U450 ( .A1(B[2]), .A2(A[2]), .ZN(n178) );
  NAND2_X1 U451 ( .A1(B[0]), .A2(A[0]), .ZN(n184) );
  NAND2_X1 U452 ( .A1(B[10]), .A2(A[10]), .ZN(n138) );
  NAND2_X1 U453 ( .A1(B[4]), .A2(A[4]), .ZN(n169) );
  NAND2_X1 U454 ( .A1(B[5]), .A2(A[5]), .ZN(n164) );
  NAND2_X1 U455 ( .A1(B[7]), .A2(A[7]), .ZN(n156) );
  NAND2_X1 U456 ( .A1(B[3]), .A2(A[3]), .ZN(n175) );
  NAND2_X1 U457 ( .A1(B[1]), .A2(A[1]), .ZN(n182) );
  NAND2_X1 U458 ( .A1(B[9]), .A2(A[9]), .ZN(n145) );
  INV_X1 U459 ( .A(n45), .ZN(n43) );
  NOR2_X1 U460 ( .A1(B[20]), .A2(A[20]), .ZN(n87) );
  NOR2_X1 U461 ( .A1(B[18]), .A2(A[18]), .ZN(n95) );
  NOR2_X1 U462 ( .A1(B[14]), .A2(A[14]), .ZN(n111) );
  NOR2_X1 U463 ( .A1(B[16]), .A2(A[16]), .ZN(n103) );
  NOR2_X1 U464 ( .A1(B[30]), .A2(A[30]), .ZN(n47) );
  NOR2_X1 U465 ( .A1(B[28]), .A2(A[28]), .ZN(n55) );
  NOR2_X1 U466 ( .A1(B[26]), .A2(A[26]), .ZN(n63) );
  NOR2_X1 U467 ( .A1(B[24]), .A2(A[24]), .ZN(n71) );
  NOR2_X1 U468 ( .A1(B[22]), .A2(A[22]), .ZN(n79) );
  OR2_X1 U469 ( .A1(B[19]), .A2(A[19]), .ZN(n396) );
  OR2_X1 U470 ( .A1(B[15]), .A2(A[15]), .ZN(n397) );
  OR2_X1 U471 ( .A1(B[17]), .A2(A[17]), .ZN(n398) );
  OR2_X1 U472 ( .A1(B[23]), .A2(A[23]), .ZN(n399) );
  NAND2_X1 U473 ( .A1(B[21]), .A2(A[21]), .ZN(n85) );
  NAND2_X1 U474 ( .A1(B[12]), .A2(A[12]), .ZN(n126) );
  NAND2_X1 U475 ( .A1(B[13]), .A2(A[13]), .ZN(n121) );
  NAND2_X1 U476 ( .A1(B[19]), .A2(A[19]), .ZN(n93) );
  NAND2_X1 U477 ( .A1(B[15]), .A2(A[15]), .ZN(n109) );
  NAND2_X1 U478 ( .A1(B[17]), .A2(A[17]), .ZN(n101) );
  NAND2_X1 U479 ( .A1(B[23]), .A2(A[23]), .ZN(n77) );
  NAND2_X1 U480 ( .A1(B[25]), .A2(A[25]), .ZN(n69) );
  NAND2_X1 U481 ( .A1(B[27]), .A2(A[27]), .ZN(n61) );
  NAND2_X1 U482 ( .A1(B[29]), .A2(A[29]), .ZN(n53) );
  NAND2_X1 U483 ( .A1(B[31]), .A2(A[31]), .ZN(n45) );
  NAND2_X1 U484 ( .A1(B[20]), .A2(A[20]), .ZN(n88) );
  NAND2_X1 U485 ( .A1(B[18]), .A2(A[18]), .ZN(n96) );
  NAND2_X1 U486 ( .A1(B[14]), .A2(A[14]), .ZN(n112) );
  NAND2_X1 U487 ( .A1(B[16]), .A2(A[16]), .ZN(n104) );
  NAND2_X1 U488 ( .A1(B[30]), .A2(A[30]), .ZN(n48) );
  NAND2_X1 U489 ( .A1(B[28]), .A2(A[28]), .ZN(n56) );
  NAND2_X1 U490 ( .A1(B[26]), .A2(A[26]), .ZN(n64) );
  NAND2_X1 U491 ( .A1(B[24]), .A2(A[24]), .ZN(n72) );
  NAND2_X1 U492 ( .A1(B[22]), .A2(A[22]), .ZN(n80) );
  OR2_X1 U493 ( .A1(B[21]), .A2(A[21]), .ZN(n400) );
  OR2_X1 U494 ( .A1(B[25]), .A2(A[25]), .ZN(n401) );
  OR2_X1 U495 ( .A1(B[27]), .A2(A[27]), .ZN(n402) );
  OR2_X1 U496 ( .A1(B[29]), .A2(A[29]), .ZN(n403) );
  OR2_X1 U497 ( .A1(B[31]), .A2(A[31]), .ZN(n404) );
  XNOR2_X1 U498 ( .A(n34), .B(n405), .ZN(SUM[39]) );
  XNOR2_X1 U499 ( .A(A[39]), .B(B[39]), .ZN(n405) );
  XNOR2_X1 U500 ( .A(n372), .B(n6), .ZN(SUM[27]) );
  XNOR2_X1 U501 ( .A(n388), .B(n12), .ZN(SUM[21]) );
  XOR2_X1 U502 ( .A(n378), .B(n7), .Z(SUM[26]) );
  AOI21_X1 U503 ( .B1(n62), .B2(n402), .A(n59), .ZN(n57) );
  OAI21_X1 U504 ( .B1(n65), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X1 U505 ( .B1(n86), .B2(n400), .A(n83), .ZN(n81) );
  XNOR2_X1 U506 ( .A(n369), .B(n16), .ZN(SUM[17]) );
  XOR2_X1 U507 ( .A(n365), .B(n13), .Z(SUM[20]) );
  OAI21_X1 U508 ( .B1(n89), .B2(n87), .A(n88), .ZN(n86) );
  XNOR2_X1 U509 ( .A(n387), .B(n4), .ZN(SUM[29]) );
  XOR2_X1 U510 ( .A(n379), .B(n5), .Z(SUM[28]) );
  XNOR2_X1 U511 ( .A(n359), .B(n14), .ZN(SUM[19]) );
  XNOR2_X1 U512 ( .A(n373), .B(n8), .ZN(SUM[25]) );
  AOI21_X1 U513 ( .B1(n54), .B2(n403), .A(n51), .ZN(n49) );
  OAI21_X1 U514 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  OAI21_X1 U515 ( .B1(n105), .B2(n103), .A(n104), .ZN(n102) );
  OAI21_X1 U516 ( .B1(n97), .B2(n95), .A(n96), .ZN(n94) );
  OAI21_X1 U517 ( .B1(n73), .B2(n71), .A(n72), .ZN(n70) );
  XNOR2_X1 U518 ( .A(n381), .B(n10), .ZN(SUM[23]) );
  XNOR2_X1 U519 ( .A(n371), .B(n18), .ZN(SUM[15]) );
  INV_X1 U520 ( .A(n41), .ZN(n185) );
  XNOR2_X1 U521 ( .A(n389), .B(n2), .ZN(SUM[31]) );
  XOR2_X1 U522 ( .A(n392), .B(n19), .Z(SUM[14]) );
  XOR2_X1 U523 ( .A(n391), .B(n11), .Z(SUM[22]) );
  XOR2_X1 U524 ( .A(n390), .B(n3), .Z(SUM[30]) );
  AOI21_X1 U525 ( .B1(n46), .B2(n404), .A(n43), .ZN(n41) );
  OAI21_X1 U526 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  OAI21_X1 U527 ( .B1(n81), .B2(n79), .A(n80), .ZN(n78) );
  OAI21_X1 U528 ( .B1(n113), .B2(n111), .A(n112), .ZN(n110) );
endmodule


module mac_1 ( clk, clear_acc, a, b, mac_out );
  input [19:0] a;
  input [19:0] b;
  output [39:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, n2, n3;
  wire   [39:0] mul;
  wire   [39:0] pipeline;
  wire   [39:0] sum;

  DFF_X1 \pipeline_reg[37]  ( .D(mul[37]), .CK(clk), .Q(pipeline[37]) );
  DFF_X1 \pipeline_reg[36]  ( .D(mul[36]), .CK(clk), .Q(pipeline[36]) );
  DFF_X1 \pipeline_reg[35]  ( .D(mul[35]), .CK(clk), .Q(pipeline[35]) );
  DFF_X1 \pipeline_reg[34]  ( .D(mul[34]), .CK(clk), .Q(pipeline[34]) );
  DFF_X1 \pipeline_reg[33]  ( .D(mul[33]), .CK(clk), .Q(pipeline[33]) );
  DFF_X1 \pipeline_reg[32]  ( .D(mul[32]), .CK(clk), .Q(pipeline[32]) );
  DFF_X1 \pipeline_reg[31]  ( .D(mul[31]), .CK(clk), .Q(pipeline[31]) );
  DFF_X1 \pipeline_reg[30]  ( .D(mul[30]), .CK(clk), .Q(pipeline[30]) );
  DFF_X1 \pipeline_reg[29]  ( .D(mul[29]), .CK(clk), .Q(pipeline[29]) );
  DFF_X1 \pipeline_reg[28]  ( .D(mul[28]), .CK(clk), .Q(pipeline[28]) );
  DFF_X1 \pipeline_reg[27]  ( .D(mul[27]), .CK(clk), .Q(pipeline[27]) );
  DFF_X1 \pipeline_reg[26]  ( .D(mul[26]), .CK(clk), .Q(pipeline[26]) );
  DFF_X1 \pipeline_reg[25]  ( .D(mul[25]), .CK(clk), .Q(pipeline[25]) );
  DFF_X1 \pipeline_reg[24]  ( .D(mul[24]), .CK(clk), .Q(pipeline[24]) );
  DFF_X1 \pipeline_reg[23]  ( .D(mul[23]), .CK(clk), .Q(pipeline[23]) );
  DFF_X1 \pipeline_reg[22]  ( .D(mul[22]), .CK(clk), .Q(pipeline[22]) );
  DFF_X1 \pipeline_reg[21]  ( .D(mul[21]), .CK(clk), .Q(pipeline[21]) );
  DFF_X1 \pipeline_reg[20]  ( .D(mul[20]), .CK(clk), .Q(pipeline[20]) );
  DFF_X1 \pipeline_reg[19]  ( .D(mul[19]), .CK(clk), .Q(pipeline[19]) );
  DFF_X1 \pipeline_reg[18]  ( .D(mul[18]), .CK(clk), .Q(pipeline[18]) );
  DFF_X1 \pipeline_reg[17]  ( .D(mul[17]), .CK(clk), .Q(pipeline[17]) );
  DFF_X1 \pipeline_reg[16]  ( .D(mul[16]), .CK(clk), .Q(pipeline[16]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \mac_out_reg[16]  ( .D(N19), .CK(clk), .Q(mac_out[16]) );
  DFF_X1 \mac_out_reg[17]  ( .D(N20), .CK(clk), .Q(mac_out[17]) );
  DFF_X1 \mac_out_reg[18]  ( .D(N21), .CK(clk), .Q(mac_out[18]) );
  DFF_X1 \mac_out_reg[19]  ( .D(N22), .CK(clk), .Q(mac_out[19]) );
  DFF_X1 \mac_out_reg[20]  ( .D(N23), .CK(clk), .Q(mac_out[20]) );
  DFF_X1 \mac_out_reg[21]  ( .D(N24), .CK(clk), .Q(mac_out[21]) );
  DFF_X1 \mac_out_reg[22]  ( .D(N25), .CK(clk), .Q(mac_out[22]) );
  DFF_X1 \mac_out_reg[23]  ( .D(N26), .CK(clk), .Q(mac_out[23]) );
  DFF_X1 \mac_out_reg[24]  ( .D(N27), .CK(clk), .Q(mac_out[24]) );
  DFF_X1 \mac_out_reg[25]  ( .D(N28), .CK(clk), .Q(mac_out[25]) );
  DFF_X1 \mac_out_reg[26]  ( .D(N29), .CK(clk), .Q(mac_out[26]) );
  DFF_X1 \mac_out_reg[27]  ( .D(N30), .CK(clk), .Q(mac_out[27]) );
  DFF_X1 \mac_out_reg[28]  ( .D(N31), .CK(clk), .Q(mac_out[28]) );
  DFF_X1 \mac_out_reg[29]  ( .D(N32), .CK(clk), .Q(mac_out[29]) );
  DFF_X1 \mac_out_reg[30]  ( .D(N33), .CK(clk), .Q(mac_out[30]) );
  DFF_X1 \mac_out_reg[31]  ( .D(N34), .CK(clk), .Q(mac_out[31]) );
  DFF_X1 \mac_out_reg[32]  ( .D(N35), .CK(clk), .Q(mac_out[32]) );
  DFF_X1 \mac_out_reg[33]  ( .D(N36), .CK(clk), .Q(mac_out[33]) );
  DFF_X1 \mac_out_reg[34]  ( .D(N37), .CK(clk), .Q(mac_out[34]) );
  DFF_X1 \mac_out_reg[35]  ( .D(N38), .CK(clk), .Q(mac_out[35]) );
  DFF_X1 \mac_out_reg[36]  ( .D(N39), .CK(clk), .Q(mac_out[36]) );
  DFF_X1 \mac_out_reg[37]  ( .D(N40), .CK(clk), .Q(mac_out[37]) );
  DFF_X1 \mac_out_reg[38]  ( .D(N41), .CK(clk), .Q(mac_out[38]) );
  DFF_X1 \mac_out_reg[39]  ( .D(N42), .CK(clk), .Q(mac_out[39]) );
  mac_1_DW_mult_tc_1 mult_355 ( .a(a), .b(b), .product(mul) );
  mac_1_DW01_add_1 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  DFF_X1 \pipeline_reg[38]  ( .D(mul[38]), .CK(clk), .Q(pipeline[38]) );
  DFF_X2 \pipeline_reg[39]  ( .D(mul[39]), .CK(clk), .Q(pipeline[39]) );
  BUF_X1 U3 ( .A(n3), .Z(n2) );
  INV_X1 U4 ( .A(clear_acc), .ZN(n3) );
  AND2_X1 U6 ( .A1(sum[39]), .A2(n2), .ZN(N42) );
  AND2_X1 U7 ( .A1(sum[38]), .A2(n2), .ZN(N41) );
  AND2_X1 U8 ( .A1(sum[37]), .A2(n2), .ZN(N40) );
  AND2_X1 U9 ( .A1(sum[36]), .A2(n2), .ZN(N39) );
  AND2_X1 U10 ( .A1(sum[35]), .A2(n2), .ZN(N38) );
  AND2_X1 U11 ( .A1(sum[34]), .A2(n2), .ZN(N37) );
  AND2_X1 U12 ( .A1(sum[33]), .A2(n2), .ZN(N36) );
  AND2_X1 U13 ( .A1(sum[32]), .A2(n2), .ZN(N35) );
  AND2_X1 U14 ( .A1(sum[31]), .A2(n2), .ZN(N34) );
  AND2_X1 U15 ( .A1(sum[30]), .A2(n2), .ZN(N33) );
  AND2_X1 U16 ( .A1(sum[29]), .A2(n2), .ZN(N32) );
  AND2_X1 U17 ( .A1(sum[28]), .A2(n3), .ZN(N31) );
  AND2_X1 U18 ( .A1(sum[27]), .A2(n3), .ZN(N30) );
  AND2_X1 U19 ( .A1(sum[26]), .A2(n3), .ZN(N29) );
  AND2_X1 U20 ( .A1(sum[25]), .A2(n3), .ZN(N28) );
  AND2_X1 U21 ( .A1(sum[24]), .A2(n3), .ZN(N27) );
  AND2_X1 U22 ( .A1(sum[23]), .A2(n3), .ZN(N26) );
  AND2_X1 U23 ( .A1(sum[22]), .A2(n3), .ZN(N25) );
  AND2_X1 U24 ( .A1(sum[21]), .A2(n3), .ZN(N24) );
  AND2_X1 U25 ( .A1(sum[20]), .A2(n3), .ZN(N23) );
  AND2_X1 U26 ( .A1(sum[19]), .A2(n3), .ZN(N22) );
  AND2_X1 U27 ( .A1(sum[18]), .A2(n3), .ZN(N21) );
  AND2_X1 U28 ( .A1(sum[17]), .A2(n3), .ZN(N20) );
  AND2_X1 U29 ( .A1(sum[16]), .A2(n3), .ZN(N19) );
  AND2_X1 U30 ( .A1(sum[15]), .A2(n3), .ZN(N18) );
  AND2_X1 U31 ( .A1(sum[14]), .A2(n3), .ZN(N17) );
  AND2_X1 U32 ( .A1(sum[13]), .A2(n3), .ZN(N16) );
  AND2_X1 U33 ( .A1(sum[12]), .A2(n3), .ZN(N15) );
  AND2_X1 U34 ( .A1(sum[11]), .A2(n3), .ZN(N14) );
  AND2_X1 U35 ( .A1(sum[10]), .A2(n3), .ZN(N13) );
  AND2_X1 U36 ( .A1(sum[9]), .A2(n3), .ZN(N12) );
  AND2_X1 U37 ( .A1(sum[8]), .A2(n3), .ZN(N11) );
  AND2_X1 U38 ( .A1(sum[7]), .A2(n3), .ZN(N10) );
  AND2_X1 U39 ( .A1(sum[6]), .A2(n3), .ZN(N9) );
  AND2_X1 U40 ( .A1(sum[5]), .A2(n3), .ZN(N8) );
  AND2_X1 U41 ( .A1(sum[4]), .A2(n3), .ZN(N7) );
  AND2_X1 U42 ( .A1(sum[3]), .A2(n3), .ZN(N6) );
  AND2_X1 U43 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U44 ( .A1(sum[1]), .A2(n3), .ZN(N4) );
  AND2_X1 U45 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
endmodule


module mac_0_DW_mult_tc_1 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n4, n7, n9, n12, n13, n18, n19, n22, n24, n25, n30, n31, n34, n36,
         n37, n42, n43, n46, n48, n49, n52, n54, n55, n58, n60, n61, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n97, n98, n99, n100, n101, n103, n105, n106, n107, n108, n109,
         n111, n113, n114, n115, n116, n117, n119, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n185, n186, n187, n188, n190, n193, n194, n195, n196, n198, n200,
         n201, n202, n203, n204, n205, n206, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n227, n228, n230, n232, n233, n234, n236, n238, n239, n240, n241,
         n242, n244, n246, n247, n248, n249, n250, n252, n254, n255, n256,
         n257, n258, n259, n260, n261, n263, n264, n266, n268, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n282, n284,
         n285, n286, n287, n291, n293, n295, n296, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n643,
         n644, n646, n647, n649, n650, n652, n653, n655, n656, n658, n659,
         n661, n664, n665, n667, n668, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1116, n1119, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1233, n1234, n1235, n1236, n1237,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599;
  assign n1 = a[1];
  assign n7 = a[3];
  assign n13 = a[5];
  assign n19 = a[7];
  assign n25 = a[9];
  assign n31 = a[11];
  assign n37 = a[13];
  assign n43 = a[15];
  assign n49 = a[17];
  assign n55 = a[19];
  assign n61 = b[0];
  assign n668 = a[0];
  assign n1090 = b[19];
  assign n1091 = b[18];
  assign n1092 = b[17];
  assign n1093 = b[16];
  assign n1094 = b[15];
  assign n1095 = b[14];
  assign n1096 = b[13];
  assign n1097 = b[12];
  assign n1098 = b[11];
  assign n1099 = b[10];
  assign n1100 = b[9];
  assign n1101 = b[8];
  assign n1102 = b[7];
  assign n1103 = b[6];
  assign n1104 = b[5];
  assign n1105 = b[4];
  assign n1106 = b[3];
  assign n1107 = b[2];
  assign n1108 = b[1];

  FA_X1 U333 ( .A(n681), .B(n304), .CI(n700), .CO(n300), .S(n301) );
  FA_X1 U334 ( .A(n305), .B(n682), .CI(n308), .CO(n302), .S(n303) );
  FA_X1 U336 ( .A(n312), .B(n683), .CI(n309), .CO(n306), .S(n307) );
  FA_X1 U337 ( .A(n701), .B(n314), .CI(n720), .CO(n308), .S(n309) );
  FA_X1 U338 ( .A(n313), .B(n320), .CI(n318), .CO(n310), .S(n311) );
  FA_X1 U339 ( .A(n684), .B(n702), .CI(n315), .CO(n312), .S(n313) );
  FA_X1 U341 ( .A(n324), .B(n321), .CI(n319), .CO(n316), .S(n317) );
  FA_X1 U342 ( .A(n328), .B(n721), .CI(n326), .CO(n318), .S(n319) );
  FA_X1 U343 ( .A(n703), .B(n685), .CI(n740), .CO(n320), .S(n321) );
  FA_X1 U344 ( .A(n325), .B(n327), .CI(n332), .CO(n322), .S(n323) );
  FA_X1 U345 ( .A(n336), .B(n329), .CI(n334), .CO(n324), .S(n325) );
  FA_X1 U346 ( .A(n686), .B(n704), .CI(n722), .CO(n326), .S(n327) );
  FA_X1 U348 ( .A(n340), .B(n342), .CI(n333), .CO(n330), .S(n331) );
  FA_X1 U349 ( .A(n335), .B(n344), .CI(n337), .CO(n332), .S(n333) );
  FA_X1 U350 ( .A(n705), .B(n346), .CI(n723), .CO(n334), .S(n335) );
  FA_X1 U351 ( .A(n741), .B(n687), .CI(n760), .CO(n336), .S(n337) );
  FA_X1 U352 ( .A(n350), .B(n343), .CI(n341), .CO(n338), .S(n339) );
  FA_X1 U353 ( .A(n345), .B(n354), .CI(n352), .CO(n340), .S(n341) );
  FA_X1 U354 ( .A(n347), .B(n724), .CI(n356), .CO(n342), .S(n343) );
  FA_X1 U355 ( .A(n742), .B(n706), .CI(n688), .CO(n344), .S(n345) );
  FA_X1 U357 ( .A(n360), .B(n353), .CI(n351), .CO(n348), .S(n349) );
  FA_X1 U358 ( .A(n357), .B(n355), .CI(n362), .CO(n350), .S(n351) );
  FA_X1 U359 ( .A(n366), .B(n743), .CI(n364), .CO(n352), .S(n353) );
  FA_X1 U360 ( .A(n707), .B(n761), .CI(n725), .CO(n354), .S(n355) );
  FA_X1 U361 ( .A(n368), .B(n689), .CI(n780), .CO(n356), .S(n357) );
  FA_X1 U362 ( .A(n372), .B(n363), .CI(n361), .CO(n358), .S(n359) );
  FA_X1 U363 ( .A(n376), .B(n365), .CI(n374), .CO(n360), .S(n361) );
  FA_X1 U364 ( .A(n378), .B(n380), .CI(n367), .CO(n362), .S(n363) );
  FA_X1 U365 ( .A(n690), .B(n708), .CI(n369), .CO(n364), .S(n365) );
  FA_X1 U366 ( .A(n762), .B(n726), .CI(n744), .CO(n366), .S(n367) );
  FA_X1 U368 ( .A(n384), .B(n375), .CI(n373), .CO(n370), .S(n371) );
  FA_X1 U369 ( .A(n377), .B(n388), .CI(n386), .CO(n372), .S(n373) );
  FA_X1 U370 ( .A(n379), .B(n390), .CI(n381), .CO(n374), .S(n375) );
  FA_X1 U371 ( .A(n727), .B(n745), .CI(n392), .CO(n376), .S(n377) );
  FA_X1 U372 ( .A(n709), .B(n781), .CI(n763), .CO(n378), .S(n379) );
  FA_X1 U373 ( .A(n394), .B(n691), .CI(n800), .CO(n380), .S(n381) );
  FA_X1 U374 ( .A(n398), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U375 ( .A(n389), .B(n402), .CI(n400), .CO(n384), .S(n385) );
  FA_X1 U376 ( .A(n391), .B(n404), .CI(n393), .CO(n386), .S(n387) );
  FA_X1 U377 ( .A(n408), .B(n395), .CI(n406), .CO(n388), .S(n389) );
  FA_X1 U378 ( .A(n746), .B(n782), .CI(n764), .CO(n390), .S(n391) );
  FA_X1 U379 ( .A(n692), .B(n728), .CI(n710), .CO(n392), .S(n393) );
  FA_X1 U381 ( .A(n401), .B(n412), .CI(n399), .CO(n396), .S(n397) );
  FA_X1 U382 ( .A(n403), .B(n416), .CI(n414), .CO(n398), .S(n399) );
  FA_X1 U384 ( .A(n420), .B(n422), .CI(n405), .CO(n402), .S(n403) );
  FA_X1 U385 ( .A(n729), .B(n765), .CI(n747), .CO(n404), .S(n405) );
  FA_X1 U386 ( .A(n711), .B(n801), .CI(n783), .CO(n406), .S(n407) );
  FA_X1 U387 ( .A(n1330), .B(n693), .CI(n820), .CO(n408), .S(n409) );
  FA_X1 U391 ( .A(n436), .B(n438), .CI(n421), .CO(n416), .S(n417) );
  FA_X1 U393 ( .A(n694), .B(n766), .CI(n712), .CO(n420), .S(n421) );
  FA_X1 U394 ( .A(n802), .B(n730), .CI(n784), .CO(n422), .S(n423) );
  FA_X1 U396 ( .A(n444), .B(n431), .CI(n429), .CO(n426), .S(n427) );
  FA_X1 U397 ( .A(n433), .B(n448), .CI(n446), .CO(n428), .S(n429) );
  FA_X1 U398 ( .A(n450), .B(n441), .CI(n435), .CO(n430), .S(n431) );
  FA_X1 U399 ( .A(n452), .B(n437), .CI(n439), .CO(n432), .S(n433) );
  FA_X1 U400 ( .A(n456), .B(n767), .CI(n454), .CO(n434), .S(n435) );
  FA_X1 U401 ( .A(n785), .B(n749), .CI(n731), .CO(n436), .S(n437) );
  FA_X1 U402 ( .A(n803), .B(n1270), .CI(n713), .CO(n438), .S(n439) );
  FA_X1 U407 ( .A(n455), .B(n470), .CI(n457), .CO(n448), .S(n449) );
  FA_X1 U408 ( .A(n472), .B(n476), .CI(n474), .CO(n450), .S(n451) );
  FA_X1 U409 ( .A(n768), .B(n786), .CI(n459), .CO(n452), .S(n453) );
  FA_X1 U416 ( .A(n473), .B(n488), .CI(n475), .CO(n466), .S(n467) );
  FA_X1 U417 ( .A(n492), .B(n477), .CI(n490), .CO(n468), .S(n469) );
  FA_X1 U418 ( .A(n805), .B(n823), .CI(n494), .CO(n470), .S(n471) );
  FA_X1 U420 ( .A(n697), .B(n860), .CI(n769), .CO(n474), .S(n475) );
  FA_X1 U423 ( .A(n498), .B(n483), .CI(n481), .CO(n478), .S(n479) );
  FA_X1 U424 ( .A(n500), .B(n487), .CI(n485), .CO(n480), .S(n481) );
  FA_X1 U426 ( .A(n489), .B(n506), .CI(n491), .CO(n484), .S(n485) );
  FA_X1 U427 ( .A(n510), .B(n495), .CI(n508), .CO(n486), .S(n487) );
  FA_X1 U428 ( .A(n770), .B(n842), .CI(n824), .CO(n488), .S(n489) );
  FA_X1 U429 ( .A(n806), .B(n752), .CI(n861), .CO(n490), .S(n491) );
  HA_X1 U431 ( .A(n716), .B(n698), .CO(n494), .S(n495) );
  FA_X1 U436 ( .A(n526), .B(n807), .CI(n524), .CO(n504), .S(n505) );
  FA_X1 U437 ( .A(n825), .B(n771), .CI(n789), .CO(n506), .S(n507) );
  FA_X1 U438 ( .A(n717), .B(n843), .CI(n753), .CO(n508), .S(n509) );
  FA_X1 U439 ( .A(n862), .B(n735), .CI(n699), .CO(n510), .S(n511) );
  FA_X1 U441 ( .A(n532), .B(n521), .CI(n519), .CO(n514), .S(n515) );
  FA_X1 U443 ( .A(n536), .B(n540), .CI(n538), .CO(n518), .S(n519) );
  FA_X1 U444 ( .A(n826), .B(n844), .CI(n527), .CO(n520), .S(n521) );
  FA_X1 U445 ( .A(n754), .B(n772), .CI(n808), .CO(n522), .S(n523) );
  FA_X1 U446 ( .A(n863), .B(n790), .CI(n671), .CO(n524), .S(n525) );
  HA_X1 U447 ( .A(n718), .B(n736), .CO(n526), .S(n527) );
  FA_X1 U450 ( .A(n537), .B(n541), .CI(n539), .CO(n532), .S(n533) );
  FA_X1 U451 ( .A(n552), .B(n554), .CI(n550), .CO(n534), .S(n535) );
  FA_X1 U453 ( .A(n845), .B(n737), .CI(n773), .CO(n538), .S(n539) );
  FA_X1 U457 ( .A(n562), .B(n564), .CI(n551), .CO(n546), .S(n547) );
  FA_X1 U458 ( .A(n555), .B(n846), .CI(n566), .CO(n548), .S(n549) );
  FA_X1 U459 ( .A(n792), .B(n865), .CI(n828), .CO(n550), .S(n551) );
  HA_X1 U461 ( .A(n738), .B(n756), .CO(n554), .S(n555) );
  FA_X1 U462 ( .A(n561), .B(n570), .CI(n559), .CO(n556), .S(n557) );
  FA_X1 U463 ( .A(n563), .B(n565), .CI(n572), .CO(n558), .S(n559) );
  FA_X1 U464 ( .A(n574), .B(n576), .CI(n567), .CO(n560), .S(n561) );
  FA_X1 U465 ( .A(n811), .B(n829), .CI(n578), .CO(n562), .S(n563) );
  FA_X1 U466 ( .A(n757), .B(n847), .CI(n793), .CO(n564), .S(n565) );
  FA_X1 U467 ( .A(n866), .B(n739), .CI(n775), .CO(n566), .S(n567) );
  FA_X1 U468 ( .A(n582), .B(n573), .CI(n571), .CO(n568), .S(n569) );
  FA_X1 U469 ( .A(n577), .B(n575), .CI(n584), .CO(n570), .S(n571) );
  FA_X1 U470 ( .A(n588), .B(n579), .CI(n586), .CO(n572), .S(n573) );
  FA_X1 U471 ( .A(n794), .B(n848), .CI(n830), .CO(n574), .S(n575) );
  FA_X1 U472 ( .A(n867), .B(n812), .CI(n673), .CO(n576), .S(n577) );
  HA_X1 U473 ( .A(n758), .B(n776), .CO(n578), .S(n579) );
  FA_X1 U474 ( .A(n585), .B(n592), .CI(n583), .CO(n580), .S(n581) );
  FA_X1 U475 ( .A(n587), .B(n589), .CI(n594), .CO(n582), .S(n583) );
  FA_X1 U476 ( .A(n598), .B(n831), .CI(n596), .CO(n584), .S(n585) );
  FA_X1 U477 ( .A(n777), .B(n849), .CI(n813), .CO(n586), .S(n587) );
  FA_X1 U478 ( .A(n795), .B(n759), .CI(n868), .CO(n588), .S(n589) );
  FA_X1 U479 ( .A(n602), .B(n595), .CI(n593), .CO(n590), .S(n591) );
  FA_X1 U480 ( .A(n604), .B(n606), .CI(n597), .CO(n592), .S(n593) );
  FA_X1 U481 ( .A(n814), .B(n850), .CI(n599), .CO(n594), .S(n595) );
  FA_X1 U482 ( .A(n869), .B(n832), .CI(n674), .CO(n596), .S(n597) );
  HA_X1 U483 ( .A(n778), .B(n796), .CO(n598), .S(n599) );
  FA_X1 U484 ( .A(n610), .B(n605), .CI(n603), .CO(n600), .S(n601) );
  FA_X1 U485 ( .A(n612), .B(n614), .CI(n607), .CO(n602), .S(n603) );
  FA_X1 U486 ( .A(n797), .B(n851), .CI(n833), .CO(n604), .S(n605) );
  FA_X1 U488 ( .A(n613), .B(n618), .CI(n611), .CO(n608), .S(n609) );
  FA_X1 U489 ( .A(n615), .B(n871), .CI(n620), .CO(n610), .S(n611) );
  FA_X1 U490 ( .A(n852), .B(n834), .CI(n675), .CO(n612), .S(n613) );
  HA_X1 U491 ( .A(n798), .B(n816), .CO(n614), .S(n615) );
  FA_X1 U492 ( .A(n621), .B(n624), .CI(n619), .CO(n616), .S(n617) );
  FA_X1 U493 ( .A(n817), .B(n853), .CI(n626), .CO(n618), .S(n619) );
  FA_X1 U494 ( .A(n835), .B(n799), .CI(n872), .CO(n620), .S(n621) );
  FA_X1 U495 ( .A(n630), .B(n627), .CI(n625), .CO(n622), .S(n623) );
  FA_X1 U496 ( .A(n854), .B(n873), .CI(n676), .CO(n624), .S(n625) );
  HA_X1 U497 ( .A(n818), .B(n836), .CO(n626), .S(n627) );
  FA_X1 U498 ( .A(n634), .B(n837), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U499 ( .A(n874), .B(n819), .CI(n855), .CO(n630), .S(n631) );
  FA_X1 U500 ( .A(n677), .B(n856), .CI(n635), .CO(n632), .S(n633) );
  HA_X1 U501 ( .A(n838), .B(n875), .CO(n634), .S(n635) );
  FA_X1 U502 ( .A(n876), .B(n839), .CI(n857), .CO(n636), .S(n637) );
  HA_X1 U503 ( .A(n858), .B(n877), .CO(n638), .S(n639) );
  CLKBUF_X3 U1025 ( .A(n9), .Z(n1552) );
  CLKBUF_X3 U1026 ( .A(n9), .Z(n1553) );
  CLKBUF_X1 U1027 ( .A(n1593), .Z(n1233) );
  CLKBUF_X1 U1028 ( .A(n1560), .Z(n1266) );
  NOR2_X2 U1029 ( .A1(n443), .A2(n460), .ZN(n161) );
  BUF_X1 U1030 ( .A(n48), .Z(n1521) );
  BUF_X2 U1031 ( .A(n1107), .Z(n1356) );
  BUF_X2 U1032 ( .A(n1094), .Z(n1595) );
  BUF_X2 U1033 ( .A(n52), .Z(n1549) );
  BUF_X1 U1034 ( .A(n13), .Z(n1349) );
  OAI22_X1 U1035 ( .A1(n24), .A2(n1327), .B1(n1015), .B2(n1547), .ZN(n1234) );
  XNOR2_X1 U1036 ( .A(n714), .B(n1235), .ZN(n455) );
  XNOR2_X1 U1037 ( .A(n732), .B(n804), .ZN(n1235) );
  BUF_X2 U1038 ( .A(n1395), .Z(n1351) );
  NOR2_X2 U1039 ( .A1(n371), .A2(n382), .ZN(n135) );
  BUF_X1 U1040 ( .A(n31), .Z(n1545) );
  BUF_X1 U1041 ( .A(n1090), .Z(n1599) );
  BUF_X1 U1042 ( .A(n1103), .Z(n1589) );
  BUF_X2 U1043 ( .A(n31), .Z(n1372) );
  BUF_X2 U1044 ( .A(n1100), .Z(n1592) );
  BUF_X2 U1045 ( .A(n1098), .Z(n1325) );
  OR2_X1 U1046 ( .A1(n1454), .A2(n1455), .ZN(n30) );
  BUF_X1 U1047 ( .A(n1101), .Z(n1591) );
  BUF_X2 U1048 ( .A(n1102), .Z(n1590) );
  BUF_X2 U1049 ( .A(n25), .Z(n1394) );
  BUF_X2 U1050 ( .A(n1103), .Z(n1334) );
  BUF_X2 U1051 ( .A(n22), .Z(n1547) );
  OAI22_X1 U1052 ( .A1(n54), .A2(n916), .B1(n915), .B2(n1549), .ZN(n714) );
  XNOR2_X1 U1053 ( .A(n1402), .B(n1403), .ZN(n419) );
  BUF_X2 U1054 ( .A(n1091), .Z(n1598) );
  BUF_X2 U1055 ( .A(n1092), .Z(n1597) );
  BUF_X2 U1056 ( .A(n1554), .Z(n1338) );
  BUF_X2 U1057 ( .A(n1093), .Z(n1596) );
  BUF_X2 U1058 ( .A(n52), .Z(n1550) );
  BUF_X2 U1059 ( .A(n1), .Z(n1357) );
  NAND2_X1 U1060 ( .A1(n569), .A2(n580), .ZN(n210) );
  INV_X1 U1061 ( .A(n1427), .ZN(n227) );
  OAI22_X1 U1062 ( .A1(n1352), .A2(n936), .B1(n935), .B2(n1365), .ZN(n1236) );
  BUF_X2 U1063 ( .A(n19), .Z(n1345) );
  OR2_X1 U1064 ( .A1(n679), .A2(n879), .ZN(n1237) );
  AND2_X1 U1065 ( .A1(n1237), .A2(n263), .ZN(product[1]) );
  XNOR2_X1 U1066 ( .A(n1333), .B(n1398), .ZN(n1239) );
  INV_X1 U1067 ( .A(n1141), .ZN(n1240) );
  CLKBUF_X3 U1068 ( .A(n49), .Z(n1411) );
  CLKBUF_X1 U1069 ( .A(n464), .Z(n1241) );
  NOR2_X1 U1070 ( .A1(n461), .A2(n478), .ZN(n1242) );
  NOR2_X1 U1071 ( .A1(n461), .A2(n478), .ZN(n166) );
  XNOR2_X1 U1072 ( .A(n1380), .B(n1371), .ZN(n1243) );
  BUF_X2 U1073 ( .A(n31), .Z(n1371) );
  BUF_X2 U1074 ( .A(n13), .Z(n1348) );
  INV_X1 U1075 ( .A(n641), .ZN(n1244) );
  CLKBUF_X3 U1076 ( .A(n58), .Z(n1341) );
  INV_X1 U1077 ( .A(n1354), .ZN(n1245) );
  CLKBUF_X1 U1078 ( .A(n58), .Z(n1551) );
  AOI21_X1 U1079 ( .B1(n221), .B2(n213), .A(n214), .ZN(n1246) );
  XOR2_X1 U1080 ( .A(n516), .B(n505), .Z(n1247) );
  XOR2_X1 U1081 ( .A(n1247), .B(n503), .Z(n499) );
  XOR2_X1 U1082 ( .A(n514), .B(n501), .Z(n1248) );
  XOR2_X1 U1083 ( .A(n1248), .B(n499), .Z(n497) );
  NAND2_X1 U1084 ( .A1(n516), .A2(n505), .ZN(n1249) );
  NAND2_X1 U1085 ( .A1(n516), .A2(n503), .ZN(n1250) );
  NAND2_X1 U1086 ( .A1(n505), .A2(n503), .ZN(n1251) );
  NAND3_X1 U1087 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n498) );
  NAND2_X1 U1088 ( .A1(n514), .A2(n501), .ZN(n1252) );
  NAND2_X1 U1089 ( .A1(n514), .A2(n499), .ZN(n1253) );
  NAND2_X1 U1090 ( .A1(n501), .A2(n499), .ZN(n1254) );
  NAND3_X1 U1091 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n496) );
  BUF_X2 U1092 ( .A(n1096), .Z(n1377) );
  AOI21_X1 U1093 ( .B1(n221), .B2(n213), .A(n214), .ZN(n212) );
  BUF_X2 U1094 ( .A(n12), .Z(n1458) );
  CLKBUF_X1 U1095 ( .A(n451), .Z(n1255) );
  XOR2_X1 U1096 ( .A(n419), .B(n423), .Z(n1256) );
  XOR2_X1 U1097 ( .A(n434), .B(n1256), .Z(n415) );
  NAND2_X1 U1098 ( .A1(n434), .A2(n419), .ZN(n1257) );
  NAND2_X1 U1099 ( .A1(n434), .A2(n423), .ZN(n1258) );
  NAND2_X1 U1100 ( .A1(n419), .A2(n423), .ZN(n1259) );
  NAND3_X1 U1101 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n414) );
  CLKBUF_X1 U1102 ( .A(n870), .Z(n1260) );
  XNOR2_X1 U1103 ( .A(n1391), .B(n535), .ZN(n1261) );
  CLKBUF_X2 U1104 ( .A(n22), .Z(n1546) );
  OR2_X2 U1105 ( .A1(n1404), .A2(n1461), .ZN(n1262) );
  NAND2_X1 U1106 ( .A1(n99), .A2(n302), .ZN(n1263) );
  NAND2_X1 U1107 ( .A1(n1397), .A2(n9), .ZN(n1264) );
  NAND2_X1 U1108 ( .A1(n1397), .A2(n9), .ZN(n1519) );
  CLKBUF_X3 U1109 ( .A(n46), .Z(n1548) );
  CLKBUF_X1 U1110 ( .A(n133), .Z(n1265) );
  BUF_X1 U1111 ( .A(n1560), .Z(n1368) );
  XNOR2_X1 U1112 ( .A(n1580), .B(a[16]), .ZN(n1267) );
  XOR2_X1 U1113 ( .A(n1580), .B(a[14]), .Z(n1268) );
  BUF_X2 U1114 ( .A(n43), .Z(n1580) );
  AOI21_X1 U1115 ( .B1(n1531), .B2(n190), .A(n1561), .ZN(n1269) );
  CLKBUF_X1 U1116 ( .A(n1560), .Z(n1367) );
  OAI22_X1 U1117 ( .A1(n1049), .A2(n1519), .B1(n1048), .B2(n1552), .ZN(n1270)
         );
  BUF_X2 U1118 ( .A(n1555), .Z(n1271) );
  BUF_X1 U1119 ( .A(n12), .Z(n1460) );
  CLKBUF_X1 U1120 ( .A(n530), .Z(n1272) );
  XOR2_X1 U1121 ( .A(n417), .B(n432), .Z(n1273) );
  XOR2_X1 U1122 ( .A(n430), .B(n1273), .Z(n413) );
  NAND2_X1 U1123 ( .A1(n430), .A2(n417), .ZN(n1274) );
  NAND2_X1 U1124 ( .A1(n430), .A2(n432), .ZN(n1275) );
  NAND2_X1 U1125 ( .A1(n417), .A2(n432), .ZN(n1276) );
  NAND3_X1 U1126 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n412) );
  XNOR2_X1 U1127 ( .A(n1277), .B(n1316), .ZN(n545) );
  XNOR2_X1 U1128 ( .A(n560), .B(n553), .ZN(n1277) );
  NAND2_X1 U1129 ( .A1(n732), .A2(n714), .ZN(n1278) );
  NAND2_X1 U1130 ( .A1(n714), .A2(n804), .ZN(n1279) );
  NAND2_X1 U1131 ( .A1(n732), .A2(n804), .ZN(n1280) );
  NAND3_X1 U1132 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n454) );
  CLKBUF_X2 U1133 ( .A(n43), .Z(n1449) );
  INV_X1 U1134 ( .A(n170), .ZN(n1281) );
  BUF_X2 U1135 ( .A(n34), .Z(n1376) );
  CLKBUF_X1 U1136 ( .A(n1466), .Z(n1282) );
  CLKBUF_X1 U1137 ( .A(n37), .Z(n1395) );
  XOR2_X1 U1138 ( .A(n750), .B(n696), .Z(n1283) );
  XOR2_X1 U1139 ( .A(n822), .B(n1283), .Z(n457) );
  NAND2_X1 U1140 ( .A1(n822), .A2(n696), .ZN(n1284) );
  NAND2_X1 U1141 ( .A1(n822), .A2(n750), .ZN(n1285) );
  NAND2_X1 U1142 ( .A1(n750), .A2(n696), .ZN(n1286) );
  NAND3_X1 U1143 ( .A1(n1285), .A2(n1284), .A3(n1286), .ZN(n456) );
  OR2_X2 U1144 ( .A1(n1543), .A2(n1544), .ZN(n1432) );
  XOR2_X1 U1145 ( .A(n468), .B(n453), .Z(n1287) );
  XOR2_X1 U1146 ( .A(n1255), .B(n1287), .Z(n447) );
  NAND2_X1 U1147 ( .A1(n451), .A2(n468), .ZN(n1288) );
  NAND2_X1 U1148 ( .A1(n451), .A2(n453), .ZN(n1289) );
  NAND2_X1 U1149 ( .A1(n468), .A2(n453), .ZN(n1290) );
  NAND3_X1 U1150 ( .A1(n1288), .A2(n1289), .A3(n1290), .ZN(n446) );
  XOR2_X1 U1151 ( .A(n407), .B(n409), .Z(n1291) );
  XOR2_X1 U1152 ( .A(n418), .B(n1291), .Z(n401) );
  NAND2_X1 U1153 ( .A1(n418), .A2(n407), .ZN(n1292) );
  NAND2_X1 U1154 ( .A1(n418), .A2(n409), .ZN(n1293) );
  NAND2_X1 U1155 ( .A1(n407), .A2(n409), .ZN(n1294) );
  NAND3_X1 U1156 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n400) );
  XOR2_X1 U1157 ( .A(n523), .B(n525), .Z(n1295) );
  XOR2_X1 U1158 ( .A(n534), .B(n1295), .Z(n517) );
  NAND2_X1 U1159 ( .A1(n534), .A2(n523), .ZN(n1296) );
  NAND2_X1 U1160 ( .A1(n534), .A2(n525), .ZN(n1297) );
  NAND2_X1 U1161 ( .A1(n523), .A2(n525), .ZN(n1298) );
  NAND3_X1 U1162 ( .A1(n1296), .A2(n1297), .A3(n1298), .ZN(n516) );
  XOR2_X1 U1163 ( .A(n520), .B(n509), .Z(n1299) );
  XOR2_X1 U1164 ( .A(n518), .B(n1299), .Z(n501) );
  NAND2_X1 U1165 ( .A1(n518), .A2(n520), .ZN(n1300) );
  NAND2_X1 U1166 ( .A1(n518), .A2(n509), .ZN(n1301) );
  NAND2_X1 U1167 ( .A1(n520), .A2(n509), .ZN(n1302) );
  NAND3_X1 U1168 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n500) );
  NOR2_X1 U1169 ( .A1(n131), .A2(n128), .ZN(n1303) );
  XOR2_X1 U1170 ( .A(n670), .B(n734), .Z(n1304) );
  XOR2_X1 U1171 ( .A(n788), .B(n1304), .Z(n493) );
  NAND2_X1 U1172 ( .A1(n788), .A2(n670), .ZN(n1305) );
  NAND2_X1 U1173 ( .A1(n788), .A2(n734), .ZN(n1306) );
  NAND2_X1 U1174 ( .A1(n670), .A2(n734), .ZN(n1307) );
  NAND3_X1 U1175 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n492) );
  CLKBUF_X1 U1176 ( .A(n1), .Z(n1308) );
  OAI22_X1 U1177 ( .A1(n1352), .A2(n936), .B1(n935), .B2(n1365), .ZN(n733) );
  XOR2_X1 U1178 ( .A(n547), .B(n558), .Z(n1309) );
  XOR2_X1 U1179 ( .A(n1309), .B(n545), .Z(n543) );
  NAND2_X1 U1180 ( .A1(n560), .A2(n553), .ZN(n1310) );
  NAND2_X1 U1181 ( .A1(n560), .A2(n549), .ZN(n1311) );
  NAND2_X1 U1182 ( .A1(n553), .A2(n549), .ZN(n1312) );
  NAND3_X1 U1183 ( .A1(n1310), .A2(n1311), .A3(n1312), .ZN(n544) );
  NAND2_X1 U1184 ( .A1(n547), .A2(n558), .ZN(n1313) );
  NAND2_X1 U1185 ( .A1(n547), .A2(n545), .ZN(n1314) );
  NAND2_X1 U1186 ( .A1(n558), .A2(n545), .ZN(n1315) );
  NAND3_X1 U1187 ( .A1(n1313), .A2(n1314), .A3(n1315), .ZN(n542) );
  CLKBUF_X1 U1188 ( .A(n549), .Z(n1316) );
  XOR2_X1 U1189 ( .A(n774), .B(n672), .Z(n1317) );
  XOR2_X1 U1190 ( .A(n810), .B(n1317), .Z(n553) );
  NAND2_X1 U1191 ( .A1(n810), .A2(n774), .ZN(n1318) );
  NAND2_X1 U1192 ( .A1(n810), .A2(n672), .ZN(n1319) );
  NAND2_X1 U1193 ( .A1(n774), .A2(n672), .ZN(n1320) );
  NAND3_X1 U1194 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n552) );
  XOR2_X1 U1195 ( .A(n809), .B(n791), .Z(n1321) );
  XOR2_X1 U1196 ( .A(n1321), .B(n827), .Z(n537) );
  NAND2_X1 U1197 ( .A1(n827), .A2(n791), .ZN(n1322) );
  NAND2_X1 U1198 ( .A1(n827), .A2(n1234), .ZN(n1323) );
  NAND2_X1 U1199 ( .A1(n791), .A2(n1234), .ZN(n1324) );
  NAND3_X1 U1200 ( .A1(n1322), .A2(n1323), .A3(n1324), .ZN(n536) );
  CLKBUF_X3 U1201 ( .A(n61), .Z(n1582) );
  CLKBUF_X1 U1202 ( .A(n840), .Z(n1326) );
  XNOR2_X1 U1203 ( .A(n1592), .B(n1345), .ZN(n1327) );
  XNOR2_X1 U1204 ( .A(n1593), .B(n1394), .ZN(n1328) );
  OAI22_X1 U1205 ( .A1(n42), .A2(n955), .B1(n954), .B2(n1559), .ZN(n1329) );
  OAI22_X1 U1206 ( .A1(n42), .A2(n955), .B1(n954), .B2(n1559), .ZN(n1366) );
  OAI22_X1 U1207 ( .A1(n18), .A2(n1028), .B1(n1027), .B2(n1271), .ZN(n1330) );
  XNOR2_X1 U1208 ( .A(n1331), .B(n482), .ZN(n463) );
  XNOR2_X1 U1209 ( .A(n467), .B(n484), .ZN(n1331) );
  INV_X1 U1210 ( .A(n1455), .ZN(n1332) );
  CLKBUF_X3 U1211 ( .A(n1530), .Z(n1382) );
  BUF_X2 U1212 ( .A(n1090), .Z(n1333) );
  OAI22_X1 U1213 ( .A1(n1519), .A2(n1050), .B1(n1049), .B2(n1553), .ZN(n1335)
         );
  NAND2_X1 U1214 ( .A1(n1527), .A2(n34), .ZN(n1336) );
  NAND2_X1 U1215 ( .A1(n1527), .A2(n34), .ZN(n1443) );
  XNOR2_X1 U1216 ( .A(n1337), .B(n1241), .ZN(n445) );
  XNOR2_X1 U1217 ( .A(n449), .B(n466), .ZN(n1337) );
  CLKBUF_X1 U1218 ( .A(n165), .Z(n1339) );
  NOR2_X1 U1219 ( .A1(n581), .A2(n590), .ZN(n1340) );
  INV_X1 U1220 ( .A(n650), .ZN(n1342) );
  NAND3_X1 U1221 ( .A1(n1263), .A2(n1466), .A3(n1468), .ZN(n1343) );
  INV_X1 U1222 ( .A(n1140), .ZN(n1344) );
  CLKBUF_X3 U1223 ( .A(n55), .Z(n1581) );
  CLKBUF_X1 U1224 ( .A(n19), .Z(n1478) );
  INV_X1 U1225 ( .A(n1554), .ZN(n1346) );
  CLKBUF_X2 U1226 ( .A(n25), .Z(n1347) );
  CLKBUF_X2 U1227 ( .A(n1395), .Z(n1350) );
  CLKBUF_X1 U1228 ( .A(n1395), .Z(n1361) );
  NAND2_X1 U1229 ( .A1(n46), .A2(n1268), .ZN(n1352) );
  INV_X1 U1230 ( .A(n1530), .ZN(n1353) );
  INV_X1 U1231 ( .A(n668), .ZN(n1354) );
  INV_X2 U1232 ( .A(n668), .ZN(n4) );
  BUF_X2 U1233 ( .A(n1105), .Z(n1355) );
  CLKBUF_X1 U1234 ( .A(n1107), .Z(n1585) );
  BUF_X2 U1235 ( .A(n7), .Z(n1578) );
  CLKBUF_X1 U1236 ( .A(n1), .Z(n1577) );
  CLKBUF_X1 U1237 ( .A(n1432), .Z(n1358) );
  XNOR2_X1 U1238 ( .A(n1599), .B(n1308), .ZN(n1359) );
  CLKBUF_X1 U1239 ( .A(n1395), .Z(n1360) );
  CLKBUF_X1 U1240 ( .A(n1395), .Z(n1362) );
  CLKBUF_X1 U1241 ( .A(n1571), .Z(n1363) );
  CLKBUF_X1 U1242 ( .A(n1570), .Z(n1364) );
  XNOR2_X2 U1243 ( .A(n1579), .B(a[14]), .ZN(n1365) );
  BUF_X2 U1244 ( .A(n37), .Z(n1579) );
  BUF_X1 U1245 ( .A(n1097), .Z(n1369) );
  BUF_X1 U1246 ( .A(n1097), .Z(n1370) );
  BUF_X1 U1247 ( .A(n1106), .Z(n1373) );
  BUF_X1 U1248 ( .A(n1106), .Z(n1374) );
  BUF_X2 U1249 ( .A(n34), .Z(n1375) );
  CLKBUF_X1 U1250 ( .A(n1598), .Z(n1378) );
  CLKBUF_X1 U1251 ( .A(n1597), .Z(n1379) );
  BUF_X2 U1252 ( .A(n1101), .Z(n1380) );
  XNOR2_X1 U1253 ( .A(n1429), .B(n31), .ZN(n1544) );
  CLKBUF_X1 U1254 ( .A(n194), .Z(n1381) );
  XNOR2_X1 U1255 ( .A(n19), .B(a[8]), .ZN(n1530) );
  CLKBUF_X1 U1256 ( .A(n176), .Z(n1383) );
  AOI21_X1 U1257 ( .B1(n1381), .B2(n175), .A(n1383), .ZN(n1384) );
  NAND2_X1 U1258 ( .A1(n1526), .A2(n1551), .ZN(n1385) );
  NAND2_X1 U1259 ( .A1(n1526), .A2(n1551), .ZN(n1386) );
  NAND2_X1 U1260 ( .A1(n1526), .A2(n1551), .ZN(n60) );
  XOR2_X1 U1261 ( .A(n1545), .B(a[10]), .Z(n1387) );
  BUF_X1 U1262 ( .A(n36), .Z(n1388) );
  BUF_X2 U1263 ( .A(n36), .Z(n1389) );
  NOR2_X1 U1264 ( .A1(n557), .A2(n568), .ZN(n1390) );
  XNOR2_X1 U1265 ( .A(n1391), .B(n535), .ZN(n531) );
  XNOR2_X1 U1266 ( .A(n546), .B(n548), .ZN(n1391) );
  NAND2_X1 U1267 ( .A1(n1116), .A2(n22), .ZN(n1392) );
  NAND2_X1 U1268 ( .A1(n1116), .A2(n22), .ZN(n1393) );
  NAND2_X1 U1269 ( .A1(n1116), .A2(n22), .ZN(n24) );
  CLKBUF_X1 U1270 ( .A(n1263), .Z(n1396) );
  BUF_X2 U1271 ( .A(n48), .Z(n1522) );
  XOR2_X1 U1272 ( .A(n1578), .B(a[2]), .Z(n1397) );
  BUF_X4 U1273 ( .A(n7), .Z(n1398) );
  XNOR2_X1 U1274 ( .A(n1399), .B(n445), .ZN(n443) );
  XNOR2_X1 U1275 ( .A(n462), .B(n447), .ZN(n1399) );
  XNOR2_X1 U1276 ( .A(n515), .B(n1400), .ZN(n513) );
  XNOR2_X1 U1277 ( .A(n530), .B(n517), .ZN(n1400) );
  INV_X1 U1278 ( .A(n139), .ZN(n1401) );
  NAND3_X1 U1279 ( .A1(n1439), .A2(n1438), .A3(n1437), .ZN(n1402) );
  NAND2_X1 U1280 ( .A1(n1387), .A2(n34), .ZN(n36) );
  XNOR2_X1 U1281 ( .A(n425), .B(n748), .ZN(n1403) );
  INV_X1 U1282 ( .A(n1555), .ZN(n1404) );
  INV_X1 U1283 ( .A(n1404), .ZN(n1405) );
  AOI21_X1 U1284 ( .B1(n1490), .B2(n1265), .A(n134), .ZN(n1406) );
  NAND3_X1 U1285 ( .A1(n1571), .A2(n1570), .A3(n1569), .ZN(n1407) );
  NAND3_X1 U1286 ( .A1(n1363), .A2(n1364), .A3(n1569), .ZN(n1408) );
  BUF_X1 U1287 ( .A(n1513), .Z(n1409) );
  BUF_X1 U1288 ( .A(n1513), .Z(n1410) );
  CLKBUF_X1 U1289 ( .A(n54), .Z(n1412) );
  XOR2_X1 U1290 ( .A(n733), .B(n1329), .Z(n1413) );
  XOR2_X1 U1291 ( .A(n1335), .B(n1413), .Z(n473) );
  NAND2_X1 U1292 ( .A1(n1335), .A2(n733), .ZN(n1414) );
  NAND2_X1 U1293 ( .A1(n841), .A2(n1366), .ZN(n1415) );
  NAND2_X1 U1294 ( .A1(n1236), .A2(n1366), .ZN(n1416) );
  NAND3_X1 U1295 ( .A1(n1414), .A2(n1416), .A3(n1415), .ZN(n472) );
  CLKBUF_X1 U1296 ( .A(n1512), .Z(n1417) );
  XNOR2_X1 U1297 ( .A(n413), .B(n1418), .ZN(n411) );
  XNOR2_X1 U1298 ( .A(n428), .B(n415), .ZN(n1418) );
  NAND2_X1 U1299 ( .A1(n449), .A2(n466), .ZN(n1419) );
  NAND2_X1 U1300 ( .A1(n449), .A2(n464), .ZN(n1420) );
  NAND2_X1 U1301 ( .A1(n466), .A2(n464), .ZN(n1421) );
  NAND3_X1 U1302 ( .A1(n1419), .A2(n1420), .A3(n1421), .ZN(n444) );
  NAND2_X1 U1303 ( .A1(n462), .A2(n447), .ZN(n1422) );
  NAND2_X1 U1304 ( .A1(n462), .A2(n445), .ZN(n1423) );
  NAND2_X1 U1305 ( .A1(n447), .A2(n445), .ZN(n1424) );
  NAND3_X1 U1306 ( .A1(n1422), .A2(n1423), .A3(n1424), .ZN(n442) );
  CLKBUF_X1 U1307 ( .A(n159), .Z(n1425) );
  AND3_X1 U1308 ( .A1(n1477), .A2(n1476), .A3(n1475), .ZN(product[39]) );
  AND2_X1 U1309 ( .A1(n601), .A2(n608), .ZN(n1427) );
  NAND2_X1 U1310 ( .A1(n1579), .A2(a[12]), .ZN(n1430) );
  NAND2_X1 U1311 ( .A1(n1428), .A2(n1429), .ZN(n1431) );
  NAND2_X1 U1312 ( .A1(n1430), .A2(n1431), .ZN(n1543) );
  INV_X1 U1313 ( .A(n1579), .ZN(n1428) );
  INV_X1 U1314 ( .A(a[12]), .ZN(n1429) );
  OR2_X1 U1315 ( .A1(n1543), .A2(n1544), .ZN(n1433) );
  OR2_X1 U1316 ( .A1(n1543), .A2(n1544), .ZN(n42) );
  XNOR2_X1 U1317 ( .A(n471), .B(n1434), .ZN(n465) );
  XNOR2_X1 U1318 ( .A(n469), .B(n486), .ZN(n1434) );
  XNOR2_X1 U1319 ( .A(n1435), .B(n463), .ZN(n461) );
  XNOR2_X1 U1320 ( .A(n480), .B(n465), .ZN(n1435) );
  XOR2_X1 U1321 ( .A(n821), .B(n695), .Z(n1436) );
  XOR2_X1 U1322 ( .A(n1436), .B(n1326), .Z(n441) );
  NAND2_X1 U1323 ( .A1(n821), .A2(n695), .ZN(n1437) );
  NAND2_X1 U1324 ( .A1(n840), .A2(n821), .ZN(n1438) );
  NAND2_X1 U1325 ( .A1(n695), .A2(n840), .ZN(n1439) );
  NAND3_X1 U1326 ( .A1(n1438), .A2(n1437), .A3(n1439), .ZN(n440) );
  NAND2_X1 U1327 ( .A1(n425), .A2(n748), .ZN(n1440) );
  NAND2_X1 U1328 ( .A1(n440), .A2(n425), .ZN(n1441) );
  NAND2_X1 U1329 ( .A1(n748), .A2(n440), .ZN(n1442) );
  NAND3_X1 U1330 ( .A1(n1442), .A2(n1441), .A3(n1440), .ZN(n418) );
  CLKBUF_X1 U1331 ( .A(n264), .Z(n1444) );
  NAND3_X1 U1332 ( .A1(n1396), .A2(n1282), .A3(n1468), .ZN(n1445) );
  NAND2_X1 U1333 ( .A1(n471), .A2(n469), .ZN(n1446) );
  NAND2_X1 U1334 ( .A1(n471), .A2(n486), .ZN(n1447) );
  NAND2_X1 U1335 ( .A1(n469), .A2(n486), .ZN(n1448) );
  NAND3_X1 U1336 ( .A1(n1446), .A2(n1447), .A3(n1448), .ZN(n464) );
  CLKBUF_X3 U1337 ( .A(n43), .Z(n1450) );
  NAND2_X1 U1338 ( .A1(n413), .A2(n428), .ZN(n1451) );
  NAND2_X1 U1339 ( .A1(n413), .A2(n415), .ZN(n1452) );
  NAND2_X1 U1340 ( .A1(n428), .A2(n415), .ZN(n1453) );
  NAND3_X1 U1341 ( .A1(n1451), .A2(n1452), .A3(n1453), .ZN(n410) );
  XNOR2_X1 U1342 ( .A(n25), .B(a[8]), .ZN(n1454) );
  XOR2_X1 U1343 ( .A(n19), .B(a[8]), .Z(n1455) );
  OR2_X2 U1344 ( .A1(n1454), .A2(n1353), .ZN(n1456) );
  OR2_X2 U1345 ( .A1(n1454), .A2(n1353), .ZN(n1457) );
  BUF_X2 U1346 ( .A(n12), .Z(n1459) );
  NAND2_X1 U1347 ( .A1(n1524), .A2(n9), .ZN(n12) );
  OR2_X1 U1348 ( .A1(n1462), .A2(n1461), .ZN(n18) );
  XNOR2_X1 U1349 ( .A(n13), .B(a[4]), .ZN(n1461) );
  XOR2_X1 U1350 ( .A(n1578), .B(a[4]), .Z(n1462) );
  OR2_X2 U1351 ( .A1(n1462), .A2(n1461), .ZN(n1463) );
  OR2_X2 U1352 ( .A1(n1346), .A2(n1461), .ZN(n1464) );
  XOR2_X1 U1353 ( .A(n301), .B(n302), .Z(n1465) );
  XOR2_X1 U1354 ( .A(n1408), .B(n1465), .Z(product[36]) );
  NAND2_X1 U1355 ( .A1(n1407), .A2(n301), .ZN(n1466) );
  NAND2_X1 U1356 ( .A1(n99), .A2(n302), .ZN(n1467) );
  NAND2_X1 U1357 ( .A1(n301), .A2(n302), .ZN(n1468) );
  NAND3_X1 U1358 ( .A1(n1466), .A2(n1467), .A3(n1468), .ZN(n98) );
  NAND3_X1 U1359 ( .A1(n1472), .A2(n1473), .A3(n1471), .ZN(n1469) );
  XOR2_X1 U1360 ( .A(n300), .B(n299), .Z(n1470) );
  XOR2_X1 U1361 ( .A(n1470), .B(n1445), .Z(product[37]) );
  NAND2_X1 U1362 ( .A1(n300), .A2(n299), .ZN(n1471) );
  NAND2_X1 U1363 ( .A1(n98), .A2(n300), .ZN(n1472) );
  NAND2_X1 U1364 ( .A1(n1343), .A2(n299), .ZN(n1473) );
  NAND3_X1 U1365 ( .A1(n1473), .A2(n1472), .A3(n1471), .ZN(n97) );
  XOR2_X1 U1366 ( .A(n680), .B(n298), .Z(n1474) );
  XOR2_X1 U1367 ( .A(n1469), .B(n1474), .Z(product[38]) );
  NAND2_X1 U1368 ( .A1(n680), .A2(n298), .ZN(n1475) );
  NAND2_X1 U1369 ( .A1(n97), .A2(n680), .ZN(n1476) );
  NAND2_X1 U1370 ( .A1(n298), .A2(n97), .ZN(n1477) );
  XNOR2_X1 U1371 ( .A(n531), .B(n1479), .ZN(n529) );
  XNOR2_X1 U1372 ( .A(n544), .B(n533), .ZN(n1479) );
  NAND2_X1 U1373 ( .A1(n546), .A2(n548), .ZN(n1480) );
  NAND2_X1 U1374 ( .A1(n546), .A2(n535), .ZN(n1481) );
  NAND2_X1 U1375 ( .A1(n548), .A2(n535), .ZN(n1482) );
  NAND3_X1 U1376 ( .A1(n1480), .A2(n1481), .A3(n1482), .ZN(n530) );
  NAND2_X1 U1377 ( .A1(n544), .A2(n533), .ZN(n1483) );
  NAND2_X1 U1378 ( .A1(n1261), .A2(n544), .ZN(n1484) );
  NAND2_X1 U1379 ( .A1(n1261), .A2(n533), .ZN(n1485) );
  NAND3_X1 U1380 ( .A1(n1483), .A2(n1484), .A3(n1485), .ZN(n528) );
  NAND2_X1 U1381 ( .A1(n515), .A2(n1272), .ZN(n1486) );
  NAND2_X1 U1382 ( .A1(n515), .A2(n517), .ZN(n1487) );
  NAND2_X1 U1383 ( .A1(n1272), .A2(n517), .ZN(n1488) );
  NAND3_X1 U1384 ( .A1(n1486), .A2(n1487), .A3(n1488), .ZN(n512) );
  XNOR2_X1 U1385 ( .A(n1489), .B(n755), .ZN(n541) );
  XNOR2_X1 U1386 ( .A(n864), .B(n719), .ZN(n1489) );
  CLKBUF_X1 U1387 ( .A(n146), .Z(n1490) );
  CLKBUF_X1 U1388 ( .A(n1385), .Z(n1491) );
  XOR2_X1 U1389 ( .A(n511), .B(n522), .Z(n1492) );
  XOR2_X1 U1390 ( .A(n1492), .B(n507), .Z(n503) );
  NAND2_X1 U1391 ( .A1(n511), .A2(n522), .ZN(n1493) );
  NAND2_X1 U1392 ( .A1(n511), .A2(n507), .ZN(n1494) );
  NAND2_X1 U1393 ( .A1(n522), .A2(n507), .ZN(n1495) );
  NAND3_X1 U1394 ( .A1(n1493), .A2(n1494), .A3(n1495), .ZN(n502) );
  XOR2_X1 U1395 ( .A(n504), .B(n493), .Z(n1496) );
  XOR2_X1 U1396 ( .A(n1496), .B(n502), .Z(n483) );
  NAND2_X1 U1397 ( .A1(n504), .A2(n493), .ZN(n1497) );
  NAND2_X1 U1398 ( .A1(n504), .A2(n502), .ZN(n1498) );
  NAND2_X1 U1399 ( .A1(n493), .A2(n502), .ZN(n1499) );
  NAND3_X1 U1400 ( .A1(n1497), .A2(n1498), .A3(n1499), .ZN(n482) );
  NAND2_X1 U1401 ( .A1(n467), .A2(n484), .ZN(n1500) );
  NAND2_X1 U1402 ( .A1(n467), .A2(n482), .ZN(n1501) );
  NAND2_X1 U1403 ( .A1(n484), .A2(n482), .ZN(n1502) );
  NAND3_X1 U1404 ( .A1(n1500), .A2(n1501), .A3(n1502), .ZN(n462) );
  NAND2_X1 U1405 ( .A1(n480), .A2(n465), .ZN(n1503) );
  NAND2_X1 U1406 ( .A1(n480), .A2(n463), .ZN(n1504) );
  NAND2_X1 U1407 ( .A1(n465), .A2(n463), .ZN(n1505) );
  NAND3_X1 U1408 ( .A1(n1503), .A2(n1504), .A3(n1505), .ZN(n460) );
  CLKBUF_X1 U1409 ( .A(n1568), .Z(n1507) );
  CLKBUF_X1 U1410 ( .A(n127), .Z(n1506) );
  CLKBUF_X1 U1411 ( .A(n106), .Z(n1508) );
  CLKBUF_X1 U1412 ( .A(n122), .Z(n1509) );
  CLKBUF_X1 U1413 ( .A(n1389), .Z(n1510) );
  AOI21_X1 U1414 ( .B1(n122), .B2(n1535), .A(n119), .ZN(n1511) );
  NOR2_X1 U1415 ( .A1(n427), .A2(n442), .ZN(n1512) );
  NAND2_X1 U1416 ( .A1(n1119), .A2(n4), .ZN(n1513) );
  NAND2_X1 U1417 ( .A1(n1119), .A2(n4), .ZN(n1514) );
  NOR2_X1 U1418 ( .A1(n497), .A2(n512), .ZN(n1515) );
  CLKBUF_X1 U1419 ( .A(n114), .Z(n1516) );
  AOI21_X1 U1420 ( .B1(n114), .B2(n1536), .A(n111), .ZN(n1517) );
  NOR2_X1 U1421 ( .A1(n410), .A2(n397), .ZN(n1518) );
  CLKBUF_X1 U1422 ( .A(n153), .Z(n1520) );
  NAND2_X1 U1423 ( .A1(n1525), .A2(n46), .ZN(n48) );
  CLKBUF_X3 U1424 ( .A(n1104), .Z(n1588) );
  XOR2_X1 U1425 ( .A(n179), .B(n1523), .Z(product[18]) );
  AND2_X1 U1426 ( .A1(n280), .A2(n178), .ZN(n1523) );
  NOR2_X1 U1427 ( .A1(n497), .A2(n512), .ZN(n177) );
  NOR2_X1 U1428 ( .A1(n359), .A2(n370), .ZN(n128) );
  NOR2_X1 U1429 ( .A1(n581), .A2(n590), .ZN(n215) );
  NOR2_X1 U1430 ( .A1(n591), .A2(n600), .ZN(n218) );
  XOR2_X1 U1431 ( .A(n1565), .B(n1444), .Z(product[34]) );
  BUF_X2 U1432 ( .A(n1095), .Z(n1594) );
  CLKBUF_X3 U1433 ( .A(n1099), .Z(n1593) );
  BUF_X2 U1434 ( .A(n1105), .Z(n1587) );
  BUF_X2 U1435 ( .A(n1108), .Z(n1584) );
  XOR2_X1 U1436 ( .A(n1578), .B(a[2]), .Z(n1524) );
  XOR2_X1 U1437 ( .A(n1580), .B(a[14]), .Z(n1525) );
  XOR2_X1 U1438 ( .A(n55), .B(a[18]), .Z(n1526) );
  XOR2_X1 U1439 ( .A(n1545), .B(a[10]), .Z(n1527) );
  NAND2_X2 U1440 ( .A1(n1528), .A2(n1267), .ZN(n54) );
  XOR2_X1 U1441 ( .A(n49), .B(a[16]), .Z(n1528) );
  AOI21_X1 U1442 ( .B1(n153), .B2(n126), .A(n127), .ZN(n1529) );
  OAI21_X1 U1443 ( .B1(n152), .B2(n143), .A(n144), .ZN(n142) );
  INV_X1 U1444 ( .A(n1520), .ZN(n152) );
  NAND2_X1 U1445 ( .A1(n145), .A2(n133), .ZN(n131) );
  XOR2_X1 U1446 ( .A(n201), .B(n81), .Z(product[15]) );
  NOR2_X1 U1447 ( .A1(n131), .A2(n128), .ZN(n126) );
  INV_X1 U1448 ( .A(n200), .ZN(n198) );
  XOR2_X1 U1449 ( .A(n137), .B(n70), .Z(product[26]) );
  NAND2_X1 U1450 ( .A1(n272), .A2(n136), .ZN(n70) );
  AOI21_X1 U1451 ( .B1(n142), .B2(n273), .A(n139), .ZN(n137) );
  INV_X1 U1452 ( .A(n135), .ZN(n272) );
  INV_X1 U1453 ( .A(n140), .ZN(n273) );
  INV_X1 U1454 ( .A(n171), .ZN(n279) );
  XOR2_X1 U1455 ( .A(n168), .B(n76), .Z(product[20]) );
  NAND2_X1 U1456 ( .A1(n278), .A2(n167), .ZN(n76) );
  AOI21_X1 U1457 ( .B1(n173), .B2(n279), .A(n170), .ZN(n168) );
  XOR2_X1 U1458 ( .A(n206), .B(n82), .Z(product[14]) );
  NAND2_X1 U1459 ( .A1(n284), .A2(n205), .ZN(n82) );
  AOI21_X1 U1460 ( .B1(n211), .B2(n285), .A(n208), .ZN(n206) );
  XOR2_X1 U1461 ( .A(n152), .B(n73), .Z(product[23]) );
  NAND2_X1 U1462 ( .A1(n275), .A2(n151), .ZN(n73) );
  XOR2_X1 U1463 ( .A(n163), .B(n75), .Z(product[21]) );
  NAND2_X1 U1464 ( .A1(n277), .A2(n162), .ZN(n75) );
  XOR2_X1 U1465 ( .A(n193), .B(n80), .Z(product[16]) );
  NAND2_X1 U1466 ( .A1(n282), .A2(n188), .ZN(n80) );
  XNOR2_X1 U1467 ( .A(n160), .B(n74), .ZN(product[22]) );
  NAND2_X1 U1468 ( .A1(n276), .A2(n1425), .ZN(n74) );
  XNOR2_X1 U1469 ( .A(n173), .B(n77), .ZN(product[19]) );
  NAND2_X1 U1470 ( .A1(n279), .A2(n1281), .ZN(n77) );
  XNOR2_X1 U1471 ( .A(n186), .B(n79), .ZN(product[17]) );
  NAND2_X1 U1472 ( .A1(n1531), .A2(n185), .ZN(n79) );
  INV_X1 U1473 ( .A(n1561), .ZN(n185) );
  XNOR2_X1 U1474 ( .A(n130), .B(n69), .ZN(product[27]) );
  NAND2_X1 U1475 ( .A1(n271), .A2(n129), .ZN(n69) );
  INV_X1 U1476 ( .A(n128), .ZN(n271) );
  INV_X1 U1477 ( .A(n1515), .ZN(n280) );
  XNOR2_X1 U1478 ( .A(n149), .B(n72), .ZN(product[24]) );
  NAND2_X1 U1479 ( .A1(n274), .A2(n148), .ZN(n72) );
  INV_X1 U1480 ( .A(n1518), .ZN(n274) );
  XNOR2_X1 U1481 ( .A(n142), .B(n71), .ZN(product[25]) );
  NAND2_X1 U1482 ( .A1(n273), .A2(n1401), .ZN(n71) );
  INV_X1 U1483 ( .A(n172), .ZN(n170) );
  NAND2_X1 U1484 ( .A1(n1531), .A2(n282), .ZN(n180) );
  INV_X1 U1485 ( .A(n141), .ZN(n139) );
  OR2_X2 U1486 ( .A1(n528), .A2(n513), .ZN(n1531) );
  INV_X1 U1487 ( .A(n113), .ZN(n111) );
  INV_X1 U1488 ( .A(n238), .ZN(n236) );
  NAND2_X1 U1489 ( .A1(n1533), .A2(n1534), .ZN(n222) );
  AOI21_X1 U1490 ( .B1(n1533), .B2(n230), .A(n1427), .ZN(n223) );
  NOR2_X1 U1491 ( .A1(n397), .A2(n410), .ZN(n147) );
  AOI21_X1 U1492 ( .B1(n1509), .B2(n1535), .A(n119), .ZN(n117) );
  INV_X1 U1493 ( .A(n121), .ZN(n119) );
  NOR2_X1 U1494 ( .A1(n557), .A2(n568), .ZN(n204) );
  NOR2_X1 U1495 ( .A1(n427), .A2(n442), .ZN(n158) );
  NOR2_X1 U1496 ( .A1(n411), .A2(n426), .ZN(n150) );
  NAND2_X1 U1497 ( .A1(n268), .A2(n116), .ZN(n66) );
  INV_X1 U1498 ( .A(n115), .ZN(n268) );
  NAND2_X1 U1499 ( .A1(n266), .A2(n108), .ZN(n64) );
  INV_X1 U1500 ( .A(n107), .ZN(n266) );
  NAND2_X1 U1501 ( .A1(n270), .A2(n124), .ZN(n68) );
  INV_X1 U1502 ( .A(n123), .ZN(n270) );
  INV_X1 U1503 ( .A(n232), .ZN(n230) );
  INV_X1 U1504 ( .A(n209), .ZN(n285) );
  NAND2_X1 U1505 ( .A1(n1535), .A2(n121), .ZN(n67) );
  NAND2_X1 U1506 ( .A1(n1537), .A2(n105), .ZN(n63) );
  NAND2_X1 U1507 ( .A1(n1536), .A2(n113), .ZN(n65) );
  NAND2_X1 U1508 ( .A1(n1538), .A2(n238), .ZN(n88) );
  XOR2_X1 U1509 ( .A(n228), .B(n86), .Z(product[10]) );
  NAND2_X1 U1510 ( .A1(n1533), .A2(n227), .ZN(n86) );
  AOI21_X1 U1511 ( .B1(n233), .B2(n1534), .A(n230), .ZN(n228) );
  XOR2_X1 U1512 ( .A(n220), .B(n85), .Z(product[11]) );
  NAND2_X1 U1513 ( .A1(n287), .A2(n219), .ZN(n85) );
  INV_X1 U1514 ( .A(n218), .ZN(n287) );
  NOR2_X1 U1515 ( .A1(n479), .A2(n496), .ZN(n171) );
  NAND2_X1 U1516 ( .A1(n371), .A2(n382), .ZN(n136) );
  NAND2_X1 U1517 ( .A1(n479), .A2(n496), .ZN(n172) );
  INV_X1 U1518 ( .A(n105), .ZN(n103) );
  XNOR2_X1 U1519 ( .A(n211), .B(n83), .ZN(product[13]) );
  NAND2_X1 U1520 ( .A1(n285), .A2(n210), .ZN(n83) );
  XNOR2_X1 U1521 ( .A(n233), .B(n87), .ZN(product[9]) );
  NAND2_X1 U1522 ( .A1(n1534), .A2(n232), .ZN(n87) );
  XNOR2_X1 U1523 ( .A(n217), .B(n84), .ZN(product[12]) );
  NAND2_X1 U1524 ( .A1(n286), .A2(n216), .ZN(n84) );
  OAI21_X1 U1525 ( .B1(n220), .B2(n218), .A(n219), .ZN(n217) );
  INV_X1 U1526 ( .A(n1340), .ZN(n286) );
  NAND2_X1 U1527 ( .A1(n383), .A2(n396), .ZN(n141) );
  NAND2_X1 U1528 ( .A1(n443), .A2(n460), .ZN(n162) );
  NAND2_X1 U1529 ( .A1(n497), .A2(n512), .ZN(n178) );
  NAND2_X1 U1530 ( .A1(n359), .A2(n370), .ZN(n129) );
  NOR2_X1 U1531 ( .A1(n1340), .A2(n218), .ZN(n213) );
  OAI21_X1 U1532 ( .B1(n215), .B2(n219), .A(n216), .ZN(n214) );
  NAND2_X1 U1533 ( .A1(n529), .A2(n542), .ZN(n188) );
  INV_X1 U1534 ( .A(n210), .ZN(n208) );
  OR2_X1 U1535 ( .A1(n543), .A2(n556), .ZN(n1532) );
  AOI21_X1 U1536 ( .B1(n1542), .B2(n255), .A(n252), .ZN(n250) );
  INV_X1 U1537 ( .A(n254), .ZN(n252) );
  OR2_X1 U1538 ( .A1(n601), .A2(n608), .ZN(n1533) );
  OAI21_X1 U1539 ( .B1(n248), .B2(n250), .A(n249), .ZN(n247) );
  NAND2_X1 U1540 ( .A1(n291), .A2(n241), .ZN(n89) );
  INV_X1 U1541 ( .A(n240), .ZN(n291) );
  AOI21_X1 U1542 ( .B1(n1541), .B2(n247), .A(n244), .ZN(n242) );
  INV_X1 U1543 ( .A(n246), .ZN(n244) );
  NAND2_X1 U1544 ( .A1(n591), .A2(n600), .ZN(n219) );
  NAND2_X1 U1545 ( .A1(n1542), .A2(n254), .ZN(n92) );
  NOR2_X1 U1546 ( .A1(n569), .A2(n580), .ZN(n209) );
  NOR2_X1 U1547 ( .A1(n349), .A2(n358), .ZN(n123) );
  NOR2_X1 U1548 ( .A1(n331), .A2(n338), .ZN(n115) );
  NOR2_X1 U1549 ( .A1(n317), .A2(n322), .ZN(n107) );
  NAND2_X1 U1550 ( .A1(n581), .A2(n590), .ZN(n216) );
  OR2_X1 U1551 ( .A1(n609), .A2(n616), .ZN(n1534) );
  OR2_X1 U1552 ( .A1(n339), .A2(n348), .ZN(n1535) );
  NAND2_X1 U1553 ( .A1(n323), .A2(n330), .ZN(n113) );
  NAND2_X1 U1554 ( .A1(n609), .A2(n616), .ZN(n232) );
  NAND2_X1 U1555 ( .A1(n311), .A2(n316), .ZN(n105) );
  NAND2_X1 U1556 ( .A1(n617), .A2(n622), .ZN(n238) );
  NAND2_X1 U1557 ( .A1(n339), .A2(n348), .ZN(n121) );
  NAND2_X1 U1558 ( .A1(n349), .A2(n358), .ZN(n124) );
  NAND2_X1 U1559 ( .A1(n331), .A2(n338), .ZN(n116) );
  NAND2_X1 U1560 ( .A1(n317), .A2(n322), .ZN(n108) );
  OR2_X1 U1561 ( .A1(n323), .A2(n330), .ZN(n1536) );
  OR2_X1 U1562 ( .A1(n311), .A2(n316), .ZN(n1537) );
  OR2_X1 U1563 ( .A1(n617), .A2(n622), .ZN(n1538) );
  INV_X1 U1564 ( .A(n259), .ZN(n258) );
  OAI21_X1 U1565 ( .B1(n260), .B2(n263), .A(n261), .ZN(n259) );
  XOR2_X1 U1566 ( .A(n94), .B(n263), .Z(product[2]) );
  NAND2_X1 U1567 ( .A1(n296), .A2(n261), .ZN(n94) );
  INV_X1 U1568 ( .A(n260), .ZN(n296) );
  XOR2_X1 U1569 ( .A(n91), .B(n250), .Z(product[5]) );
  NAND2_X1 U1570 ( .A1(n293), .A2(n249), .ZN(n91) );
  INV_X1 U1571 ( .A(n248), .ZN(n293) );
  XNOR2_X1 U1572 ( .A(n90), .B(n247), .ZN(product[6]) );
  NAND2_X1 U1573 ( .A1(n1541), .A2(n246), .ZN(n90) );
  XOR2_X1 U1574 ( .A(n93), .B(n258), .Z(product[3]) );
  INV_X1 U1575 ( .A(n256), .ZN(n295) );
  XNOR2_X1 U1576 ( .A(n1333), .B(n1371), .ZN(n964) );
  XNOR2_X1 U1577 ( .A(n1355), .B(n1371), .ZN(n979) );
  XNOR2_X1 U1578 ( .A(n1588), .B(n1371), .ZN(n978) );
  XNOR2_X1 U1579 ( .A(n1369), .B(n1372), .ZN(n971) );
  XNOR2_X1 U1580 ( .A(n1373), .B(n1371), .ZN(n980) );
  XNOR2_X1 U1581 ( .A(n1593), .B(n1372), .ZN(n973) );
  XNOR2_X1 U1582 ( .A(n1380), .B(n1371), .ZN(n975) );
  XNOR2_X1 U1583 ( .A(n1377), .B(n1372), .ZN(n970) );
  XNOR2_X1 U1584 ( .A(n1325), .B(n1372), .ZN(n972) );
  XNOR2_X1 U1585 ( .A(n1584), .B(n1371), .ZN(n982) );
  XNOR2_X1 U1586 ( .A(n1597), .B(n1371), .ZN(n966) );
  NOR2_X1 U1587 ( .A1(n633), .A2(n636), .ZN(n248) );
  NOR2_X1 U1588 ( .A1(n878), .A2(n859), .ZN(n260) );
  XNOR2_X1 U1589 ( .A(n1539), .B(n1564), .ZN(product[35]) );
  XNOR2_X1 U1590 ( .A(n303), .B(n306), .ZN(n1539) );
  NAND2_X1 U1591 ( .A1(n679), .A2(n879), .ZN(n263) );
  XNOR2_X1 U1592 ( .A(n1592), .B(n1372), .ZN(n974) );
  XNOR2_X1 U1593 ( .A(n1334), .B(n1371), .ZN(n977) );
  XNOR2_X1 U1594 ( .A(n1590), .B(n1371), .ZN(n976) );
  XNOR2_X1 U1595 ( .A(n1356), .B(n1371), .ZN(n981) );
  XNOR2_X1 U1596 ( .A(n1594), .B(n1371), .ZN(n969) );
  XNOR2_X1 U1597 ( .A(n1598), .B(n1372), .ZN(n965) );
  XNOR2_X1 U1598 ( .A(n1596), .B(n1372), .ZN(n967) );
  XNOR2_X1 U1599 ( .A(n1595), .B(n1372), .ZN(n968) );
  NAND2_X1 U1600 ( .A1(n878), .A2(n859), .ZN(n261) );
  INV_X1 U1601 ( .A(n394), .ZN(n395) );
  INV_X1 U1602 ( .A(n328), .ZN(n329) );
  XNOR2_X1 U1603 ( .A(n815), .B(n1540), .ZN(n607) );
  XNOR2_X1 U1604 ( .A(n870), .B(n779), .ZN(n1540) );
  NOR2_X1 U1605 ( .A1(n623), .A2(n628), .ZN(n240) );
  NOR2_X1 U1606 ( .A1(n639), .A2(n678), .ZN(n256) );
  NAND2_X1 U1607 ( .A1(n633), .A2(n636), .ZN(n249) );
  INV_X1 U1608 ( .A(n1372), .ZN(n1144) );
  INV_X1 U1609 ( .A(n298), .ZN(n299) );
  OR2_X1 U1610 ( .A1(n629), .A2(n632), .ZN(n1541) );
  NAND2_X1 U1611 ( .A1(n629), .A2(n632), .ZN(n246) );
  OR2_X1 U1612 ( .A1(n637), .A2(n638), .ZN(n1542) );
  NAND2_X1 U1613 ( .A1(n623), .A2(n628), .ZN(n241) );
  OAI22_X1 U1614 ( .A1(n1410), .A2(n1086), .B1(n1085), .B2(n1354), .ZN(n877)
         );
  OAI22_X1 U1615 ( .A1(n1514), .A2(n1088), .B1(n1087), .B2(n1354), .ZN(n879)
         );
  OAI22_X1 U1616 ( .A1(n1409), .A2(n1149), .B1(n1089), .B2(n4), .ZN(n679) );
  OR2_X1 U1617 ( .A1(n1583), .A2(n1149), .ZN(n1089) );
  OAI22_X1 U1618 ( .A1(n1514), .A2(n1087), .B1(n1086), .B2(n1354), .ZN(n878)
         );
  OAI22_X1 U1619 ( .A1(n1514), .A2(n1074), .B1(n1073), .B2(n4), .ZN(n865) );
  XNOR2_X1 U1620 ( .A(n1582), .B(n1372), .ZN(n983) );
  OAI22_X1 U1621 ( .A1(n1514), .A2(n1082), .B1(n1081), .B2(n1354), .ZN(n873)
         );
  OAI22_X1 U1622 ( .A1(n1513), .A2(n1359), .B1(n1069), .B2(n4), .ZN(n667) );
  OR2_X1 U1623 ( .A1(n1583), .A2(n1147), .ZN(n1047) );
  XNOR2_X1 U1624 ( .A(n1582), .B(n1450), .ZN(n941) );
  XNOR2_X1 U1625 ( .A(n1582), .B(n1411), .ZN(n920) );
  OAI22_X1 U1626 ( .A1(n1410), .A2(n1084), .B1(n1083), .B2(n1354), .ZN(n875)
         );
  INV_X1 U1627 ( .A(n1544), .ZN(n1559) );
  XNOR2_X1 U1628 ( .A(n1333), .B(n1450), .ZN(n922) );
  XNOR2_X1 U1629 ( .A(n1333), .B(n1240), .ZN(n901) );
  XNOR2_X1 U1630 ( .A(n1333), .B(n1478), .ZN(n1006) );
  INV_X1 U1631 ( .A(n1382), .ZN(n656) );
  BUF_X1 U1632 ( .A(n1106), .Z(n1586) );
  XNOR2_X1 U1633 ( .A(n1325), .B(n1449), .ZN(n930) );
  XNOR2_X1 U1634 ( .A(n1374), .B(n1450), .ZN(n938) );
  XNOR2_X1 U1635 ( .A(n1585), .B(n1450), .ZN(n939) );
  XNOR2_X1 U1636 ( .A(n1595), .B(n1450), .ZN(n926) );
  XNOR2_X1 U1637 ( .A(n1584), .B(n1449), .ZN(n940) );
  XNOR2_X1 U1638 ( .A(n1589), .B(n1450), .ZN(n935) );
  XNOR2_X1 U1639 ( .A(n1594), .B(n1450), .ZN(n927) );
  XNOR2_X1 U1640 ( .A(n1593), .B(n1449), .ZN(n931) );
  XNOR2_X1 U1641 ( .A(n1587), .B(n1449), .ZN(n937) );
  XNOR2_X1 U1642 ( .A(n1369), .B(n1450), .ZN(n929) );
  XNOR2_X1 U1643 ( .A(n1588), .B(n1449), .ZN(n936) );
  XNOR2_X1 U1644 ( .A(n1596), .B(n1449), .ZN(n925) );
  XNOR2_X1 U1645 ( .A(n1592), .B(n1450), .ZN(n932) );
  XNOR2_X1 U1646 ( .A(n1590), .B(n1450), .ZN(n934) );
  XNOR2_X1 U1647 ( .A(n1377), .B(n1449), .ZN(n928) );
  XNOR2_X1 U1648 ( .A(n1380), .B(n1449), .ZN(n933) );
  XNOR2_X1 U1649 ( .A(n1379), .B(n1449), .ZN(n924) );
  XNOR2_X1 U1650 ( .A(n1378), .B(n1449), .ZN(n923) );
  INV_X1 U1651 ( .A(n304), .ZN(n305) );
  XNOR2_X1 U1652 ( .A(n1374), .B(n1411), .ZN(n917) );
  XNOR2_X1 U1653 ( .A(n1355), .B(n1411), .ZN(n916) );
  XNOR2_X1 U1654 ( .A(n1356), .B(n1411), .ZN(n918) );
  XNOR2_X1 U1655 ( .A(n1584), .B(n1411), .ZN(n919) );
  XNOR2_X1 U1656 ( .A(n1588), .B(n1411), .ZN(n915) );
  XNOR2_X1 U1657 ( .A(n1334), .B(n1411), .ZN(n914) );
  XNOR2_X1 U1658 ( .A(n1594), .B(n1240), .ZN(n906) );
  XNOR2_X1 U1659 ( .A(n1233), .B(n1411), .ZN(n910) );
  XNOR2_X1 U1660 ( .A(n1377), .B(n1240), .ZN(n907) );
  XNOR2_X1 U1661 ( .A(n1380), .B(n1411), .ZN(n912) );
  XNOR2_X1 U1662 ( .A(n1370), .B(n1411), .ZN(n908) );
  XNOR2_X1 U1663 ( .A(n1592), .B(n1411), .ZN(n911) );
  XNOR2_X1 U1664 ( .A(n1590), .B(n1411), .ZN(n913) );
  XNOR2_X1 U1665 ( .A(n1325), .B(n1411), .ZN(n909) );
  XNOR2_X1 U1666 ( .A(n1595), .B(n1240), .ZN(n905) );
  XNOR2_X1 U1667 ( .A(n1596), .B(n1240), .ZN(n904) );
  XNOR2_X1 U1668 ( .A(n1379), .B(n1240), .ZN(n903) );
  XNOR2_X1 U1669 ( .A(n1378), .B(n1240), .ZN(n902) );
  XNOR2_X1 U1670 ( .A(n1369), .B(n1345), .ZN(n1013) );
  XNOR2_X1 U1671 ( .A(n1325), .B(n1345), .ZN(n1014) );
  XNOR2_X1 U1672 ( .A(n1377), .B(n1478), .ZN(n1012) );
  XNOR2_X1 U1673 ( .A(n1594), .B(n1345), .ZN(n1011) );
  XNOR2_X1 U1674 ( .A(n1591), .B(n1478), .ZN(n1017) );
  XNOR2_X1 U1675 ( .A(n1598), .B(n1345), .ZN(n1007) );
  XNOR2_X1 U1676 ( .A(n1593), .B(n1478), .ZN(n1015) );
  XNOR2_X1 U1677 ( .A(n1595), .B(n1345), .ZN(n1010) );
  XNOR2_X1 U1678 ( .A(n1590), .B(n1345), .ZN(n1018) );
  XNOR2_X1 U1679 ( .A(n1592), .B(n1478), .ZN(n1016) );
  XNOR2_X1 U1680 ( .A(n1334), .B(n1345), .ZN(n1019) );
  XNOR2_X1 U1681 ( .A(n1596), .B(n1345), .ZN(n1009) );
  XNOR2_X1 U1682 ( .A(n1588), .B(n1478), .ZN(n1020) );
  XNOR2_X1 U1683 ( .A(n1355), .B(n1345), .ZN(n1021) );
  XNOR2_X1 U1684 ( .A(n1373), .B(n1345), .ZN(n1022) );
  XNOR2_X1 U1685 ( .A(n1356), .B(n1345), .ZN(n1023) );
  XNOR2_X1 U1686 ( .A(n1584), .B(n1345), .ZN(n1024) );
  XNOR2_X1 U1687 ( .A(n1597), .B(n1345), .ZN(n1008) );
  AND2_X1 U1688 ( .A1(n1583), .A2(n665), .ZN(n859) );
  INV_X1 U1689 ( .A(n655), .ZN(n780) );
  INV_X1 U1690 ( .A(n314), .ZN(n315) );
  AND2_X1 U1691 ( .A1(n1583), .A2(n641), .ZN(n699) );
  OAI22_X1 U1692 ( .A1(n1513), .A2(n1071), .B1(n1070), .B2(n4), .ZN(n862) );
  OAI22_X1 U1693 ( .A1(n1514), .A2(n1072), .B1(n1071), .B2(n4), .ZN(n863) );
  INV_X1 U1694 ( .A(n649), .ZN(n740) );
  INV_X1 U1695 ( .A(n643), .ZN(n700) );
  INV_X1 U1696 ( .A(n346), .ZN(n347) );
  AND2_X1 U1697 ( .A1(n1583), .A2(n650), .ZN(n759) );
  OAI22_X1 U1698 ( .A1(n1514), .A2(n1077), .B1(n1076), .B2(n4), .ZN(n868) );
  AND2_X1 U1699 ( .A1(n1583), .A2(n1346), .ZN(n839) );
  OAI22_X1 U1700 ( .A1(n1409), .A2(n1085), .B1(n1084), .B2(n4), .ZN(n876) );
  INV_X1 U1701 ( .A(n667), .ZN(n860) );
  INV_X1 U1702 ( .A(n652), .ZN(n760) );
  INV_X1 U1703 ( .A(n646), .ZN(n720) );
  INV_X1 U1704 ( .A(n424), .ZN(n425) );
  OAI22_X1 U1705 ( .A1(n1409), .A2(n1080), .B1(n1079), .B2(n1354), .ZN(n871)
         );
  AND2_X1 U1706 ( .A1(n1583), .A2(n647), .ZN(n739) );
  OAI22_X1 U1707 ( .A1(n1514), .A2(n1075), .B1(n1074), .B2(n4), .ZN(n866) );
  OAI22_X1 U1708 ( .A1(n1514), .A2(n1078), .B1(n1077), .B2(n1354), .ZN(n869)
         );
  AND2_X1 U1709 ( .A1(n1583), .A2(n659), .ZN(n819) );
  OAI22_X1 U1710 ( .A1(n1410), .A2(n1083), .B1(n1082), .B2(n4), .ZN(n874) );
  OAI22_X1 U1711 ( .A1(n1514), .A2(n1076), .B1(n1075), .B2(n4), .ZN(n867) );
  INV_X1 U1712 ( .A(n458), .ZN(n459) );
  INV_X1 U1713 ( .A(n1450), .ZN(n1142) );
  OAI22_X1 U1714 ( .A1(n1409), .A2(n1070), .B1(n1359), .B2(n4), .ZN(n861) );
  AND2_X1 U1715 ( .A1(n1583), .A2(n656), .ZN(n799) );
  OAI22_X1 U1716 ( .A1(n1514), .A2(n1081), .B1(n1080), .B2(n1354), .ZN(n872)
         );
  INV_X1 U1717 ( .A(n640), .ZN(n680) );
  INV_X1 U1718 ( .A(n368), .ZN(n369) );
  XNOR2_X1 U1719 ( .A(n1582), .B(n1478), .ZN(n1025) );
  INV_X1 U1720 ( .A(n658), .ZN(n800) );
  INV_X1 U1721 ( .A(n1411), .ZN(n1141) );
  INV_X1 U1722 ( .A(n1345), .ZN(n1146) );
  OR2_X1 U1723 ( .A1(n1582), .A2(n1142), .ZN(n942) );
  OR2_X1 U1724 ( .A1(n1582), .A2(n1145), .ZN(n1005) );
  OR2_X1 U1725 ( .A1(n1582), .A2(n1141), .ZN(n921) );
  OR2_X1 U1726 ( .A1(n1583), .A2(n1143), .ZN(n963) );
  OR2_X1 U1727 ( .A1(n1583), .A2(n1144), .ZN(n984) );
  OR2_X1 U1728 ( .A1(n1583), .A2(n1140), .ZN(n900) );
  OR2_X1 U1729 ( .A1(n1583), .A2(n1146), .ZN(n1026) );
  BUF_X2 U1730 ( .A(n61), .Z(n1583) );
  XOR2_X1 U1731 ( .A(n19), .B(a[6]), .Z(n1116) );
  AND2_X1 U1732 ( .A1(n1583), .A2(n1245), .ZN(product[0]) );
  XNOR2_X1 U1733 ( .A(n13), .B(a[6]), .ZN(n22) );
  XNOR2_X1 U1734 ( .A(n1579), .B(a[14]), .ZN(n46) );
  XNOR2_X1 U1735 ( .A(n1580), .B(a[16]), .ZN(n52) );
  XNOR2_X1 U1736 ( .A(n25), .B(a[10]), .ZN(n34) );
  XNOR2_X1 U1737 ( .A(n49), .B(a[18]), .ZN(n58) );
  XNOR2_X1 U1738 ( .A(n1), .B(a[2]), .ZN(n9) );
  XNOR2_X1 U1739 ( .A(n1578), .B(a[4]), .ZN(n1554) );
  XNOR2_X1 U1740 ( .A(n1578), .B(a[4]), .ZN(n1555) );
  INV_X1 U1741 ( .A(n1490), .ZN(n144) );
  NAND2_X1 U1742 ( .A1(n397), .A2(n410), .ZN(n148) );
  NAND2_X1 U1743 ( .A1(n815), .A2(n1260), .ZN(n1556) );
  NAND2_X1 U1744 ( .A1(n815), .A2(n779), .ZN(n1557) );
  NAND2_X1 U1745 ( .A1(n1260), .A2(n779), .ZN(n1558) );
  NAND3_X1 U1746 ( .A1(n1556), .A2(n1557), .A3(n1558), .ZN(n606) );
  AND2_X1 U1747 ( .A1(n1583), .A2(n653), .ZN(n779) );
  OAI22_X1 U1748 ( .A1(n1410), .A2(n1079), .B1(n1078), .B2(n4), .ZN(n870) );
  INV_X1 U1749 ( .A(n1544), .ZN(n1560) );
  NAND2_X1 U1750 ( .A1(n461), .A2(n478), .ZN(n167) );
  XNOR2_X1 U1751 ( .A(n92), .B(n255), .ZN(product[4]) );
  OAI21_X1 U1752 ( .B1(n256), .B2(n258), .A(n257), .ZN(n255) );
  NAND2_X1 U1753 ( .A1(n295), .A2(n257), .ZN(n93) );
  INV_X1 U1754 ( .A(n234), .ZN(n233) );
  OAI21_X1 U1755 ( .B1(n141), .B2(n135), .A(n136), .ZN(n134) );
  XNOR2_X1 U1756 ( .A(n1333), .B(n1344), .ZN(n880) );
  XNOR2_X1 U1757 ( .A(n1378), .B(n1344), .ZN(n881) );
  XNOR2_X1 U1758 ( .A(n1379), .B(n1344), .ZN(n882) );
  XNOR2_X1 U1759 ( .A(n1596), .B(n1344), .ZN(n883) );
  XNOR2_X1 U1760 ( .A(n1594), .B(n1344), .ZN(n885) );
  XNOR2_X1 U1761 ( .A(n1595), .B(n1344), .ZN(n884) );
  XNOR2_X1 U1762 ( .A(n1377), .B(n1344), .ZN(n886) );
  XNOR2_X1 U1763 ( .A(n1369), .B(n1344), .ZN(n887) );
  XNOR2_X1 U1764 ( .A(n1325), .B(n1344), .ZN(n888) );
  XNOR2_X1 U1765 ( .A(n1233), .B(n1581), .ZN(n889) );
  XNOR2_X1 U1766 ( .A(n1592), .B(n1581), .ZN(n890) );
  XNOR2_X1 U1767 ( .A(n1380), .B(n1581), .ZN(n891) );
  XNOR2_X1 U1768 ( .A(n1590), .B(n1581), .ZN(n892) );
  XNOR2_X1 U1769 ( .A(n1582), .B(n1581), .ZN(n899) );
  XNOR2_X1 U1770 ( .A(n1588), .B(n1581), .ZN(n894) );
  XNOR2_X1 U1771 ( .A(n1334), .B(n1581), .ZN(n893) );
  XNOR2_X1 U1772 ( .A(n1108), .B(n1581), .ZN(n898) );
  INV_X1 U1773 ( .A(n1581), .ZN(n1140) );
  XNOR2_X1 U1774 ( .A(n1587), .B(n1581), .ZN(n895) );
  XNOR2_X1 U1775 ( .A(n1585), .B(n1581), .ZN(n897) );
  XNOR2_X1 U1776 ( .A(n1586), .B(n1581), .ZN(n896) );
  INV_X1 U1777 ( .A(n187), .ZN(n282) );
  OAI21_X1 U1778 ( .B1(n193), .B2(n187), .A(n188), .ZN(n186) );
  NOR2_X1 U1779 ( .A1(n529), .A2(n542), .ZN(n187) );
  XNOR2_X1 U1780 ( .A(n1595), .B(n1348), .ZN(n1031) );
  XNOR2_X1 U1781 ( .A(n1356), .B(n1349), .ZN(n1044) );
  INV_X1 U1782 ( .A(n1348), .ZN(n1147) );
  XNOR2_X1 U1783 ( .A(n1380), .B(n1348), .ZN(n1038) );
  XNOR2_X1 U1784 ( .A(n1334), .B(n1348), .ZN(n1040) );
  XNOR2_X1 U1785 ( .A(n1590), .B(n1348), .ZN(n1039) );
  XNOR2_X1 U1786 ( .A(n1377), .B(n1348), .ZN(n1033) );
  XNOR2_X1 U1787 ( .A(n1594), .B(n13), .ZN(n1032) );
  XNOR2_X1 U1788 ( .A(n1596), .B(n1349), .ZN(n1030) );
  XNOR2_X1 U1789 ( .A(n1582), .B(n1348), .ZN(n1046) );
  XNOR2_X1 U1790 ( .A(n1374), .B(n1349), .ZN(n1043) );
  XNOR2_X1 U1791 ( .A(n1355), .B(n1348), .ZN(n1042) );
  XNOR2_X1 U1792 ( .A(n1588), .B(n1349), .ZN(n1041) );
  XNOR2_X1 U1793 ( .A(n1592), .B(n1349), .ZN(n1037) );
  XNOR2_X1 U1794 ( .A(n1333), .B(n1348), .ZN(n1027) );
  XNOR2_X1 U1795 ( .A(n1597), .B(n1349), .ZN(n1029) );
  XNOR2_X1 U1796 ( .A(n1369), .B(n1348), .ZN(n1034) );
  XNOR2_X1 U1797 ( .A(n1598), .B(n1348), .ZN(n1028) );
  XNOR2_X1 U1798 ( .A(n1584), .B(n1348), .ZN(n1045) );
  XNOR2_X1 U1799 ( .A(n1593), .B(n1348), .ZN(n1036) );
  XNOR2_X1 U1800 ( .A(n1325), .B(n1349), .ZN(n1035) );
  AND2_X1 U1801 ( .A1(n513), .A2(n528), .ZN(n1561) );
  OR2_X1 U1802 ( .A1(n1583), .A2(n1148), .ZN(n1068) );
  CLKBUF_X1 U1803 ( .A(n1567), .Z(n1562) );
  NAND3_X1 U1804 ( .A1(n1567), .A2(n1568), .A3(n1566), .ZN(n1563) );
  NAND3_X1 U1805 ( .A1(n1507), .A2(n1562), .A3(n1566), .ZN(n1564) );
  XOR2_X1 U1806 ( .A(n307), .B(n310), .Z(n1565) );
  NAND2_X1 U1807 ( .A1(n307), .A2(n310), .ZN(n1566) );
  NAND2_X1 U1808 ( .A1(n264), .A2(n307), .ZN(n1567) );
  NAND2_X1 U1809 ( .A1(n264), .A2(n310), .ZN(n1568) );
  NAND3_X1 U1810 ( .A1(n1568), .A2(n1567), .A3(n1566), .ZN(n100) );
  NAND2_X1 U1811 ( .A1(n303), .A2(n306), .ZN(n1569) );
  NAND2_X1 U1812 ( .A1(n1563), .A2(n303), .ZN(n1570) );
  NAND2_X1 U1813 ( .A1(n306), .A2(n100), .ZN(n1571) );
  NAND3_X1 U1814 ( .A1(n1571), .A2(n1570), .A3(n1569), .ZN(n99) );
  INV_X1 U1815 ( .A(n664), .ZN(n840) );
  AOI21_X1 U1816 ( .B1(n146), .B2(n133), .A(n134), .ZN(n132) );
  NAND2_X1 U1817 ( .A1(n156), .A2(n164), .ZN(n154) );
  XNOR2_X1 U1818 ( .A(n1333), .B(n1360), .ZN(n943) );
  XNOR2_X1 U1819 ( .A(n1378), .B(n1362), .ZN(n944) );
  XNOR2_X1 U1820 ( .A(n1596), .B(n1350), .ZN(n946) );
  XNOR2_X1 U1821 ( .A(n1379), .B(n1351), .ZN(n945) );
  XNOR2_X1 U1822 ( .A(n1595), .B(n1350), .ZN(n947) );
  XNOR2_X1 U1823 ( .A(n1594), .B(n1351), .ZN(n948) );
  XNOR2_X1 U1824 ( .A(n1593), .B(n1350), .ZN(n952) );
  XNOR2_X1 U1825 ( .A(n1325), .B(n1350), .ZN(n951) );
  XNOR2_X1 U1826 ( .A(n1589), .B(n1351), .ZN(n956) );
  XNOR2_X1 U1827 ( .A(n1590), .B(n1361), .ZN(n955) );
  INV_X1 U1828 ( .A(n1360), .ZN(n1143) );
  XNOR2_X1 U1829 ( .A(n1370), .B(n1362), .ZN(n950) );
  XNOR2_X1 U1830 ( .A(n1377), .B(n1351), .ZN(n949) );
  XNOR2_X1 U1831 ( .A(n1588), .B(n1362), .ZN(n957) );
  XNOR2_X1 U1832 ( .A(n1356), .B(n1360), .ZN(n960) );
  XNOR2_X1 U1833 ( .A(n1592), .B(n1361), .ZN(n953) );
  XNOR2_X1 U1834 ( .A(n1591), .B(n1361), .ZN(n954) );
  XNOR2_X1 U1835 ( .A(n1582), .B(n1351), .ZN(n962) );
  XNOR2_X1 U1836 ( .A(n1584), .B(n1350), .ZN(n961) );
  INV_X1 U1837 ( .A(n1390), .ZN(n284) );
  NOR2_X1 U1838 ( .A1(n1390), .A2(n209), .ZN(n202) );
  OAI21_X1 U1839 ( .B1(n204), .B2(n210), .A(n205), .ZN(n203) );
  NAND2_X1 U1840 ( .A1(n557), .A2(n568), .ZN(n205) );
  XNOR2_X1 U1841 ( .A(n1333), .B(n1394), .ZN(n985) );
  XNOR2_X1 U1842 ( .A(n1598), .B(n1347), .ZN(n986) );
  XNOR2_X1 U1843 ( .A(n1377), .B(n1394), .ZN(n991) );
  XNOR2_X1 U1844 ( .A(n1594), .B(n1394), .ZN(n990) );
  XNOR2_X1 U1845 ( .A(n1595), .B(n1394), .ZN(n989) );
  XNOR2_X1 U1846 ( .A(n1596), .B(n1347), .ZN(n988) );
  XNOR2_X1 U1847 ( .A(n1582), .B(n1394), .ZN(n1004) );
  XNOR2_X1 U1848 ( .A(n1597), .B(n1347), .ZN(n987) );
  XNOR2_X1 U1849 ( .A(n1370), .B(n1347), .ZN(n992) );
  XNOR2_X1 U1850 ( .A(n1588), .B(n1394), .ZN(n999) );
  INV_X1 U1851 ( .A(n1347), .ZN(n1145) );
  XNOR2_X1 U1852 ( .A(n1584), .B(n1347), .ZN(n1003) );
  XNOR2_X1 U1853 ( .A(n1592), .B(n1347), .ZN(n995) );
  XNOR2_X1 U1854 ( .A(n1325), .B(n1394), .ZN(n993) );
  XNOR2_X1 U1855 ( .A(n1593), .B(n1394), .ZN(n994) );
  XNOR2_X1 U1856 ( .A(n1356), .B(n1394), .ZN(n1002) );
  XNOR2_X1 U1857 ( .A(n1589), .B(n1347), .ZN(n998) );
  XNOR2_X1 U1858 ( .A(n1590), .B(n1347), .ZN(n997) );
  XNOR2_X1 U1859 ( .A(n1587), .B(n1394), .ZN(n1000) );
  XNOR2_X1 U1860 ( .A(n1373), .B(n1347), .ZN(n1001) );
  XNOR2_X1 U1861 ( .A(n1591), .B(n1347), .ZN(n996) );
  XNOR2_X1 U1862 ( .A(n1588), .B(n1398), .ZN(n1062) );
  XNOR2_X1 U1863 ( .A(n1380), .B(n1398), .ZN(n1059) );
  INV_X1 U1864 ( .A(n1398), .ZN(n1148) );
  XNOR2_X1 U1865 ( .A(n1597), .B(n1398), .ZN(n1050) );
  XNOR2_X1 U1866 ( .A(n1598), .B(n1398), .ZN(n1049) );
  XNOR2_X1 U1867 ( .A(n1595), .B(n1398), .ZN(n1052) );
  XNOR2_X1 U1868 ( .A(n1596), .B(n1398), .ZN(n1051) );
  XNOR2_X1 U1869 ( .A(n1374), .B(n1398), .ZN(n1064) );
  XNOR2_X1 U1870 ( .A(n1334), .B(n1398), .ZN(n1061) );
  XNOR2_X1 U1871 ( .A(n1590), .B(n1398), .ZN(n1060) );
  XNOR2_X1 U1872 ( .A(n1355), .B(n1398), .ZN(n1063) );
  XNOR2_X1 U1873 ( .A(n1325), .B(n1398), .ZN(n1056) );
  XNOR2_X1 U1874 ( .A(n1370), .B(n1398), .ZN(n1055) );
  XNOR2_X1 U1875 ( .A(n1377), .B(n1398), .ZN(n1054) );
  XNOR2_X1 U1876 ( .A(n1582), .B(n1398), .ZN(n1067) );
  XNOR2_X1 U1877 ( .A(n1584), .B(n1398), .ZN(n1066) );
  XNOR2_X1 U1878 ( .A(n1594), .B(n1398), .ZN(n1053) );
  XNOR2_X1 U1879 ( .A(n1356), .B(n1398), .ZN(n1065) );
  XNOR2_X1 U1880 ( .A(n1592), .B(n1398), .ZN(n1058) );
  XNOR2_X1 U1881 ( .A(n1593), .B(n1398), .ZN(n1057) );
  XNOR2_X1 U1882 ( .A(n1333), .B(n1398), .ZN(n1048) );
  NAND2_X1 U1883 ( .A1(n755), .A2(n864), .ZN(n1572) );
  NAND2_X1 U1884 ( .A1(n755), .A2(n719), .ZN(n1573) );
  NAND2_X1 U1885 ( .A1(n864), .A2(n719), .ZN(n1574) );
  NAND3_X1 U1886 ( .A1(n1572), .A2(n1573), .A3(n1574), .ZN(n540) );
  OR2_X1 U1887 ( .A1(n1432), .A2(n959), .ZN(n1575) );
  OR2_X1 U1888 ( .A1(n958), .A2(n1368), .ZN(n1576) );
  NAND2_X1 U1889 ( .A1(n1575), .A2(n1576), .ZN(n755) );
  AND2_X1 U1890 ( .A1(n1583), .A2(n644), .ZN(n719) );
  OAI22_X1 U1891 ( .A1(n1514), .A2(n1073), .B1(n1072), .B2(n4), .ZN(n864) );
  XNOR2_X1 U1892 ( .A(n1586), .B(n1351), .ZN(n959) );
  XNOR2_X1 U1893 ( .A(n1587), .B(n1350), .ZN(n958) );
  NOR2_X1 U1894 ( .A1(n140), .A2(n135), .ZN(n133) );
  NOR2_X1 U1895 ( .A1(n383), .A2(n396), .ZN(n140) );
  INV_X1 U1896 ( .A(n661), .ZN(n820) );
  XNOR2_X1 U1897 ( .A(n239), .B(n88), .ZN(product[8]) );
  AOI21_X1 U1898 ( .B1(n239), .B2(n1538), .A(n236), .ZN(n234) );
  NAND2_X1 U1899 ( .A1(n637), .A2(n638), .ZN(n254) );
  XOR2_X1 U1900 ( .A(n242), .B(n89), .Z(product[7]) );
  OAI21_X1 U1901 ( .B1(n242), .B2(n240), .A(n241), .ZN(n239) );
  XNOR2_X1 U1902 ( .A(n1380), .B(n1577), .ZN(n1080) );
  XNOR2_X1 U1903 ( .A(n1590), .B(n1577), .ZN(n1081) );
  XNOR2_X1 U1904 ( .A(n1377), .B(n1357), .ZN(n1075) );
  XNOR2_X1 U1905 ( .A(n1597), .B(n1357), .ZN(n1071) );
  XNOR2_X1 U1906 ( .A(n1592), .B(n1357), .ZN(n1079) );
  XNOR2_X1 U1907 ( .A(n1598), .B(n1357), .ZN(n1070) );
  XNOR2_X1 U1908 ( .A(n1593), .B(n1357), .ZN(n1078) );
  XNOR2_X1 U1909 ( .A(n1594), .B(n1357), .ZN(n1074) );
  XNOR2_X1 U1910 ( .A(n1369), .B(n1357), .ZN(n1076) );
  XNOR2_X1 U1911 ( .A(n1596), .B(n1357), .ZN(n1072) );
  XNOR2_X1 U1912 ( .A(n1325), .B(n1577), .ZN(n1077) );
  XNOR2_X1 U1913 ( .A(n1595), .B(n1357), .ZN(n1073) );
  XNOR2_X1 U1914 ( .A(n1334), .B(n1357), .ZN(n1082) );
  XNOR2_X1 U1915 ( .A(n1588), .B(n1357), .ZN(n1083) );
  XNOR2_X1 U1916 ( .A(n1599), .B(n1308), .ZN(n1069) );
  XNOR2_X1 U1917 ( .A(n1582), .B(n1577), .ZN(n1088) );
  XNOR2_X1 U1918 ( .A(n1356), .B(n1577), .ZN(n1086) );
  XNOR2_X1 U1919 ( .A(n1373), .B(n1577), .ZN(n1085) );
  XNOR2_X1 U1920 ( .A(n1584), .B(n1577), .ZN(n1087) );
  XNOR2_X1 U1921 ( .A(n1587), .B(n1577), .ZN(n1084) );
  INV_X1 U1922 ( .A(n1357), .ZN(n1149) );
  XOR2_X1 U1923 ( .A(n1), .B(n668), .Z(n1119) );
  OAI21_X1 U1924 ( .B1(n152), .B2(n131), .A(n1406), .ZN(n130) );
  NAND2_X1 U1925 ( .A1(n1532), .A2(n200), .ZN(n81) );
  NAND2_X1 U1926 ( .A1(n202), .A2(n1532), .ZN(n195) );
  NAND2_X1 U1927 ( .A1(n543), .A2(n556), .ZN(n200) );
  OAI21_X1 U1928 ( .B1(n152), .B2(n150), .A(n151), .ZN(n149) );
  INV_X1 U1929 ( .A(n150), .ZN(n275) );
  NOR2_X1 U1930 ( .A1(n1518), .A2(n150), .ZN(n145) );
  NAND2_X1 U1931 ( .A1(n411), .A2(n426), .ZN(n151) );
  INV_X1 U1932 ( .A(n1417), .ZN(n276) );
  OAI21_X1 U1933 ( .B1(n158), .B2(n162), .A(n159), .ZN(n157) );
  NAND2_X1 U1934 ( .A1(n427), .A2(n442), .ZN(n159) );
  OAI21_X1 U1935 ( .B1(n222), .B2(n234), .A(n223), .ZN(n221) );
  AOI21_X1 U1936 ( .B1(n1531), .B2(n190), .A(n1561), .ZN(n181) );
  INV_X1 U1937 ( .A(n188), .ZN(n190) );
  OAI21_X1 U1938 ( .B1(n163), .B2(n161), .A(n162), .ZN(n160) );
  INV_X1 U1939 ( .A(n161), .ZN(n277) );
  NOR2_X1 U1940 ( .A1(n1512), .A2(n161), .ZN(n156) );
  OR2_X1 U1941 ( .A1(n787), .A2(n715), .ZN(n476) );
  XNOR2_X1 U1942 ( .A(n715), .B(n787), .ZN(n477) );
  INV_X1 U1943 ( .A(n1246), .ZN(n211) );
  NOR2_X1 U1944 ( .A1(n1515), .A2(n180), .ZN(n175) );
  OAI22_X1 U1945 ( .A1(n880), .A2(n1491), .B1(n880), .B2(n1244), .ZN(n640) );
  OAI22_X1 U1946 ( .A1(n1491), .A2(n881), .B1(n880), .B2(n1244), .ZN(n298) );
  OAI22_X1 U1947 ( .A1(n1491), .A2(n882), .B1(n881), .B2(n1244), .ZN(n681) );
  OAI22_X1 U1948 ( .A1(n1491), .A2(n883), .B1(n882), .B2(n1244), .ZN(n682) );
  OAI22_X1 U1949 ( .A1(n1491), .A2(n884), .B1(n883), .B2(n1244), .ZN(n683) );
  OAI22_X1 U1950 ( .A1(n1491), .A2(n886), .B1(n885), .B2(n1341), .ZN(n685) );
  OAI22_X1 U1951 ( .A1(n1491), .A2(n885), .B1(n884), .B2(n1244), .ZN(n684) );
  OAI22_X1 U1952 ( .A1(n1491), .A2(n887), .B1(n886), .B2(n1341), .ZN(n686) );
  OAI22_X1 U1953 ( .A1(n1491), .A2(n888), .B1(n887), .B2(n1341), .ZN(n687) );
  OAI22_X1 U1954 ( .A1(n1385), .A2(n889), .B1(n888), .B2(n1341), .ZN(n688) );
  OAI22_X1 U1955 ( .A1(n1386), .A2(n890), .B1(n889), .B2(n1341), .ZN(n689) );
  OAI22_X1 U1956 ( .A1(n1386), .A2(n891), .B1(n890), .B2(n1341), .ZN(n690) );
  OAI22_X1 U1957 ( .A1(n1385), .A2(n892), .B1(n891), .B2(n1341), .ZN(n691) );
  OAI22_X1 U1958 ( .A1(n1385), .A2(n894), .B1(n893), .B2(n1341), .ZN(n693) );
  OAI22_X1 U1959 ( .A1(n1385), .A2(n893), .B1(n892), .B2(n1341), .ZN(n692) );
  OAI22_X1 U1960 ( .A1(n1386), .A2(n895), .B1(n894), .B2(n1341), .ZN(n694) );
  OAI22_X1 U1961 ( .A1(n1386), .A2(n899), .B1(n898), .B2(n1341), .ZN(n698) );
  OAI22_X1 U1962 ( .A1(n1386), .A2(n896), .B1(n895), .B2(n1341), .ZN(n695) );
  OAI22_X1 U1963 ( .A1(n1386), .A2(n1140), .B1(n900), .B2(n1341), .ZN(n670) );
  INV_X1 U1964 ( .A(n1341), .ZN(n641) );
  OAI22_X1 U1965 ( .A1(n60), .A2(n898), .B1(n897), .B2(n1341), .ZN(n697) );
  OAI22_X1 U1966 ( .A1(n60), .A2(n897), .B1(n896), .B2(n1341), .ZN(n696) );
  AOI21_X1 U1967 ( .B1(n1520), .B2(n1303), .A(n1506), .ZN(n125) );
  OAI21_X1 U1968 ( .B1(n132), .B2(n128), .A(n129), .ZN(n127) );
  INV_X1 U1969 ( .A(n221), .ZN(n220) );
  INV_X1 U1970 ( .A(n1381), .ZN(n193) );
  AOI21_X1 U1971 ( .B1(n194), .B2(n175), .A(n176), .ZN(n174) );
  NAND2_X1 U1972 ( .A1(n639), .A2(n678), .ZN(n257) );
  OAI22_X1 U1973 ( .A1(n1459), .A2(n1055), .B1(n1054), .B2(n1552), .ZN(n846)
         );
  OAI22_X1 U1974 ( .A1(n1264), .A2(n1053), .B1(n1052), .B2(n1553), .ZN(n844)
         );
  OAI22_X1 U1975 ( .A1(n1459), .A2(n1059), .B1(n1058), .B2(n1552), .ZN(n850)
         );
  OAI22_X1 U1976 ( .A1(n1264), .A2(n1062), .B1(n1061), .B2(n1553), .ZN(n853)
         );
  OAI22_X1 U1977 ( .A1(n1519), .A2(n1051), .B1(n1050), .B2(n1552), .ZN(n842)
         );
  OAI22_X1 U1978 ( .A1(n1264), .A2(n1060), .B1(n1059), .B2(n1553), .ZN(n851)
         );
  OAI22_X1 U1979 ( .A1(n1264), .A2(n1063), .B1(n1062), .B2(n1552), .ZN(n854)
         );
  OAI22_X1 U1980 ( .A1(n1264), .A2(n1057), .B1(n1056), .B2(n1553), .ZN(n848)
         );
  OAI22_X1 U1981 ( .A1(n1459), .A2(n1052), .B1(n1051), .B2(n1552), .ZN(n843)
         );
  OAI22_X1 U1982 ( .A1(n1458), .A2(n1058), .B1(n1057), .B2(n1552), .ZN(n849)
         );
  OAI22_X1 U1983 ( .A1(n1519), .A2(n1049), .B1(n1239), .B2(n1552), .ZN(n458)
         );
  OAI22_X1 U1984 ( .A1(n1264), .A2(n1056), .B1(n1055), .B2(n1553), .ZN(n847)
         );
  OAI22_X1 U1985 ( .A1(n1458), .A2(n1065), .B1(n1064), .B2(n1553), .ZN(n856)
         );
  OAI22_X1 U1986 ( .A1(n1459), .A2(n1054), .B1(n1053), .B2(n1553), .ZN(n845)
         );
  OAI22_X1 U1987 ( .A1(n1519), .A2(n1050), .B1(n1049), .B2(n1553), .ZN(n841)
         );
  OAI22_X1 U1988 ( .A1(n1458), .A2(n1148), .B1(n1068), .B2(n1552), .ZN(n678)
         );
  OAI22_X1 U1989 ( .A1(n1458), .A2(n1061), .B1(n1060), .B2(n1553), .ZN(n852)
         );
  OAI22_X1 U1990 ( .A1(n1459), .A2(n1064), .B1(n1063), .B2(n1552), .ZN(n855)
         );
  OAI22_X1 U1991 ( .A1(n1460), .A2(n1239), .B1(n1048), .B2(n1553), .ZN(n664)
         );
  INV_X1 U1992 ( .A(n1552), .ZN(n665) );
  OAI22_X1 U1993 ( .A1(n1264), .A2(n1066), .B1(n1065), .B2(n1552), .ZN(n857)
         );
  OAI22_X1 U1994 ( .A1(n1458), .A2(n1067), .B1(n1066), .B2(n1553), .ZN(n858)
         );
  INV_X1 U1995 ( .A(n145), .ZN(n143) );
  OAI22_X1 U1996 ( .A1(n901), .A2(n1412), .B1(n901), .B2(n1549), .ZN(n643) );
  OAI22_X1 U1997 ( .A1(n1412), .A2(n902), .B1(n901), .B2(n1550), .ZN(n304) );
  OAI22_X1 U1998 ( .A1(n1412), .A2(n903), .B1(n902), .B2(n1549), .ZN(n701) );
  OAI22_X1 U1999 ( .A1(n1412), .A2(n905), .B1(n904), .B2(n1550), .ZN(n703) );
  OAI22_X1 U2000 ( .A1(n1412), .A2(n904), .B1(n903), .B2(n1549), .ZN(n702) );
  OAI22_X1 U2001 ( .A1(n1412), .A2(n906), .B1(n905), .B2(n1550), .ZN(n704) );
  OAI22_X1 U2002 ( .A1(n1412), .A2(n907), .B1(n906), .B2(n1549), .ZN(n705) );
  OAI22_X1 U2003 ( .A1(n1412), .A2(n908), .B1(n907), .B2(n1550), .ZN(n706) );
  OAI22_X1 U2004 ( .A1(n1412), .A2(n909), .B1(n908), .B2(n1549), .ZN(n707) );
  OAI22_X1 U2005 ( .A1(n54), .A2(n910), .B1(n909), .B2(n1550), .ZN(n708) );
  OAI22_X1 U2006 ( .A1(n54), .A2(n911), .B1(n910), .B2(n1549), .ZN(n709) );
  OAI22_X1 U2007 ( .A1(n54), .A2(n1141), .B1(n921), .B2(n1550), .ZN(n671) );
  OAI22_X1 U2008 ( .A1(n54), .A2(n915), .B1(n914), .B2(n1549), .ZN(n713) );
  OAI22_X1 U2009 ( .A1(n54), .A2(n914), .B1(n913), .B2(n1550), .ZN(n712) );
  OAI22_X1 U2010 ( .A1(n54), .A2(n919), .B1(n918), .B2(n1549), .ZN(n717) );
  OAI22_X1 U2011 ( .A1(n54), .A2(n920), .B1(n919), .B2(n1550), .ZN(n718) );
  OAI22_X1 U2012 ( .A1(n54), .A2(n918), .B1(n917), .B2(n1550), .ZN(n716) );
  OAI22_X1 U2013 ( .A1(n54), .A2(n912), .B1(n911), .B2(n1550), .ZN(n710) );
  OAI22_X1 U2014 ( .A1(n54), .A2(n913), .B1(n912), .B2(n1549), .ZN(n711) );
  INV_X1 U2015 ( .A(n1549), .ZN(n644) );
  OAI22_X1 U2016 ( .A1(n54), .A2(n917), .B1(n916), .B2(n1550), .ZN(n715) );
  OAI21_X1 U2017 ( .B1(n193), .B2(n180), .A(n1269), .ZN(n179) );
  OAI21_X1 U2018 ( .B1(n181), .B2(n177), .A(n178), .ZN(n176) );
  OAI22_X1 U2019 ( .A1(n943), .A2(n1358), .B1(n943), .B2(n1342), .ZN(n649) );
  OAI22_X1 U2020 ( .A1(n1433), .A2(n944), .B1(n943), .B2(n1367), .ZN(n328) );
  OAI22_X1 U2021 ( .A1(n1358), .A2(n945), .B1(n944), .B2(n1342), .ZN(n741) );
  OAI22_X1 U2022 ( .A1(n1433), .A2(n947), .B1(n946), .B2(n1266), .ZN(n743) );
  OAI22_X1 U2023 ( .A1(n1358), .A2(n946), .B1(n945), .B2(n1342), .ZN(n742) );
  OAI22_X1 U2024 ( .A1(n1433), .A2(n948), .B1(n947), .B2(n1342), .ZN(n744) );
  OAI22_X1 U2025 ( .A1(n1358), .A2(n949), .B1(n948), .B2(n1342), .ZN(n745) );
  OAI22_X1 U2026 ( .A1(n1433), .A2(n952), .B1(n951), .B2(n1367), .ZN(n748) );
  OAI22_X1 U2027 ( .A1(n957), .A2(n1432), .B1(n956), .B2(n1559), .ZN(n753) );
  OAI22_X1 U2028 ( .A1(n1432), .A2(n958), .B1(n957), .B2(n1266), .ZN(n754) );
  OAI22_X1 U2029 ( .A1(n1432), .A2(n953), .B1(n952), .B2(n1368), .ZN(n749) );
  OAI22_X1 U2030 ( .A1(n1433), .A2(n1143), .B1(n963), .B2(n1367), .ZN(n673) );
  OAI22_X1 U2031 ( .A1(n956), .A2(n1432), .B1(n955), .B2(n1266), .ZN(n752) );
  OAI22_X1 U2032 ( .A1(n1433), .A2(n951), .B1(n950), .B2(n1559), .ZN(n747) );
  INV_X1 U2033 ( .A(n1559), .ZN(n650) );
  OAI22_X1 U2034 ( .A1(n1433), .A2(n960), .B1(n959), .B2(n1367), .ZN(n756) );
  OAI22_X1 U2035 ( .A1(n1432), .A2(n950), .B1(n949), .B2(n1559), .ZN(n746) );
  OAI22_X1 U2036 ( .A1(n1433), .A2(n961), .B1(n960), .B2(n1266), .ZN(n757) );
  OAI22_X1 U2037 ( .A1(n42), .A2(n954), .B1(n953), .B2(n1368), .ZN(n750) );
  OAI22_X1 U2038 ( .A1(n42), .A2(n962), .B1(n961), .B2(n1559), .ZN(n758) );
  AOI21_X1 U2039 ( .B1(n211), .B2(n202), .A(n203), .ZN(n201) );
  OAI21_X1 U2040 ( .B1(n195), .B2(n212), .A(n196), .ZN(n194) );
  AOI21_X1 U2041 ( .B1(n203), .B2(n1532), .A(n198), .ZN(n196) );
  OAI22_X1 U2042 ( .A1(n1510), .A2(n965), .B1(n964), .B2(n1376), .ZN(n346) );
  OAI22_X1 U2043 ( .A1(n964), .A2(n1510), .B1(n964), .B2(n1375), .ZN(n652) );
  OAI22_X1 U2044 ( .A1(n1510), .A2(n966), .B1(n965), .B2(n1375), .ZN(n761) );
  OAI22_X1 U2045 ( .A1(n1510), .A2(n967), .B1(n966), .B2(n1376), .ZN(n762) );
  OAI22_X1 U2046 ( .A1(n1389), .A2(n968), .B1(n967), .B2(n1375), .ZN(n763) );
  OAI22_X1 U2047 ( .A1(n1388), .A2(n1243), .B1(n974), .B2(n1376), .ZN(n770) );
  OAI22_X1 U2048 ( .A1(n1389), .A2(n973), .B1(n972), .B2(n1376), .ZN(n768) );
  OAI22_X1 U2049 ( .A1(n1510), .A2(n972), .B1(n971), .B2(n1376), .ZN(n767) );
  OAI22_X1 U2050 ( .A1(n1389), .A2(n977), .B1(n976), .B2(n1376), .ZN(n772) );
  OAI22_X1 U2051 ( .A1(n1389), .A2(n971), .B1(n970), .B2(n1375), .ZN(n766) );
  OAI22_X1 U2052 ( .A1(n1336), .A2(n976), .B1(n975), .B2(n1376), .ZN(n771) );
  OAI22_X1 U2053 ( .A1(n1388), .A2(n970), .B1(n969), .B2(n1375), .ZN(n765) );
  OAI22_X1 U2054 ( .A1(n1388), .A2(n969), .B1(n968), .B2(n1376), .ZN(n764) );
  OAI22_X1 U2055 ( .A1(n1389), .A2(n1144), .B1(n984), .B2(n1375), .ZN(n674) );
  OAI22_X1 U2056 ( .A1(n1336), .A2(n983), .B1(n982), .B2(n1375), .ZN(n778) );
  OAI22_X1 U2057 ( .A1(n1389), .A2(n978), .B1(n977), .B2(n1376), .ZN(n773) );
  OAI22_X1 U2058 ( .A1(n1443), .A2(n974), .B1(n973), .B2(n1376), .ZN(n769) );
  OAI22_X1 U2059 ( .A1(n1336), .A2(n982), .B1(n981), .B2(n1375), .ZN(n777) );
  OAI22_X1 U2060 ( .A1(n1443), .A2(n979), .B1(n978), .B2(n1375), .ZN(n774) );
  OAI22_X1 U2061 ( .A1(n1443), .A2(n980), .B1(n979), .B2(n1376), .ZN(n775) );
  OAI22_X1 U2062 ( .A1(n1336), .A2(n981), .B1(n980), .B2(n1375), .ZN(n776) );
  INV_X1 U2063 ( .A(n1375), .ZN(n653) );
  OAI21_X1 U2064 ( .B1(n151), .B2(n147), .A(n148), .ZN(n146) );
  INV_X1 U2065 ( .A(n1242), .ZN(n278) );
  AOI21_X1 U2066 ( .B1(n173), .B2(n164), .A(n1339), .ZN(n163) );
  OAI22_X1 U2067 ( .A1(n922), .A2(n1522), .B1(n922), .B2(n1548), .ZN(n646) );
  AOI21_X1 U2068 ( .B1(n165), .B2(n156), .A(n157), .ZN(n155) );
  NOR2_X1 U2069 ( .A1(n171), .A2(n1242), .ZN(n164) );
  OAI22_X1 U2070 ( .A1(n1522), .A2(n924), .B1(n923), .B2(n1365), .ZN(n721) );
  OAI21_X1 U2071 ( .B1(n166), .B2(n172), .A(n167), .ZN(n165) );
  OAI22_X1 U2072 ( .A1(n1522), .A2(n923), .B1(n922), .B2(n1548), .ZN(n314) );
  OAI22_X1 U2073 ( .A1(n1522), .A2(n925), .B1(n924), .B2(n1365), .ZN(n722) );
  OAI22_X1 U2074 ( .A1(n1522), .A2(n927), .B1(n926), .B2(n1548), .ZN(n724) );
  OAI22_X1 U2075 ( .A1(n1522), .A2(n926), .B1(n925), .B2(n1365), .ZN(n723) );
  OAI22_X1 U2076 ( .A1(n1522), .A2(n928), .B1(n927), .B2(n1548), .ZN(n725) );
  OAI22_X1 U2077 ( .A1(n1522), .A2(n929), .B1(n928), .B2(n1365), .ZN(n726) );
  OAI22_X1 U2078 ( .A1(n1522), .A2(n930), .B1(n929), .B2(n1548), .ZN(n727) );
  OAI22_X1 U2079 ( .A1(n1521), .A2(n931), .B1(n930), .B2(n1365), .ZN(n728) );
  OAI22_X1 U2080 ( .A1(n1522), .A2(n933), .B1(n932), .B2(n1548), .ZN(n730) );
  OAI22_X1 U2081 ( .A1(n1521), .A2(n934), .B1(n933), .B2(n1548), .ZN(n731) );
  OAI22_X1 U2082 ( .A1(n1521), .A2(n932), .B1(n931), .B2(n1365), .ZN(n729) );
  OAI22_X1 U2083 ( .A1(n1522), .A2(n941), .B1(n940), .B2(n1365), .ZN(n738) );
  OAI22_X1 U2084 ( .A1(n1352), .A2(n1142), .B1(n942), .B2(n1365), .ZN(n672) );
  OAI22_X1 U2085 ( .A1(n1522), .A2(n939), .B1(n938), .B2(n1548), .ZN(n736) );
  OAI22_X1 U2086 ( .A1(n1521), .A2(n940), .B1(n939), .B2(n1548), .ZN(n737) );
  OAI22_X1 U2087 ( .A1(n1352), .A2(n937), .B1(n936), .B2(n1365), .ZN(n734) );
  OAI22_X1 U2088 ( .A1(n1352), .A2(n935), .B1(n934), .B2(n1548), .ZN(n732) );
  OAI22_X1 U2089 ( .A1(n1352), .A2(n938), .B1(n937), .B2(n1365), .ZN(n735) );
  INV_X1 U2090 ( .A(n1548), .ZN(n647) );
  INV_X1 U2091 ( .A(n1384), .ZN(n173) );
  OAI22_X1 U2092 ( .A1(n985), .A2(n1457), .B1(n985), .B2(n1332), .ZN(n655) );
  OAI22_X1 U2093 ( .A1(n1457), .A2(n986), .B1(n985), .B2(n1332), .ZN(n368) );
  OAI22_X1 U2094 ( .A1(n1457), .A2(n987), .B1(n986), .B2(n1332), .ZN(n781) );
  OAI22_X1 U2095 ( .A1(n1457), .A2(n1003), .B1(n1002), .B2(n1332), .ZN(n797)
         );
  OAI22_X1 U2096 ( .A1(n1457), .A2(n992), .B1(n991), .B2(n1382), .ZN(n786) );
  OAI22_X1 U2097 ( .A1(n1457), .A2(n989), .B1(n988), .B2(n1382), .ZN(n783) );
  OAI22_X1 U2098 ( .A1(n1457), .A2(n990), .B1(n989), .B2(n1332), .ZN(n784) );
  OAI22_X1 U2099 ( .A1(n1456), .A2(n991), .B1(n990), .B2(n1382), .ZN(n785) );
  OAI22_X1 U2100 ( .A1(n1456), .A2(n988), .B1(n987), .B2(n1382), .ZN(n782) );
  OAI22_X1 U2101 ( .A1(n1457), .A2(n999), .B1(n998), .B2(n1332), .ZN(n793) );
  OAI22_X1 U2102 ( .A1(n1457), .A2(n996), .B1(n995), .B2(n1382), .ZN(n790) );
  OAI22_X1 U2103 ( .A1(n1457), .A2(n1000), .B1(n999), .B2(n1382), .ZN(n794) );
  OAI22_X1 U2104 ( .A1(n1457), .A2(n993), .B1(n992), .B2(n1382), .ZN(n787) );
  OAI22_X1 U2105 ( .A1(n1457), .A2(n1004), .B1(n1003), .B2(n1332), .ZN(n798)
         );
  OAI22_X1 U2106 ( .A1(n1456), .A2(n995), .B1(n1328), .B2(n1382), .ZN(n789) );
  OAI22_X1 U2107 ( .A1(n1457), .A2(n1002), .B1(n1001), .B2(n1382), .ZN(n796)
         );
  OAI22_X1 U2108 ( .A1(n30), .A2(n994), .B1(n993), .B2(n1382), .ZN(n788) );
  OAI22_X1 U2109 ( .A1(n1457), .A2(n1145), .B1(n1005), .B2(n1332), .ZN(n675)
         );
  OAI22_X1 U2110 ( .A1(n1456), .A2(n998), .B1(n997), .B2(n1382), .ZN(n792) );
  OAI22_X1 U2111 ( .A1(n30), .A2(n997), .B1(n996), .B2(n1382), .ZN(n791) );
  OAI22_X1 U2112 ( .A1(n30), .A2(n1001), .B1(n1000), .B2(n1382), .ZN(n795) );
  AOI21_X1 U2113 ( .B1(n1516), .B2(n1536), .A(n111), .ZN(n109) );
  OAI21_X1 U2114 ( .B1(n174), .B2(n154), .A(n155), .ZN(n153) );
  XNOR2_X1 U2115 ( .A(n1509), .B(n67), .ZN(product[29]) );
  XOR2_X1 U2116 ( .A(n109), .B(n64), .Z(product[32]) );
  XOR2_X1 U2117 ( .A(n125), .B(n68), .Z(product[28]) );
  OAI21_X1 U2118 ( .B1(n1529), .B2(n123), .A(n124), .ZN(n122) );
  OAI22_X1 U2119 ( .A1(n1392), .A2(n1014), .B1(n1013), .B2(n1546), .ZN(n807)
         );
  OAI22_X1 U2120 ( .A1(n1392), .A2(n1007), .B1(n1006), .B2(n1546), .ZN(n394)
         );
  OAI22_X1 U2121 ( .A1(n1392), .A2(n1012), .B1(n1011), .B2(n1546), .ZN(n805)
         );
  OAI22_X1 U2122 ( .A1(n1006), .A2(n1392), .B1(n1006), .B2(n1546), .ZN(n658)
         );
  OAI22_X1 U2123 ( .A1(n24), .A2(n1024), .B1(n1023), .B2(n1547), .ZN(n817) );
  OAI22_X1 U2124 ( .A1(n1392), .A2(n1021), .B1(n1020), .B2(n1546), .ZN(n814)
         );
  OAI22_X1 U2125 ( .A1(n1392), .A2(n1008), .B1(n1007), .B2(n1546), .ZN(n801)
         );
  OAI22_X1 U2126 ( .A1(n1010), .A2(n1393), .B1(n1009), .B2(n1547), .ZN(n803)
         );
  OAI22_X1 U2127 ( .A1(n1393), .A2(n1009), .B1(n1008), .B2(n1547), .ZN(n802)
         );
  OAI22_X1 U2128 ( .A1(n1392), .A2(n1146), .B1(n1026), .B2(n1547), .ZN(n676)
         );
  OAI22_X1 U2129 ( .A1(n1393), .A2(n1015), .B1(n1014), .B2(n1547), .ZN(n808)
         );
  OAI22_X1 U2130 ( .A1(n1013), .A2(n24), .B1(n1012), .B2(n1546), .ZN(n806) );
  OAI22_X1 U2131 ( .A1(n1393), .A2(n1025), .B1(n1024), .B2(n1547), .ZN(n818)
         );
  OAI22_X1 U2132 ( .A1(n1392), .A2(n1019), .B1(n1018), .B2(n1546), .ZN(n812)
         );
  OAI22_X1 U2133 ( .A1(n1020), .A2(n1392), .B1(n1019), .B2(n1547), .ZN(n813)
         );
  OAI22_X1 U2134 ( .A1(n1392), .A2(n1018), .B1(n1017), .B2(n1546), .ZN(n811)
         );
  OAI22_X1 U2135 ( .A1(n1393), .A2(n1023), .B1(n1022), .B2(n1546), .ZN(n816)
         );
  OAI22_X1 U2136 ( .A1(n24), .A2(n1011), .B1(n1010), .B2(n1547), .ZN(n804) );
  OAI22_X1 U2137 ( .A1(n1017), .A2(n24), .B1(n1016), .B2(n1546), .ZN(n810) );
  OAI22_X1 U2138 ( .A1(n24), .A2(n1327), .B1(n1015), .B2(n1547), .ZN(n809) );
  OAI22_X1 U2139 ( .A1(n1393), .A2(n1022), .B1(n1021), .B2(n1547), .ZN(n815)
         );
  INV_X1 U2140 ( .A(n1547), .ZN(n659) );
  XNOR2_X1 U2141 ( .A(n1516), .B(n65), .ZN(product[31]) );
  XNOR2_X1 U2142 ( .A(n1508), .B(n63), .ZN(product[33]) );
  XOR2_X1 U2143 ( .A(n117), .B(n66), .Z(product[30]) );
  INV_X1 U2144 ( .A(n101), .ZN(n264) );
  AOI21_X1 U2145 ( .B1(n106), .B2(n1537), .A(n103), .ZN(n101) );
  OAI21_X1 U2146 ( .B1(n1511), .B2(n115), .A(n116), .ZN(n114) );
  OAI22_X1 U2147 ( .A1(n1464), .A2(n1039), .B1(n1038), .B2(n1338), .ZN(n831)
         );
  OAI22_X1 U2148 ( .A1(n1262), .A2(n1031), .B1(n1030), .B2(n1271), .ZN(n823)
         );
  OAI22_X1 U2149 ( .A1(n1464), .A2(n1041), .B1(n1040), .B2(n1405), .ZN(n833)
         );
  OAI22_X1 U2150 ( .A1(n1464), .A2(n1032), .B1(n1031), .B2(n1338), .ZN(n824)
         );
  OAI22_X1 U2151 ( .A1(n1262), .A2(n1034), .B1(n1033), .B2(n1338), .ZN(n826)
         );
  OAI22_X1 U2152 ( .A1(n18), .A2(n1045), .B1(n1044), .B2(n1271), .ZN(n837) );
  OAI22_X1 U2153 ( .A1(n1464), .A2(n1038), .B1(n1037), .B2(n1405), .ZN(n830)
         );
  OAI22_X1 U2154 ( .A1(n1464), .A2(n1044), .B1(n1043), .B2(n1338), .ZN(n836)
         );
  OAI22_X1 U2155 ( .A1(n1262), .A2(n1028), .B1(n1027), .B2(n1271), .ZN(n424)
         );
  OAI22_X1 U2156 ( .A1(n1464), .A2(n1040), .B1(n1039), .B2(n1338), .ZN(n832)
         );
  OAI22_X1 U2157 ( .A1(n1463), .A2(n1033), .B1(n1032), .B2(n1271), .ZN(n825)
         );
  OAI22_X1 U2158 ( .A1(n1262), .A2(n1037), .B1(n1036), .B2(n1338), .ZN(n829)
         );
  OAI22_X1 U2159 ( .A1(n18), .A2(n1147), .B1(n1047), .B2(n1338), .ZN(n677) );
  OAI22_X1 U2160 ( .A1(n1027), .A2(n1463), .B1(n1027), .B2(n1338), .ZN(n661)
         );
  OAI22_X1 U2161 ( .A1(n1463), .A2(n1030), .B1(n1029), .B2(n1405), .ZN(n822)
         );
  OAI22_X1 U2162 ( .A1(n18), .A2(n1029), .B1(n1028), .B2(n1271), .ZN(n821) );
  OAI22_X1 U2163 ( .A1(n1463), .A2(n1036), .B1(n1035), .B2(n1338), .ZN(n828)
         );
  OAI22_X1 U2164 ( .A1(n1464), .A2(n1043), .B1(n1042), .B2(n1405), .ZN(n835)
         );
  OAI22_X1 U2165 ( .A1(n1464), .A2(n1042), .B1(n1041), .B2(n1338), .ZN(n834)
         );
  OAI22_X1 U2166 ( .A1(n1035), .A2(n1262), .B1(n1034), .B2(n1405), .ZN(n827)
         );
  OAI22_X1 U2167 ( .A1(n1262), .A2(n1046), .B1(n1045), .B2(n1271), .ZN(n838)
         );
  OAI21_X1 U2168 ( .B1(n1517), .B2(n107), .A(n108), .ZN(n106) );
endmodule


module mac_0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n34, n35, n36, n37, n38, n39, n40, n41, n43, n45, n46, n47,
         n48, n49, n51, n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65,
         n67, n69, n70, n71, n72, n73, n75, n77, n78, n79, n80, n81, n83, n85,
         n86, n87, n88, n89, n91, n93, n94, n95, n96, n97, n99, n101, n102,
         n103, n104, n105, n107, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n119, n121, n122, n124, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n184, n185, n187, n189, n191,
         n193, n195, n197, n199, n201, n203, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409;

  FA_X1 U3 ( .A(B[38]), .B(A[38]), .CI(n35), .CO(n34), .S(SUM[38]) );
  FA_X1 U7 ( .A(B[34]), .B(A[34]), .CI(n39), .CO(n38), .S(SUM[34]) );
  FA_X1 U9 ( .A(B[32]), .B(A[32]), .CI(n185), .CO(n40), .S(SUM[32]) );
  NAND2_X1 U254 ( .A1(B[36]), .A2(A[36]), .ZN(n381) );
  NAND2_X1 U255 ( .A1(B[8]), .A2(A[8]), .ZN(n148) );
  OR2_X1 U256 ( .A1(B[11]), .A2(A[11]), .ZN(n344) );
  OR2_X1 U257 ( .A1(B[0]), .A2(A[0]), .ZN(n345) );
  CLKBUF_X1 U258 ( .A(n40), .Z(n346) );
  CLKBUF_X1 U259 ( .A(n38), .Z(n347) );
  CLKBUF_X1 U260 ( .A(n376), .Z(n348) );
  CLKBUF_X1 U261 ( .A(n382), .Z(n349) );
  CLKBUF_X1 U262 ( .A(n150), .Z(n350) );
  CLKBUF_X1 U263 ( .A(n115), .Z(n351) );
  NAND3_X1 U264 ( .A1(n383), .A2(n382), .A3(n381), .ZN(n352) );
  NAND3_X1 U265 ( .A1(n375), .A2(n376), .A3(n377), .ZN(n353) );
  NAND3_X1 U266 ( .A1(n375), .A2(n348), .A3(n377), .ZN(n354) );
  AOI21_X1 U267 ( .B1(n350), .B2(n114), .A(n351), .ZN(n355) );
  AOI21_X1 U268 ( .B1(n150), .B2(n114), .A(n115), .ZN(n113) );
  CLKBUF_X1 U269 ( .A(n70), .Z(n356) );
  AOI21_X1 U270 ( .B1(n356), .B2(n407), .A(n67), .ZN(n357) );
  AOI21_X1 U271 ( .B1(n70), .B2(n407), .A(n67), .ZN(n65) );
  AOI21_X1 U272 ( .B1(n362), .B2(n130), .A(n131), .ZN(n358) );
  CLKBUF_X1 U273 ( .A(n173), .Z(n359) );
  NOR2_X1 U274 ( .A1(B[5]), .A2(A[5]), .ZN(n360) );
  NOR2_X1 U275 ( .A1(B[7]), .A2(A[7]), .ZN(n361) );
  CLKBUF_X1 U276 ( .A(n143), .Z(n362) );
  CLKBUF_X1 U277 ( .A(n110), .Z(n363) );
  AOI21_X1 U278 ( .B1(n363), .B2(n402), .A(n107), .ZN(n364) );
  CLKBUF_X1 U279 ( .A(n78), .Z(n365) );
  AOI21_X1 U280 ( .B1(n365), .B2(n405), .A(n75), .ZN(n366) );
  CLKBUF_X1 U281 ( .A(n102), .Z(n367) );
  XOR2_X1 U282 ( .A(B[33]), .B(A[33]), .Z(n368) );
  XOR2_X1 U283 ( .A(n346), .B(n368), .Z(SUM[33]) );
  NAND2_X1 U284 ( .A1(n40), .A2(B[33]), .ZN(n369) );
  NAND2_X1 U285 ( .A1(n40), .A2(A[33]), .ZN(n370) );
  NAND2_X1 U286 ( .A1(B[33]), .A2(A[33]), .ZN(n371) );
  NAND3_X1 U287 ( .A1(n369), .A2(n370), .A3(n371), .ZN(n39) );
  AOI21_X1 U288 ( .B1(n172), .B2(n180), .A(n359), .ZN(n372) );
  CLKBUF_X1 U289 ( .A(n86), .Z(n373) );
  NOR2_X2 U290 ( .A1(B[3]), .A2(A[3]), .ZN(n174) );
  XOR2_X1 U291 ( .A(B[35]), .B(A[35]), .Z(n374) );
  XOR2_X1 U292 ( .A(n347), .B(n374), .Z(SUM[35]) );
  NAND2_X1 U293 ( .A1(n38), .A2(B[35]), .ZN(n375) );
  NAND2_X1 U294 ( .A1(n38), .A2(A[35]), .ZN(n376) );
  NAND2_X1 U295 ( .A1(B[35]), .A2(A[35]), .ZN(n377) );
  NAND3_X1 U296 ( .A1(n375), .A2(n376), .A3(n377), .ZN(n37) );
  NOR2_X1 U297 ( .A1(B[11]), .A2(A[11]), .ZN(n378) );
  NAND3_X1 U298 ( .A1(n383), .A2(n349), .A3(n381), .ZN(n379) );
  NOR2_X1 U299 ( .A1(B[11]), .A2(A[11]), .ZN(n132) );
  XOR2_X1 U300 ( .A(B[36]), .B(A[36]), .Z(n380) );
  XOR2_X1 U301 ( .A(n380), .B(n354), .Z(SUM[36]) );
  NAND2_X1 U302 ( .A1(B[36]), .A2(n37), .ZN(n382) );
  NAND2_X1 U303 ( .A1(A[36]), .A2(n353), .ZN(n383) );
  NAND3_X1 U304 ( .A1(n383), .A2(n382), .A3(n381), .ZN(n36) );
  XOR2_X1 U305 ( .A(B[37]), .B(A[37]), .Z(n384) );
  XOR2_X1 U306 ( .A(n384), .B(n379), .Z(SUM[37]) );
  NAND2_X1 U307 ( .A1(B[37]), .A2(A[37]), .ZN(n385) );
  NAND2_X1 U308 ( .A1(B[37]), .A2(n352), .ZN(n386) );
  NAND2_X1 U309 ( .A1(A[37]), .A2(n36), .ZN(n387) );
  NAND3_X1 U310 ( .A1(n385), .A2(n386), .A3(n387), .ZN(n35) );
  CLKBUF_X1 U311 ( .A(n54), .Z(n388) );
  AOI21_X1 U312 ( .B1(n373), .B2(n400), .A(n83), .ZN(n389) );
  CLKBUF_X1 U313 ( .A(n62), .Z(n390) );
  CLKBUF_X1 U314 ( .A(n94), .Z(n391) );
  AOI21_X1 U315 ( .B1(n367), .B2(n403), .A(n99), .ZN(n392) );
  AOI21_X1 U316 ( .B1(n391), .B2(n401), .A(n91), .ZN(n393) );
  CLKBUF_X1 U317 ( .A(n46), .Z(n394) );
  AOI21_X1 U318 ( .B1(n388), .B2(n404), .A(n51), .ZN(n395) );
  AOI21_X1 U319 ( .B1(n390), .B2(n406), .A(n59), .ZN(n396) );
  NOR2_X2 U320 ( .A1(B[9]), .A2(A[9]), .ZN(n144) );
  INV_X1 U321 ( .A(n350), .ZN(n149) );
  OAI21_X1 U322 ( .B1(n149), .B2(n140), .A(n141), .ZN(n139) );
  INV_X1 U323 ( .A(n362), .ZN(n141) );
  INV_X1 U324 ( .A(n142), .ZN(n140) );
  NAND2_X1 U325 ( .A1(n142), .A2(n130), .ZN(n128) );
  AOI21_X1 U326 ( .B1(n170), .B2(n161), .A(n162), .ZN(n160) );
  INV_X1 U327 ( .A(n372), .ZN(n170) );
  INV_X1 U328 ( .A(n180), .ZN(n179) );
  INV_X1 U329 ( .A(n77), .ZN(n75) );
  INV_X1 U330 ( .A(n69), .ZN(n67) );
  AOI21_X1 U331 ( .B1(n86), .B2(n400), .A(n83), .ZN(n81) );
  INV_X1 U332 ( .A(n85), .ZN(n83) );
  AOI21_X1 U333 ( .B1(n62), .B2(n406), .A(n59), .ZN(n57) );
  INV_X1 U334 ( .A(n61), .ZN(n59) );
  AOI21_X1 U335 ( .B1(n54), .B2(n404), .A(n51), .ZN(n49) );
  INV_X1 U336 ( .A(n53), .ZN(n51) );
  NOR2_X1 U337 ( .A1(n128), .A2(n116), .ZN(n114) );
  NAND2_X1 U338 ( .A1(n398), .A2(n399), .ZN(n116) );
  OAI21_X1 U339 ( .B1(n163), .B2(n169), .A(n164), .ZN(n162) );
  AOI21_X1 U340 ( .B1(n172), .B2(n180), .A(n173), .ZN(n171) );
  AOI21_X1 U341 ( .B1(n94), .B2(n401), .A(n91), .ZN(n89) );
  INV_X1 U342 ( .A(n93), .ZN(n91) );
  AOI21_X1 U343 ( .B1(n110), .B2(n402), .A(n107), .ZN(n105) );
  INV_X1 U344 ( .A(n109), .ZN(n107) );
  AOI21_X1 U345 ( .B1(n102), .B2(n403), .A(n99), .ZN(n97) );
  INV_X1 U346 ( .A(n101), .ZN(n99) );
  OAI21_X1 U347 ( .B1(n144), .B2(n148), .A(n145), .ZN(n143) );
  NOR2_X1 U348 ( .A1(n168), .A2(n360), .ZN(n161) );
  OAI21_X1 U349 ( .B1(n181), .B2(n184), .A(n182), .ZN(n180) );
  NOR2_X1 U350 ( .A1(n137), .A2(n378), .ZN(n130) );
  NAND2_X1 U351 ( .A1(n199), .A2(n96), .ZN(n15) );
  INV_X1 U352 ( .A(n95), .ZN(n199) );
  NAND2_X1 U353 ( .A1(n201), .A2(n104), .ZN(n17) );
  INV_X1 U354 ( .A(n103), .ZN(n201) );
  NOR2_X1 U355 ( .A1(n147), .A2(n144), .ZN(n142) );
  OAI21_X1 U356 ( .B1(n171), .B2(n151), .A(n152), .ZN(n150) );
  NAND2_X1 U357 ( .A1(n161), .A2(n153), .ZN(n151) );
  AOI21_X1 U358 ( .B1(n153), .B2(n162), .A(n154), .ZN(n152) );
  NOR2_X1 U359 ( .A1(n158), .A2(n361), .ZN(n153) );
  AOI21_X1 U360 ( .B1(n143), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U361 ( .B1(n132), .B2(n138), .A(n133), .ZN(n131) );
  INV_X1 U362 ( .A(n126), .ZN(n124) );
  OAI21_X1 U363 ( .B1(n155), .B2(n159), .A(n156), .ZN(n154) );
  AOI21_X1 U364 ( .B1(n399), .B2(n124), .A(n119), .ZN(n117) );
  INV_X1 U365 ( .A(n121), .ZN(n119) );
  NAND2_X1 U366 ( .A1(n191), .A2(n64), .ZN(n7) );
  INV_X1 U367 ( .A(n63), .ZN(n191) );
  NAND2_X1 U368 ( .A1(n193), .A2(n72), .ZN(n9) );
  INV_X1 U369 ( .A(n71), .ZN(n193) );
  NAND2_X1 U370 ( .A1(n197), .A2(n88), .ZN(n13) );
  INV_X1 U371 ( .A(n87), .ZN(n197) );
  NAND2_X1 U372 ( .A1(n408), .A2(n45), .ZN(n2) );
  XOR2_X1 U373 ( .A(n395), .B(n3), .Z(SUM[30]) );
  NAND2_X1 U374 ( .A1(n187), .A2(n48), .ZN(n3) );
  INV_X1 U375 ( .A(n47), .ZN(n187) );
  NAND2_X1 U376 ( .A1(n404), .A2(n53), .ZN(n4) );
  XOR2_X1 U377 ( .A(n396), .B(n5), .Z(SUM[28]) );
  NAND2_X1 U378 ( .A1(n189), .A2(n56), .ZN(n5) );
  INV_X1 U379 ( .A(n55), .ZN(n189) );
  NAND2_X1 U380 ( .A1(n406), .A2(n61), .ZN(n6) );
  NAND2_X1 U381 ( .A1(n407), .A2(n69), .ZN(n8) );
  NAND2_X1 U382 ( .A1(n405), .A2(n77), .ZN(n10) );
  XOR2_X1 U383 ( .A(n389), .B(n11), .Z(SUM[22]) );
  NAND2_X1 U384 ( .A1(n195), .A2(n80), .ZN(n11) );
  INV_X1 U385 ( .A(n79), .ZN(n195) );
  NAND2_X1 U386 ( .A1(n400), .A2(n85), .ZN(n12) );
  XNOR2_X1 U387 ( .A(n391), .B(n14), .ZN(SUM[19]) );
  NAND2_X1 U388 ( .A1(n401), .A2(n93), .ZN(n14) );
  NAND2_X1 U389 ( .A1(n403), .A2(n101), .ZN(n16) );
  XOR2_X1 U390 ( .A(n122), .B(n20), .Z(SUM[13]) );
  NAND2_X1 U391 ( .A1(n399), .A2(n121), .ZN(n20) );
  AOI21_X1 U392 ( .B1(n127), .B2(n398), .A(n124), .ZN(n122) );
  XNOR2_X1 U393 ( .A(n127), .B(n21), .ZN(SUM[12]) );
  NAND2_X1 U394 ( .A1(n398), .A2(n126), .ZN(n21) );
  XOR2_X1 U395 ( .A(n134), .B(n22), .Z(SUM[11]) );
  NAND2_X1 U396 ( .A1(n344), .A2(n133), .ZN(n22) );
  AOI21_X1 U397 ( .B1(n139), .B2(n207), .A(n136), .ZN(n134) );
  XOR2_X1 U398 ( .A(n165), .B(n28), .Z(SUM[5]) );
  NAND2_X1 U399 ( .A1(n212), .A2(n164), .ZN(n28) );
  AOI21_X1 U400 ( .B1(n170), .B2(n213), .A(n167), .ZN(n165) );
  INV_X1 U401 ( .A(n137), .ZN(n207) );
  INV_X1 U402 ( .A(n168), .ZN(n213) );
  XOR2_X1 U403 ( .A(n149), .B(n25), .Z(SUM[8]) );
  NAND2_X1 U404 ( .A1(n209), .A2(n148), .ZN(n25) );
  INV_X1 U405 ( .A(n147), .ZN(n209) );
  XNOR2_X1 U406 ( .A(n146), .B(n24), .ZN(SUM[9]) );
  NAND2_X1 U407 ( .A1(n208), .A2(n145), .ZN(n24) );
  OAI21_X1 U408 ( .B1(n149), .B2(n147), .A(n148), .ZN(n146) );
  INV_X1 U409 ( .A(n138), .ZN(n136) );
  INV_X1 U410 ( .A(n169), .ZN(n167) );
  INV_X1 U411 ( .A(n144), .ZN(n208) );
  INV_X1 U412 ( .A(n361), .ZN(n210) );
  INV_X1 U413 ( .A(n360), .ZN(n212) );
  XOR2_X1 U414 ( .A(n160), .B(n27), .Z(SUM[6]) );
  NAND2_X1 U415 ( .A1(n211), .A2(n159), .ZN(n27) );
  INV_X1 U416 ( .A(n158), .ZN(n211) );
  XNOR2_X1 U417 ( .A(n170), .B(n29), .ZN(SUM[4]) );
  NAND2_X1 U418 ( .A1(n213), .A2(n169), .ZN(n29) );
  XNOR2_X1 U419 ( .A(n176), .B(n30), .ZN(SUM[3]) );
  NAND2_X1 U420 ( .A1(n214), .A2(n175), .ZN(n30) );
  OAI21_X1 U421 ( .B1(n179), .B2(n177), .A(n178), .ZN(n176) );
  XOR2_X1 U422 ( .A(n179), .B(n31), .Z(SUM[2]) );
  NAND2_X1 U423 ( .A1(n215), .A2(n178), .ZN(n31) );
  INV_X1 U424 ( .A(n177), .ZN(n215) );
  XOR2_X1 U425 ( .A(n32), .B(n184), .Z(SUM[1]) );
  NAND2_X1 U426 ( .A1(n216), .A2(n182), .ZN(n32) );
  INV_X1 U427 ( .A(n181), .ZN(n216) );
  AND2_X1 U428 ( .A1(n345), .A2(n184), .ZN(SUM[0]) );
  NAND2_X1 U429 ( .A1(n402), .A2(n109), .ZN(n18) );
  XOR2_X1 U430 ( .A(n355), .B(n19), .Z(SUM[14]) );
  NAND2_X1 U431 ( .A1(n203), .A2(n112), .ZN(n19) );
  INV_X1 U432 ( .A(n111), .ZN(n203) );
  XNOR2_X1 U433 ( .A(n139), .B(n23), .ZN(SUM[10]) );
  NAND2_X1 U434 ( .A1(n207), .A2(n138), .ZN(n23) );
  XNOR2_X1 U435 ( .A(n157), .B(n26), .ZN(SUM[7]) );
  NAND2_X1 U436 ( .A1(n210), .A2(n156), .ZN(n26) );
  OAI21_X1 U437 ( .B1(n160), .B2(n158), .A(n159), .ZN(n157) );
  NOR2_X1 U438 ( .A1(B[6]), .A2(A[6]), .ZN(n158) );
  NOR2_X1 U439 ( .A1(B[8]), .A2(A[8]), .ZN(n147) );
  NOR2_X1 U440 ( .A1(B[5]), .A2(A[5]), .ZN(n163) );
  NOR2_X1 U441 ( .A1(B[7]), .A2(A[7]), .ZN(n155) );
  OR2_X1 U442 ( .A1(B[12]), .A2(A[12]), .ZN(n398) );
  OR2_X1 U443 ( .A1(B[13]), .A2(A[13]), .ZN(n399) );
  NOR2_X1 U444 ( .A1(B[2]), .A2(A[2]), .ZN(n177) );
  NAND2_X1 U445 ( .A1(B[11]), .A2(A[11]), .ZN(n133) );
  NOR2_X1 U446 ( .A1(B[10]), .A2(A[10]), .ZN(n137) );
  NOR2_X1 U447 ( .A1(B[4]), .A2(A[4]), .ZN(n168) );
  NOR2_X1 U448 ( .A1(B[1]), .A2(A[1]), .ZN(n181) );
  NAND2_X1 U449 ( .A1(B[6]), .A2(A[6]), .ZN(n159) );
  NAND2_X1 U450 ( .A1(B[0]), .A2(A[0]), .ZN(n184) );
  NAND2_X1 U451 ( .A1(B[4]), .A2(A[4]), .ZN(n169) );
  NAND2_X1 U452 ( .A1(B[10]), .A2(A[10]), .ZN(n138) );
  NAND2_X1 U453 ( .A1(B[2]), .A2(A[2]), .ZN(n178) );
  NAND2_X1 U454 ( .A1(B[1]), .A2(A[1]), .ZN(n182) );
  NAND2_X1 U455 ( .A1(B[5]), .A2(A[5]), .ZN(n164) );
  NAND2_X1 U456 ( .A1(B[7]), .A2(A[7]), .ZN(n156) );
  NAND2_X1 U457 ( .A1(B[9]), .A2(A[9]), .ZN(n145) );
  INV_X1 U458 ( .A(n45), .ZN(n43) );
  NOR2_X1 U459 ( .A1(B[20]), .A2(A[20]), .ZN(n87) );
  NOR2_X1 U460 ( .A1(B[18]), .A2(A[18]), .ZN(n95) );
  NOR2_X1 U461 ( .A1(B[14]), .A2(A[14]), .ZN(n111) );
  NOR2_X1 U462 ( .A1(B[16]), .A2(A[16]), .ZN(n103) );
  NOR2_X1 U463 ( .A1(B[30]), .A2(A[30]), .ZN(n47) );
  NOR2_X1 U464 ( .A1(B[28]), .A2(A[28]), .ZN(n55) );
  NOR2_X1 U465 ( .A1(B[26]), .A2(A[26]), .ZN(n63) );
  NOR2_X1 U466 ( .A1(B[24]), .A2(A[24]), .ZN(n71) );
  NOR2_X1 U467 ( .A1(B[22]), .A2(A[22]), .ZN(n79) );
  OR2_X1 U468 ( .A1(B[21]), .A2(A[21]), .ZN(n400) );
  OR2_X1 U469 ( .A1(B[19]), .A2(A[19]), .ZN(n401) );
  OR2_X1 U470 ( .A1(B[15]), .A2(A[15]), .ZN(n402) );
  OR2_X1 U471 ( .A1(B[17]), .A2(A[17]), .ZN(n403) );
  OR2_X1 U472 ( .A1(B[29]), .A2(A[29]), .ZN(n404) );
  NAND2_X1 U473 ( .A1(B[21]), .A2(A[21]), .ZN(n85) );
  NAND2_X1 U474 ( .A1(B[12]), .A2(A[12]), .ZN(n126) );
  NAND2_X1 U475 ( .A1(B[19]), .A2(A[19]), .ZN(n93) );
  NAND2_X1 U476 ( .A1(B[13]), .A2(A[13]), .ZN(n121) );
  NAND2_X1 U477 ( .A1(B[15]), .A2(A[15]), .ZN(n109) );
  NAND2_X1 U478 ( .A1(B[17]), .A2(A[17]), .ZN(n101) );
  NAND2_X1 U479 ( .A1(B[23]), .A2(A[23]), .ZN(n77) );
  NAND2_X1 U480 ( .A1(B[25]), .A2(A[25]), .ZN(n69) );
  NAND2_X1 U481 ( .A1(B[27]), .A2(A[27]), .ZN(n61) );
  NAND2_X1 U482 ( .A1(B[29]), .A2(A[29]), .ZN(n53) );
  NAND2_X1 U483 ( .A1(B[31]), .A2(A[31]), .ZN(n45) );
  NAND2_X1 U484 ( .A1(B[20]), .A2(A[20]), .ZN(n88) );
  NAND2_X1 U485 ( .A1(B[18]), .A2(A[18]), .ZN(n96) );
  NAND2_X1 U486 ( .A1(B[14]), .A2(A[14]), .ZN(n112) );
  NAND2_X1 U487 ( .A1(B[16]), .A2(A[16]), .ZN(n104) );
  NAND2_X1 U488 ( .A1(B[30]), .A2(A[30]), .ZN(n48) );
  NAND2_X1 U489 ( .A1(B[28]), .A2(A[28]), .ZN(n56) );
  NAND2_X1 U490 ( .A1(B[26]), .A2(A[26]), .ZN(n64) );
  NAND2_X1 U491 ( .A1(B[24]), .A2(A[24]), .ZN(n72) );
  NAND2_X1 U492 ( .A1(B[22]), .A2(A[22]), .ZN(n80) );
  OR2_X1 U493 ( .A1(B[23]), .A2(A[23]), .ZN(n405) );
  OR2_X1 U494 ( .A1(B[27]), .A2(A[27]), .ZN(n406) );
  OR2_X1 U495 ( .A1(B[25]), .A2(A[25]), .ZN(n407) );
  OR2_X1 U496 ( .A1(B[31]), .A2(A[31]), .ZN(n408) );
  XNOR2_X1 U497 ( .A(n34), .B(n409), .ZN(SUM[39]) );
  XNOR2_X1 U498 ( .A(A[39]), .B(B[39]), .ZN(n409) );
  OAI21_X1 U499 ( .B1(n97), .B2(n95), .A(n96), .ZN(n94) );
  XOR2_X1 U500 ( .A(n392), .B(n15), .Z(SUM[18]) );
  XNOR2_X1 U501 ( .A(n373), .B(n12), .ZN(SUM[21]) );
  XNOR2_X1 U502 ( .A(n367), .B(n16), .ZN(SUM[17]) );
  XNOR2_X1 U503 ( .A(n394), .B(n2), .ZN(SUM[31]) );
  XOR2_X1 U504 ( .A(n364), .B(n17), .Z(SUM[16]) );
  INV_X1 U505 ( .A(n41), .ZN(n185) );
  OAI21_X1 U506 ( .B1(n105), .B2(n103), .A(n104), .ZN(n102) );
  AOI21_X1 U507 ( .B1(n46), .B2(n408), .A(n43), .ZN(n41) );
  OAI21_X1 U508 ( .B1(n49), .B2(n47), .A(n48), .ZN(n46) );
  XNOR2_X1 U509 ( .A(n365), .B(n10), .ZN(SUM[23]) );
  XNOR2_X1 U510 ( .A(n388), .B(n4), .ZN(SUM[29]) );
  XNOR2_X1 U511 ( .A(n363), .B(n18), .ZN(SUM[15]) );
  XOR2_X1 U512 ( .A(n393), .B(n13), .Z(SUM[20]) );
  AOI21_X1 U513 ( .B1(n78), .B2(n405), .A(n75), .ZN(n73) );
  OAI21_X1 U514 ( .B1(n89), .B2(n87), .A(n88), .ZN(n86) );
  OAI21_X1 U515 ( .B1(n113), .B2(n111), .A(n112), .ZN(n110) );
  OAI21_X1 U516 ( .B1(n81), .B2(n79), .A(n80), .ZN(n78) );
  OAI21_X1 U517 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  XNOR2_X1 U518 ( .A(n390), .B(n6), .ZN(SUM[27]) );
  XNOR2_X1 U519 ( .A(n356), .B(n8), .ZN(SUM[25]) );
  INV_X1 U520 ( .A(n174), .ZN(n214) );
  NOR2_X1 U521 ( .A1(n177), .A2(n174), .ZN(n172) );
  OAI21_X1 U522 ( .B1(n174), .B2(n178), .A(n175), .ZN(n173) );
  NAND2_X1 U523 ( .A1(B[3]), .A2(A[3]), .ZN(n175) );
  XOR2_X1 U524 ( .A(n357), .B(n7), .Z(SUM[26]) );
  XOR2_X1 U525 ( .A(n366), .B(n9), .Z(SUM[24]) );
  OAI21_X1 U526 ( .B1(n149), .B2(n128), .A(n358), .ZN(n127) );
  OAI21_X1 U527 ( .B1(n65), .B2(n63), .A(n64), .ZN(n62) );
  OAI21_X1 U528 ( .B1(n73), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U529 ( .B1(n129), .B2(n116), .A(n117), .ZN(n115) );
endmodule


module mac_0 ( clk, clear_acc, a, b, mac_out );
  input [19:0] a;
  input [19:0] b;
  output [39:0] mac_out;
  input clk, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, n2, n3;
  wire   [39:0] mul;
  wire   [39:0] pipeline;
  wire   [39:0] sum;

  DFF_X1 \pipeline_reg[37]  ( .D(mul[37]), .CK(clk), .Q(pipeline[37]) );
  DFF_X1 \pipeline_reg[36]  ( .D(mul[36]), .CK(clk), .Q(pipeline[36]) );
  DFF_X1 \pipeline_reg[35]  ( .D(mul[35]), .CK(clk), .Q(pipeline[35]) );
  DFF_X1 \pipeline_reg[34]  ( .D(mul[34]), .CK(clk), .Q(pipeline[34]) );
  DFF_X1 \pipeline_reg[33]  ( .D(mul[33]), .CK(clk), .Q(pipeline[33]) );
  DFF_X1 \pipeline_reg[32]  ( .D(mul[32]), .CK(clk), .Q(pipeline[32]) );
  DFF_X1 \pipeline_reg[31]  ( .D(mul[31]), .CK(clk), .Q(pipeline[31]) );
  DFF_X1 \pipeline_reg[30]  ( .D(mul[30]), .CK(clk), .Q(pipeline[30]) );
  DFF_X1 \pipeline_reg[29]  ( .D(mul[29]), .CK(clk), .Q(pipeline[29]) );
  DFF_X1 \pipeline_reg[28]  ( .D(mul[28]), .CK(clk), .Q(pipeline[28]) );
  DFF_X1 \pipeline_reg[27]  ( .D(mul[27]), .CK(clk), .Q(pipeline[27]) );
  DFF_X1 \pipeline_reg[26]  ( .D(mul[26]), .CK(clk), .Q(pipeline[26]) );
  DFF_X1 \pipeline_reg[25]  ( .D(mul[25]), .CK(clk), .Q(pipeline[25]) );
  DFF_X1 \pipeline_reg[24]  ( .D(mul[24]), .CK(clk), .Q(pipeline[24]) );
  DFF_X1 \pipeline_reg[23]  ( .D(mul[23]), .CK(clk), .Q(pipeline[23]) );
  DFF_X1 \pipeline_reg[22]  ( .D(mul[22]), .CK(clk), .Q(pipeline[22]) );
  DFF_X1 \pipeline_reg[21]  ( .D(mul[21]), .CK(clk), .Q(pipeline[21]) );
  DFF_X1 \pipeline_reg[20]  ( .D(mul[20]), .CK(clk), .Q(pipeline[20]) );
  DFF_X1 \pipeline_reg[19]  ( .D(mul[19]), .CK(clk), .Q(pipeline[19]) );
  DFF_X1 \pipeline_reg[18]  ( .D(mul[18]), .CK(clk), .Q(pipeline[18]) );
  DFF_X1 \pipeline_reg[17]  ( .D(mul[17]), .CK(clk), .Q(pipeline[17]) );
  DFF_X1 \pipeline_reg[16]  ( .D(mul[16]), .CK(clk), .Q(pipeline[16]) );
  DFF_X1 \pipeline_reg[15]  ( .D(mul[15]), .CK(clk), .Q(pipeline[15]) );
  DFF_X1 \pipeline_reg[14]  ( .D(mul[14]), .CK(clk), .Q(pipeline[14]) );
  DFF_X1 \pipeline_reg[13]  ( .D(mul[13]), .CK(clk), .Q(pipeline[13]) );
  DFF_X1 \pipeline_reg[12]  ( .D(mul[12]), .CK(clk), .Q(pipeline[12]) );
  DFF_X1 \pipeline_reg[11]  ( .D(mul[11]), .CK(clk), .Q(pipeline[11]) );
  DFF_X1 \pipeline_reg[10]  ( .D(mul[10]), .CK(clk), .Q(pipeline[10]) );
  DFF_X1 \pipeline_reg[9]  ( .D(mul[9]), .CK(clk), .Q(pipeline[9]) );
  DFF_X1 \pipeline_reg[8]  ( .D(mul[8]), .CK(clk), .Q(pipeline[8]) );
  DFF_X1 \pipeline_reg[7]  ( .D(mul[7]), .CK(clk), .Q(pipeline[7]) );
  DFF_X1 \pipeline_reg[6]  ( .D(mul[6]), .CK(clk), .Q(pipeline[6]) );
  DFF_X1 \pipeline_reg[5]  ( .D(mul[5]), .CK(clk), .Q(pipeline[5]) );
  DFF_X1 \pipeline_reg[4]  ( .D(mul[4]), .CK(clk), .Q(pipeline[4]) );
  DFF_X1 \pipeline_reg[3]  ( .D(mul[3]), .CK(clk), .Q(pipeline[3]) );
  DFF_X1 \pipeline_reg[2]  ( .D(mul[2]), .CK(clk), .Q(pipeline[2]) );
  DFF_X1 \pipeline_reg[1]  ( .D(mul[1]), .CK(clk), .Q(pipeline[1]) );
  DFF_X1 \pipeline_reg[0]  ( .D(mul[0]), .CK(clk), .Q(pipeline[0]) );
  DFF_X1 \mac_out_reg[0]  ( .D(N3), .CK(clk), .Q(mac_out[0]) );
  DFF_X1 \mac_out_reg[1]  ( .D(N4), .CK(clk), .Q(mac_out[1]) );
  DFF_X1 \mac_out_reg[2]  ( .D(N5), .CK(clk), .Q(mac_out[2]) );
  DFF_X1 \mac_out_reg[3]  ( .D(N6), .CK(clk), .Q(mac_out[3]) );
  DFF_X1 \mac_out_reg[4]  ( .D(N7), .CK(clk), .Q(mac_out[4]) );
  DFF_X1 \mac_out_reg[5]  ( .D(N8), .CK(clk), .Q(mac_out[5]) );
  DFF_X1 \mac_out_reg[6]  ( .D(N9), .CK(clk), .Q(mac_out[6]) );
  DFF_X1 \mac_out_reg[7]  ( .D(N10), .CK(clk), .Q(mac_out[7]) );
  DFF_X1 \mac_out_reg[8]  ( .D(N11), .CK(clk), .Q(mac_out[8]) );
  DFF_X1 \mac_out_reg[9]  ( .D(N12), .CK(clk), .Q(mac_out[9]) );
  DFF_X1 \mac_out_reg[10]  ( .D(N13), .CK(clk), .Q(mac_out[10]) );
  DFF_X1 \mac_out_reg[11]  ( .D(N14), .CK(clk), .Q(mac_out[11]) );
  DFF_X1 \mac_out_reg[12]  ( .D(N15), .CK(clk), .Q(mac_out[12]) );
  DFF_X1 \mac_out_reg[13]  ( .D(N16), .CK(clk), .Q(mac_out[13]) );
  DFF_X1 \mac_out_reg[14]  ( .D(N17), .CK(clk), .Q(mac_out[14]) );
  DFF_X1 \mac_out_reg[15]  ( .D(N18), .CK(clk), .Q(mac_out[15]) );
  DFF_X1 \mac_out_reg[16]  ( .D(N19), .CK(clk), .Q(mac_out[16]) );
  DFF_X1 \mac_out_reg[17]  ( .D(N20), .CK(clk), .Q(mac_out[17]) );
  DFF_X1 \mac_out_reg[18]  ( .D(N21), .CK(clk), .Q(mac_out[18]) );
  DFF_X1 \mac_out_reg[19]  ( .D(N22), .CK(clk), .Q(mac_out[19]) );
  DFF_X1 \mac_out_reg[20]  ( .D(N23), .CK(clk), .Q(mac_out[20]) );
  DFF_X1 \mac_out_reg[21]  ( .D(N24), .CK(clk), .Q(mac_out[21]) );
  DFF_X1 \mac_out_reg[22]  ( .D(N25), .CK(clk), .Q(mac_out[22]) );
  DFF_X1 \mac_out_reg[23]  ( .D(N26), .CK(clk), .Q(mac_out[23]) );
  DFF_X1 \mac_out_reg[24]  ( .D(N27), .CK(clk), .Q(mac_out[24]) );
  DFF_X1 \mac_out_reg[25]  ( .D(N28), .CK(clk), .Q(mac_out[25]) );
  DFF_X1 \mac_out_reg[26]  ( .D(N29), .CK(clk), .Q(mac_out[26]) );
  DFF_X1 \mac_out_reg[27]  ( .D(N30), .CK(clk), .Q(mac_out[27]) );
  DFF_X1 \mac_out_reg[28]  ( .D(N31), .CK(clk), .Q(mac_out[28]) );
  DFF_X1 \mac_out_reg[29]  ( .D(N32), .CK(clk), .Q(mac_out[29]) );
  DFF_X1 \mac_out_reg[30]  ( .D(N33), .CK(clk), .Q(mac_out[30]) );
  DFF_X1 \mac_out_reg[31]  ( .D(N34), .CK(clk), .Q(mac_out[31]) );
  DFF_X1 \mac_out_reg[32]  ( .D(N35), .CK(clk), .Q(mac_out[32]) );
  DFF_X1 \mac_out_reg[33]  ( .D(N36), .CK(clk), .Q(mac_out[33]) );
  DFF_X1 \mac_out_reg[34]  ( .D(N37), .CK(clk), .Q(mac_out[34]) );
  DFF_X1 \mac_out_reg[35]  ( .D(N38), .CK(clk), .Q(mac_out[35]) );
  DFF_X1 \mac_out_reg[36]  ( .D(N39), .CK(clk), .Q(mac_out[36]) );
  DFF_X1 \mac_out_reg[37]  ( .D(N40), .CK(clk), .Q(mac_out[37]) );
  DFF_X1 \mac_out_reg[38]  ( .D(N41), .CK(clk), .Q(mac_out[38]) );
  DFF_X1 \mac_out_reg[39]  ( .D(N42), .CK(clk), .Q(mac_out[39]) );
  mac_0_DW_mult_tc_1 mult_355 ( .a(a), .b(b), .product(mul) );
  mac_0_DW01_add_1 add_356 ( .A(pipeline), .B(mac_out), .CI(1'b0), .SUM(sum)
         );
  DFF_X1 \pipeline_reg[38]  ( .D(mul[38]), .CK(clk), .Q(pipeline[38]) );
  DFF_X1 \pipeline_reg[39]  ( .D(mul[39]), .CK(clk), .Q(pipeline[39]) );
  BUF_X1 U3 ( .A(n3), .Z(n2) );
  INV_X1 U4 ( .A(clear_acc), .ZN(n3) );
  AND2_X1 U6 ( .A1(sum[39]), .A2(n2), .ZN(N42) );
  AND2_X1 U7 ( .A1(sum[38]), .A2(n2), .ZN(N41) );
  AND2_X1 U8 ( .A1(sum[37]), .A2(n2), .ZN(N40) );
  AND2_X1 U9 ( .A1(sum[36]), .A2(n2), .ZN(N39) );
  AND2_X1 U10 ( .A1(sum[35]), .A2(n2), .ZN(N38) );
  AND2_X1 U11 ( .A1(sum[34]), .A2(n2), .ZN(N37) );
  AND2_X1 U12 ( .A1(sum[33]), .A2(n2), .ZN(N36) );
  AND2_X1 U13 ( .A1(sum[32]), .A2(n2), .ZN(N35) );
  AND2_X1 U14 ( .A1(sum[31]), .A2(n2), .ZN(N34) );
  AND2_X1 U15 ( .A1(sum[30]), .A2(n2), .ZN(N33) );
  AND2_X1 U16 ( .A1(sum[29]), .A2(n2), .ZN(N32) );
  AND2_X1 U17 ( .A1(sum[28]), .A2(n3), .ZN(N31) );
  AND2_X1 U18 ( .A1(sum[27]), .A2(n3), .ZN(N30) );
  AND2_X1 U19 ( .A1(sum[26]), .A2(n3), .ZN(N29) );
  AND2_X1 U20 ( .A1(sum[25]), .A2(n3), .ZN(N28) );
  AND2_X1 U21 ( .A1(sum[24]), .A2(n3), .ZN(N27) );
  AND2_X1 U22 ( .A1(sum[23]), .A2(n3), .ZN(N26) );
  AND2_X1 U23 ( .A1(sum[22]), .A2(n3), .ZN(N25) );
  AND2_X1 U24 ( .A1(sum[21]), .A2(n3), .ZN(N24) );
  AND2_X1 U25 ( .A1(sum[20]), .A2(n3), .ZN(N23) );
  AND2_X1 U26 ( .A1(sum[19]), .A2(n3), .ZN(N22) );
  AND2_X1 U27 ( .A1(sum[18]), .A2(n3), .ZN(N21) );
  AND2_X1 U28 ( .A1(sum[17]), .A2(n3), .ZN(N20) );
  AND2_X1 U29 ( .A1(sum[16]), .A2(n3), .ZN(N19) );
  AND2_X1 U30 ( .A1(sum[15]), .A2(n3), .ZN(N18) );
  AND2_X1 U31 ( .A1(sum[14]), .A2(n3), .ZN(N17) );
  AND2_X1 U32 ( .A1(sum[13]), .A2(n3), .ZN(N16) );
  AND2_X1 U33 ( .A1(sum[12]), .A2(n3), .ZN(N15) );
  AND2_X1 U34 ( .A1(sum[11]), .A2(n3), .ZN(N14) );
  AND2_X1 U35 ( .A1(sum[10]), .A2(n3), .ZN(N13) );
  AND2_X1 U36 ( .A1(sum[9]), .A2(n3), .ZN(N12) );
  AND2_X1 U37 ( .A1(sum[8]), .A2(n3), .ZN(N11) );
  AND2_X1 U38 ( .A1(sum[7]), .A2(n3), .ZN(N10) );
  AND2_X1 U39 ( .A1(sum[6]), .A2(n3), .ZN(N9) );
  AND2_X1 U40 ( .A1(sum[5]), .A2(n3), .ZN(N8) );
  AND2_X1 U41 ( .A1(sum[4]), .A2(n3), .ZN(N7) );
  AND2_X1 U42 ( .A1(sum[3]), .A2(n3), .ZN(N6) );
  AND2_X1 U43 ( .A1(sum[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U44 ( .A1(sum[1]), .A2(n3), .ZN(N4) );
  AND2_X1 U45 ( .A1(sum[0]), .A2(n2), .ZN(N3) );
endmodule


module memory_WIDTH40_SIZE1_LOGSIZE4_7 ( clk, data_in, data_out, addr, wr_en
 );
  input [39:0] data_in;
  output [39:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   \mem[0][39] , \mem[0][38] , \mem[0][37] , \mem[0][36] , \mem[0][35] ,
         \mem[0][34] , \mem[0][33] , \mem[0][32] , \mem[0][31] , \mem[0][30] ,
         \mem[0][29] , \mem[0][28] , \mem[0][27] , \mem[0][26] , \mem[0][25] ,
         \mem[0][24] , \mem[0][23] , \mem[0][22] , \mem[0][21] , \mem[0][20] ,
         \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] , \mem[0][15] ,
         \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] ,
         \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , n43,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n85, n86;

  DFF_X1 \mem_reg[0][39]  ( .D(n5), .CK(clk), .Q(\mem[0][39] ) );
  DFF_X1 \mem_reg[0][38]  ( .D(n6), .CK(clk), .Q(\mem[0][38] ) );
  DFF_X1 \mem_reg[0][37]  ( .D(n7), .CK(clk), .Q(\mem[0][37] ) );
  DFF_X1 \mem_reg[0][36]  ( .D(n8), .CK(clk), .Q(\mem[0][36] ) );
  DFF_X1 \mem_reg[0][35]  ( .D(n9), .CK(clk), .Q(\mem[0][35] ) );
  DFF_X1 \mem_reg[0][34]  ( .D(n10), .CK(clk), .Q(\mem[0][34] ) );
  DFF_X1 \mem_reg[0][33]  ( .D(n11), .CK(clk), .Q(\mem[0][33] ) );
  DFF_X1 \mem_reg[0][32]  ( .D(n12), .CK(clk), .Q(\mem[0][32] ) );
  DFF_X1 \mem_reg[0][31]  ( .D(n13), .CK(clk), .Q(\mem[0][31] ) );
  DFF_X1 \mem_reg[0][30]  ( .D(n14), .CK(clk), .Q(\mem[0][30] ) );
  DFF_X1 \mem_reg[0][29]  ( .D(n15), .CK(clk), .Q(\mem[0][29] ) );
  DFF_X1 \mem_reg[0][28]  ( .D(n16), .CK(clk), .Q(\mem[0][28] ) );
  DFF_X1 \mem_reg[0][27]  ( .D(n17), .CK(clk), .Q(\mem[0][27] ) );
  DFF_X1 \mem_reg[0][26]  ( .D(n18), .CK(clk), .Q(\mem[0][26] ) );
  DFF_X1 \mem_reg[0][25]  ( .D(n19), .CK(clk), .Q(\mem[0][25] ) );
  DFF_X1 \mem_reg[0][24]  ( .D(n20), .CK(clk), .Q(\mem[0][24] ) );
  DFF_X1 \mem_reg[0][23]  ( .D(n21), .CK(clk), .Q(\mem[0][23] ) );
  DFF_X1 \mem_reg[0][22]  ( .D(n22), .CK(clk), .Q(\mem[0][22] ) );
  DFF_X1 \mem_reg[0][21]  ( .D(n23), .CK(clk), .Q(\mem[0][21] ) );
  DFF_X1 \mem_reg[0][20]  ( .D(n24), .CK(clk), .Q(\mem[0][20] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n25), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n26), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n27), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n28), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n29), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n30), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n31), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n32), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n33), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n34), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n35), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n36), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n37), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n38), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n39), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n40), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n41), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n42), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n44), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n85), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[39]  ( .D(\mem[0][39] ), .CK(clk), .Q(data_out[39]) );
  DFF_X1 \data_out_reg[38]  ( .D(\mem[0][38] ), .CK(clk), .Q(data_out[38]) );
  DFF_X1 \data_out_reg[37]  ( .D(\mem[0][37] ), .CK(clk), .Q(data_out[37]) );
  DFF_X1 \data_out_reg[36]  ( .D(\mem[0][36] ), .CK(clk), .Q(data_out[36]) );
  DFF_X1 \data_out_reg[35]  ( .D(\mem[0][35] ), .CK(clk), .Q(data_out[35]) );
  DFF_X1 \data_out_reg[34]  ( .D(\mem[0][34] ), .CK(clk), .Q(data_out[34]) );
  DFF_X1 \data_out_reg[33]  ( .D(\mem[0][33] ), .CK(clk), .Q(data_out[33]) );
  DFF_X1 \data_out_reg[32]  ( .D(\mem[0][32] ), .CK(clk), .Q(data_out[32]) );
  DFF_X1 \data_out_reg[31]  ( .D(\mem[0][31] ), .CK(clk), .Q(data_out[31]) );
  DFF_X1 \data_out_reg[30]  ( .D(\mem[0][30] ), .CK(clk), .Q(data_out[30]) );
  DFF_X1 \data_out_reg[29]  ( .D(\mem[0][29] ), .CK(clk), .Q(data_out[29]) );
  DFF_X1 \data_out_reg[28]  ( .D(\mem[0][28] ), .CK(clk), .Q(data_out[28]) );
  DFF_X1 \data_out_reg[27]  ( .D(\mem[0][27] ), .CK(clk), .Q(data_out[27]) );
  DFF_X1 \data_out_reg[26]  ( .D(\mem[0][26] ), .CK(clk), .Q(data_out[26]) );
  DFF_X1 \data_out_reg[25]  ( .D(\mem[0][25] ), .CK(clk), .Q(data_out[25]) );
  DFF_X1 \data_out_reg[24]  ( .D(\mem[0][24] ), .CK(clk), .Q(data_out[24]) );
  DFF_X1 \data_out_reg[23]  ( .D(\mem[0][23] ), .CK(clk), .Q(data_out[23]) );
  DFF_X1 \data_out_reg[22]  ( .D(\mem[0][22] ), .CK(clk), .Q(data_out[22]) );
  DFF_X1 \data_out_reg[21]  ( .D(\mem[0][21] ), .CK(clk), .Q(data_out[21]) );
  DFF_X1 \data_out_reg[20]  ( .D(\mem[0][20] ), .CK(clk), .Q(data_out[20]) );
  DFF_X1 \data_out_reg[19]  ( .D(\mem[0][19] ), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(\mem[0][18] ), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[17]  ( .D(\mem[0][17] ), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \data_out_reg[16]  ( .D(\mem[0][16] ), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  AND3_X1 U3 ( .A1(wr_en), .A2(n86), .A3(n84), .ZN(n1) );
  INV_X1 U4 ( .A(n1), .ZN(n3) );
  INV_X1 U5 ( .A(n1), .ZN(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n4) );
  INV_X1 U7 ( .A(addr[0]), .ZN(n86) );
  NOR3_X1 U8 ( .A1(addr[1]), .A2(addr[3]), .A3(addr[2]), .ZN(n84) );
  INV_X1 U9 ( .A(n43), .ZN(n85) );
  AOI22_X1 U10 ( .A1(\mem[0][0] ), .A2(n3), .B1(data_in[0]), .B2(n4), .ZN(n43)
         );
  INV_X1 U11 ( .A(n45), .ZN(n44) );
  AOI22_X1 U12 ( .A1(\mem[0][1] ), .A2(n2), .B1(data_in[1]), .B2(n4), .ZN(n45)
         );
  INV_X1 U13 ( .A(n46), .ZN(n42) );
  AOI22_X1 U14 ( .A1(\mem[0][2] ), .A2(n2), .B1(data_in[2]), .B2(n1), .ZN(n46)
         );
  INV_X1 U15 ( .A(n47), .ZN(n41) );
  AOI22_X1 U16 ( .A1(\mem[0][3] ), .A2(n3), .B1(data_in[3]), .B2(n4), .ZN(n47)
         );
  INV_X1 U17 ( .A(n48), .ZN(n40) );
  AOI22_X1 U18 ( .A1(\mem[0][4] ), .A2(n3), .B1(data_in[4]), .B2(n1), .ZN(n48)
         );
  INV_X1 U19 ( .A(n49), .ZN(n39) );
  AOI22_X1 U20 ( .A1(\mem[0][5] ), .A2(n3), .B1(data_in[5]), .B2(n1), .ZN(n49)
         );
  INV_X1 U21 ( .A(n50), .ZN(n38) );
  AOI22_X1 U22 ( .A1(\mem[0][6] ), .A2(n3), .B1(data_in[6]), .B2(n4), .ZN(n50)
         );
  INV_X1 U23 ( .A(n51), .ZN(n37) );
  AOI22_X1 U24 ( .A1(\mem[0][7] ), .A2(n3), .B1(data_in[7]), .B2(n1), .ZN(n51)
         );
  INV_X1 U25 ( .A(n52), .ZN(n36) );
  AOI22_X1 U26 ( .A1(\mem[0][8] ), .A2(n3), .B1(data_in[8]), .B2(n1), .ZN(n52)
         );
  INV_X1 U27 ( .A(n53), .ZN(n35) );
  AOI22_X1 U28 ( .A1(\mem[0][9] ), .A2(n3), .B1(data_in[9]), .B2(n1), .ZN(n53)
         );
  INV_X1 U29 ( .A(n54), .ZN(n34) );
  AOI22_X1 U30 ( .A1(\mem[0][10] ), .A2(n3), .B1(data_in[10]), .B2(n4), .ZN(
        n54) );
  INV_X1 U31 ( .A(n55), .ZN(n33) );
  AOI22_X1 U32 ( .A1(\mem[0][11] ), .A2(n3), .B1(data_in[11]), .B2(n1), .ZN(
        n55) );
  INV_X1 U33 ( .A(n56), .ZN(n32) );
  AOI22_X1 U34 ( .A1(\mem[0][12] ), .A2(n3), .B1(data_in[12]), .B2(n4), .ZN(
        n56) );
  INV_X1 U35 ( .A(n57), .ZN(n31) );
  AOI22_X1 U36 ( .A1(\mem[0][13] ), .A2(n3), .B1(data_in[13]), .B2(n4), .ZN(
        n57) );
  INV_X1 U37 ( .A(n58), .ZN(n30) );
  AOI22_X1 U38 ( .A1(\mem[0][14] ), .A2(n3), .B1(data_in[14]), .B2(n4), .ZN(
        n58) );
  INV_X1 U39 ( .A(n59), .ZN(n29) );
  AOI22_X1 U40 ( .A1(\mem[0][15] ), .A2(n3), .B1(data_in[15]), .B2(n4), .ZN(
        n59) );
  INV_X1 U41 ( .A(n60), .ZN(n28) );
  AOI22_X1 U42 ( .A1(\mem[0][16] ), .A2(n2), .B1(data_in[16]), .B2(n1), .ZN(
        n60) );
  INV_X1 U43 ( .A(n61), .ZN(n27) );
  AOI22_X1 U44 ( .A1(\mem[0][17] ), .A2(n2), .B1(data_in[17]), .B2(n1), .ZN(
        n61) );
  INV_X1 U45 ( .A(n62), .ZN(n26) );
  AOI22_X1 U46 ( .A1(\mem[0][18] ), .A2(n2), .B1(data_in[18]), .B2(n1), .ZN(
        n62) );
  INV_X1 U47 ( .A(n63), .ZN(n25) );
  AOI22_X1 U48 ( .A1(\mem[0][19] ), .A2(n2), .B1(data_in[19]), .B2(n1), .ZN(
        n63) );
  INV_X1 U49 ( .A(n64), .ZN(n24) );
  AOI22_X1 U50 ( .A1(\mem[0][20] ), .A2(n2), .B1(data_in[20]), .B2(n4), .ZN(
        n64) );
  INV_X1 U51 ( .A(n65), .ZN(n23) );
  AOI22_X1 U52 ( .A1(\mem[0][21] ), .A2(n2), .B1(data_in[21]), .B2(n1), .ZN(
        n65) );
  INV_X1 U53 ( .A(n66), .ZN(n22) );
  AOI22_X1 U54 ( .A1(\mem[0][22] ), .A2(n2), .B1(data_in[22]), .B2(n4), .ZN(
        n66) );
  INV_X1 U55 ( .A(n67), .ZN(n21) );
  AOI22_X1 U56 ( .A1(\mem[0][23] ), .A2(n2), .B1(data_in[23]), .B2(n1), .ZN(
        n67) );
  INV_X1 U57 ( .A(n68), .ZN(n20) );
  AOI22_X1 U58 ( .A1(\mem[0][24] ), .A2(n2), .B1(data_in[24]), .B2(n1), .ZN(
        n68) );
  INV_X1 U59 ( .A(n69), .ZN(n19) );
  AOI22_X1 U60 ( .A1(\mem[0][25] ), .A2(n2), .B1(data_in[25]), .B2(n4), .ZN(
        n69) );
  INV_X1 U61 ( .A(n70), .ZN(n18) );
  AOI22_X1 U62 ( .A1(\mem[0][26] ), .A2(n2), .B1(data_in[26]), .B2(n1), .ZN(
        n70) );
  INV_X1 U63 ( .A(n71), .ZN(n17) );
  AOI22_X1 U64 ( .A1(\mem[0][27] ), .A2(n2), .B1(data_in[27]), .B2(n1), .ZN(
        n71) );
  INV_X1 U65 ( .A(n72), .ZN(n16) );
  AOI22_X1 U66 ( .A1(\mem[0][28] ), .A2(n3), .B1(data_in[28]), .B2(n1), .ZN(
        n72) );
  INV_X1 U67 ( .A(n73), .ZN(n15) );
  AOI22_X1 U68 ( .A1(\mem[0][29] ), .A2(n2), .B1(data_in[29]), .B2(n4), .ZN(
        n73) );
  INV_X1 U69 ( .A(n74), .ZN(n14) );
  AOI22_X1 U70 ( .A1(\mem[0][30] ), .A2(n3), .B1(data_in[30]), .B2(n4), .ZN(
        n74) );
  INV_X1 U71 ( .A(n75), .ZN(n13) );
  AOI22_X1 U72 ( .A1(\mem[0][31] ), .A2(n2), .B1(data_in[31]), .B2(n1), .ZN(
        n75) );
  INV_X1 U73 ( .A(n76), .ZN(n12) );
  AOI22_X1 U74 ( .A1(\mem[0][32] ), .A2(n3), .B1(data_in[32]), .B2(n1), .ZN(
        n76) );
  INV_X1 U75 ( .A(n77), .ZN(n11) );
  AOI22_X1 U76 ( .A1(\mem[0][33] ), .A2(n2), .B1(data_in[33]), .B2(n4), .ZN(
        n77) );
  INV_X1 U77 ( .A(n78), .ZN(n10) );
  AOI22_X1 U78 ( .A1(\mem[0][34] ), .A2(n3), .B1(data_in[34]), .B2(n1), .ZN(
        n78) );
  INV_X1 U79 ( .A(n79), .ZN(n9) );
  AOI22_X1 U80 ( .A1(\mem[0][35] ), .A2(n2), .B1(data_in[35]), .B2(n1), .ZN(
        n79) );
  INV_X1 U81 ( .A(n80), .ZN(n8) );
  AOI22_X1 U82 ( .A1(\mem[0][36] ), .A2(n3), .B1(data_in[36]), .B2(n4), .ZN(
        n80) );
  INV_X1 U83 ( .A(n81), .ZN(n7) );
  AOI22_X1 U84 ( .A1(\mem[0][37] ), .A2(n2), .B1(data_in[37]), .B2(n4), .ZN(
        n81) );
  INV_X1 U85 ( .A(n82), .ZN(n6) );
  AOI22_X1 U86 ( .A1(\mem[0][38] ), .A2(n3), .B1(data_in[38]), .B2(n1), .ZN(
        n82) );
  INV_X1 U87 ( .A(n83), .ZN(n5) );
  AOI22_X1 U88 ( .A1(\mem[0][39] ), .A2(n2), .B1(data_in[39]), .B2(n1), .ZN(
        n83) );
endmodule


module memory_WIDTH40_SIZE1_LOGSIZE4_6 ( clk, data_in, data_out, addr, wr_en
 );
  input [39:0] data_in;
  output [39:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   \mem[0][39] , \mem[0][38] , \mem[0][37] , \mem[0][36] , \mem[0][35] ,
         \mem[0][34] , \mem[0][33] , \mem[0][32] , \mem[0][31] , \mem[0][30] ,
         \mem[0][29] , \mem[0][28] , \mem[0][27] , \mem[0][26] , \mem[0][25] ,
         \mem[0][24] , \mem[0][23] , \mem[0][22] , \mem[0][21] , \mem[0][20] ,
         \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] , \mem[0][15] ,
         \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] ,
         \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  DFF_X1 \mem_reg[0][39]  ( .D(n5), .CK(clk), .Q(\mem[0][39] ) );
  DFF_X1 \data_out_reg[39]  ( .D(\mem[0][39] ), .CK(clk), .Q(data_out[39]) );
  DFF_X1 \mem_reg[0][38]  ( .D(n6), .CK(clk), .Q(\mem[0][38] ) );
  DFF_X1 \data_out_reg[38]  ( .D(\mem[0][38] ), .CK(clk), .Q(data_out[38]) );
  DFF_X1 \mem_reg[0][37]  ( .D(n7), .CK(clk), .Q(\mem[0][37] ) );
  DFF_X1 \data_out_reg[37]  ( .D(\mem[0][37] ), .CK(clk), .Q(data_out[37]) );
  DFF_X1 \mem_reg[0][36]  ( .D(n8), .CK(clk), .Q(\mem[0][36] ) );
  DFF_X1 \data_out_reg[36]  ( .D(\mem[0][36] ), .CK(clk), .Q(data_out[36]) );
  DFF_X1 \mem_reg[0][35]  ( .D(n9), .CK(clk), .Q(\mem[0][35] ) );
  DFF_X1 \data_out_reg[35]  ( .D(\mem[0][35] ), .CK(clk), .Q(data_out[35]) );
  DFF_X1 \mem_reg[0][34]  ( .D(n10), .CK(clk), .Q(\mem[0][34] ) );
  DFF_X1 \data_out_reg[34]  ( .D(\mem[0][34] ), .CK(clk), .Q(data_out[34]) );
  DFF_X1 \mem_reg[0][33]  ( .D(n11), .CK(clk), .Q(\mem[0][33] ) );
  DFF_X1 \data_out_reg[33]  ( .D(\mem[0][33] ), .CK(clk), .Q(data_out[33]) );
  DFF_X1 \mem_reg[0][32]  ( .D(n12), .CK(clk), .Q(\mem[0][32] ) );
  DFF_X1 \data_out_reg[32]  ( .D(\mem[0][32] ), .CK(clk), .Q(data_out[32]) );
  DFF_X1 \mem_reg[0][31]  ( .D(n13), .CK(clk), .Q(\mem[0][31] ) );
  DFF_X1 \data_out_reg[31]  ( .D(\mem[0][31] ), .CK(clk), .Q(data_out[31]) );
  DFF_X1 \mem_reg[0][30]  ( .D(n14), .CK(clk), .Q(\mem[0][30] ) );
  DFF_X1 \data_out_reg[30]  ( .D(\mem[0][30] ), .CK(clk), .Q(data_out[30]) );
  DFF_X1 \mem_reg[0][29]  ( .D(n15), .CK(clk), .Q(\mem[0][29] ) );
  DFF_X1 \data_out_reg[29]  ( .D(\mem[0][29] ), .CK(clk), .Q(data_out[29]) );
  DFF_X1 \mem_reg[0][28]  ( .D(n16), .CK(clk), .Q(\mem[0][28] ) );
  DFF_X1 \data_out_reg[28]  ( .D(\mem[0][28] ), .CK(clk), .Q(data_out[28]) );
  DFF_X1 \mem_reg[0][27]  ( .D(n17), .CK(clk), .Q(\mem[0][27] ) );
  DFF_X1 \data_out_reg[27]  ( .D(\mem[0][27] ), .CK(clk), .Q(data_out[27]) );
  DFF_X1 \mem_reg[0][26]  ( .D(n18), .CK(clk), .Q(\mem[0][26] ) );
  DFF_X1 \data_out_reg[26]  ( .D(\mem[0][26] ), .CK(clk), .Q(data_out[26]) );
  DFF_X1 \mem_reg[0][25]  ( .D(n19), .CK(clk), .Q(\mem[0][25] ) );
  DFF_X1 \data_out_reg[25]  ( .D(\mem[0][25] ), .CK(clk), .Q(data_out[25]) );
  DFF_X1 \mem_reg[0][24]  ( .D(n20), .CK(clk), .Q(\mem[0][24] ) );
  DFF_X1 \data_out_reg[24]  ( .D(\mem[0][24] ), .CK(clk), .Q(data_out[24]) );
  DFF_X1 \mem_reg[0][23]  ( .D(n21), .CK(clk), .Q(\mem[0][23] ) );
  DFF_X1 \data_out_reg[23]  ( .D(\mem[0][23] ), .CK(clk), .Q(data_out[23]) );
  DFF_X1 \mem_reg[0][22]  ( .D(n22), .CK(clk), .Q(\mem[0][22] ) );
  DFF_X1 \data_out_reg[22]  ( .D(\mem[0][22] ), .CK(clk), .Q(data_out[22]) );
  DFF_X1 \mem_reg[0][21]  ( .D(n23), .CK(clk), .Q(\mem[0][21] ) );
  DFF_X1 \data_out_reg[21]  ( .D(\mem[0][21] ), .CK(clk), .Q(data_out[21]) );
  DFF_X1 \mem_reg[0][20]  ( .D(n24), .CK(clk), .Q(\mem[0][20] ) );
  DFF_X1 \data_out_reg[20]  ( .D(\mem[0][20] ), .CK(clk), .Q(data_out[20]) );
  DFF_X1 \mem_reg[0][19]  ( .D(n25), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \data_out_reg[19]  ( .D(\mem[0][19] ), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \mem_reg[0][18]  ( .D(n26), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \data_out_reg[18]  ( .D(\mem[0][18] ), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \mem_reg[0][17]  ( .D(n27), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \data_out_reg[17]  ( .D(\mem[0][17] ), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \mem_reg[0][16]  ( .D(n28), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \data_out_reg[16]  ( .D(\mem[0][16] ), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \mem_reg[0][15]  ( .D(n29), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n30), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n31), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n32), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n33), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n34), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n35), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n36), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n37), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n38), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n39), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n40), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n41), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n42), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n44), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n85), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  AND3_X1 U3 ( .A1(wr_en), .A2(n86), .A3(n87), .ZN(n1) );
  INV_X1 U4 ( .A(n1), .ZN(n3) );
  INV_X1 U5 ( .A(n1), .ZN(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n4) );
  INV_X1 U7 ( .A(addr[0]), .ZN(n86) );
  NOR3_X1 U8 ( .A1(addr[1]), .A2(addr[3]), .A3(addr[2]), .ZN(n87) );
  INV_X1 U9 ( .A(n127), .ZN(n85) );
  AOI22_X1 U10 ( .A1(\mem[0][0] ), .A2(n3), .B1(data_in[0]), .B2(n4), .ZN(n127) );
  INV_X1 U11 ( .A(n126), .ZN(n44) );
  AOI22_X1 U12 ( .A1(\mem[0][1] ), .A2(n2), .B1(data_in[1]), .B2(n1), .ZN(n126) );
  INV_X1 U13 ( .A(n125), .ZN(n42) );
  AOI22_X1 U14 ( .A1(\mem[0][2] ), .A2(n2), .B1(data_in[2]), .B2(n4), .ZN(n125) );
  INV_X1 U15 ( .A(n124), .ZN(n41) );
  AOI22_X1 U16 ( .A1(\mem[0][3] ), .A2(n3), .B1(data_in[3]), .B2(n4), .ZN(n124) );
  INV_X1 U17 ( .A(n123), .ZN(n40) );
  AOI22_X1 U18 ( .A1(\mem[0][4] ), .A2(n3), .B1(data_in[4]), .B2(n1), .ZN(n123) );
  INV_X1 U19 ( .A(n122), .ZN(n39) );
  AOI22_X1 U20 ( .A1(\mem[0][5] ), .A2(n3), .B1(data_in[5]), .B2(n4), .ZN(n122) );
  INV_X1 U21 ( .A(n121), .ZN(n38) );
  AOI22_X1 U22 ( .A1(\mem[0][6] ), .A2(n3), .B1(data_in[6]), .B2(n1), .ZN(n121) );
  INV_X1 U23 ( .A(n120), .ZN(n37) );
  AOI22_X1 U24 ( .A1(\mem[0][7] ), .A2(n3), .B1(data_in[7]), .B2(n1), .ZN(n120) );
  INV_X1 U25 ( .A(n119), .ZN(n36) );
  AOI22_X1 U26 ( .A1(\mem[0][8] ), .A2(n3), .B1(data_in[8]), .B2(n1), .ZN(n119) );
  INV_X1 U27 ( .A(n118), .ZN(n35) );
  AOI22_X1 U28 ( .A1(\mem[0][9] ), .A2(n3), .B1(data_in[9]), .B2(n4), .ZN(n118) );
  INV_X1 U29 ( .A(n117), .ZN(n34) );
  AOI22_X1 U30 ( .A1(\mem[0][10] ), .A2(n3), .B1(data_in[10]), .B2(n4), .ZN(
        n117) );
  INV_X1 U31 ( .A(n115), .ZN(n32) );
  AOI22_X1 U32 ( .A1(\mem[0][12] ), .A2(n3), .B1(data_in[12]), .B2(n1), .ZN(
        n115) );
  INV_X1 U33 ( .A(n114), .ZN(n31) );
  AOI22_X1 U34 ( .A1(\mem[0][13] ), .A2(n3), .B1(data_in[13]), .B2(n1), .ZN(
        n114) );
  INV_X1 U35 ( .A(n113), .ZN(n30) );
  AOI22_X1 U36 ( .A1(\mem[0][14] ), .A2(n3), .B1(data_in[14]), .B2(n1), .ZN(
        n113) );
  INV_X1 U37 ( .A(n112), .ZN(n29) );
  AOI22_X1 U38 ( .A1(\mem[0][15] ), .A2(n3), .B1(data_in[15]), .B2(n4), .ZN(
        n112) );
  INV_X1 U39 ( .A(n111), .ZN(n28) );
  AOI22_X1 U40 ( .A1(\mem[0][16] ), .A2(n2), .B1(data_in[16]), .B2(n4), .ZN(
        n111) );
  INV_X1 U41 ( .A(n110), .ZN(n27) );
  AOI22_X1 U42 ( .A1(\mem[0][17] ), .A2(n2), .B1(data_in[17]), .B2(n4), .ZN(
        n110) );
  INV_X1 U43 ( .A(n109), .ZN(n26) );
  AOI22_X1 U44 ( .A1(\mem[0][18] ), .A2(n2), .B1(data_in[18]), .B2(n4), .ZN(
        n109) );
  INV_X1 U45 ( .A(n108), .ZN(n25) );
  AOI22_X1 U46 ( .A1(\mem[0][19] ), .A2(n2), .B1(data_in[19]), .B2(n4), .ZN(
        n108) );
  INV_X1 U47 ( .A(n107), .ZN(n24) );
  AOI22_X1 U48 ( .A1(\mem[0][20] ), .A2(n2), .B1(data_in[20]), .B2(n1), .ZN(
        n107) );
  INV_X1 U49 ( .A(n106), .ZN(n23) );
  AOI22_X1 U50 ( .A1(\mem[0][21] ), .A2(n2), .B1(data_in[21]), .B2(n1), .ZN(
        n106) );
  INV_X1 U51 ( .A(n105), .ZN(n22) );
  AOI22_X1 U52 ( .A1(\mem[0][22] ), .A2(n2), .B1(data_in[22]), .B2(n1), .ZN(
        n105) );
  INV_X1 U53 ( .A(n104), .ZN(n21) );
  AOI22_X1 U54 ( .A1(\mem[0][23] ), .A2(n2), .B1(data_in[23]), .B2(n1), .ZN(
        n104) );
  INV_X1 U55 ( .A(n103), .ZN(n20) );
  AOI22_X1 U56 ( .A1(\mem[0][24] ), .A2(n2), .B1(data_in[24]), .B2(n1), .ZN(
        n103) );
  INV_X1 U57 ( .A(n102), .ZN(n19) );
  AOI22_X1 U58 ( .A1(\mem[0][25] ), .A2(n2), .B1(data_in[25]), .B2(n4), .ZN(
        n102) );
  INV_X1 U59 ( .A(n101), .ZN(n18) );
  AOI22_X1 U60 ( .A1(\mem[0][26] ), .A2(n2), .B1(data_in[26]), .B2(n1), .ZN(
        n101) );
  INV_X1 U61 ( .A(n100), .ZN(n17) );
  AOI22_X1 U62 ( .A1(\mem[0][27] ), .A2(n2), .B1(data_in[27]), .B2(n1), .ZN(
        n100) );
  INV_X1 U63 ( .A(n99), .ZN(n16) );
  AOI22_X1 U64 ( .A1(\mem[0][28] ), .A2(n3), .B1(data_in[28]), .B2(n4), .ZN(
        n99) );
  INV_X1 U65 ( .A(n98), .ZN(n15) );
  AOI22_X1 U66 ( .A1(\mem[0][29] ), .A2(n2), .B1(data_in[29]), .B2(n1), .ZN(
        n98) );
  INV_X1 U67 ( .A(n97), .ZN(n14) );
  AOI22_X1 U68 ( .A1(\mem[0][30] ), .A2(n3), .B1(data_in[30]), .B2(n1), .ZN(
        n97) );
  INV_X1 U69 ( .A(n96), .ZN(n13) );
  AOI22_X1 U70 ( .A1(\mem[0][31] ), .A2(n2), .B1(data_in[31]), .B2(n4), .ZN(
        n96) );
  INV_X1 U71 ( .A(n116), .ZN(n33) );
  AOI22_X1 U72 ( .A1(\mem[0][11] ), .A2(n3), .B1(data_in[11]), .B2(n1), .ZN(
        n116) );
  INV_X1 U73 ( .A(n95), .ZN(n12) );
  AOI22_X1 U74 ( .A1(\mem[0][32] ), .A2(n3), .B1(data_in[32]), .B2(n1), .ZN(
        n95) );
  INV_X1 U75 ( .A(n94), .ZN(n11) );
  AOI22_X1 U76 ( .A1(\mem[0][33] ), .A2(n2), .B1(data_in[33]), .B2(n1), .ZN(
        n94) );
  INV_X1 U77 ( .A(n93), .ZN(n10) );
  AOI22_X1 U78 ( .A1(\mem[0][34] ), .A2(n3), .B1(data_in[34]), .B2(n4), .ZN(
        n93) );
  INV_X1 U79 ( .A(n92), .ZN(n9) );
  AOI22_X1 U80 ( .A1(\mem[0][35] ), .A2(n2), .B1(data_in[35]), .B2(n1), .ZN(
        n92) );
  INV_X1 U81 ( .A(n91), .ZN(n8) );
  AOI22_X1 U82 ( .A1(\mem[0][36] ), .A2(n3), .B1(data_in[36]), .B2(n4), .ZN(
        n91) );
  INV_X1 U83 ( .A(n90), .ZN(n7) );
  AOI22_X1 U84 ( .A1(\mem[0][37] ), .A2(n2), .B1(data_in[37]), .B2(n1), .ZN(
        n90) );
  INV_X1 U85 ( .A(n89), .ZN(n6) );
  AOI22_X1 U86 ( .A1(\mem[0][38] ), .A2(n3), .B1(data_in[38]), .B2(n1), .ZN(
        n89) );
  INV_X1 U87 ( .A(n88), .ZN(n5) );
  AOI22_X1 U88 ( .A1(\mem[0][39] ), .A2(n2), .B1(data_in[39]), .B2(n4), .ZN(
        n88) );
endmodule


module memory_WIDTH40_SIZE1_LOGSIZE4_5 ( clk, data_in, data_out, addr, wr_en
 );
  input [39:0] data_in;
  output [39:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   \mem[0][39] , \mem[0][38] , \mem[0][37] , \mem[0][36] , \mem[0][35] ,
         \mem[0][34] , \mem[0][33] , \mem[0][32] , \mem[0][31] , \mem[0][30] ,
         \mem[0][29] , \mem[0][28] , \mem[0][27] , \mem[0][26] , \mem[0][25] ,
         \mem[0][24] , \mem[0][23] , \mem[0][22] , \mem[0][21] , \mem[0][20] ,
         \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] , \mem[0][15] ,
         \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] ,
         \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  DFF_X1 \mem_reg[0][39]  ( .D(n5), .CK(clk), .Q(\mem[0][39] ) );
  DFF_X1 \data_out_reg[39]  ( .D(\mem[0][39] ), .CK(clk), .Q(data_out[39]) );
  DFF_X1 \mem_reg[0][38]  ( .D(n6), .CK(clk), .Q(\mem[0][38] ) );
  DFF_X1 \data_out_reg[38]  ( .D(\mem[0][38] ), .CK(clk), .Q(data_out[38]) );
  DFF_X1 \mem_reg[0][37]  ( .D(n7), .CK(clk), .Q(\mem[0][37] ) );
  DFF_X1 \data_out_reg[37]  ( .D(\mem[0][37] ), .CK(clk), .Q(data_out[37]) );
  DFF_X1 \mem_reg[0][36]  ( .D(n8), .CK(clk), .Q(\mem[0][36] ) );
  DFF_X1 \data_out_reg[36]  ( .D(\mem[0][36] ), .CK(clk), .Q(data_out[36]) );
  DFF_X1 \mem_reg[0][35]  ( .D(n9), .CK(clk), .Q(\mem[0][35] ) );
  DFF_X1 \data_out_reg[35]  ( .D(\mem[0][35] ), .CK(clk), .Q(data_out[35]) );
  DFF_X1 \mem_reg[0][34]  ( .D(n10), .CK(clk), .Q(\mem[0][34] ) );
  DFF_X1 \data_out_reg[34]  ( .D(\mem[0][34] ), .CK(clk), .Q(data_out[34]) );
  DFF_X1 \mem_reg[0][33]  ( .D(n11), .CK(clk), .Q(\mem[0][33] ) );
  DFF_X1 \data_out_reg[33]  ( .D(\mem[0][33] ), .CK(clk), .Q(data_out[33]) );
  DFF_X1 \mem_reg[0][32]  ( .D(n12), .CK(clk), .Q(\mem[0][32] ) );
  DFF_X1 \data_out_reg[32]  ( .D(\mem[0][32] ), .CK(clk), .Q(data_out[32]) );
  DFF_X1 \mem_reg[0][31]  ( .D(n13), .CK(clk), .Q(\mem[0][31] ) );
  DFF_X1 \data_out_reg[31]  ( .D(\mem[0][31] ), .CK(clk), .Q(data_out[31]) );
  DFF_X1 \mem_reg[0][30]  ( .D(n14), .CK(clk), .Q(\mem[0][30] ) );
  DFF_X1 \data_out_reg[30]  ( .D(\mem[0][30] ), .CK(clk), .Q(data_out[30]) );
  DFF_X1 \mem_reg[0][29]  ( .D(n15), .CK(clk), .Q(\mem[0][29] ) );
  DFF_X1 \data_out_reg[29]  ( .D(\mem[0][29] ), .CK(clk), .Q(data_out[29]) );
  DFF_X1 \mem_reg[0][28]  ( .D(n16), .CK(clk), .Q(\mem[0][28] ) );
  DFF_X1 \data_out_reg[28]  ( .D(\mem[0][28] ), .CK(clk), .Q(data_out[28]) );
  DFF_X1 \mem_reg[0][27]  ( .D(n17), .CK(clk), .Q(\mem[0][27] ) );
  DFF_X1 \data_out_reg[27]  ( .D(\mem[0][27] ), .CK(clk), .Q(data_out[27]) );
  DFF_X1 \mem_reg[0][26]  ( .D(n18), .CK(clk), .Q(\mem[0][26] ) );
  DFF_X1 \data_out_reg[26]  ( .D(\mem[0][26] ), .CK(clk), .Q(data_out[26]) );
  DFF_X1 \mem_reg[0][25]  ( .D(n19), .CK(clk), .Q(\mem[0][25] ) );
  DFF_X1 \data_out_reg[25]  ( .D(\mem[0][25] ), .CK(clk), .Q(data_out[25]) );
  DFF_X1 \mem_reg[0][24]  ( .D(n20), .CK(clk), .Q(\mem[0][24] ) );
  DFF_X1 \data_out_reg[24]  ( .D(\mem[0][24] ), .CK(clk), .Q(data_out[24]) );
  DFF_X1 \mem_reg[0][23]  ( .D(n21), .CK(clk), .Q(\mem[0][23] ) );
  DFF_X1 \data_out_reg[23]  ( .D(\mem[0][23] ), .CK(clk), .Q(data_out[23]) );
  DFF_X1 \mem_reg[0][22]  ( .D(n22), .CK(clk), .Q(\mem[0][22] ) );
  DFF_X1 \data_out_reg[22]  ( .D(\mem[0][22] ), .CK(clk), .Q(data_out[22]) );
  DFF_X1 \mem_reg[0][21]  ( .D(n23), .CK(clk), .Q(\mem[0][21] ) );
  DFF_X1 \data_out_reg[21]  ( .D(\mem[0][21] ), .CK(clk), .Q(data_out[21]) );
  DFF_X1 \mem_reg[0][20]  ( .D(n24), .CK(clk), .Q(\mem[0][20] ) );
  DFF_X1 \data_out_reg[20]  ( .D(\mem[0][20] ), .CK(clk), .Q(data_out[20]) );
  DFF_X1 \mem_reg[0][19]  ( .D(n25), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \data_out_reg[19]  ( .D(\mem[0][19] ), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \mem_reg[0][18]  ( .D(n26), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \data_out_reg[18]  ( .D(\mem[0][18] ), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \mem_reg[0][17]  ( .D(n27), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \data_out_reg[17]  ( .D(\mem[0][17] ), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \mem_reg[0][16]  ( .D(n28), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \data_out_reg[16]  ( .D(\mem[0][16] ), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \mem_reg[0][15]  ( .D(n29), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n30), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n31), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n32), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n33), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n34), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n35), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n36), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n37), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n38), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n39), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n40), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n41), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n42), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n44), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n85), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  AND3_X1 U3 ( .A1(wr_en), .A2(n86), .A3(n87), .ZN(n1) );
  INV_X1 U4 ( .A(n1), .ZN(n3) );
  INV_X1 U5 ( .A(n1), .ZN(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n4) );
  INV_X1 U7 ( .A(addr[0]), .ZN(n86) );
  NOR3_X1 U8 ( .A1(addr[1]), .A2(addr[3]), .A3(addr[2]), .ZN(n87) );
  INV_X1 U9 ( .A(n127), .ZN(n85) );
  AOI22_X1 U10 ( .A1(\mem[0][0] ), .A2(n3), .B1(data_in[0]), .B2(n4), .ZN(n127) );
  INV_X1 U11 ( .A(n126), .ZN(n44) );
  AOI22_X1 U12 ( .A1(\mem[0][1] ), .A2(n2), .B1(data_in[1]), .B2(n4), .ZN(n126) );
  INV_X1 U13 ( .A(n125), .ZN(n42) );
  AOI22_X1 U14 ( .A1(\mem[0][2] ), .A2(n2), .B1(data_in[2]), .B2(n1), .ZN(n125) );
  INV_X1 U15 ( .A(n124), .ZN(n41) );
  AOI22_X1 U16 ( .A1(\mem[0][3] ), .A2(n3), .B1(data_in[3]), .B2(n4), .ZN(n124) );
  INV_X1 U17 ( .A(n123), .ZN(n40) );
  AOI22_X1 U18 ( .A1(\mem[0][4] ), .A2(n3), .B1(data_in[4]), .B2(n4), .ZN(n123) );
  INV_X1 U19 ( .A(n122), .ZN(n39) );
  AOI22_X1 U20 ( .A1(\mem[0][5] ), .A2(n3), .B1(data_in[5]), .B2(n4), .ZN(n122) );
  INV_X1 U21 ( .A(n121), .ZN(n38) );
  AOI22_X1 U22 ( .A1(\mem[0][6] ), .A2(n3), .B1(data_in[6]), .B2(n4), .ZN(n121) );
  INV_X1 U23 ( .A(n120), .ZN(n37) );
  AOI22_X1 U24 ( .A1(\mem[0][7] ), .A2(n3), .B1(data_in[7]), .B2(n4), .ZN(n120) );
  INV_X1 U25 ( .A(n119), .ZN(n36) );
  AOI22_X1 U26 ( .A1(\mem[0][8] ), .A2(n3), .B1(data_in[8]), .B2(n1), .ZN(n119) );
  INV_X1 U27 ( .A(n118), .ZN(n35) );
  AOI22_X1 U28 ( .A1(\mem[0][9] ), .A2(n3), .B1(data_in[9]), .B2(n1), .ZN(n118) );
  INV_X1 U29 ( .A(n117), .ZN(n34) );
  AOI22_X1 U30 ( .A1(\mem[0][10] ), .A2(n3), .B1(data_in[10]), .B2(n1), .ZN(
        n117) );
  INV_X1 U31 ( .A(n115), .ZN(n32) );
  AOI22_X1 U32 ( .A1(\mem[0][12] ), .A2(n3), .B1(data_in[12]), .B2(n1), .ZN(
        n115) );
  INV_X1 U33 ( .A(n114), .ZN(n31) );
  AOI22_X1 U34 ( .A1(\mem[0][13] ), .A2(n3), .B1(data_in[13]), .B2(n4), .ZN(
        n114) );
  INV_X1 U35 ( .A(n113), .ZN(n30) );
  AOI22_X1 U36 ( .A1(\mem[0][14] ), .A2(n3), .B1(data_in[14]), .B2(n1), .ZN(
        n113) );
  INV_X1 U37 ( .A(n112), .ZN(n29) );
  AOI22_X1 U38 ( .A1(\mem[0][15] ), .A2(n3), .B1(data_in[15]), .B2(n4), .ZN(
        n112) );
  INV_X1 U39 ( .A(n111), .ZN(n28) );
  AOI22_X1 U40 ( .A1(\mem[0][16] ), .A2(n2), .B1(data_in[16]), .B2(n1), .ZN(
        n111) );
  INV_X1 U41 ( .A(n110), .ZN(n27) );
  AOI22_X1 U42 ( .A1(\mem[0][17] ), .A2(n2), .B1(data_in[17]), .B2(n1), .ZN(
        n110) );
  INV_X1 U43 ( .A(n109), .ZN(n26) );
  AOI22_X1 U44 ( .A1(\mem[0][18] ), .A2(n2), .B1(data_in[18]), .B2(n4), .ZN(
        n109) );
  INV_X1 U45 ( .A(n108), .ZN(n25) );
  AOI22_X1 U46 ( .A1(\mem[0][19] ), .A2(n2), .B1(data_in[19]), .B2(n1), .ZN(
        n108) );
  INV_X1 U47 ( .A(n107), .ZN(n24) );
  AOI22_X1 U48 ( .A1(\mem[0][20] ), .A2(n2), .B1(data_in[20]), .B2(n4), .ZN(
        n107) );
  INV_X1 U49 ( .A(n106), .ZN(n23) );
  AOI22_X1 U50 ( .A1(\mem[0][21] ), .A2(n2), .B1(data_in[21]), .B2(n1), .ZN(
        n106) );
  INV_X1 U51 ( .A(n105), .ZN(n22) );
  AOI22_X1 U52 ( .A1(\mem[0][22] ), .A2(n2), .B1(data_in[22]), .B2(n1), .ZN(
        n105) );
  INV_X1 U53 ( .A(n104), .ZN(n21) );
  AOI22_X1 U54 ( .A1(\mem[0][23] ), .A2(n2), .B1(data_in[23]), .B2(n1), .ZN(
        n104) );
  INV_X1 U55 ( .A(n103), .ZN(n20) );
  AOI22_X1 U56 ( .A1(\mem[0][24] ), .A2(n2), .B1(data_in[24]), .B2(n4), .ZN(
        n103) );
  INV_X1 U57 ( .A(n102), .ZN(n19) );
  AOI22_X1 U58 ( .A1(\mem[0][25] ), .A2(n2), .B1(data_in[25]), .B2(n4), .ZN(
        n102) );
  INV_X1 U59 ( .A(n101), .ZN(n18) );
  AOI22_X1 U60 ( .A1(\mem[0][26] ), .A2(n2), .B1(data_in[26]), .B2(n4), .ZN(
        n101) );
  INV_X1 U61 ( .A(n100), .ZN(n17) );
  AOI22_X1 U62 ( .A1(\mem[0][27] ), .A2(n2), .B1(data_in[27]), .B2(n1), .ZN(
        n100) );
  INV_X1 U63 ( .A(n99), .ZN(n16) );
  AOI22_X1 U64 ( .A1(\mem[0][28] ), .A2(n3), .B1(data_in[28]), .B2(n1), .ZN(
        n99) );
  INV_X1 U65 ( .A(n98), .ZN(n15) );
  AOI22_X1 U66 ( .A1(\mem[0][29] ), .A2(n2), .B1(data_in[29]), .B2(n1), .ZN(
        n98) );
  INV_X1 U67 ( .A(n97), .ZN(n14) );
  AOI22_X1 U68 ( .A1(\mem[0][30] ), .A2(n3), .B1(data_in[30]), .B2(n4), .ZN(
        n97) );
  INV_X1 U69 ( .A(n96), .ZN(n13) );
  AOI22_X1 U70 ( .A1(\mem[0][31] ), .A2(n2), .B1(data_in[31]), .B2(n1), .ZN(
        n96) );
  INV_X1 U71 ( .A(n116), .ZN(n33) );
  AOI22_X1 U72 ( .A1(\mem[0][11] ), .A2(n3), .B1(data_in[11]), .B2(n1), .ZN(
        n116) );
  INV_X1 U73 ( .A(n95), .ZN(n12) );
  AOI22_X1 U74 ( .A1(\mem[0][32] ), .A2(n3), .B1(data_in[32]), .B2(n4), .ZN(
        n95) );
  INV_X1 U75 ( .A(n94), .ZN(n11) );
  AOI22_X1 U76 ( .A1(\mem[0][33] ), .A2(n2), .B1(data_in[33]), .B2(n1), .ZN(
        n94) );
  INV_X1 U77 ( .A(n93), .ZN(n10) );
  AOI22_X1 U78 ( .A1(\mem[0][34] ), .A2(n3), .B1(data_in[34]), .B2(n1), .ZN(
        n93) );
  INV_X1 U79 ( .A(n92), .ZN(n9) );
  AOI22_X1 U80 ( .A1(\mem[0][35] ), .A2(n2), .B1(data_in[35]), .B2(n1), .ZN(
        n92) );
  INV_X1 U81 ( .A(n91), .ZN(n8) );
  AOI22_X1 U82 ( .A1(\mem[0][36] ), .A2(n3), .B1(data_in[36]), .B2(n1), .ZN(
        n91) );
  INV_X1 U83 ( .A(n90), .ZN(n7) );
  AOI22_X1 U84 ( .A1(\mem[0][37] ), .A2(n2), .B1(data_in[37]), .B2(n1), .ZN(
        n90) );
  INV_X1 U85 ( .A(n89), .ZN(n6) );
  AOI22_X1 U86 ( .A1(\mem[0][38] ), .A2(n3), .B1(data_in[38]), .B2(n1), .ZN(
        n89) );
  INV_X1 U87 ( .A(n88), .ZN(n5) );
  AOI22_X1 U88 ( .A1(\mem[0][39] ), .A2(n2), .B1(data_in[39]), .B2(n4), .ZN(
        n88) );
endmodule


module memory_WIDTH40_SIZE1_LOGSIZE4_4 ( clk, data_in, data_out, addr, wr_en
 );
  input [39:0] data_in;
  output [39:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   \mem[0][39] , \mem[0][38] , \mem[0][37] , \mem[0][36] , \mem[0][35] ,
         \mem[0][34] , \mem[0][33] , \mem[0][32] , \mem[0][31] , \mem[0][30] ,
         \mem[0][29] , \mem[0][28] , \mem[0][27] , \mem[0][26] , \mem[0][25] ,
         \mem[0][24] , \mem[0][23] , \mem[0][22] , \mem[0][21] , \mem[0][20] ,
         \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] , \mem[0][15] ,
         \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] ,
         \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  DFF_X1 \mem_reg[0][39]  ( .D(n5), .CK(clk), .Q(\mem[0][39] ) );
  DFF_X1 \data_out_reg[39]  ( .D(\mem[0][39] ), .CK(clk), .Q(data_out[39]) );
  DFF_X1 \mem_reg[0][38]  ( .D(n6), .CK(clk), .Q(\mem[0][38] ) );
  DFF_X1 \data_out_reg[38]  ( .D(\mem[0][38] ), .CK(clk), .Q(data_out[38]) );
  DFF_X1 \mem_reg[0][37]  ( .D(n7), .CK(clk), .Q(\mem[0][37] ) );
  DFF_X1 \data_out_reg[37]  ( .D(\mem[0][37] ), .CK(clk), .Q(data_out[37]) );
  DFF_X1 \mem_reg[0][36]  ( .D(n8), .CK(clk), .Q(\mem[0][36] ) );
  DFF_X1 \data_out_reg[36]  ( .D(\mem[0][36] ), .CK(clk), .Q(data_out[36]) );
  DFF_X1 \mem_reg[0][35]  ( .D(n9), .CK(clk), .Q(\mem[0][35] ) );
  DFF_X1 \data_out_reg[35]  ( .D(\mem[0][35] ), .CK(clk), .Q(data_out[35]) );
  DFF_X1 \mem_reg[0][34]  ( .D(n10), .CK(clk), .Q(\mem[0][34] ) );
  DFF_X1 \data_out_reg[34]  ( .D(\mem[0][34] ), .CK(clk), .Q(data_out[34]) );
  DFF_X1 \mem_reg[0][33]  ( .D(n11), .CK(clk), .Q(\mem[0][33] ) );
  DFF_X1 \data_out_reg[33]  ( .D(\mem[0][33] ), .CK(clk), .Q(data_out[33]) );
  DFF_X1 \mem_reg[0][32]  ( .D(n12), .CK(clk), .Q(\mem[0][32] ) );
  DFF_X1 \data_out_reg[32]  ( .D(\mem[0][32] ), .CK(clk), .Q(data_out[32]) );
  DFF_X1 \mem_reg[0][31]  ( .D(n13), .CK(clk), .Q(\mem[0][31] ) );
  DFF_X1 \data_out_reg[31]  ( .D(\mem[0][31] ), .CK(clk), .Q(data_out[31]) );
  DFF_X1 \mem_reg[0][30]  ( .D(n14), .CK(clk), .Q(\mem[0][30] ) );
  DFF_X1 \data_out_reg[30]  ( .D(\mem[0][30] ), .CK(clk), .Q(data_out[30]) );
  DFF_X1 \mem_reg[0][29]  ( .D(n15), .CK(clk), .Q(\mem[0][29] ) );
  DFF_X1 \data_out_reg[29]  ( .D(\mem[0][29] ), .CK(clk), .Q(data_out[29]) );
  DFF_X1 \mem_reg[0][28]  ( .D(n16), .CK(clk), .Q(\mem[0][28] ) );
  DFF_X1 \data_out_reg[28]  ( .D(\mem[0][28] ), .CK(clk), .Q(data_out[28]) );
  DFF_X1 \mem_reg[0][27]  ( .D(n17), .CK(clk), .Q(\mem[0][27] ) );
  DFF_X1 \data_out_reg[27]  ( .D(\mem[0][27] ), .CK(clk), .Q(data_out[27]) );
  DFF_X1 \mem_reg[0][26]  ( .D(n18), .CK(clk), .Q(\mem[0][26] ) );
  DFF_X1 \data_out_reg[26]  ( .D(\mem[0][26] ), .CK(clk), .Q(data_out[26]) );
  DFF_X1 \mem_reg[0][25]  ( .D(n19), .CK(clk), .Q(\mem[0][25] ) );
  DFF_X1 \data_out_reg[25]  ( .D(\mem[0][25] ), .CK(clk), .Q(data_out[25]) );
  DFF_X1 \mem_reg[0][24]  ( .D(n20), .CK(clk), .Q(\mem[0][24] ) );
  DFF_X1 \data_out_reg[24]  ( .D(\mem[0][24] ), .CK(clk), .Q(data_out[24]) );
  DFF_X1 \mem_reg[0][23]  ( .D(n21), .CK(clk), .Q(\mem[0][23] ) );
  DFF_X1 \data_out_reg[23]  ( .D(\mem[0][23] ), .CK(clk), .Q(data_out[23]) );
  DFF_X1 \mem_reg[0][22]  ( .D(n22), .CK(clk), .Q(\mem[0][22] ) );
  DFF_X1 \data_out_reg[22]  ( .D(\mem[0][22] ), .CK(clk), .Q(data_out[22]) );
  DFF_X1 \mem_reg[0][21]  ( .D(n23), .CK(clk), .Q(\mem[0][21] ) );
  DFF_X1 \data_out_reg[21]  ( .D(\mem[0][21] ), .CK(clk), .Q(data_out[21]) );
  DFF_X1 \mem_reg[0][20]  ( .D(n24), .CK(clk), .Q(\mem[0][20] ) );
  DFF_X1 \data_out_reg[20]  ( .D(\mem[0][20] ), .CK(clk), .Q(data_out[20]) );
  DFF_X1 \mem_reg[0][19]  ( .D(n25), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \data_out_reg[19]  ( .D(\mem[0][19] ), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \mem_reg[0][18]  ( .D(n26), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \data_out_reg[18]  ( .D(\mem[0][18] ), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \mem_reg[0][17]  ( .D(n27), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \data_out_reg[17]  ( .D(\mem[0][17] ), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \mem_reg[0][16]  ( .D(n28), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \data_out_reg[16]  ( .D(\mem[0][16] ), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \mem_reg[0][15]  ( .D(n29), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n30), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n31), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n32), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n33), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n34), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n35), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n36), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n37), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n38), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n39), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n40), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n41), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n42), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n44), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n85), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  AND3_X1 U3 ( .A1(wr_en), .A2(n86), .A3(n87), .ZN(n1) );
  INV_X1 U4 ( .A(n1), .ZN(n3) );
  INV_X1 U5 ( .A(n1), .ZN(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n4) );
  INV_X1 U7 ( .A(addr[0]), .ZN(n86) );
  NOR3_X1 U8 ( .A1(addr[1]), .A2(addr[3]), .A3(addr[2]), .ZN(n87) );
  INV_X1 U9 ( .A(n127), .ZN(n85) );
  INV_X1 U10 ( .A(n126), .ZN(n44) );
  AOI22_X1 U11 ( .A1(\mem[0][1] ), .A2(n3), .B1(data_in[1]), .B2(n1), .ZN(n126) );
  INV_X1 U12 ( .A(n125), .ZN(n42) );
  AOI22_X1 U13 ( .A1(\mem[0][2] ), .A2(n2), .B1(data_in[2]), .B2(n1), .ZN(n125) );
  INV_X1 U14 ( .A(n123), .ZN(n40) );
  AOI22_X1 U15 ( .A1(\mem[0][4] ), .A2(n3), .B1(data_in[4]), .B2(n4), .ZN(n123) );
  INV_X1 U16 ( .A(n121), .ZN(n38) );
  AOI22_X1 U17 ( .A1(\mem[0][6] ), .A2(n3), .B1(data_in[6]), .B2(n4), .ZN(n121) );
  INV_X1 U18 ( .A(n119), .ZN(n36) );
  AOI22_X1 U19 ( .A1(\mem[0][8] ), .A2(n3), .B1(data_in[8]), .B2(n4), .ZN(n119) );
  INV_X1 U20 ( .A(n118), .ZN(n35) );
  AOI22_X1 U21 ( .A1(\mem[0][9] ), .A2(n3), .B1(data_in[9]), .B2(n4), .ZN(n118) );
  INV_X1 U22 ( .A(n117), .ZN(n34) );
  AOI22_X1 U23 ( .A1(\mem[0][10] ), .A2(n3), .B1(data_in[10]), .B2(n1), .ZN(
        n117) );
  INV_X1 U24 ( .A(n115), .ZN(n32) );
  AOI22_X1 U25 ( .A1(\mem[0][12] ), .A2(n3), .B1(data_in[12]), .B2(n4), .ZN(
        n115) );
  INV_X1 U26 ( .A(n114), .ZN(n31) );
  AOI22_X1 U27 ( .A1(\mem[0][13] ), .A2(n3), .B1(data_in[13]), .B2(n4), .ZN(
        n114) );
  INV_X1 U28 ( .A(n113), .ZN(n30) );
  AOI22_X1 U29 ( .A1(\mem[0][14] ), .A2(n3), .B1(data_in[14]), .B2(n4), .ZN(
        n113) );
  INV_X1 U30 ( .A(n112), .ZN(n29) );
  AOI22_X1 U31 ( .A1(\mem[0][15] ), .A2(n3), .B1(data_in[15]), .B2(n1), .ZN(
        n112) );
  INV_X1 U32 ( .A(n111), .ZN(n28) );
  AOI22_X1 U33 ( .A1(\mem[0][16] ), .A2(n2), .B1(data_in[16]), .B2(n4), .ZN(
        n111) );
  INV_X1 U34 ( .A(n110), .ZN(n27) );
  AOI22_X1 U35 ( .A1(\mem[0][17] ), .A2(n2), .B1(data_in[17]), .B2(n1), .ZN(
        n110) );
  INV_X1 U36 ( .A(n109), .ZN(n26) );
  AOI22_X1 U37 ( .A1(\mem[0][18] ), .A2(n2), .B1(data_in[18]), .B2(n1), .ZN(
        n109) );
  INV_X1 U38 ( .A(n108), .ZN(n25) );
  AOI22_X1 U39 ( .A1(\mem[0][19] ), .A2(n2), .B1(data_in[19]), .B2(n1), .ZN(
        n108) );
  INV_X1 U40 ( .A(n107), .ZN(n24) );
  AOI22_X1 U41 ( .A1(\mem[0][20] ), .A2(n2), .B1(data_in[20]), .B2(n4), .ZN(
        n107) );
  INV_X1 U42 ( .A(n106), .ZN(n23) );
  AOI22_X1 U43 ( .A1(\mem[0][21] ), .A2(n2), .B1(data_in[21]), .B2(n1), .ZN(
        n106) );
  INV_X1 U44 ( .A(n105), .ZN(n22) );
  AOI22_X1 U45 ( .A1(\mem[0][22] ), .A2(n2), .B1(data_in[22]), .B2(n4), .ZN(
        n105) );
  INV_X1 U46 ( .A(n104), .ZN(n21) );
  AOI22_X1 U47 ( .A1(\mem[0][23] ), .A2(n2), .B1(data_in[23]), .B2(n1), .ZN(
        n104) );
  INV_X1 U48 ( .A(n103), .ZN(n20) );
  AOI22_X1 U49 ( .A1(\mem[0][24] ), .A2(n2), .B1(data_in[24]), .B2(n4), .ZN(
        n103) );
  INV_X1 U50 ( .A(n102), .ZN(n19) );
  AOI22_X1 U51 ( .A1(\mem[0][25] ), .A2(n2), .B1(data_in[25]), .B2(n4), .ZN(
        n102) );
  INV_X1 U52 ( .A(n101), .ZN(n18) );
  AOI22_X1 U53 ( .A1(\mem[0][26] ), .A2(n2), .B1(data_in[26]), .B2(n1), .ZN(
        n101) );
  INV_X1 U54 ( .A(n100), .ZN(n17) );
  AOI22_X1 U55 ( .A1(\mem[0][27] ), .A2(n2), .B1(data_in[27]), .B2(n1), .ZN(
        n100) );
  INV_X1 U56 ( .A(n99), .ZN(n16) );
  AOI22_X1 U57 ( .A1(\mem[0][28] ), .A2(n3), .B1(data_in[28]), .B2(n4), .ZN(
        n99) );
  INV_X1 U58 ( .A(n98), .ZN(n15) );
  AOI22_X1 U59 ( .A1(\mem[0][29] ), .A2(n2), .B1(data_in[29]), .B2(n4), .ZN(
        n98) );
  INV_X1 U60 ( .A(n97), .ZN(n14) );
  AOI22_X1 U61 ( .A1(\mem[0][30] ), .A2(n3), .B1(data_in[30]), .B2(n4), .ZN(
        n97) );
  INV_X1 U62 ( .A(n96), .ZN(n13) );
  AOI22_X1 U63 ( .A1(\mem[0][31] ), .A2(n2), .B1(data_in[31]), .B2(n1), .ZN(
        n96) );
  INV_X1 U64 ( .A(n122), .ZN(n39) );
  AOI22_X1 U65 ( .A1(\mem[0][5] ), .A2(n3), .B1(data_in[5]), .B2(n4), .ZN(n122) );
  INV_X1 U66 ( .A(n120), .ZN(n37) );
  AOI22_X1 U67 ( .A1(\mem[0][7] ), .A2(n3), .B1(data_in[7]), .B2(n1), .ZN(n120) );
  INV_X1 U68 ( .A(n116), .ZN(n33) );
  AOI22_X1 U69 ( .A1(\mem[0][11] ), .A2(n3), .B1(data_in[11]), .B2(n1), .ZN(
        n116) );
  INV_X1 U70 ( .A(n95), .ZN(n12) );
  AOI22_X1 U71 ( .A1(\mem[0][32] ), .A2(n3), .B1(data_in[32]), .B2(n4), .ZN(
        n95) );
  INV_X1 U72 ( .A(n94), .ZN(n11) );
  AOI22_X1 U73 ( .A1(\mem[0][33] ), .A2(n2), .B1(data_in[33]), .B2(n1), .ZN(
        n94) );
  INV_X1 U74 ( .A(n93), .ZN(n10) );
  AOI22_X1 U75 ( .A1(\mem[0][34] ), .A2(n3), .B1(data_in[34]), .B2(n1), .ZN(
        n93) );
  INV_X1 U76 ( .A(n92), .ZN(n9) );
  AOI22_X1 U77 ( .A1(\mem[0][35] ), .A2(n2), .B1(data_in[35]), .B2(n1), .ZN(
        n92) );
  INV_X1 U78 ( .A(n91), .ZN(n8) );
  AOI22_X1 U79 ( .A1(\mem[0][36] ), .A2(n3), .B1(data_in[36]), .B2(n4), .ZN(
        n91) );
  INV_X1 U80 ( .A(n90), .ZN(n7) );
  AOI22_X1 U81 ( .A1(\mem[0][37] ), .A2(n2), .B1(data_in[37]), .B2(n4), .ZN(
        n90) );
  INV_X1 U82 ( .A(n89), .ZN(n6) );
  AOI22_X1 U83 ( .A1(\mem[0][38] ), .A2(n3), .B1(data_in[38]), .B2(n4), .ZN(
        n89) );
  INV_X1 U84 ( .A(n88), .ZN(n5) );
  AOI22_X1 U85 ( .A1(\mem[0][39] ), .A2(n2), .B1(data_in[39]), .B2(n4), .ZN(
        n88) );
  INV_X1 U86 ( .A(n124), .ZN(n41) );
  AOI22_X1 U87 ( .A1(\mem[0][3] ), .A2(n2), .B1(data_in[3]), .B2(n1), .ZN(n124) );
  AOI22_X1 U88 ( .A1(\mem[0][0] ), .A2(n3), .B1(data_in[0]), .B2(n1), .ZN(n127) );
endmodule


module memory_WIDTH40_SIZE1_LOGSIZE4_3 ( clk, data_in, data_out, addr, wr_en
 );
  input [39:0] data_in;
  output [39:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   \mem[0][39] , \mem[0][38] , \mem[0][37] , \mem[0][36] , \mem[0][35] ,
         \mem[0][34] , \mem[0][33] , \mem[0][32] , \mem[0][31] , \mem[0][30] ,
         \mem[0][29] , \mem[0][28] , \mem[0][27] , \mem[0][26] , \mem[0][25] ,
         \mem[0][24] , \mem[0][23] , \mem[0][22] , \mem[0][21] , \mem[0][20] ,
         \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] , \mem[0][15] ,
         \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] ,
         \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  DFF_X1 \mem_reg[0][39]  ( .D(n5), .CK(clk), .Q(\mem[0][39] ) );
  DFF_X1 \data_out_reg[39]  ( .D(\mem[0][39] ), .CK(clk), .Q(data_out[39]) );
  DFF_X1 \mem_reg[0][38]  ( .D(n6), .CK(clk), .Q(\mem[0][38] ) );
  DFF_X1 \data_out_reg[38]  ( .D(\mem[0][38] ), .CK(clk), .Q(data_out[38]) );
  DFF_X1 \mem_reg[0][37]  ( .D(n7), .CK(clk), .Q(\mem[0][37] ) );
  DFF_X1 \data_out_reg[37]  ( .D(\mem[0][37] ), .CK(clk), .Q(data_out[37]) );
  DFF_X1 \mem_reg[0][36]  ( .D(n8), .CK(clk), .Q(\mem[0][36] ) );
  DFF_X1 \data_out_reg[36]  ( .D(\mem[0][36] ), .CK(clk), .Q(data_out[36]) );
  DFF_X1 \mem_reg[0][35]  ( .D(n9), .CK(clk), .Q(\mem[0][35] ) );
  DFF_X1 \data_out_reg[35]  ( .D(\mem[0][35] ), .CK(clk), .Q(data_out[35]) );
  DFF_X1 \mem_reg[0][34]  ( .D(n10), .CK(clk), .Q(\mem[0][34] ) );
  DFF_X1 \data_out_reg[34]  ( .D(\mem[0][34] ), .CK(clk), .Q(data_out[34]) );
  DFF_X1 \mem_reg[0][33]  ( .D(n11), .CK(clk), .Q(\mem[0][33] ) );
  DFF_X1 \data_out_reg[33]  ( .D(\mem[0][33] ), .CK(clk), .Q(data_out[33]) );
  DFF_X1 \mem_reg[0][32]  ( .D(n12), .CK(clk), .Q(\mem[0][32] ) );
  DFF_X1 \data_out_reg[32]  ( .D(\mem[0][32] ), .CK(clk), .Q(data_out[32]) );
  DFF_X1 \mem_reg[0][31]  ( .D(n13), .CK(clk), .Q(\mem[0][31] ) );
  DFF_X1 \data_out_reg[31]  ( .D(\mem[0][31] ), .CK(clk), .Q(data_out[31]) );
  DFF_X1 \mem_reg[0][30]  ( .D(n14), .CK(clk), .Q(\mem[0][30] ) );
  DFF_X1 \data_out_reg[30]  ( .D(\mem[0][30] ), .CK(clk), .Q(data_out[30]) );
  DFF_X1 \mem_reg[0][29]  ( .D(n15), .CK(clk), .Q(\mem[0][29] ) );
  DFF_X1 \data_out_reg[29]  ( .D(\mem[0][29] ), .CK(clk), .Q(data_out[29]) );
  DFF_X1 \mem_reg[0][28]  ( .D(n16), .CK(clk), .Q(\mem[0][28] ) );
  DFF_X1 \data_out_reg[28]  ( .D(\mem[0][28] ), .CK(clk), .Q(data_out[28]) );
  DFF_X1 \mem_reg[0][27]  ( .D(n17), .CK(clk), .Q(\mem[0][27] ) );
  DFF_X1 \data_out_reg[27]  ( .D(\mem[0][27] ), .CK(clk), .Q(data_out[27]) );
  DFF_X1 \mem_reg[0][26]  ( .D(n18), .CK(clk), .Q(\mem[0][26] ) );
  DFF_X1 \data_out_reg[26]  ( .D(\mem[0][26] ), .CK(clk), .Q(data_out[26]) );
  DFF_X1 \mem_reg[0][25]  ( .D(n19), .CK(clk), .Q(\mem[0][25] ) );
  DFF_X1 \data_out_reg[25]  ( .D(\mem[0][25] ), .CK(clk), .Q(data_out[25]) );
  DFF_X1 \mem_reg[0][24]  ( .D(n20), .CK(clk), .Q(\mem[0][24] ) );
  DFF_X1 \data_out_reg[24]  ( .D(\mem[0][24] ), .CK(clk), .Q(data_out[24]) );
  DFF_X1 \mem_reg[0][23]  ( .D(n21), .CK(clk), .Q(\mem[0][23] ) );
  DFF_X1 \data_out_reg[23]  ( .D(\mem[0][23] ), .CK(clk), .Q(data_out[23]) );
  DFF_X1 \mem_reg[0][22]  ( .D(n22), .CK(clk), .Q(\mem[0][22] ) );
  DFF_X1 \data_out_reg[22]  ( .D(\mem[0][22] ), .CK(clk), .Q(data_out[22]) );
  DFF_X1 \mem_reg[0][21]  ( .D(n23), .CK(clk), .Q(\mem[0][21] ) );
  DFF_X1 \data_out_reg[21]  ( .D(\mem[0][21] ), .CK(clk), .Q(data_out[21]) );
  DFF_X1 \mem_reg[0][20]  ( .D(n24), .CK(clk), .Q(\mem[0][20] ) );
  DFF_X1 \data_out_reg[20]  ( .D(\mem[0][20] ), .CK(clk), .Q(data_out[20]) );
  DFF_X1 \mem_reg[0][19]  ( .D(n25), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \data_out_reg[19]  ( .D(\mem[0][19] ), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \mem_reg[0][18]  ( .D(n26), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \data_out_reg[18]  ( .D(\mem[0][18] ), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \mem_reg[0][17]  ( .D(n27), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \data_out_reg[17]  ( .D(\mem[0][17] ), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \mem_reg[0][16]  ( .D(n28), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \data_out_reg[16]  ( .D(\mem[0][16] ), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \mem_reg[0][15]  ( .D(n29), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n30), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n31), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n32), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n33), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n34), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n35), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n36), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n37), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n38), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n39), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n40), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n41), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n42), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n44), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n85), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  AND3_X1 U3 ( .A1(wr_en), .A2(n86), .A3(n87), .ZN(n1) );
  INV_X1 U4 ( .A(n1), .ZN(n3) );
  INV_X1 U5 ( .A(n1), .ZN(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n4) );
  INV_X1 U7 ( .A(addr[0]), .ZN(n86) );
  NOR3_X1 U8 ( .A1(addr[1]), .A2(addr[3]), .A3(addr[2]), .ZN(n87) );
  INV_X1 U9 ( .A(n127), .ZN(n85) );
  AOI22_X1 U10 ( .A1(\mem[0][0] ), .A2(n3), .B1(data_in[0]), .B2(n4), .ZN(n127) );
  INV_X1 U11 ( .A(n126), .ZN(n44) );
  AOI22_X1 U12 ( .A1(\mem[0][1] ), .A2(n2), .B1(data_in[1]), .B2(n4), .ZN(n126) );
  INV_X1 U13 ( .A(n125), .ZN(n42) );
  AOI22_X1 U14 ( .A1(\mem[0][2] ), .A2(n2), .B1(data_in[2]), .B2(n4), .ZN(n125) );
  INV_X1 U15 ( .A(n124), .ZN(n41) );
  AOI22_X1 U16 ( .A1(\mem[0][3] ), .A2(n3), .B1(data_in[3]), .B2(n4), .ZN(n124) );
  INV_X1 U17 ( .A(n123), .ZN(n40) );
  AOI22_X1 U18 ( .A1(\mem[0][4] ), .A2(n3), .B1(data_in[4]), .B2(n1), .ZN(n123) );
  INV_X1 U19 ( .A(n122), .ZN(n39) );
  AOI22_X1 U20 ( .A1(\mem[0][5] ), .A2(n3), .B1(data_in[5]), .B2(n1), .ZN(n122) );
  INV_X1 U21 ( .A(n121), .ZN(n38) );
  AOI22_X1 U22 ( .A1(\mem[0][6] ), .A2(n3), .B1(data_in[6]), .B2(n1), .ZN(n121) );
  INV_X1 U23 ( .A(n120), .ZN(n37) );
  AOI22_X1 U24 ( .A1(\mem[0][7] ), .A2(n3), .B1(data_in[7]), .B2(n4), .ZN(n120) );
  INV_X1 U25 ( .A(n119), .ZN(n36) );
  AOI22_X1 U26 ( .A1(\mem[0][8] ), .A2(n3), .B1(data_in[8]), .B2(n1), .ZN(n119) );
  INV_X1 U27 ( .A(n117), .ZN(n34) );
  AOI22_X1 U28 ( .A1(\mem[0][10] ), .A2(n3), .B1(data_in[10]), .B2(n1), .ZN(
        n117) );
  INV_X1 U29 ( .A(n115), .ZN(n32) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n3), .B1(data_in[12]), .B2(n4), .ZN(
        n115) );
  INV_X1 U31 ( .A(n114), .ZN(n31) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n3), .B1(data_in[13]), .B2(n1), .ZN(
        n114) );
  INV_X1 U33 ( .A(n113), .ZN(n30) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n3), .B1(data_in[14]), .B2(n1), .ZN(
        n113) );
  INV_X1 U35 ( .A(n112), .ZN(n29) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n3), .B1(data_in[15]), .B2(n4), .ZN(
        n112) );
  INV_X1 U37 ( .A(n111), .ZN(n28) );
  AOI22_X1 U38 ( .A1(\mem[0][16] ), .A2(n2), .B1(data_in[16]), .B2(n1), .ZN(
        n111) );
  INV_X1 U39 ( .A(n110), .ZN(n27) );
  AOI22_X1 U40 ( .A1(\mem[0][17] ), .A2(n2), .B1(data_in[17]), .B2(n4), .ZN(
        n110) );
  INV_X1 U41 ( .A(n109), .ZN(n26) );
  AOI22_X1 U42 ( .A1(\mem[0][18] ), .A2(n2), .B1(data_in[18]), .B2(n1), .ZN(
        n109) );
  INV_X1 U43 ( .A(n108), .ZN(n25) );
  AOI22_X1 U44 ( .A1(\mem[0][19] ), .A2(n2), .B1(data_in[19]), .B2(n1), .ZN(
        n108) );
  INV_X1 U45 ( .A(n107), .ZN(n24) );
  AOI22_X1 U46 ( .A1(\mem[0][20] ), .A2(n2), .B1(data_in[20]), .B2(n4), .ZN(
        n107) );
  INV_X1 U47 ( .A(n106), .ZN(n23) );
  AOI22_X1 U48 ( .A1(\mem[0][21] ), .A2(n2), .B1(data_in[21]), .B2(n4), .ZN(
        n106) );
  INV_X1 U49 ( .A(n105), .ZN(n22) );
  AOI22_X1 U50 ( .A1(\mem[0][22] ), .A2(n2), .B1(data_in[22]), .B2(n4), .ZN(
        n105) );
  INV_X1 U51 ( .A(n104), .ZN(n21) );
  AOI22_X1 U52 ( .A1(\mem[0][23] ), .A2(n2), .B1(data_in[23]), .B2(n4), .ZN(
        n104) );
  INV_X1 U53 ( .A(n103), .ZN(n20) );
  AOI22_X1 U54 ( .A1(\mem[0][24] ), .A2(n2), .B1(data_in[24]), .B2(n1), .ZN(
        n103) );
  INV_X1 U55 ( .A(n102), .ZN(n19) );
  AOI22_X1 U56 ( .A1(\mem[0][25] ), .A2(n2), .B1(data_in[25]), .B2(n1), .ZN(
        n102) );
  INV_X1 U57 ( .A(n101), .ZN(n18) );
  AOI22_X1 U58 ( .A1(\mem[0][26] ), .A2(n2), .B1(data_in[26]), .B2(n1), .ZN(
        n101) );
  INV_X1 U59 ( .A(n100), .ZN(n17) );
  AOI22_X1 U60 ( .A1(\mem[0][27] ), .A2(n2), .B1(data_in[27]), .B2(n1), .ZN(
        n100) );
  INV_X1 U61 ( .A(n99), .ZN(n16) );
  AOI22_X1 U62 ( .A1(\mem[0][28] ), .A2(n3), .B1(data_in[28]), .B2(n4), .ZN(
        n99) );
  INV_X1 U63 ( .A(n98), .ZN(n15) );
  AOI22_X1 U64 ( .A1(\mem[0][29] ), .A2(n2), .B1(data_in[29]), .B2(n1), .ZN(
        n98) );
  INV_X1 U65 ( .A(n97), .ZN(n14) );
  AOI22_X1 U66 ( .A1(\mem[0][30] ), .A2(n3), .B1(data_in[30]), .B2(n1), .ZN(
        n97) );
  INV_X1 U67 ( .A(n96), .ZN(n13) );
  AOI22_X1 U68 ( .A1(\mem[0][31] ), .A2(n2), .B1(data_in[31]), .B2(n1), .ZN(
        n96) );
  INV_X1 U69 ( .A(n118), .ZN(n35) );
  AOI22_X1 U70 ( .A1(\mem[0][9] ), .A2(n3), .B1(data_in[9]), .B2(n4), .ZN(n118) );
  INV_X1 U71 ( .A(n116), .ZN(n33) );
  AOI22_X1 U72 ( .A1(\mem[0][11] ), .A2(n3), .B1(data_in[11]), .B2(n1), .ZN(
        n116) );
  INV_X1 U73 ( .A(n95), .ZN(n12) );
  AOI22_X1 U74 ( .A1(\mem[0][32] ), .A2(n3), .B1(data_in[32]), .B2(n1), .ZN(
        n95) );
  INV_X1 U75 ( .A(n94), .ZN(n11) );
  AOI22_X1 U76 ( .A1(\mem[0][33] ), .A2(n2), .B1(data_in[33]), .B2(n1), .ZN(
        n94) );
  INV_X1 U77 ( .A(n93), .ZN(n10) );
  AOI22_X1 U78 ( .A1(\mem[0][34] ), .A2(n3), .B1(data_in[34]), .B2(n4), .ZN(
        n93) );
  INV_X1 U79 ( .A(n92), .ZN(n9) );
  AOI22_X1 U80 ( .A1(\mem[0][35] ), .A2(n2), .B1(data_in[35]), .B2(n1), .ZN(
        n92) );
  INV_X1 U81 ( .A(n91), .ZN(n8) );
  AOI22_X1 U82 ( .A1(\mem[0][36] ), .A2(n3), .B1(data_in[36]), .B2(n4), .ZN(
        n91) );
  INV_X1 U83 ( .A(n90), .ZN(n7) );
  AOI22_X1 U84 ( .A1(\mem[0][37] ), .A2(n2), .B1(data_in[37]), .B2(n1), .ZN(
        n90) );
  INV_X1 U85 ( .A(n89), .ZN(n6) );
  AOI22_X1 U86 ( .A1(\mem[0][38] ), .A2(n3), .B1(data_in[38]), .B2(n1), .ZN(
        n89) );
  INV_X1 U87 ( .A(n88), .ZN(n5) );
  AOI22_X1 U88 ( .A1(\mem[0][39] ), .A2(n2), .B1(data_in[39]), .B2(n4), .ZN(
        n88) );
endmodule


module memory_WIDTH40_SIZE1_LOGSIZE4_2 ( clk, data_in, data_out, addr, wr_en
 );
  input [39:0] data_in;
  output [39:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   \mem[0][39] , \mem[0][38] , \mem[0][37] , \mem[0][36] , \mem[0][35] ,
         \mem[0][34] , \mem[0][33] , \mem[0][32] , \mem[0][31] , \mem[0][30] ,
         \mem[0][29] , \mem[0][28] , \mem[0][27] , \mem[0][26] , \mem[0][25] ,
         \mem[0][24] , \mem[0][23] , \mem[0][22] , \mem[0][21] , \mem[0][20] ,
         \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] , \mem[0][15] ,
         \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] ,
         \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  DFF_X1 \mem_reg[0][39]  ( .D(n5), .CK(clk), .Q(\mem[0][39] ) );
  DFF_X1 \data_out_reg[39]  ( .D(\mem[0][39] ), .CK(clk), .Q(data_out[39]) );
  DFF_X1 \mem_reg[0][38]  ( .D(n6), .CK(clk), .Q(\mem[0][38] ) );
  DFF_X1 \data_out_reg[38]  ( .D(\mem[0][38] ), .CK(clk), .Q(data_out[38]) );
  DFF_X1 \mem_reg[0][37]  ( .D(n7), .CK(clk), .Q(\mem[0][37] ) );
  DFF_X1 \data_out_reg[37]  ( .D(\mem[0][37] ), .CK(clk), .Q(data_out[37]) );
  DFF_X1 \mem_reg[0][36]  ( .D(n8), .CK(clk), .Q(\mem[0][36] ) );
  DFF_X1 \data_out_reg[36]  ( .D(\mem[0][36] ), .CK(clk), .Q(data_out[36]) );
  DFF_X1 \mem_reg[0][35]  ( .D(n9), .CK(clk), .Q(\mem[0][35] ) );
  DFF_X1 \data_out_reg[35]  ( .D(\mem[0][35] ), .CK(clk), .Q(data_out[35]) );
  DFF_X1 \mem_reg[0][34]  ( .D(n10), .CK(clk), .Q(\mem[0][34] ) );
  DFF_X1 \data_out_reg[34]  ( .D(\mem[0][34] ), .CK(clk), .Q(data_out[34]) );
  DFF_X1 \mem_reg[0][33]  ( .D(n11), .CK(clk), .Q(\mem[0][33] ) );
  DFF_X1 \data_out_reg[33]  ( .D(\mem[0][33] ), .CK(clk), .Q(data_out[33]) );
  DFF_X1 \mem_reg[0][32]  ( .D(n12), .CK(clk), .Q(\mem[0][32] ) );
  DFF_X1 \data_out_reg[32]  ( .D(\mem[0][32] ), .CK(clk), .Q(data_out[32]) );
  DFF_X1 \mem_reg[0][31]  ( .D(n13), .CK(clk), .Q(\mem[0][31] ) );
  DFF_X1 \data_out_reg[31]  ( .D(\mem[0][31] ), .CK(clk), .Q(data_out[31]) );
  DFF_X1 \mem_reg[0][30]  ( .D(n14), .CK(clk), .Q(\mem[0][30] ) );
  DFF_X1 \data_out_reg[30]  ( .D(\mem[0][30] ), .CK(clk), .Q(data_out[30]) );
  DFF_X1 \mem_reg[0][29]  ( .D(n15), .CK(clk), .Q(\mem[0][29] ) );
  DFF_X1 \data_out_reg[29]  ( .D(\mem[0][29] ), .CK(clk), .Q(data_out[29]) );
  DFF_X1 \mem_reg[0][28]  ( .D(n16), .CK(clk), .Q(\mem[0][28] ) );
  DFF_X1 \data_out_reg[28]  ( .D(\mem[0][28] ), .CK(clk), .Q(data_out[28]) );
  DFF_X1 \mem_reg[0][27]  ( .D(n17), .CK(clk), .Q(\mem[0][27] ) );
  DFF_X1 \data_out_reg[27]  ( .D(\mem[0][27] ), .CK(clk), .Q(data_out[27]) );
  DFF_X1 \mem_reg[0][26]  ( .D(n18), .CK(clk), .Q(\mem[0][26] ) );
  DFF_X1 \data_out_reg[26]  ( .D(\mem[0][26] ), .CK(clk), .Q(data_out[26]) );
  DFF_X1 \mem_reg[0][25]  ( .D(n19), .CK(clk), .Q(\mem[0][25] ) );
  DFF_X1 \data_out_reg[25]  ( .D(\mem[0][25] ), .CK(clk), .Q(data_out[25]) );
  DFF_X1 \mem_reg[0][24]  ( .D(n20), .CK(clk), .Q(\mem[0][24] ) );
  DFF_X1 \data_out_reg[24]  ( .D(\mem[0][24] ), .CK(clk), .Q(data_out[24]) );
  DFF_X1 \mem_reg[0][23]  ( .D(n21), .CK(clk), .Q(\mem[0][23] ) );
  DFF_X1 \data_out_reg[23]  ( .D(\mem[0][23] ), .CK(clk), .Q(data_out[23]) );
  DFF_X1 \mem_reg[0][22]  ( .D(n22), .CK(clk), .Q(\mem[0][22] ) );
  DFF_X1 \data_out_reg[22]  ( .D(\mem[0][22] ), .CK(clk), .Q(data_out[22]) );
  DFF_X1 \mem_reg[0][21]  ( .D(n23), .CK(clk), .Q(\mem[0][21] ) );
  DFF_X1 \data_out_reg[21]  ( .D(\mem[0][21] ), .CK(clk), .Q(data_out[21]) );
  DFF_X1 \mem_reg[0][20]  ( .D(n24), .CK(clk), .Q(\mem[0][20] ) );
  DFF_X1 \data_out_reg[20]  ( .D(\mem[0][20] ), .CK(clk), .Q(data_out[20]) );
  DFF_X1 \mem_reg[0][19]  ( .D(n25), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \data_out_reg[19]  ( .D(\mem[0][19] ), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \mem_reg[0][18]  ( .D(n26), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \data_out_reg[18]  ( .D(\mem[0][18] ), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \mem_reg[0][17]  ( .D(n27), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \data_out_reg[17]  ( .D(\mem[0][17] ), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \mem_reg[0][16]  ( .D(n28), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \data_out_reg[16]  ( .D(\mem[0][16] ), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \mem_reg[0][15]  ( .D(n29), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n30), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n31), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n32), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n33), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n34), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n35), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n36), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n37), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n38), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n39), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n40), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n41), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n42), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n44), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n85), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  AND3_X1 U3 ( .A1(wr_en), .A2(n86), .A3(n87), .ZN(n1) );
  INV_X1 U4 ( .A(n1), .ZN(n3) );
  INV_X1 U5 ( .A(n1), .ZN(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n4) );
  INV_X1 U7 ( .A(addr[0]), .ZN(n86) );
  NOR3_X1 U8 ( .A1(addr[1]), .A2(addr[3]), .A3(addr[2]), .ZN(n87) );
  INV_X1 U9 ( .A(n127), .ZN(n85) );
  AOI22_X1 U10 ( .A1(\mem[0][0] ), .A2(n3), .B1(data_in[0]), .B2(n4), .ZN(n127) );
  INV_X1 U11 ( .A(n126), .ZN(n44) );
  AOI22_X1 U12 ( .A1(\mem[0][1] ), .A2(n2), .B1(data_in[1]), .B2(n4), .ZN(n126) );
  INV_X1 U13 ( .A(n125), .ZN(n42) );
  AOI22_X1 U14 ( .A1(\mem[0][2] ), .A2(n2), .B1(data_in[2]), .B2(n4), .ZN(n125) );
  INV_X1 U15 ( .A(n124), .ZN(n41) );
  AOI22_X1 U16 ( .A1(\mem[0][3] ), .A2(n3), .B1(data_in[3]), .B2(n1), .ZN(n124) );
  INV_X1 U17 ( .A(n123), .ZN(n40) );
  AOI22_X1 U18 ( .A1(\mem[0][4] ), .A2(n3), .B1(data_in[4]), .B2(n4), .ZN(n123) );
  INV_X1 U19 ( .A(n122), .ZN(n39) );
  AOI22_X1 U20 ( .A1(\mem[0][5] ), .A2(n3), .B1(data_in[5]), .B2(n4), .ZN(n122) );
  INV_X1 U21 ( .A(n121), .ZN(n38) );
  AOI22_X1 U22 ( .A1(\mem[0][6] ), .A2(n3), .B1(data_in[6]), .B2(n4), .ZN(n121) );
  INV_X1 U23 ( .A(n120), .ZN(n37) );
  AOI22_X1 U24 ( .A1(\mem[0][7] ), .A2(n3), .B1(data_in[7]), .B2(n1), .ZN(n120) );
  INV_X1 U25 ( .A(n119), .ZN(n36) );
  AOI22_X1 U26 ( .A1(\mem[0][8] ), .A2(n3), .B1(data_in[8]), .B2(n4), .ZN(n119) );
  INV_X1 U27 ( .A(n118), .ZN(n35) );
  AOI22_X1 U28 ( .A1(\mem[0][9] ), .A2(n3), .B1(data_in[9]), .B2(n4), .ZN(n118) );
  INV_X1 U29 ( .A(n117), .ZN(n34) );
  AOI22_X1 U30 ( .A1(\mem[0][10] ), .A2(n3), .B1(data_in[10]), .B2(n4), .ZN(
        n117) );
  INV_X1 U31 ( .A(n115), .ZN(n32) );
  AOI22_X1 U32 ( .A1(\mem[0][12] ), .A2(n3), .B1(data_in[12]), .B2(n1), .ZN(
        n115) );
  INV_X1 U33 ( .A(n114), .ZN(n31) );
  AOI22_X1 U34 ( .A1(\mem[0][13] ), .A2(n3), .B1(data_in[13]), .B2(n1), .ZN(
        n114) );
  INV_X1 U35 ( .A(n113), .ZN(n30) );
  AOI22_X1 U36 ( .A1(\mem[0][14] ), .A2(n3), .B1(data_in[14]), .B2(n1), .ZN(
        n113) );
  INV_X1 U37 ( .A(n112), .ZN(n29) );
  AOI22_X1 U38 ( .A1(\mem[0][15] ), .A2(n3), .B1(data_in[15]), .B2(n1), .ZN(
        n112) );
  INV_X1 U39 ( .A(n111), .ZN(n28) );
  AOI22_X1 U40 ( .A1(\mem[0][16] ), .A2(n2), .B1(data_in[16]), .B2(n1), .ZN(
        n111) );
  INV_X1 U41 ( .A(n110), .ZN(n27) );
  AOI22_X1 U42 ( .A1(\mem[0][17] ), .A2(n2), .B1(data_in[17]), .B2(n4), .ZN(
        n110) );
  INV_X1 U43 ( .A(n109), .ZN(n26) );
  AOI22_X1 U44 ( .A1(\mem[0][18] ), .A2(n2), .B1(data_in[18]), .B2(n1), .ZN(
        n109) );
  INV_X1 U45 ( .A(n108), .ZN(n25) );
  AOI22_X1 U46 ( .A1(\mem[0][19] ), .A2(n2), .B1(data_in[19]), .B2(n4), .ZN(
        n108) );
  INV_X1 U47 ( .A(n107), .ZN(n24) );
  AOI22_X1 U48 ( .A1(\mem[0][20] ), .A2(n2), .B1(data_in[20]), .B2(n1), .ZN(
        n107) );
  INV_X1 U49 ( .A(n106), .ZN(n23) );
  AOI22_X1 U50 ( .A1(\mem[0][21] ), .A2(n2), .B1(data_in[21]), .B2(n1), .ZN(
        n106) );
  INV_X1 U51 ( .A(n105), .ZN(n22) );
  AOI22_X1 U52 ( .A1(\mem[0][22] ), .A2(n2), .B1(data_in[22]), .B2(n4), .ZN(
        n105) );
  INV_X1 U53 ( .A(n104), .ZN(n21) );
  AOI22_X1 U54 ( .A1(\mem[0][23] ), .A2(n2), .B1(data_in[23]), .B2(n1), .ZN(
        n104) );
  INV_X1 U55 ( .A(n103), .ZN(n20) );
  AOI22_X1 U56 ( .A1(\mem[0][24] ), .A2(n2), .B1(data_in[24]), .B2(n1), .ZN(
        n103) );
  INV_X1 U57 ( .A(n102), .ZN(n19) );
  AOI22_X1 U58 ( .A1(\mem[0][25] ), .A2(n2), .B1(data_in[25]), .B2(n1), .ZN(
        n102) );
  INV_X1 U59 ( .A(n101), .ZN(n18) );
  AOI22_X1 U60 ( .A1(\mem[0][26] ), .A2(n2), .B1(data_in[26]), .B2(n1), .ZN(
        n101) );
  INV_X1 U61 ( .A(n100), .ZN(n17) );
  AOI22_X1 U62 ( .A1(\mem[0][27] ), .A2(n2), .B1(data_in[27]), .B2(n4), .ZN(
        n100) );
  INV_X1 U63 ( .A(n99), .ZN(n16) );
  AOI22_X1 U64 ( .A1(\mem[0][28] ), .A2(n3), .B1(data_in[28]), .B2(n1), .ZN(
        n99) );
  INV_X1 U65 ( .A(n98), .ZN(n15) );
  AOI22_X1 U66 ( .A1(\mem[0][29] ), .A2(n2), .B1(data_in[29]), .B2(n4), .ZN(
        n98) );
  INV_X1 U67 ( .A(n97), .ZN(n14) );
  AOI22_X1 U68 ( .A1(\mem[0][30] ), .A2(n3), .B1(data_in[30]), .B2(n1), .ZN(
        n97) );
  INV_X1 U69 ( .A(n96), .ZN(n13) );
  AOI22_X1 U70 ( .A1(\mem[0][31] ), .A2(n2), .B1(data_in[31]), .B2(n1), .ZN(
        n96) );
  INV_X1 U71 ( .A(n116), .ZN(n33) );
  AOI22_X1 U72 ( .A1(\mem[0][11] ), .A2(n3), .B1(data_in[11]), .B2(n4), .ZN(
        n116) );
  INV_X1 U73 ( .A(n95), .ZN(n12) );
  AOI22_X1 U74 ( .A1(\mem[0][32] ), .A2(n3), .B1(data_in[32]), .B2(n1), .ZN(
        n95) );
  INV_X1 U75 ( .A(n94), .ZN(n11) );
  AOI22_X1 U76 ( .A1(\mem[0][33] ), .A2(n2), .B1(data_in[33]), .B2(n4), .ZN(
        n94) );
  INV_X1 U77 ( .A(n93), .ZN(n10) );
  AOI22_X1 U78 ( .A1(\mem[0][34] ), .A2(n3), .B1(data_in[34]), .B2(n1), .ZN(
        n93) );
  INV_X1 U79 ( .A(n92), .ZN(n9) );
  AOI22_X1 U80 ( .A1(\mem[0][35] ), .A2(n2), .B1(data_in[35]), .B2(n1), .ZN(
        n92) );
  INV_X1 U81 ( .A(n91), .ZN(n8) );
  AOI22_X1 U82 ( .A1(\mem[0][36] ), .A2(n3), .B1(data_in[36]), .B2(n1), .ZN(
        n91) );
  INV_X1 U83 ( .A(n90), .ZN(n7) );
  AOI22_X1 U84 ( .A1(\mem[0][37] ), .A2(n2), .B1(data_in[37]), .B2(n1), .ZN(
        n90) );
  INV_X1 U85 ( .A(n89), .ZN(n6) );
  AOI22_X1 U86 ( .A1(\mem[0][38] ), .A2(n3), .B1(data_in[38]), .B2(n1), .ZN(
        n89) );
  INV_X1 U87 ( .A(n88), .ZN(n5) );
  AOI22_X1 U88 ( .A1(\mem[0][39] ), .A2(n2), .B1(data_in[39]), .B2(n4), .ZN(
        n88) );
endmodule


module memory_WIDTH40_SIZE1_LOGSIZE4_1 ( clk, data_in, data_out, addr, wr_en
 );
  input [39:0] data_in;
  output [39:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   \mem[0][39] , \mem[0][38] , \mem[0][37] , \mem[0][36] , \mem[0][35] ,
         \mem[0][34] , \mem[0][33] , \mem[0][32] , \mem[0][31] , \mem[0][30] ,
         \mem[0][29] , \mem[0][28] , \mem[0][27] , \mem[0][26] , \mem[0][25] ,
         \mem[0][24] , \mem[0][23] , \mem[0][22] , \mem[0][21] , \mem[0][20] ,
         \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] , \mem[0][15] ,
         \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] ,
         \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  DFF_X1 \mem_reg[0][39]  ( .D(n5), .CK(clk), .Q(\mem[0][39] ) );
  DFF_X1 \data_out_reg[39]  ( .D(\mem[0][39] ), .CK(clk), .Q(data_out[39]) );
  DFF_X1 \mem_reg[0][38]  ( .D(n6), .CK(clk), .Q(\mem[0][38] ) );
  DFF_X1 \data_out_reg[38]  ( .D(\mem[0][38] ), .CK(clk), .Q(data_out[38]) );
  DFF_X1 \mem_reg[0][37]  ( .D(n7), .CK(clk), .Q(\mem[0][37] ) );
  DFF_X1 \data_out_reg[37]  ( .D(\mem[0][37] ), .CK(clk), .Q(data_out[37]) );
  DFF_X1 \mem_reg[0][36]  ( .D(n8), .CK(clk), .Q(\mem[0][36] ) );
  DFF_X1 \data_out_reg[36]  ( .D(\mem[0][36] ), .CK(clk), .Q(data_out[36]) );
  DFF_X1 \mem_reg[0][35]  ( .D(n9), .CK(clk), .Q(\mem[0][35] ) );
  DFF_X1 \data_out_reg[35]  ( .D(\mem[0][35] ), .CK(clk), .Q(data_out[35]) );
  DFF_X1 \mem_reg[0][34]  ( .D(n10), .CK(clk), .Q(\mem[0][34] ) );
  DFF_X1 \data_out_reg[34]  ( .D(\mem[0][34] ), .CK(clk), .Q(data_out[34]) );
  DFF_X1 \mem_reg[0][33]  ( .D(n11), .CK(clk), .Q(\mem[0][33] ) );
  DFF_X1 \data_out_reg[33]  ( .D(\mem[0][33] ), .CK(clk), .Q(data_out[33]) );
  DFF_X1 \mem_reg[0][32]  ( .D(n12), .CK(clk), .Q(\mem[0][32] ) );
  DFF_X1 \data_out_reg[32]  ( .D(\mem[0][32] ), .CK(clk), .Q(data_out[32]) );
  DFF_X1 \mem_reg[0][31]  ( .D(n13), .CK(clk), .Q(\mem[0][31] ) );
  DFF_X1 \data_out_reg[31]  ( .D(\mem[0][31] ), .CK(clk), .Q(data_out[31]) );
  DFF_X1 \mem_reg[0][30]  ( .D(n14), .CK(clk), .Q(\mem[0][30] ) );
  DFF_X1 \data_out_reg[30]  ( .D(\mem[0][30] ), .CK(clk), .Q(data_out[30]) );
  DFF_X1 \mem_reg[0][29]  ( .D(n15), .CK(clk), .Q(\mem[0][29] ) );
  DFF_X1 \data_out_reg[29]  ( .D(\mem[0][29] ), .CK(clk), .Q(data_out[29]) );
  DFF_X1 \mem_reg[0][28]  ( .D(n16), .CK(clk), .Q(\mem[0][28] ) );
  DFF_X1 \data_out_reg[28]  ( .D(\mem[0][28] ), .CK(clk), .Q(data_out[28]) );
  DFF_X1 \mem_reg[0][27]  ( .D(n17), .CK(clk), .Q(\mem[0][27] ) );
  DFF_X1 \data_out_reg[27]  ( .D(\mem[0][27] ), .CK(clk), .Q(data_out[27]) );
  DFF_X1 \mem_reg[0][26]  ( .D(n18), .CK(clk), .Q(\mem[0][26] ) );
  DFF_X1 \data_out_reg[26]  ( .D(\mem[0][26] ), .CK(clk), .Q(data_out[26]) );
  DFF_X1 \mem_reg[0][25]  ( .D(n19), .CK(clk), .Q(\mem[0][25] ) );
  DFF_X1 \data_out_reg[25]  ( .D(\mem[0][25] ), .CK(clk), .Q(data_out[25]) );
  DFF_X1 \mem_reg[0][24]  ( .D(n20), .CK(clk), .Q(\mem[0][24] ) );
  DFF_X1 \data_out_reg[24]  ( .D(\mem[0][24] ), .CK(clk), .Q(data_out[24]) );
  DFF_X1 \mem_reg[0][23]  ( .D(n21), .CK(clk), .Q(\mem[0][23] ) );
  DFF_X1 \data_out_reg[23]  ( .D(\mem[0][23] ), .CK(clk), .Q(data_out[23]) );
  DFF_X1 \mem_reg[0][22]  ( .D(n22), .CK(clk), .Q(\mem[0][22] ) );
  DFF_X1 \data_out_reg[22]  ( .D(\mem[0][22] ), .CK(clk), .Q(data_out[22]) );
  DFF_X1 \mem_reg[0][21]  ( .D(n23), .CK(clk), .Q(\mem[0][21] ) );
  DFF_X1 \data_out_reg[21]  ( .D(\mem[0][21] ), .CK(clk), .Q(data_out[21]) );
  DFF_X1 \mem_reg[0][20]  ( .D(n24), .CK(clk), .Q(\mem[0][20] ) );
  DFF_X1 \data_out_reg[20]  ( .D(\mem[0][20] ), .CK(clk), .Q(data_out[20]) );
  DFF_X1 \mem_reg[0][19]  ( .D(n25), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \data_out_reg[19]  ( .D(\mem[0][19] ), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \mem_reg[0][18]  ( .D(n26), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \data_out_reg[18]  ( .D(\mem[0][18] ), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \mem_reg[0][17]  ( .D(n27), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \data_out_reg[17]  ( .D(\mem[0][17] ), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \mem_reg[0][16]  ( .D(n28), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \data_out_reg[16]  ( .D(\mem[0][16] ), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \mem_reg[0][15]  ( .D(n29), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n30), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n31), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n32), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n33), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n34), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n35), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n36), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n37), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n38), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n39), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n40), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n41), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n42), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n44), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n85), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  AND3_X1 U3 ( .A1(wr_en), .A2(n86), .A3(n87), .ZN(n1) );
  INV_X1 U4 ( .A(n1), .ZN(n3) );
  INV_X1 U5 ( .A(n1), .ZN(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n4) );
  INV_X1 U7 ( .A(addr[0]), .ZN(n86) );
  NOR3_X1 U8 ( .A1(addr[1]), .A2(addr[3]), .A3(addr[2]), .ZN(n87) );
  INV_X1 U9 ( .A(n127), .ZN(n85) );
  AOI22_X1 U10 ( .A1(\mem[0][0] ), .A2(n3), .B1(data_in[0]), .B2(n1), .ZN(n127) );
  INV_X1 U11 ( .A(n126), .ZN(n44) );
  AOI22_X1 U12 ( .A1(\mem[0][1] ), .A2(n2), .B1(data_in[1]), .B2(n4), .ZN(n126) );
  INV_X1 U13 ( .A(n125), .ZN(n42) );
  AOI22_X1 U14 ( .A1(\mem[0][2] ), .A2(n2), .B1(data_in[2]), .B2(n1), .ZN(n125) );
  INV_X1 U15 ( .A(n124), .ZN(n41) );
  AOI22_X1 U16 ( .A1(\mem[0][3] ), .A2(n3), .B1(data_in[3]), .B2(n1), .ZN(n124) );
  INV_X1 U17 ( .A(n123), .ZN(n40) );
  AOI22_X1 U18 ( .A1(\mem[0][4] ), .A2(n3), .B1(data_in[4]), .B2(n4), .ZN(n123) );
  INV_X1 U19 ( .A(n122), .ZN(n39) );
  AOI22_X1 U20 ( .A1(\mem[0][5] ), .A2(n3), .B1(data_in[5]), .B2(n4), .ZN(n122) );
  INV_X1 U21 ( .A(n121), .ZN(n38) );
  AOI22_X1 U22 ( .A1(\mem[0][6] ), .A2(n3), .B1(data_in[6]), .B2(n1), .ZN(n121) );
  INV_X1 U23 ( .A(n120), .ZN(n37) );
  AOI22_X1 U24 ( .A1(\mem[0][7] ), .A2(n3), .B1(data_in[7]), .B2(n4), .ZN(n120) );
  INV_X1 U25 ( .A(n119), .ZN(n36) );
  AOI22_X1 U26 ( .A1(\mem[0][8] ), .A2(n3), .B1(data_in[8]), .B2(n1), .ZN(n119) );
  INV_X1 U27 ( .A(n118), .ZN(n35) );
  AOI22_X1 U28 ( .A1(\mem[0][9] ), .A2(n3), .B1(data_in[9]), .B2(n1), .ZN(n118) );
  INV_X1 U29 ( .A(n117), .ZN(n34) );
  AOI22_X1 U30 ( .A1(\mem[0][10] ), .A2(n3), .B1(data_in[10]), .B2(n4), .ZN(
        n117) );
  INV_X1 U31 ( .A(n115), .ZN(n32) );
  AOI22_X1 U32 ( .A1(\mem[0][12] ), .A2(n3), .B1(data_in[12]), .B2(n1), .ZN(
        n115) );
  INV_X1 U33 ( .A(n114), .ZN(n31) );
  AOI22_X1 U34 ( .A1(\mem[0][13] ), .A2(n3), .B1(data_in[13]), .B2(n4), .ZN(
        n114) );
  INV_X1 U35 ( .A(n113), .ZN(n30) );
  AOI22_X1 U36 ( .A1(\mem[0][14] ), .A2(n3), .B1(data_in[14]), .B2(n1), .ZN(
        n113) );
  INV_X1 U37 ( .A(n112), .ZN(n29) );
  AOI22_X1 U38 ( .A1(\mem[0][15] ), .A2(n3), .B1(data_in[15]), .B2(n4), .ZN(
        n112) );
  INV_X1 U39 ( .A(n111), .ZN(n28) );
  AOI22_X1 U40 ( .A1(\mem[0][16] ), .A2(n2), .B1(data_in[16]), .B2(n1), .ZN(
        n111) );
  INV_X1 U41 ( .A(n110), .ZN(n27) );
  AOI22_X1 U42 ( .A1(\mem[0][17] ), .A2(n2), .B1(data_in[17]), .B2(n4), .ZN(
        n110) );
  INV_X1 U43 ( .A(n109), .ZN(n26) );
  AOI22_X1 U44 ( .A1(\mem[0][18] ), .A2(n2), .B1(data_in[18]), .B2(n1), .ZN(
        n109) );
  INV_X1 U45 ( .A(n108), .ZN(n25) );
  AOI22_X1 U46 ( .A1(\mem[0][19] ), .A2(n2), .B1(data_in[19]), .B2(n1), .ZN(
        n108) );
  INV_X1 U47 ( .A(n107), .ZN(n24) );
  AOI22_X1 U48 ( .A1(\mem[0][20] ), .A2(n2), .B1(data_in[20]), .B2(n4), .ZN(
        n107) );
  INV_X1 U49 ( .A(n106), .ZN(n23) );
  AOI22_X1 U50 ( .A1(\mem[0][21] ), .A2(n2), .B1(data_in[21]), .B2(n4), .ZN(
        n106) );
  INV_X1 U51 ( .A(n105), .ZN(n22) );
  AOI22_X1 U52 ( .A1(\mem[0][22] ), .A2(n2), .B1(data_in[22]), .B2(n1), .ZN(
        n105) );
  INV_X1 U53 ( .A(n104), .ZN(n21) );
  AOI22_X1 U54 ( .A1(\mem[0][23] ), .A2(n2), .B1(data_in[23]), .B2(n4), .ZN(
        n104) );
  INV_X1 U55 ( .A(n103), .ZN(n20) );
  AOI22_X1 U56 ( .A1(\mem[0][24] ), .A2(n2), .B1(data_in[24]), .B2(n1), .ZN(
        n103) );
  INV_X1 U57 ( .A(n102), .ZN(n19) );
  AOI22_X1 U58 ( .A1(\mem[0][25] ), .A2(n2), .B1(data_in[25]), .B2(n1), .ZN(
        n102) );
  INV_X1 U59 ( .A(n101), .ZN(n18) );
  AOI22_X1 U60 ( .A1(\mem[0][26] ), .A2(n2), .B1(data_in[26]), .B2(n4), .ZN(
        n101) );
  INV_X1 U61 ( .A(n100), .ZN(n17) );
  AOI22_X1 U62 ( .A1(\mem[0][27] ), .A2(n2), .B1(data_in[27]), .B2(n1), .ZN(
        n100) );
  INV_X1 U63 ( .A(n99), .ZN(n16) );
  AOI22_X1 U64 ( .A1(\mem[0][28] ), .A2(n3), .B1(data_in[28]), .B2(n4), .ZN(
        n99) );
  INV_X1 U65 ( .A(n98), .ZN(n15) );
  AOI22_X1 U66 ( .A1(\mem[0][29] ), .A2(n2), .B1(data_in[29]), .B2(n4), .ZN(
        n98) );
  INV_X1 U67 ( .A(n97), .ZN(n14) );
  AOI22_X1 U68 ( .A1(\mem[0][30] ), .A2(n3), .B1(data_in[30]), .B2(n4), .ZN(
        n97) );
  INV_X1 U69 ( .A(n96), .ZN(n13) );
  AOI22_X1 U70 ( .A1(\mem[0][31] ), .A2(n2), .B1(data_in[31]), .B2(n4), .ZN(
        n96) );
  INV_X1 U71 ( .A(n116), .ZN(n33) );
  AOI22_X1 U72 ( .A1(\mem[0][11] ), .A2(n3), .B1(data_in[11]), .B2(n1), .ZN(
        n116) );
  INV_X1 U73 ( .A(n95), .ZN(n12) );
  AOI22_X1 U74 ( .A1(\mem[0][32] ), .A2(n3), .B1(data_in[32]), .B2(n1), .ZN(
        n95) );
  INV_X1 U75 ( .A(n94), .ZN(n11) );
  AOI22_X1 U76 ( .A1(\mem[0][33] ), .A2(n2), .B1(data_in[33]), .B2(n1), .ZN(
        n94) );
  INV_X1 U77 ( .A(n93), .ZN(n10) );
  AOI22_X1 U78 ( .A1(\mem[0][34] ), .A2(n3), .B1(data_in[34]), .B2(n1), .ZN(
        n93) );
  INV_X1 U79 ( .A(n92), .ZN(n9) );
  AOI22_X1 U80 ( .A1(\mem[0][35] ), .A2(n2), .B1(data_in[35]), .B2(n4), .ZN(
        n92) );
  INV_X1 U81 ( .A(n91), .ZN(n8) );
  AOI22_X1 U82 ( .A1(\mem[0][36] ), .A2(n3), .B1(data_in[36]), .B2(n4), .ZN(
        n91) );
  INV_X1 U83 ( .A(n90), .ZN(n7) );
  AOI22_X1 U84 ( .A1(\mem[0][37] ), .A2(n2), .B1(data_in[37]), .B2(n4), .ZN(
        n90) );
  INV_X1 U85 ( .A(n89), .ZN(n6) );
  AOI22_X1 U86 ( .A1(\mem[0][38] ), .A2(n3), .B1(data_in[38]), .B2(n4), .ZN(
        n89) );
  INV_X1 U87 ( .A(n88), .ZN(n5) );
  AOI22_X1 U88 ( .A1(\mem[0][39] ), .A2(n2), .B1(data_in[39]), .B2(n4), .ZN(
        n88) );
endmodule


module memory_WIDTH40_SIZE1_LOGSIZE4_0 ( clk, data_in, data_out, addr, wr_en
 );
  input [39:0] data_in;
  output [39:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   \mem[0][39] , \mem[0][38] , \mem[0][37] , \mem[0][36] , \mem[0][35] ,
         \mem[0][34] , \mem[0][33] , \mem[0][32] , \mem[0][31] , \mem[0][30] ,
         \mem[0][29] , \mem[0][28] , \mem[0][27] , \mem[0][26] , \mem[0][25] ,
         \mem[0][24] , \mem[0][23] , \mem[0][22] , \mem[0][21] , \mem[0][20] ,
         \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] , \mem[0][15] ,
         \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] ,
         \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  DFF_X1 \mem_reg[0][39]  ( .D(n5), .CK(clk), .Q(\mem[0][39] ) );
  DFF_X1 \data_out_reg[39]  ( .D(\mem[0][39] ), .CK(clk), .Q(data_out[39]) );
  DFF_X1 \mem_reg[0][38]  ( .D(n6), .CK(clk), .Q(\mem[0][38] ) );
  DFF_X1 \data_out_reg[38]  ( .D(\mem[0][38] ), .CK(clk), .Q(data_out[38]) );
  DFF_X1 \mem_reg[0][37]  ( .D(n7), .CK(clk), .Q(\mem[0][37] ) );
  DFF_X1 \data_out_reg[37]  ( .D(\mem[0][37] ), .CK(clk), .Q(data_out[37]) );
  DFF_X1 \mem_reg[0][36]  ( .D(n8), .CK(clk), .Q(\mem[0][36] ) );
  DFF_X1 \data_out_reg[36]  ( .D(\mem[0][36] ), .CK(clk), .Q(data_out[36]) );
  DFF_X1 \mem_reg[0][35]  ( .D(n9), .CK(clk), .Q(\mem[0][35] ) );
  DFF_X1 \data_out_reg[35]  ( .D(\mem[0][35] ), .CK(clk), .Q(data_out[35]) );
  DFF_X1 \mem_reg[0][34]  ( .D(n10), .CK(clk), .Q(\mem[0][34] ) );
  DFF_X1 \data_out_reg[34]  ( .D(\mem[0][34] ), .CK(clk), .Q(data_out[34]) );
  DFF_X1 \mem_reg[0][33]  ( .D(n11), .CK(clk), .Q(\mem[0][33] ) );
  DFF_X1 \data_out_reg[33]  ( .D(\mem[0][33] ), .CK(clk), .Q(data_out[33]) );
  DFF_X1 \mem_reg[0][32]  ( .D(n12), .CK(clk), .Q(\mem[0][32] ) );
  DFF_X1 \data_out_reg[32]  ( .D(\mem[0][32] ), .CK(clk), .Q(data_out[32]) );
  DFF_X1 \mem_reg[0][31]  ( .D(n13), .CK(clk), .Q(\mem[0][31] ) );
  DFF_X1 \data_out_reg[31]  ( .D(\mem[0][31] ), .CK(clk), .Q(data_out[31]) );
  DFF_X1 \mem_reg[0][30]  ( .D(n14), .CK(clk), .Q(\mem[0][30] ) );
  DFF_X1 \data_out_reg[30]  ( .D(\mem[0][30] ), .CK(clk), .Q(data_out[30]) );
  DFF_X1 \mem_reg[0][29]  ( .D(n15), .CK(clk), .Q(\mem[0][29] ) );
  DFF_X1 \data_out_reg[29]  ( .D(\mem[0][29] ), .CK(clk), .Q(data_out[29]) );
  DFF_X1 \mem_reg[0][28]  ( .D(n16), .CK(clk), .Q(\mem[0][28] ) );
  DFF_X1 \data_out_reg[28]  ( .D(\mem[0][28] ), .CK(clk), .Q(data_out[28]) );
  DFF_X1 \mem_reg[0][27]  ( .D(n17), .CK(clk), .Q(\mem[0][27] ) );
  DFF_X1 \data_out_reg[27]  ( .D(\mem[0][27] ), .CK(clk), .Q(data_out[27]) );
  DFF_X1 \mem_reg[0][26]  ( .D(n18), .CK(clk), .Q(\mem[0][26] ) );
  DFF_X1 \data_out_reg[26]  ( .D(\mem[0][26] ), .CK(clk), .Q(data_out[26]) );
  DFF_X1 \mem_reg[0][25]  ( .D(n19), .CK(clk), .Q(\mem[0][25] ) );
  DFF_X1 \data_out_reg[25]  ( .D(\mem[0][25] ), .CK(clk), .Q(data_out[25]) );
  DFF_X1 \mem_reg[0][24]  ( .D(n20), .CK(clk), .Q(\mem[0][24] ) );
  DFF_X1 \data_out_reg[24]  ( .D(\mem[0][24] ), .CK(clk), .Q(data_out[24]) );
  DFF_X1 \mem_reg[0][23]  ( .D(n21), .CK(clk), .Q(\mem[0][23] ) );
  DFF_X1 \data_out_reg[23]  ( .D(\mem[0][23] ), .CK(clk), .Q(data_out[23]) );
  DFF_X1 \mem_reg[0][22]  ( .D(n22), .CK(clk), .Q(\mem[0][22] ) );
  DFF_X1 \data_out_reg[22]  ( .D(\mem[0][22] ), .CK(clk), .Q(data_out[22]) );
  DFF_X1 \mem_reg[0][21]  ( .D(n23), .CK(clk), .Q(\mem[0][21] ) );
  DFF_X1 \data_out_reg[21]  ( .D(\mem[0][21] ), .CK(clk), .Q(data_out[21]) );
  DFF_X1 \mem_reg[0][20]  ( .D(n24), .CK(clk), .Q(\mem[0][20] ) );
  DFF_X1 \data_out_reg[20]  ( .D(\mem[0][20] ), .CK(clk), .Q(data_out[20]) );
  DFF_X1 \mem_reg[0][19]  ( .D(n25), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \data_out_reg[19]  ( .D(\mem[0][19] ), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \mem_reg[0][18]  ( .D(n26), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \data_out_reg[18]  ( .D(\mem[0][18] ), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \mem_reg[0][17]  ( .D(n27), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \data_out_reg[17]  ( .D(\mem[0][17] ), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \mem_reg[0][16]  ( .D(n28), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \data_out_reg[16]  ( .D(\mem[0][16] ), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \mem_reg[0][15]  ( .D(n29), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \data_out_reg[15]  ( .D(\mem[0][15] ), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \mem_reg[0][14]  ( .D(n30), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \data_out_reg[14]  ( .D(\mem[0][14] ), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \mem_reg[0][13]  ( .D(n31), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \data_out_reg[13]  ( .D(\mem[0][13] ), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \mem_reg[0][12]  ( .D(n32), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \data_out_reg[12]  ( .D(\mem[0][12] ), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \mem_reg[0][11]  ( .D(n33), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \data_out_reg[11]  ( .D(\mem[0][11] ), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \mem_reg[0][10]  ( .D(n34), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \data_out_reg[10]  ( .D(\mem[0][10] ), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[0][9]  ( .D(n35), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \data_out_reg[9]  ( .D(\mem[0][9] ), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \mem_reg[0][8]  ( .D(n36), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \data_out_reg[8]  ( .D(\mem[0][8] ), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \mem_reg[0][7]  ( .D(n37), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \data_out_reg[7]  ( .D(\mem[0][7] ), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \mem_reg[0][6]  ( .D(n38), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \data_out_reg[6]  ( .D(\mem[0][6] ), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[0][5]  ( .D(n39), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \data_out_reg[5]  ( .D(\mem[0][5] ), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \mem_reg[0][4]  ( .D(n40), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \data_out_reg[4]  ( .D(\mem[0][4] ), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[0][3]  ( .D(n41), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \data_out_reg[3]  ( .D(\mem[0][3] ), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[0][2]  ( .D(n42), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \data_out_reg[2]  ( .D(\mem[0][2] ), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[0][1]  ( .D(n44), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \data_out_reg[1]  ( .D(\mem[0][1] ), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[0][0]  ( .D(n85), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[0]  ( .D(\mem[0][0] ), .CK(clk), .Q(data_out[0]) );
  AND3_X1 U3 ( .A1(wr_en), .A2(n86), .A3(n87), .ZN(n1) );
  INV_X1 U4 ( .A(n1), .ZN(n3) );
  INV_X1 U5 ( .A(n1), .ZN(n2) );
  BUF_X1 U6 ( .A(n1), .Z(n4) );
  INV_X1 U7 ( .A(addr[0]), .ZN(n86) );
  NOR3_X1 U8 ( .A1(addr[1]), .A2(addr[3]), .A3(addr[2]), .ZN(n87) );
  INV_X1 U9 ( .A(n127), .ZN(n85) );
  AOI22_X1 U10 ( .A1(\mem[0][0] ), .A2(n3), .B1(data_in[0]), .B2(n4), .ZN(n127) );
  INV_X1 U11 ( .A(n126), .ZN(n44) );
  AOI22_X1 U12 ( .A1(\mem[0][1] ), .A2(n2), .B1(data_in[1]), .B2(n4), .ZN(n126) );
  INV_X1 U13 ( .A(n125), .ZN(n42) );
  AOI22_X1 U14 ( .A1(\mem[0][2] ), .A2(n2), .B1(data_in[2]), .B2(n1), .ZN(n125) );
  INV_X1 U15 ( .A(n123), .ZN(n40) );
  AOI22_X1 U16 ( .A1(\mem[0][4] ), .A2(n3), .B1(data_in[4]), .B2(n1), .ZN(n123) );
  INV_X1 U17 ( .A(n122), .ZN(n39) );
  AOI22_X1 U18 ( .A1(\mem[0][5] ), .A2(n3), .B1(data_in[5]), .B2(n1), .ZN(n122) );
  INV_X1 U19 ( .A(n121), .ZN(n38) );
  AOI22_X1 U20 ( .A1(\mem[0][6] ), .A2(n3), .B1(data_in[6]), .B2(n4), .ZN(n121) );
  INV_X1 U21 ( .A(n120), .ZN(n37) );
  AOI22_X1 U22 ( .A1(\mem[0][7] ), .A2(n3), .B1(data_in[7]), .B2(n4), .ZN(n120) );
  INV_X1 U23 ( .A(n119), .ZN(n36) );
  AOI22_X1 U24 ( .A1(\mem[0][8] ), .A2(n3), .B1(data_in[8]), .B2(n4), .ZN(n119) );
  INV_X1 U25 ( .A(n118), .ZN(n35) );
  AOI22_X1 U26 ( .A1(\mem[0][9] ), .A2(n3), .B1(data_in[9]), .B2(n1), .ZN(n118) );
  INV_X1 U27 ( .A(n117), .ZN(n34) );
  AOI22_X1 U28 ( .A1(\mem[0][10] ), .A2(n3), .B1(data_in[10]), .B2(n1), .ZN(
        n117) );
  INV_X1 U29 ( .A(n115), .ZN(n32) );
  AOI22_X1 U30 ( .A1(\mem[0][12] ), .A2(n3), .B1(data_in[12]), .B2(n1), .ZN(
        n115) );
  INV_X1 U31 ( .A(n114), .ZN(n31) );
  AOI22_X1 U32 ( .A1(\mem[0][13] ), .A2(n3), .B1(data_in[13]), .B2(n4), .ZN(
        n114) );
  INV_X1 U33 ( .A(n113), .ZN(n30) );
  AOI22_X1 U34 ( .A1(\mem[0][14] ), .A2(n3), .B1(data_in[14]), .B2(n4), .ZN(
        n113) );
  INV_X1 U35 ( .A(n112), .ZN(n29) );
  AOI22_X1 U36 ( .A1(\mem[0][15] ), .A2(n3), .B1(data_in[15]), .B2(n4), .ZN(
        n112) );
  INV_X1 U37 ( .A(n111), .ZN(n28) );
  AOI22_X1 U38 ( .A1(\mem[0][16] ), .A2(n2), .B1(data_in[16]), .B2(n4), .ZN(
        n111) );
  INV_X1 U39 ( .A(n110), .ZN(n27) );
  AOI22_X1 U40 ( .A1(\mem[0][17] ), .A2(n2), .B1(data_in[17]), .B2(n1), .ZN(
        n110) );
  INV_X1 U41 ( .A(n109), .ZN(n26) );
  AOI22_X1 U42 ( .A1(\mem[0][18] ), .A2(n2), .B1(data_in[18]), .B2(n1), .ZN(
        n109) );
  INV_X1 U43 ( .A(n108), .ZN(n25) );
  AOI22_X1 U44 ( .A1(\mem[0][19] ), .A2(n2), .B1(data_in[19]), .B2(n4), .ZN(
        n108) );
  INV_X1 U45 ( .A(n107), .ZN(n24) );
  AOI22_X1 U46 ( .A1(\mem[0][20] ), .A2(n2), .B1(data_in[20]), .B2(n1), .ZN(
        n107) );
  INV_X1 U47 ( .A(n106), .ZN(n23) );
  AOI22_X1 U48 ( .A1(\mem[0][21] ), .A2(n2), .B1(data_in[21]), .B2(n1), .ZN(
        n106) );
  INV_X1 U49 ( .A(n105), .ZN(n22) );
  AOI22_X1 U50 ( .A1(\mem[0][22] ), .A2(n2), .B1(data_in[22]), .B2(n1), .ZN(
        n105) );
  INV_X1 U51 ( .A(n104), .ZN(n21) );
  AOI22_X1 U52 ( .A1(\mem[0][23] ), .A2(n2), .B1(data_in[23]), .B2(n1), .ZN(
        n104) );
  INV_X1 U53 ( .A(n103), .ZN(n20) );
  AOI22_X1 U54 ( .A1(\mem[0][24] ), .A2(n2), .B1(data_in[24]), .B2(n4), .ZN(
        n103) );
  INV_X1 U55 ( .A(n102), .ZN(n19) );
  AOI22_X1 U56 ( .A1(\mem[0][25] ), .A2(n2), .B1(data_in[25]), .B2(n4), .ZN(
        n102) );
  INV_X1 U57 ( .A(n101), .ZN(n18) );
  AOI22_X1 U58 ( .A1(\mem[0][26] ), .A2(n2), .B1(data_in[26]), .B2(n4), .ZN(
        n101) );
  INV_X1 U59 ( .A(n100), .ZN(n17) );
  AOI22_X1 U60 ( .A1(\mem[0][27] ), .A2(n2), .B1(data_in[27]), .B2(n4), .ZN(
        n100) );
  INV_X1 U61 ( .A(n99), .ZN(n16) );
  AOI22_X1 U62 ( .A1(\mem[0][28] ), .A2(n3), .B1(data_in[28]), .B2(n1), .ZN(
        n99) );
  INV_X1 U63 ( .A(n98), .ZN(n15) );
  AOI22_X1 U64 ( .A1(\mem[0][29] ), .A2(n2), .B1(data_in[29]), .B2(n1), .ZN(
        n98) );
  INV_X1 U65 ( .A(n97), .ZN(n14) );
  AOI22_X1 U66 ( .A1(\mem[0][30] ), .A2(n3), .B1(data_in[30]), .B2(n1), .ZN(
        n97) );
  INV_X1 U67 ( .A(n96), .ZN(n13) );
  AOI22_X1 U68 ( .A1(\mem[0][31] ), .A2(n2), .B1(data_in[31]), .B2(n1), .ZN(
        n96) );
  INV_X1 U69 ( .A(n116), .ZN(n33) );
  AOI22_X1 U70 ( .A1(\mem[0][11] ), .A2(n3), .B1(data_in[11]), .B2(n1), .ZN(
        n116) );
  INV_X1 U71 ( .A(n95), .ZN(n12) );
  AOI22_X1 U72 ( .A1(\mem[0][32] ), .A2(n3), .B1(data_in[32]), .B2(n1), .ZN(
        n95) );
  INV_X1 U73 ( .A(n94), .ZN(n11) );
  AOI22_X1 U74 ( .A1(\mem[0][33] ), .A2(n2), .B1(data_in[33]), .B2(n1), .ZN(
        n94) );
  INV_X1 U75 ( .A(n93), .ZN(n10) );
  AOI22_X1 U76 ( .A1(\mem[0][34] ), .A2(n3), .B1(data_in[34]), .B2(n1), .ZN(
        n93) );
  INV_X1 U77 ( .A(n92), .ZN(n9) );
  AOI22_X1 U78 ( .A1(\mem[0][35] ), .A2(n2), .B1(data_in[35]), .B2(n1), .ZN(
        n92) );
  INV_X1 U79 ( .A(n91), .ZN(n8) );
  AOI22_X1 U80 ( .A1(\mem[0][36] ), .A2(n3), .B1(data_in[36]), .B2(n4), .ZN(
        n91) );
  INV_X1 U81 ( .A(n90), .ZN(n7) );
  AOI22_X1 U82 ( .A1(\mem[0][37] ), .A2(n2), .B1(data_in[37]), .B2(n1), .ZN(
        n90) );
  INV_X1 U83 ( .A(n89), .ZN(n6) );
  AOI22_X1 U84 ( .A1(\mem[0][38] ), .A2(n3), .B1(data_in[38]), .B2(n1), .ZN(
        n89) );
  INV_X1 U85 ( .A(n88), .ZN(n5) );
  AOI22_X1 U86 ( .A1(\mem[0][39] ), .A2(n2), .B1(data_in[39]), .B2(n4), .ZN(
        n88) );
  INV_X1 U87 ( .A(n124), .ZN(n41) );
  AOI22_X1 U88 ( .A1(\mem[0][3] ), .A2(n3), .B1(data_in[3]), .B2(n4), .ZN(n124) );
endmodule


module datapath ( clk, wr_en_x, clear_acc, wr_en_y, addr_x, addr_y, .addr_a({
        \addr_a[7][3] , \addr_a[7][2] , \addr_a[7][1] , \addr_a[7][0] , 
        \addr_a[6][3] , \addr_a[6][2] , \addr_a[6][1] , \addr_a[6][0] , 
        \addr_a[5][3] , \addr_a[5][2] , \addr_a[5][1] , \addr_a[5][0] , 
        \addr_a[4][3] , \addr_a[4][2] , \addr_a[4][1] , \addr_a[4][0] , 
        \addr_a[3][3] , \addr_a[3][2] , \addr_a[3][1] , \addr_a[3][0] , 
        \addr_a[2][3] , \addr_a[2][2] , \addr_a[2][1] , \addr_a[2][0] , 
        \addr_a[1][3] , \addr_a[1][2] , \addr_a[1][1] , \addr_a[1][0] , 
        \addr_a[0][3] , \addr_a[0][2] , \addr_a[0][1] , \addr_a[0][0] }), 
        data_in, wr_en_a, data_out );
  input [3:0] addr_x;
  input [3:0] addr_y;
  input [19:0] data_in;
  input [7:0] wr_en_a;
  output [39:0] data_out;
  input clk, wr_en_x, clear_acc, wr_en_y, \addr_a[7][3] , \addr_a[7][2] ,
         \addr_a[7][1] , \addr_a[7][0] , \addr_a[6][3] , \addr_a[6][2] ,
         \addr_a[6][1] , \addr_a[6][0] , \addr_a[5][3] , \addr_a[5][2] ,
         \addr_a[5][1] , \addr_a[5][0] , \addr_a[4][3] , \addr_a[4][2] ,
         \addr_a[4][1] , \addr_a[4][0] , \addr_a[3][3] , \addr_a[3][2] ,
         \addr_a[3][1] , \addr_a[3][0] , \addr_a[2][3] , \addr_a[2][2] ,
         \addr_a[2][1] , \addr_a[2][0] , \addr_a[1][3] , \addr_a[1][2] ,
         \addr_a[1][1] , \addr_a[1][0] , \addr_a[0][3] , \addr_a[0][2] ,
         \addr_a[0][1] , \addr_a[0][0] ;
  wire   \matrix_out[7][19] , \matrix_out[7][18] , \matrix_out[7][17] ,
         \matrix_out[7][16] , \matrix_out[7][15] , \matrix_out[7][14] ,
         \matrix_out[7][13] , \matrix_out[7][12] , \matrix_out[7][11] ,
         \matrix_out[7][10] , \matrix_out[7][9] , \matrix_out[7][8] ,
         \matrix_out[7][7] , \matrix_out[7][6] , \matrix_out[7][5] ,
         \matrix_out[7][4] , \matrix_out[7][3] , \matrix_out[7][2] ,
         \matrix_out[7][1] , \matrix_out[7][0] , \matrix_out[6][19] ,
         \matrix_out[6][18] , \matrix_out[6][17] , \matrix_out[6][16] ,
         \matrix_out[6][15] , \matrix_out[6][14] , \matrix_out[6][13] ,
         \matrix_out[6][12] , \matrix_out[6][11] , \matrix_out[6][10] ,
         \matrix_out[6][9] , \matrix_out[6][8] , \matrix_out[6][7] ,
         \matrix_out[6][6] , \matrix_out[6][5] , \matrix_out[6][4] ,
         \matrix_out[6][3] , \matrix_out[6][2] , \matrix_out[6][1] ,
         \matrix_out[6][0] , \matrix_out[5][19] , \matrix_out[5][18] ,
         \matrix_out[5][17] , \matrix_out[5][16] , \matrix_out[5][15] ,
         \matrix_out[5][14] , \matrix_out[5][13] , \matrix_out[5][12] ,
         \matrix_out[5][11] , \matrix_out[5][10] , \matrix_out[5][9] ,
         \matrix_out[5][8] , \matrix_out[5][7] , \matrix_out[5][6] ,
         \matrix_out[5][5] , \matrix_out[5][4] , \matrix_out[5][3] ,
         \matrix_out[5][2] , \matrix_out[5][1] , \matrix_out[5][0] ,
         \matrix_out[4][19] , \matrix_out[4][18] , \matrix_out[4][17] ,
         \matrix_out[4][16] , \matrix_out[4][15] , \matrix_out[4][14] ,
         \matrix_out[4][13] , \matrix_out[4][12] , \matrix_out[4][11] ,
         \matrix_out[4][10] , \matrix_out[4][9] , \matrix_out[4][8] ,
         \matrix_out[4][7] , \matrix_out[4][6] , \matrix_out[4][5] ,
         \matrix_out[4][4] , \matrix_out[4][3] , \matrix_out[4][2] ,
         \matrix_out[4][1] , \matrix_out[4][0] , \matrix_out[3][19] ,
         \matrix_out[3][18] , \matrix_out[3][17] , \matrix_out[3][16] ,
         \matrix_out[3][15] , \matrix_out[3][14] , \matrix_out[3][13] ,
         \matrix_out[3][12] , \matrix_out[3][11] , \matrix_out[3][10] ,
         \matrix_out[3][9] , \matrix_out[3][8] , \matrix_out[3][7] ,
         \matrix_out[3][6] , \matrix_out[3][5] , \matrix_out[3][4] ,
         \matrix_out[3][3] , \matrix_out[3][2] , \matrix_out[3][1] ,
         \matrix_out[3][0] , \matrix_out[2][19] , \matrix_out[2][18] ,
         \matrix_out[2][17] , \matrix_out[2][16] , \matrix_out[2][15] ,
         \matrix_out[2][14] , \matrix_out[2][13] , \matrix_out[2][12] ,
         \matrix_out[2][11] , \matrix_out[2][10] , \matrix_out[2][9] ,
         \matrix_out[2][8] , \matrix_out[2][7] , \matrix_out[2][6] ,
         \matrix_out[2][5] , \matrix_out[2][4] , \matrix_out[2][3] ,
         \matrix_out[2][2] , \matrix_out[2][1] , \matrix_out[2][0] ,
         \matrix_out[1][19] , \matrix_out[1][18] , \matrix_out[1][17] ,
         \matrix_out[1][16] , \matrix_out[1][15] , \matrix_out[1][14] ,
         \matrix_out[1][13] , \matrix_out[1][12] , \matrix_out[1][11] ,
         \matrix_out[1][10] , \matrix_out[1][9] , \matrix_out[1][8] ,
         \matrix_out[1][7] , \matrix_out[1][6] , \matrix_out[1][5] ,
         \matrix_out[1][4] , \matrix_out[1][3] , \matrix_out[1][2] ,
         \matrix_out[1][1] , \matrix_out[1][0] , \matrix_out[0][19] ,
         \matrix_out[0][18] , \matrix_out[0][17] , \matrix_out[0][16] ,
         \matrix_out[0][15] , \matrix_out[0][14] , \matrix_out[0][13] ,
         \matrix_out[0][12] , \matrix_out[0][11] , \matrix_out[0][10] ,
         \matrix_out[0][9] , \matrix_out[0][8] , \matrix_out[0][7] ,
         \matrix_out[0][6] , \matrix_out[0][5] , \matrix_out[0][4] ,
         \matrix_out[0][3] , \matrix_out[0][2] , \matrix_out[0][1] ,
         \matrix_out[0][0] , \mac_out[7][39] , \mac_out[7][38] ,
         \mac_out[7][37] , \mac_out[7][36] , \mac_out[7][35] ,
         \mac_out[7][34] , \mac_out[7][33] , \mac_out[7][32] ,
         \mac_out[7][31] , \mac_out[7][30] , \mac_out[7][29] ,
         \mac_out[7][28] , \mac_out[7][27] , \mac_out[7][26] ,
         \mac_out[7][25] , \mac_out[7][24] , \mac_out[7][23] ,
         \mac_out[7][22] , \mac_out[7][21] , \mac_out[7][20] ,
         \mac_out[7][19] , \mac_out[7][18] , \mac_out[7][17] ,
         \mac_out[7][16] , \mac_out[7][15] , \mac_out[7][14] ,
         \mac_out[7][13] , \mac_out[7][12] , \mac_out[7][11] ,
         \mac_out[7][10] , \mac_out[7][9] , \mac_out[7][8] , \mac_out[7][7] ,
         \mac_out[7][6] , \mac_out[7][5] , \mac_out[7][4] , \mac_out[7][3] ,
         \mac_out[7][2] , \mac_out[7][1] , \mac_out[7][0] , \mac_out[6][39] ,
         \mac_out[6][38] , \mac_out[6][37] , \mac_out[6][36] ,
         \mac_out[6][35] , \mac_out[6][34] , \mac_out[6][33] ,
         \mac_out[6][32] , \mac_out[6][31] , \mac_out[6][30] ,
         \mac_out[6][29] , \mac_out[6][28] , \mac_out[6][27] ,
         \mac_out[6][26] , \mac_out[6][25] , \mac_out[6][24] ,
         \mac_out[6][23] , \mac_out[6][22] , \mac_out[6][21] ,
         \mac_out[6][20] , \mac_out[6][19] , \mac_out[6][18] ,
         \mac_out[6][17] , \mac_out[6][16] , \mac_out[6][15] ,
         \mac_out[6][14] , \mac_out[6][13] , \mac_out[6][12] ,
         \mac_out[6][11] , \mac_out[6][10] , \mac_out[6][9] , \mac_out[6][8] ,
         \mac_out[6][7] , \mac_out[6][6] , \mac_out[6][5] , \mac_out[6][4] ,
         \mac_out[6][3] , \mac_out[6][2] , \mac_out[6][1] , \mac_out[6][0] ,
         \mac_out[5][39] , \mac_out[5][38] , \mac_out[5][37] ,
         \mac_out[5][36] , \mac_out[5][35] , \mac_out[5][34] ,
         \mac_out[5][33] , \mac_out[5][32] , \mac_out[5][31] ,
         \mac_out[5][30] , \mac_out[5][29] , \mac_out[5][28] ,
         \mac_out[5][27] , \mac_out[5][26] , \mac_out[5][25] ,
         \mac_out[5][24] , \mac_out[5][23] , \mac_out[5][22] ,
         \mac_out[5][21] , \mac_out[5][20] , \mac_out[5][19] ,
         \mac_out[5][18] , \mac_out[5][17] , \mac_out[5][16] ,
         \mac_out[5][15] , \mac_out[5][14] , \mac_out[5][13] ,
         \mac_out[5][12] , \mac_out[5][11] , \mac_out[5][10] , \mac_out[5][9] ,
         \mac_out[5][8] , \mac_out[5][7] , \mac_out[5][6] , \mac_out[5][5] ,
         \mac_out[5][4] , \mac_out[5][3] , \mac_out[5][2] , \mac_out[5][1] ,
         \mac_out[5][0] , \mac_out[4][39] , \mac_out[4][38] , \mac_out[4][37] ,
         \mac_out[4][36] , \mac_out[4][35] , \mac_out[4][34] ,
         \mac_out[4][33] , \mac_out[4][32] , \mac_out[4][31] ,
         \mac_out[4][30] , \mac_out[4][29] , \mac_out[4][28] ,
         \mac_out[4][27] , \mac_out[4][26] , \mac_out[4][25] ,
         \mac_out[4][24] , \mac_out[4][23] , \mac_out[4][22] ,
         \mac_out[4][21] , \mac_out[4][20] , \mac_out[4][19] ,
         \mac_out[4][18] , \mac_out[4][17] , \mac_out[4][16] ,
         \mac_out[4][15] , \mac_out[4][14] , \mac_out[4][13] ,
         \mac_out[4][12] , \mac_out[4][11] , \mac_out[4][10] , \mac_out[4][9] ,
         \mac_out[4][8] , \mac_out[4][7] , \mac_out[4][6] , \mac_out[4][5] ,
         \mac_out[4][4] , \mac_out[4][3] , \mac_out[4][2] , \mac_out[4][1] ,
         \mac_out[4][0] , \mac_out[3][39] , \mac_out[3][38] , \mac_out[3][37] ,
         \mac_out[3][36] , \mac_out[3][35] , \mac_out[3][34] ,
         \mac_out[3][33] , \mac_out[3][32] , \mac_out[3][31] ,
         \mac_out[3][30] , \mac_out[3][29] , \mac_out[3][28] ,
         \mac_out[3][27] , \mac_out[3][26] , \mac_out[3][25] ,
         \mac_out[3][24] , \mac_out[3][23] , \mac_out[3][22] ,
         \mac_out[3][21] , \mac_out[3][20] , \mac_out[3][19] ,
         \mac_out[3][18] , \mac_out[3][17] , \mac_out[3][16] ,
         \mac_out[3][15] , \mac_out[3][14] , \mac_out[3][13] ,
         \mac_out[3][12] , \mac_out[3][11] , \mac_out[3][10] , \mac_out[3][9] ,
         \mac_out[3][8] , \mac_out[3][7] , \mac_out[3][6] , \mac_out[3][5] ,
         \mac_out[3][4] , \mac_out[3][3] , \mac_out[3][2] , \mac_out[3][1] ,
         \mac_out[3][0] , \mac_out[2][39] , \mac_out[2][38] , \mac_out[2][37] ,
         \mac_out[2][36] , \mac_out[2][35] , \mac_out[2][34] ,
         \mac_out[2][33] , \mac_out[2][32] , \mac_out[2][31] ,
         \mac_out[2][30] , \mac_out[2][29] , \mac_out[2][28] ,
         \mac_out[2][27] , \mac_out[2][26] , \mac_out[2][25] ,
         \mac_out[2][24] , \mac_out[2][23] , \mac_out[2][22] ,
         \mac_out[2][21] , \mac_out[2][20] , \mac_out[2][19] ,
         \mac_out[2][18] , \mac_out[2][17] , \mac_out[2][16] ,
         \mac_out[2][15] , \mac_out[2][14] , \mac_out[2][13] ,
         \mac_out[2][12] , \mac_out[2][11] , \mac_out[2][10] , \mac_out[2][9] ,
         \mac_out[2][8] , \mac_out[2][7] , \mac_out[2][6] , \mac_out[2][5] ,
         \mac_out[2][4] , \mac_out[2][3] , \mac_out[2][2] , \mac_out[2][1] ,
         \mac_out[2][0] , \mac_out[1][39] , \mac_out[1][38] , \mac_out[1][37] ,
         \mac_out[1][36] , \mac_out[1][35] , \mac_out[1][34] ,
         \mac_out[1][33] , \mac_out[1][32] , \mac_out[1][31] ,
         \mac_out[1][30] , \mac_out[1][29] , \mac_out[1][28] ,
         \mac_out[1][27] , \mac_out[1][26] , \mac_out[1][25] ,
         \mac_out[1][24] , \mac_out[1][23] , \mac_out[1][22] ,
         \mac_out[1][21] , \mac_out[1][20] , \mac_out[1][19] ,
         \mac_out[1][18] , \mac_out[1][17] , \mac_out[1][16] ,
         \mac_out[1][15] , \mac_out[1][14] , \mac_out[1][13] ,
         \mac_out[1][12] , \mac_out[1][11] , \mac_out[1][10] , \mac_out[1][9] ,
         \mac_out[1][8] , \mac_out[1][7] , \mac_out[1][6] , \mac_out[1][5] ,
         \mac_out[1][4] , \mac_out[1][3] , \mac_out[1][2] , \mac_out[1][1] ,
         \mac_out[1][0] , \mac_out[0][39] , \mac_out[0][38] , \mac_out[0][37] ,
         \mac_out[0][36] , \mac_out[0][35] , \mac_out[0][34] ,
         \mac_out[0][33] , \mac_out[0][32] , \mac_out[0][31] ,
         \mac_out[0][30] , \mac_out[0][29] , \mac_out[0][28] ,
         \mac_out[0][27] , \mac_out[0][26] , \mac_out[0][25] ,
         \mac_out[0][24] , \mac_out[0][23] , \mac_out[0][22] ,
         \mac_out[0][21] , \mac_out[0][20] , \mac_out[0][19] ,
         \mac_out[0][18] , \mac_out[0][17] , \mac_out[0][16] ,
         \mac_out[0][15] , \mac_out[0][14] , \mac_out[0][13] ,
         \mac_out[0][12] , \mac_out[0][11] , \mac_out[0][10] , \mac_out[0][9] ,
         \mac_out[0][8] , \mac_out[0][7] , \mac_out[0][6] , \mac_out[0][5] ,
         \mac_out[0][4] , \mac_out[0][3] , \mac_out[0][2] , \mac_out[0][1] ,
         \mac_out[0][0] , \mux[7][39] , \mux[7][38] , \mux[7][37] ,
         \mux[7][36] , \mux[7][35] , \mux[7][34] , \mux[7][33] , \mux[7][32] ,
         \mux[7][31] , \mux[7][30] , \mux[7][29] , \mux[7][28] , \mux[7][27] ,
         \mux[7][26] , \mux[7][25] , \mux[7][24] , \mux[7][23] , \mux[7][22] ,
         \mux[7][21] , \mux[7][20] , \mux[7][19] , \mux[7][18] , \mux[7][17] ,
         \mux[7][16] , \mux[7][15] , \mux[7][14] , \mux[7][13] , \mux[7][12] ,
         \mux[7][11] , \mux[7][10] , \mux[7][9] , \mux[7][8] , \mux[7][7] ,
         \mux[7][6] , \mux[7][5] , \mux[7][4] , \mux[7][3] , \mux[7][2] ,
         \mux[7][1] , \mux[7][0] , \mux[6][39] , \mux[6][38] , \mux[6][37] ,
         \mux[6][36] , \mux[6][35] , \mux[6][34] , \mux[6][33] , \mux[6][32] ,
         \mux[6][31] , \mux[6][30] , \mux[6][29] , \mux[6][28] , \mux[6][27] ,
         \mux[6][26] , \mux[6][25] , \mux[6][24] , \mux[6][23] , \mux[6][22] ,
         \mux[6][21] , \mux[6][20] , \mux[6][19] , \mux[6][18] , \mux[6][17] ,
         \mux[6][16] , \mux[6][15] , \mux[6][14] , \mux[6][13] , \mux[6][12] ,
         \mux[6][11] , \mux[6][10] , \mux[6][9] , \mux[6][8] , \mux[6][7] ,
         \mux[6][6] , \mux[6][5] , \mux[6][4] , \mux[6][3] , \mux[6][2] ,
         \mux[6][1] , \mux[6][0] , \mux[5][39] , \mux[5][38] , \mux[5][37] ,
         \mux[5][36] , \mux[5][35] , \mux[5][34] , \mux[5][33] , \mux[5][32] ,
         \mux[5][31] , \mux[5][30] , \mux[5][29] , \mux[5][28] , \mux[5][27] ,
         \mux[5][26] , \mux[5][25] , \mux[5][24] , \mux[5][23] , \mux[5][22] ,
         \mux[5][21] , \mux[5][20] , \mux[5][19] , \mux[5][18] , \mux[5][17] ,
         \mux[5][16] , \mux[5][15] , \mux[5][14] , \mux[5][13] , \mux[5][12] ,
         \mux[5][11] , \mux[5][10] , \mux[5][9] , \mux[5][8] , \mux[5][7] ,
         \mux[5][6] , \mux[5][5] , \mux[5][4] , \mux[5][3] , \mux[5][2] ,
         \mux[5][1] , \mux[5][0] , \mux[4][39] , \mux[4][38] , \mux[4][37] ,
         \mux[4][36] , \mux[4][35] , \mux[4][34] , \mux[4][33] , \mux[4][32] ,
         \mux[4][31] , \mux[4][30] , \mux[4][29] , \mux[4][28] , \mux[4][27] ,
         \mux[4][26] , \mux[4][25] , \mux[4][24] , \mux[4][23] , \mux[4][22] ,
         \mux[4][21] , \mux[4][20] , \mux[4][19] , \mux[4][18] , \mux[4][17] ,
         \mux[4][16] , \mux[4][15] , \mux[4][14] , \mux[4][13] , \mux[4][12] ,
         \mux[4][11] , \mux[4][10] , \mux[4][9] , \mux[4][8] , \mux[4][7] ,
         \mux[4][6] , \mux[4][5] , \mux[4][4] , \mux[4][3] , \mux[4][2] ,
         \mux[4][1] , \mux[4][0] , \mux[3][39] , \mux[3][38] , \mux[3][37] ,
         \mux[3][36] , \mux[3][35] , \mux[3][34] , \mux[3][33] , \mux[3][32] ,
         \mux[3][31] , \mux[3][30] , \mux[3][29] , \mux[3][28] , \mux[3][27] ,
         \mux[3][26] , \mux[3][25] , \mux[3][24] , \mux[3][23] , \mux[3][22] ,
         \mux[3][21] , \mux[3][20] , \mux[3][19] , \mux[3][18] , \mux[3][17] ,
         \mux[3][16] , \mux[3][15] , \mux[3][14] , \mux[3][13] , \mux[3][12] ,
         \mux[3][11] , \mux[3][10] , \mux[3][9] , \mux[3][8] , \mux[3][7] ,
         \mux[3][6] , \mux[3][5] , \mux[3][4] , \mux[3][3] , \mux[3][2] ,
         \mux[3][1] , \mux[3][0] , \mux[2][39] , \mux[2][38] , \mux[2][37] ,
         \mux[2][36] , \mux[2][35] , \mux[2][34] , \mux[2][33] , \mux[2][32] ,
         \mux[2][31] , \mux[2][30] , \mux[2][29] , \mux[2][28] , \mux[2][27] ,
         \mux[2][26] , \mux[2][25] , \mux[2][24] , \mux[2][23] , \mux[2][22] ,
         \mux[2][21] , \mux[2][20] , \mux[2][19] , \mux[2][18] , \mux[2][17] ,
         \mux[2][16] , \mux[2][15] , \mux[2][14] , \mux[2][13] , \mux[2][12] ,
         \mux[2][11] , \mux[2][10] , \mux[2][9] , \mux[2][8] , \mux[2][7] ,
         \mux[2][6] , \mux[2][5] , \mux[2][4] , \mux[2][3] , \mux[2][2] ,
         \mux[2][1] , \mux[2][0] , \mux[1][39] , \mux[1][38] , \mux[1][37] ,
         \mux[1][36] , \mux[1][35] , \mux[1][34] , \mux[1][33] , \mux[1][32] ,
         \mux[1][31] , \mux[1][30] , \mux[1][29] , \mux[1][28] , \mux[1][27] ,
         \mux[1][26] , \mux[1][25] , \mux[1][24] , \mux[1][23] , \mux[1][22] ,
         \mux[1][21] , \mux[1][20] , \mux[1][19] , \mux[1][18] , \mux[1][17] ,
         \mux[1][16] , \mux[1][15] , \mux[1][14] , \mux[1][13] , \mux[1][12] ,
         \mux[1][11] , \mux[1][10] , \mux[1][9] , \mux[1][8] , \mux[1][7] ,
         \mux[1][6] , \mux[1][5] , \mux[1][4] , \mux[1][3] , \mux[1][2] ,
         \mux[1][1] , \mux[1][0] , \mux[0][39] , \mux[0][38] , \mux[0][37] ,
         \mux[0][36] , \mux[0][35] , \mux[0][34] , \mux[0][33] , \mux[0][32] ,
         \mux[0][31] , \mux[0][30] , \mux[0][29] , \mux[0][28] , \mux[0][27] ,
         \mux[0][26] , \mux[0][25] , \mux[0][24] , \mux[0][23] , \mux[0][22] ,
         \mux[0][21] , \mux[0][20] , \mux[0][19] , \mux[0][18] , \mux[0][17] ,
         \mux[0][16] , \mux[0][15] , \mux[0][14] , \mux[0][13] , \mux[0][12] ,
         \mux[0][11] , \mux[0][10] , \mux[0][9] , \mux[0][8] , \mux[0][7] ,
         \mux[0][6] , \mux[0][5] , \mux[0][4] , \mux[0][3] , \mux[0][2] ,
         \mux[0][1] , \mux[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305;
  wire   [19:0] vector_out;

  memory_WIDTH20_SIZE8_LOGSIZE4_8 \matrix[0]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[0][19] , \matrix_out[0][18] , 
        \matrix_out[0][17] , \matrix_out[0][16] , \matrix_out[0][15] , 
        \matrix_out[0][14] , \matrix_out[0][13] , \matrix_out[0][12] , 
        \matrix_out[0][11] , \matrix_out[0][10] , \matrix_out[0][9] , 
        \matrix_out[0][8] , \matrix_out[0][7] , \matrix_out[0][6] , 
        \matrix_out[0][5] , \matrix_out[0][4] , \matrix_out[0][3] , 
        \matrix_out[0][2] , \matrix_out[0][1] , \matrix_out[0][0] }), .addr({
        \addr_a[0][3] , \addr_a[0][2] , \addr_a[0][1] , \addr_a[0][0] }), 
        .wr_en(wr_en_a[0]) );
  memory_WIDTH20_SIZE8_LOGSIZE4_7 \matrix[1]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[1][19] , \matrix_out[1][18] , 
        \matrix_out[1][17] , \matrix_out[1][16] , \matrix_out[1][15] , 
        \matrix_out[1][14] , \matrix_out[1][13] , \matrix_out[1][12] , 
        \matrix_out[1][11] , \matrix_out[1][10] , \matrix_out[1][9] , 
        \matrix_out[1][8] , \matrix_out[1][7] , \matrix_out[1][6] , 
        \matrix_out[1][5] , \matrix_out[1][4] , \matrix_out[1][3] , 
        \matrix_out[1][2] , \matrix_out[1][1] , \matrix_out[1][0] }), .addr({
        \addr_a[1][3] , \addr_a[1][2] , \addr_a[1][1] , \addr_a[1][0] }), 
        .wr_en(wr_en_a[1]) );
  memory_WIDTH20_SIZE8_LOGSIZE4_6 \matrix[2]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[2][19] , \matrix_out[2][18] , 
        \matrix_out[2][17] , \matrix_out[2][16] , \matrix_out[2][15] , 
        \matrix_out[2][14] , \matrix_out[2][13] , \matrix_out[2][12] , 
        \matrix_out[2][11] , \matrix_out[2][10] , \matrix_out[2][9] , 
        \matrix_out[2][8] , \matrix_out[2][7] , \matrix_out[2][6] , 
        \matrix_out[2][5] , \matrix_out[2][4] , \matrix_out[2][3] , 
        \matrix_out[2][2] , \matrix_out[2][1] , \matrix_out[2][0] }), .addr({
        \addr_a[2][3] , \addr_a[2][2] , \addr_a[2][1] , \addr_a[2][0] }), 
        .wr_en(wr_en_a[2]) );
  memory_WIDTH20_SIZE8_LOGSIZE4_5 \matrix[3]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[3][19] , \matrix_out[3][18] , 
        \matrix_out[3][17] , \matrix_out[3][16] , \matrix_out[3][15] , 
        \matrix_out[3][14] , \matrix_out[3][13] , \matrix_out[3][12] , 
        \matrix_out[3][11] , \matrix_out[3][10] , \matrix_out[3][9] , 
        \matrix_out[3][8] , \matrix_out[3][7] , \matrix_out[3][6] , 
        \matrix_out[3][5] , \matrix_out[3][4] , \matrix_out[3][3] , 
        \matrix_out[3][2] , \matrix_out[3][1] , \matrix_out[3][0] }), .addr({
        \addr_a[3][3] , \addr_a[3][2] , \addr_a[3][1] , \addr_a[3][0] }), 
        .wr_en(wr_en_a[3]) );
  memory_WIDTH20_SIZE8_LOGSIZE4_4 \matrix[4]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[4][19] , \matrix_out[4][18] , 
        \matrix_out[4][17] , \matrix_out[4][16] , \matrix_out[4][15] , 
        \matrix_out[4][14] , \matrix_out[4][13] , \matrix_out[4][12] , 
        \matrix_out[4][11] , \matrix_out[4][10] , \matrix_out[4][9] , 
        \matrix_out[4][8] , \matrix_out[4][7] , \matrix_out[4][6] , 
        \matrix_out[4][5] , \matrix_out[4][4] , \matrix_out[4][3] , 
        \matrix_out[4][2] , \matrix_out[4][1] , \matrix_out[4][0] }), .addr({
        \addr_a[4][3] , \addr_a[4][2] , \addr_a[4][1] , \addr_a[4][0] }), 
        .wr_en(wr_en_a[4]) );
  memory_WIDTH20_SIZE8_LOGSIZE4_3 \matrix[5]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[5][19] , \matrix_out[5][18] , 
        \matrix_out[5][17] , \matrix_out[5][16] , \matrix_out[5][15] , 
        \matrix_out[5][14] , \matrix_out[5][13] , \matrix_out[5][12] , 
        \matrix_out[5][11] , \matrix_out[5][10] , \matrix_out[5][9] , 
        \matrix_out[5][8] , \matrix_out[5][7] , \matrix_out[5][6] , 
        \matrix_out[5][5] , \matrix_out[5][4] , \matrix_out[5][3] , 
        \matrix_out[5][2] , \matrix_out[5][1] , \matrix_out[5][0] }), .addr({
        \addr_a[5][3] , \addr_a[5][2] , \addr_a[5][1] , \addr_a[5][0] }), 
        .wr_en(wr_en_a[5]) );
  memory_WIDTH20_SIZE8_LOGSIZE4_2 \matrix[6]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[6][19] , \matrix_out[6][18] , 
        \matrix_out[6][17] , \matrix_out[6][16] , \matrix_out[6][15] , 
        \matrix_out[6][14] , \matrix_out[6][13] , \matrix_out[6][12] , 
        \matrix_out[6][11] , \matrix_out[6][10] , \matrix_out[6][9] , 
        \matrix_out[6][8] , \matrix_out[6][7] , \matrix_out[6][6] , 
        \matrix_out[6][5] , \matrix_out[6][4] , \matrix_out[6][3] , 
        \matrix_out[6][2] , \matrix_out[6][1] , \matrix_out[6][0] }), .addr({
        \addr_a[6][3] , \addr_a[6][2] , \addr_a[6][1] , \addr_a[6][0] }), 
        .wr_en(wr_en_a[6]) );
  memory_WIDTH20_SIZE8_LOGSIZE4_1 \matrix[7]  ( .clk(clk), .data_in(data_in), 
        .data_out({\matrix_out[7][19] , \matrix_out[7][18] , 
        \matrix_out[7][17] , \matrix_out[7][16] , \matrix_out[7][15] , 
        \matrix_out[7][14] , \matrix_out[7][13] , \matrix_out[7][12] , 
        \matrix_out[7][11] , \matrix_out[7][10] , \matrix_out[7][9] , 
        \matrix_out[7][8] , \matrix_out[7][7] , \matrix_out[7][6] , 
        \matrix_out[7][5] , \matrix_out[7][4] , \matrix_out[7][3] , 
        \matrix_out[7][2] , \matrix_out[7][1] , \matrix_out[7][0] }), .addr({
        \addr_a[7][3] , \addr_a[7][2] , \addr_a[7][1] , \addr_a[7][0] }), 
        .wr_en(wr_en_a[7]) );
  memory_WIDTH20_SIZE8_LOGSIZE4_0 vector ( .clk(clk), .data_in(data_in), 
        .data_out(vector_out), .addr(addr_x), .wr_en(wr_en_x) );
  mac_7 \mac_mod[0]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[0][19] , \matrix_out[0][18] , \matrix_out[0][17] , 
        \matrix_out[0][16] , \matrix_out[0][15] , \matrix_out[0][14] , 
        \matrix_out[0][13] , \matrix_out[0][12] , \matrix_out[0][11] , 
        \matrix_out[0][10] , \matrix_out[0][9] , \matrix_out[0][8] , 
        \matrix_out[0][7] , \matrix_out[0][6] , \matrix_out[0][5] , 
        \matrix_out[0][4] , \matrix_out[0][3] , \matrix_out[0][2] , 
        \matrix_out[0][1] , \matrix_out[0][0] }), .b({n305, n302, 
        vector_out[17], n299, n295, n294, n291, n290, n287, n284, n281, n278, 
        n275, n272, n3, n270, n7, n267, n263, n9}), .mac_out({\mac_out[0][39] , 
        \mac_out[0][38] , \mac_out[0][37] , \mac_out[0][36] , \mac_out[0][35] , 
        \mac_out[0][34] , \mac_out[0][33] , \mac_out[0][32] , \mac_out[0][31] , 
        \mac_out[0][30] , \mac_out[0][29] , \mac_out[0][28] , \mac_out[0][27] , 
        \mac_out[0][26] , \mac_out[0][25] , \mac_out[0][24] , \mac_out[0][23] , 
        \mac_out[0][22] , \mac_out[0][21] , \mac_out[0][20] , \mac_out[0][19] , 
        \mac_out[0][18] , \mac_out[0][17] , \mac_out[0][16] , \mac_out[0][15] , 
        \mac_out[0][14] , \mac_out[0][13] , \mac_out[0][12] , \mac_out[0][11] , 
        \mac_out[0][10] , \mac_out[0][9] , \mac_out[0][8] , \mac_out[0][7] , 
        \mac_out[0][6] , \mac_out[0][5] , \mac_out[0][4] , \mac_out[0][3] , 
        \mac_out[0][2] , \mac_out[0][1] , \mac_out[0][0] }) );
  mac_6 \mac_mod[1]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[1][19] , \matrix_out[1][18] , \matrix_out[1][17] , 
        \matrix_out[1][16] , \matrix_out[1][15] , \matrix_out[1][14] , 
        \matrix_out[1][13] , \matrix_out[1][12] , \matrix_out[1][11] , 
        \matrix_out[1][10] , \matrix_out[1][9] , \matrix_out[1][8] , 
        \matrix_out[1][7] , \matrix_out[1][6] , \matrix_out[1][5] , 
        \matrix_out[1][4] , \matrix_out[1][3] , \matrix_out[1][2] , 
        \matrix_out[1][1] , \matrix_out[1][0] }), .b({n303, n300, 
        vector_out[17], n297, n295, n293, n292, n288, n285, n282, n279, n276, 
        n273, n271, n2, n5, n268, n267, n4, n9}), .mac_out({\mac_out[1][39] , 
        \mac_out[1][38] , \mac_out[1][37] , \mac_out[1][36] , \mac_out[1][35] , 
        \mac_out[1][34] , \mac_out[1][33] , \mac_out[1][32] , \mac_out[1][31] , 
        \mac_out[1][30] , \mac_out[1][29] , \mac_out[1][28] , \mac_out[1][27] , 
        \mac_out[1][26] , \mac_out[1][25] , \mac_out[1][24] , \mac_out[1][23] , 
        \mac_out[1][22] , \mac_out[1][21] , \mac_out[1][20] , \mac_out[1][19] , 
        \mac_out[1][18] , \mac_out[1][17] , \mac_out[1][16] , \mac_out[1][15] , 
        \mac_out[1][14] , \mac_out[1][13] , \mac_out[1][12] , \mac_out[1][11] , 
        \mac_out[1][10] , \mac_out[1][9] , \mac_out[1][8] , \mac_out[1][7] , 
        \mac_out[1][6] , \mac_out[1][5] , \mac_out[1][4] , \mac_out[1][3] , 
        \mac_out[1][2] , \mac_out[1][1] , \mac_out[1][0] }) );
  mac_5 \mac_mod[2]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[2][19] , \matrix_out[2][18] , \matrix_out[2][17] , 
        \matrix_out[2][16] , \matrix_out[2][15] , \matrix_out[2][14] , 
        \matrix_out[2][13] , \matrix_out[2][12] , \matrix_out[2][11] , 
        \matrix_out[2][10] , \matrix_out[2][9] , \matrix_out[2][8] , 
        \matrix_out[2][7] , \matrix_out[2][6] , \matrix_out[2][5] , 
        \matrix_out[2][4] , \matrix_out[2][3] , \matrix_out[2][2] , 
        \matrix_out[2][1] , \matrix_out[2][0] }), .b({n303, n300, 
        vector_out[17], n297, n295, n293, n291, n288, n285, n282, n279, n276, 
        n273, n271, n3, n270, n7, n266, n4, n9}), .mac_out({\mac_out[2][39] , 
        \mac_out[2][38] , \mac_out[2][37] , \mac_out[2][36] , \mac_out[2][35] , 
        \mac_out[2][34] , \mac_out[2][33] , \mac_out[2][32] , \mac_out[2][31] , 
        \mac_out[2][30] , \mac_out[2][29] , \mac_out[2][28] , \mac_out[2][27] , 
        \mac_out[2][26] , \mac_out[2][25] , \mac_out[2][24] , \mac_out[2][23] , 
        \mac_out[2][22] , \mac_out[2][21] , \mac_out[2][20] , \mac_out[2][19] , 
        \mac_out[2][18] , \mac_out[2][17] , \mac_out[2][16] , \mac_out[2][15] , 
        \mac_out[2][14] , \mac_out[2][13] , \mac_out[2][12] , \mac_out[2][11] , 
        \mac_out[2][10] , \mac_out[2][9] , \mac_out[2][8] , \mac_out[2][7] , 
        \mac_out[2][6] , \mac_out[2][5] , \mac_out[2][4] , \mac_out[2][3] , 
        \mac_out[2][2] , \mac_out[2][1] , \mac_out[2][0] }) );
  mac_4 \mac_mod[3]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[3][19] , \matrix_out[3][18] , \matrix_out[3][17] , 
        \matrix_out[3][16] , \matrix_out[3][15] , \matrix_out[3][14] , 
        \matrix_out[3][13] , \matrix_out[3][12] , \matrix_out[3][11] , 
        \matrix_out[3][10] , \matrix_out[3][9] , \matrix_out[3][8] , 
        \matrix_out[3][7] , \matrix_out[3][6] , \matrix_out[3][5] , 
        \matrix_out[3][4] , \matrix_out[3][3] , \matrix_out[3][2] , 
        \matrix_out[3][1] , \matrix_out[3][0] }), .b({n303, n300, 
        vector_out[17], n297, n295, n293, n292, n288, n285, n282, n279, n277, 
        n273, n271, n2, n5, n268, n266, n265, n8}), .mac_out({\mac_out[3][39] , 
        \mac_out[3][38] , \mac_out[3][37] , \mac_out[3][36] , \mac_out[3][35] , 
        \mac_out[3][34] , \mac_out[3][33] , \mac_out[3][32] , \mac_out[3][31] , 
        \mac_out[3][30] , \mac_out[3][29] , \mac_out[3][28] , \mac_out[3][27] , 
        \mac_out[3][26] , \mac_out[3][25] , \mac_out[3][24] , \mac_out[3][23] , 
        \mac_out[3][22] , \mac_out[3][21] , \mac_out[3][20] , \mac_out[3][19] , 
        \mac_out[3][18] , \mac_out[3][17] , \mac_out[3][16] , \mac_out[3][15] , 
        \mac_out[3][14] , \mac_out[3][13] , \mac_out[3][12] , \mac_out[3][11] , 
        \mac_out[3][10] , \mac_out[3][9] , \mac_out[3][8] , \mac_out[3][7] , 
        \mac_out[3][6] , \mac_out[3][5] , \mac_out[3][4] , \mac_out[3][3] , 
        \mac_out[3][2] , \mac_out[3][1] , \mac_out[3][0] }) );
  mac_3 \mac_mod[4]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[4][19] , \matrix_out[4][18] , \matrix_out[4][17] , 
        \matrix_out[4][16] , \matrix_out[4][15] , \matrix_out[4][14] , 
        \matrix_out[4][13] , \matrix_out[4][12] , \matrix_out[4][11] , 
        \matrix_out[4][10] , \matrix_out[4][9] , \matrix_out[4][8] , 
        \matrix_out[4][7] , \matrix_out[4][6] , \matrix_out[4][5] , 
        \matrix_out[4][4] , \matrix_out[4][3] , \matrix_out[4][2] , 
        \matrix_out[4][1] , \matrix_out[4][0] }), .b({n304, n301, 
        vector_out[17], n298, n296, n294, n291, n289, n286, n283, n280, n278, 
        n274, n271, n2, vector_out[4], n7, n267, n263, n8}), .mac_out({
        \mac_out[4][39] , \mac_out[4][38] , \mac_out[4][37] , \mac_out[4][36] , 
        \mac_out[4][35] , \mac_out[4][34] , \mac_out[4][33] , \mac_out[4][32] , 
        \mac_out[4][31] , \mac_out[4][30] , \mac_out[4][29] , \mac_out[4][28] , 
        \mac_out[4][27] , \mac_out[4][26] , \mac_out[4][25] , \mac_out[4][24] , 
        \mac_out[4][23] , \mac_out[4][22] , \mac_out[4][21] , \mac_out[4][20] , 
        \mac_out[4][19] , \mac_out[4][18] , \mac_out[4][17] , \mac_out[4][16] , 
        \mac_out[4][15] , \mac_out[4][14] , \mac_out[4][13] , \mac_out[4][12] , 
        \mac_out[4][11] , \mac_out[4][10] , \mac_out[4][9] , \mac_out[4][8] , 
        \mac_out[4][7] , \mac_out[4][6] , \mac_out[4][5] , \mac_out[4][4] , 
        \mac_out[4][3] , \mac_out[4][2] , \mac_out[4][1] , \mac_out[4][0] })
         );
  mac_2 \mac_mod[5]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[5][19] , \matrix_out[5][18] , \matrix_out[5][17] , 
        \matrix_out[5][16] , \matrix_out[5][15] , \matrix_out[5][14] , 
        \matrix_out[5][13] , \matrix_out[5][12] , \matrix_out[5][11] , 
        \matrix_out[5][10] , \matrix_out[5][9] , \matrix_out[5][8] , 
        \matrix_out[5][7] , \matrix_out[5][6] , \matrix_out[5][5] , 
        \matrix_out[5][4] , \matrix_out[5][3] , \matrix_out[5][2] , 
        \matrix_out[5][1] , \matrix_out[5][0] }), .b({n304, n301, 
        vector_out[17], n298, n296, n294, n292, n289, n286, n283, n280, n277, 
        n275, n271, n1, vector_out[4], n7, n266, n264, n9}), .mac_out({
        \mac_out[5][39] , \mac_out[5][38] , \mac_out[5][37] , \mac_out[5][36] , 
        \mac_out[5][35] , \mac_out[5][34] , \mac_out[5][33] , \mac_out[5][32] , 
        \mac_out[5][31] , \mac_out[5][30] , \mac_out[5][29] , \mac_out[5][28] , 
        \mac_out[5][27] , \mac_out[5][26] , \mac_out[5][25] , \mac_out[5][24] , 
        \mac_out[5][23] , \mac_out[5][22] , \mac_out[5][21] , \mac_out[5][20] , 
        \mac_out[5][19] , \mac_out[5][18] , \mac_out[5][17] , \mac_out[5][16] , 
        \mac_out[5][15] , \mac_out[5][14] , \mac_out[5][13] , \mac_out[5][12] , 
        \mac_out[5][11] , \mac_out[5][10] , \mac_out[5][9] , \mac_out[5][8] , 
        \mac_out[5][7] , \mac_out[5][6] , \mac_out[5][5] , \mac_out[5][4] , 
        \mac_out[5][3] , \mac_out[5][2] , \mac_out[5][1] , \mac_out[5][0] })
         );
  mac_1 \mac_mod[6]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[6][19] , \matrix_out[6][18] , \matrix_out[6][17] , 
        \matrix_out[6][16] , \matrix_out[6][15] , \matrix_out[6][14] , 
        \matrix_out[6][13] , \matrix_out[6][12] , \matrix_out[6][11] , 
        \matrix_out[6][10] , \matrix_out[6][9] , \matrix_out[6][8] , 
        \matrix_out[6][7] , \matrix_out[6][6] , \matrix_out[6][5] , 
        \matrix_out[6][4] , \matrix_out[6][3] , \matrix_out[6][2] , 
        \matrix_out[6][1] , \matrix_out[6][0] }), .b({n303, n301, 
        vector_out[17], n298, n296, n294, n291, n289, n286, n283, n280, n6, 
        n274, n272, n1, n5, n269, n267, vector_out[1], n8}), .mac_out({
        \mac_out[6][39] , \mac_out[6][38] , \mac_out[6][37] , \mac_out[6][36] , 
        \mac_out[6][35] , \mac_out[6][34] , \mac_out[6][33] , \mac_out[6][32] , 
        \mac_out[6][31] , \mac_out[6][30] , \mac_out[6][29] , \mac_out[6][28] , 
        \mac_out[6][27] , \mac_out[6][26] , \mac_out[6][25] , \mac_out[6][24] , 
        \mac_out[6][23] , \mac_out[6][22] , \mac_out[6][21] , \mac_out[6][20] , 
        \mac_out[6][19] , \mac_out[6][18] , \mac_out[6][17] , \mac_out[6][16] , 
        \mac_out[6][15] , \mac_out[6][14] , \mac_out[6][13] , \mac_out[6][12] , 
        \mac_out[6][11] , \mac_out[6][10] , \mac_out[6][9] , \mac_out[6][8] , 
        \mac_out[6][7] , \mac_out[6][6] , \mac_out[6][5] , \mac_out[6][4] , 
        \mac_out[6][3] , \mac_out[6][2] , \mac_out[6][1] , \mac_out[6][0] })
         );
  mac_0 \mac_mod[7]  ( .clk(clk), .clear_acc(clear_acc), .a({
        \matrix_out[7][19] , \matrix_out[7][18] , \matrix_out[7][17] , 
        \matrix_out[7][16] , \matrix_out[7][15] , \matrix_out[7][14] , 
        \matrix_out[7][13] , \matrix_out[7][12] , \matrix_out[7][11] , 
        \matrix_out[7][10] , \matrix_out[7][9] , \matrix_out[7][8] , 
        \matrix_out[7][7] , \matrix_out[7][6] , \matrix_out[7][5] , 
        \matrix_out[7][4] , \matrix_out[7][3] , \matrix_out[7][2] , 
        \matrix_out[7][1] , \matrix_out[7][0] }), .b({n305, n302, 
        vector_out[17], n299, n295, n294, n292, n290, n287, n284, n281, n6, 
        n275, n272, n1, n5, n269, n267, n264, n8}), .mac_out({\mac_out[7][39] , 
        \mac_out[7][38] , \mac_out[7][37] , \mac_out[7][36] , \mac_out[7][35] , 
        \mac_out[7][34] , \mac_out[7][33] , \mac_out[7][32] , \mac_out[7][31] , 
        \mac_out[7][30] , \mac_out[7][29] , \mac_out[7][28] , \mac_out[7][27] , 
        \mac_out[7][26] , \mac_out[7][25] , \mac_out[7][24] , \mac_out[7][23] , 
        \mac_out[7][22] , \mac_out[7][21] , \mac_out[7][20] , \mac_out[7][19] , 
        \mac_out[7][18] , \mac_out[7][17] , \mac_out[7][16] , \mac_out[7][15] , 
        \mac_out[7][14] , \mac_out[7][13] , \mac_out[7][12] , \mac_out[7][11] , 
        \mac_out[7][10] , \mac_out[7][9] , \mac_out[7][8] , \mac_out[7][7] , 
        \mac_out[7][6] , \mac_out[7][5] , \mac_out[7][4] , \mac_out[7][3] , 
        \mac_out[7][2] , \mac_out[7][1] , \mac_out[7][0] }) );
  memory_WIDTH40_SIZE1_LOGSIZE4_7 \y[0]  ( .clk(clk), .data_in({
        \mac_out[0][39] , \mac_out[0][38] , \mac_out[0][37] , \mac_out[0][36] , 
        \mac_out[0][35] , \mac_out[0][34] , \mac_out[0][33] , \mac_out[0][32] , 
        \mac_out[0][31] , \mac_out[0][30] , \mac_out[0][29] , \mac_out[0][28] , 
        \mac_out[0][27] , \mac_out[0][26] , \mac_out[0][25] , \mac_out[0][24] , 
        \mac_out[0][23] , \mac_out[0][22] , \mac_out[0][21] , \mac_out[0][20] , 
        \mac_out[0][19] , \mac_out[0][18] , \mac_out[0][17] , \mac_out[0][16] , 
        \mac_out[0][15] , \mac_out[0][14] , \mac_out[0][13] , \mac_out[0][12] , 
        \mac_out[0][11] , \mac_out[0][10] , \mac_out[0][9] , \mac_out[0][8] , 
        \mac_out[0][7] , \mac_out[0][6] , \mac_out[0][5] , \mac_out[0][4] , 
        \mac_out[0][3] , \mac_out[0][2] , \mac_out[0][1] , \mac_out[0][0] }), 
        .data_out({\mux[0][39] , \mux[0][38] , \mux[0][37] , \mux[0][36] , 
        \mux[0][35] , \mux[0][34] , \mux[0][33] , \mux[0][32] , \mux[0][31] , 
        \mux[0][30] , \mux[0][29] , \mux[0][28] , \mux[0][27] , \mux[0][26] , 
        \mux[0][25] , \mux[0][24] , \mux[0][23] , \mux[0][22] , \mux[0][21] , 
        \mux[0][20] , \mux[0][19] , \mux[0][18] , \mux[0][17] , \mux[0][16] , 
        \mux[0][15] , \mux[0][14] , \mux[0][13] , \mux[0][12] , \mux[0][11] , 
        \mux[0][10] , \mux[0][9] , \mux[0][8] , \mux[0][7] , \mux[0][6] , 
        \mux[0][5] , \mux[0][4] , \mux[0][3] , \mux[0][2] , \mux[0][1] , 
        \mux[0][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(wr_en_y) );
  memory_WIDTH40_SIZE1_LOGSIZE4_6 \y[1]  ( .clk(clk), .data_in({
        \mac_out[1][39] , \mac_out[1][38] , \mac_out[1][37] , \mac_out[1][36] , 
        \mac_out[1][35] , \mac_out[1][34] , \mac_out[1][33] , \mac_out[1][32] , 
        \mac_out[1][31] , \mac_out[1][30] , \mac_out[1][29] , \mac_out[1][28] , 
        \mac_out[1][27] , \mac_out[1][26] , \mac_out[1][25] , \mac_out[1][24] , 
        \mac_out[1][23] , \mac_out[1][22] , \mac_out[1][21] , \mac_out[1][20] , 
        \mac_out[1][19] , \mac_out[1][18] , \mac_out[1][17] , \mac_out[1][16] , 
        \mac_out[1][15] , \mac_out[1][14] , \mac_out[1][13] , \mac_out[1][12] , 
        \mac_out[1][11] , \mac_out[1][10] , \mac_out[1][9] , \mac_out[1][8] , 
        \mac_out[1][7] , \mac_out[1][6] , \mac_out[1][5] , \mac_out[1][4] , 
        \mac_out[1][3] , \mac_out[1][2] , \mac_out[1][1] , \mac_out[1][0] }), 
        .data_out({\mux[1][39] , \mux[1][38] , \mux[1][37] , \mux[1][36] , 
        \mux[1][35] , \mux[1][34] , \mux[1][33] , \mux[1][32] , \mux[1][31] , 
        \mux[1][30] , \mux[1][29] , \mux[1][28] , \mux[1][27] , \mux[1][26] , 
        \mux[1][25] , \mux[1][24] , \mux[1][23] , \mux[1][22] , \mux[1][21] , 
        \mux[1][20] , \mux[1][19] , \mux[1][18] , \mux[1][17] , \mux[1][16] , 
        \mux[1][15] , \mux[1][14] , \mux[1][13] , \mux[1][12] , \mux[1][11] , 
        \mux[1][10] , \mux[1][9] , \mux[1][8] , \mux[1][7] , \mux[1][6] , 
        \mux[1][5] , \mux[1][4] , \mux[1][3] , \mux[1][2] , \mux[1][1] , 
        \mux[1][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(wr_en_y) );
  memory_WIDTH40_SIZE1_LOGSIZE4_5 \y[2]  ( .clk(clk), .data_in({
        \mac_out[2][39] , \mac_out[2][38] , \mac_out[2][37] , \mac_out[2][36] , 
        \mac_out[2][35] , \mac_out[2][34] , \mac_out[2][33] , \mac_out[2][32] , 
        \mac_out[2][31] , \mac_out[2][30] , \mac_out[2][29] , \mac_out[2][28] , 
        \mac_out[2][27] , \mac_out[2][26] , \mac_out[2][25] , \mac_out[2][24] , 
        \mac_out[2][23] , \mac_out[2][22] , \mac_out[2][21] , \mac_out[2][20] , 
        \mac_out[2][19] , \mac_out[2][18] , \mac_out[2][17] , \mac_out[2][16] , 
        \mac_out[2][15] , \mac_out[2][14] , \mac_out[2][13] , \mac_out[2][12] , 
        \mac_out[2][11] , \mac_out[2][10] , \mac_out[2][9] , \mac_out[2][8] , 
        \mac_out[2][7] , \mac_out[2][6] , \mac_out[2][5] , \mac_out[2][4] , 
        \mac_out[2][3] , \mac_out[2][2] , \mac_out[2][1] , \mac_out[2][0] }), 
        .data_out({\mux[2][39] , \mux[2][38] , \mux[2][37] , \mux[2][36] , 
        \mux[2][35] , \mux[2][34] , \mux[2][33] , \mux[2][32] , \mux[2][31] , 
        \mux[2][30] , \mux[2][29] , \mux[2][28] , \mux[2][27] , \mux[2][26] , 
        \mux[2][25] , \mux[2][24] , \mux[2][23] , \mux[2][22] , \mux[2][21] , 
        \mux[2][20] , \mux[2][19] , \mux[2][18] , \mux[2][17] , \mux[2][16] , 
        \mux[2][15] , \mux[2][14] , \mux[2][13] , \mux[2][12] , \mux[2][11] , 
        \mux[2][10] , \mux[2][9] , \mux[2][8] , \mux[2][7] , \mux[2][6] , 
        \mux[2][5] , \mux[2][4] , \mux[2][3] , \mux[2][2] , \mux[2][1] , 
        \mux[2][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(wr_en_y) );
  memory_WIDTH40_SIZE1_LOGSIZE4_4 \y[3]  ( .clk(clk), .data_in({
        \mac_out[3][39] , \mac_out[3][38] , \mac_out[3][37] , \mac_out[3][36] , 
        \mac_out[3][35] , \mac_out[3][34] , \mac_out[3][33] , \mac_out[3][32] , 
        \mac_out[3][31] , \mac_out[3][30] , \mac_out[3][29] , \mac_out[3][28] , 
        \mac_out[3][27] , \mac_out[3][26] , \mac_out[3][25] , \mac_out[3][24] , 
        \mac_out[3][23] , \mac_out[3][22] , \mac_out[3][21] , \mac_out[3][20] , 
        \mac_out[3][19] , \mac_out[3][18] , \mac_out[3][17] , \mac_out[3][16] , 
        \mac_out[3][15] , \mac_out[3][14] , \mac_out[3][13] , \mac_out[3][12] , 
        \mac_out[3][11] , \mac_out[3][10] , \mac_out[3][9] , \mac_out[3][8] , 
        \mac_out[3][7] , \mac_out[3][6] , \mac_out[3][5] , \mac_out[3][4] , 
        \mac_out[3][3] , \mac_out[3][2] , \mac_out[3][1] , \mac_out[3][0] }), 
        .data_out({\mux[3][39] , \mux[3][38] , \mux[3][37] , \mux[3][36] , 
        \mux[3][35] , \mux[3][34] , \mux[3][33] , \mux[3][32] , \mux[3][31] , 
        \mux[3][30] , \mux[3][29] , \mux[3][28] , \mux[3][27] , \mux[3][26] , 
        \mux[3][25] , \mux[3][24] , \mux[3][23] , \mux[3][22] , \mux[3][21] , 
        \mux[3][20] , \mux[3][19] , \mux[3][18] , \mux[3][17] , \mux[3][16] , 
        \mux[3][15] , \mux[3][14] , \mux[3][13] , \mux[3][12] , \mux[3][11] , 
        \mux[3][10] , \mux[3][9] , \mux[3][8] , \mux[3][7] , \mux[3][6] , 
        \mux[3][5] , \mux[3][4] , \mux[3][3] , \mux[3][2] , \mux[3][1] , 
        \mux[3][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(wr_en_y) );
  memory_WIDTH40_SIZE1_LOGSIZE4_3 \y[4]  ( .clk(clk), .data_in({
        \mac_out[4][39] , \mac_out[4][38] , \mac_out[4][37] , \mac_out[4][36] , 
        \mac_out[4][35] , \mac_out[4][34] , \mac_out[4][33] , \mac_out[4][32] , 
        \mac_out[4][31] , \mac_out[4][30] , \mac_out[4][29] , \mac_out[4][28] , 
        \mac_out[4][27] , \mac_out[4][26] , \mac_out[4][25] , \mac_out[4][24] , 
        \mac_out[4][23] , \mac_out[4][22] , \mac_out[4][21] , \mac_out[4][20] , 
        \mac_out[4][19] , \mac_out[4][18] , \mac_out[4][17] , \mac_out[4][16] , 
        \mac_out[4][15] , \mac_out[4][14] , \mac_out[4][13] , \mac_out[4][12] , 
        \mac_out[4][11] , \mac_out[4][10] , \mac_out[4][9] , \mac_out[4][8] , 
        \mac_out[4][7] , \mac_out[4][6] , \mac_out[4][5] , \mac_out[4][4] , 
        \mac_out[4][3] , \mac_out[4][2] , \mac_out[4][1] , \mac_out[4][0] }), 
        .data_out({\mux[4][39] , \mux[4][38] , \mux[4][37] , \mux[4][36] , 
        \mux[4][35] , \mux[4][34] , \mux[4][33] , \mux[4][32] , \mux[4][31] , 
        \mux[4][30] , \mux[4][29] , \mux[4][28] , \mux[4][27] , \mux[4][26] , 
        \mux[4][25] , \mux[4][24] , \mux[4][23] , \mux[4][22] , \mux[4][21] , 
        \mux[4][20] , \mux[4][19] , \mux[4][18] , \mux[4][17] , \mux[4][16] , 
        \mux[4][15] , \mux[4][14] , \mux[4][13] , \mux[4][12] , \mux[4][11] , 
        \mux[4][10] , \mux[4][9] , \mux[4][8] , \mux[4][7] , \mux[4][6] , 
        \mux[4][5] , \mux[4][4] , \mux[4][3] , \mux[4][2] , \mux[4][1] , 
        \mux[4][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(wr_en_y) );
  memory_WIDTH40_SIZE1_LOGSIZE4_2 \y[5]  ( .clk(clk), .data_in({
        \mac_out[5][39] , \mac_out[5][38] , \mac_out[5][37] , \mac_out[5][36] , 
        \mac_out[5][35] , \mac_out[5][34] , \mac_out[5][33] , \mac_out[5][32] , 
        \mac_out[5][31] , \mac_out[5][30] , \mac_out[5][29] , \mac_out[5][28] , 
        \mac_out[5][27] , \mac_out[5][26] , \mac_out[5][25] , \mac_out[5][24] , 
        \mac_out[5][23] , \mac_out[5][22] , \mac_out[5][21] , \mac_out[5][20] , 
        \mac_out[5][19] , \mac_out[5][18] , \mac_out[5][17] , \mac_out[5][16] , 
        \mac_out[5][15] , \mac_out[5][14] , \mac_out[5][13] , \mac_out[5][12] , 
        \mac_out[5][11] , \mac_out[5][10] , \mac_out[5][9] , \mac_out[5][8] , 
        \mac_out[5][7] , \mac_out[5][6] , \mac_out[5][5] , \mac_out[5][4] , 
        \mac_out[5][3] , \mac_out[5][2] , \mac_out[5][1] , \mac_out[5][0] }), 
        .data_out({\mux[5][39] , \mux[5][38] , \mux[5][37] , \mux[5][36] , 
        \mux[5][35] , \mux[5][34] , \mux[5][33] , \mux[5][32] , \mux[5][31] , 
        \mux[5][30] , \mux[5][29] , \mux[5][28] , \mux[5][27] , \mux[5][26] , 
        \mux[5][25] , \mux[5][24] , \mux[5][23] , \mux[5][22] , \mux[5][21] , 
        \mux[5][20] , \mux[5][19] , \mux[5][18] , \mux[5][17] , \mux[5][16] , 
        \mux[5][15] , \mux[5][14] , \mux[5][13] , \mux[5][12] , \mux[5][11] , 
        \mux[5][10] , \mux[5][9] , \mux[5][8] , \mux[5][7] , \mux[5][6] , 
        \mux[5][5] , \mux[5][4] , \mux[5][3] , \mux[5][2] , \mux[5][1] , 
        \mux[5][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(wr_en_y) );
  memory_WIDTH40_SIZE1_LOGSIZE4_1 \y[6]  ( .clk(clk), .data_in({
        \mac_out[6][39] , \mac_out[6][38] , \mac_out[6][37] , \mac_out[6][36] , 
        \mac_out[6][35] , \mac_out[6][34] , \mac_out[6][33] , \mac_out[6][32] , 
        \mac_out[6][31] , \mac_out[6][30] , \mac_out[6][29] , \mac_out[6][28] , 
        \mac_out[6][27] , \mac_out[6][26] , \mac_out[6][25] , \mac_out[6][24] , 
        \mac_out[6][23] , \mac_out[6][22] , \mac_out[6][21] , \mac_out[6][20] , 
        \mac_out[6][19] , \mac_out[6][18] , \mac_out[6][17] , \mac_out[6][16] , 
        \mac_out[6][15] , \mac_out[6][14] , \mac_out[6][13] , \mac_out[6][12] , 
        \mac_out[6][11] , \mac_out[6][10] , \mac_out[6][9] , \mac_out[6][8] , 
        \mac_out[6][7] , \mac_out[6][6] , \mac_out[6][5] , \mac_out[6][4] , 
        \mac_out[6][3] , \mac_out[6][2] , \mac_out[6][1] , \mac_out[6][0] }), 
        .data_out({\mux[6][39] , \mux[6][38] , \mux[6][37] , \mux[6][36] , 
        \mux[6][35] , \mux[6][34] , \mux[6][33] , \mux[6][32] , \mux[6][31] , 
        \mux[6][30] , \mux[6][29] , \mux[6][28] , \mux[6][27] , \mux[6][26] , 
        \mux[6][25] , \mux[6][24] , \mux[6][23] , \mux[6][22] , \mux[6][21] , 
        \mux[6][20] , \mux[6][19] , \mux[6][18] , \mux[6][17] , \mux[6][16] , 
        \mux[6][15] , \mux[6][14] , \mux[6][13] , \mux[6][12] , \mux[6][11] , 
        \mux[6][10] , \mux[6][9] , \mux[6][8] , \mux[6][7] , \mux[6][6] , 
        \mux[6][5] , \mux[6][4] , \mux[6][3] , \mux[6][2] , \mux[6][1] , 
        \mux[6][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(wr_en_y) );
  memory_WIDTH40_SIZE1_LOGSIZE4_0 \y[7]  ( .clk(clk), .data_in({
        \mac_out[7][39] , \mac_out[7][38] , \mac_out[7][37] , \mac_out[7][36] , 
        \mac_out[7][35] , \mac_out[7][34] , \mac_out[7][33] , \mac_out[7][32] , 
        \mac_out[7][31] , \mac_out[7][30] , \mac_out[7][29] , \mac_out[7][28] , 
        \mac_out[7][27] , \mac_out[7][26] , \mac_out[7][25] , \mac_out[7][24] , 
        \mac_out[7][23] , \mac_out[7][22] , \mac_out[7][21] , \mac_out[7][20] , 
        \mac_out[7][19] , \mac_out[7][18] , \mac_out[7][17] , \mac_out[7][16] , 
        \mac_out[7][15] , \mac_out[7][14] , \mac_out[7][13] , \mac_out[7][12] , 
        \mac_out[7][11] , \mac_out[7][10] , \mac_out[7][9] , \mac_out[7][8] , 
        \mac_out[7][7] , \mac_out[7][6] , \mac_out[7][5] , \mac_out[7][4] , 
        \mac_out[7][3] , \mac_out[7][2] , \mac_out[7][1] , \mac_out[7][0] }), 
        .data_out({\mux[7][39] , \mux[7][38] , \mux[7][37] , \mux[7][36] , 
        \mux[7][35] , \mux[7][34] , \mux[7][33] , \mux[7][32] , \mux[7][31] , 
        \mux[7][30] , \mux[7][29] , \mux[7][28] , \mux[7][27] , \mux[7][26] , 
        \mux[7][25] , \mux[7][24] , \mux[7][23] , \mux[7][22] , \mux[7][21] , 
        \mux[7][20] , \mux[7][19] , \mux[7][18] , \mux[7][17] , \mux[7][16] , 
        \mux[7][15] , \mux[7][14] , \mux[7][13] , \mux[7][12] , \mux[7][11] , 
        \mux[7][10] , \mux[7][9] , \mux[7][8] , \mux[7][7] , \mux[7][6] , 
        \mux[7][5] , \mux[7][4] , \mux[7][3] , \mux[7][2] , \mux[7][1] , 
        \mux[7][0] }), .addr({1'b0, 1'b0, 1'b0, 1'b0}), .wr_en(wr_en_y) );
  CLKBUF_X3 U2 ( .A(vector_out[10]), .Z(n283) );
  BUF_X2 U3 ( .A(vector_out[15]), .Z(n295) );
  BUF_X1 U4 ( .A(vector_out[12]), .Z(n290) );
  BUF_X1 U5 ( .A(vector_out[1]), .Z(n265) );
  BUF_X1 U6 ( .A(vector_out[11]), .Z(n287) );
  BUF_X2 U7 ( .A(vector_out[16]), .Z(n297) );
  BUF_X2 U8 ( .A(vector_out[10]), .Z(n282) );
  BUF_X1 U9 ( .A(vector_out[7]), .Z(n273) );
  BUF_X1 U10 ( .A(vector_out[18]), .Z(n301) );
  BUF_X1 U11 ( .A(vector_out[12]), .Z(n289) );
  BUF_X2 U12 ( .A(vector_out[4]), .Z(n5) );
  BUF_X1 U13 ( .A(vector_out[18]), .Z(n300) );
  BUF_X1 U14 ( .A(vector_out[1]), .Z(n264) );
  BUF_X2 U15 ( .A(vector_out[5]), .Z(n2) );
  BUF_X2 U16 ( .A(vector_out[0]), .Z(n9) );
  BUF_X1 U17 ( .A(vector_out[5]), .Z(n1) );
  BUF_X1 U18 ( .A(vector_out[5]), .Z(n3) );
  BUF_X1 U19 ( .A(vector_out[19]), .Z(n305) );
  BUF_X1 U20 ( .A(vector_out[9]), .Z(n280) );
  BUF_X1 U21 ( .A(vector_out[13]), .Z(n292) );
  BUF_X2 U22 ( .A(vector_out[2]), .Z(n266) );
  BUF_X1 U23 ( .A(vector_out[1]), .Z(n4) );
  BUF_X1 U24 ( .A(vector_out[3]), .Z(n268) );
  BUF_X1 U25 ( .A(vector_out[11]), .Z(n286) );
  CLKBUF_X1 U26 ( .A(vector_out[3]), .Z(n269) );
  CLKBUF_X3 U27 ( .A(vector_out[3]), .Z(n7) );
  BUF_X1 U28 ( .A(vector_out[1]), .Z(n263) );
  CLKBUF_X1 U29 ( .A(vector_out[8]), .Z(n6) );
  CLKBUF_X1 U30 ( .A(vector_out[8]), .Z(n278) );
  CLKBUF_X3 U31 ( .A(vector_out[2]), .Z(n267) );
  BUF_X1 U32 ( .A(vector_out[7]), .Z(n274) );
  BUF_X2 U33 ( .A(vector_out[0]), .Z(n8) );
  BUF_X1 U34 ( .A(vector_out[7]), .Z(n275) );
  BUF_X1 U35 ( .A(vector_out[10]), .Z(n284) );
  BUF_X2 U36 ( .A(vector_out[6]), .Z(n271) );
  BUF_X1 U37 ( .A(vector_out[14]), .Z(n293) );
  BUF_X2 U38 ( .A(vector_out[4]), .Z(n270) );
  BUF_X2 U39 ( .A(vector_out[19]), .Z(n303) );
  BUF_X1 U40 ( .A(vector_out[12]), .Z(n288) );
  BUF_X2 U41 ( .A(vector_out[9]), .Z(n279) );
  BUF_X1 U42 ( .A(vector_out[8]), .Z(n276) );
  CLKBUF_X1 U43 ( .A(vector_out[18]), .Z(n302) );
  BUF_X1 U44 ( .A(vector_out[15]), .Z(n296) );
  BUF_X1 U45 ( .A(vector_out[11]), .Z(n285) );
  BUF_X1 U46 ( .A(vector_out[16]), .Z(n298) );
  BUF_X1 U47 ( .A(vector_out[13]), .Z(n291) );
  BUF_X1 U48 ( .A(n262), .Z(n259) );
  BUF_X1 U49 ( .A(n262), .Z(n260) );
  BUF_X1 U50 ( .A(n262), .Z(n261) );
  BUF_X1 U51 ( .A(addr_y[1]), .Z(n252) );
  BUF_X1 U52 ( .A(addr_y[1]), .Z(n253) );
  BUF_X1 U53 ( .A(addr_y[1]), .Z(n254) );
  BUF_X1 U54 ( .A(addr_y[1]), .Z(n255) );
  BUF_X1 U55 ( .A(n262), .Z(n256) );
  BUF_X1 U56 ( .A(n262), .Z(n257) );
  BUF_X1 U57 ( .A(n262), .Z(n258) );
  BUF_X1 U58 ( .A(n251), .Z(n250) );
  BUF_X1 U59 ( .A(addr_y[0]), .Z(n262) );
  BUF_X1 U60 ( .A(addr_y[2]), .Z(n251) );
  BUF_X1 U61 ( .A(vector_out[19]), .Z(n304) );
  BUF_X1 U62 ( .A(vector_out[8]), .Z(n277) );
  BUF_X1 U63 ( .A(vector_out[14]), .Z(n294) );
  BUF_X1 U64 ( .A(vector_out[6]), .Z(n272) );
  CLKBUF_X1 U65 ( .A(vector_out[9]), .Z(n281) );
  BUF_X1 U66 ( .A(vector_out[16]), .Z(n299) );
  MUX2_X1 U67 ( .A(\mux[6][0] ), .B(\mux[7][0] ), .S(n259), .Z(n10) );
  MUX2_X1 U68 ( .A(\mux[4][0] ), .B(\mux[5][0] ), .S(n258), .Z(n11) );
  MUX2_X1 U69 ( .A(n11), .B(n10), .S(addr_y[1]), .Z(n12) );
  MUX2_X1 U70 ( .A(\mux[2][0] ), .B(\mux[3][0] ), .S(n262), .Z(n13) );
  MUX2_X1 U71 ( .A(\mux[0][0] ), .B(\mux[1][0] ), .S(n259), .Z(n14) );
  MUX2_X1 U72 ( .A(n14), .B(n13), .S(addr_y[1]), .Z(n15) );
  MUX2_X1 U73 ( .A(n15), .B(n12), .S(n250), .Z(data_out[0]) );
  MUX2_X1 U74 ( .A(\mux[6][1] ), .B(\mux[7][1] ), .S(n257), .Z(n16) );
  MUX2_X1 U75 ( .A(\mux[4][1] ), .B(\mux[5][1] ), .S(n258), .Z(n17) );
  MUX2_X1 U76 ( .A(n17), .B(n16), .S(addr_y[1]), .Z(n18) );
  MUX2_X1 U77 ( .A(\mux[2][1] ), .B(\mux[3][1] ), .S(n259), .Z(n19) );
  MUX2_X1 U78 ( .A(\mux[0][1] ), .B(\mux[1][1] ), .S(n262), .Z(n20) );
  MUX2_X1 U79 ( .A(n20), .B(n19), .S(addr_y[1]), .Z(n21) );
  MUX2_X1 U80 ( .A(n21), .B(n18), .S(n251), .Z(data_out[1]) );
  MUX2_X1 U81 ( .A(\mux[6][2] ), .B(\mux[7][2] ), .S(n260), .Z(n22) );
  MUX2_X1 U82 ( .A(\mux[4][2] ), .B(\mux[5][2] ), .S(n259), .Z(n23) );
  MUX2_X1 U83 ( .A(n23), .B(n22), .S(addr_y[1]), .Z(n24) );
  MUX2_X1 U84 ( .A(\mux[2][2] ), .B(\mux[3][2] ), .S(n260), .Z(n25) );
  MUX2_X1 U85 ( .A(\mux[0][2] ), .B(\mux[1][2] ), .S(n261), .Z(n26) );
  MUX2_X1 U86 ( .A(n26), .B(n25), .S(addr_y[1]), .Z(n27) );
  MUX2_X1 U87 ( .A(n27), .B(n24), .S(n250), .Z(data_out[2]) );
  MUX2_X1 U88 ( .A(\mux[6][3] ), .B(\mux[7][3] ), .S(n256), .Z(n28) );
  MUX2_X1 U89 ( .A(\mux[4][3] ), .B(\mux[5][3] ), .S(n257), .Z(n29) );
  MUX2_X1 U90 ( .A(n29), .B(n28), .S(addr_y[1]), .Z(n30) );
  MUX2_X1 U91 ( .A(\mux[2][3] ), .B(\mux[3][3] ), .S(n258), .Z(n31) );
  MUX2_X1 U92 ( .A(\mux[0][3] ), .B(\mux[1][3] ), .S(n262), .Z(n32) );
  MUX2_X1 U93 ( .A(n32), .B(n31), .S(n252), .Z(n33) );
  MUX2_X1 U94 ( .A(n33), .B(n30), .S(n251), .Z(data_out[3]) );
  MUX2_X1 U95 ( .A(\mux[6][4] ), .B(\mux[7][4] ), .S(n259), .Z(n34) );
  MUX2_X1 U96 ( .A(\mux[4][4] ), .B(\mux[5][4] ), .S(n260), .Z(n35) );
  MUX2_X1 U97 ( .A(n35), .B(n34), .S(n252), .Z(n36) );
  MUX2_X1 U98 ( .A(\mux[2][4] ), .B(\mux[3][4] ), .S(n257), .Z(n37) );
  MUX2_X1 U99 ( .A(\mux[0][4] ), .B(\mux[1][4] ), .S(n262), .Z(n38) );
  MUX2_X1 U100 ( .A(n38), .B(n37), .S(n252), .Z(n39) );
  MUX2_X1 U101 ( .A(n39), .B(n36), .S(n250), .Z(data_out[4]) );
  MUX2_X1 U102 ( .A(\mux[6][5] ), .B(\mux[7][5] ), .S(addr_y[0]), .Z(n40) );
  MUX2_X1 U103 ( .A(\mux[4][5] ), .B(\mux[5][5] ), .S(n258), .Z(n41) );
  MUX2_X1 U104 ( .A(n41), .B(n40), .S(n252), .Z(n42) );
  MUX2_X1 U105 ( .A(\mux[2][5] ), .B(\mux[3][5] ), .S(n262), .Z(n43) );
  MUX2_X1 U106 ( .A(\mux[0][5] ), .B(\mux[1][5] ), .S(n261), .Z(n44) );
  MUX2_X1 U107 ( .A(n44), .B(n43), .S(n252), .Z(n45) );
  MUX2_X1 U108 ( .A(n45), .B(n42), .S(n250), .Z(data_out[5]) );
  MUX2_X1 U109 ( .A(\mux[6][6] ), .B(\mux[7][6] ), .S(n262), .Z(n46) );
  MUX2_X1 U110 ( .A(\mux[4][6] ), .B(\mux[5][6] ), .S(addr_y[0]), .Z(n47) );
  MUX2_X1 U111 ( .A(n47), .B(n46), .S(n252), .Z(n48) );
  MUX2_X1 U112 ( .A(\mux[2][6] ), .B(\mux[3][6] ), .S(n262), .Z(n49) );
  MUX2_X1 U113 ( .A(\mux[0][6] ), .B(\mux[1][6] ), .S(n259), .Z(n50) );
  MUX2_X1 U114 ( .A(n50), .B(n49), .S(n252), .Z(n51) );
  MUX2_X1 U115 ( .A(n51), .B(n48), .S(n250), .Z(data_out[6]) );
  MUX2_X1 U116 ( .A(\mux[6][7] ), .B(\mux[7][7] ), .S(n259), .Z(n52) );
  MUX2_X1 U117 ( .A(\mux[4][7] ), .B(\mux[5][7] ), .S(addr_y[0]), .Z(n53) );
  MUX2_X1 U118 ( .A(n53), .B(n52), .S(n252), .Z(n54) );
  MUX2_X1 U119 ( .A(\mux[2][7] ), .B(\mux[3][7] ), .S(n256), .Z(n55) );
  MUX2_X1 U120 ( .A(\mux[0][7] ), .B(\mux[1][7] ), .S(n260), .Z(n56) );
  MUX2_X1 U121 ( .A(n56), .B(n55), .S(n252), .Z(n57) );
  MUX2_X1 U122 ( .A(n57), .B(n54), .S(n250), .Z(data_out[7]) );
  MUX2_X1 U123 ( .A(\mux[6][8] ), .B(\mux[7][8] ), .S(n260), .Z(n58) );
  MUX2_X1 U124 ( .A(\mux[4][8] ), .B(\mux[5][8] ), .S(n262), .Z(n59) );
  MUX2_X1 U125 ( .A(n59), .B(n58), .S(n252), .Z(n60) );
  MUX2_X1 U126 ( .A(\mux[2][8] ), .B(\mux[3][8] ), .S(addr_y[0]), .Z(n61) );
  MUX2_X1 U127 ( .A(\mux[0][8] ), .B(\mux[1][8] ), .S(n257), .Z(n62) );
  MUX2_X1 U128 ( .A(n62), .B(n61), .S(n252), .Z(n63) );
  MUX2_X1 U129 ( .A(n63), .B(n60), .S(n250), .Z(data_out[8]) );
  MUX2_X1 U130 ( .A(\mux[6][9] ), .B(\mux[7][9] ), .S(n261), .Z(n64) );
  MUX2_X1 U131 ( .A(\mux[4][9] ), .B(\mux[5][9] ), .S(n261), .Z(n65) );
  MUX2_X1 U132 ( .A(n65), .B(n64), .S(n252), .Z(n66) );
  MUX2_X1 U133 ( .A(\mux[2][9] ), .B(\mux[3][9] ), .S(n262), .Z(n67) );
  MUX2_X1 U134 ( .A(\mux[0][9] ), .B(\mux[1][9] ), .S(addr_y[0]), .Z(n68) );
  MUX2_X1 U135 ( .A(n68), .B(n67), .S(n252), .Z(n69) );
  MUX2_X1 U136 ( .A(n69), .B(n66), .S(n250), .Z(data_out[9]) );
  MUX2_X1 U137 ( .A(\mux[6][10] ), .B(\mux[7][10] ), .S(n256), .Z(n70) );
  MUX2_X1 U138 ( .A(\mux[4][10] ), .B(\mux[5][10] ), .S(addr_y[0]), .Z(n71) );
  MUX2_X1 U139 ( .A(n71), .B(n70), .S(n253), .Z(n72) );
  MUX2_X1 U140 ( .A(\mux[2][10] ), .B(\mux[3][10] ), .S(n257), .Z(n73) );
  MUX2_X1 U141 ( .A(\mux[0][10] ), .B(\mux[1][10] ), .S(addr_y[0]), .Z(n74) );
  MUX2_X1 U142 ( .A(n74), .B(n73), .S(n253), .Z(n75) );
  MUX2_X1 U143 ( .A(n75), .B(n72), .S(n250), .Z(data_out[10]) );
  MUX2_X1 U144 ( .A(\mux[6][11] ), .B(\mux[7][11] ), .S(n256), .Z(n76) );
  MUX2_X1 U145 ( .A(\mux[4][11] ), .B(\mux[5][11] ), .S(n258), .Z(n77) );
  MUX2_X1 U146 ( .A(n77), .B(n76), .S(n253), .Z(n78) );
  MUX2_X1 U147 ( .A(\mux[2][11] ), .B(\mux[3][11] ), .S(n262), .Z(n79) );
  MUX2_X1 U148 ( .A(\mux[0][11] ), .B(\mux[1][11] ), .S(addr_y[0]), .Z(n80) );
  MUX2_X1 U149 ( .A(n80), .B(n79), .S(n253), .Z(n81) );
  MUX2_X1 U150 ( .A(n81), .B(n78), .S(n250), .Z(data_out[11]) );
  MUX2_X1 U151 ( .A(\mux[6][12] ), .B(\mux[7][12] ), .S(n258), .Z(n82) );
  MUX2_X1 U152 ( .A(\mux[4][12] ), .B(\mux[5][12] ), .S(n257), .Z(n83) );
  MUX2_X1 U153 ( .A(n83), .B(n82), .S(n253), .Z(n84) );
  MUX2_X1 U154 ( .A(\mux[2][12] ), .B(\mux[3][12] ), .S(n262), .Z(n85) );
  MUX2_X1 U155 ( .A(\mux[0][12] ), .B(\mux[1][12] ), .S(n262), .Z(n86) );
  MUX2_X1 U156 ( .A(n86), .B(n85), .S(n253), .Z(n87) );
  MUX2_X1 U157 ( .A(n87), .B(n84), .S(n250), .Z(data_out[12]) );
  MUX2_X1 U158 ( .A(\mux[6][13] ), .B(\mux[7][13] ), .S(n262), .Z(n88) );
  MUX2_X1 U159 ( .A(\mux[4][13] ), .B(\mux[5][13] ), .S(n259), .Z(n89) );
  MUX2_X1 U160 ( .A(n89), .B(n88), .S(n253), .Z(n90) );
  MUX2_X1 U161 ( .A(\mux[2][13] ), .B(\mux[3][13] ), .S(n260), .Z(n91) );
  MUX2_X1 U162 ( .A(\mux[0][13] ), .B(\mux[1][13] ), .S(n261), .Z(n92) );
  MUX2_X1 U163 ( .A(n92), .B(n91), .S(n253), .Z(n93) );
  MUX2_X1 U164 ( .A(n93), .B(n90), .S(n250), .Z(data_out[13]) );
  MUX2_X1 U165 ( .A(\mux[6][14] ), .B(\mux[7][14] ), .S(n256), .Z(n94) );
  MUX2_X1 U166 ( .A(\mux[4][14] ), .B(\mux[5][14] ), .S(n257), .Z(n95) );
  MUX2_X1 U167 ( .A(n95), .B(n94), .S(n253), .Z(n96) );
  MUX2_X1 U168 ( .A(\mux[2][14] ), .B(\mux[3][14] ), .S(n258), .Z(n97) );
  MUX2_X1 U169 ( .A(\mux[0][14] ), .B(\mux[1][14] ), .S(n260), .Z(n98) );
  MUX2_X1 U170 ( .A(n98), .B(n97), .S(n253), .Z(n99) );
  MUX2_X1 U171 ( .A(n99), .B(n96), .S(n250), .Z(data_out[14]) );
  MUX2_X1 U172 ( .A(\mux[6][15] ), .B(\mux[7][15] ), .S(n261), .Z(n100) );
  MUX2_X1 U173 ( .A(\mux[4][15] ), .B(\mux[5][15] ), .S(n260), .Z(n101) );
  MUX2_X1 U174 ( .A(n101), .B(n100), .S(n253), .Z(n102) );
  MUX2_X1 U175 ( .A(\mux[2][15] ), .B(\mux[3][15] ), .S(addr_y[0]), .Z(n103)
         );
  MUX2_X1 U176 ( .A(\mux[0][15] ), .B(\mux[1][15] ), .S(n262), .Z(n104) );
  MUX2_X1 U177 ( .A(n104), .B(n103), .S(n253), .Z(n105) );
  MUX2_X1 U178 ( .A(n105), .B(n102), .S(n250), .Z(data_out[15]) );
  MUX2_X1 U179 ( .A(\mux[6][16] ), .B(\mux[7][16] ), .S(n261), .Z(n106) );
  MUX2_X1 U180 ( .A(\mux[4][16] ), .B(\mux[5][16] ), .S(n259), .Z(n107) );
  MUX2_X1 U181 ( .A(n107), .B(n106), .S(n254), .Z(n108) );
  MUX2_X1 U182 ( .A(\mux[2][16] ), .B(\mux[3][16] ), .S(n259), .Z(n109) );
  MUX2_X1 U183 ( .A(\mux[0][16] ), .B(\mux[1][16] ), .S(n260), .Z(n110) );
  MUX2_X1 U184 ( .A(n110), .B(n109), .S(n254), .Z(n111) );
  MUX2_X1 U185 ( .A(n111), .B(n108), .S(addr_y[2]), .Z(data_out[16]) );
  MUX2_X1 U186 ( .A(\mux[6][17] ), .B(\mux[7][17] ), .S(n261), .Z(n112) );
  MUX2_X1 U187 ( .A(\mux[4][17] ), .B(\mux[5][17] ), .S(n256), .Z(n113) );
  MUX2_X1 U188 ( .A(n113), .B(n112), .S(n254), .Z(n114) );
  MUX2_X1 U189 ( .A(\mux[2][17] ), .B(\mux[3][17] ), .S(n257), .Z(n115) );
  MUX2_X1 U190 ( .A(\mux[0][17] ), .B(\mux[1][17] ), .S(n258), .Z(n116) );
  MUX2_X1 U191 ( .A(n116), .B(n115), .S(n254), .Z(n117) );
  MUX2_X1 U192 ( .A(n117), .B(n114), .S(addr_y[2]), .Z(data_out[17]) );
  MUX2_X1 U193 ( .A(\mux[6][18] ), .B(\mux[7][18] ), .S(n261), .Z(n118) );
  MUX2_X1 U194 ( .A(\mux[4][18] ), .B(\mux[5][18] ), .S(n258), .Z(n119) );
  MUX2_X1 U195 ( .A(n119), .B(n118), .S(n254), .Z(n120) );
  MUX2_X1 U196 ( .A(\mux[2][18] ), .B(\mux[3][18] ), .S(n260), .Z(n121) );
  MUX2_X1 U197 ( .A(\mux[0][18] ), .B(\mux[1][18] ), .S(n256), .Z(n122) );
  MUX2_X1 U198 ( .A(n122), .B(n121), .S(n254), .Z(n123) );
  MUX2_X1 U199 ( .A(n123), .B(n120), .S(n251), .Z(data_out[18]) );
  MUX2_X1 U200 ( .A(\mux[6][19] ), .B(\mux[7][19] ), .S(n256), .Z(n124) );
  MUX2_X1 U201 ( .A(\mux[4][19] ), .B(\mux[5][19] ), .S(n257), .Z(n125) );
  MUX2_X1 U202 ( .A(n125), .B(n124), .S(n254), .Z(n126) );
  MUX2_X1 U203 ( .A(\mux[2][19] ), .B(\mux[3][19] ), .S(n262), .Z(n127) );
  MUX2_X1 U204 ( .A(\mux[0][19] ), .B(\mux[1][19] ), .S(addr_y[0]), .Z(n128)
         );
  MUX2_X1 U205 ( .A(n128), .B(n127), .S(n254), .Z(n129) );
  MUX2_X1 U206 ( .A(n129), .B(n126), .S(n251), .Z(data_out[19]) );
  MUX2_X1 U207 ( .A(\mux[6][20] ), .B(\mux[7][20] ), .S(n257), .Z(n130) );
  MUX2_X1 U208 ( .A(\mux[4][20] ), .B(\mux[5][20] ), .S(n261), .Z(n131) );
  MUX2_X1 U209 ( .A(n131), .B(n130), .S(n254), .Z(n132) );
  MUX2_X1 U210 ( .A(\mux[2][20] ), .B(\mux[3][20] ), .S(n258), .Z(n133) );
  MUX2_X1 U211 ( .A(\mux[0][20] ), .B(\mux[1][20] ), .S(n262), .Z(n134) );
  MUX2_X1 U212 ( .A(n134), .B(n133), .S(n254), .Z(n135) );
  MUX2_X1 U213 ( .A(n135), .B(n132), .S(addr_y[2]), .Z(data_out[20]) );
  MUX2_X1 U214 ( .A(\mux[6][21] ), .B(\mux[7][21] ), .S(n262), .Z(n136) );
  MUX2_X1 U215 ( .A(\mux[4][21] ), .B(\mux[5][21] ), .S(n256), .Z(n137) );
  MUX2_X1 U216 ( .A(n137), .B(n136), .S(n254), .Z(n138) );
  MUX2_X1 U217 ( .A(\mux[2][21] ), .B(\mux[3][21] ), .S(n256), .Z(n139) );
  MUX2_X1 U218 ( .A(\mux[0][21] ), .B(\mux[1][21] ), .S(n262), .Z(n140) );
  MUX2_X1 U219 ( .A(n140), .B(n139), .S(n254), .Z(n141) );
  MUX2_X1 U220 ( .A(n141), .B(n138), .S(n251), .Z(data_out[21]) );
  MUX2_X1 U221 ( .A(\mux[6][22] ), .B(\mux[7][22] ), .S(n256), .Z(n142) );
  MUX2_X1 U222 ( .A(\mux[4][22] ), .B(\mux[5][22] ), .S(n256), .Z(n143) );
  MUX2_X1 U223 ( .A(n143), .B(n142), .S(n255), .Z(n144) );
  MUX2_X1 U224 ( .A(\mux[2][22] ), .B(\mux[3][22] ), .S(n256), .Z(n145) );
  MUX2_X1 U225 ( .A(\mux[0][22] ), .B(\mux[1][22] ), .S(n256), .Z(n146) );
  MUX2_X1 U226 ( .A(n146), .B(n145), .S(n255), .Z(n147) );
  MUX2_X1 U227 ( .A(n147), .B(n144), .S(addr_y[2]), .Z(data_out[22]) );
  MUX2_X1 U228 ( .A(\mux[6][23] ), .B(\mux[7][23] ), .S(n256), .Z(n148) );
  MUX2_X1 U229 ( .A(\mux[4][23] ), .B(\mux[5][23] ), .S(n256), .Z(n149) );
  MUX2_X1 U230 ( .A(n149), .B(n148), .S(n255), .Z(n150) );
  MUX2_X1 U231 ( .A(\mux[2][23] ), .B(\mux[3][23] ), .S(n256), .Z(n151) );
  MUX2_X1 U232 ( .A(\mux[0][23] ), .B(\mux[1][23] ), .S(n256), .Z(n152) );
  MUX2_X1 U233 ( .A(n152), .B(n151), .S(n255), .Z(n153) );
  MUX2_X1 U234 ( .A(n153), .B(n150), .S(addr_y[2]), .Z(data_out[23]) );
  MUX2_X1 U235 ( .A(\mux[6][24] ), .B(\mux[7][24] ), .S(n256), .Z(n154) );
  MUX2_X1 U236 ( .A(\mux[4][24] ), .B(\mux[5][24] ), .S(n256), .Z(n155) );
  MUX2_X1 U237 ( .A(n155), .B(n154), .S(n255), .Z(n156) );
  MUX2_X1 U238 ( .A(\mux[2][24] ), .B(\mux[3][24] ), .S(n256), .Z(n157) );
  MUX2_X1 U239 ( .A(\mux[0][24] ), .B(\mux[1][24] ), .S(n256), .Z(n158) );
  MUX2_X1 U240 ( .A(n158), .B(n157), .S(n255), .Z(n159) );
  MUX2_X1 U241 ( .A(n159), .B(n156), .S(addr_y[2]), .Z(data_out[24]) );
  MUX2_X1 U242 ( .A(\mux[6][25] ), .B(\mux[7][25] ), .S(n257), .Z(n160) );
  MUX2_X1 U243 ( .A(\mux[4][25] ), .B(\mux[5][25] ), .S(n257), .Z(n161) );
  MUX2_X1 U244 ( .A(n161), .B(n160), .S(n255), .Z(n162) );
  MUX2_X1 U245 ( .A(\mux[2][25] ), .B(\mux[3][25] ), .S(n257), .Z(n163) );
  MUX2_X1 U246 ( .A(\mux[0][25] ), .B(\mux[1][25] ), .S(n257), .Z(n164) );
  MUX2_X1 U247 ( .A(n164), .B(n163), .S(n255), .Z(n165) );
  MUX2_X1 U248 ( .A(n165), .B(n162), .S(n251), .Z(data_out[25]) );
  MUX2_X1 U249 ( .A(\mux[6][26] ), .B(\mux[7][26] ), .S(n257), .Z(n166) );
  MUX2_X1 U250 ( .A(\mux[4][26] ), .B(\mux[5][26] ), .S(n257), .Z(n167) );
  MUX2_X1 U251 ( .A(n167), .B(n166), .S(n255), .Z(n168) );
  MUX2_X1 U252 ( .A(\mux[2][26] ), .B(\mux[3][26] ), .S(n257), .Z(n169) );
  MUX2_X1 U253 ( .A(\mux[0][26] ), .B(\mux[1][26] ), .S(n257), .Z(n170) );
  MUX2_X1 U254 ( .A(n170), .B(n169), .S(n255), .Z(n171) );
  MUX2_X1 U255 ( .A(n171), .B(n168), .S(n251), .Z(data_out[26]) );
  MUX2_X1 U256 ( .A(\mux[6][27] ), .B(\mux[7][27] ), .S(n257), .Z(n172) );
  MUX2_X1 U257 ( .A(\mux[4][27] ), .B(\mux[5][27] ), .S(n257), .Z(n173) );
  MUX2_X1 U258 ( .A(n173), .B(n172), .S(n255), .Z(n174) );
  MUX2_X1 U259 ( .A(\mux[2][27] ), .B(\mux[3][27] ), .S(n257), .Z(n175) );
  MUX2_X1 U260 ( .A(\mux[0][27] ), .B(\mux[1][27] ), .S(n257), .Z(n176) );
  MUX2_X1 U261 ( .A(n176), .B(n175), .S(n255), .Z(n177) );
  MUX2_X1 U262 ( .A(n177), .B(n174), .S(n251), .Z(data_out[27]) );
  MUX2_X1 U263 ( .A(\mux[6][28] ), .B(\mux[7][28] ), .S(n258), .Z(n178) );
  MUX2_X1 U264 ( .A(\mux[4][28] ), .B(\mux[5][28] ), .S(n258), .Z(n179) );
  MUX2_X1 U265 ( .A(n179), .B(n178), .S(addr_y[1]), .Z(n180) );
  MUX2_X1 U266 ( .A(\mux[2][28] ), .B(\mux[3][28] ), .S(n258), .Z(n181) );
  MUX2_X1 U267 ( .A(\mux[0][28] ), .B(\mux[1][28] ), .S(n258), .Z(n182) );
  MUX2_X1 U268 ( .A(n182), .B(n181), .S(n255), .Z(n183) );
  MUX2_X1 U269 ( .A(n183), .B(n180), .S(n251), .Z(data_out[28]) );
  MUX2_X1 U270 ( .A(\mux[6][29] ), .B(\mux[7][29] ), .S(n258), .Z(n184) );
  MUX2_X1 U271 ( .A(\mux[4][29] ), .B(\mux[5][29] ), .S(n258), .Z(n185) );
  MUX2_X1 U272 ( .A(n185), .B(n184), .S(n252), .Z(n186) );
  MUX2_X1 U273 ( .A(\mux[2][29] ), .B(\mux[3][29] ), .S(n258), .Z(n187) );
  MUX2_X1 U274 ( .A(\mux[0][29] ), .B(\mux[1][29] ), .S(n258), .Z(n188) );
  MUX2_X1 U275 ( .A(n188), .B(n187), .S(n253), .Z(n189) );
  MUX2_X1 U276 ( .A(n189), .B(n186), .S(n251), .Z(data_out[29]) );
  MUX2_X1 U277 ( .A(\mux[6][30] ), .B(\mux[7][30] ), .S(n258), .Z(n190) );
  MUX2_X1 U278 ( .A(\mux[4][30] ), .B(\mux[5][30] ), .S(n258), .Z(n191) );
  MUX2_X1 U279 ( .A(n191), .B(n190), .S(n254), .Z(n192) );
  MUX2_X1 U280 ( .A(\mux[2][30] ), .B(\mux[3][30] ), .S(n258), .Z(n193) );
  MUX2_X1 U281 ( .A(\mux[0][30] ), .B(\mux[1][30] ), .S(n258), .Z(n194) );
  MUX2_X1 U282 ( .A(n194), .B(n193), .S(n255), .Z(n195) );
  MUX2_X1 U283 ( .A(n195), .B(n192), .S(addr_y[2]), .Z(data_out[30]) );
  MUX2_X1 U284 ( .A(\mux[6][31] ), .B(\mux[7][31] ), .S(n259), .Z(n196) );
  MUX2_X1 U285 ( .A(\mux[4][31] ), .B(\mux[5][31] ), .S(n259), .Z(n197) );
  MUX2_X1 U286 ( .A(n197), .B(n196), .S(n252), .Z(n198) );
  MUX2_X1 U287 ( .A(\mux[2][31] ), .B(\mux[3][31] ), .S(n259), .Z(n199) );
  MUX2_X1 U288 ( .A(\mux[0][31] ), .B(\mux[1][31] ), .S(n259), .Z(n200) );
  MUX2_X1 U289 ( .A(n200), .B(n199), .S(n253), .Z(n201) );
  MUX2_X1 U290 ( .A(n201), .B(n198), .S(addr_y[2]), .Z(data_out[31]) );
  MUX2_X1 U291 ( .A(\mux[6][32] ), .B(\mux[7][32] ), .S(n259), .Z(n202) );
  MUX2_X1 U292 ( .A(\mux[4][32] ), .B(\mux[5][32] ), .S(n259), .Z(n203) );
  MUX2_X1 U293 ( .A(n203), .B(n202), .S(n254), .Z(n204) );
  MUX2_X1 U294 ( .A(\mux[2][32] ), .B(\mux[3][32] ), .S(n259), .Z(n205) );
  MUX2_X1 U295 ( .A(\mux[0][32] ), .B(\mux[1][32] ), .S(n259), .Z(n206) );
  MUX2_X1 U296 ( .A(n206), .B(n205), .S(n255), .Z(n207) );
  MUX2_X1 U297 ( .A(n207), .B(n204), .S(n251), .Z(data_out[32]) );
  MUX2_X1 U298 ( .A(\mux[6][33] ), .B(\mux[7][33] ), .S(n259), .Z(n208) );
  MUX2_X1 U299 ( .A(\mux[4][33] ), .B(\mux[5][33] ), .S(n259), .Z(n209) );
  MUX2_X1 U300 ( .A(n209), .B(n208), .S(n252), .Z(n210) );
  MUX2_X1 U301 ( .A(\mux[2][33] ), .B(\mux[3][33] ), .S(n259), .Z(n211) );
  MUX2_X1 U302 ( .A(\mux[0][33] ), .B(\mux[1][33] ), .S(n259), .Z(n212) );
  MUX2_X1 U303 ( .A(n212), .B(n211), .S(n253), .Z(n213) );
  MUX2_X1 U304 ( .A(n213), .B(n210), .S(addr_y[2]), .Z(data_out[33]) );
  MUX2_X1 U305 ( .A(\mux[6][34] ), .B(\mux[7][34] ), .S(n260), .Z(n214) );
  MUX2_X1 U306 ( .A(\mux[4][34] ), .B(\mux[5][34] ), .S(n260), .Z(n215) );
  MUX2_X1 U307 ( .A(n215), .B(n214), .S(n253), .Z(n216) );
  MUX2_X1 U308 ( .A(\mux[2][34] ), .B(\mux[3][34] ), .S(n260), .Z(n217) );
  MUX2_X1 U309 ( .A(\mux[0][34] ), .B(\mux[1][34] ), .S(n260), .Z(n218) );
  MUX2_X1 U310 ( .A(n218), .B(n217), .S(n254), .Z(n219) );
  MUX2_X1 U311 ( .A(n219), .B(n216), .S(n250), .Z(data_out[34]) );
  MUX2_X1 U312 ( .A(\mux[6][35] ), .B(\mux[7][35] ), .S(n260), .Z(n220) );
  MUX2_X1 U313 ( .A(\mux[4][35] ), .B(\mux[5][35] ), .S(n260), .Z(n221) );
  MUX2_X1 U314 ( .A(n221), .B(n220), .S(n255), .Z(n222) );
  MUX2_X1 U315 ( .A(\mux[2][35] ), .B(\mux[3][35] ), .S(n260), .Z(n223) );
  MUX2_X1 U316 ( .A(\mux[0][35] ), .B(\mux[1][35] ), .S(n260), .Z(n224) );
  MUX2_X1 U317 ( .A(n224), .B(n223), .S(n254), .Z(n225) );
  MUX2_X1 U318 ( .A(n225), .B(n222), .S(n251), .Z(data_out[35]) );
  MUX2_X1 U319 ( .A(\mux[6][36] ), .B(\mux[7][36] ), .S(n260), .Z(n226) );
  MUX2_X1 U320 ( .A(\mux[4][36] ), .B(\mux[5][36] ), .S(n260), .Z(n227) );
  MUX2_X1 U321 ( .A(n227), .B(n226), .S(n252), .Z(n228) );
  MUX2_X1 U322 ( .A(\mux[2][36] ), .B(\mux[3][36] ), .S(n260), .Z(n229) );
  MUX2_X1 U323 ( .A(\mux[0][36] ), .B(\mux[1][36] ), .S(n260), .Z(n230) );
  MUX2_X1 U324 ( .A(n230), .B(n229), .S(n253), .Z(n231) );
  MUX2_X1 U325 ( .A(n231), .B(n228), .S(addr_y[2]), .Z(data_out[36]) );
  MUX2_X1 U326 ( .A(\mux[6][37] ), .B(\mux[7][37] ), .S(n261), .Z(n232) );
  MUX2_X1 U327 ( .A(\mux[4][37] ), .B(\mux[5][37] ), .S(n261), .Z(n233) );
  MUX2_X1 U328 ( .A(n233), .B(n232), .S(n254), .Z(n234) );
  MUX2_X1 U329 ( .A(\mux[2][37] ), .B(\mux[3][37] ), .S(n261), .Z(n235) );
  MUX2_X1 U330 ( .A(\mux[0][37] ), .B(\mux[1][37] ), .S(n261), .Z(n236) );
  MUX2_X1 U331 ( .A(n236), .B(n235), .S(n255), .Z(n237) );
  MUX2_X1 U332 ( .A(n237), .B(n234), .S(n251), .Z(data_out[37]) );
  MUX2_X1 U333 ( .A(\mux[6][38] ), .B(\mux[7][38] ), .S(n261), .Z(n238) );
  MUX2_X1 U334 ( .A(\mux[4][38] ), .B(\mux[5][38] ), .S(n261), .Z(n239) );
  MUX2_X1 U335 ( .A(n239), .B(n238), .S(n255), .Z(n240) );
  MUX2_X1 U336 ( .A(\mux[2][38] ), .B(\mux[3][38] ), .S(n261), .Z(n241) );
  MUX2_X1 U337 ( .A(\mux[0][38] ), .B(\mux[1][38] ), .S(n261), .Z(n242) );
  MUX2_X1 U338 ( .A(n242), .B(n241), .S(n252), .Z(n243) );
  MUX2_X1 U339 ( .A(n243), .B(n240), .S(n251), .Z(data_out[38]) );
  MUX2_X1 U340 ( .A(\mux[6][39] ), .B(\mux[7][39] ), .S(n261), .Z(n244) );
  MUX2_X1 U341 ( .A(\mux[4][39] ), .B(\mux[5][39] ), .S(n261), .Z(n245) );
  MUX2_X1 U342 ( .A(n245), .B(n244), .S(n253), .Z(n246) );
  MUX2_X1 U343 ( .A(\mux[2][39] ), .B(\mux[3][39] ), .S(n261), .Z(n247) );
  MUX2_X1 U344 ( .A(\mux[0][39] ), .B(\mux[1][39] ), .S(n261), .Z(n248) );
  MUX2_X1 U345 ( .A(n248), .B(n247), .S(n254), .Z(n249) );
  MUX2_X1 U346 ( .A(n249), .B(n246), .S(n251), .Z(data_out[39]) );
endmodule


module mvm_8_8_20_1 ( clk, reset, loadMatrix, loadVector, start, done, data_in, 
        data_out );
  input [19:0] data_in;
  output [39:0] data_out;
  input clk, reset, loadMatrix, loadVector, start;
  output done;
  wire   wr_en_x, clear_acc, wr_en_y, \addr_a[7][2] , \addr_a[7][1] ,
         \addr_a[7][0] , \addr_a[6][2] , \addr_a[6][1] , \addr_a[6][0] ,
         \addr_a[5][2] , \addr_a[5][1] , \addr_a[5][0] , \addr_a[4][2] ,
         \addr_a[4][1] , \addr_a[4][0] , \addr_a[3][2] , \addr_a[3][1] ,
         \addr_a[3][0] , \addr_a[2][2] , \addr_a[2][1] , \addr_a[2][0] ,
         \addr_a[1][2] , \addr_a[1][1] , \addr_a[1][0] , \addr_a[0][2] ,
         \addr_a[0][1] , \addr_a[0][0] ;
  wire   [3:0] addr_x;
  wire   [3:0] addr_y;
  wire   [7:0] wr_en_a;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9;

  controlpath c ( .clk(clk), .reset(reset), .start(start), .loadMatrix(
        loadMatrix), .loadVector(loadVector), .wr_en_x(wr_en_x), .clear_acc(
        clear_acc), .wr_en_y(wr_en_y), .done(done), .addr_x({
        SYNOPSYS_UNCONNECTED__0, addr_x[2:0]}), .addr_y({
        SYNOPSYS_UNCONNECTED__1, addr_y[2:0]}), .addr_a({
        SYNOPSYS_UNCONNECTED__2, \addr_a[7][2] , \addr_a[7][1] , 
        \addr_a[7][0] , SYNOPSYS_UNCONNECTED__3, \addr_a[6][2] , 
        \addr_a[6][1] , \addr_a[6][0] , SYNOPSYS_UNCONNECTED__4, 
        \addr_a[5][2] , \addr_a[5][1] , \addr_a[5][0] , 
        SYNOPSYS_UNCONNECTED__5, \addr_a[4][2] , \addr_a[4][1] , 
        \addr_a[4][0] , SYNOPSYS_UNCONNECTED__6, \addr_a[3][2] , 
        \addr_a[3][1] , \addr_a[3][0] , SYNOPSYS_UNCONNECTED__7, 
        \addr_a[2][2] , \addr_a[2][1] , \addr_a[2][0] , 
        SYNOPSYS_UNCONNECTED__8, \addr_a[1][2] , \addr_a[1][1] , 
        \addr_a[1][0] , SYNOPSYS_UNCONNECTED__9, \addr_a[0][2] , 
        \addr_a[0][1] , \addr_a[0][0] }), .wr_en_a(wr_en_a) );
  datapath d ( .clk(clk), .wr_en_x(wr_en_x), .clear_acc(clear_acc), .wr_en_y(
        wr_en_y), .addr_x({1'b0, addr_x[2:0]}), .addr_y({1'b0, addr_y[2:0]}), 
        .addr_a({1'b0, \addr_a[7][2] , \addr_a[7][1] , \addr_a[7][0] , 1'b0, 
        \addr_a[6][2] , \addr_a[6][1] , \addr_a[6][0] , 1'b0, \addr_a[5][2] , 
        \addr_a[5][1] , \addr_a[5][0] , 1'b0, \addr_a[4][2] , \addr_a[4][1] , 
        \addr_a[4][0] , 1'b0, \addr_a[3][2] , \addr_a[3][1] , \addr_a[3][0] , 
        1'b0, \addr_a[2][2] , \addr_a[2][1] , \addr_a[2][0] , 1'b0, 
        \addr_a[1][2] , \addr_a[1][1] , \addr_a[1][0] , 1'b0, \addr_a[0][2] , 
        \addr_a[0][1] , \addr_a[0][0] }), .data_in(data_in), .wr_en_a(wr_en_a), 
        .data_out(data_out) );
endmodule

