
module control_K32_logK6_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[11]), .B(A[11]), .Z(SUM[11]) );
endmodule


module control_K32_logK6_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(carry[6]), .B(A[6]), .Z(SUM[6]) );
endmodule


module control_K32_logK6_DW01_inc_2 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(carry[12]), .B(A[12]), .Z(SUM[12]) );
endmodule


module control_K32_logK6_DW01_inc_3 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[6]), .B(A[6]), .Z(SUM[6]) );
endmodule


module control_K32_logK6 ( clk, start, reset, loadMatrix, loadVector, addr_x, 
        wr_en_x, addr_a, wr_en_a, clear_acc, addr_y, wr_en_y, done );
  output [5:0] addr_x;
  output [11:0] addr_a;
  output [5:0] addr_y;
  input clk, start, reset, loadMatrix, loadVector;
  output wr_en_x, wr_en_a, clear_acc, wr_en_y, done;
  wire   N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N65, N66,
         N67, N68, N69, N70, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81,
         N82, N83, N84, N85, N86, N87, N89, N90, N91, N92, N93, N94, N95, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N173, N174, N175, N176, N177, N178, N217, N218, N219, N220, N221,
         N222, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N292, n3, n21, n22, n23, n24, n25, n26, n29, n33, n37, n38, n39, n40,
         n41, n42, n44, n46, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, N299, N298,
         N297, N296, N295, N294, N293, \add_162/carry[11] ,
         \add_162/carry[10] , \add_162/carry[9] , \add_162/carry[8] ,
         \add_162/carry[7] , \add_162/carry[6] , n1, n2, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n27, n28,
         n30, n31, n32, n34, n35, n36, n43, n45;
  wire   [2:0] state;
  wire   [12:0] counter;
  wire   [6:0] counter2;
  wire   [6:0] multiplier;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign addr_x[5] = 1'b0;

  DFF_X1 \counter_reg[6]  ( .D(N81), .CK(clk), .Q(counter[6]) );
  DFF_X1 \counter_reg[7]  ( .D(N82), .CK(clk), .Q(counter[7]) );
  DFF_X1 \counter_reg[8]  ( .D(N83), .CK(clk), .Q(counter[8]) );
  DFF_X1 \counter_reg[9]  ( .D(N84), .CK(clk), .Q(counter[9]) );
  DFF_X1 \counter_reg[10]  ( .D(N85), .CK(clk), .Q(counter[10]) );
  DFF_X1 \counter_reg[11]  ( .D(N86), .CK(clk), .Q(counter[11]) );
  DFF_X1 \counter_reg[12]  ( .D(N87), .CK(clk), .Q(counter[12]) );
  DFF_X1 \state_reg[0]  ( .D(N72), .CK(clk), .Q(state[0]) );
  DLH_X1 \addr_x_reg[4]  ( .G(N217), .D(N222), .Q(addr_x[4]) );
  DLH_X1 \addr_x_reg[3]  ( .G(N217), .D(N221), .Q(addr_x[3]) );
  DLH_X1 \addr_x_reg[2]  ( .G(N217), .D(N220), .Q(addr_x[2]) );
  DLH_X1 \addr_x_reg[1]  ( .G(N217), .D(N219), .Q(addr_x[1]) );
  DLH_X1 \addr_x_reg[0]  ( .G(N217), .D(N218), .Q(addr_x[0]) );
  DLH_X1 \addr_a_reg[0]  ( .G(N217), .D(N224), .Q(addr_a[0]) );
  DLH_X1 \addr_a_reg[1]  ( .G(N217), .D(N225), .Q(addr_a[1]) );
  DLH_X1 \addr_a_reg[2]  ( .G(N217), .D(N226), .Q(addr_a[2]) );
  DLH_X1 \addr_a_reg[3]  ( .G(N217), .D(N227), .Q(addr_a[3]) );
  DLH_X1 \addr_a_reg[4]  ( .G(N217), .D(N228), .Q(addr_a[4]) );
  DLH_X1 \addr_a_reg[5]  ( .G(N217), .D(N229), .Q(addr_a[5]) );
  DLH_X1 \addr_a_reg[6]  ( .G(N217), .D(N230), .Q(addr_a[6]) );
  DLH_X1 \addr_a_reg[7]  ( .G(N217), .D(N231), .Q(addr_a[7]) );
  DLH_X1 \addr_a_reg[8]  ( .G(N217), .D(N232), .Q(addr_a[8]) );
  DLH_X1 \addr_a_reg[9]  ( .G(N217), .D(N233), .Q(addr_a[9]) );
  DLH_X1 \addr_a_reg[10]  ( .G(N217), .D(n8), .Q(addr_a[10]) );
  DLH_X1 \addr_a_reg[11]  ( .G(N217), .D(n7), .Q(addr_a[11]) );
  OAI22_X2 U34 ( .A1(n34), .A2(n22), .B1(n70), .B2(n38), .ZN(addr_y[4]) );
  NOR2_X2 U108 ( .A1(n87), .A2(n34), .ZN(n91) );
  NAND3_X1 U146 ( .A1(n108), .A2(n17), .A3(n71), .ZN(N217) );
  NAND3_X1 U147 ( .A1(n33), .A2(n29), .A3(state[0]), .ZN(n79) );
  NAND3_X1 U149 ( .A1(n76), .A2(n87), .A3(n86), .ZN(n108) );
  control_K32_logK6_DW01_inc_0 add_154 ( .A(addr_a), .SUM({N164, N163, N162, 
        N161, N160, N159, N158, N157, N156, N155, N154, N153}) );
  control_K32_logK6_DW01_inc_1 add_85 ( .A(multiplier), .SUM({N70, N69, N68, 
        N67, N66, N65, SYNOPSYS_UNCONNECTED__0}) );
  control_K32_logK6_DW01_inc_2 add_82 ( .A(counter), .SUM({N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, SYNOPSYS_UNCONNECTED__1}) );
  control_K32_logK6_DW01_inc_3 add_88_aco ( .A({N299, N298, N297, N296, N295, 
        N294, N293}), .SUM({N95, N94, N93, N92, N91, N90, N89}) );
  FA_X1 \add_162/U1_6  ( .A(multiplier[1]), .B(counter2[6]), .CI(
        \add_162/carry[6] ), .CO(\add_162/carry[7] ), .S(N173) );
  DFF_X1 \counter_reg[0]  ( .D(N75), .CK(clk), .Q(counter[0]), .QN(n42) );
  DFF_X1 \counter_reg[1]  ( .D(N76), .CK(clk), .Q(counter[1]), .QN(n41) );
  DFF_X1 \counter_reg[2]  ( .D(N77), .CK(clk), .Q(counter[2]), .QN(n40) );
  DFF_X1 \counter_reg[3]  ( .D(N78), .CK(clk), .Q(counter[3]), .QN(n39) );
  DFF_X1 \counter_reg[4]  ( .D(N79), .CK(clk), .Q(counter[4]), .QN(n38) );
  DFF_X1 \counter2_reg[0]  ( .D(n119), .CK(clk), .Q(counter2[0]), .QN(n19) );
  DFF_X1 \counter_reg[5]  ( .D(N80), .CK(clk), .Q(counter[5]), .QN(n37) );
  DFF_X1 \counter2_reg[1]  ( .D(n120), .CK(clk), .Q(counter2[1]), .QN(n6) );
  DFF_X1 \multiplier_reg[5]  ( .D(n112), .CK(clk), .Q(multiplier[5]), .QN(n21)
         );
  DFF_X1 \multiplier_reg[4]  ( .D(n113), .CK(clk), .Q(multiplier[4]), .QN(n22)
         );
  DFF_X1 \multiplier_reg[3]  ( .D(n114), .CK(clk), .Q(multiplier[3]), .QN(n23)
         );
  DFF_X1 \multiplier_reg[2]  ( .D(n115), .CK(clk), .Q(multiplier[2]), .QN(n24)
         );
  DFF_X1 \multiplier_reg[1]  ( .D(n116), .CK(clk), .Q(multiplier[1]), .QN(n25)
         );
  DFF_X1 \multiplier_reg[0]  ( .D(n117), .CK(clk), .Q(multiplier[0]), .QN(n26)
         );
  DFF_X1 \multiplier_reg[6]  ( .D(n118), .CK(clk), .Q(multiplier[6]), .QN(n3)
         );
  DFF_X1 \state_reg[2]  ( .D(N74), .CK(clk), .Q(state[2]), .QN(n29) );
  DFF_X1 \counter2_reg[2]  ( .D(n121), .CK(clk), .Q(counter2[2]), .QN(n5) );
  DFF_X1 \state_reg[1]  ( .D(N73), .CK(clk), .Q(state[1]), .QN(n33) );
  DFF_X1 \counter2_reg[3]  ( .D(n122), .CK(clk), .Q(counter2[3]), .QN(n4) );
  DFF_X1 \counter2_reg[4]  ( .D(n123), .CK(clk), .Q(counter2[4]), .QN(n2) );
  DFF_X1 \counter2_reg[5]  ( .D(n124), .CK(clk), .Q(counter2[5]), .QN(n46) );
  DFF_X1 \counter2_reg[6]  ( .D(n125), .CK(clk), .Q(counter2[6]), .QN(n44) );
  OAI22_X1 U4 ( .A1(n34), .A2(n24), .B1(n70), .B2(n40), .ZN(addr_y[2]) );
  XNOR2_X1 U5 ( .A(counter2[5]), .B(multiplier[0]), .ZN(n1) );
  INV_X1 U6 ( .A(n90), .ZN(n15) );
  INV_X1 U7 ( .A(wr_en_a), .ZN(n12) );
  INV_X1 U8 ( .A(wr_en_x), .ZN(n10) );
  OAI21_X1 U9 ( .B1(n59), .B2(n36), .A(n60), .ZN(n56) );
  NOR2_X1 U10 ( .A1(n79), .A2(n13), .ZN(wr_en_a) );
  NAND2_X1 U11 ( .A1(n71), .A2(n18), .ZN(clear_acc) );
  INV_X1 U12 ( .A(wr_en_y), .ZN(n18) );
  NAND2_X1 U13 ( .A1(n58), .A2(n56), .ZN(n57) );
  INV_X1 U14 ( .A(n76), .ZN(n34) );
  NOR2_X1 U15 ( .A1(n34), .A2(n59), .ZN(wr_en_y) );
  NOR2_X1 U16 ( .A1(n81), .A2(n11), .ZN(wr_en_x) );
  INV_X1 U17 ( .A(n80), .ZN(n11) );
  AND2_X1 U18 ( .A1(n59), .A2(n58), .ZN(N292) );
  INV_X1 U19 ( .A(n73), .ZN(n9) );
  INV_X1 U20 ( .A(n78), .ZN(n13) );
  AND2_X1 U21 ( .A1(N62), .A2(n58), .ZN(N86) );
  AND2_X1 U22 ( .A1(N61), .A2(n58), .ZN(N85) );
  AND2_X1 U23 ( .A1(N60), .A2(n58), .ZN(N84) );
  AND2_X1 U24 ( .A1(N59), .A2(n58), .ZN(N83) );
  AND2_X1 U25 ( .A1(N58), .A2(n58), .ZN(N82) );
  AND2_X1 U26 ( .A1(N57), .A2(n58), .ZN(N81) );
  INV_X1 U27 ( .A(n87), .ZN(n16) );
  AND2_X1 U28 ( .A1(N56), .A2(n58), .ZN(N80) );
  AND2_X1 U29 ( .A1(N55), .A2(n58), .ZN(N79) );
  AND2_X1 U30 ( .A1(N54), .A2(n58), .ZN(N78) );
  AND2_X1 U31 ( .A1(N53), .A2(n58), .ZN(N77) );
  AND2_X1 U32 ( .A1(N52), .A2(n58), .ZN(N76) );
  INV_X1 U33 ( .A(n91), .ZN(n17) );
  NOR2_X1 U35 ( .A1(n109), .A2(n108), .ZN(n90) );
  NOR2_X1 U36 ( .A1(n108), .A2(n14), .ZN(n92) );
  INV_X1 U37 ( .A(n109), .ZN(n14) );
  NAND2_X1 U38 ( .A1(n60), .A2(n36), .ZN(n61) );
  INV_X1 U39 ( .A(n58), .ZN(n36) );
  NOR4_X1 U40 ( .A1(counter[5]), .A2(counter[6]), .A3(n13), .A4(n110), .ZN(n80) );
  OR3_X1 U41 ( .A1(counter[7]), .A2(counter[9]), .A3(counter[8]), .ZN(n110) );
  OAI221_X1 U42 ( .B1(n78), .B2(n79), .C1(n80), .C2(n81), .A(n82), .ZN(n73) );
  AOI21_X1 U43 ( .B1(n83), .B2(n84), .A(n85), .ZN(n82) );
  NOR3_X1 U44 ( .A1(n42), .A2(n40), .A3(n41), .ZN(n83) );
  NOR3_X1 U45 ( .A1(n34), .A2(n16), .A3(n86), .ZN(n85) );
  NAND3_X1 U46 ( .A1(state[1]), .A2(n29), .A3(state[0]), .ZN(n70) );
  NOR4_X1 U47 ( .A1(n11), .A2(n70), .A3(n38), .A4(n39), .ZN(n84) );
  NOR3_X1 U48 ( .A1(counter[12]), .A2(counter[11]), .A3(counter[10]), .ZN(n78)
         );
  OAI221_X1 U49 ( .B1(n70), .B2(n41), .C1(n34), .C2(n25), .A(n29), .ZN(
        addr_y[1]) );
  OAI221_X1 U50 ( .B1(n70), .B2(n42), .C1(n34), .C2(n26), .A(n29), .ZN(
        addr_y[0]) );
  NOR2_X1 U51 ( .A1(n74), .A2(state[2]), .ZN(n76) );
  OAI22_X1 U52 ( .A1(n56), .A2(n21), .B1(n57), .B2(n27), .ZN(n112) );
  INV_X1 U53 ( .A(N69), .ZN(n27) );
  OAI22_X1 U54 ( .A1(n56), .A2(n22), .B1(n57), .B2(n28), .ZN(n113) );
  INV_X1 U55 ( .A(N68), .ZN(n28) );
  OAI22_X1 U56 ( .A1(n56), .A2(n23), .B1(n57), .B2(n30), .ZN(n114) );
  INV_X1 U57 ( .A(N67), .ZN(n30) );
  OAI22_X1 U58 ( .A1(n56), .A2(n24), .B1(n57), .B2(n31), .ZN(n115) );
  INV_X1 U59 ( .A(N66), .ZN(n31) );
  OAI22_X1 U60 ( .A1(n56), .A2(n25), .B1(n57), .B2(n32), .ZN(n116) );
  INV_X1 U61 ( .A(N65), .ZN(n32) );
  OAI22_X1 U62 ( .A1(n56), .A2(n26), .B1(n57), .B2(multiplier[0]), .ZN(n117)
         );
  OAI22_X1 U63 ( .A1(n56), .A2(n3), .B1(n57), .B2(n20), .ZN(n118) );
  INV_X1 U64 ( .A(N70), .ZN(n20) );
  OAI22_X1 U65 ( .A1(n34), .A2(n21), .B1(n70), .B2(n37), .ZN(addr_y[5]) );
  OAI22_X1 U66 ( .A1(reset), .A2(n43), .B1(n77), .B2(n36), .ZN(N72) );
  AOI22_X1 U67 ( .A1(n9), .A2(state[0]), .B1(n76), .B2(n73), .ZN(n77) );
  NAND2_X1 U68 ( .A1(n88), .A2(n19), .ZN(n87) );
  OAI22_X1 U69 ( .A1(n34), .A2(n23), .B1(n70), .B2(n39), .ZN(addr_y[3]) );
  OAI21_X1 U70 ( .B1(n75), .B2(n36), .A(n60), .ZN(N73) );
  AOI21_X1 U71 ( .B1(n9), .B2(state[1]), .A(n76), .ZN(n75) );
  OAI21_X1 U72 ( .B1(n72), .B2(n36), .A(n35), .ZN(N74) );
  AOI21_X1 U73 ( .B1(n73), .B2(n74), .A(state[2]), .ZN(n72) );
  OAI21_X1 U74 ( .B1(n61), .B2(n6), .A(n63), .ZN(n120) );
  NAND2_X1 U75 ( .A1(N90), .A2(n61), .ZN(n63) );
  OAI21_X1 U76 ( .B1(n61), .B2(n5), .A(n64), .ZN(n121) );
  NAND2_X1 U77 ( .A1(N91), .A2(n61), .ZN(n64) );
  OAI21_X1 U78 ( .B1(n61), .B2(n4), .A(n65), .ZN(n122) );
  NAND2_X1 U79 ( .A1(N92), .A2(n61), .ZN(n65) );
  OAI21_X1 U80 ( .B1(n61), .B2(n2), .A(n66), .ZN(n123) );
  NAND2_X1 U81 ( .A1(N93), .A2(n61), .ZN(n66) );
  OAI21_X1 U82 ( .B1(n61), .B2(n44), .A(n68), .ZN(n125) );
  NAND2_X1 U83 ( .A1(N95), .A2(n61), .ZN(n68) );
  NAND2_X1 U84 ( .A1(counter2[0]), .A2(n88), .ZN(n59) );
  OAI21_X1 U85 ( .B1(n46), .B2(n61), .A(n67), .ZN(n124) );
  NAND2_X1 U86 ( .A1(N94), .A2(n61), .ZN(n67) );
  OR3_X1 U87 ( .A1(state[1]), .A2(state[2]), .A3(state[0]), .ZN(n81) );
  OAI21_X1 U88 ( .B1(n19), .B2(n61), .A(n62), .ZN(n119) );
  NAND2_X1 U89 ( .A1(N89), .A2(n61), .ZN(n62) );
  OR2_X1 U90 ( .A1(n33), .A2(state[0]), .ZN(n74) );
  AND4_X1 U91 ( .A1(n6), .A2(n5), .A3(counter2[5]), .A4(n111), .ZN(n88) );
  NOR3_X1 U92 ( .A1(counter2[3]), .A2(counter2[6]), .A3(counter2[4]), .ZN(n111) );
  AND2_X1 U93 ( .A1(N63), .A2(n58), .ZN(N87) );
  NOR2_X1 U94 ( .A1(multiplier[6]), .A2(multiplier[5]), .ZN(n86) );
  OAI21_X1 U95 ( .B1(n36), .B2(counter[0]), .A(n60), .ZN(N75) );
  AND4_X1 U96 ( .A1(n70), .A2(n79), .A3(n81), .A4(n29), .ZN(n71) );
  NAND4_X1 U97 ( .A1(start), .A2(n43), .A3(n45), .A4(n35), .ZN(n60) );
  INV_X1 U98 ( .A(loadVector), .ZN(n45) );
  OAI221_X1 U99 ( .B1(n15), .B2(n1), .C1(n37), .C2(n12), .A(n102), .ZN(N229)
         );
  AOI22_X1 U100 ( .A1(N158), .A2(n91), .B1(addr_a[5]), .B2(n92), .ZN(n102) );
  OAI221_X1 U101 ( .B1(n15), .B2(n2), .C1(n38), .C2(n12), .A(n103), .ZN(N228)
         );
  AOI22_X1 U102 ( .A1(N157), .A2(n91), .B1(addr_a[4]), .B2(n92), .ZN(n103) );
  OAI221_X1 U103 ( .B1(n15), .B2(n4), .C1(n39), .C2(n12), .A(n104), .ZN(N227)
         );
  AOI22_X1 U104 ( .A1(N156), .A2(n91), .B1(addr_a[3]), .B2(n92), .ZN(n104) );
  OAI221_X1 U105 ( .B1(n15), .B2(n5), .C1(n40), .C2(n12), .A(n105), .ZN(N226)
         );
  AOI22_X1 U106 ( .A1(N155), .A2(n91), .B1(addr_a[2]), .B2(n92), .ZN(n105) );
  OAI221_X1 U107 ( .B1(n15), .B2(n6), .C1(n41), .C2(n12), .A(n106), .ZN(N225)
         );
  AOI22_X1 U109 ( .A1(N154), .A2(n91), .B1(addr_a[1]), .B2(n92), .ZN(n106) );
  OAI221_X1 U110 ( .B1(n15), .B2(n19), .C1(n42), .C2(n12), .A(n107), .ZN(N224)
         );
  AOI22_X1 U111 ( .A1(N153), .A2(n91), .B1(addr_a[0]), .B2(n92), .ZN(n107) );
  NOR4_X1 U112 ( .A1(n69), .A2(n70), .A3(counter[0]), .A4(n11), .ZN(done) );
  NAND4_X1 U113 ( .A1(n41), .A2(n40), .A3(n39), .A4(n38), .ZN(n69) );
  OAI22_X1 U114 ( .A1(n42), .A2(n10), .B1(n19), .B2(n15), .ZN(N218) );
  OAI22_X1 U115 ( .A1(n41), .A2(n10), .B1(n6), .B2(n15), .ZN(N219) );
  OAI22_X1 U116 ( .A1(n40), .A2(n10), .B1(n5), .B2(n15), .ZN(N220) );
  OAI22_X1 U117 ( .A1(n39), .A2(n10), .B1(n4), .B2(n15), .ZN(N221) );
  OAI22_X1 U118 ( .A1(n38), .A2(n10), .B1(n2), .B2(n15), .ZN(N222) );
  NAND2_X1 U119 ( .A1(n44), .A2(n46), .ZN(n109) );
  NAND2_X1 U120 ( .A1(n96), .A2(n97), .ZN(N232) );
  AOI22_X1 U121 ( .A1(N175), .A2(n90), .B1(counter[8]), .B2(wr_en_a), .ZN(n96)
         );
  AOI22_X1 U122 ( .A1(N161), .A2(n91), .B1(addr_a[8]), .B2(n92), .ZN(n97) );
  INV_X1 U123 ( .A(reset), .ZN(n35) );
  NAND2_X1 U124 ( .A1(n94), .A2(n95), .ZN(N233) );
  AOI22_X1 U125 ( .A1(N176), .A2(n90), .B1(counter[9]), .B2(wr_en_a), .ZN(n94)
         );
  AOI22_X1 U126 ( .A1(N162), .A2(n91), .B1(addr_a[9]), .B2(n92), .ZN(n95) );
  INV_X1 U127 ( .A(loadMatrix), .ZN(n43) );
  NAND2_X1 U128 ( .A1(n98), .A2(n99), .ZN(N231) );
  AOI22_X1 U129 ( .A1(N174), .A2(n90), .B1(counter[7]), .B2(wr_en_a), .ZN(n98)
         );
  AOI22_X1 U130 ( .A1(N160), .A2(n91), .B1(addr_a[7]), .B2(n92), .ZN(n99) );
  NAND2_X1 U131 ( .A1(n100), .A2(n101), .ZN(N230) );
  AOI22_X1 U132 ( .A1(N173), .A2(n90), .B1(counter[6]), .B2(wr_en_a), .ZN(n100) );
  AOI22_X1 U133 ( .A1(N159), .A2(n91), .B1(addr_a[6]), .B2(n92), .ZN(n101) );
  INV_X1 U134 ( .A(n89), .ZN(n7) );
  AOI222_X1 U135 ( .A1(N178), .A2(n90), .B1(N164), .B2(n91), .C1(addr_a[11]), 
        .C2(n92), .ZN(n89) );
  INV_X1 U136 ( .A(n93), .ZN(n8) );
  AOI222_X1 U137 ( .A1(N177), .A2(n90), .B1(N163), .B2(n91), .C1(addr_a[10]), 
        .C2(n92), .ZN(n93) );
  NOR4_X4 U138 ( .A1(loadMatrix), .A2(loadVector), .A3(reset), .A4(start), 
        .ZN(n58) );
  XOR2_X1 U139 ( .A(multiplier[6]), .B(\add_162/carry[11] ), .Z(N178) );
  AND2_X1 U140 ( .A1(\add_162/carry[10] ), .A2(multiplier[5]), .ZN(
        \add_162/carry[11] ) );
  XOR2_X1 U141 ( .A(multiplier[5]), .B(\add_162/carry[10] ), .Z(N177) );
  AND2_X1 U142 ( .A1(\add_162/carry[9] ), .A2(multiplier[4]), .ZN(
        \add_162/carry[10] ) );
  XOR2_X1 U143 ( .A(multiplier[4]), .B(\add_162/carry[9] ), .Z(N176) );
  AND2_X1 U144 ( .A1(\add_162/carry[8] ), .A2(multiplier[3]), .ZN(
        \add_162/carry[9] ) );
  XOR2_X1 U145 ( .A(multiplier[3]), .B(\add_162/carry[8] ), .Z(N175) );
  AND2_X1 U148 ( .A1(\add_162/carry[7] ), .A2(multiplier[2]), .ZN(
        \add_162/carry[8] ) );
  XOR2_X1 U150 ( .A(multiplier[2]), .B(\add_162/carry[7] ), .Z(N174) );
  AND2_X1 U151 ( .A1(multiplier[0]), .A2(counter2[5]), .ZN(\add_162/carry[6] )
         );
  AND2_X1 U152 ( .A1(counter2[0]), .A2(N292), .ZN(N293) );
  AND2_X1 U153 ( .A1(counter2[1]), .A2(N292), .ZN(N294) );
  AND2_X1 U154 ( .A1(counter2[2]), .A2(N292), .ZN(N295) );
  AND2_X1 U155 ( .A1(counter2[3]), .A2(N292), .ZN(N296) );
  AND2_X1 U156 ( .A1(counter2[4]), .A2(N292), .ZN(N297) );
  AND2_X1 U157 ( .A1(counter2[5]), .A2(N292), .ZN(N298) );
  AND2_X1 U158 ( .A1(N292), .A2(counter2[6]), .ZN(N299) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE6 ( clk, data_in, data_out, addr, wr_en );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N16, N17, N18, N19, N20, N22,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n625), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n626), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n627), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n628), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n629), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n630), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n631), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n632), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n633), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n634), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n635), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n636), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n637), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n638), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n639), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n640), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n641), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n642), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n643), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n644), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n645), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n646), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n647), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n648), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n649), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n650), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n651), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n652), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n653), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n654), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n655), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n656), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n657), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n658), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n659), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n660), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n661), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n662), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n663), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n664), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n665), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n666), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n667), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n668), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n669), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n670), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n671), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n672), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n673), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n674), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n675), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n676), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n677), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n678), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n679), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n680), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n681), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n682), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n683), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n684), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n685), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n686), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n687), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n688), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n689), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n690), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n691), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n692), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n693), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n694), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n695), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n696), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n697), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n698), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n699), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n700), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n701), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n702), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n703), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n704), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n705), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n706), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n707), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n708), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n709), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n710), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n711), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n712), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n713), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n714), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n715), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n716), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n717), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n718), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n719), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n720), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n721), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n722), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n723), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n724), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n725), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n726), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n727), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n728), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n729), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n730), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n731), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n732), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n733), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n734), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n735), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n736), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n737), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n738), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n739), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n740), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n741), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n742), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n743), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n744), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n745), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n746), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n747), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n748), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n749), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n750), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n751), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n752), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n753), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n754), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n755), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n756), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n757), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n758), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n759), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n760), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n761), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n762), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n763), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n764), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n765), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n766), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n767), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n768), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n769), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n770), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n771), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n772), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n773), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n774), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n775), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n776), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n777), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n778), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n779), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n780), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n781), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n782), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n783), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n784), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n785), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n786), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n787), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n788), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n789), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n790), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n791), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n792), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n793), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n794), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n795), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n796), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n797), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n798), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n799), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n800), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n801), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n802), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n803), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n804), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n805), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n806), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n807), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n808), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n809), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n810), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n811), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n812), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n813), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n814), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n815), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n816), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n594), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n593), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n592), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n591), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n590), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n589), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n588), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n587), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n586), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n585), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n584), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n583), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n582), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n581), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n580), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n579), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n578), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n577), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n576), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n575), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n574), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n573), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n572), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n571), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n570), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n569), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n568), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n567), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n566), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n565), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n564), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n563), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n562), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n561), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n560), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n559), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n558), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n557), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n556), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n555), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n554), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n553), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n552), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n551), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n550), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n549), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n548), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n547), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n546), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n545), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n544), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n543), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n542), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n541), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n540), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n539), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n538), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n537), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n536), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n535), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n534), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n533), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n532), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n531), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n61), .SI(n46), .SE(N14), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n606), .SI(n226), .SE(N14), .CK(clk), .Q(
        data_out[7]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  CLKBUF_X1 U3 ( .A(N11), .Z(n609) );
  BUF_X1 U4 ( .A(n614), .Z(n613) );
  BUF_X1 U5 ( .A(N10), .Z(n612) );
  BUF_X1 U6 ( .A(n614), .Z(n611) );
  INV_X1 U7 ( .A(n313), .ZN(n840) );
  INV_X1 U8 ( .A(n323), .ZN(n839) );
  INV_X1 U9 ( .A(n332), .ZN(n838) );
  INV_X1 U10 ( .A(n341), .ZN(n837) );
  INV_X1 U11 ( .A(n386), .ZN(n832) );
  INV_X1 U12 ( .A(n396), .ZN(n831) );
  INV_X1 U13 ( .A(n405), .ZN(n830) );
  INV_X1 U14 ( .A(n414), .ZN(n829) );
  INV_X1 U15 ( .A(n459), .ZN(n824) );
  INV_X1 U16 ( .A(n469), .ZN(n823) );
  INV_X1 U17 ( .A(n478), .ZN(n822) );
  INV_X1 U18 ( .A(n487), .ZN(n821) );
  INV_X1 U19 ( .A(n350), .ZN(n836) );
  INV_X1 U20 ( .A(n359), .ZN(n835) );
  INV_X1 U21 ( .A(n368), .ZN(n834) );
  INV_X1 U22 ( .A(n377), .ZN(n833) );
  INV_X1 U23 ( .A(n496), .ZN(n820) );
  INV_X1 U24 ( .A(n505), .ZN(n819) );
  INV_X1 U25 ( .A(n514), .ZN(n818) );
  INV_X1 U26 ( .A(n523), .ZN(n817) );
  INV_X1 U27 ( .A(n423), .ZN(n828) );
  INV_X1 U28 ( .A(n432), .ZN(n827) );
  INV_X1 U29 ( .A(n441), .ZN(n826) );
  INV_X1 U30 ( .A(n450), .ZN(n825) );
  BUF_X1 U31 ( .A(N11), .Z(n608) );
  BUF_X1 U32 ( .A(N10), .Z(n614) );
  NAND2_X1 U33 ( .A1(n250), .A2(n240), .ZN(n241) );
  NAND2_X1 U34 ( .A1(n260), .A2(n240), .ZN(n251) );
  NAND2_X1 U35 ( .A1(n270), .A2(n240), .ZN(n261) );
  NAND2_X1 U36 ( .A1(n280), .A2(n240), .ZN(n271) );
  NAND2_X1 U37 ( .A1(n290), .A2(n240), .ZN(n281) );
  NAND2_X1 U38 ( .A1(n300), .A2(n240), .ZN(n291) );
  NAND2_X1 U39 ( .A1(n310), .A2(n240), .ZN(n301) );
  NAND2_X1 U40 ( .A1(n239), .A2(n240), .ZN(n230) );
  NAND2_X1 U41 ( .A1(n321), .A2(n239), .ZN(n313) );
  NAND2_X1 U42 ( .A1(n321), .A2(n250), .ZN(n323) );
  NAND2_X1 U43 ( .A1(n321), .A2(n260), .ZN(n332) );
  NAND2_X1 U44 ( .A1(n321), .A2(n270), .ZN(n341) );
  NAND2_X1 U45 ( .A1(n394), .A2(n239), .ZN(n386) );
  NAND2_X1 U46 ( .A1(n394), .A2(n250), .ZN(n396) );
  NAND2_X1 U47 ( .A1(n394), .A2(n260), .ZN(n405) );
  NAND2_X1 U48 ( .A1(n394), .A2(n270), .ZN(n414) );
  NAND2_X1 U49 ( .A1(n467), .A2(n239), .ZN(n459) );
  NAND2_X1 U50 ( .A1(n467), .A2(n250), .ZN(n469) );
  NAND2_X1 U51 ( .A1(n467), .A2(n260), .ZN(n478) );
  NAND2_X1 U52 ( .A1(n467), .A2(n270), .ZN(n487) );
  NAND2_X1 U53 ( .A1(n321), .A2(n280), .ZN(n350) );
  NAND2_X1 U54 ( .A1(n321), .A2(n290), .ZN(n359) );
  NAND2_X1 U55 ( .A1(n321), .A2(n300), .ZN(n368) );
  NAND2_X1 U56 ( .A1(n321), .A2(n310), .ZN(n377) );
  NAND2_X1 U57 ( .A1(n394), .A2(n280), .ZN(n423) );
  NAND2_X1 U58 ( .A1(n394), .A2(n290), .ZN(n432) );
  NAND2_X1 U59 ( .A1(n394), .A2(n300), .ZN(n441) );
  NAND2_X1 U60 ( .A1(n394), .A2(n310), .ZN(n450) );
  NAND2_X1 U61 ( .A1(n467), .A2(n280), .ZN(n496) );
  NAND2_X1 U62 ( .A1(n467), .A2(n290), .ZN(n505) );
  NAND2_X1 U63 ( .A1(n467), .A2(n300), .ZN(n514) );
  NAND2_X1 U64 ( .A1(n467), .A2(n310), .ZN(n523) );
  AND3_X1 U65 ( .A1(n843), .A2(n842), .A3(n311), .ZN(n240) );
  AND3_X1 U66 ( .A1(N13), .A2(n311), .A3(N14), .ZN(n467) );
  AND3_X1 U67 ( .A1(n311), .A2(n842), .A3(N13), .ZN(n321) );
  AND3_X1 U68 ( .A1(n311), .A2(n843), .A3(N14), .ZN(n394) );
  NOR2_X1 U69 ( .A1(n841), .A2(addr[5]), .ZN(n311) );
  INV_X1 U70 ( .A(wr_en), .ZN(n841) );
  OAI21_X1 U71 ( .B1(n230), .B2(n617), .A(n231), .ZN(n531) );
  NAND2_X1 U72 ( .A1(\mem[0][0] ), .A2(n230), .ZN(n231) );
  OAI21_X1 U73 ( .B1(n230), .B2(n618), .A(n232), .ZN(n532) );
  NAND2_X1 U74 ( .A1(\mem[0][1] ), .A2(n230), .ZN(n232) );
  OAI21_X1 U75 ( .B1(n230), .B2(n619), .A(n233), .ZN(n533) );
  NAND2_X1 U76 ( .A1(\mem[0][2] ), .A2(n230), .ZN(n233) );
  OAI21_X1 U77 ( .B1(n230), .B2(n620), .A(n234), .ZN(n534) );
  NAND2_X1 U78 ( .A1(\mem[0][3] ), .A2(n230), .ZN(n234) );
  OAI21_X1 U79 ( .B1(n230), .B2(n621), .A(n235), .ZN(n535) );
  NAND2_X1 U80 ( .A1(\mem[0][4] ), .A2(n230), .ZN(n235) );
  OAI21_X1 U81 ( .B1(n230), .B2(n622), .A(n236), .ZN(n536) );
  NAND2_X1 U82 ( .A1(\mem[0][5] ), .A2(n230), .ZN(n236) );
  OAI21_X1 U83 ( .B1(n230), .B2(n623), .A(n237), .ZN(n537) );
  NAND2_X1 U84 ( .A1(\mem[0][6] ), .A2(n230), .ZN(n237) );
  OAI21_X1 U85 ( .B1(n230), .B2(n624), .A(n238), .ZN(n538) );
  NAND2_X1 U86 ( .A1(\mem[0][7] ), .A2(n230), .ZN(n238) );
  OAI21_X1 U87 ( .B1(n617), .B2(n241), .A(n242), .ZN(n539) );
  NAND2_X1 U88 ( .A1(\mem[1][0] ), .A2(n241), .ZN(n242) );
  OAI21_X1 U89 ( .B1(n618), .B2(n241), .A(n243), .ZN(n540) );
  NAND2_X1 U90 ( .A1(\mem[1][1] ), .A2(n241), .ZN(n243) );
  OAI21_X1 U91 ( .B1(n619), .B2(n241), .A(n244), .ZN(n541) );
  NAND2_X1 U92 ( .A1(\mem[1][2] ), .A2(n241), .ZN(n244) );
  OAI21_X1 U93 ( .B1(n620), .B2(n241), .A(n245), .ZN(n542) );
  NAND2_X1 U94 ( .A1(\mem[1][3] ), .A2(n241), .ZN(n245) );
  OAI21_X1 U95 ( .B1(n621), .B2(n241), .A(n246), .ZN(n543) );
  NAND2_X1 U96 ( .A1(\mem[1][4] ), .A2(n241), .ZN(n246) );
  OAI21_X1 U97 ( .B1(n622), .B2(n241), .A(n247), .ZN(n544) );
  NAND2_X1 U98 ( .A1(\mem[1][5] ), .A2(n241), .ZN(n247) );
  OAI21_X1 U99 ( .B1(n623), .B2(n241), .A(n248), .ZN(n545) );
  NAND2_X1 U100 ( .A1(\mem[1][6] ), .A2(n241), .ZN(n248) );
  OAI21_X1 U101 ( .B1(n624), .B2(n241), .A(n249), .ZN(n546) );
  NAND2_X1 U102 ( .A1(\mem[1][7] ), .A2(n241), .ZN(n249) );
  OAI21_X1 U103 ( .B1(n617), .B2(n251), .A(n252), .ZN(n547) );
  NAND2_X1 U104 ( .A1(\mem[2][0] ), .A2(n251), .ZN(n252) );
  OAI21_X1 U105 ( .B1(n618), .B2(n251), .A(n253), .ZN(n548) );
  NAND2_X1 U106 ( .A1(\mem[2][1] ), .A2(n251), .ZN(n253) );
  OAI21_X1 U107 ( .B1(n619), .B2(n251), .A(n254), .ZN(n549) );
  NAND2_X1 U108 ( .A1(\mem[2][2] ), .A2(n251), .ZN(n254) );
  OAI21_X1 U109 ( .B1(n620), .B2(n251), .A(n255), .ZN(n550) );
  NAND2_X1 U110 ( .A1(\mem[2][3] ), .A2(n251), .ZN(n255) );
  OAI21_X1 U111 ( .B1(n621), .B2(n251), .A(n256), .ZN(n551) );
  NAND2_X1 U112 ( .A1(\mem[2][4] ), .A2(n251), .ZN(n256) );
  OAI21_X1 U113 ( .B1(n622), .B2(n251), .A(n257), .ZN(n552) );
  NAND2_X1 U114 ( .A1(\mem[2][5] ), .A2(n251), .ZN(n257) );
  OAI21_X1 U115 ( .B1(n623), .B2(n251), .A(n258), .ZN(n553) );
  NAND2_X1 U116 ( .A1(\mem[2][6] ), .A2(n251), .ZN(n258) );
  OAI21_X1 U117 ( .B1(n624), .B2(n251), .A(n259), .ZN(n554) );
  NAND2_X1 U118 ( .A1(\mem[2][7] ), .A2(n251), .ZN(n259) );
  OAI21_X1 U119 ( .B1(n617), .B2(n261), .A(n262), .ZN(n555) );
  NAND2_X1 U120 ( .A1(\mem[3][0] ), .A2(n261), .ZN(n262) );
  OAI21_X1 U121 ( .B1(n618), .B2(n261), .A(n263), .ZN(n556) );
  NAND2_X1 U122 ( .A1(\mem[3][1] ), .A2(n261), .ZN(n263) );
  OAI21_X1 U123 ( .B1(n619), .B2(n261), .A(n264), .ZN(n557) );
  NAND2_X1 U124 ( .A1(\mem[3][2] ), .A2(n261), .ZN(n264) );
  OAI21_X1 U125 ( .B1(n620), .B2(n261), .A(n265), .ZN(n558) );
  NAND2_X1 U126 ( .A1(\mem[3][3] ), .A2(n261), .ZN(n265) );
  OAI21_X1 U127 ( .B1(n621), .B2(n261), .A(n266), .ZN(n559) );
  NAND2_X1 U128 ( .A1(\mem[3][4] ), .A2(n261), .ZN(n266) );
  OAI21_X1 U129 ( .B1(n622), .B2(n261), .A(n267), .ZN(n560) );
  NAND2_X1 U130 ( .A1(\mem[3][5] ), .A2(n261), .ZN(n267) );
  OAI21_X1 U131 ( .B1(n623), .B2(n261), .A(n268), .ZN(n561) );
  NAND2_X1 U132 ( .A1(\mem[3][6] ), .A2(n261), .ZN(n268) );
  OAI21_X1 U133 ( .B1(n624), .B2(n261), .A(n269), .ZN(n562) );
  NAND2_X1 U134 ( .A1(\mem[3][7] ), .A2(n261), .ZN(n269) );
  OAI21_X1 U135 ( .B1(n617), .B2(n271), .A(n272), .ZN(n563) );
  NAND2_X1 U136 ( .A1(\mem[4][0] ), .A2(n271), .ZN(n272) );
  OAI21_X1 U137 ( .B1(n618), .B2(n271), .A(n273), .ZN(n564) );
  NAND2_X1 U138 ( .A1(\mem[4][1] ), .A2(n271), .ZN(n273) );
  OAI21_X1 U139 ( .B1(n619), .B2(n271), .A(n274), .ZN(n565) );
  NAND2_X1 U140 ( .A1(\mem[4][2] ), .A2(n271), .ZN(n274) );
  OAI21_X1 U141 ( .B1(n620), .B2(n271), .A(n275), .ZN(n566) );
  NAND2_X1 U142 ( .A1(\mem[4][3] ), .A2(n271), .ZN(n275) );
  OAI21_X1 U143 ( .B1(n621), .B2(n271), .A(n276), .ZN(n567) );
  NAND2_X1 U144 ( .A1(\mem[4][4] ), .A2(n271), .ZN(n276) );
  OAI21_X1 U145 ( .B1(n622), .B2(n271), .A(n277), .ZN(n568) );
  NAND2_X1 U146 ( .A1(\mem[4][5] ), .A2(n271), .ZN(n277) );
  OAI21_X1 U147 ( .B1(n623), .B2(n271), .A(n278), .ZN(n569) );
  NAND2_X1 U148 ( .A1(\mem[4][6] ), .A2(n271), .ZN(n278) );
  OAI21_X1 U149 ( .B1(n624), .B2(n271), .A(n279), .ZN(n570) );
  NAND2_X1 U150 ( .A1(\mem[4][7] ), .A2(n271), .ZN(n279) );
  OAI21_X1 U151 ( .B1(n617), .B2(n291), .A(n292), .ZN(n579) );
  NAND2_X1 U152 ( .A1(\mem[6][0] ), .A2(n291), .ZN(n292) );
  OAI21_X1 U153 ( .B1(n618), .B2(n291), .A(n293), .ZN(n580) );
  NAND2_X1 U154 ( .A1(\mem[6][1] ), .A2(n291), .ZN(n293) );
  OAI21_X1 U155 ( .B1(n619), .B2(n291), .A(n294), .ZN(n581) );
  NAND2_X1 U156 ( .A1(\mem[6][2] ), .A2(n291), .ZN(n294) );
  OAI21_X1 U157 ( .B1(n620), .B2(n291), .A(n295), .ZN(n582) );
  NAND2_X1 U158 ( .A1(\mem[6][3] ), .A2(n291), .ZN(n295) );
  OAI21_X1 U159 ( .B1(n621), .B2(n291), .A(n296), .ZN(n583) );
  NAND2_X1 U160 ( .A1(\mem[6][4] ), .A2(n291), .ZN(n296) );
  OAI21_X1 U161 ( .B1(n622), .B2(n291), .A(n297), .ZN(n584) );
  NAND2_X1 U162 ( .A1(\mem[6][5] ), .A2(n291), .ZN(n297) );
  OAI21_X1 U163 ( .B1(n623), .B2(n291), .A(n298), .ZN(n585) );
  NAND2_X1 U164 ( .A1(\mem[6][6] ), .A2(n291), .ZN(n298) );
  OAI21_X1 U165 ( .B1(n624), .B2(n291), .A(n299), .ZN(n586) );
  NAND2_X1 U166 ( .A1(\mem[6][7] ), .A2(n291), .ZN(n299) );
  OAI21_X1 U167 ( .B1(n617), .B2(n301), .A(n302), .ZN(n587) );
  NAND2_X1 U168 ( .A1(\mem[7][0] ), .A2(n301), .ZN(n302) );
  OAI21_X1 U169 ( .B1(n618), .B2(n301), .A(n303), .ZN(n588) );
  NAND2_X1 U170 ( .A1(\mem[7][1] ), .A2(n301), .ZN(n303) );
  OAI21_X1 U171 ( .B1(n619), .B2(n301), .A(n304), .ZN(n589) );
  NAND2_X1 U172 ( .A1(\mem[7][2] ), .A2(n301), .ZN(n304) );
  OAI21_X1 U173 ( .B1(n620), .B2(n301), .A(n305), .ZN(n590) );
  NAND2_X1 U174 ( .A1(\mem[7][3] ), .A2(n301), .ZN(n305) );
  OAI21_X1 U175 ( .B1(n621), .B2(n301), .A(n306), .ZN(n591) );
  NAND2_X1 U176 ( .A1(\mem[7][4] ), .A2(n301), .ZN(n306) );
  OAI21_X1 U177 ( .B1(n622), .B2(n301), .A(n307), .ZN(n592) );
  NAND2_X1 U178 ( .A1(\mem[7][5] ), .A2(n301), .ZN(n307) );
  OAI21_X1 U179 ( .B1(n623), .B2(n301), .A(n308), .ZN(n593) );
  NAND2_X1 U180 ( .A1(\mem[7][6] ), .A2(n301), .ZN(n308) );
  OAI21_X1 U181 ( .B1(n624), .B2(n301), .A(n309), .ZN(n594) );
  NAND2_X1 U182 ( .A1(\mem[7][7] ), .A2(n301), .ZN(n309) );
  OAI21_X1 U183 ( .B1(n617), .B2(n281), .A(n282), .ZN(n571) );
  NAND2_X1 U184 ( .A1(\mem[5][0] ), .A2(n281), .ZN(n282) );
  OAI21_X1 U185 ( .B1(n618), .B2(n281), .A(n283), .ZN(n572) );
  NAND2_X1 U186 ( .A1(\mem[5][1] ), .A2(n281), .ZN(n283) );
  OAI21_X1 U187 ( .B1(n619), .B2(n281), .A(n284), .ZN(n573) );
  NAND2_X1 U188 ( .A1(\mem[5][2] ), .A2(n281), .ZN(n284) );
  OAI21_X1 U189 ( .B1(n620), .B2(n281), .A(n285), .ZN(n574) );
  NAND2_X1 U190 ( .A1(\mem[5][3] ), .A2(n281), .ZN(n285) );
  OAI21_X1 U191 ( .B1(n621), .B2(n281), .A(n286), .ZN(n575) );
  NAND2_X1 U192 ( .A1(\mem[5][4] ), .A2(n281), .ZN(n286) );
  OAI21_X1 U193 ( .B1(n622), .B2(n281), .A(n287), .ZN(n576) );
  NAND2_X1 U194 ( .A1(\mem[5][5] ), .A2(n281), .ZN(n287) );
  OAI21_X1 U195 ( .B1(n623), .B2(n281), .A(n288), .ZN(n577) );
  NAND2_X1 U196 ( .A1(\mem[5][6] ), .A2(n281), .ZN(n288) );
  OAI21_X1 U197 ( .B1(n624), .B2(n281), .A(n289), .ZN(n578) );
  NAND2_X1 U198 ( .A1(\mem[5][7] ), .A2(n281), .ZN(n289) );
  INV_X1 U199 ( .A(n312), .ZN(n816) );
  AOI22_X1 U200 ( .A1(data_in[0]), .A2(n840), .B1(n313), .B2(\mem[8][0] ), 
        .ZN(n312) );
  INV_X1 U201 ( .A(n314), .ZN(n815) );
  AOI22_X1 U202 ( .A1(data_in[1]), .A2(n840), .B1(n313), .B2(\mem[8][1] ), 
        .ZN(n314) );
  INV_X1 U203 ( .A(n315), .ZN(n814) );
  AOI22_X1 U204 ( .A1(data_in[2]), .A2(n840), .B1(n313), .B2(\mem[8][2] ), 
        .ZN(n315) );
  INV_X1 U205 ( .A(n316), .ZN(n813) );
  AOI22_X1 U206 ( .A1(data_in[3]), .A2(n840), .B1(n313), .B2(\mem[8][3] ), 
        .ZN(n316) );
  INV_X1 U207 ( .A(n317), .ZN(n812) );
  AOI22_X1 U208 ( .A1(data_in[4]), .A2(n840), .B1(n313), .B2(\mem[8][4] ), 
        .ZN(n317) );
  INV_X1 U209 ( .A(n318), .ZN(n811) );
  AOI22_X1 U210 ( .A1(data_in[5]), .A2(n840), .B1(n313), .B2(\mem[8][5] ), 
        .ZN(n318) );
  INV_X1 U211 ( .A(n319), .ZN(n810) );
  AOI22_X1 U212 ( .A1(data_in[6]), .A2(n840), .B1(n313), .B2(\mem[8][6] ), 
        .ZN(n319) );
  INV_X1 U213 ( .A(n320), .ZN(n809) );
  AOI22_X1 U214 ( .A1(data_in[7]), .A2(n840), .B1(n313), .B2(\mem[8][7] ), 
        .ZN(n320) );
  INV_X1 U215 ( .A(n322), .ZN(n808) );
  AOI22_X1 U216 ( .A1(data_in[0]), .A2(n839), .B1(n323), .B2(\mem[9][0] ), 
        .ZN(n322) );
  INV_X1 U217 ( .A(n324), .ZN(n807) );
  AOI22_X1 U218 ( .A1(data_in[1]), .A2(n839), .B1(n323), .B2(\mem[9][1] ), 
        .ZN(n324) );
  INV_X1 U219 ( .A(n325), .ZN(n806) );
  AOI22_X1 U220 ( .A1(data_in[2]), .A2(n839), .B1(n323), .B2(\mem[9][2] ), 
        .ZN(n325) );
  INV_X1 U221 ( .A(n326), .ZN(n805) );
  AOI22_X1 U222 ( .A1(data_in[3]), .A2(n839), .B1(n323), .B2(\mem[9][3] ), 
        .ZN(n326) );
  INV_X1 U223 ( .A(n327), .ZN(n804) );
  AOI22_X1 U224 ( .A1(data_in[4]), .A2(n839), .B1(n323), .B2(\mem[9][4] ), 
        .ZN(n327) );
  INV_X1 U225 ( .A(n328), .ZN(n803) );
  AOI22_X1 U226 ( .A1(data_in[5]), .A2(n839), .B1(n323), .B2(\mem[9][5] ), 
        .ZN(n328) );
  INV_X1 U227 ( .A(n329), .ZN(n802) );
  AOI22_X1 U228 ( .A1(data_in[6]), .A2(n839), .B1(n323), .B2(\mem[9][6] ), 
        .ZN(n329) );
  INV_X1 U229 ( .A(n330), .ZN(n801) );
  AOI22_X1 U230 ( .A1(data_in[7]), .A2(n839), .B1(n323), .B2(\mem[9][7] ), 
        .ZN(n330) );
  INV_X1 U231 ( .A(n331), .ZN(n800) );
  AOI22_X1 U232 ( .A1(data_in[0]), .A2(n838), .B1(n332), .B2(\mem[10][0] ), 
        .ZN(n331) );
  INV_X1 U233 ( .A(n333), .ZN(n799) );
  AOI22_X1 U234 ( .A1(data_in[1]), .A2(n838), .B1(n332), .B2(\mem[10][1] ), 
        .ZN(n333) );
  INV_X1 U235 ( .A(n334), .ZN(n798) );
  AOI22_X1 U236 ( .A1(data_in[2]), .A2(n838), .B1(n332), .B2(\mem[10][2] ), 
        .ZN(n334) );
  INV_X1 U237 ( .A(n335), .ZN(n797) );
  AOI22_X1 U238 ( .A1(data_in[3]), .A2(n838), .B1(n332), .B2(\mem[10][3] ), 
        .ZN(n335) );
  INV_X1 U239 ( .A(n336), .ZN(n796) );
  AOI22_X1 U240 ( .A1(data_in[4]), .A2(n838), .B1(n332), .B2(\mem[10][4] ), 
        .ZN(n336) );
  INV_X1 U241 ( .A(n337), .ZN(n795) );
  AOI22_X1 U242 ( .A1(data_in[5]), .A2(n838), .B1(n332), .B2(\mem[10][5] ), 
        .ZN(n337) );
  INV_X1 U243 ( .A(n338), .ZN(n794) );
  AOI22_X1 U244 ( .A1(data_in[6]), .A2(n838), .B1(n332), .B2(\mem[10][6] ), 
        .ZN(n338) );
  INV_X1 U245 ( .A(n339), .ZN(n793) );
  AOI22_X1 U246 ( .A1(data_in[7]), .A2(n838), .B1(n332), .B2(\mem[10][7] ), 
        .ZN(n339) );
  INV_X1 U247 ( .A(n340), .ZN(n792) );
  AOI22_X1 U248 ( .A1(data_in[0]), .A2(n837), .B1(n341), .B2(\mem[11][0] ), 
        .ZN(n340) );
  INV_X1 U249 ( .A(n342), .ZN(n791) );
  AOI22_X1 U250 ( .A1(data_in[1]), .A2(n837), .B1(n341), .B2(\mem[11][1] ), 
        .ZN(n342) );
  INV_X1 U251 ( .A(n343), .ZN(n790) );
  AOI22_X1 U252 ( .A1(data_in[2]), .A2(n837), .B1(n341), .B2(\mem[11][2] ), 
        .ZN(n343) );
  INV_X1 U253 ( .A(n344), .ZN(n789) );
  AOI22_X1 U254 ( .A1(data_in[3]), .A2(n837), .B1(n341), .B2(\mem[11][3] ), 
        .ZN(n344) );
  INV_X1 U255 ( .A(n345), .ZN(n788) );
  AOI22_X1 U256 ( .A1(data_in[4]), .A2(n837), .B1(n341), .B2(\mem[11][4] ), 
        .ZN(n345) );
  INV_X1 U257 ( .A(n346), .ZN(n787) );
  AOI22_X1 U258 ( .A1(data_in[5]), .A2(n837), .B1(n341), .B2(\mem[11][5] ), 
        .ZN(n346) );
  INV_X1 U259 ( .A(n347), .ZN(n786) );
  AOI22_X1 U260 ( .A1(data_in[6]), .A2(n837), .B1(n341), .B2(\mem[11][6] ), 
        .ZN(n347) );
  INV_X1 U261 ( .A(n348), .ZN(n785) );
  AOI22_X1 U262 ( .A1(data_in[7]), .A2(n837), .B1(n341), .B2(\mem[11][7] ), 
        .ZN(n348) );
  INV_X1 U263 ( .A(n349), .ZN(n784) );
  AOI22_X1 U264 ( .A1(data_in[0]), .A2(n836), .B1(n350), .B2(\mem[12][0] ), 
        .ZN(n349) );
  INV_X1 U265 ( .A(n351), .ZN(n783) );
  AOI22_X1 U266 ( .A1(data_in[1]), .A2(n836), .B1(n350), .B2(\mem[12][1] ), 
        .ZN(n351) );
  INV_X1 U267 ( .A(n352), .ZN(n782) );
  AOI22_X1 U268 ( .A1(data_in[2]), .A2(n836), .B1(n350), .B2(\mem[12][2] ), 
        .ZN(n352) );
  INV_X1 U269 ( .A(n353), .ZN(n781) );
  AOI22_X1 U270 ( .A1(data_in[3]), .A2(n836), .B1(n350), .B2(\mem[12][3] ), 
        .ZN(n353) );
  INV_X1 U271 ( .A(n354), .ZN(n780) );
  AOI22_X1 U272 ( .A1(data_in[4]), .A2(n836), .B1(n350), .B2(\mem[12][4] ), 
        .ZN(n354) );
  INV_X1 U273 ( .A(n355), .ZN(n779) );
  AOI22_X1 U274 ( .A1(data_in[5]), .A2(n836), .B1(n350), .B2(\mem[12][5] ), 
        .ZN(n355) );
  INV_X1 U275 ( .A(n356), .ZN(n778) );
  AOI22_X1 U276 ( .A1(data_in[6]), .A2(n836), .B1(n350), .B2(\mem[12][6] ), 
        .ZN(n356) );
  INV_X1 U277 ( .A(n357), .ZN(n777) );
  AOI22_X1 U278 ( .A1(data_in[7]), .A2(n836), .B1(n350), .B2(\mem[12][7] ), 
        .ZN(n357) );
  INV_X1 U279 ( .A(n358), .ZN(n776) );
  AOI22_X1 U280 ( .A1(data_in[0]), .A2(n835), .B1(n359), .B2(\mem[13][0] ), 
        .ZN(n358) );
  INV_X1 U281 ( .A(n360), .ZN(n775) );
  AOI22_X1 U282 ( .A1(data_in[1]), .A2(n835), .B1(n359), .B2(\mem[13][1] ), 
        .ZN(n360) );
  INV_X1 U283 ( .A(n361), .ZN(n774) );
  AOI22_X1 U284 ( .A1(data_in[2]), .A2(n835), .B1(n359), .B2(\mem[13][2] ), 
        .ZN(n361) );
  INV_X1 U285 ( .A(n362), .ZN(n773) );
  AOI22_X1 U286 ( .A1(data_in[3]), .A2(n835), .B1(n359), .B2(\mem[13][3] ), 
        .ZN(n362) );
  INV_X1 U287 ( .A(n363), .ZN(n772) );
  AOI22_X1 U288 ( .A1(data_in[4]), .A2(n835), .B1(n359), .B2(\mem[13][4] ), 
        .ZN(n363) );
  INV_X1 U289 ( .A(n364), .ZN(n771) );
  AOI22_X1 U290 ( .A1(data_in[5]), .A2(n835), .B1(n359), .B2(\mem[13][5] ), 
        .ZN(n364) );
  INV_X1 U291 ( .A(n365), .ZN(n770) );
  AOI22_X1 U292 ( .A1(data_in[6]), .A2(n835), .B1(n359), .B2(\mem[13][6] ), 
        .ZN(n365) );
  INV_X1 U293 ( .A(n366), .ZN(n769) );
  AOI22_X1 U294 ( .A1(data_in[7]), .A2(n835), .B1(n359), .B2(\mem[13][7] ), 
        .ZN(n366) );
  INV_X1 U295 ( .A(n367), .ZN(n768) );
  AOI22_X1 U296 ( .A1(data_in[0]), .A2(n834), .B1(n368), .B2(\mem[14][0] ), 
        .ZN(n367) );
  INV_X1 U297 ( .A(n369), .ZN(n767) );
  AOI22_X1 U298 ( .A1(data_in[1]), .A2(n834), .B1(n368), .B2(\mem[14][1] ), 
        .ZN(n369) );
  INV_X1 U299 ( .A(n370), .ZN(n766) );
  AOI22_X1 U300 ( .A1(data_in[2]), .A2(n834), .B1(n368), .B2(\mem[14][2] ), 
        .ZN(n370) );
  INV_X1 U301 ( .A(n371), .ZN(n765) );
  AOI22_X1 U302 ( .A1(data_in[3]), .A2(n834), .B1(n368), .B2(\mem[14][3] ), 
        .ZN(n371) );
  INV_X1 U303 ( .A(n372), .ZN(n764) );
  AOI22_X1 U304 ( .A1(data_in[4]), .A2(n834), .B1(n368), .B2(\mem[14][4] ), 
        .ZN(n372) );
  INV_X1 U305 ( .A(n373), .ZN(n763) );
  AOI22_X1 U306 ( .A1(data_in[5]), .A2(n834), .B1(n368), .B2(\mem[14][5] ), 
        .ZN(n373) );
  INV_X1 U307 ( .A(n374), .ZN(n762) );
  AOI22_X1 U308 ( .A1(data_in[6]), .A2(n834), .B1(n368), .B2(\mem[14][6] ), 
        .ZN(n374) );
  INV_X1 U309 ( .A(n375), .ZN(n761) );
  AOI22_X1 U310 ( .A1(data_in[7]), .A2(n834), .B1(n368), .B2(\mem[14][7] ), 
        .ZN(n375) );
  INV_X1 U311 ( .A(n376), .ZN(n760) );
  AOI22_X1 U312 ( .A1(data_in[0]), .A2(n833), .B1(n377), .B2(\mem[15][0] ), 
        .ZN(n376) );
  INV_X1 U313 ( .A(n378), .ZN(n759) );
  AOI22_X1 U314 ( .A1(data_in[1]), .A2(n833), .B1(n377), .B2(\mem[15][1] ), 
        .ZN(n378) );
  INV_X1 U315 ( .A(n379), .ZN(n758) );
  AOI22_X1 U316 ( .A1(data_in[2]), .A2(n833), .B1(n377), .B2(\mem[15][2] ), 
        .ZN(n379) );
  INV_X1 U317 ( .A(n380), .ZN(n757) );
  AOI22_X1 U318 ( .A1(data_in[3]), .A2(n833), .B1(n377), .B2(\mem[15][3] ), 
        .ZN(n380) );
  INV_X1 U319 ( .A(n381), .ZN(n756) );
  AOI22_X1 U320 ( .A1(data_in[4]), .A2(n833), .B1(n377), .B2(\mem[15][4] ), 
        .ZN(n381) );
  INV_X1 U321 ( .A(n382), .ZN(n755) );
  AOI22_X1 U322 ( .A1(data_in[5]), .A2(n833), .B1(n377), .B2(\mem[15][5] ), 
        .ZN(n382) );
  INV_X1 U323 ( .A(n383), .ZN(n754) );
  AOI22_X1 U324 ( .A1(data_in[6]), .A2(n833), .B1(n377), .B2(\mem[15][6] ), 
        .ZN(n383) );
  INV_X1 U325 ( .A(n384), .ZN(n753) );
  AOI22_X1 U326 ( .A1(data_in[7]), .A2(n833), .B1(n377), .B2(\mem[15][7] ), 
        .ZN(n384) );
  INV_X1 U327 ( .A(n385), .ZN(n752) );
  AOI22_X1 U328 ( .A1(data_in[0]), .A2(n832), .B1(n386), .B2(\mem[16][0] ), 
        .ZN(n385) );
  INV_X1 U329 ( .A(n387), .ZN(n751) );
  AOI22_X1 U330 ( .A1(data_in[1]), .A2(n832), .B1(n386), .B2(\mem[16][1] ), 
        .ZN(n387) );
  INV_X1 U331 ( .A(n388), .ZN(n750) );
  AOI22_X1 U332 ( .A1(data_in[2]), .A2(n832), .B1(n386), .B2(\mem[16][2] ), 
        .ZN(n388) );
  INV_X1 U333 ( .A(n389), .ZN(n749) );
  AOI22_X1 U334 ( .A1(data_in[3]), .A2(n832), .B1(n386), .B2(\mem[16][3] ), 
        .ZN(n389) );
  INV_X1 U335 ( .A(n390), .ZN(n748) );
  AOI22_X1 U336 ( .A1(data_in[4]), .A2(n832), .B1(n386), .B2(\mem[16][4] ), 
        .ZN(n390) );
  INV_X1 U337 ( .A(n391), .ZN(n747) );
  AOI22_X1 U338 ( .A1(data_in[5]), .A2(n832), .B1(n386), .B2(\mem[16][5] ), 
        .ZN(n391) );
  INV_X1 U339 ( .A(n392), .ZN(n746) );
  AOI22_X1 U340 ( .A1(data_in[6]), .A2(n832), .B1(n386), .B2(\mem[16][6] ), 
        .ZN(n392) );
  INV_X1 U341 ( .A(n393), .ZN(n745) );
  AOI22_X1 U342 ( .A1(data_in[7]), .A2(n832), .B1(n386), .B2(\mem[16][7] ), 
        .ZN(n393) );
  INV_X1 U343 ( .A(n395), .ZN(n744) );
  AOI22_X1 U344 ( .A1(data_in[0]), .A2(n831), .B1(n396), .B2(\mem[17][0] ), 
        .ZN(n395) );
  INV_X1 U345 ( .A(n397), .ZN(n743) );
  AOI22_X1 U346 ( .A1(data_in[1]), .A2(n831), .B1(n396), .B2(\mem[17][1] ), 
        .ZN(n397) );
  INV_X1 U347 ( .A(n398), .ZN(n742) );
  AOI22_X1 U348 ( .A1(data_in[2]), .A2(n831), .B1(n396), .B2(\mem[17][2] ), 
        .ZN(n398) );
  INV_X1 U349 ( .A(n399), .ZN(n741) );
  AOI22_X1 U350 ( .A1(data_in[3]), .A2(n831), .B1(n396), .B2(\mem[17][3] ), 
        .ZN(n399) );
  INV_X1 U351 ( .A(n400), .ZN(n740) );
  AOI22_X1 U352 ( .A1(data_in[4]), .A2(n831), .B1(n396), .B2(\mem[17][4] ), 
        .ZN(n400) );
  INV_X1 U353 ( .A(n401), .ZN(n739) );
  AOI22_X1 U354 ( .A1(data_in[5]), .A2(n831), .B1(n396), .B2(\mem[17][5] ), 
        .ZN(n401) );
  INV_X1 U355 ( .A(n402), .ZN(n738) );
  AOI22_X1 U356 ( .A1(data_in[6]), .A2(n831), .B1(n396), .B2(\mem[17][6] ), 
        .ZN(n402) );
  INV_X1 U357 ( .A(n403), .ZN(n737) );
  AOI22_X1 U358 ( .A1(data_in[7]), .A2(n831), .B1(n396), .B2(\mem[17][7] ), 
        .ZN(n403) );
  INV_X1 U359 ( .A(n404), .ZN(n736) );
  AOI22_X1 U360 ( .A1(data_in[0]), .A2(n830), .B1(n405), .B2(\mem[18][0] ), 
        .ZN(n404) );
  INV_X1 U361 ( .A(n406), .ZN(n735) );
  AOI22_X1 U362 ( .A1(data_in[1]), .A2(n830), .B1(n405), .B2(\mem[18][1] ), 
        .ZN(n406) );
  INV_X1 U363 ( .A(n407), .ZN(n734) );
  AOI22_X1 U364 ( .A1(data_in[2]), .A2(n830), .B1(n405), .B2(\mem[18][2] ), 
        .ZN(n407) );
  INV_X1 U365 ( .A(n408), .ZN(n733) );
  AOI22_X1 U366 ( .A1(data_in[3]), .A2(n830), .B1(n405), .B2(\mem[18][3] ), 
        .ZN(n408) );
  INV_X1 U367 ( .A(n409), .ZN(n732) );
  AOI22_X1 U368 ( .A1(data_in[4]), .A2(n830), .B1(n405), .B2(\mem[18][4] ), 
        .ZN(n409) );
  INV_X1 U369 ( .A(n410), .ZN(n731) );
  AOI22_X1 U370 ( .A1(data_in[5]), .A2(n830), .B1(n405), .B2(\mem[18][5] ), 
        .ZN(n410) );
  INV_X1 U371 ( .A(n411), .ZN(n730) );
  AOI22_X1 U372 ( .A1(data_in[6]), .A2(n830), .B1(n405), .B2(\mem[18][6] ), 
        .ZN(n411) );
  INV_X1 U373 ( .A(n412), .ZN(n729) );
  AOI22_X1 U374 ( .A1(data_in[7]), .A2(n830), .B1(n405), .B2(\mem[18][7] ), 
        .ZN(n412) );
  INV_X1 U375 ( .A(n413), .ZN(n728) );
  AOI22_X1 U376 ( .A1(data_in[0]), .A2(n829), .B1(n414), .B2(\mem[19][0] ), 
        .ZN(n413) );
  INV_X1 U377 ( .A(n415), .ZN(n727) );
  AOI22_X1 U378 ( .A1(data_in[1]), .A2(n829), .B1(n414), .B2(\mem[19][1] ), 
        .ZN(n415) );
  INV_X1 U379 ( .A(n416), .ZN(n726) );
  AOI22_X1 U380 ( .A1(data_in[2]), .A2(n829), .B1(n414), .B2(\mem[19][2] ), 
        .ZN(n416) );
  INV_X1 U381 ( .A(n417), .ZN(n725) );
  AOI22_X1 U382 ( .A1(data_in[3]), .A2(n829), .B1(n414), .B2(\mem[19][3] ), 
        .ZN(n417) );
  INV_X1 U383 ( .A(n418), .ZN(n724) );
  AOI22_X1 U384 ( .A1(data_in[4]), .A2(n829), .B1(n414), .B2(\mem[19][4] ), 
        .ZN(n418) );
  INV_X1 U385 ( .A(n419), .ZN(n723) );
  AOI22_X1 U386 ( .A1(data_in[5]), .A2(n829), .B1(n414), .B2(\mem[19][5] ), 
        .ZN(n419) );
  INV_X1 U387 ( .A(n420), .ZN(n722) );
  AOI22_X1 U388 ( .A1(data_in[6]), .A2(n829), .B1(n414), .B2(\mem[19][6] ), 
        .ZN(n420) );
  INV_X1 U389 ( .A(n421), .ZN(n721) );
  AOI22_X1 U390 ( .A1(data_in[7]), .A2(n829), .B1(n414), .B2(\mem[19][7] ), 
        .ZN(n421) );
  INV_X1 U391 ( .A(n422), .ZN(n720) );
  AOI22_X1 U392 ( .A1(data_in[0]), .A2(n828), .B1(n423), .B2(\mem[20][0] ), 
        .ZN(n422) );
  INV_X1 U393 ( .A(n424), .ZN(n719) );
  AOI22_X1 U394 ( .A1(data_in[1]), .A2(n828), .B1(n423), .B2(\mem[20][1] ), 
        .ZN(n424) );
  INV_X1 U395 ( .A(n425), .ZN(n718) );
  AOI22_X1 U396 ( .A1(data_in[2]), .A2(n828), .B1(n423), .B2(\mem[20][2] ), 
        .ZN(n425) );
  INV_X1 U397 ( .A(n426), .ZN(n717) );
  AOI22_X1 U398 ( .A1(data_in[3]), .A2(n828), .B1(n423), .B2(\mem[20][3] ), 
        .ZN(n426) );
  INV_X1 U399 ( .A(n427), .ZN(n716) );
  AOI22_X1 U400 ( .A1(data_in[4]), .A2(n828), .B1(n423), .B2(\mem[20][4] ), 
        .ZN(n427) );
  INV_X1 U401 ( .A(n428), .ZN(n715) );
  AOI22_X1 U402 ( .A1(data_in[5]), .A2(n828), .B1(n423), .B2(\mem[20][5] ), 
        .ZN(n428) );
  INV_X1 U403 ( .A(n429), .ZN(n714) );
  AOI22_X1 U404 ( .A1(data_in[6]), .A2(n828), .B1(n423), .B2(\mem[20][6] ), 
        .ZN(n429) );
  INV_X1 U405 ( .A(n430), .ZN(n713) );
  AOI22_X1 U406 ( .A1(data_in[7]), .A2(n828), .B1(n423), .B2(\mem[20][7] ), 
        .ZN(n430) );
  INV_X1 U407 ( .A(n431), .ZN(n712) );
  AOI22_X1 U408 ( .A1(data_in[0]), .A2(n827), .B1(n432), .B2(\mem[21][0] ), 
        .ZN(n431) );
  INV_X1 U409 ( .A(n433), .ZN(n711) );
  AOI22_X1 U410 ( .A1(data_in[1]), .A2(n827), .B1(n432), .B2(\mem[21][1] ), 
        .ZN(n433) );
  INV_X1 U411 ( .A(n434), .ZN(n710) );
  AOI22_X1 U412 ( .A1(data_in[2]), .A2(n827), .B1(n432), .B2(\mem[21][2] ), 
        .ZN(n434) );
  INV_X1 U413 ( .A(n435), .ZN(n709) );
  AOI22_X1 U414 ( .A1(data_in[3]), .A2(n827), .B1(n432), .B2(\mem[21][3] ), 
        .ZN(n435) );
  INV_X1 U415 ( .A(n436), .ZN(n708) );
  AOI22_X1 U416 ( .A1(data_in[4]), .A2(n827), .B1(n432), .B2(\mem[21][4] ), 
        .ZN(n436) );
  INV_X1 U417 ( .A(n437), .ZN(n707) );
  AOI22_X1 U418 ( .A1(data_in[5]), .A2(n827), .B1(n432), .B2(\mem[21][5] ), 
        .ZN(n437) );
  INV_X1 U419 ( .A(n438), .ZN(n706) );
  AOI22_X1 U420 ( .A1(data_in[6]), .A2(n827), .B1(n432), .B2(\mem[21][6] ), 
        .ZN(n438) );
  INV_X1 U421 ( .A(n439), .ZN(n705) );
  AOI22_X1 U422 ( .A1(data_in[7]), .A2(n827), .B1(n432), .B2(\mem[21][7] ), 
        .ZN(n439) );
  INV_X1 U423 ( .A(n440), .ZN(n704) );
  AOI22_X1 U424 ( .A1(data_in[0]), .A2(n826), .B1(n441), .B2(\mem[22][0] ), 
        .ZN(n440) );
  INV_X1 U425 ( .A(n442), .ZN(n703) );
  AOI22_X1 U426 ( .A1(data_in[1]), .A2(n826), .B1(n441), .B2(\mem[22][1] ), 
        .ZN(n442) );
  INV_X1 U427 ( .A(n443), .ZN(n702) );
  AOI22_X1 U428 ( .A1(data_in[2]), .A2(n826), .B1(n441), .B2(\mem[22][2] ), 
        .ZN(n443) );
  INV_X1 U429 ( .A(n444), .ZN(n701) );
  AOI22_X1 U430 ( .A1(data_in[3]), .A2(n826), .B1(n441), .B2(\mem[22][3] ), 
        .ZN(n444) );
  INV_X1 U431 ( .A(n445), .ZN(n700) );
  AOI22_X1 U432 ( .A1(data_in[4]), .A2(n826), .B1(n441), .B2(\mem[22][4] ), 
        .ZN(n445) );
  INV_X1 U433 ( .A(n446), .ZN(n699) );
  AOI22_X1 U434 ( .A1(data_in[5]), .A2(n826), .B1(n441), .B2(\mem[22][5] ), 
        .ZN(n446) );
  INV_X1 U435 ( .A(n447), .ZN(n698) );
  AOI22_X1 U436 ( .A1(data_in[6]), .A2(n826), .B1(n441), .B2(\mem[22][6] ), 
        .ZN(n447) );
  INV_X1 U437 ( .A(n448), .ZN(n697) );
  AOI22_X1 U438 ( .A1(data_in[7]), .A2(n826), .B1(n441), .B2(\mem[22][7] ), 
        .ZN(n448) );
  INV_X1 U439 ( .A(n449), .ZN(n696) );
  AOI22_X1 U440 ( .A1(data_in[0]), .A2(n825), .B1(n450), .B2(\mem[23][0] ), 
        .ZN(n449) );
  INV_X1 U441 ( .A(n451), .ZN(n695) );
  AOI22_X1 U442 ( .A1(data_in[1]), .A2(n825), .B1(n450), .B2(\mem[23][1] ), 
        .ZN(n451) );
  INV_X1 U443 ( .A(n452), .ZN(n694) );
  AOI22_X1 U444 ( .A1(data_in[2]), .A2(n825), .B1(n450), .B2(\mem[23][2] ), 
        .ZN(n452) );
  INV_X1 U445 ( .A(n453), .ZN(n693) );
  AOI22_X1 U446 ( .A1(data_in[3]), .A2(n825), .B1(n450), .B2(\mem[23][3] ), 
        .ZN(n453) );
  INV_X1 U447 ( .A(n454), .ZN(n692) );
  AOI22_X1 U448 ( .A1(data_in[4]), .A2(n825), .B1(n450), .B2(\mem[23][4] ), 
        .ZN(n454) );
  INV_X1 U449 ( .A(n455), .ZN(n691) );
  AOI22_X1 U450 ( .A1(data_in[5]), .A2(n825), .B1(n450), .B2(\mem[23][5] ), 
        .ZN(n455) );
  INV_X1 U451 ( .A(n456), .ZN(n690) );
  AOI22_X1 U452 ( .A1(data_in[6]), .A2(n825), .B1(n450), .B2(\mem[23][6] ), 
        .ZN(n456) );
  INV_X1 U453 ( .A(n457), .ZN(n689) );
  AOI22_X1 U454 ( .A1(data_in[7]), .A2(n825), .B1(n450), .B2(\mem[23][7] ), 
        .ZN(n457) );
  INV_X1 U455 ( .A(n458), .ZN(n688) );
  AOI22_X1 U456 ( .A1(data_in[0]), .A2(n824), .B1(n459), .B2(\mem[24][0] ), 
        .ZN(n458) );
  INV_X1 U457 ( .A(n460), .ZN(n687) );
  AOI22_X1 U458 ( .A1(data_in[1]), .A2(n824), .B1(n459), .B2(\mem[24][1] ), 
        .ZN(n460) );
  INV_X1 U459 ( .A(n461), .ZN(n686) );
  AOI22_X1 U460 ( .A1(data_in[2]), .A2(n824), .B1(n459), .B2(\mem[24][2] ), 
        .ZN(n461) );
  INV_X1 U461 ( .A(n462), .ZN(n685) );
  AOI22_X1 U462 ( .A1(data_in[3]), .A2(n824), .B1(n459), .B2(\mem[24][3] ), 
        .ZN(n462) );
  INV_X1 U463 ( .A(n463), .ZN(n684) );
  AOI22_X1 U464 ( .A1(data_in[4]), .A2(n824), .B1(n459), .B2(\mem[24][4] ), 
        .ZN(n463) );
  INV_X1 U465 ( .A(n464), .ZN(n683) );
  AOI22_X1 U466 ( .A1(data_in[5]), .A2(n824), .B1(n459), .B2(\mem[24][5] ), 
        .ZN(n464) );
  INV_X1 U467 ( .A(n465), .ZN(n682) );
  AOI22_X1 U468 ( .A1(data_in[6]), .A2(n824), .B1(n459), .B2(\mem[24][6] ), 
        .ZN(n465) );
  INV_X1 U469 ( .A(n466), .ZN(n681) );
  AOI22_X1 U470 ( .A1(data_in[7]), .A2(n824), .B1(n459), .B2(\mem[24][7] ), 
        .ZN(n466) );
  INV_X1 U471 ( .A(n468), .ZN(n680) );
  AOI22_X1 U472 ( .A1(data_in[0]), .A2(n823), .B1(n469), .B2(\mem[25][0] ), 
        .ZN(n468) );
  INV_X1 U473 ( .A(n470), .ZN(n679) );
  AOI22_X1 U474 ( .A1(data_in[1]), .A2(n823), .B1(n469), .B2(\mem[25][1] ), 
        .ZN(n470) );
  INV_X1 U475 ( .A(n471), .ZN(n678) );
  AOI22_X1 U476 ( .A1(data_in[2]), .A2(n823), .B1(n469), .B2(\mem[25][2] ), 
        .ZN(n471) );
  INV_X1 U477 ( .A(n472), .ZN(n677) );
  AOI22_X1 U478 ( .A1(data_in[3]), .A2(n823), .B1(n469), .B2(\mem[25][3] ), 
        .ZN(n472) );
  INV_X1 U479 ( .A(n473), .ZN(n676) );
  AOI22_X1 U480 ( .A1(data_in[4]), .A2(n823), .B1(n469), .B2(\mem[25][4] ), 
        .ZN(n473) );
  INV_X1 U481 ( .A(n474), .ZN(n675) );
  AOI22_X1 U482 ( .A1(data_in[5]), .A2(n823), .B1(n469), .B2(\mem[25][5] ), 
        .ZN(n474) );
  INV_X1 U483 ( .A(n475), .ZN(n674) );
  AOI22_X1 U484 ( .A1(data_in[6]), .A2(n823), .B1(n469), .B2(\mem[25][6] ), 
        .ZN(n475) );
  INV_X1 U485 ( .A(n476), .ZN(n673) );
  AOI22_X1 U486 ( .A1(data_in[7]), .A2(n823), .B1(n469), .B2(\mem[25][7] ), 
        .ZN(n476) );
  INV_X1 U487 ( .A(n477), .ZN(n672) );
  AOI22_X1 U488 ( .A1(data_in[0]), .A2(n822), .B1(n478), .B2(\mem[26][0] ), 
        .ZN(n477) );
  INV_X1 U489 ( .A(n479), .ZN(n671) );
  AOI22_X1 U490 ( .A1(data_in[1]), .A2(n822), .B1(n478), .B2(\mem[26][1] ), 
        .ZN(n479) );
  INV_X1 U491 ( .A(n480), .ZN(n670) );
  AOI22_X1 U492 ( .A1(data_in[2]), .A2(n822), .B1(n478), .B2(\mem[26][2] ), 
        .ZN(n480) );
  INV_X1 U493 ( .A(n481), .ZN(n669) );
  AOI22_X1 U494 ( .A1(data_in[3]), .A2(n822), .B1(n478), .B2(\mem[26][3] ), 
        .ZN(n481) );
  INV_X1 U495 ( .A(n482), .ZN(n668) );
  AOI22_X1 U496 ( .A1(data_in[4]), .A2(n822), .B1(n478), .B2(\mem[26][4] ), 
        .ZN(n482) );
  INV_X1 U497 ( .A(n483), .ZN(n667) );
  AOI22_X1 U498 ( .A1(data_in[5]), .A2(n822), .B1(n478), .B2(\mem[26][5] ), 
        .ZN(n483) );
  INV_X1 U499 ( .A(n484), .ZN(n666) );
  AOI22_X1 U500 ( .A1(data_in[6]), .A2(n822), .B1(n478), .B2(\mem[26][6] ), 
        .ZN(n484) );
  INV_X1 U501 ( .A(n485), .ZN(n665) );
  AOI22_X1 U502 ( .A1(data_in[7]), .A2(n822), .B1(n478), .B2(\mem[26][7] ), 
        .ZN(n485) );
  INV_X1 U503 ( .A(n486), .ZN(n664) );
  AOI22_X1 U504 ( .A1(data_in[0]), .A2(n821), .B1(n487), .B2(\mem[27][0] ), 
        .ZN(n486) );
  INV_X1 U505 ( .A(n488), .ZN(n663) );
  AOI22_X1 U506 ( .A1(data_in[1]), .A2(n821), .B1(n487), .B2(\mem[27][1] ), 
        .ZN(n488) );
  INV_X1 U507 ( .A(n489), .ZN(n662) );
  AOI22_X1 U508 ( .A1(data_in[2]), .A2(n821), .B1(n487), .B2(\mem[27][2] ), 
        .ZN(n489) );
  INV_X1 U509 ( .A(n490), .ZN(n661) );
  AOI22_X1 U510 ( .A1(data_in[3]), .A2(n821), .B1(n487), .B2(\mem[27][3] ), 
        .ZN(n490) );
  INV_X1 U511 ( .A(n491), .ZN(n660) );
  AOI22_X1 U512 ( .A1(data_in[4]), .A2(n821), .B1(n487), .B2(\mem[27][4] ), 
        .ZN(n491) );
  INV_X1 U513 ( .A(n492), .ZN(n659) );
  AOI22_X1 U514 ( .A1(data_in[5]), .A2(n821), .B1(n487), .B2(\mem[27][5] ), 
        .ZN(n492) );
  INV_X1 U515 ( .A(n493), .ZN(n658) );
  AOI22_X1 U516 ( .A1(data_in[6]), .A2(n821), .B1(n487), .B2(\mem[27][6] ), 
        .ZN(n493) );
  INV_X1 U517 ( .A(n494), .ZN(n657) );
  AOI22_X1 U518 ( .A1(data_in[7]), .A2(n821), .B1(n487), .B2(\mem[27][7] ), 
        .ZN(n494) );
  INV_X1 U519 ( .A(n495), .ZN(n656) );
  AOI22_X1 U520 ( .A1(data_in[0]), .A2(n820), .B1(n496), .B2(\mem[28][0] ), 
        .ZN(n495) );
  INV_X1 U521 ( .A(n497), .ZN(n655) );
  AOI22_X1 U522 ( .A1(data_in[1]), .A2(n820), .B1(n496), .B2(\mem[28][1] ), 
        .ZN(n497) );
  INV_X1 U523 ( .A(n498), .ZN(n654) );
  AOI22_X1 U524 ( .A1(data_in[2]), .A2(n820), .B1(n496), .B2(\mem[28][2] ), 
        .ZN(n498) );
  INV_X1 U525 ( .A(n499), .ZN(n653) );
  AOI22_X1 U526 ( .A1(data_in[3]), .A2(n820), .B1(n496), .B2(\mem[28][3] ), 
        .ZN(n499) );
  INV_X1 U527 ( .A(n500), .ZN(n652) );
  AOI22_X1 U528 ( .A1(data_in[4]), .A2(n820), .B1(n496), .B2(\mem[28][4] ), 
        .ZN(n500) );
  INV_X1 U529 ( .A(n501), .ZN(n651) );
  AOI22_X1 U530 ( .A1(data_in[5]), .A2(n820), .B1(n496), .B2(\mem[28][5] ), 
        .ZN(n501) );
  INV_X1 U531 ( .A(n502), .ZN(n650) );
  AOI22_X1 U532 ( .A1(data_in[6]), .A2(n820), .B1(n496), .B2(\mem[28][6] ), 
        .ZN(n502) );
  INV_X1 U533 ( .A(n503), .ZN(n649) );
  AOI22_X1 U534 ( .A1(data_in[7]), .A2(n820), .B1(n496), .B2(\mem[28][7] ), 
        .ZN(n503) );
  INV_X1 U535 ( .A(n504), .ZN(n648) );
  AOI22_X1 U536 ( .A1(data_in[0]), .A2(n819), .B1(n505), .B2(\mem[29][0] ), 
        .ZN(n504) );
  INV_X1 U537 ( .A(n506), .ZN(n647) );
  AOI22_X1 U538 ( .A1(data_in[1]), .A2(n819), .B1(n505), .B2(\mem[29][1] ), 
        .ZN(n506) );
  INV_X1 U539 ( .A(n507), .ZN(n646) );
  AOI22_X1 U540 ( .A1(data_in[2]), .A2(n819), .B1(n505), .B2(\mem[29][2] ), 
        .ZN(n507) );
  INV_X1 U541 ( .A(n508), .ZN(n645) );
  AOI22_X1 U542 ( .A1(data_in[3]), .A2(n819), .B1(n505), .B2(\mem[29][3] ), 
        .ZN(n508) );
  INV_X1 U543 ( .A(n509), .ZN(n644) );
  AOI22_X1 U544 ( .A1(data_in[4]), .A2(n819), .B1(n505), .B2(\mem[29][4] ), 
        .ZN(n509) );
  INV_X1 U545 ( .A(n510), .ZN(n643) );
  AOI22_X1 U546 ( .A1(data_in[5]), .A2(n819), .B1(n505), .B2(\mem[29][5] ), 
        .ZN(n510) );
  INV_X1 U547 ( .A(n511), .ZN(n642) );
  AOI22_X1 U548 ( .A1(data_in[6]), .A2(n819), .B1(n505), .B2(\mem[29][6] ), 
        .ZN(n511) );
  INV_X1 U549 ( .A(n512), .ZN(n641) );
  AOI22_X1 U550 ( .A1(data_in[7]), .A2(n819), .B1(n505), .B2(\mem[29][7] ), 
        .ZN(n512) );
  INV_X1 U551 ( .A(n513), .ZN(n640) );
  AOI22_X1 U552 ( .A1(data_in[0]), .A2(n818), .B1(n514), .B2(\mem[30][0] ), 
        .ZN(n513) );
  INV_X1 U553 ( .A(n515), .ZN(n639) );
  AOI22_X1 U554 ( .A1(data_in[1]), .A2(n818), .B1(n514), .B2(\mem[30][1] ), 
        .ZN(n515) );
  INV_X1 U555 ( .A(n516), .ZN(n638) );
  AOI22_X1 U556 ( .A1(data_in[2]), .A2(n818), .B1(n514), .B2(\mem[30][2] ), 
        .ZN(n516) );
  INV_X1 U557 ( .A(n517), .ZN(n637) );
  AOI22_X1 U558 ( .A1(data_in[3]), .A2(n818), .B1(n514), .B2(\mem[30][3] ), 
        .ZN(n517) );
  INV_X1 U559 ( .A(n518), .ZN(n636) );
  AOI22_X1 U560 ( .A1(data_in[4]), .A2(n818), .B1(n514), .B2(\mem[30][4] ), 
        .ZN(n518) );
  INV_X1 U561 ( .A(n519), .ZN(n635) );
  AOI22_X1 U562 ( .A1(data_in[5]), .A2(n818), .B1(n514), .B2(\mem[30][5] ), 
        .ZN(n519) );
  INV_X1 U563 ( .A(n520), .ZN(n634) );
  AOI22_X1 U564 ( .A1(data_in[6]), .A2(n818), .B1(n514), .B2(\mem[30][6] ), 
        .ZN(n520) );
  INV_X1 U565 ( .A(n521), .ZN(n633) );
  AOI22_X1 U566 ( .A1(data_in[7]), .A2(n818), .B1(n514), .B2(\mem[30][7] ), 
        .ZN(n521) );
  INV_X1 U567 ( .A(n522), .ZN(n632) );
  AOI22_X1 U568 ( .A1(data_in[0]), .A2(n817), .B1(n523), .B2(\mem[31][0] ), 
        .ZN(n522) );
  INV_X1 U569 ( .A(n524), .ZN(n631) );
  AOI22_X1 U570 ( .A1(data_in[1]), .A2(n817), .B1(n523), .B2(\mem[31][1] ), 
        .ZN(n524) );
  INV_X1 U571 ( .A(n525), .ZN(n630) );
  AOI22_X1 U572 ( .A1(data_in[2]), .A2(n817), .B1(n523), .B2(\mem[31][2] ), 
        .ZN(n525) );
  INV_X1 U573 ( .A(n526), .ZN(n629) );
  AOI22_X1 U574 ( .A1(data_in[3]), .A2(n817), .B1(n523), .B2(\mem[31][3] ), 
        .ZN(n526) );
  INV_X1 U575 ( .A(n527), .ZN(n628) );
  AOI22_X1 U576 ( .A1(data_in[4]), .A2(n817), .B1(n523), .B2(\mem[31][4] ), 
        .ZN(n527) );
  INV_X1 U577 ( .A(n528), .ZN(n627) );
  AOI22_X1 U578 ( .A1(data_in[5]), .A2(n817), .B1(n523), .B2(\mem[31][5] ), 
        .ZN(n528) );
  INV_X1 U579 ( .A(n529), .ZN(n626) );
  AOI22_X1 U580 ( .A1(data_in[6]), .A2(n817), .B1(n523), .B2(\mem[31][6] ), 
        .ZN(n529) );
  INV_X1 U581 ( .A(n530), .ZN(n625) );
  AOI22_X1 U582 ( .A1(data_in[7]), .A2(n817), .B1(n523), .B2(\mem[31][7] ), 
        .ZN(n530) );
  NOR3_X1 U583 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n239) );
  NOR3_X1 U584 ( .A1(N11), .A2(N12), .A3(n615), .ZN(n250) );
  NOR3_X1 U585 ( .A1(N10), .A2(N12), .A3(n616), .ZN(n260) );
  NOR3_X1 U586 ( .A1(n615), .A2(N12), .A3(n616), .ZN(n270) );
  AND3_X1 U587 ( .A1(N11), .A2(n615), .A3(N12), .ZN(n300) );
  AND3_X1 U588 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n310) );
  AND3_X1 U589 ( .A1(n615), .A2(n616), .A3(N12), .ZN(n280) );
  AND3_X1 U590 ( .A1(N10), .A2(n616), .A3(N12), .ZN(n290) );
  INV_X1 U591 ( .A(N13), .ZN(n843) );
  BUF_X1 U592 ( .A(N12), .Z(n607) );
  INV_X1 U593 ( .A(N14), .ZN(n842) );
  MUX2_X1 U594 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n610), .Z(n2) );
  MUX2_X1 U595 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n610), .Z(n3) );
  MUX2_X1 U596 ( .A(n3), .B(n2), .S(N11), .Z(n4) );
  MUX2_X1 U597 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n610), .Z(n5) );
  MUX2_X1 U598 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n610), .Z(n6) );
  MUX2_X1 U599 ( .A(n6), .B(n5), .S(N11), .Z(n7) );
  MUX2_X1 U600 ( .A(n7), .B(n4), .S(n607), .Z(n8) );
  MUX2_X1 U601 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n610), .Z(n9) );
  MUX2_X1 U602 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n610), .Z(n10) );
  MUX2_X1 U603 ( .A(n10), .B(n9), .S(N11), .Z(n11) );
  MUX2_X1 U604 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n610), .Z(n12) );
  MUX2_X1 U605 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n610), .Z(n13) );
  MUX2_X1 U606 ( .A(n13), .B(n12), .S(N11), .Z(n14) );
  MUX2_X1 U607 ( .A(n14), .B(n11), .S(n607), .Z(n15) );
  MUX2_X1 U608 ( .A(n15), .B(n8), .S(N13), .Z(n16) );
  MUX2_X1 U609 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n614), .Z(n17) );
  MUX2_X1 U610 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(N10), .Z(n18) );
  MUX2_X1 U611 ( .A(n18), .B(n17), .S(n608), .Z(n19) );
  MUX2_X1 U612 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n614), .Z(n20) );
  MUX2_X1 U613 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n610), .Z(n21) );
  MUX2_X1 U614 ( .A(n21), .B(n20), .S(n608), .Z(n22) );
  MUX2_X1 U615 ( .A(n22), .B(n19), .S(n607), .Z(n23) );
  MUX2_X1 U616 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(N10), .Z(n24) );
  MUX2_X1 U617 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n614), .Z(n25) );
  MUX2_X1 U618 ( .A(n25), .B(n24), .S(n608), .Z(n26) );
  MUX2_X1 U619 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n613), .Z(n27) );
  MUX2_X1 U620 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n612), .Z(n28) );
  MUX2_X1 U621 ( .A(n28), .B(n27), .S(n608), .Z(n29) );
  MUX2_X1 U622 ( .A(n29), .B(n26), .S(n607), .Z(n30) );
  MUX2_X1 U623 ( .A(n30), .B(n23), .S(N13), .Z(n31) );
  MUX2_X1 U624 ( .A(n31), .B(n16), .S(N14), .Z(N22) );
  MUX2_X1 U625 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n612), .Z(n32) );
  MUX2_X1 U626 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n612), .Z(n33) );
  MUX2_X1 U627 ( .A(n33), .B(n32), .S(n608), .Z(n34) );
  MUX2_X1 U628 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n614), .Z(n35) );
  MUX2_X1 U629 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n612), .Z(n36) );
  MUX2_X1 U630 ( .A(n36), .B(n35), .S(n608), .Z(n37) );
  MUX2_X1 U631 ( .A(n37), .B(n34), .S(n607), .Z(n38) );
  MUX2_X1 U632 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n614), .Z(n39) );
  MUX2_X1 U633 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n611), .Z(n40) );
  MUX2_X1 U634 ( .A(n40), .B(n39), .S(n608), .Z(n41) );
  MUX2_X1 U635 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n610), .Z(n42) );
  MUX2_X1 U636 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(N10), .Z(n43) );
  MUX2_X1 U637 ( .A(n43), .B(n42), .S(n608), .Z(n44) );
  MUX2_X1 U638 ( .A(n44), .B(n41), .S(n607), .Z(n45) );
  MUX2_X1 U639 ( .A(n45), .B(n38), .S(N13), .Z(n46) );
  MUX2_X1 U640 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n614), .Z(n47) );
  MUX2_X1 U641 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n613), .Z(n48) );
  MUX2_X1 U642 ( .A(n48), .B(n47), .S(n608), .Z(n49) );
  MUX2_X1 U643 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n612), .Z(n50) );
  MUX2_X1 U644 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n613), .Z(n51) );
  MUX2_X1 U645 ( .A(n51), .B(n50), .S(n608), .Z(n52) );
  MUX2_X1 U646 ( .A(n52), .B(n49), .S(n607), .Z(n53) );
  MUX2_X1 U647 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n613), .Z(n54) );
  MUX2_X1 U648 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n55) );
  MUX2_X1 U649 ( .A(n55), .B(n54), .S(n608), .Z(n56) );
  MUX2_X1 U650 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n613), .Z(n57) );
  MUX2_X1 U651 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n611), .Z(n58) );
  MUX2_X1 U652 ( .A(n58), .B(n57), .S(n608), .Z(n59) );
  MUX2_X1 U653 ( .A(n59), .B(n56), .S(n607), .Z(n60) );
  MUX2_X1 U654 ( .A(n60), .B(n53), .S(N13), .Z(n61) );
  MUX2_X1 U655 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n614), .Z(n62) );
  MUX2_X1 U656 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n614), .Z(n63) );
  MUX2_X1 U657 ( .A(n63), .B(n62), .S(n609), .Z(n64) );
  MUX2_X1 U658 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(N10), .Z(n65) );
  MUX2_X1 U659 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n614), .Z(n66) );
  MUX2_X1 U660 ( .A(n66), .B(n65), .S(n609), .Z(n67) );
  MUX2_X1 U661 ( .A(n67), .B(n64), .S(N12), .Z(n68) );
  MUX2_X1 U662 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(N10), .Z(n69) );
  MUX2_X1 U663 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(N10), .Z(n70) );
  MUX2_X1 U664 ( .A(n70), .B(n69), .S(n609), .Z(n71) );
  MUX2_X1 U665 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n614), .Z(n72) );
  MUX2_X1 U666 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n610), .Z(n73) );
  MUX2_X1 U667 ( .A(n73), .B(n72), .S(n609), .Z(n74) );
  MUX2_X1 U668 ( .A(n74), .B(n71), .S(n607), .Z(n75) );
  MUX2_X1 U669 ( .A(n75), .B(n68), .S(N13), .Z(n76) );
  MUX2_X1 U670 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(N10), .Z(n77) );
  MUX2_X1 U671 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n614), .Z(n78) );
  MUX2_X1 U672 ( .A(n78), .B(n77), .S(n609), .Z(n79) );
  MUX2_X1 U673 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n610), .Z(n80) );
  MUX2_X1 U674 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n610), .Z(n81) );
  MUX2_X1 U675 ( .A(n81), .B(n80), .S(n609), .Z(n82) );
  MUX2_X1 U676 ( .A(n82), .B(n79), .S(N12), .Z(n83) );
  MUX2_X1 U677 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n611), .Z(n84) );
  MUX2_X1 U678 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n611), .Z(n85) );
  MUX2_X1 U679 ( .A(n85), .B(n84), .S(n609), .Z(n86) );
  MUX2_X1 U680 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n611), .Z(n87) );
  MUX2_X1 U681 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n611), .Z(n88) );
  MUX2_X1 U682 ( .A(n88), .B(n87), .S(n609), .Z(n89) );
  MUX2_X1 U683 ( .A(n89), .B(n86), .S(n607), .Z(n90) );
  MUX2_X1 U684 ( .A(n90), .B(n83), .S(N13), .Z(n91) );
  MUX2_X1 U685 ( .A(n91), .B(n76), .S(N14), .Z(N20) );
  MUX2_X1 U686 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n611), .Z(n92) );
  MUX2_X1 U687 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n611), .Z(n93) );
  MUX2_X1 U688 ( .A(n93), .B(n92), .S(n609), .Z(n94) );
  MUX2_X1 U689 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n611), .Z(n95) );
  MUX2_X1 U690 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n611), .Z(n96) );
  MUX2_X1 U691 ( .A(n96), .B(n95), .S(n609), .Z(n97) );
  MUX2_X1 U692 ( .A(n97), .B(n94), .S(N12), .Z(n98) );
  MUX2_X1 U693 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n611), .Z(n99) );
  MUX2_X1 U694 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n611), .Z(n100) );
  MUX2_X1 U695 ( .A(n100), .B(n99), .S(n609), .Z(n101) );
  MUX2_X1 U696 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n611), .Z(n102) );
  MUX2_X1 U697 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n611), .Z(n103) );
  MUX2_X1 U698 ( .A(n103), .B(n102), .S(n609), .Z(n104) );
  MUX2_X1 U699 ( .A(n104), .B(n101), .S(n607), .Z(n105) );
  MUX2_X1 U700 ( .A(n105), .B(n98), .S(N13), .Z(n106) );
  MUX2_X1 U701 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n612), .Z(n107) );
  MUX2_X1 U702 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n612), .Z(n108) );
  MUX2_X1 U703 ( .A(n108), .B(n107), .S(N11), .Z(n109) );
  MUX2_X1 U704 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n612), .Z(n110) );
  MUX2_X1 U705 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n612), .Z(n111) );
  MUX2_X1 U706 ( .A(n111), .B(n110), .S(N11), .Z(n112) );
  MUX2_X1 U707 ( .A(n112), .B(n109), .S(N12), .Z(n113) );
  MUX2_X1 U708 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n612), .Z(n114) );
  MUX2_X1 U709 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n612), .Z(n115) );
  MUX2_X1 U710 ( .A(n115), .B(n114), .S(n608), .Z(n116) );
  MUX2_X1 U711 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n612), .Z(n117) );
  MUX2_X1 U712 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n612), .Z(n118) );
  MUX2_X1 U713 ( .A(n118), .B(n117), .S(n609), .Z(n119) );
  MUX2_X1 U714 ( .A(n119), .B(n116), .S(n607), .Z(n120) );
  MUX2_X1 U715 ( .A(n120), .B(n113), .S(N13), .Z(n121) );
  MUX2_X1 U716 ( .A(n121), .B(n106), .S(N14), .Z(N19) );
  MUX2_X1 U717 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n612), .Z(n122) );
  MUX2_X1 U718 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n612), .Z(n123) );
  MUX2_X1 U719 ( .A(n123), .B(n122), .S(N11), .Z(n124) );
  MUX2_X1 U720 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n612), .Z(n125) );
  MUX2_X1 U721 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n612), .Z(n126) );
  MUX2_X1 U722 ( .A(n126), .B(n125), .S(n608), .Z(n127) );
  MUX2_X1 U723 ( .A(n127), .B(n124), .S(N12), .Z(n128) );
  MUX2_X1 U724 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n610), .Z(n129) );
  MUX2_X1 U725 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(N10), .Z(n130) );
  MUX2_X1 U726 ( .A(n130), .B(n129), .S(n609), .Z(n131) );
  MUX2_X1 U727 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n614), .Z(n132) );
  MUX2_X1 U728 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n613), .Z(n133) );
  MUX2_X1 U729 ( .A(n133), .B(n132), .S(N11), .Z(n134) );
  MUX2_X1 U730 ( .A(n134), .B(n131), .S(n607), .Z(n135) );
  MUX2_X1 U731 ( .A(n135), .B(n128), .S(N13), .Z(n136) );
  MUX2_X1 U732 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n612), .Z(n137) );
  MUX2_X1 U733 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n614), .Z(n138) );
  MUX2_X1 U734 ( .A(n138), .B(n137), .S(n608), .Z(n139) );
  MUX2_X1 U735 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n614), .Z(n140) );
  MUX2_X1 U736 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n610), .Z(n141) );
  MUX2_X1 U737 ( .A(n141), .B(n140), .S(n609), .Z(n142) );
  MUX2_X1 U738 ( .A(n142), .B(n139), .S(N12), .Z(n143) );
  MUX2_X1 U739 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n611), .Z(n144) );
  MUX2_X1 U740 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n610), .Z(n145) );
  MUX2_X1 U741 ( .A(n145), .B(n144), .S(N11), .Z(n146) );
  MUX2_X1 U742 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n147) );
  MUX2_X1 U743 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n614), .Z(n148) );
  MUX2_X1 U744 ( .A(n148), .B(n147), .S(n608), .Z(n149) );
  MUX2_X1 U745 ( .A(n149), .B(n146), .S(n607), .Z(n150) );
  MUX2_X1 U746 ( .A(n150), .B(n143), .S(N13), .Z(n151) );
  MUX2_X1 U747 ( .A(n151), .B(n136), .S(N14), .Z(N18) );
  MUX2_X1 U748 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n613), .Z(n152) );
  MUX2_X1 U749 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n612), .Z(n153) );
  MUX2_X1 U750 ( .A(n153), .B(n152), .S(n608), .Z(n154) );
  MUX2_X1 U751 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n611), .Z(n155) );
  MUX2_X1 U752 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n610), .Z(n156) );
  MUX2_X1 U753 ( .A(n156), .B(n155), .S(n609), .Z(n157) );
  MUX2_X1 U754 ( .A(n157), .B(n154), .S(N12), .Z(n158) );
  MUX2_X1 U755 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(N10), .Z(n159) );
  MUX2_X1 U756 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n614), .Z(n160) );
  MUX2_X1 U757 ( .A(n160), .B(n159), .S(n609), .Z(n161) );
  MUX2_X1 U758 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n613), .Z(n162) );
  MUX2_X1 U759 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n612), .Z(n163) );
  MUX2_X1 U760 ( .A(n163), .B(n162), .S(N11), .Z(n164) );
  MUX2_X1 U761 ( .A(n164), .B(n161), .S(n607), .Z(n165) );
  MUX2_X1 U762 ( .A(n165), .B(n158), .S(N13), .Z(n166) );
  MUX2_X1 U763 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n611), .Z(n167) );
  MUX2_X1 U764 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n610), .Z(n168) );
  MUX2_X1 U765 ( .A(n168), .B(n167), .S(n608), .Z(n169) );
  MUX2_X1 U766 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(N10), .Z(n170) );
  MUX2_X1 U767 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n614), .Z(n171) );
  MUX2_X1 U768 ( .A(n171), .B(n170), .S(n609), .Z(n172) );
  MUX2_X1 U769 ( .A(n172), .B(n169), .S(N12), .Z(n173) );
  MUX2_X1 U770 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n613), .Z(n174) );
  MUX2_X1 U771 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n613), .Z(n175) );
  MUX2_X1 U772 ( .A(n175), .B(n174), .S(N11), .Z(n176) );
  MUX2_X1 U773 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n613), .Z(n177) );
  MUX2_X1 U774 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n613), .Z(n178) );
  MUX2_X1 U775 ( .A(n178), .B(n177), .S(N11), .Z(n179) );
  MUX2_X1 U776 ( .A(n179), .B(n176), .S(n607), .Z(n180) );
  MUX2_X1 U777 ( .A(n180), .B(n173), .S(N13), .Z(n181) );
  MUX2_X1 U778 ( .A(n181), .B(n166), .S(N14), .Z(N17) );
  MUX2_X1 U779 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n613), .Z(n182) );
  MUX2_X1 U780 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n613), .Z(n183) );
  MUX2_X1 U781 ( .A(n183), .B(n182), .S(n608), .Z(n184) );
  MUX2_X1 U782 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n613), .Z(n185) );
  MUX2_X1 U783 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n613), .Z(n186) );
  MUX2_X1 U784 ( .A(n186), .B(n185), .S(n609), .Z(n187) );
  MUX2_X1 U785 ( .A(n187), .B(n184), .S(N12), .Z(n188) );
  MUX2_X1 U786 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n613), .Z(n189) );
  MUX2_X1 U787 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n613), .Z(n190) );
  MUX2_X1 U788 ( .A(n190), .B(n189), .S(n608), .Z(n191) );
  MUX2_X1 U789 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n613), .Z(n192) );
  MUX2_X1 U790 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n613), .Z(n193) );
  MUX2_X1 U791 ( .A(n193), .B(n192), .S(N11), .Z(n194) );
  MUX2_X1 U792 ( .A(n194), .B(n191), .S(n607), .Z(n195) );
  MUX2_X1 U793 ( .A(n195), .B(n188), .S(N13), .Z(n196) );
  MUX2_X1 U794 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n614), .Z(n197) );
  MUX2_X1 U795 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n613), .Z(n198) );
  MUX2_X1 U796 ( .A(n198), .B(n197), .S(N11), .Z(n199) );
  MUX2_X1 U797 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n612), .Z(n200) );
  MUX2_X1 U798 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n201) );
  MUX2_X1 U799 ( .A(n201), .B(n200), .S(N11), .Z(n202) );
  MUX2_X1 U800 ( .A(n202), .B(n199), .S(N12), .Z(n203) );
  MUX2_X1 U801 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n611), .Z(n204) );
  MUX2_X1 U802 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n610), .Z(n205) );
  MUX2_X1 U803 ( .A(n205), .B(n204), .S(n608), .Z(n206) );
  MUX2_X1 U804 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n207) );
  MUX2_X1 U805 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n614), .Z(n208) );
  MUX2_X1 U806 ( .A(n208), .B(n207), .S(n609), .Z(n209) );
  MUX2_X1 U807 ( .A(n209), .B(n206), .S(n607), .Z(n210) );
  MUX2_X1 U808 ( .A(n210), .B(n203), .S(N13), .Z(n211) );
  MUX2_X1 U809 ( .A(n211), .B(n196), .S(N14), .Z(N16) );
  MUX2_X1 U810 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n613), .Z(n212) );
  MUX2_X1 U811 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n612), .Z(n213) );
  MUX2_X1 U812 ( .A(n213), .B(n212), .S(n609), .Z(n214) );
  MUX2_X1 U813 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n611), .Z(n215) );
  MUX2_X1 U814 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n611), .Z(n216) );
  MUX2_X1 U815 ( .A(n216), .B(n215), .S(n608), .Z(n217) );
  MUX2_X1 U816 ( .A(n217), .B(n214), .S(N12), .Z(n218) );
  MUX2_X1 U817 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n614), .Z(n219) );
  MUX2_X1 U818 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n610), .Z(n220) );
  MUX2_X1 U819 ( .A(n220), .B(n219), .S(N11), .Z(n221) );
  MUX2_X1 U820 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n610), .Z(n222) );
  MUX2_X1 U821 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n611), .Z(n223) );
  MUX2_X1 U822 ( .A(n223), .B(n222), .S(n608), .Z(n224) );
  MUX2_X1 U823 ( .A(n224), .B(n221), .S(N12), .Z(n225) );
  MUX2_X1 U824 ( .A(n225), .B(n218), .S(N13), .Z(n226) );
  MUX2_X1 U825 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n610), .Z(n227) );
  MUX2_X1 U826 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n228) );
  MUX2_X1 U827 ( .A(n228), .B(n227), .S(n609), .Z(n229) );
  MUX2_X1 U828 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n614), .Z(n595) );
  MUX2_X1 U829 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n613), .Z(n596) );
  MUX2_X1 U830 ( .A(n596), .B(n595), .S(N11), .Z(n597) );
  MUX2_X1 U831 ( .A(n597), .B(n229), .S(n607), .Z(n598) );
  MUX2_X1 U832 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n612), .Z(n599) );
  MUX2_X1 U833 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n600) );
  MUX2_X1 U834 ( .A(n600), .B(n599), .S(n609), .Z(n601) );
  MUX2_X1 U835 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n602) );
  MUX2_X1 U836 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n611), .Z(n603) );
  MUX2_X1 U837 ( .A(n603), .B(n602), .S(N11), .Z(n604) );
  MUX2_X1 U838 ( .A(n604), .B(n601), .S(N12), .Z(n605) );
  MUX2_X1 U839 ( .A(n605), .B(n598), .S(N13), .Z(n606) );
  CLKBUF_X1 U840 ( .A(n614), .Z(n610) );
  INV_X1 U841 ( .A(N10), .ZN(n615) );
  INV_X1 U842 ( .A(N11), .ZN(n616) );
  INV_X1 U843 ( .A(data_in[0]), .ZN(n617) );
  INV_X1 U844 ( .A(data_in[1]), .ZN(n618) );
  INV_X1 U845 ( .A(data_in[2]), .ZN(n619) );
  INV_X1 U846 ( .A(data_in[3]), .ZN(n620) );
  INV_X1 U847 ( .A(data_in[4]), .ZN(n621) );
  INV_X1 U848 ( .A(data_in[5]), .ZN(n622) );
  INV_X1 U849 ( .A(data_in[6]), .ZN(n623) );
  INV_X1 U850 ( .A(data_in[7]), .ZN(n624) );
endmodule


module memory_WIDTH8_SIZE1024_LOGSIZE12 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [11:0] addr;
  input clk, wr_en;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, \mem[1023][7] ,
         \mem[1023][6] , \mem[1023][5] , \mem[1023][4] , \mem[1023][3] ,
         \mem[1023][2] , \mem[1023][1] , \mem[1023][0] , \mem[1022][7] ,
         \mem[1022][6] , \mem[1022][5] , \mem[1022][4] , \mem[1022][3] ,
         \mem[1022][2] , \mem[1022][1] , \mem[1022][0] , \mem[1021][7] ,
         \mem[1021][6] , \mem[1021][5] , \mem[1021][4] , \mem[1021][3] ,
         \mem[1021][2] , \mem[1021][1] , \mem[1021][0] , \mem[1020][7] ,
         \mem[1020][6] , \mem[1020][5] , \mem[1020][4] , \mem[1020][3] ,
         \mem[1020][2] , \mem[1020][1] , \mem[1020][0] , \mem[1019][7] ,
         \mem[1019][6] , \mem[1019][5] , \mem[1019][4] , \mem[1019][3] ,
         \mem[1019][2] , \mem[1019][1] , \mem[1019][0] , \mem[1018][7] ,
         \mem[1018][6] , \mem[1018][5] , \mem[1018][4] , \mem[1018][3] ,
         \mem[1018][2] , \mem[1018][1] , \mem[1018][0] , \mem[1017][7] ,
         \mem[1017][6] , \mem[1017][5] , \mem[1017][4] , \mem[1017][3] ,
         \mem[1017][2] , \mem[1017][1] , \mem[1017][0] , \mem[1016][7] ,
         \mem[1016][6] , \mem[1016][5] , \mem[1016][4] , \mem[1016][3] ,
         \mem[1016][2] , \mem[1016][1] , \mem[1016][0] , \mem[1015][7] ,
         \mem[1015][6] , \mem[1015][5] , \mem[1015][4] , \mem[1015][3] ,
         \mem[1015][2] , \mem[1015][1] , \mem[1015][0] , \mem[1014][7] ,
         \mem[1014][6] , \mem[1014][5] , \mem[1014][4] , \mem[1014][3] ,
         \mem[1014][2] , \mem[1014][1] , \mem[1014][0] , \mem[1013][7] ,
         \mem[1013][6] , \mem[1013][5] , \mem[1013][4] , \mem[1013][3] ,
         \mem[1013][2] , \mem[1013][1] , \mem[1013][0] , \mem[1012][7] ,
         \mem[1012][6] , \mem[1012][5] , \mem[1012][4] , \mem[1012][3] ,
         \mem[1012][2] , \mem[1012][1] , \mem[1012][0] , \mem[1011][7] ,
         \mem[1011][6] , \mem[1011][5] , \mem[1011][4] , \mem[1011][3] ,
         \mem[1011][2] , \mem[1011][1] , \mem[1011][0] , \mem[1010][7] ,
         \mem[1010][6] , \mem[1010][5] , \mem[1010][4] , \mem[1010][3] ,
         \mem[1010][2] , \mem[1010][1] , \mem[1010][0] , \mem[1009][7] ,
         \mem[1009][6] , \mem[1009][5] , \mem[1009][4] , \mem[1009][3] ,
         \mem[1009][2] , \mem[1009][1] , \mem[1009][0] , \mem[1008][7] ,
         \mem[1008][6] , \mem[1008][5] , \mem[1008][4] , \mem[1008][3] ,
         \mem[1008][2] , \mem[1008][1] , \mem[1008][0] , \mem[1007][7] ,
         \mem[1007][6] , \mem[1007][5] , \mem[1007][4] , \mem[1007][3] ,
         \mem[1007][2] , \mem[1007][1] , \mem[1007][0] , \mem[1006][7] ,
         \mem[1006][6] , \mem[1006][5] , \mem[1006][4] , \mem[1006][3] ,
         \mem[1006][2] , \mem[1006][1] , \mem[1006][0] , \mem[1005][7] ,
         \mem[1005][6] , \mem[1005][5] , \mem[1005][4] , \mem[1005][3] ,
         \mem[1005][2] , \mem[1005][1] , \mem[1005][0] , \mem[1004][7] ,
         \mem[1004][6] , \mem[1004][5] , \mem[1004][4] , \mem[1004][3] ,
         \mem[1004][2] , \mem[1004][1] , \mem[1004][0] , \mem[1003][7] ,
         \mem[1003][6] , \mem[1003][5] , \mem[1003][4] , \mem[1003][3] ,
         \mem[1003][2] , \mem[1003][1] , \mem[1003][0] , \mem[1002][7] ,
         \mem[1002][6] , \mem[1002][5] , \mem[1002][4] , \mem[1002][3] ,
         \mem[1002][2] , \mem[1002][1] , \mem[1002][0] , \mem[1001][7] ,
         \mem[1001][6] , \mem[1001][5] , \mem[1001][4] , \mem[1001][3] ,
         \mem[1001][2] , \mem[1001][1] , \mem[1001][0] , \mem[1000][7] ,
         \mem[1000][6] , \mem[1000][5] , \mem[1000][4] , \mem[1000][3] ,
         \mem[1000][2] , \mem[1000][1] , \mem[1000][0] , \mem[999][7] ,
         \mem[999][6] , \mem[999][5] , \mem[999][4] , \mem[999][3] ,
         \mem[999][2] , \mem[999][1] , \mem[999][0] , \mem[998][7] ,
         \mem[998][6] , \mem[998][5] , \mem[998][4] , \mem[998][3] ,
         \mem[998][2] , \mem[998][1] , \mem[998][0] , \mem[997][7] ,
         \mem[997][6] , \mem[997][5] , \mem[997][4] , \mem[997][3] ,
         \mem[997][2] , \mem[997][1] , \mem[997][0] , \mem[996][7] ,
         \mem[996][6] , \mem[996][5] , \mem[996][4] , \mem[996][3] ,
         \mem[996][2] , \mem[996][1] , \mem[996][0] , \mem[995][7] ,
         \mem[995][6] , \mem[995][5] , \mem[995][4] , \mem[995][3] ,
         \mem[995][2] , \mem[995][1] , \mem[995][0] , \mem[994][7] ,
         \mem[994][6] , \mem[994][5] , \mem[994][4] , \mem[994][3] ,
         \mem[994][2] , \mem[994][1] , \mem[994][0] , \mem[993][7] ,
         \mem[993][6] , \mem[993][5] , \mem[993][4] , \mem[993][3] ,
         \mem[993][2] , \mem[993][1] , \mem[993][0] , \mem[992][7] ,
         \mem[992][6] , \mem[992][5] , \mem[992][4] , \mem[992][3] ,
         \mem[992][2] , \mem[992][1] , \mem[992][0] , \mem[991][7] ,
         \mem[991][6] , \mem[991][5] , \mem[991][4] , \mem[991][3] ,
         \mem[991][2] , \mem[991][1] , \mem[991][0] , \mem[990][7] ,
         \mem[990][6] , \mem[990][5] , \mem[990][4] , \mem[990][3] ,
         \mem[990][2] , \mem[990][1] , \mem[990][0] , \mem[989][7] ,
         \mem[989][6] , \mem[989][5] , \mem[989][4] , \mem[989][3] ,
         \mem[989][2] , \mem[989][1] , \mem[989][0] , \mem[988][7] ,
         \mem[988][6] , \mem[988][5] , \mem[988][4] , \mem[988][3] ,
         \mem[988][2] , \mem[988][1] , \mem[988][0] , \mem[987][7] ,
         \mem[987][6] , \mem[987][5] , \mem[987][4] , \mem[987][3] ,
         \mem[987][2] , \mem[987][1] , \mem[987][0] , \mem[986][7] ,
         \mem[986][6] , \mem[986][5] , \mem[986][4] , \mem[986][3] ,
         \mem[986][2] , \mem[986][1] , \mem[986][0] , \mem[985][7] ,
         \mem[985][6] , \mem[985][5] , \mem[985][4] , \mem[985][3] ,
         \mem[985][2] , \mem[985][1] , \mem[985][0] , \mem[984][7] ,
         \mem[984][6] , \mem[984][5] , \mem[984][4] , \mem[984][3] ,
         \mem[984][2] , \mem[984][1] , \mem[984][0] , \mem[983][7] ,
         \mem[983][6] , \mem[983][5] , \mem[983][4] , \mem[983][3] ,
         \mem[983][2] , \mem[983][1] , \mem[983][0] , \mem[982][7] ,
         \mem[982][6] , \mem[982][5] , \mem[982][4] , \mem[982][3] ,
         \mem[982][2] , \mem[982][1] , \mem[982][0] , \mem[981][7] ,
         \mem[981][6] , \mem[981][5] , \mem[981][4] , \mem[981][3] ,
         \mem[981][2] , \mem[981][1] , \mem[981][0] , \mem[980][7] ,
         \mem[980][6] , \mem[980][5] , \mem[980][4] , \mem[980][3] ,
         \mem[980][2] , \mem[980][1] , \mem[980][0] , \mem[979][7] ,
         \mem[979][6] , \mem[979][5] , \mem[979][4] , \mem[979][3] ,
         \mem[979][2] , \mem[979][1] , \mem[979][0] , \mem[978][7] ,
         \mem[978][6] , \mem[978][5] , \mem[978][4] , \mem[978][3] ,
         \mem[978][2] , \mem[978][1] , \mem[978][0] , \mem[977][7] ,
         \mem[977][6] , \mem[977][5] , \mem[977][4] , \mem[977][3] ,
         \mem[977][2] , \mem[977][1] , \mem[977][0] , \mem[976][7] ,
         \mem[976][6] , \mem[976][5] , \mem[976][4] , \mem[976][3] ,
         \mem[976][2] , \mem[976][1] , \mem[976][0] , \mem[975][7] ,
         \mem[975][6] , \mem[975][5] , \mem[975][4] , \mem[975][3] ,
         \mem[975][2] , \mem[975][1] , \mem[975][0] , \mem[974][7] ,
         \mem[974][6] , \mem[974][5] , \mem[974][4] , \mem[974][3] ,
         \mem[974][2] , \mem[974][1] , \mem[974][0] , \mem[973][7] ,
         \mem[973][6] , \mem[973][5] , \mem[973][4] , \mem[973][3] ,
         \mem[973][2] , \mem[973][1] , \mem[973][0] , \mem[972][7] ,
         \mem[972][6] , \mem[972][5] , \mem[972][4] , \mem[972][3] ,
         \mem[972][2] , \mem[972][1] , \mem[972][0] , \mem[971][7] ,
         \mem[971][6] , \mem[971][5] , \mem[971][4] , \mem[971][3] ,
         \mem[971][2] , \mem[971][1] , \mem[971][0] , \mem[970][7] ,
         \mem[970][6] , \mem[970][5] , \mem[970][4] , \mem[970][3] ,
         \mem[970][2] , \mem[970][1] , \mem[970][0] , \mem[969][7] ,
         \mem[969][6] , \mem[969][5] , \mem[969][4] , \mem[969][3] ,
         \mem[969][2] , \mem[969][1] , \mem[969][0] , \mem[968][7] ,
         \mem[968][6] , \mem[968][5] , \mem[968][4] , \mem[968][3] ,
         \mem[968][2] , \mem[968][1] , \mem[968][0] , \mem[967][7] ,
         \mem[967][6] , \mem[967][5] , \mem[967][4] , \mem[967][3] ,
         \mem[967][2] , \mem[967][1] , \mem[967][0] , \mem[966][7] ,
         \mem[966][6] , \mem[966][5] , \mem[966][4] , \mem[966][3] ,
         \mem[966][2] , \mem[966][1] , \mem[966][0] , \mem[965][7] ,
         \mem[965][6] , \mem[965][5] , \mem[965][4] , \mem[965][3] ,
         \mem[965][2] , \mem[965][1] , \mem[965][0] , \mem[964][7] ,
         \mem[964][6] , \mem[964][5] , \mem[964][4] , \mem[964][3] ,
         \mem[964][2] , \mem[964][1] , \mem[964][0] , \mem[963][7] ,
         \mem[963][6] , \mem[963][5] , \mem[963][4] , \mem[963][3] ,
         \mem[963][2] , \mem[963][1] , \mem[963][0] , \mem[962][7] ,
         \mem[962][6] , \mem[962][5] , \mem[962][4] , \mem[962][3] ,
         \mem[962][2] , \mem[962][1] , \mem[962][0] , \mem[961][7] ,
         \mem[961][6] , \mem[961][5] , \mem[961][4] , \mem[961][3] ,
         \mem[961][2] , \mem[961][1] , \mem[961][0] , \mem[960][7] ,
         \mem[960][6] , \mem[960][5] , \mem[960][4] , \mem[960][3] ,
         \mem[960][2] , \mem[960][1] , \mem[960][0] , \mem[959][7] ,
         \mem[959][6] , \mem[959][5] , \mem[959][4] , \mem[959][3] ,
         \mem[959][2] , \mem[959][1] , \mem[959][0] , \mem[958][7] ,
         \mem[958][6] , \mem[958][5] , \mem[958][4] , \mem[958][3] ,
         \mem[958][2] , \mem[958][1] , \mem[958][0] , \mem[957][7] ,
         \mem[957][6] , \mem[957][5] , \mem[957][4] , \mem[957][3] ,
         \mem[957][2] , \mem[957][1] , \mem[957][0] , \mem[956][7] ,
         \mem[956][6] , \mem[956][5] , \mem[956][4] , \mem[956][3] ,
         \mem[956][2] , \mem[956][1] , \mem[956][0] , \mem[955][7] ,
         \mem[955][6] , \mem[955][5] , \mem[955][4] , \mem[955][3] ,
         \mem[955][2] , \mem[955][1] , \mem[955][0] , \mem[954][7] ,
         \mem[954][6] , \mem[954][5] , \mem[954][4] , \mem[954][3] ,
         \mem[954][2] , \mem[954][1] , \mem[954][0] , \mem[953][7] ,
         \mem[953][6] , \mem[953][5] , \mem[953][4] , \mem[953][3] ,
         \mem[953][2] , \mem[953][1] , \mem[953][0] , \mem[952][7] ,
         \mem[952][6] , \mem[952][5] , \mem[952][4] , \mem[952][3] ,
         \mem[952][2] , \mem[952][1] , \mem[952][0] , \mem[951][7] ,
         \mem[951][6] , \mem[951][5] , \mem[951][4] , \mem[951][3] ,
         \mem[951][2] , \mem[951][1] , \mem[951][0] , \mem[950][7] ,
         \mem[950][6] , \mem[950][5] , \mem[950][4] , \mem[950][3] ,
         \mem[950][2] , \mem[950][1] , \mem[950][0] , \mem[949][7] ,
         \mem[949][6] , \mem[949][5] , \mem[949][4] , \mem[949][3] ,
         \mem[949][2] , \mem[949][1] , \mem[949][0] , \mem[948][7] ,
         \mem[948][6] , \mem[948][5] , \mem[948][4] , \mem[948][3] ,
         \mem[948][2] , \mem[948][1] , \mem[948][0] , \mem[947][7] ,
         \mem[947][6] , \mem[947][5] , \mem[947][4] , \mem[947][3] ,
         \mem[947][2] , \mem[947][1] , \mem[947][0] , \mem[946][7] ,
         \mem[946][6] , \mem[946][5] , \mem[946][4] , \mem[946][3] ,
         \mem[946][2] , \mem[946][1] , \mem[946][0] , \mem[945][7] ,
         \mem[945][6] , \mem[945][5] , \mem[945][4] , \mem[945][3] ,
         \mem[945][2] , \mem[945][1] , \mem[945][0] , \mem[944][7] ,
         \mem[944][6] , \mem[944][5] , \mem[944][4] , \mem[944][3] ,
         \mem[944][2] , \mem[944][1] , \mem[944][0] , \mem[943][7] ,
         \mem[943][6] , \mem[943][5] , \mem[943][4] , \mem[943][3] ,
         \mem[943][2] , \mem[943][1] , \mem[943][0] , \mem[942][7] ,
         \mem[942][6] , \mem[942][5] , \mem[942][4] , \mem[942][3] ,
         \mem[942][2] , \mem[942][1] , \mem[942][0] , \mem[941][7] ,
         \mem[941][6] , \mem[941][5] , \mem[941][4] , \mem[941][3] ,
         \mem[941][2] , \mem[941][1] , \mem[941][0] , \mem[940][7] ,
         \mem[940][6] , \mem[940][5] , \mem[940][4] , \mem[940][3] ,
         \mem[940][2] , \mem[940][1] , \mem[940][0] , \mem[939][7] ,
         \mem[939][6] , \mem[939][5] , \mem[939][4] , \mem[939][3] ,
         \mem[939][2] , \mem[939][1] , \mem[939][0] , \mem[938][7] ,
         \mem[938][6] , \mem[938][5] , \mem[938][4] , \mem[938][3] ,
         \mem[938][2] , \mem[938][1] , \mem[938][0] , \mem[937][7] ,
         \mem[937][6] , \mem[937][5] , \mem[937][4] , \mem[937][3] ,
         \mem[937][2] , \mem[937][1] , \mem[937][0] , \mem[936][7] ,
         \mem[936][6] , \mem[936][5] , \mem[936][4] , \mem[936][3] ,
         \mem[936][2] , \mem[936][1] , \mem[936][0] , \mem[935][7] ,
         \mem[935][6] , \mem[935][5] , \mem[935][4] , \mem[935][3] ,
         \mem[935][2] , \mem[935][1] , \mem[935][0] , \mem[934][7] ,
         \mem[934][6] , \mem[934][5] , \mem[934][4] , \mem[934][3] ,
         \mem[934][2] , \mem[934][1] , \mem[934][0] , \mem[933][7] ,
         \mem[933][6] , \mem[933][5] , \mem[933][4] , \mem[933][3] ,
         \mem[933][2] , \mem[933][1] , \mem[933][0] , \mem[932][7] ,
         \mem[932][6] , \mem[932][5] , \mem[932][4] , \mem[932][3] ,
         \mem[932][2] , \mem[932][1] , \mem[932][0] , \mem[931][7] ,
         \mem[931][6] , \mem[931][5] , \mem[931][4] , \mem[931][3] ,
         \mem[931][2] , \mem[931][1] , \mem[931][0] , \mem[930][7] ,
         \mem[930][6] , \mem[930][5] , \mem[930][4] , \mem[930][3] ,
         \mem[930][2] , \mem[930][1] , \mem[930][0] , \mem[929][7] ,
         \mem[929][6] , \mem[929][5] , \mem[929][4] , \mem[929][3] ,
         \mem[929][2] , \mem[929][1] , \mem[929][0] , \mem[928][7] ,
         \mem[928][6] , \mem[928][5] , \mem[928][4] , \mem[928][3] ,
         \mem[928][2] , \mem[928][1] , \mem[928][0] , \mem[927][7] ,
         \mem[927][6] , \mem[927][5] , \mem[927][4] , \mem[927][3] ,
         \mem[927][2] , \mem[927][1] , \mem[927][0] , \mem[926][7] ,
         \mem[926][6] , \mem[926][5] , \mem[926][4] , \mem[926][3] ,
         \mem[926][2] , \mem[926][1] , \mem[926][0] , \mem[925][7] ,
         \mem[925][6] , \mem[925][5] , \mem[925][4] , \mem[925][3] ,
         \mem[925][2] , \mem[925][1] , \mem[925][0] , \mem[924][7] ,
         \mem[924][6] , \mem[924][5] , \mem[924][4] , \mem[924][3] ,
         \mem[924][2] , \mem[924][1] , \mem[924][0] , \mem[923][7] ,
         \mem[923][6] , \mem[923][5] , \mem[923][4] , \mem[923][3] ,
         \mem[923][2] , \mem[923][1] , \mem[923][0] , \mem[922][7] ,
         \mem[922][6] , \mem[922][5] , \mem[922][4] , \mem[922][3] ,
         \mem[922][2] , \mem[922][1] , \mem[922][0] , \mem[921][7] ,
         \mem[921][6] , \mem[921][5] , \mem[921][4] , \mem[921][3] ,
         \mem[921][2] , \mem[921][1] , \mem[921][0] , \mem[920][7] ,
         \mem[920][6] , \mem[920][5] , \mem[920][4] , \mem[920][3] ,
         \mem[920][2] , \mem[920][1] , \mem[920][0] , \mem[919][7] ,
         \mem[919][6] , \mem[919][5] , \mem[919][4] , \mem[919][3] ,
         \mem[919][2] , \mem[919][1] , \mem[919][0] , \mem[918][7] ,
         \mem[918][6] , \mem[918][5] , \mem[918][4] , \mem[918][3] ,
         \mem[918][2] , \mem[918][1] , \mem[918][0] , \mem[917][7] ,
         \mem[917][6] , \mem[917][5] , \mem[917][4] , \mem[917][3] ,
         \mem[917][2] , \mem[917][1] , \mem[917][0] , \mem[916][7] ,
         \mem[916][6] , \mem[916][5] , \mem[916][4] , \mem[916][3] ,
         \mem[916][2] , \mem[916][1] , \mem[916][0] , \mem[915][7] ,
         \mem[915][6] , \mem[915][5] , \mem[915][4] , \mem[915][3] ,
         \mem[915][2] , \mem[915][1] , \mem[915][0] , \mem[914][7] ,
         \mem[914][6] , \mem[914][5] , \mem[914][4] , \mem[914][3] ,
         \mem[914][2] , \mem[914][1] , \mem[914][0] , \mem[913][7] ,
         \mem[913][6] , \mem[913][5] , \mem[913][4] , \mem[913][3] ,
         \mem[913][2] , \mem[913][1] , \mem[913][0] , \mem[912][7] ,
         \mem[912][6] , \mem[912][5] , \mem[912][4] , \mem[912][3] ,
         \mem[912][2] , \mem[912][1] , \mem[912][0] , \mem[911][7] ,
         \mem[911][6] , \mem[911][5] , \mem[911][4] , \mem[911][3] ,
         \mem[911][2] , \mem[911][1] , \mem[911][0] , \mem[910][7] ,
         \mem[910][6] , \mem[910][5] , \mem[910][4] , \mem[910][3] ,
         \mem[910][2] , \mem[910][1] , \mem[910][0] , \mem[909][7] ,
         \mem[909][6] , \mem[909][5] , \mem[909][4] , \mem[909][3] ,
         \mem[909][2] , \mem[909][1] , \mem[909][0] , \mem[908][7] ,
         \mem[908][6] , \mem[908][5] , \mem[908][4] , \mem[908][3] ,
         \mem[908][2] , \mem[908][1] , \mem[908][0] , \mem[907][7] ,
         \mem[907][6] , \mem[907][5] , \mem[907][4] , \mem[907][3] ,
         \mem[907][2] , \mem[907][1] , \mem[907][0] , \mem[906][7] ,
         \mem[906][6] , \mem[906][5] , \mem[906][4] , \mem[906][3] ,
         \mem[906][2] , \mem[906][1] , \mem[906][0] , \mem[905][7] ,
         \mem[905][6] , \mem[905][5] , \mem[905][4] , \mem[905][3] ,
         \mem[905][2] , \mem[905][1] , \mem[905][0] , \mem[904][7] ,
         \mem[904][6] , \mem[904][5] , \mem[904][4] , \mem[904][3] ,
         \mem[904][2] , \mem[904][1] , \mem[904][0] , \mem[903][7] ,
         \mem[903][6] , \mem[903][5] , \mem[903][4] , \mem[903][3] ,
         \mem[903][2] , \mem[903][1] , \mem[903][0] , \mem[902][7] ,
         \mem[902][6] , \mem[902][5] , \mem[902][4] , \mem[902][3] ,
         \mem[902][2] , \mem[902][1] , \mem[902][0] , \mem[901][7] ,
         \mem[901][6] , \mem[901][5] , \mem[901][4] , \mem[901][3] ,
         \mem[901][2] , \mem[901][1] , \mem[901][0] , \mem[900][7] ,
         \mem[900][6] , \mem[900][5] , \mem[900][4] , \mem[900][3] ,
         \mem[900][2] , \mem[900][1] , \mem[900][0] , \mem[899][7] ,
         \mem[899][6] , \mem[899][5] , \mem[899][4] , \mem[899][3] ,
         \mem[899][2] , \mem[899][1] , \mem[899][0] , \mem[898][7] ,
         \mem[898][6] , \mem[898][5] , \mem[898][4] , \mem[898][3] ,
         \mem[898][2] , \mem[898][1] , \mem[898][0] , \mem[897][7] ,
         \mem[897][6] , \mem[897][5] , \mem[897][4] , \mem[897][3] ,
         \mem[897][2] , \mem[897][1] , \mem[897][0] , \mem[896][7] ,
         \mem[896][6] , \mem[896][5] , \mem[896][4] , \mem[896][3] ,
         \mem[896][2] , \mem[896][1] , \mem[896][0] , \mem[895][7] ,
         \mem[895][6] , \mem[895][5] , \mem[895][4] , \mem[895][3] ,
         \mem[895][2] , \mem[895][1] , \mem[895][0] , \mem[894][7] ,
         \mem[894][6] , \mem[894][5] , \mem[894][4] , \mem[894][3] ,
         \mem[894][2] , \mem[894][1] , \mem[894][0] , \mem[893][7] ,
         \mem[893][6] , \mem[893][5] , \mem[893][4] , \mem[893][3] ,
         \mem[893][2] , \mem[893][1] , \mem[893][0] , \mem[892][7] ,
         \mem[892][6] , \mem[892][5] , \mem[892][4] , \mem[892][3] ,
         \mem[892][2] , \mem[892][1] , \mem[892][0] , \mem[891][7] ,
         \mem[891][6] , \mem[891][5] , \mem[891][4] , \mem[891][3] ,
         \mem[891][2] , \mem[891][1] , \mem[891][0] , \mem[890][7] ,
         \mem[890][6] , \mem[890][5] , \mem[890][4] , \mem[890][3] ,
         \mem[890][2] , \mem[890][1] , \mem[890][0] , \mem[889][7] ,
         \mem[889][6] , \mem[889][5] , \mem[889][4] , \mem[889][3] ,
         \mem[889][2] , \mem[889][1] , \mem[889][0] , \mem[888][7] ,
         \mem[888][6] , \mem[888][5] , \mem[888][4] , \mem[888][3] ,
         \mem[888][2] , \mem[888][1] , \mem[888][0] , \mem[887][7] ,
         \mem[887][6] , \mem[887][5] , \mem[887][4] , \mem[887][3] ,
         \mem[887][2] , \mem[887][1] , \mem[887][0] , \mem[886][7] ,
         \mem[886][6] , \mem[886][5] , \mem[886][4] , \mem[886][3] ,
         \mem[886][2] , \mem[886][1] , \mem[886][0] , \mem[885][7] ,
         \mem[885][6] , \mem[885][5] , \mem[885][4] , \mem[885][3] ,
         \mem[885][2] , \mem[885][1] , \mem[885][0] , \mem[884][7] ,
         \mem[884][6] , \mem[884][5] , \mem[884][4] , \mem[884][3] ,
         \mem[884][2] , \mem[884][1] , \mem[884][0] , \mem[883][7] ,
         \mem[883][6] , \mem[883][5] , \mem[883][4] , \mem[883][3] ,
         \mem[883][2] , \mem[883][1] , \mem[883][0] , \mem[882][7] ,
         \mem[882][6] , \mem[882][5] , \mem[882][4] , \mem[882][3] ,
         \mem[882][2] , \mem[882][1] , \mem[882][0] , \mem[881][7] ,
         \mem[881][6] , \mem[881][5] , \mem[881][4] , \mem[881][3] ,
         \mem[881][2] , \mem[881][1] , \mem[881][0] , \mem[880][7] ,
         \mem[880][6] , \mem[880][5] , \mem[880][4] , \mem[880][3] ,
         \mem[880][2] , \mem[880][1] , \mem[880][0] , \mem[879][7] ,
         \mem[879][6] , \mem[879][5] , \mem[879][4] , \mem[879][3] ,
         \mem[879][2] , \mem[879][1] , \mem[879][0] , \mem[878][7] ,
         \mem[878][6] , \mem[878][5] , \mem[878][4] , \mem[878][3] ,
         \mem[878][2] , \mem[878][1] , \mem[878][0] , \mem[877][7] ,
         \mem[877][6] , \mem[877][5] , \mem[877][4] , \mem[877][3] ,
         \mem[877][2] , \mem[877][1] , \mem[877][0] , \mem[876][7] ,
         \mem[876][6] , \mem[876][5] , \mem[876][4] , \mem[876][3] ,
         \mem[876][2] , \mem[876][1] , \mem[876][0] , \mem[875][7] ,
         \mem[875][6] , \mem[875][5] , \mem[875][4] , \mem[875][3] ,
         \mem[875][2] , \mem[875][1] , \mem[875][0] , \mem[874][7] ,
         \mem[874][6] , \mem[874][5] , \mem[874][4] , \mem[874][3] ,
         \mem[874][2] , \mem[874][1] , \mem[874][0] , \mem[873][7] ,
         \mem[873][6] , \mem[873][5] , \mem[873][4] , \mem[873][3] ,
         \mem[873][2] , \mem[873][1] , \mem[873][0] , \mem[872][7] ,
         \mem[872][6] , \mem[872][5] , \mem[872][4] , \mem[872][3] ,
         \mem[872][2] , \mem[872][1] , \mem[872][0] , \mem[871][7] ,
         \mem[871][6] , \mem[871][5] , \mem[871][4] , \mem[871][3] ,
         \mem[871][2] , \mem[871][1] , \mem[871][0] , \mem[870][7] ,
         \mem[870][6] , \mem[870][5] , \mem[870][4] , \mem[870][3] ,
         \mem[870][2] , \mem[870][1] , \mem[870][0] , \mem[869][7] ,
         \mem[869][6] , \mem[869][5] , \mem[869][4] , \mem[869][3] ,
         \mem[869][2] , \mem[869][1] , \mem[869][0] , \mem[868][7] ,
         \mem[868][6] , \mem[868][5] , \mem[868][4] , \mem[868][3] ,
         \mem[868][2] , \mem[868][1] , \mem[868][0] , \mem[867][7] ,
         \mem[867][6] , \mem[867][5] , \mem[867][4] , \mem[867][3] ,
         \mem[867][2] , \mem[867][1] , \mem[867][0] , \mem[866][7] ,
         \mem[866][6] , \mem[866][5] , \mem[866][4] , \mem[866][3] ,
         \mem[866][2] , \mem[866][1] , \mem[866][0] , \mem[865][7] ,
         \mem[865][6] , \mem[865][5] , \mem[865][4] , \mem[865][3] ,
         \mem[865][2] , \mem[865][1] , \mem[865][0] , \mem[864][7] ,
         \mem[864][6] , \mem[864][5] , \mem[864][4] , \mem[864][3] ,
         \mem[864][2] , \mem[864][1] , \mem[864][0] , \mem[863][7] ,
         \mem[863][6] , \mem[863][5] , \mem[863][4] , \mem[863][3] ,
         \mem[863][2] , \mem[863][1] , \mem[863][0] , \mem[862][7] ,
         \mem[862][6] , \mem[862][5] , \mem[862][4] , \mem[862][3] ,
         \mem[862][2] , \mem[862][1] , \mem[862][0] , \mem[861][7] ,
         \mem[861][6] , \mem[861][5] , \mem[861][4] , \mem[861][3] ,
         \mem[861][2] , \mem[861][1] , \mem[861][0] , \mem[860][7] ,
         \mem[860][6] , \mem[860][5] , \mem[860][4] , \mem[860][3] ,
         \mem[860][2] , \mem[860][1] , \mem[860][0] , \mem[859][7] ,
         \mem[859][6] , \mem[859][5] , \mem[859][4] , \mem[859][3] ,
         \mem[859][2] , \mem[859][1] , \mem[859][0] , \mem[858][7] ,
         \mem[858][6] , \mem[858][5] , \mem[858][4] , \mem[858][3] ,
         \mem[858][2] , \mem[858][1] , \mem[858][0] , \mem[857][7] ,
         \mem[857][6] , \mem[857][5] , \mem[857][4] , \mem[857][3] ,
         \mem[857][2] , \mem[857][1] , \mem[857][0] , \mem[856][7] ,
         \mem[856][6] , \mem[856][5] , \mem[856][4] , \mem[856][3] ,
         \mem[856][2] , \mem[856][1] , \mem[856][0] , \mem[855][7] ,
         \mem[855][6] , \mem[855][5] , \mem[855][4] , \mem[855][3] ,
         \mem[855][2] , \mem[855][1] , \mem[855][0] , \mem[854][7] ,
         \mem[854][6] , \mem[854][5] , \mem[854][4] , \mem[854][3] ,
         \mem[854][2] , \mem[854][1] , \mem[854][0] , \mem[853][7] ,
         \mem[853][6] , \mem[853][5] , \mem[853][4] , \mem[853][3] ,
         \mem[853][2] , \mem[853][1] , \mem[853][0] , \mem[852][7] ,
         \mem[852][6] , \mem[852][5] , \mem[852][4] , \mem[852][3] ,
         \mem[852][2] , \mem[852][1] , \mem[852][0] , \mem[851][7] ,
         \mem[851][6] , \mem[851][5] , \mem[851][4] , \mem[851][3] ,
         \mem[851][2] , \mem[851][1] , \mem[851][0] , \mem[850][7] ,
         \mem[850][6] , \mem[850][5] , \mem[850][4] , \mem[850][3] ,
         \mem[850][2] , \mem[850][1] , \mem[850][0] , \mem[849][7] ,
         \mem[849][6] , \mem[849][5] , \mem[849][4] , \mem[849][3] ,
         \mem[849][2] , \mem[849][1] , \mem[849][0] , \mem[848][7] ,
         \mem[848][6] , \mem[848][5] , \mem[848][4] , \mem[848][3] ,
         \mem[848][2] , \mem[848][1] , \mem[848][0] , \mem[847][7] ,
         \mem[847][6] , \mem[847][5] , \mem[847][4] , \mem[847][3] ,
         \mem[847][2] , \mem[847][1] , \mem[847][0] , \mem[846][7] ,
         \mem[846][6] , \mem[846][5] , \mem[846][4] , \mem[846][3] ,
         \mem[846][2] , \mem[846][1] , \mem[846][0] , \mem[845][7] ,
         \mem[845][6] , \mem[845][5] , \mem[845][4] , \mem[845][3] ,
         \mem[845][2] , \mem[845][1] , \mem[845][0] , \mem[844][7] ,
         \mem[844][6] , \mem[844][5] , \mem[844][4] , \mem[844][3] ,
         \mem[844][2] , \mem[844][1] , \mem[844][0] , \mem[843][7] ,
         \mem[843][6] , \mem[843][5] , \mem[843][4] , \mem[843][3] ,
         \mem[843][2] , \mem[843][1] , \mem[843][0] , \mem[842][7] ,
         \mem[842][6] , \mem[842][5] , \mem[842][4] , \mem[842][3] ,
         \mem[842][2] , \mem[842][1] , \mem[842][0] , \mem[841][7] ,
         \mem[841][6] , \mem[841][5] , \mem[841][4] , \mem[841][3] ,
         \mem[841][2] , \mem[841][1] , \mem[841][0] , \mem[840][7] ,
         \mem[840][6] , \mem[840][5] , \mem[840][4] , \mem[840][3] ,
         \mem[840][2] , \mem[840][1] , \mem[840][0] , \mem[839][7] ,
         \mem[839][6] , \mem[839][5] , \mem[839][4] , \mem[839][3] ,
         \mem[839][2] , \mem[839][1] , \mem[839][0] , \mem[838][7] ,
         \mem[838][6] , \mem[838][5] , \mem[838][4] , \mem[838][3] ,
         \mem[838][2] , \mem[838][1] , \mem[838][0] , \mem[837][7] ,
         \mem[837][6] , \mem[837][5] , \mem[837][4] , \mem[837][3] ,
         \mem[837][2] , \mem[837][1] , \mem[837][0] , \mem[836][7] ,
         \mem[836][6] , \mem[836][5] , \mem[836][4] , \mem[836][3] ,
         \mem[836][2] , \mem[836][1] , \mem[836][0] , \mem[835][7] ,
         \mem[835][6] , \mem[835][5] , \mem[835][4] , \mem[835][3] ,
         \mem[835][2] , \mem[835][1] , \mem[835][0] , \mem[834][7] ,
         \mem[834][6] , \mem[834][5] , \mem[834][4] , \mem[834][3] ,
         \mem[834][2] , \mem[834][1] , \mem[834][0] , \mem[833][7] ,
         \mem[833][6] , \mem[833][5] , \mem[833][4] , \mem[833][3] ,
         \mem[833][2] , \mem[833][1] , \mem[833][0] , \mem[832][7] ,
         \mem[832][6] , \mem[832][5] , \mem[832][4] , \mem[832][3] ,
         \mem[832][2] , \mem[832][1] , \mem[832][0] , \mem[831][7] ,
         \mem[831][6] , \mem[831][5] , \mem[831][4] , \mem[831][3] ,
         \mem[831][2] , \mem[831][1] , \mem[831][0] , \mem[830][7] ,
         \mem[830][6] , \mem[830][5] , \mem[830][4] , \mem[830][3] ,
         \mem[830][2] , \mem[830][1] , \mem[830][0] , \mem[829][7] ,
         \mem[829][6] , \mem[829][5] , \mem[829][4] , \mem[829][3] ,
         \mem[829][2] , \mem[829][1] , \mem[829][0] , \mem[828][7] ,
         \mem[828][6] , \mem[828][5] , \mem[828][4] , \mem[828][3] ,
         \mem[828][2] , \mem[828][1] , \mem[828][0] , \mem[827][7] ,
         \mem[827][6] , \mem[827][5] , \mem[827][4] , \mem[827][3] ,
         \mem[827][2] , \mem[827][1] , \mem[827][0] , \mem[826][7] ,
         \mem[826][6] , \mem[826][5] , \mem[826][4] , \mem[826][3] ,
         \mem[826][2] , \mem[826][1] , \mem[826][0] , \mem[825][7] ,
         \mem[825][6] , \mem[825][5] , \mem[825][4] , \mem[825][3] ,
         \mem[825][2] , \mem[825][1] , \mem[825][0] , \mem[824][7] ,
         \mem[824][6] , \mem[824][5] , \mem[824][4] , \mem[824][3] ,
         \mem[824][2] , \mem[824][1] , \mem[824][0] , \mem[823][7] ,
         \mem[823][6] , \mem[823][5] , \mem[823][4] , \mem[823][3] ,
         \mem[823][2] , \mem[823][1] , \mem[823][0] , \mem[822][7] ,
         \mem[822][6] , \mem[822][5] , \mem[822][4] , \mem[822][3] ,
         \mem[822][2] , \mem[822][1] , \mem[822][0] , \mem[821][7] ,
         \mem[821][6] , \mem[821][5] , \mem[821][4] , \mem[821][3] ,
         \mem[821][2] , \mem[821][1] , \mem[821][0] , \mem[820][7] ,
         \mem[820][6] , \mem[820][5] , \mem[820][4] , \mem[820][3] ,
         \mem[820][2] , \mem[820][1] , \mem[820][0] , \mem[819][7] ,
         \mem[819][6] , \mem[819][5] , \mem[819][4] , \mem[819][3] ,
         \mem[819][2] , \mem[819][1] , \mem[819][0] , \mem[818][7] ,
         \mem[818][6] , \mem[818][5] , \mem[818][4] , \mem[818][3] ,
         \mem[818][2] , \mem[818][1] , \mem[818][0] , \mem[817][7] ,
         \mem[817][6] , \mem[817][5] , \mem[817][4] , \mem[817][3] ,
         \mem[817][2] , \mem[817][1] , \mem[817][0] , \mem[816][7] ,
         \mem[816][6] , \mem[816][5] , \mem[816][4] , \mem[816][3] ,
         \mem[816][2] , \mem[816][1] , \mem[816][0] , \mem[815][7] ,
         \mem[815][6] , \mem[815][5] , \mem[815][4] , \mem[815][3] ,
         \mem[815][2] , \mem[815][1] , \mem[815][0] , \mem[814][7] ,
         \mem[814][6] , \mem[814][5] , \mem[814][4] , \mem[814][3] ,
         \mem[814][2] , \mem[814][1] , \mem[814][0] , \mem[813][7] ,
         \mem[813][6] , \mem[813][5] , \mem[813][4] , \mem[813][3] ,
         \mem[813][2] , \mem[813][1] , \mem[813][0] , \mem[812][7] ,
         \mem[812][6] , \mem[812][5] , \mem[812][4] , \mem[812][3] ,
         \mem[812][2] , \mem[812][1] , \mem[812][0] , \mem[811][7] ,
         \mem[811][6] , \mem[811][5] , \mem[811][4] , \mem[811][3] ,
         \mem[811][2] , \mem[811][1] , \mem[811][0] , \mem[810][7] ,
         \mem[810][6] , \mem[810][5] , \mem[810][4] , \mem[810][3] ,
         \mem[810][2] , \mem[810][1] , \mem[810][0] , \mem[809][7] ,
         \mem[809][6] , \mem[809][5] , \mem[809][4] , \mem[809][3] ,
         \mem[809][2] , \mem[809][1] , \mem[809][0] , \mem[808][7] ,
         \mem[808][6] , \mem[808][5] , \mem[808][4] , \mem[808][3] ,
         \mem[808][2] , \mem[808][1] , \mem[808][0] , \mem[807][7] ,
         \mem[807][6] , \mem[807][5] , \mem[807][4] , \mem[807][3] ,
         \mem[807][2] , \mem[807][1] , \mem[807][0] , \mem[806][7] ,
         \mem[806][6] , \mem[806][5] , \mem[806][4] , \mem[806][3] ,
         \mem[806][2] , \mem[806][1] , \mem[806][0] , \mem[805][7] ,
         \mem[805][6] , \mem[805][5] , \mem[805][4] , \mem[805][3] ,
         \mem[805][2] , \mem[805][1] , \mem[805][0] , \mem[804][7] ,
         \mem[804][6] , \mem[804][5] , \mem[804][4] , \mem[804][3] ,
         \mem[804][2] , \mem[804][1] , \mem[804][0] , \mem[803][7] ,
         \mem[803][6] , \mem[803][5] , \mem[803][4] , \mem[803][3] ,
         \mem[803][2] , \mem[803][1] , \mem[803][0] , \mem[802][7] ,
         \mem[802][6] , \mem[802][5] , \mem[802][4] , \mem[802][3] ,
         \mem[802][2] , \mem[802][1] , \mem[802][0] , \mem[801][7] ,
         \mem[801][6] , \mem[801][5] , \mem[801][4] , \mem[801][3] ,
         \mem[801][2] , \mem[801][1] , \mem[801][0] , \mem[800][7] ,
         \mem[800][6] , \mem[800][5] , \mem[800][4] , \mem[800][3] ,
         \mem[800][2] , \mem[800][1] , \mem[800][0] , \mem[799][7] ,
         \mem[799][6] , \mem[799][5] , \mem[799][4] , \mem[799][3] ,
         \mem[799][2] , \mem[799][1] , \mem[799][0] , \mem[798][7] ,
         \mem[798][6] , \mem[798][5] , \mem[798][4] , \mem[798][3] ,
         \mem[798][2] , \mem[798][1] , \mem[798][0] , \mem[797][7] ,
         \mem[797][6] , \mem[797][5] , \mem[797][4] , \mem[797][3] ,
         \mem[797][2] , \mem[797][1] , \mem[797][0] , \mem[796][7] ,
         \mem[796][6] , \mem[796][5] , \mem[796][4] , \mem[796][3] ,
         \mem[796][2] , \mem[796][1] , \mem[796][0] , \mem[795][7] ,
         \mem[795][6] , \mem[795][5] , \mem[795][4] , \mem[795][3] ,
         \mem[795][2] , \mem[795][1] , \mem[795][0] , \mem[794][7] ,
         \mem[794][6] , \mem[794][5] , \mem[794][4] , \mem[794][3] ,
         \mem[794][2] , \mem[794][1] , \mem[794][0] , \mem[793][7] ,
         \mem[793][6] , \mem[793][5] , \mem[793][4] , \mem[793][3] ,
         \mem[793][2] , \mem[793][1] , \mem[793][0] , \mem[792][7] ,
         \mem[792][6] , \mem[792][5] , \mem[792][4] , \mem[792][3] ,
         \mem[792][2] , \mem[792][1] , \mem[792][0] , \mem[791][7] ,
         \mem[791][6] , \mem[791][5] , \mem[791][4] , \mem[791][3] ,
         \mem[791][2] , \mem[791][1] , \mem[791][0] , \mem[790][7] ,
         \mem[790][6] , \mem[790][5] , \mem[790][4] , \mem[790][3] ,
         \mem[790][2] , \mem[790][1] , \mem[790][0] , \mem[789][7] ,
         \mem[789][6] , \mem[789][5] , \mem[789][4] , \mem[789][3] ,
         \mem[789][2] , \mem[789][1] , \mem[789][0] , \mem[788][7] ,
         \mem[788][6] , \mem[788][5] , \mem[788][4] , \mem[788][3] ,
         \mem[788][2] , \mem[788][1] , \mem[788][0] , \mem[787][7] ,
         \mem[787][6] , \mem[787][5] , \mem[787][4] , \mem[787][3] ,
         \mem[787][2] , \mem[787][1] , \mem[787][0] , \mem[786][7] ,
         \mem[786][6] , \mem[786][5] , \mem[786][4] , \mem[786][3] ,
         \mem[786][2] , \mem[786][1] , \mem[786][0] , \mem[785][7] ,
         \mem[785][6] , \mem[785][5] , \mem[785][4] , \mem[785][3] ,
         \mem[785][2] , \mem[785][1] , \mem[785][0] , \mem[784][7] ,
         \mem[784][6] , \mem[784][5] , \mem[784][4] , \mem[784][3] ,
         \mem[784][2] , \mem[784][1] , \mem[784][0] , \mem[783][7] ,
         \mem[783][6] , \mem[783][5] , \mem[783][4] , \mem[783][3] ,
         \mem[783][2] , \mem[783][1] , \mem[783][0] , \mem[782][7] ,
         \mem[782][6] , \mem[782][5] , \mem[782][4] , \mem[782][3] ,
         \mem[782][2] , \mem[782][1] , \mem[782][0] , \mem[781][7] ,
         \mem[781][6] , \mem[781][5] , \mem[781][4] , \mem[781][3] ,
         \mem[781][2] , \mem[781][1] , \mem[781][0] , \mem[780][7] ,
         \mem[780][6] , \mem[780][5] , \mem[780][4] , \mem[780][3] ,
         \mem[780][2] , \mem[780][1] , \mem[780][0] , \mem[779][7] ,
         \mem[779][6] , \mem[779][5] , \mem[779][4] , \mem[779][3] ,
         \mem[779][2] , \mem[779][1] , \mem[779][0] , \mem[778][7] ,
         \mem[778][6] , \mem[778][5] , \mem[778][4] , \mem[778][3] ,
         \mem[778][2] , \mem[778][1] , \mem[778][0] , \mem[777][7] ,
         \mem[777][6] , \mem[777][5] , \mem[777][4] , \mem[777][3] ,
         \mem[777][2] , \mem[777][1] , \mem[777][0] , \mem[776][7] ,
         \mem[776][6] , \mem[776][5] , \mem[776][4] , \mem[776][3] ,
         \mem[776][2] , \mem[776][1] , \mem[776][0] , \mem[775][7] ,
         \mem[775][6] , \mem[775][5] , \mem[775][4] , \mem[775][3] ,
         \mem[775][2] , \mem[775][1] , \mem[775][0] , \mem[774][7] ,
         \mem[774][6] , \mem[774][5] , \mem[774][4] , \mem[774][3] ,
         \mem[774][2] , \mem[774][1] , \mem[774][0] , \mem[773][7] ,
         \mem[773][6] , \mem[773][5] , \mem[773][4] , \mem[773][3] ,
         \mem[773][2] , \mem[773][1] , \mem[773][0] , \mem[772][7] ,
         \mem[772][6] , \mem[772][5] , \mem[772][4] , \mem[772][3] ,
         \mem[772][2] , \mem[772][1] , \mem[772][0] , \mem[771][7] ,
         \mem[771][6] , \mem[771][5] , \mem[771][4] , \mem[771][3] ,
         \mem[771][2] , \mem[771][1] , \mem[771][0] , \mem[770][7] ,
         \mem[770][6] , \mem[770][5] , \mem[770][4] , \mem[770][3] ,
         \mem[770][2] , \mem[770][1] , \mem[770][0] , \mem[769][7] ,
         \mem[769][6] , \mem[769][5] , \mem[769][4] , \mem[769][3] ,
         \mem[769][2] , \mem[769][1] , \mem[769][0] , \mem[768][7] ,
         \mem[768][6] , \mem[768][5] , \mem[768][4] , \mem[768][3] ,
         \mem[768][2] , \mem[768][1] , \mem[768][0] , \mem[767][7] ,
         \mem[767][6] , \mem[767][5] , \mem[767][4] , \mem[767][3] ,
         \mem[767][2] , \mem[767][1] , \mem[767][0] , \mem[766][7] ,
         \mem[766][6] , \mem[766][5] , \mem[766][4] , \mem[766][3] ,
         \mem[766][2] , \mem[766][1] , \mem[766][0] , \mem[765][7] ,
         \mem[765][6] , \mem[765][5] , \mem[765][4] , \mem[765][3] ,
         \mem[765][2] , \mem[765][1] , \mem[765][0] , \mem[764][7] ,
         \mem[764][6] , \mem[764][5] , \mem[764][4] , \mem[764][3] ,
         \mem[764][2] , \mem[764][1] , \mem[764][0] , \mem[763][7] ,
         \mem[763][6] , \mem[763][5] , \mem[763][4] , \mem[763][3] ,
         \mem[763][2] , \mem[763][1] , \mem[763][0] , \mem[762][7] ,
         \mem[762][6] , \mem[762][5] , \mem[762][4] , \mem[762][3] ,
         \mem[762][2] , \mem[762][1] , \mem[762][0] , \mem[761][7] ,
         \mem[761][6] , \mem[761][5] , \mem[761][4] , \mem[761][3] ,
         \mem[761][2] , \mem[761][1] , \mem[761][0] , \mem[760][7] ,
         \mem[760][6] , \mem[760][5] , \mem[760][4] , \mem[760][3] ,
         \mem[760][2] , \mem[760][1] , \mem[760][0] , \mem[759][7] ,
         \mem[759][6] , \mem[759][5] , \mem[759][4] , \mem[759][3] ,
         \mem[759][2] , \mem[759][1] , \mem[759][0] , \mem[758][7] ,
         \mem[758][6] , \mem[758][5] , \mem[758][4] , \mem[758][3] ,
         \mem[758][2] , \mem[758][1] , \mem[758][0] , \mem[757][7] ,
         \mem[757][6] , \mem[757][5] , \mem[757][4] , \mem[757][3] ,
         \mem[757][2] , \mem[757][1] , \mem[757][0] , \mem[756][7] ,
         \mem[756][6] , \mem[756][5] , \mem[756][4] , \mem[756][3] ,
         \mem[756][2] , \mem[756][1] , \mem[756][0] , \mem[755][7] ,
         \mem[755][6] , \mem[755][5] , \mem[755][4] , \mem[755][3] ,
         \mem[755][2] , \mem[755][1] , \mem[755][0] , \mem[754][7] ,
         \mem[754][6] , \mem[754][5] , \mem[754][4] , \mem[754][3] ,
         \mem[754][2] , \mem[754][1] , \mem[754][0] , \mem[753][7] ,
         \mem[753][6] , \mem[753][5] , \mem[753][4] , \mem[753][3] ,
         \mem[753][2] , \mem[753][1] , \mem[753][0] , \mem[752][7] ,
         \mem[752][6] , \mem[752][5] , \mem[752][4] , \mem[752][3] ,
         \mem[752][2] , \mem[752][1] , \mem[752][0] , \mem[751][7] ,
         \mem[751][6] , \mem[751][5] , \mem[751][4] , \mem[751][3] ,
         \mem[751][2] , \mem[751][1] , \mem[751][0] , \mem[750][7] ,
         \mem[750][6] , \mem[750][5] , \mem[750][4] , \mem[750][3] ,
         \mem[750][2] , \mem[750][1] , \mem[750][0] , \mem[749][7] ,
         \mem[749][6] , \mem[749][5] , \mem[749][4] , \mem[749][3] ,
         \mem[749][2] , \mem[749][1] , \mem[749][0] , \mem[748][7] ,
         \mem[748][6] , \mem[748][5] , \mem[748][4] , \mem[748][3] ,
         \mem[748][2] , \mem[748][1] , \mem[748][0] , \mem[747][7] ,
         \mem[747][6] , \mem[747][5] , \mem[747][4] , \mem[747][3] ,
         \mem[747][2] , \mem[747][1] , \mem[747][0] , \mem[746][7] ,
         \mem[746][6] , \mem[746][5] , \mem[746][4] , \mem[746][3] ,
         \mem[746][2] , \mem[746][1] , \mem[746][0] , \mem[745][7] ,
         \mem[745][6] , \mem[745][5] , \mem[745][4] , \mem[745][3] ,
         \mem[745][2] , \mem[745][1] , \mem[745][0] , \mem[744][7] ,
         \mem[744][6] , \mem[744][5] , \mem[744][4] , \mem[744][3] ,
         \mem[744][2] , \mem[744][1] , \mem[744][0] , \mem[743][7] ,
         \mem[743][6] , \mem[743][5] , \mem[743][4] , \mem[743][3] ,
         \mem[743][2] , \mem[743][1] , \mem[743][0] , \mem[742][7] ,
         \mem[742][6] , \mem[742][5] , \mem[742][4] , \mem[742][3] ,
         \mem[742][2] , \mem[742][1] , \mem[742][0] , \mem[741][7] ,
         \mem[741][6] , \mem[741][5] , \mem[741][4] , \mem[741][3] ,
         \mem[741][2] , \mem[741][1] , \mem[741][0] , \mem[740][7] ,
         \mem[740][6] , \mem[740][5] , \mem[740][4] , \mem[740][3] ,
         \mem[740][2] , \mem[740][1] , \mem[740][0] , \mem[739][7] ,
         \mem[739][6] , \mem[739][5] , \mem[739][4] , \mem[739][3] ,
         \mem[739][2] , \mem[739][1] , \mem[739][0] , \mem[738][7] ,
         \mem[738][6] , \mem[738][5] , \mem[738][4] , \mem[738][3] ,
         \mem[738][2] , \mem[738][1] , \mem[738][0] , \mem[737][7] ,
         \mem[737][6] , \mem[737][5] , \mem[737][4] , \mem[737][3] ,
         \mem[737][2] , \mem[737][1] , \mem[737][0] , \mem[736][7] ,
         \mem[736][6] , \mem[736][5] , \mem[736][4] , \mem[736][3] ,
         \mem[736][2] , \mem[736][1] , \mem[736][0] , \mem[735][7] ,
         \mem[735][6] , \mem[735][5] , \mem[735][4] , \mem[735][3] ,
         \mem[735][2] , \mem[735][1] , \mem[735][0] , \mem[734][7] ,
         \mem[734][6] , \mem[734][5] , \mem[734][4] , \mem[734][3] ,
         \mem[734][2] , \mem[734][1] , \mem[734][0] , \mem[733][7] ,
         \mem[733][6] , \mem[733][5] , \mem[733][4] , \mem[733][3] ,
         \mem[733][2] , \mem[733][1] , \mem[733][0] , \mem[732][7] ,
         \mem[732][6] , \mem[732][5] , \mem[732][4] , \mem[732][3] ,
         \mem[732][2] , \mem[732][1] , \mem[732][0] , \mem[731][7] ,
         \mem[731][6] , \mem[731][5] , \mem[731][4] , \mem[731][3] ,
         \mem[731][2] , \mem[731][1] , \mem[731][0] , \mem[730][7] ,
         \mem[730][6] , \mem[730][5] , \mem[730][4] , \mem[730][3] ,
         \mem[730][2] , \mem[730][1] , \mem[730][0] , \mem[729][7] ,
         \mem[729][6] , \mem[729][5] , \mem[729][4] , \mem[729][3] ,
         \mem[729][2] , \mem[729][1] , \mem[729][0] , \mem[728][7] ,
         \mem[728][6] , \mem[728][5] , \mem[728][4] , \mem[728][3] ,
         \mem[728][2] , \mem[728][1] , \mem[728][0] , \mem[727][7] ,
         \mem[727][6] , \mem[727][5] , \mem[727][4] , \mem[727][3] ,
         \mem[727][2] , \mem[727][1] , \mem[727][0] , \mem[726][7] ,
         \mem[726][6] , \mem[726][5] , \mem[726][4] , \mem[726][3] ,
         \mem[726][2] , \mem[726][1] , \mem[726][0] , \mem[725][7] ,
         \mem[725][6] , \mem[725][5] , \mem[725][4] , \mem[725][3] ,
         \mem[725][2] , \mem[725][1] , \mem[725][0] , \mem[724][7] ,
         \mem[724][6] , \mem[724][5] , \mem[724][4] , \mem[724][3] ,
         \mem[724][2] , \mem[724][1] , \mem[724][0] , \mem[723][7] ,
         \mem[723][6] , \mem[723][5] , \mem[723][4] , \mem[723][3] ,
         \mem[723][2] , \mem[723][1] , \mem[723][0] , \mem[722][7] ,
         \mem[722][6] , \mem[722][5] , \mem[722][4] , \mem[722][3] ,
         \mem[722][2] , \mem[722][1] , \mem[722][0] , \mem[721][7] ,
         \mem[721][6] , \mem[721][5] , \mem[721][4] , \mem[721][3] ,
         \mem[721][2] , \mem[721][1] , \mem[721][0] , \mem[720][7] ,
         \mem[720][6] , \mem[720][5] , \mem[720][4] , \mem[720][3] ,
         \mem[720][2] , \mem[720][1] , \mem[720][0] , \mem[719][7] ,
         \mem[719][6] , \mem[719][5] , \mem[719][4] , \mem[719][3] ,
         \mem[719][2] , \mem[719][1] , \mem[719][0] , \mem[718][7] ,
         \mem[718][6] , \mem[718][5] , \mem[718][4] , \mem[718][3] ,
         \mem[718][2] , \mem[718][1] , \mem[718][0] , \mem[717][7] ,
         \mem[717][6] , \mem[717][5] , \mem[717][4] , \mem[717][3] ,
         \mem[717][2] , \mem[717][1] , \mem[717][0] , \mem[716][7] ,
         \mem[716][6] , \mem[716][5] , \mem[716][4] , \mem[716][3] ,
         \mem[716][2] , \mem[716][1] , \mem[716][0] , \mem[715][7] ,
         \mem[715][6] , \mem[715][5] , \mem[715][4] , \mem[715][3] ,
         \mem[715][2] , \mem[715][1] , \mem[715][0] , \mem[714][7] ,
         \mem[714][6] , \mem[714][5] , \mem[714][4] , \mem[714][3] ,
         \mem[714][2] , \mem[714][1] , \mem[714][0] , \mem[713][7] ,
         \mem[713][6] , \mem[713][5] , \mem[713][4] , \mem[713][3] ,
         \mem[713][2] , \mem[713][1] , \mem[713][0] , \mem[712][7] ,
         \mem[712][6] , \mem[712][5] , \mem[712][4] , \mem[712][3] ,
         \mem[712][2] , \mem[712][1] , \mem[712][0] , \mem[711][7] ,
         \mem[711][6] , \mem[711][5] , \mem[711][4] , \mem[711][3] ,
         \mem[711][2] , \mem[711][1] , \mem[711][0] , \mem[710][7] ,
         \mem[710][6] , \mem[710][5] , \mem[710][4] , \mem[710][3] ,
         \mem[710][2] , \mem[710][1] , \mem[710][0] , \mem[709][7] ,
         \mem[709][6] , \mem[709][5] , \mem[709][4] , \mem[709][3] ,
         \mem[709][2] , \mem[709][1] , \mem[709][0] , \mem[708][7] ,
         \mem[708][6] , \mem[708][5] , \mem[708][4] , \mem[708][3] ,
         \mem[708][2] , \mem[708][1] , \mem[708][0] , \mem[707][7] ,
         \mem[707][6] , \mem[707][5] , \mem[707][4] , \mem[707][3] ,
         \mem[707][2] , \mem[707][1] , \mem[707][0] , \mem[706][7] ,
         \mem[706][6] , \mem[706][5] , \mem[706][4] , \mem[706][3] ,
         \mem[706][2] , \mem[706][1] , \mem[706][0] , \mem[705][7] ,
         \mem[705][6] , \mem[705][5] , \mem[705][4] , \mem[705][3] ,
         \mem[705][2] , \mem[705][1] , \mem[705][0] , \mem[704][7] ,
         \mem[704][6] , \mem[704][5] , \mem[704][4] , \mem[704][3] ,
         \mem[704][2] , \mem[704][1] , \mem[704][0] , \mem[703][7] ,
         \mem[703][6] , \mem[703][5] , \mem[703][4] , \mem[703][3] ,
         \mem[703][2] , \mem[703][1] , \mem[703][0] , \mem[702][7] ,
         \mem[702][6] , \mem[702][5] , \mem[702][4] , \mem[702][3] ,
         \mem[702][2] , \mem[702][1] , \mem[702][0] , \mem[701][7] ,
         \mem[701][6] , \mem[701][5] , \mem[701][4] , \mem[701][3] ,
         \mem[701][2] , \mem[701][1] , \mem[701][0] , \mem[700][7] ,
         \mem[700][6] , \mem[700][5] , \mem[700][4] , \mem[700][3] ,
         \mem[700][2] , \mem[700][1] , \mem[700][0] , \mem[699][7] ,
         \mem[699][6] , \mem[699][5] , \mem[699][4] , \mem[699][3] ,
         \mem[699][2] , \mem[699][1] , \mem[699][0] , \mem[698][7] ,
         \mem[698][6] , \mem[698][5] , \mem[698][4] , \mem[698][3] ,
         \mem[698][2] , \mem[698][1] , \mem[698][0] , \mem[697][7] ,
         \mem[697][6] , \mem[697][5] , \mem[697][4] , \mem[697][3] ,
         \mem[697][2] , \mem[697][1] , \mem[697][0] , \mem[696][7] ,
         \mem[696][6] , \mem[696][5] , \mem[696][4] , \mem[696][3] ,
         \mem[696][2] , \mem[696][1] , \mem[696][0] , \mem[695][7] ,
         \mem[695][6] , \mem[695][5] , \mem[695][4] , \mem[695][3] ,
         \mem[695][2] , \mem[695][1] , \mem[695][0] , \mem[694][7] ,
         \mem[694][6] , \mem[694][5] , \mem[694][4] , \mem[694][3] ,
         \mem[694][2] , \mem[694][1] , \mem[694][0] , \mem[693][7] ,
         \mem[693][6] , \mem[693][5] , \mem[693][4] , \mem[693][3] ,
         \mem[693][2] , \mem[693][1] , \mem[693][0] , \mem[692][7] ,
         \mem[692][6] , \mem[692][5] , \mem[692][4] , \mem[692][3] ,
         \mem[692][2] , \mem[692][1] , \mem[692][0] , \mem[691][7] ,
         \mem[691][6] , \mem[691][5] , \mem[691][4] , \mem[691][3] ,
         \mem[691][2] , \mem[691][1] , \mem[691][0] , \mem[690][7] ,
         \mem[690][6] , \mem[690][5] , \mem[690][4] , \mem[690][3] ,
         \mem[690][2] , \mem[690][1] , \mem[690][0] , \mem[689][7] ,
         \mem[689][6] , \mem[689][5] , \mem[689][4] , \mem[689][3] ,
         \mem[689][2] , \mem[689][1] , \mem[689][0] , \mem[688][7] ,
         \mem[688][6] , \mem[688][5] , \mem[688][4] , \mem[688][3] ,
         \mem[688][2] , \mem[688][1] , \mem[688][0] , \mem[687][7] ,
         \mem[687][6] , \mem[687][5] , \mem[687][4] , \mem[687][3] ,
         \mem[687][2] , \mem[687][1] , \mem[687][0] , \mem[686][7] ,
         \mem[686][6] , \mem[686][5] , \mem[686][4] , \mem[686][3] ,
         \mem[686][2] , \mem[686][1] , \mem[686][0] , \mem[685][7] ,
         \mem[685][6] , \mem[685][5] , \mem[685][4] , \mem[685][3] ,
         \mem[685][2] , \mem[685][1] , \mem[685][0] , \mem[684][7] ,
         \mem[684][6] , \mem[684][5] , \mem[684][4] , \mem[684][3] ,
         \mem[684][2] , \mem[684][1] , \mem[684][0] , \mem[683][7] ,
         \mem[683][6] , \mem[683][5] , \mem[683][4] , \mem[683][3] ,
         \mem[683][2] , \mem[683][1] , \mem[683][0] , \mem[682][7] ,
         \mem[682][6] , \mem[682][5] , \mem[682][4] , \mem[682][3] ,
         \mem[682][2] , \mem[682][1] , \mem[682][0] , \mem[681][7] ,
         \mem[681][6] , \mem[681][5] , \mem[681][4] , \mem[681][3] ,
         \mem[681][2] , \mem[681][1] , \mem[681][0] , \mem[680][7] ,
         \mem[680][6] , \mem[680][5] , \mem[680][4] , \mem[680][3] ,
         \mem[680][2] , \mem[680][1] , \mem[680][0] , \mem[679][7] ,
         \mem[679][6] , \mem[679][5] , \mem[679][4] , \mem[679][3] ,
         \mem[679][2] , \mem[679][1] , \mem[679][0] , \mem[678][7] ,
         \mem[678][6] , \mem[678][5] , \mem[678][4] , \mem[678][3] ,
         \mem[678][2] , \mem[678][1] , \mem[678][0] , \mem[677][7] ,
         \mem[677][6] , \mem[677][5] , \mem[677][4] , \mem[677][3] ,
         \mem[677][2] , \mem[677][1] , \mem[677][0] , \mem[676][7] ,
         \mem[676][6] , \mem[676][5] , \mem[676][4] , \mem[676][3] ,
         \mem[676][2] , \mem[676][1] , \mem[676][0] , \mem[675][7] ,
         \mem[675][6] , \mem[675][5] , \mem[675][4] , \mem[675][3] ,
         \mem[675][2] , \mem[675][1] , \mem[675][0] , \mem[674][7] ,
         \mem[674][6] , \mem[674][5] , \mem[674][4] , \mem[674][3] ,
         \mem[674][2] , \mem[674][1] , \mem[674][0] , \mem[673][7] ,
         \mem[673][6] , \mem[673][5] , \mem[673][4] , \mem[673][3] ,
         \mem[673][2] , \mem[673][1] , \mem[673][0] , \mem[672][7] ,
         \mem[672][6] , \mem[672][5] , \mem[672][4] , \mem[672][3] ,
         \mem[672][2] , \mem[672][1] , \mem[672][0] , \mem[671][7] ,
         \mem[671][6] , \mem[671][5] , \mem[671][4] , \mem[671][3] ,
         \mem[671][2] , \mem[671][1] , \mem[671][0] , \mem[670][7] ,
         \mem[670][6] , \mem[670][5] , \mem[670][4] , \mem[670][3] ,
         \mem[670][2] , \mem[670][1] , \mem[670][0] , \mem[669][7] ,
         \mem[669][6] , \mem[669][5] , \mem[669][4] , \mem[669][3] ,
         \mem[669][2] , \mem[669][1] , \mem[669][0] , \mem[668][7] ,
         \mem[668][6] , \mem[668][5] , \mem[668][4] , \mem[668][3] ,
         \mem[668][2] , \mem[668][1] , \mem[668][0] , \mem[667][7] ,
         \mem[667][6] , \mem[667][5] , \mem[667][4] , \mem[667][3] ,
         \mem[667][2] , \mem[667][1] , \mem[667][0] , \mem[666][7] ,
         \mem[666][6] , \mem[666][5] , \mem[666][4] , \mem[666][3] ,
         \mem[666][2] , \mem[666][1] , \mem[666][0] , \mem[665][7] ,
         \mem[665][6] , \mem[665][5] , \mem[665][4] , \mem[665][3] ,
         \mem[665][2] , \mem[665][1] , \mem[665][0] , \mem[664][7] ,
         \mem[664][6] , \mem[664][5] , \mem[664][4] , \mem[664][3] ,
         \mem[664][2] , \mem[664][1] , \mem[664][0] , \mem[663][7] ,
         \mem[663][6] , \mem[663][5] , \mem[663][4] , \mem[663][3] ,
         \mem[663][2] , \mem[663][1] , \mem[663][0] , \mem[662][7] ,
         \mem[662][6] , \mem[662][5] , \mem[662][4] , \mem[662][3] ,
         \mem[662][2] , \mem[662][1] , \mem[662][0] , \mem[661][7] ,
         \mem[661][6] , \mem[661][5] , \mem[661][4] , \mem[661][3] ,
         \mem[661][2] , \mem[661][1] , \mem[661][0] , \mem[660][7] ,
         \mem[660][6] , \mem[660][5] , \mem[660][4] , \mem[660][3] ,
         \mem[660][2] , \mem[660][1] , \mem[660][0] , \mem[659][7] ,
         \mem[659][6] , \mem[659][5] , \mem[659][4] , \mem[659][3] ,
         \mem[659][2] , \mem[659][1] , \mem[659][0] , \mem[658][7] ,
         \mem[658][6] , \mem[658][5] , \mem[658][4] , \mem[658][3] ,
         \mem[658][2] , \mem[658][1] , \mem[658][0] , \mem[657][7] ,
         \mem[657][6] , \mem[657][5] , \mem[657][4] , \mem[657][3] ,
         \mem[657][2] , \mem[657][1] , \mem[657][0] , \mem[656][7] ,
         \mem[656][6] , \mem[656][5] , \mem[656][4] , \mem[656][3] ,
         \mem[656][2] , \mem[656][1] , \mem[656][0] , \mem[655][7] ,
         \mem[655][6] , \mem[655][5] , \mem[655][4] , \mem[655][3] ,
         \mem[655][2] , \mem[655][1] , \mem[655][0] , \mem[654][7] ,
         \mem[654][6] , \mem[654][5] , \mem[654][4] , \mem[654][3] ,
         \mem[654][2] , \mem[654][1] , \mem[654][0] , \mem[653][7] ,
         \mem[653][6] , \mem[653][5] , \mem[653][4] , \mem[653][3] ,
         \mem[653][2] , \mem[653][1] , \mem[653][0] , \mem[652][7] ,
         \mem[652][6] , \mem[652][5] , \mem[652][4] , \mem[652][3] ,
         \mem[652][2] , \mem[652][1] , \mem[652][0] , \mem[651][7] ,
         \mem[651][6] , \mem[651][5] , \mem[651][4] , \mem[651][3] ,
         \mem[651][2] , \mem[651][1] , \mem[651][0] , \mem[650][7] ,
         \mem[650][6] , \mem[650][5] , \mem[650][4] , \mem[650][3] ,
         \mem[650][2] , \mem[650][1] , \mem[650][0] , \mem[649][7] ,
         \mem[649][6] , \mem[649][5] , \mem[649][4] , \mem[649][3] ,
         \mem[649][2] , \mem[649][1] , \mem[649][0] , \mem[648][7] ,
         \mem[648][6] , \mem[648][5] , \mem[648][4] , \mem[648][3] ,
         \mem[648][2] , \mem[648][1] , \mem[648][0] , \mem[647][7] ,
         \mem[647][6] , \mem[647][5] , \mem[647][4] , \mem[647][3] ,
         \mem[647][2] , \mem[647][1] , \mem[647][0] , \mem[646][7] ,
         \mem[646][6] , \mem[646][5] , \mem[646][4] , \mem[646][3] ,
         \mem[646][2] , \mem[646][1] , \mem[646][0] , \mem[645][7] ,
         \mem[645][6] , \mem[645][5] , \mem[645][4] , \mem[645][3] ,
         \mem[645][2] , \mem[645][1] , \mem[645][0] , \mem[644][7] ,
         \mem[644][6] , \mem[644][5] , \mem[644][4] , \mem[644][3] ,
         \mem[644][2] , \mem[644][1] , \mem[644][0] , \mem[643][7] ,
         \mem[643][6] , \mem[643][5] , \mem[643][4] , \mem[643][3] ,
         \mem[643][2] , \mem[643][1] , \mem[643][0] , \mem[642][7] ,
         \mem[642][6] , \mem[642][5] , \mem[642][4] , \mem[642][3] ,
         \mem[642][2] , \mem[642][1] , \mem[642][0] , \mem[641][7] ,
         \mem[641][6] , \mem[641][5] , \mem[641][4] , \mem[641][3] ,
         \mem[641][2] , \mem[641][1] , \mem[641][0] , \mem[640][7] ,
         \mem[640][6] , \mem[640][5] , \mem[640][4] , \mem[640][3] ,
         \mem[640][2] , \mem[640][1] , \mem[640][0] , \mem[639][7] ,
         \mem[639][6] , \mem[639][5] , \mem[639][4] , \mem[639][3] ,
         \mem[639][2] , \mem[639][1] , \mem[639][0] , \mem[638][7] ,
         \mem[638][6] , \mem[638][5] , \mem[638][4] , \mem[638][3] ,
         \mem[638][2] , \mem[638][1] , \mem[638][0] , \mem[637][7] ,
         \mem[637][6] , \mem[637][5] , \mem[637][4] , \mem[637][3] ,
         \mem[637][2] , \mem[637][1] , \mem[637][0] , \mem[636][7] ,
         \mem[636][6] , \mem[636][5] , \mem[636][4] , \mem[636][3] ,
         \mem[636][2] , \mem[636][1] , \mem[636][0] , \mem[635][7] ,
         \mem[635][6] , \mem[635][5] , \mem[635][4] , \mem[635][3] ,
         \mem[635][2] , \mem[635][1] , \mem[635][0] , \mem[634][7] ,
         \mem[634][6] , \mem[634][5] , \mem[634][4] , \mem[634][3] ,
         \mem[634][2] , \mem[634][1] , \mem[634][0] , \mem[633][7] ,
         \mem[633][6] , \mem[633][5] , \mem[633][4] , \mem[633][3] ,
         \mem[633][2] , \mem[633][1] , \mem[633][0] , \mem[632][7] ,
         \mem[632][6] , \mem[632][5] , \mem[632][4] , \mem[632][3] ,
         \mem[632][2] , \mem[632][1] , \mem[632][0] , \mem[631][7] ,
         \mem[631][6] , \mem[631][5] , \mem[631][4] , \mem[631][3] ,
         \mem[631][2] , \mem[631][1] , \mem[631][0] , \mem[630][7] ,
         \mem[630][6] , \mem[630][5] , \mem[630][4] , \mem[630][3] ,
         \mem[630][2] , \mem[630][1] , \mem[630][0] , \mem[629][7] ,
         \mem[629][6] , \mem[629][5] , \mem[629][4] , \mem[629][3] ,
         \mem[629][2] , \mem[629][1] , \mem[629][0] , \mem[628][7] ,
         \mem[628][6] , \mem[628][5] , \mem[628][4] , \mem[628][3] ,
         \mem[628][2] , \mem[628][1] , \mem[628][0] , \mem[627][7] ,
         \mem[627][6] , \mem[627][5] , \mem[627][4] , \mem[627][3] ,
         \mem[627][2] , \mem[627][1] , \mem[627][0] , \mem[626][7] ,
         \mem[626][6] , \mem[626][5] , \mem[626][4] , \mem[626][3] ,
         \mem[626][2] , \mem[626][1] , \mem[626][0] , \mem[625][7] ,
         \mem[625][6] , \mem[625][5] , \mem[625][4] , \mem[625][3] ,
         \mem[625][2] , \mem[625][1] , \mem[625][0] , \mem[624][7] ,
         \mem[624][6] , \mem[624][5] , \mem[624][4] , \mem[624][3] ,
         \mem[624][2] , \mem[624][1] , \mem[624][0] , \mem[623][7] ,
         \mem[623][6] , \mem[623][5] , \mem[623][4] , \mem[623][3] ,
         \mem[623][2] , \mem[623][1] , \mem[623][0] , \mem[622][7] ,
         \mem[622][6] , \mem[622][5] , \mem[622][4] , \mem[622][3] ,
         \mem[622][2] , \mem[622][1] , \mem[622][0] , \mem[621][7] ,
         \mem[621][6] , \mem[621][5] , \mem[621][4] , \mem[621][3] ,
         \mem[621][2] , \mem[621][1] , \mem[621][0] , \mem[620][7] ,
         \mem[620][6] , \mem[620][5] , \mem[620][4] , \mem[620][3] ,
         \mem[620][2] , \mem[620][1] , \mem[620][0] , \mem[619][7] ,
         \mem[619][6] , \mem[619][5] , \mem[619][4] , \mem[619][3] ,
         \mem[619][2] , \mem[619][1] , \mem[619][0] , \mem[618][7] ,
         \mem[618][6] , \mem[618][5] , \mem[618][4] , \mem[618][3] ,
         \mem[618][2] , \mem[618][1] , \mem[618][0] , \mem[617][7] ,
         \mem[617][6] , \mem[617][5] , \mem[617][4] , \mem[617][3] ,
         \mem[617][2] , \mem[617][1] , \mem[617][0] , \mem[616][7] ,
         \mem[616][6] , \mem[616][5] , \mem[616][4] , \mem[616][3] ,
         \mem[616][2] , \mem[616][1] , \mem[616][0] , \mem[615][7] ,
         \mem[615][6] , \mem[615][5] , \mem[615][4] , \mem[615][3] ,
         \mem[615][2] , \mem[615][1] , \mem[615][0] , \mem[614][7] ,
         \mem[614][6] , \mem[614][5] , \mem[614][4] , \mem[614][3] ,
         \mem[614][2] , \mem[614][1] , \mem[614][0] , \mem[613][7] ,
         \mem[613][6] , \mem[613][5] , \mem[613][4] , \mem[613][3] ,
         \mem[613][2] , \mem[613][1] , \mem[613][0] , \mem[612][7] ,
         \mem[612][6] , \mem[612][5] , \mem[612][4] , \mem[612][3] ,
         \mem[612][2] , \mem[612][1] , \mem[612][0] , \mem[611][7] ,
         \mem[611][6] , \mem[611][5] , \mem[611][4] , \mem[611][3] ,
         \mem[611][2] , \mem[611][1] , \mem[611][0] , \mem[610][7] ,
         \mem[610][6] , \mem[610][5] , \mem[610][4] , \mem[610][3] ,
         \mem[610][2] , \mem[610][1] , \mem[610][0] , \mem[609][7] ,
         \mem[609][6] , \mem[609][5] , \mem[609][4] , \mem[609][3] ,
         \mem[609][2] , \mem[609][1] , \mem[609][0] , \mem[608][7] ,
         \mem[608][6] , \mem[608][5] , \mem[608][4] , \mem[608][3] ,
         \mem[608][2] , \mem[608][1] , \mem[608][0] , \mem[607][7] ,
         \mem[607][6] , \mem[607][5] , \mem[607][4] , \mem[607][3] ,
         \mem[607][2] , \mem[607][1] , \mem[607][0] , \mem[606][7] ,
         \mem[606][6] , \mem[606][5] , \mem[606][4] , \mem[606][3] ,
         \mem[606][2] , \mem[606][1] , \mem[606][0] , \mem[605][7] ,
         \mem[605][6] , \mem[605][5] , \mem[605][4] , \mem[605][3] ,
         \mem[605][2] , \mem[605][1] , \mem[605][0] , \mem[604][7] ,
         \mem[604][6] , \mem[604][5] , \mem[604][4] , \mem[604][3] ,
         \mem[604][2] , \mem[604][1] , \mem[604][0] , \mem[603][7] ,
         \mem[603][6] , \mem[603][5] , \mem[603][4] , \mem[603][3] ,
         \mem[603][2] , \mem[603][1] , \mem[603][0] , \mem[602][7] ,
         \mem[602][6] , \mem[602][5] , \mem[602][4] , \mem[602][3] ,
         \mem[602][2] , \mem[602][1] , \mem[602][0] , \mem[601][7] ,
         \mem[601][6] , \mem[601][5] , \mem[601][4] , \mem[601][3] ,
         \mem[601][2] , \mem[601][1] , \mem[601][0] , \mem[600][7] ,
         \mem[600][6] , \mem[600][5] , \mem[600][4] , \mem[600][3] ,
         \mem[600][2] , \mem[600][1] , \mem[600][0] , \mem[599][7] ,
         \mem[599][6] , \mem[599][5] , \mem[599][4] , \mem[599][3] ,
         \mem[599][2] , \mem[599][1] , \mem[599][0] , \mem[598][7] ,
         \mem[598][6] , \mem[598][5] , \mem[598][4] , \mem[598][3] ,
         \mem[598][2] , \mem[598][1] , \mem[598][0] , \mem[597][7] ,
         \mem[597][6] , \mem[597][5] , \mem[597][4] , \mem[597][3] ,
         \mem[597][2] , \mem[597][1] , \mem[597][0] , \mem[596][7] ,
         \mem[596][6] , \mem[596][5] , \mem[596][4] , \mem[596][3] ,
         \mem[596][2] , \mem[596][1] , \mem[596][0] , \mem[595][7] ,
         \mem[595][6] , \mem[595][5] , \mem[595][4] , \mem[595][3] ,
         \mem[595][2] , \mem[595][1] , \mem[595][0] , \mem[594][7] ,
         \mem[594][6] , \mem[594][5] , \mem[594][4] , \mem[594][3] ,
         \mem[594][2] , \mem[594][1] , \mem[594][0] , \mem[593][7] ,
         \mem[593][6] , \mem[593][5] , \mem[593][4] , \mem[593][3] ,
         \mem[593][2] , \mem[593][1] , \mem[593][0] , \mem[592][7] ,
         \mem[592][6] , \mem[592][5] , \mem[592][4] , \mem[592][3] ,
         \mem[592][2] , \mem[592][1] , \mem[592][0] , \mem[591][7] ,
         \mem[591][6] , \mem[591][5] , \mem[591][4] , \mem[591][3] ,
         \mem[591][2] , \mem[591][1] , \mem[591][0] , \mem[590][7] ,
         \mem[590][6] , \mem[590][5] , \mem[590][4] , \mem[590][3] ,
         \mem[590][2] , \mem[590][1] , \mem[590][0] , \mem[589][7] ,
         \mem[589][6] , \mem[589][5] , \mem[589][4] , \mem[589][3] ,
         \mem[589][2] , \mem[589][1] , \mem[589][0] , \mem[588][7] ,
         \mem[588][6] , \mem[588][5] , \mem[588][4] , \mem[588][3] ,
         \mem[588][2] , \mem[588][1] , \mem[588][0] , \mem[587][7] ,
         \mem[587][6] , \mem[587][5] , \mem[587][4] , \mem[587][3] ,
         \mem[587][2] , \mem[587][1] , \mem[587][0] , \mem[586][7] ,
         \mem[586][6] , \mem[586][5] , \mem[586][4] , \mem[586][3] ,
         \mem[586][2] , \mem[586][1] , \mem[586][0] , \mem[585][7] ,
         \mem[585][6] , \mem[585][5] , \mem[585][4] , \mem[585][3] ,
         \mem[585][2] , \mem[585][1] , \mem[585][0] , \mem[584][7] ,
         \mem[584][6] , \mem[584][5] , \mem[584][4] , \mem[584][3] ,
         \mem[584][2] , \mem[584][1] , \mem[584][0] , \mem[583][7] ,
         \mem[583][6] , \mem[583][5] , \mem[583][4] , \mem[583][3] ,
         \mem[583][2] , \mem[583][1] , \mem[583][0] , \mem[582][7] ,
         \mem[582][6] , \mem[582][5] , \mem[582][4] , \mem[582][3] ,
         \mem[582][2] , \mem[582][1] , \mem[582][0] , \mem[581][7] ,
         \mem[581][6] , \mem[581][5] , \mem[581][4] , \mem[581][3] ,
         \mem[581][2] , \mem[581][1] , \mem[581][0] , \mem[580][7] ,
         \mem[580][6] , \mem[580][5] , \mem[580][4] , \mem[580][3] ,
         \mem[580][2] , \mem[580][1] , \mem[580][0] , \mem[579][7] ,
         \mem[579][6] , \mem[579][5] , \mem[579][4] , \mem[579][3] ,
         \mem[579][2] , \mem[579][1] , \mem[579][0] , \mem[578][7] ,
         \mem[578][6] , \mem[578][5] , \mem[578][4] , \mem[578][3] ,
         \mem[578][2] , \mem[578][1] , \mem[578][0] , \mem[577][7] ,
         \mem[577][6] , \mem[577][5] , \mem[577][4] , \mem[577][3] ,
         \mem[577][2] , \mem[577][1] , \mem[577][0] , \mem[576][7] ,
         \mem[576][6] , \mem[576][5] , \mem[576][4] , \mem[576][3] ,
         \mem[576][2] , \mem[576][1] , \mem[576][0] , \mem[575][7] ,
         \mem[575][6] , \mem[575][5] , \mem[575][4] , \mem[575][3] ,
         \mem[575][2] , \mem[575][1] , \mem[575][0] , \mem[574][7] ,
         \mem[574][6] , \mem[574][5] , \mem[574][4] , \mem[574][3] ,
         \mem[574][2] , \mem[574][1] , \mem[574][0] , \mem[573][7] ,
         \mem[573][6] , \mem[573][5] , \mem[573][4] , \mem[573][3] ,
         \mem[573][2] , \mem[573][1] , \mem[573][0] , \mem[572][7] ,
         \mem[572][6] , \mem[572][5] , \mem[572][4] , \mem[572][3] ,
         \mem[572][2] , \mem[572][1] , \mem[572][0] , \mem[571][7] ,
         \mem[571][6] , \mem[571][5] , \mem[571][4] , \mem[571][3] ,
         \mem[571][2] , \mem[571][1] , \mem[571][0] , \mem[570][7] ,
         \mem[570][6] , \mem[570][5] , \mem[570][4] , \mem[570][3] ,
         \mem[570][2] , \mem[570][1] , \mem[570][0] , \mem[569][7] ,
         \mem[569][6] , \mem[569][5] , \mem[569][4] , \mem[569][3] ,
         \mem[569][2] , \mem[569][1] , \mem[569][0] , \mem[568][7] ,
         \mem[568][6] , \mem[568][5] , \mem[568][4] , \mem[568][3] ,
         \mem[568][2] , \mem[568][1] , \mem[568][0] , \mem[567][7] ,
         \mem[567][6] , \mem[567][5] , \mem[567][4] , \mem[567][3] ,
         \mem[567][2] , \mem[567][1] , \mem[567][0] , \mem[566][7] ,
         \mem[566][6] , \mem[566][5] , \mem[566][4] , \mem[566][3] ,
         \mem[566][2] , \mem[566][1] , \mem[566][0] , \mem[565][7] ,
         \mem[565][6] , \mem[565][5] , \mem[565][4] , \mem[565][3] ,
         \mem[565][2] , \mem[565][1] , \mem[565][0] , \mem[564][7] ,
         \mem[564][6] , \mem[564][5] , \mem[564][4] , \mem[564][3] ,
         \mem[564][2] , \mem[564][1] , \mem[564][0] , \mem[563][7] ,
         \mem[563][6] , \mem[563][5] , \mem[563][4] , \mem[563][3] ,
         \mem[563][2] , \mem[563][1] , \mem[563][0] , \mem[562][7] ,
         \mem[562][6] , \mem[562][5] , \mem[562][4] , \mem[562][3] ,
         \mem[562][2] , \mem[562][1] , \mem[562][0] , \mem[561][7] ,
         \mem[561][6] , \mem[561][5] , \mem[561][4] , \mem[561][3] ,
         \mem[561][2] , \mem[561][1] , \mem[561][0] , \mem[560][7] ,
         \mem[560][6] , \mem[560][5] , \mem[560][4] , \mem[560][3] ,
         \mem[560][2] , \mem[560][1] , \mem[560][0] , \mem[559][7] ,
         \mem[559][6] , \mem[559][5] , \mem[559][4] , \mem[559][3] ,
         \mem[559][2] , \mem[559][1] , \mem[559][0] , \mem[558][7] ,
         \mem[558][6] , \mem[558][5] , \mem[558][4] , \mem[558][3] ,
         \mem[558][2] , \mem[558][1] , \mem[558][0] , \mem[557][7] ,
         \mem[557][6] , \mem[557][5] , \mem[557][4] , \mem[557][3] ,
         \mem[557][2] , \mem[557][1] , \mem[557][0] , \mem[556][7] ,
         \mem[556][6] , \mem[556][5] , \mem[556][4] , \mem[556][3] ,
         \mem[556][2] , \mem[556][1] , \mem[556][0] , \mem[555][7] ,
         \mem[555][6] , \mem[555][5] , \mem[555][4] , \mem[555][3] ,
         \mem[555][2] , \mem[555][1] , \mem[555][0] , \mem[554][7] ,
         \mem[554][6] , \mem[554][5] , \mem[554][4] , \mem[554][3] ,
         \mem[554][2] , \mem[554][1] , \mem[554][0] , \mem[553][7] ,
         \mem[553][6] , \mem[553][5] , \mem[553][4] , \mem[553][3] ,
         \mem[553][2] , \mem[553][1] , \mem[553][0] , \mem[552][7] ,
         \mem[552][6] , \mem[552][5] , \mem[552][4] , \mem[552][3] ,
         \mem[552][2] , \mem[552][1] , \mem[552][0] , \mem[551][7] ,
         \mem[551][6] , \mem[551][5] , \mem[551][4] , \mem[551][3] ,
         \mem[551][2] , \mem[551][1] , \mem[551][0] , \mem[550][7] ,
         \mem[550][6] , \mem[550][5] , \mem[550][4] , \mem[550][3] ,
         \mem[550][2] , \mem[550][1] , \mem[550][0] , \mem[549][7] ,
         \mem[549][6] , \mem[549][5] , \mem[549][4] , \mem[549][3] ,
         \mem[549][2] , \mem[549][1] , \mem[549][0] , \mem[548][7] ,
         \mem[548][6] , \mem[548][5] , \mem[548][4] , \mem[548][3] ,
         \mem[548][2] , \mem[548][1] , \mem[548][0] , \mem[547][7] ,
         \mem[547][6] , \mem[547][5] , \mem[547][4] , \mem[547][3] ,
         \mem[547][2] , \mem[547][1] , \mem[547][0] , \mem[546][7] ,
         \mem[546][6] , \mem[546][5] , \mem[546][4] , \mem[546][3] ,
         \mem[546][2] , \mem[546][1] , \mem[546][0] , \mem[545][7] ,
         \mem[545][6] , \mem[545][5] , \mem[545][4] , \mem[545][3] ,
         \mem[545][2] , \mem[545][1] , \mem[545][0] , \mem[544][7] ,
         \mem[544][6] , \mem[544][5] , \mem[544][4] , \mem[544][3] ,
         \mem[544][2] , \mem[544][1] , \mem[544][0] , \mem[543][7] ,
         \mem[543][6] , \mem[543][5] , \mem[543][4] , \mem[543][3] ,
         \mem[543][2] , \mem[543][1] , \mem[543][0] , \mem[542][7] ,
         \mem[542][6] , \mem[542][5] , \mem[542][4] , \mem[542][3] ,
         \mem[542][2] , \mem[542][1] , \mem[542][0] , \mem[541][7] ,
         \mem[541][6] , \mem[541][5] , \mem[541][4] , \mem[541][3] ,
         \mem[541][2] , \mem[541][1] , \mem[541][0] , \mem[540][7] ,
         \mem[540][6] , \mem[540][5] , \mem[540][4] , \mem[540][3] ,
         \mem[540][2] , \mem[540][1] , \mem[540][0] , \mem[539][7] ,
         \mem[539][6] , \mem[539][5] , \mem[539][4] , \mem[539][3] ,
         \mem[539][2] , \mem[539][1] , \mem[539][0] , \mem[538][7] ,
         \mem[538][6] , \mem[538][5] , \mem[538][4] , \mem[538][3] ,
         \mem[538][2] , \mem[538][1] , \mem[538][0] , \mem[537][7] ,
         \mem[537][6] , \mem[537][5] , \mem[537][4] , \mem[537][3] ,
         \mem[537][2] , \mem[537][1] , \mem[537][0] , \mem[536][7] ,
         \mem[536][6] , \mem[536][5] , \mem[536][4] , \mem[536][3] ,
         \mem[536][2] , \mem[536][1] , \mem[536][0] , \mem[535][7] ,
         \mem[535][6] , \mem[535][5] , \mem[535][4] , \mem[535][3] ,
         \mem[535][2] , \mem[535][1] , \mem[535][0] , \mem[534][7] ,
         \mem[534][6] , \mem[534][5] , \mem[534][4] , \mem[534][3] ,
         \mem[534][2] , \mem[534][1] , \mem[534][0] , \mem[533][7] ,
         \mem[533][6] , \mem[533][5] , \mem[533][4] , \mem[533][3] ,
         \mem[533][2] , \mem[533][1] , \mem[533][0] , \mem[532][7] ,
         \mem[532][6] , \mem[532][5] , \mem[532][4] , \mem[532][3] ,
         \mem[532][2] , \mem[532][1] , \mem[532][0] , \mem[531][7] ,
         \mem[531][6] , \mem[531][5] , \mem[531][4] , \mem[531][3] ,
         \mem[531][2] , \mem[531][1] , \mem[531][0] , \mem[530][7] ,
         \mem[530][6] , \mem[530][5] , \mem[530][4] , \mem[530][3] ,
         \mem[530][2] , \mem[530][1] , \mem[530][0] , \mem[529][7] ,
         \mem[529][6] , \mem[529][5] , \mem[529][4] , \mem[529][3] ,
         \mem[529][2] , \mem[529][1] , \mem[529][0] , \mem[528][7] ,
         \mem[528][6] , \mem[528][5] , \mem[528][4] , \mem[528][3] ,
         \mem[528][2] , \mem[528][1] , \mem[528][0] , \mem[527][7] ,
         \mem[527][6] , \mem[527][5] , \mem[527][4] , \mem[527][3] ,
         \mem[527][2] , \mem[527][1] , \mem[527][0] , \mem[526][7] ,
         \mem[526][6] , \mem[526][5] , \mem[526][4] , \mem[526][3] ,
         \mem[526][2] , \mem[526][1] , \mem[526][0] , \mem[525][7] ,
         \mem[525][6] , \mem[525][5] , \mem[525][4] , \mem[525][3] ,
         \mem[525][2] , \mem[525][1] , \mem[525][0] , \mem[524][7] ,
         \mem[524][6] , \mem[524][5] , \mem[524][4] , \mem[524][3] ,
         \mem[524][2] , \mem[524][1] , \mem[524][0] , \mem[523][7] ,
         \mem[523][6] , \mem[523][5] , \mem[523][4] , \mem[523][3] ,
         \mem[523][2] , \mem[523][1] , \mem[523][0] , \mem[522][7] ,
         \mem[522][6] , \mem[522][5] , \mem[522][4] , \mem[522][3] ,
         \mem[522][2] , \mem[522][1] , \mem[522][0] , \mem[521][7] ,
         \mem[521][6] , \mem[521][5] , \mem[521][4] , \mem[521][3] ,
         \mem[521][2] , \mem[521][1] , \mem[521][0] , \mem[520][7] ,
         \mem[520][6] , \mem[520][5] , \mem[520][4] , \mem[520][3] ,
         \mem[520][2] , \mem[520][1] , \mem[520][0] , \mem[519][7] ,
         \mem[519][6] , \mem[519][5] , \mem[519][4] , \mem[519][3] ,
         \mem[519][2] , \mem[519][1] , \mem[519][0] , \mem[518][7] ,
         \mem[518][6] , \mem[518][5] , \mem[518][4] , \mem[518][3] ,
         \mem[518][2] , \mem[518][1] , \mem[518][0] , \mem[517][7] ,
         \mem[517][6] , \mem[517][5] , \mem[517][4] , \mem[517][3] ,
         \mem[517][2] , \mem[517][1] , \mem[517][0] , \mem[516][7] ,
         \mem[516][6] , \mem[516][5] , \mem[516][4] , \mem[516][3] ,
         \mem[516][2] , \mem[516][1] , \mem[516][0] , \mem[515][7] ,
         \mem[515][6] , \mem[515][5] , \mem[515][4] , \mem[515][3] ,
         \mem[515][2] , \mem[515][1] , \mem[515][0] , \mem[514][7] ,
         \mem[514][6] , \mem[514][5] , \mem[514][4] , \mem[514][3] ,
         \mem[514][2] , \mem[514][1] , \mem[514][0] , \mem[513][7] ,
         \mem[513][6] , \mem[513][5] , \mem[513][4] , \mem[513][3] ,
         \mem[513][2] , \mem[513][1] , \mem[513][0] , \mem[512][7] ,
         \mem[512][6] , \mem[512][5] , \mem[512][4] , \mem[512][3] ,
         \mem[512][2] , \mem[512][1] , \mem[512][0] , \mem[511][7] ,
         \mem[511][6] , \mem[511][5] , \mem[511][4] , \mem[511][3] ,
         \mem[511][2] , \mem[511][1] , \mem[511][0] , \mem[510][7] ,
         \mem[510][6] , \mem[510][5] , \mem[510][4] , \mem[510][3] ,
         \mem[510][2] , \mem[510][1] , \mem[510][0] , \mem[509][7] ,
         \mem[509][6] , \mem[509][5] , \mem[509][4] , \mem[509][3] ,
         \mem[509][2] , \mem[509][1] , \mem[509][0] , \mem[508][7] ,
         \mem[508][6] , \mem[508][5] , \mem[508][4] , \mem[508][3] ,
         \mem[508][2] , \mem[508][1] , \mem[508][0] , \mem[507][7] ,
         \mem[507][6] , \mem[507][5] , \mem[507][4] , \mem[507][3] ,
         \mem[507][2] , \mem[507][1] , \mem[507][0] , \mem[506][7] ,
         \mem[506][6] , \mem[506][5] , \mem[506][4] , \mem[506][3] ,
         \mem[506][2] , \mem[506][1] , \mem[506][0] , \mem[505][7] ,
         \mem[505][6] , \mem[505][5] , \mem[505][4] , \mem[505][3] ,
         \mem[505][2] , \mem[505][1] , \mem[505][0] , \mem[504][7] ,
         \mem[504][6] , \mem[504][5] , \mem[504][4] , \mem[504][3] ,
         \mem[504][2] , \mem[504][1] , \mem[504][0] , \mem[503][7] ,
         \mem[503][6] , \mem[503][5] , \mem[503][4] , \mem[503][3] ,
         \mem[503][2] , \mem[503][1] , \mem[503][0] , \mem[502][7] ,
         \mem[502][6] , \mem[502][5] , \mem[502][4] , \mem[502][3] ,
         \mem[502][2] , \mem[502][1] , \mem[502][0] , \mem[501][7] ,
         \mem[501][6] , \mem[501][5] , \mem[501][4] , \mem[501][3] ,
         \mem[501][2] , \mem[501][1] , \mem[501][0] , \mem[500][7] ,
         \mem[500][6] , \mem[500][5] , \mem[500][4] , \mem[500][3] ,
         \mem[500][2] , \mem[500][1] , \mem[500][0] , \mem[499][7] ,
         \mem[499][6] , \mem[499][5] , \mem[499][4] , \mem[499][3] ,
         \mem[499][2] , \mem[499][1] , \mem[499][0] , \mem[498][7] ,
         \mem[498][6] , \mem[498][5] , \mem[498][4] , \mem[498][3] ,
         \mem[498][2] , \mem[498][1] , \mem[498][0] , \mem[497][7] ,
         \mem[497][6] , \mem[497][5] , \mem[497][4] , \mem[497][3] ,
         \mem[497][2] , \mem[497][1] , \mem[497][0] , \mem[496][7] ,
         \mem[496][6] , \mem[496][5] , \mem[496][4] , \mem[496][3] ,
         \mem[496][2] , \mem[496][1] , \mem[496][0] , \mem[495][7] ,
         \mem[495][6] , \mem[495][5] , \mem[495][4] , \mem[495][3] ,
         \mem[495][2] , \mem[495][1] , \mem[495][0] , \mem[494][7] ,
         \mem[494][6] , \mem[494][5] , \mem[494][4] , \mem[494][3] ,
         \mem[494][2] , \mem[494][1] , \mem[494][0] , \mem[493][7] ,
         \mem[493][6] , \mem[493][5] , \mem[493][4] , \mem[493][3] ,
         \mem[493][2] , \mem[493][1] , \mem[493][0] , \mem[492][7] ,
         \mem[492][6] , \mem[492][5] , \mem[492][4] , \mem[492][3] ,
         \mem[492][2] , \mem[492][1] , \mem[492][0] , \mem[491][7] ,
         \mem[491][6] , \mem[491][5] , \mem[491][4] , \mem[491][3] ,
         \mem[491][2] , \mem[491][1] , \mem[491][0] , \mem[490][7] ,
         \mem[490][6] , \mem[490][5] , \mem[490][4] , \mem[490][3] ,
         \mem[490][2] , \mem[490][1] , \mem[490][0] , \mem[489][7] ,
         \mem[489][6] , \mem[489][5] , \mem[489][4] , \mem[489][3] ,
         \mem[489][2] , \mem[489][1] , \mem[489][0] , \mem[488][7] ,
         \mem[488][6] , \mem[488][5] , \mem[488][4] , \mem[488][3] ,
         \mem[488][2] , \mem[488][1] , \mem[488][0] , \mem[487][7] ,
         \mem[487][6] , \mem[487][5] , \mem[487][4] , \mem[487][3] ,
         \mem[487][2] , \mem[487][1] , \mem[487][0] , \mem[486][7] ,
         \mem[486][6] , \mem[486][5] , \mem[486][4] , \mem[486][3] ,
         \mem[486][2] , \mem[486][1] , \mem[486][0] , \mem[485][7] ,
         \mem[485][6] , \mem[485][5] , \mem[485][4] , \mem[485][3] ,
         \mem[485][2] , \mem[485][1] , \mem[485][0] , \mem[484][7] ,
         \mem[484][6] , \mem[484][5] , \mem[484][4] , \mem[484][3] ,
         \mem[484][2] , \mem[484][1] , \mem[484][0] , \mem[483][7] ,
         \mem[483][6] , \mem[483][5] , \mem[483][4] , \mem[483][3] ,
         \mem[483][2] , \mem[483][1] , \mem[483][0] , \mem[482][7] ,
         \mem[482][6] , \mem[482][5] , \mem[482][4] , \mem[482][3] ,
         \mem[482][2] , \mem[482][1] , \mem[482][0] , \mem[481][7] ,
         \mem[481][6] , \mem[481][5] , \mem[481][4] , \mem[481][3] ,
         \mem[481][2] , \mem[481][1] , \mem[481][0] , \mem[480][7] ,
         \mem[480][6] , \mem[480][5] , \mem[480][4] , \mem[480][3] ,
         \mem[480][2] , \mem[480][1] , \mem[480][0] , \mem[479][7] ,
         \mem[479][6] , \mem[479][5] , \mem[479][4] , \mem[479][3] ,
         \mem[479][2] , \mem[479][1] , \mem[479][0] , \mem[478][7] ,
         \mem[478][6] , \mem[478][5] , \mem[478][4] , \mem[478][3] ,
         \mem[478][2] , \mem[478][1] , \mem[478][0] , \mem[477][7] ,
         \mem[477][6] , \mem[477][5] , \mem[477][4] , \mem[477][3] ,
         \mem[477][2] , \mem[477][1] , \mem[477][0] , \mem[476][7] ,
         \mem[476][6] , \mem[476][5] , \mem[476][4] , \mem[476][3] ,
         \mem[476][2] , \mem[476][1] , \mem[476][0] , \mem[475][7] ,
         \mem[475][6] , \mem[475][5] , \mem[475][4] , \mem[475][3] ,
         \mem[475][2] , \mem[475][1] , \mem[475][0] , \mem[474][7] ,
         \mem[474][6] , \mem[474][5] , \mem[474][4] , \mem[474][3] ,
         \mem[474][2] , \mem[474][1] , \mem[474][0] , \mem[473][7] ,
         \mem[473][6] , \mem[473][5] , \mem[473][4] , \mem[473][3] ,
         \mem[473][2] , \mem[473][1] , \mem[473][0] , \mem[472][7] ,
         \mem[472][6] , \mem[472][5] , \mem[472][4] , \mem[472][3] ,
         \mem[472][2] , \mem[472][1] , \mem[472][0] , \mem[471][7] ,
         \mem[471][6] , \mem[471][5] , \mem[471][4] , \mem[471][3] ,
         \mem[471][2] , \mem[471][1] , \mem[471][0] , \mem[470][7] ,
         \mem[470][6] , \mem[470][5] , \mem[470][4] , \mem[470][3] ,
         \mem[470][2] , \mem[470][1] , \mem[470][0] , \mem[469][7] ,
         \mem[469][6] , \mem[469][5] , \mem[469][4] , \mem[469][3] ,
         \mem[469][2] , \mem[469][1] , \mem[469][0] , \mem[468][7] ,
         \mem[468][6] , \mem[468][5] , \mem[468][4] , \mem[468][3] ,
         \mem[468][2] , \mem[468][1] , \mem[468][0] , \mem[467][7] ,
         \mem[467][6] , \mem[467][5] , \mem[467][4] , \mem[467][3] ,
         \mem[467][2] , \mem[467][1] , \mem[467][0] , \mem[466][7] ,
         \mem[466][6] , \mem[466][5] , \mem[466][4] , \mem[466][3] ,
         \mem[466][2] , \mem[466][1] , \mem[466][0] , \mem[465][7] ,
         \mem[465][6] , \mem[465][5] , \mem[465][4] , \mem[465][3] ,
         \mem[465][2] , \mem[465][1] , \mem[465][0] , \mem[464][7] ,
         \mem[464][6] , \mem[464][5] , \mem[464][4] , \mem[464][3] ,
         \mem[464][2] , \mem[464][1] , \mem[464][0] , \mem[463][7] ,
         \mem[463][6] , \mem[463][5] , \mem[463][4] , \mem[463][3] ,
         \mem[463][2] , \mem[463][1] , \mem[463][0] , \mem[462][7] ,
         \mem[462][6] , \mem[462][5] , \mem[462][4] , \mem[462][3] ,
         \mem[462][2] , \mem[462][1] , \mem[462][0] , \mem[461][7] ,
         \mem[461][6] , \mem[461][5] , \mem[461][4] , \mem[461][3] ,
         \mem[461][2] , \mem[461][1] , \mem[461][0] , \mem[460][7] ,
         \mem[460][6] , \mem[460][5] , \mem[460][4] , \mem[460][3] ,
         \mem[460][2] , \mem[460][1] , \mem[460][0] , \mem[459][7] ,
         \mem[459][6] , \mem[459][5] , \mem[459][4] , \mem[459][3] ,
         \mem[459][2] , \mem[459][1] , \mem[459][0] , \mem[458][7] ,
         \mem[458][6] , \mem[458][5] , \mem[458][4] , \mem[458][3] ,
         \mem[458][2] , \mem[458][1] , \mem[458][0] , \mem[457][7] ,
         \mem[457][6] , \mem[457][5] , \mem[457][4] , \mem[457][3] ,
         \mem[457][2] , \mem[457][1] , \mem[457][0] , \mem[456][7] ,
         \mem[456][6] , \mem[456][5] , \mem[456][4] , \mem[456][3] ,
         \mem[456][2] , \mem[456][1] , \mem[456][0] , \mem[455][7] ,
         \mem[455][6] , \mem[455][5] , \mem[455][4] , \mem[455][3] ,
         \mem[455][2] , \mem[455][1] , \mem[455][0] , \mem[454][7] ,
         \mem[454][6] , \mem[454][5] , \mem[454][4] , \mem[454][3] ,
         \mem[454][2] , \mem[454][1] , \mem[454][0] , \mem[453][7] ,
         \mem[453][6] , \mem[453][5] , \mem[453][4] , \mem[453][3] ,
         \mem[453][2] , \mem[453][1] , \mem[453][0] , \mem[452][7] ,
         \mem[452][6] , \mem[452][5] , \mem[452][4] , \mem[452][3] ,
         \mem[452][2] , \mem[452][1] , \mem[452][0] , \mem[451][7] ,
         \mem[451][6] , \mem[451][5] , \mem[451][4] , \mem[451][3] ,
         \mem[451][2] , \mem[451][1] , \mem[451][0] , \mem[450][7] ,
         \mem[450][6] , \mem[450][5] , \mem[450][4] , \mem[450][3] ,
         \mem[450][2] , \mem[450][1] , \mem[450][0] , \mem[449][7] ,
         \mem[449][6] , \mem[449][5] , \mem[449][4] , \mem[449][3] ,
         \mem[449][2] , \mem[449][1] , \mem[449][0] , \mem[448][7] ,
         \mem[448][6] , \mem[448][5] , \mem[448][4] , \mem[448][3] ,
         \mem[448][2] , \mem[448][1] , \mem[448][0] , \mem[447][7] ,
         \mem[447][6] , \mem[447][5] , \mem[447][4] , \mem[447][3] ,
         \mem[447][2] , \mem[447][1] , \mem[447][0] , \mem[446][7] ,
         \mem[446][6] , \mem[446][5] , \mem[446][4] , \mem[446][3] ,
         \mem[446][2] , \mem[446][1] , \mem[446][0] , \mem[445][7] ,
         \mem[445][6] , \mem[445][5] , \mem[445][4] , \mem[445][3] ,
         \mem[445][2] , \mem[445][1] , \mem[445][0] , \mem[444][7] ,
         \mem[444][6] , \mem[444][5] , \mem[444][4] , \mem[444][3] ,
         \mem[444][2] , \mem[444][1] , \mem[444][0] , \mem[443][7] ,
         \mem[443][6] , \mem[443][5] , \mem[443][4] , \mem[443][3] ,
         \mem[443][2] , \mem[443][1] , \mem[443][0] , \mem[442][7] ,
         \mem[442][6] , \mem[442][5] , \mem[442][4] , \mem[442][3] ,
         \mem[442][2] , \mem[442][1] , \mem[442][0] , \mem[441][7] ,
         \mem[441][6] , \mem[441][5] , \mem[441][4] , \mem[441][3] ,
         \mem[441][2] , \mem[441][1] , \mem[441][0] , \mem[440][7] ,
         \mem[440][6] , \mem[440][5] , \mem[440][4] , \mem[440][3] ,
         \mem[440][2] , \mem[440][1] , \mem[440][0] , \mem[439][7] ,
         \mem[439][6] , \mem[439][5] , \mem[439][4] , \mem[439][3] ,
         \mem[439][2] , \mem[439][1] , \mem[439][0] , \mem[438][7] ,
         \mem[438][6] , \mem[438][5] , \mem[438][4] , \mem[438][3] ,
         \mem[438][2] , \mem[438][1] , \mem[438][0] , \mem[437][7] ,
         \mem[437][6] , \mem[437][5] , \mem[437][4] , \mem[437][3] ,
         \mem[437][2] , \mem[437][1] , \mem[437][0] , \mem[436][7] ,
         \mem[436][6] , \mem[436][5] , \mem[436][4] , \mem[436][3] ,
         \mem[436][2] , \mem[436][1] , \mem[436][0] , \mem[435][7] ,
         \mem[435][6] , \mem[435][5] , \mem[435][4] , \mem[435][3] ,
         \mem[435][2] , \mem[435][1] , \mem[435][0] , \mem[434][7] ,
         \mem[434][6] , \mem[434][5] , \mem[434][4] , \mem[434][3] ,
         \mem[434][2] , \mem[434][1] , \mem[434][0] , \mem[433][7] ,
         \mem[433][6] , \mem[433][5] , \mem[433][4] , \mem[433][3] ,
         \mem[433][2] , \mem[433][1] , \mem[433][0] , \mem[432][7] ,
         \mem[432][6] , \mem[432][5] , \mem[432][4] , \mem[432][3] ,
         \mem[432][2] , \mem[432][1] , \mem[432][0] , \mem[431][7] ,
         \mem[431][6] , \mem[431][5] , \mem[431][4] , \mem[431][3] ,
         \mem[431][2] , \mem[431][1] , \mem[431][0] , \mem[430][7] ,
         \mem[430][6] , \mem[430][5] , \mem[430][4] , \mem[430][3] ,
         \mem[430][2] , \mem[430][1] , \mem[430][0] , \mem[429][7] ,
         \mem[429][6] , \mem[429][5] , \mem[429][4] , \mem[429][3] ,
         \mem[429][2] , \mem[429][1] , \mem[429][0] , \mem[428][7] ,
         \mem[428][6] , \mem[428][5] , \mem[428][4] , \mem[428][3] ,
         \mem[428][2] , \mem[428][1] , \mem[428][0] , \mem[427][7] ,
         \mem[427][6] , \mem[427][5] , \mem[427][4] , \mem[427][3] ,
         \mem[427][2] , \mem[427][1] , \mem[427][0] , \mem[426][7] ,
         \mem[426][6] , \mem[426][5] , \mem[426][4] , \mem[426][3] ,
         \mem[426][2] , \mem[426][1] , \mem[426][0] , \mem[425][7] ,
         \mem[425][6] , \mem[425][5] , \mem[425][4] , \mem[425][3] ,
         \mem[425][2] , \mem[425][1] , \mem[425][0] , \mem[424][7] ,
         \mem[424][6] , \mem[424][5] , \mem[424][4] , \mem[424][3] ,
         \mem[424][2] , \mem[424][1] , \mem[424][0] , \mem[423][7] ,
         \mem[423][6] , \mem[423][5] , \mem[423][4] , \mem[423][3] ,
         \mem[423][2] , \mem[423][1] , \mem[423][0] , \mem[422][7] ,
         \mem[422][6] , \mem[422][5] , \mem[422][4] , \mem[422][3] ,
         \mem[422][2] , \mem[422][1] , \mem[422][0] , \mem[421][7] ,
         \mem[421][6] , \mem[421][5] , \mem[421][4] , \mem[421][3] ,
         \mem[421][2] , \mem[421][1] , \mem[421][0] , \mem[420][7] ,
         \mem[420][6] , \mem[420][5] , \mem[420][4] , \mem[420][3] ,
         \mem[420][2] , \mem[420][1] , \mem[420][0] , \mem[419][7] ,
         \mem[419][6] , \mem[419][5] , \mem[419][4] , \mem[419][3] ,
         \mem[419][2] , \mem[419][1] , \mem[419][0] , \mem[418][7] ,
         \mem[418][6] , \mem[418][5] , \mem[418][4] , \mem[418][3] ,
         \mem[418][2] , \mem[418][1] , \mem[418][0] , \mem[417][7] ,
         \mem[417][6] , \mem[417][5] , \mem[417][4] , \mem[417][3] ,
         \mem[417][2] , \mem[417][1] , \mem[417][0] , \mem[416][7] ,
         \mem[416][6] , \mem[416][5] , \mem[416][4] , \mem[416][3] ,
         \mem[416][2] , \mem[416][1] , \mem[416][0] , \mem[415][7] ,
         \mem[415][6] , \mem[415][5] , \mem[415][4] , \mem[415][3] ,
         \mem[415][2] , \mem[415][1] , \mem[415][0] , \mem[414][7] ,
         \mem[414][6] , \mem[414][5] , \mem[414][4] , \mem[414][3] ,
         \mem[414][2] , \mem[414][1] , \mem[414][0] , \mem[413][7] ,
         \mem[413][6] , \mem[413][5] , \mem[413][4] , \mem[413][3] ,
         \mem[413][2] , \mem[413][1] , \mem[413][0] , \mem[412][7] ,
         \mem[412][6] , \mem[412][5] , \mem[412][4] , \mem[412][3] ,
         \mem[412][2] , \mem[412][1] , \mem[412][0] , \mem[411][7] ,
         \mem[411][6] , \mem[411][5] , \mem[411][4] , \mem[411][3] ,
         \mem[411][2] , \mem[411][1] , \mem[411][0] , \mem[410][7] ,
         \mem[410][6] , \mem[410][5] , \mem[410][4] , \mem[410][3] ,
         \mem[410][2] , \mem[410][1] , \mem[410][0] , \mem[409][7] ,
         \mem[409][6] , \mem[409][5] , \mem[409][4] , \mem[409][3] ,
         \mem[409][2] , \mem[409][1] , \mem[409][0] , \mem[408][7] ,
         \mem[408][6] , \mem[408][5] , \mem[408][4] , \mem[408][3] ,
         \mem[408][2] , \mem[408][1] , \mem[408][0] , \mem[407][7] ,
         \mem[407][6] , \mem[407][5] , \mem[407][4] , \mem[407][3] ,
         \mem[407][2] , \mem[407][1] , \mem[407][0] , \mem[406][7] ,
         \mem[406][6] , \mem[406][5] , \mem[406][4] , \mem[406][3] ,
         \mem[406][2] , \mem[406][1] , \mem[406][0] , \mem[405][7] ,
         \mem[405][6] , \mem[405][5] , \mem[405][4] , \mem[405][3] ,
         \mem[405][2] , \mem[405][1] , \mem[405][0] , \mem[404][7] ,
         \mem[404][6] , \mem[404][5] , \mem[404][4] , \mem[404][3] ,
         \mem[404][2] , \mem[404][1] , \mem[404][0] , \mem[403][7] ,
         \mem[403][6] , \mem[403][5] , \mem[403][4] , \mem[403][3] ,
         \mem[403][2] , \mem[403][1] , \mem[403][0] , \mem[402][7] ,
         \mem[402][6] , \mem[402][5] , \mem[402][4] , \mem[402][3] ,
         \mem[402][2] , \mem[402][1] , \mem[402][0] , \mem[401][7] ,
         \mem[401][6] , \mem[401][5] , \mem[401][4] , \mem[401][3] ,
         \mem[401][2] , \mem[401][1] , \mem[401][0] , \mem[400][7] ,
         \mem[400][6] , \mem[400][5] , \mem[400][4] , \mem[400][3] ,
         \mem[400][2] , \mem[400][1] , \mem[400][0] , \mem[399][7] ,
         \mem[399][6] , \mem[399][5] , \mem[399][4] , \mem[399][3] ,
         \mem[399][2] , \mem[399][1] , \mem[399][0] , \mem[398][7] ,
         \mem[398][6] , \mem[398][5] , \mem[398][4] , \mem[398][3] ,
         \mem[398][2] , \mem[398][1] , \mem[398][0] , \mem[397][7] ,
         \mem[397][6] , \mem[397][5] , \mem[397][4] , \mem[397][3] ,
         \mem[397][2] , \mem[397][1] , \mem[397][0] , \mem[396][7] ,
         \mem[396][6] , \mem[396][5] , \mem[396][4] , \mem[396][3] ,
         \mem[396][2] , \mem[396][1] , \mem[396][0] , \mem[395][7] ,
         \mem[395][6] , \mem[395][5] , \mem[395][4] , \mem[395][3] ,
         \mem[395][2] , \mem[395][1] , \mem[395][0] , \mem[394][7] ,
         \mem[394][6] , \mem[394][5] , \mem[394][4] , \mem[394][3] ,
         \mem[394][2] , \mem[394][1] , \mem[394][0] , \mem[393][7] ,
         \mem[393][6] , \mem[393][5] , \mem[393][4] , \mem[393][3] ,
         \mem[393][2] , \mem[393][1] , \mem[393][0] , \mem[392][7] ,
         \mem[392][6] , \mem[392][5] , \mem[392][4] , \mem[392][3] ,
         \mem[392][2] , \mem[392][1] , \mem[392][0] , \mem[391][7] ,
         \mem[391][6] , \mem[391][5] , \mem[391][4] , \mem[391][3] ,
         \mem[391][2] , \mem[391][1] , \mem[391][0] , \mem[390][7] ,
         \mem[390][6] , \mem[390][5] , \mem[390][4] , \mem[390][3] ,
         \mem[390][2] , \mem[390][1] , \mem[390][0] , \mem[389][7] ,
         \mem[389][6] , \mem[389][5] , \mem[389][4] , \mem[389][3] ,
         \mem[389][2] , \mem[389][1] , \mem[389][0] , \mem[388][7] ,
         \mem[388][6] , \mem[388][5] , \mem[388][4] , \mem[388][3] ,
         \mem[388][2] , \mem[388][1] , \mem[388][0] , \mem[387][7] ,
         \mem[387][6] , \mem[387][5] , \mem[387][4] , \mem[387][3] ,
         \mem[387][2] , \mem[387][1] , \mem[387][0] , \mem[386][7] ,
         \mem[386][6] , \mem[386][5] , \mem[386][4] , \mem[386][3] ,
         \mem[386][2] , \mem[386][1] , \mem[386][0] , \mem[385][7] ,
         \mem[385][6] , \mem[385][5] , \mem[385][4] , \mem[385][3] ,
         \mem[385][2] , \mem[385][1] , \mem[385][0] , \mem[384][7] ,
         \mem[384][6] , \mem[384][5] , \mem[384][4] , \mem[384][3] ,
         \mem[384][2] , \mem[384][1] , \mem[384][0] , \mem[383][7] ,
         \mem[383][6] , \mem[383][5] , \mem[383][4] , \mem[383][3] ,
         \mem[383][2] , \mem[383][1] , \mem[383][0] , \mem[382][7] ,
         \mem[382][6] , \mem[382][5] , \mem[382][4] , \mem[382][3] ,
         \mem[382][2] , \mem[382][1] , \mem[382][0] , \mem[381][7] ,
         \mem[381][6] , \mem[381][5] , \mem[381][4] , \mem[381][3] ,
         \mem[381][2] , \mem[381][1] , \mem[381][0] , \mem[380][7] ,
         \mem[380][6] , \mem[380][5] , \mem[380][4] , \mem[380][3] ,
         \mem[380][2] , \mem[380][1] , \mem[380][0] , \mem[379][7] ,
         \mem[379][6] , \mem[379][5] , \mem[379][4] , \mem[379][3] ,
         \mem[379][2] , \mem[379][1] , \mem[379][0] , \mem[378][7] ,
         \mem[378][6] , \mem[378][5] , \mem[378][4] , \mem[378][3] ,
         \mem[378][2] , \mem[378][1] , \mem[378][0] , \mem[377][7] ,
         \mem[377][6] , \mem[377][5] , \mem[377][4] , \mem[377][3] ,
         \mem[377][2] , \mem[377][1] , \mem[377][0] , \mem[376][7] ,
         \mem[376][6] , \mem[376][5] , \mem[376][4] , \mem[376][3] ,
         \mem[376][2] , \mem[376][1] , \mem[376][0] , \mem[375][7] ,
         \mem[375][6] , \mem[375][5] , \mem[375][4] , \mem[375][3] ,
         \mem[375][2] , \mem[375][1] , \mem[375][0] , \mem[374][7] ,
         \mem[374][6] , \mem[374][5] , \mem[374][4] , \mem[374][3] ,
         \mem[374][2] , \mem[374][1] , \mem[374][0] , \mem[373][7] ,
         \mem[373][6] , \mem[373][5] , \mem[373][4] , \mem[373][3] ,
         \mem[373][2] , \mem[373][1] , \mem[373][0] , \mem[372][7] ,
         \mem[372][6] , \mem[372][5] , \mem[372][4] , \mem[372][3] ,
         \mem[372][2] , \mem[372][1] , \mem[372][0] , \mem[371][7] ,
         \mem[371][6] , \mem[371][5] , \mem[371][4] , \mem[371][3] ,
         \mem[371][2] , \mem[371][1] , \mem[371][0] , \mem[370][7] ,
         \mem[370][6] , \mem[370][5] , \mem[370][4] , \mem[370][3] ,
         \mem[370][2] , \mem[370][1] , \mem[370][0] , \mem[369][7] ,
         \mem[369][6] , \mem[369][5] , \mem[369][4] , \mem[369][3] ,
         \mem[369][2] , \mem[369][1] , \mem[369][0] , \mem[368][7] ,
         \mem[368][6] , \mem[368][5] , \mem[368][4] , \mem[368][3] ,
         \mem[368][2] , \mem[368][1] , \mem[368][0] , \mem[367][7] ,
         \mem[367][6] , \mem[367][5] , \mem[367][4] , \mem[367][3] ,
         \mem[367][2] , \mem[367][1] , \mem[367][0] , \mem[366][7] ,
         \mem[366][6] , \mem[366][5] , \mem[366][4] , \mem[366][3] ,
         \mem[366][2] , \mem[366][1] , \mem[366][0] , \mem[365][7] ,
         \mem[365][6] , \mem[365][5] , \mem[365][4] , \mem[365][3] ,
         \mem[365][2] , \mem[365][1] , \mem[365][0] , \mem[364][7] ,
         \mem[364][6] , \mem[364][5] , \mem[364][4] , \mem[364][3] ,
         \mem[364][2] , \mem[364][1] , \mem[364][0] , \mem[363][7] ,
         \mem[363][6] , \mem[363][5] , \mem[363][4] , \mem[363][3] ,
         \mem[363][2] , \mem[363][1] , \mem[363][0] , \mem[362][7] ,
         \mem[362][6] , \mem[362][5] , \mem[362][4] , \mem[362][3] ,
         \mem[362][2] , \mem[362][1] , \mem[362][0] , \mem[361][7] ,
         \mem[361][6] , \mem[361][5] , \mem[361][4] , \mem[361][3] ,
         \mem[361][2] , \mem[361][1] , \mem[361][0] , \mem[360][7] ,
         \mem[360][6] , \mem[360][5] , \mem[360][4] , \mem[360][3] ,
         \mem[360][2] , \mem[360][1] , \mem[360][0] , \mem[359][7] ,
         \mem[359][6] , \mem[359][5] , \mem[359][4] , \mem[359][3] ,
         \mem[359][2] , \mem[359][1] , \mem[359][0] , \mem[358][7] ,
         \mem[358][6] , \mem[358][5] , \mem[358][4] , \mem[358][3] ,
         \mem[358][2] , \mem[358][1] , \mem[358][0] , \mem[357][7] ,
         \mem[357][6] , \mem[357][5] , \mem[357][4] , \mem[357][3] ,
         \mem[357][2] , \mem[357][1] , \mem[357][0] , \mem[356][7] ,
         \mem[356][6] , \mem[356][5] , \mem[356][4] , \mem[356][3] ,
         \mem[356][2] , \mem[356][1] , \mem[356][0] , \mem[355][7] ,
         \mem[355][6] , \mem[355][5] , \mem[355][4] , \mem[355][3] ,
         \mem[355][2] , \mem[355][1] , \mem[355][0] , \mem[354][7] ,
         \mem[354][6] , \mem[354][5] , \mem[354][4] , \mem[354][3] ,
         \mem[354][2] , \mem[354][1] , \mem[354][0] , \mem[353][7] ,
         \mem[353][6] , \mem[353][5] , \mem[353][4] , \mem[353][3] ,
         \mem[353][2] , \mem[353][1] , \mem[353][0] , \mem[352][7] ,
         \mem[352][6] , \mem[352][5] , \mem[352][4] , \mem[352][3] ,
         \mem[352][2] , \mem[352][1] , \mem[352][0] , \mem[351][7] ,
         \mem[351][6] , \mem[351][5] , \mem[351][4] , \mem[351][3] ,
         \mem[351][2] , \mem[351][1] , \mem[351][0] , \mem[350][7] ,
         \mem[350][6] , \mem[350][5] , \mem[350][4] , \mem[350][3] ,
         \mem[350][2] , \mem[350][1] , \mem[350][0] , \mem[349][7] ,
         \mem[349][6] , \mem[349][5] , \mem[349][4] , \mem[349][3] ,
         \mem[349][2] , \mem[349][1] , \mem[349][0] , \mem[348][7] ,
         \mem[348][6] , \mem[348][5] , \mem[348][4] , \mem[348][3] ,
         \mem[348][2] , \mem[348][1] , \mem[348][0] , \mem[347][7] ,
         \mem[347][6] , \mem[347][5] , \mem[347][4] , \mem[347][3] ,
         \mem[347][2] , \mem[347][1] , \mem[347][0] , \mem[346][7] ,
         \mem[346][6] , \mem[346][5] , \mem[346][4] , \mem[346][3] ,
         \mem[346][2] , \mem[346][1] , \mem[346][0] , \mem[345][7] ,
         \mem[345][6] , \mem[345][5] , \mem[345][4] , \mem[345][3] ,
         \mem[345][2] , \mem[345][1] , \mem[345][0] , \mem[344][7] ,
         \mem[344][6] , \mem[344][5] , \mem[344][4] , \mem[344][3] ,
         \mem[344][2] , \mem[344][1] , \mem[344][0] , \mem[343][7] ,
         \mem[343][6] , \mem[343][5] , \mem[343][4] , \mem[343][3] ,
         \mem[343][2] , \mem[343][1] , \mem[343][0] , \mem[342][7] ,
         \mem[342][6] , \mem[342][5] , \mem[342][4] , \mem[342][3] ,
         \mem[342][2] , \mem[342][1] , \mem[342][0] , \mem[341][7] ,
         \mem[341][6] , \mem[341][5] , \mem[341][4] , \mem[341][3] ,
         \mem[341][2] , \mem[341][1] , \mem[341][0] , \mem[340][7] ,
         \mem[340][6] , \mem[340][5] , \mem[340][4] , \mem[340][3] ,
         \mem[340][2] , \mem[340][1] , \mem[340][0] , \mem[339][7] ,
         \mem[339][6] , \mem[339][5] , \mem[339][4] , \mem[339][3] ,
         \mem[339][2] , \mem[339][1] , \mem[339][0] , \mem[338][7] ,
         \mem[338][6] , \mem[338][5] , \mem[338][4] , \mem[338][3] ,
         \mem[338][2] , \mem[338][1] , \mem[338][0] , \mem[337][7] ,
         \mem[337][6] , \mem[337][5] , \mem[337][4] , \mem[337][3] ,
         \mem[337][2] , \mem[337][1] , \mem[337][0] , \mem[336][7] ,
         \mem[336][6] , \mem[336][5] , \mem[336][4] , \mem[336][3] ,
         \mem[336][2] , \mem[336][1] , \mem[336][0] , \mem[335][7] ,
         \mem[335][6] , \mem[335][5] , \mem[335][4] , \mem[335][3] ,
         \mem[335][2] , \mem[335][1] , \mem[335][0] , \mem[334][7] ,
         \mem[334][6] , \mem[334][5] , \mem[334][4] , \mem[334][3] ,
         \mem[334][2] , \mem[334][1] , \mem[334][0] , \mem[333][7] ,
         \mem[333][6] , \mem[333][5] , \mem[333][4] , \mem[333][3] ,
         \mem[333][2] , \mem[333][1] , \mem[333][0] , \mem[332][7] ,
         \mem[332][6] , \mem[332][5] , \mem[332][4] , \mem[332][3] ,
         \mem[332][2] , \mem[332][1] , \mem[332][0] , \mem[331][7] ,
         \mem[331][6] , \mem[331][5] , \mem[331][4] , \mem[331][3] ,
         \mem[331][2] , \mem[331][1] , \mem[331][0] , \mem[330][7] ,
         \mem[330][6] , \mem[330][5] , \mem[330][4] , \mem[330][3] ,
         \mem[330][2] , \mem[330][1] , \mem[330][0] , \mem[329][7] ,
         \mem[329][6] , \mem[329][5] , \mem[329][4] , \mem[329][3] ,
         \mem[329][2] , \mem[329][1] , \mem[329][0] , \mem[328][7] ,
         \mem[328][6] , \mem[328][5] , \mem[328][4] , \mem[328][3] ,
         \mem[328][2] , \mem[328][1] , \mem[328][0] , \mem[327][7] ,
         \mem[327][6] , \mem[327][5] , \mem[327][4] , \mem[327][3] ,
         \mem[327][2] , \mem[327][1] , \mem[327][0] , \mem[326][7] ,
         \mem[326][6] , \mem[326][5] , \mem[326][4] , \mem[326][3] ,
         \mem[326][2] , \mem[326][1] , \mem[326][0] , \mem[325][7] ,
         \mem[325][6] , \mem[325][5] , \mem[325][4] , \mem[325][3] ,
         \mem[325][2] , \mem[325][1] , \mem[325][0] , \mem[324][7] ,
         \mem[324][6] , \mem[324][5] , \mem[324][4] , \mem[324][3] ,
         \mem[324][2] , \mem[324][1] , \mem[324][0] , \mem[323][7] ,
         \mem[323][6] , \mem[323][5] , \mem[323][4] , \mem[323][3] ,
         \mem[323][2] , \mem[323][1] , \mem[323][0] , \mem[322][7] ,
         \mem[322][6] , \mem[322][5] , \mem[322][4] , \mem[322][3] ,
         \mem[322][2] , \mem[322][1] , \mem[322][0] , \mem[321][7] ,
         \mem[321][6] , \mem[321][5] , \mem[321][4] , \mem[321][3] ,
         \mem[321][2] , \mem[321][1] , \mem[321][0] , \mem[320][7] ,
         \mem[320][6] , \mem[320][5] , \mem[320][4] , \mem[320][3] ,
         \mem[320][2] , \mem[320][1] , \mem[320][0] , \mem[319][7] ,
         \mem[319][6] , \mem[319][5] , \mem[319][4] , \mem[319][3] ,
         \mem[319][2] , \mem[319][1] , \mem[319][0] , \mem[318][7] ,
         \mem[318][6] , \mem[318][5] , \mem[318][4] , \mem[318][3] ,
         \mem[318][2] , \mem[318][1] , \mem[318][0] , \mem[317][7] ,
         \mem[317][6] , \mem[317][5] , \mem[317][4] , \mem[317][3] ,
         \mem[317][2] , \mem[317][1] , \mem[317][0] , \mem[316][7] ,
         \mem[316][6] , \mem[316][5] , \mem[316][4] , \mem[316][3] ,
         \mem[316][2] , \mem[316][1] , \mem[316][0] , \mem[315][7] ,
         \mem[315][6] , \mem[315][5] , \mem[315][4] , \mem[315][3] ,
         \mem[315][2] , \mem[315][1] , \mem[315][0] , \mem[314][7] ,
         \mem[314][6] , \mem[314][5] , \mem[314][4] , \mem[314][3] ,
         \mem[314][2] , \mem[314][1] , \mem[314][0] , \mem[313][7] ,
         \mem[313][6] , \mem[313][5] , \mem[313][4] , \mem[313][3] ,
         \mem[313][2] , \mem[313][1] , \mem[313][0] , \mem[312][7] ,
         \mem[312][6] , \mem[312][5] , \mem[312][4] , \mem[312][3] ,
         \mem[312][2] , \mem[312][1] , \mem[312][0] , \mem[311][7] ,
         \mem[311][6] , \mem[311][5] , \mem[311][4] , \mem[311][3] ,
         \mem[311][2] , \mem[311][1] , \mem[311][0] , \mem[310][7] ,
         \mem[310][6] , \mem[310][5] , \mem[310][4] , \mem[310][3] ,
         \mem[310][2] , \mem[310][1] , \mem[310][0] , \mem[309][7] ,
         \mem[309][6] , \mem[309][5] , \mem[309][4] , \mem[309][3] ,
         \mem[309][2] , \mem[309][1] , \mem[309][0] , \mem[308][7] ,
         \mem[308][6] , \mem[308][5] , \mem[308][4] , \mem[308][3] ,
         \mem[308][2] , \mem[308][1] , \mem[308][0] , \mem[307][7] ,
         \mem[307][6] , \mem[307][5] , \mem[307][4] , \mem[307][3] ,
         \mem[307][2] , \mem[307][1] , \mem[307][0] , \mem[306][7] ,
         \mem[306][6] , \mem[306][5] , \mem[306][4] , \mem[306][3] ,
         \mem[306][2] , \mem[306][1] , \mem[306][0] , \mem[305][7] ,
         \mem[305][6] , \mem[305][5] , \mem[305][4] , \mem[305][3] ,
         \mem[305][2] , \mem[305][1] , \mem[305][0] , \mem[304][7] ,
         \mem[304][6] , \mem[304][5] , \mem[304][4] , \mem[304][3] ,
         \mem[304][2] , \mem[304][1] , \mem[304][0] , \mem[303][7] ,
         \mem[303][6] , \mem[303][5] , \mem[303][4] , \mem[303][3] ,
         \mem[303][2] , \mem[303][1] , \mem[303][0] , \mem[302][7] ,
         \mem[302][6] , \mem[302][5] , \mem[302][4] , \mem[302][3] ,
         \mem[302][2] , \mem[302][1] , \mem[302][0] , \mem[301][7] ,
         \mem[301][6] , \mem[301][5] , \mem[301][4] , \mem[301][3] ,
         \mem[301][2] , \mem[301][1] , \mem[301][0] , \mem[300][7] ,
         \mem[300][6] , \mem[300][5] , \mem[300][4] , \mem[300][3] ,
         \mem[300][2] , \mem[300][1] , \mem[300][0] , \mem[299][7] ,
         \mem[299][6] , \mem[299][5] , \mem[299][4] , \mem[299][3] ,
         \mem[299][2] , \mem[299][1] , \mem[299][0] , \mem[298][7] ,
         \mem[298][6] , \mem[298][5] , \mem[298][4] , \mem[298][3] ,
         \mem[298][2] , \mem[298][1] , \mem[298][0] , \mem[297][7] ,
         \mem[297][6] , \mem[297][5] , \mem[297][4] , \mem[297][3] ,
         \mem[297][2] , \mem[297][1] , \mem[297][0] , \mem[296][7] ,
         \mem[296][6] , \mem[296][5] , \mem[296][4] , \mem[296][3] ,
         \mem[296][2] , \mem[296][1] , \mem[296][0] , \mem[295][7] ,
         \mem[295][6] , \mem[295][5] , \mem[295][4] , \mem[295][3] ,
         \mem[295][2] , \mem[295][1] , \mem[295][0] , \mem[294][7] ,
         \mem[294][6] , \mem[294][5] , \mem[294][4] , \mem[294][3] ,
         \mem[294][2] , \mem[294][1] , \mem[294][0] , \mem[293][7] ,
         \mem[293][6] , \mem[293][5] , \mem[293][4] , \mem[293][3] ,
         \mem[293][2] , \mem[293][1] , \mem[293][0] , \mem[292][7] ,
         \mem[292][6] , \mem[292][5] , \mem[292][4] , \mem[292][3] ,
         \mem[292][2] , \mem[292][1] , \mem[292][0] , \mem[291][7] ,
         \mem[291][6] , \mem[291][5] , \mem[291][4] , \mem[291][3] ,
         \mem[291][2] , \mem[291][1] , \mem[291][0] , \mem[290][7] ,
         \mem[290][6] , \mem[290][5] , \mem[290][4] , \mem[290][3] ,
         \mem[290][2] , \mem[290][1] , \mem[290][0] , \mem[289][7] ,
         \mem[289][6] , \mem[289][5] , \mem[289][4] , \mem[289][3] ,
         \mem[289][2] , \mem[289][1] , \mem[289][0] , \mem[288][7] ,
         \mem[288][6] , \mem[288][5] , \mem[288][4] , \mem[288][3] ,
         \mem[288][2] , \mem[288][1] , \mem[288][0] , \mem[287][7] ,
         \mem[287][6] , \mem[287][5] , \mem[287][4] , \mem[287][3] ,
         \mem[287][2] , \mem[287][1] , \mem[287][0] , \mem[286][7] ,
         \mem[286][6] , \mem[286][5] , \mem[286][4] , \mem[286][3] ,
         \mem[286][2] , \mem[286][1] , \mem[286][0] , \mem[285][7] ,
         \mem[285][6] , \mem[285][5] , \mem[285][4] , \mem[285][3] ,
         \mem[285][2] , \mem[285][1] , \mem[285][0] , \mem[284][7] ,
         \mem[284][6] , \mem[284][5] , \mem[284][4] , \mem[284][3] ,
         \mem[284][2] , \mem[284][1] , \mem[284][0] , \mem[283][7] ,
         \mem[283][6] , \mem[283][5] , \mem[283][4] , \mem[283][3] ,
         \mem[283][2] , \mem[283][1] , \mem[283][0] , \mem[282][7] ,
         \mem[282][6] , \mem[282][5] , \mem[282][4] , \mem[282][3] ,
         \mem[282][2] , \mem[282][1] , \mem[282][0] , \mem[281][7] ,
         \mem[281][6] , \mem[281][5] , \mem[281][4] , \mem[281][3] ,
         \mem[281][2] , \mem[281][1] , \mem[281][0] , \mem[280][7] ,
         \mem[280][6] , \mem[280][5] , \mem[280][4] , \mem[280][3] ,
         \mem[280][2] , \mem[280][1] , \mem[280][0] , \mem[279][7] ,
         \mem[279][6] , \mem[279][5] , \mem[279][4] , \mem[279][3] ,
         \mem[279][2] , \mem[279][1] , \mem[279][0] , \mem[278][7] ,
         \mem[278][6] , \mem[278][5] , \mem[278][4] , \mem[278][3] ,
         \mem[278][2] , \mem[278][1] , \mem[278][0] , \mem[277][7] ,
         \mem[277][6] , \mem[277][5] , \mem[277][4] , \mem[277][3] ,
         \mem[277][2] , \mem[277][1] , \mem[277][0] , \mem[276][7] ,
         \mem[276][6] , \mem[276][5] , \mem[276][4] , \mem[276][3] ,
         \mem[276][2] , \mem[276][1] , \mem[276][0] , \mem[275][7] ,
         \mem[275][6] , \mem[275][5] , \mem[275][4] , \mem[275][3] ,
         \mem[275][2] , \mem[275][1] , \mem[275][0] , \mem[274][7] ,
         \mem[274][6] , \mem[274][5] , \mem[274][4] , \mem[274][3] ,
         \mem[274][2] , \mem[274][1] , \mem[274][0] , \mem[273][7] ,
         \mem[273][6] , \mem[273][5] , \mem[273][4] , \mem[273][3] ,
         \mem[273][2] , \mem[273][1] , \mem[273][0] , \mem[272][7] ,
         \mem[272][6] , \mem[272][5] , \mem[272][4] , \mem[272][3] ,
         \mem[272][2] , \mem[272][1] , \mem[272][0] , \mem[271][7] ,
         \mem[271][6] , \mem[271][5] , \mem[271][4] , \mem[271][3] ,
         \mem[271][2] , \mem[271][1] , \mem[271][0] , \mem[270][7] ,
         \mem[270][6] , \mem[270][5] , \mem[270][4] , \mem[270][3] ,
         \mem[270][2] , \mem[270][1] , \mem[270][0] , \mem[269][7] ,
         \mem[269][6] , \mem[269][5] , \mem[269][4] , \mem[269][3] ,
         \mem[269][2] , \mem[269][1] , \mem[269][0] , \mem[268][7] ,
         \mem[268][6] , \mem[268][5] , \mem[268][4] , \mem[268][3] ,
         \mem[268][2] , \mem[268][1] , \mem[268][0] , \mem[267][7] ,
         \mem[267][6] , \mem[267][5] , \mem[267][4] , \mem[267][3] ,
         \mem[267][2] , \mem[267][1] , \mem[267][0] , \mem[266][7] ,
         \mem[266][6] , \mem[266][5] , \mem[266][4] , \mem[266][3] ,
         \mem[266][2] , \mem[266][1] , \mem[266][0] , \mem[265][7] ,
         \mem[265][6] , \mem[265][5] , \mem[265][4] , \mem[265][3] ,
         \mem[265][2] , \mem[265][1] , \mem[265][0] , \mem[264][7] ,
         \mem[264][6] , \mem[264][5] , \mem[264][4] , \mem[264][3] ,
         \mem[264][2] , \mem[264][1] , \mem[264][0] , \mem[263][7] ,
         \mem[263][6] , \mem[263][5] , \mem[263][4] , \mem[263][3] ,
         \mem[263][2] , \mem[263][1] , \mem[263][0] , \mem[262][7] ,
         \mem[262][6] , \mem[262][5] , \mem[262][4] , \mem[262][3] ,
         \mem[262][2] , \mem[262][1] , \mem[262][0] , \mem[261][7] ,
         \mem[261][6] , \mem[261][5] , \mem[261][4] , \mem[261][3] ,
         \mem[261][2] , \mem[261][1] , \mem[261][0] , \mem[260][7] ,
         \mem[260][6] , \mem[260][5] , \mem[260][4] , \mem[260][3] ,
         \mem[260][2] , \mem[260][1] , \mem[260][0] , \mem[259][7] ,
         \mem[259][6] , \mem[259][5] , \mem[259][4] , \mem[259][3] ,
         \mem[259][2] , \mem[259][1] , \mem[259][0] , \mem[258][7] ,
         \mem[258][6] , \mem[258][5] , \mem[258][4] , \mem[258][3] ,
         \mem[258][2] , \mem[258][1] , \mem[258][0] , \mem[257][7] ,
         \mem[257][6] , \mem[257][5] , \mem[257][4] , \mem[257][3] ,
         \mem[257][2] , \mem[257][1] , \mem[257][0] , \mem[256][7] ,
         \mem[256][6] , \mem[256][5] , \mem[256][4] , \mem[256][3] ,
         \mem[256][2] , \mem[256][1] , \mem[256][0] , \mem[255][7] ,
         \mem[255][6] , \mem[255][5] , \mem[255][4] , \mem[255][3] ,
         \mem[255][2] , \mem[255][1] , \mem[255][0] , \mem[254][7] ,
         \mem[254][6] , \mem[254][5] , \mem[254][4] , \mem[254][3] ,
         \mem[254][2] , \mem[254][1] , \mem[254][0] , \mem[253][7] ,
         \mem[253][6] , \mem[253][5] , \mem[253][4] , \mem[253][3] ,
         \mem[253][2] , \mem[253][1] , \mem[253][0] , \mem[252][7] ,
         \mem[252][6] , \mem[252][5] , \mem[252][4] , \mem[252][3] ,
         \mem[252][2] , \mem[252][1] , \mem[252][0] , \mem[251][7] ,
         \mem[251][6] , \mem[251][5] , \mem[251][4] , \mem[251][3] ,
         \mem[251][2] , \mem[251][1] , \mem[251][0] , \mem[250][7] ,
         \mem[250][6] , \mem[250][5] , \mem[250][4] , \mem[250][3] ,
         \mem[250][2] , \mem[250][1] , \mem[250][0] , \mem[249][7] ,
         \mem[249][6] , \mem[249][5] , \mem[249][4] , \mem[249][3] ,
         \mem[249][2] , \mem[249][1] , \mem[249][0] , \mem[248][7] ,
         \mem[248][6] , \mem[248][5] , \mem[248][4] , \mem[248][3] ,
         \mem[248][2] , \mem[248][1] , \mem[248][0] , \mem[247][7] ,
         \mem[247][6] , \mem[247][5] , \mem[247][4] , \mem[247][3] ,
         \mem[247][2] , \mem[247][1] , \mem[247][0] , \mem[246][7] ,
         \mem[246][6] , \mem[246][5] , \mem[246][4] , \mem[246][3] ,
         \mem[246][2] , \mem[246][1] , \mem[246][0] , \mem[245][7] ,
         \mem[245][6] , \mem[245][5] , \mem[245][4] , \mem[245][3] ,
         \mem[245][2] , \mem[245][1] , \mem[245][0] , \mem[244][7] ,
         \mem[244][6] , \mem[244][5] , \mem[244][4] , \mem[244][3] ,
         \mem[244][2] , \mem[244][1] , \mem[244][0] , \mem[243][7] ,
         \mem[243][6] , \mem[243][5] , \mem[243][4] , \mem[243][3] ,
         \mem[243][2] , \mem[243][1] , \mem[243][0] , \mem[242][7] ,
         \mem[242][6] , \mem[242][5] , \mem[242][4] , \mem[242][3] ,
         \mem[242][2] , \mem[242][1] , \mem[242][0] , \mem[241][7] ,
         \mem[241][6] , \mem[241][5] , \mem[241][4] , \mem[241][3] ,
         \mem[241][2] , \mem[241][1] , \mem[241][0] , \mem[240][7] ,
         \mem[240][6] , \mem[240][5] , \mem[240][4] , \mem[240][3] ,
         \mem[240][2] , \mem[240][1] , \mem[240][0] , \mem[239][7] ,
         \mem[239][6] , \mem[239][5] , \mem[239][4] , \mem[239][3] ,
         \mem[239][2] , \mem[239][1] , \mem[239][0] , \mem[238][7] ,
         \mem[238][6] , \mem[238][5] , \mem[238][4] , \mem[238][3] ,
         \mem[238][2] , \mem[238][1] , \mem[238][0] , \mem[237][7] ,
         \mem[237][6] , \mem[237][5] , \mem[237][4] , \mem[237][3] ,
         \mem[237][2] , \mem[237][1] , \mem[237][0] , \mem[236][7] ,
         \mem[236][6] , \mem[236][5] , \mem[236][4] , \mem[236][3] ,
         \mem[236][2] , \mem[236][1] , \mem[236][0] , \mem[235][7] ,
         \mem[235][6] , \mem[235][5] , \mem[235][4] , \mem[235][3] ,
         \mem[235][2] , \mem[235][1] , \mem[235][0] , \mem[234][7] ,
         \mem[234][6] , \mem[234][5] , \mem[234][4] , \mem[234][3] ,
         \mem[234][2] , \mem[234][1] , \mem[234][0] , \mem[233][7] ,
         \mem[233][6] , \mem[233][5] , \mem[233][4] , \mem[233][3] ,
         \mem[233][2] , \mem[233][1] , \mem[233][0] , \mem[232][7] ,
         \mem[232][6] , \mem[232][5] , \mem[232][4] , \mem[232][3] ,
         \mem[232][2] , \mem[232][1] , \mem[232][0] , \mem[231][7] ,
         \mem[231][6] , \mem[231][5] , \mem[231][4] , \mem[231][3] ,
         \mem[231][2] , \mem[231][1] , \mem[231][0] , \mem[230][7] ,
         \mem[230][6] , \mem[230][5] , \mem[230][4] , \mem[230][3] ,
         \mem[230][2] , \mem[230][1] , \mem[230][0] , \mem[229][7] ,
         \mem[229][6] , \mem[229][5] , \mem[229][4] , \mem[229][3] ,
         \mem[229][2] , \mem[229][1] , \mem[229][0] , \mem[228][7] ,
         \mem[228][6] , \mem[228][5] , \mem[228][4] , \mem[228][3] ,
         \mem[228][2] , \mem[228][1] , \mem[228][0] , \mem[227][7] ,
         \mem[227][6] , \mem[227][5] , \mem[227][4] , \mem[227][3] ,
         \mem[227][2] , \mem[227][1] , \mem[227][0] , \mem[226][7] ,
         \mem[226][6] , \mem[226][5] , \mem[226][4] , \mem[226][3] ,
         \mem[226][2] , \mem[226][1] , \mem[226][0] , \mem[225][7] ,
         \mem[225][6] , \mem[225][5] , \mem[225][4] , \mem[225][3] ,
         \mem[225][2] , \mem[225][1] , \mem[225][0] , \mem[224][7] ,
         \mem[224][6] , \mem[224][5] , \mem[224][4] , \mem[224][3] ,
         \mem[224][2] , \mem[224][1] , \mem[224][0] , \mem[223][7] ,
         \mem[223][6] , \mem[223][5] , \mem[223][4] , \mem[223][3] ,
         \mem[223][2] , \mem[223][1] , \mem[223][0] , \mem[222][7] ,
         \mem[222][6] , \mem[222][5] , \mem[222][4] , \mem[222][3] ,
         \mem[222][2] , \mem[222][1] , \mem[222][0] , \mem[221][7] ,
         \mem[221][6] , \mem[221][5] , \mem[221][4] , \mem[221][3] ,
         \mem[221][2] , \mem[221][1] , \mem[221][0] , \mem[220][7] ,
         \mem[220][6] , \mem[220][5] , \mem[220][4] , \mem[220][3] ,
         \mem[220][2] , \mem[220][1] , \mem[220][0] , \mem[219][7] ,
         \mem[219][6] , \mem[219][5] , \mem[219][4] , \mem[219][3] ,
         \mem[219][2] , \mem[219][1] , \mem[219][0] , \mem[218][7] ,
         \mem[218][6] , \mem[218][5] , \mem[218][4] , \mem[218][3] ,
         \mem[218][2] , \mem[218][1] , \mem[218][0] , \mem[217][7] ,
         \mem[217][6] , \mem[217][5] , \mem[217][4] , \mem[217][3] ,
         \mem[217][2] , \mem[217][1] , \mem[217][0] , \mem[216][7] ,
         \mem[216][6] , \mem[216][5] , \mem[216][4] , \mem[216][3] ,
         \mem[216][2] , \mem[216][1] , \mem[216][0] , \mem[215][7] ,
         \mem[215][6] , \mem[215][5] , \mem[215][4] , \mem[215][3] ,
         \mem[215][2] , \mem[215][1] , \mem[215][0] , \mem[214][7] ,
         \mem[214][6] , \mem[214][5] , \mem[214][4] , \mem[214][3] ,
         \mem[214][2] , \mem[214][1] , \mem[214][0] , \mem[213][7] ,
         \mem[213][6] , \mem[213][5] , \mem[213][4] , \mem[213][3] ,
         \mem[213][2] , \mem[213][1] , \mem[213][0] , \mem[212][7] ,
         \mem[212][6] , \mem[212][5] , \mem[212][4] , \mem[212][3] ,
         \mem[212][2] , \mem[212][1] , \mem[212][0] , \mem[211][7] ,
         \mem[211][6] , \mem[211][5] , \mem[211][4] , \mem[211][3] ,
         \mem[211][2] , \mem[211][1] , \mem[211][0] , \mem[210][7] ,
         \mem[210][6] , \mem[210][5] , \mem[210][4] , \mem[210][3] ,
         \mem[210][2] , \mem[210][1] , \mem[210][0] , \mem[209][7] ,
         \mem[209][6] , \mem[209][5] , \mem[209][4] , \mem[209][3] ,
         \mem[209][2] , \mem[209][1] , \mem[209][0] , \mem[208][7] ,
         \mem[208][6] , \mem[208][5] , \mem[208][4] , \mem[208][3] ,
         \mem[208][2] , \mem[208][1] , \mem[208][0] , \mem[207][7] ,
         \mem[207][6] , \mem[207][5] , \mem[207][4] , \mem[207][3] ,
         \mem[207][2] , \mem[207][1] , \mem[207][0] , \mem[206][7] ,
         \mem[206][6] , \mem[206][5] , \mem[206][4] , \mem[206][3] ,
         \mem[206][2] , \mem[206][1] , \mem[206][0] , \mem[205][7] ,
         \mem[205][6] , \mem[205][5] , \mem[205][4] , \mem[205][3] ,
         \mem[205][2] , \mem[205][1] , \mem[205][0] , \mem[204][7] ,
         \mem[204][6] , \mem[204][5] , \mem[204][4] , \mem[204][3] ,
         \mem[204][2] , \mem[204][1] , \mem[204][0] , \mem[203][7] ,
         \mem[203][6] , \mem[203][5] , \mem[203][4] , \mem[203][3] ,
         \mem[203][2] , \mem[203][1] , \mem[203][0] , \mem[202][7] ,
         \mem[202][6] , \mem[202][5] , \mem[202][4] , \mem[202][3] ,
         \mem[202][2] , \mem[202][1] , \mem[202][0] , \mem[201][7] ,
         \mem[201][6] , \mem[201][5] , \mem[201][4] , \mem[201][3] ,
         \mem[201][2] , \mem[201][1] , \mem[201][0] , \mem[200][7] ,
         \mem[200][6] , \mem[200][5] , \mem[200][4] , \mem[200][3] ,
         \mem[200][2] , \mem[200][1] , \mem[200][0] , \mem[199][7] ,
         \mem[199][6] , \mem[199][5] , \mem[199][4] , \mem[199][3] ,
         \mem[199][2] , \mem[199][1] , \mem[199][0] , \mem[198][7] ,
         \mem[198][6] , \mem[198][5] , \mem[198][4] , \mem[198][3] ,
         \mem[198][2] , \mem[198][1] , \mem[198][0] , \mem[197][7] ,
         \mem[197][6] , \mem[197][5] , \mem[197][4] , \mem[197][3] ,
         \mem[197][2] , \mem[197][1] , \mem[197][0] , \mem[196][7] ,
         \mem[196][6] , \mem[196][5] , \mem[196][4] , \mem[196][3] ,
         \mem[196][2] , \mem[196][1] , \mem[196][0] , \mem[195][7] ,
         \mem[195][6] , \mem[195][5] , \mem[195][4] , \mem[195][3] ,
         \mem[195][2] , \mem[195][1] , \mem[195][0] , \mem[194][7] ,
         \mem[194][6] , \mem[194][5] , \mem[194][4] , \mem[194][3] ,
         \mem[194][2] , \mem[194][1] , \mem[194][0] , \mem[193][7] ,
         \mem[193][6] , \mem[193][5] , \mem[193][4] , \mem[193][3] ,
         \mem[193][2] , \mem[193][1] , \mem[193][0] , \mem[192][7] ,
         \mem[192][6] , \mem[192][5] , \mem[192][4] , \mem[192][3] ,
         \mem[192][2] , \mem[192][1] , \mem[192][0] , \mem[191][7] ,
         \mem[191][6] , \mem[191][5] , \mem[191][4] , \mem[191][3] ,
         \mem[191][2] , \mem[191][1] , \mem[191][0] , \mem[190][7] ,
         \mem[190][6] , \mem[190][5] , \mem[190][4] , \mem[190][3] ,
         \mem[190][2] , \mem[190][1] , \mem[190][0] , \mem[189][7] ,
         \mem[189][6] , \mem[189][5] , \mem[189][4] , \mem[189][3] ,
         \mem[189][2] , \mem[189][1] , \mem[189][0] , \mem[188][7] ,
         \mem[188][6] , \mem[188][5] , \mem[188][4] , \mem[188][3] ,
         \mem[188][2] , \mem[188][1] , \mem[188][0] , \mem[187][7] ,
         \mem[187][6] , \mem[187][5] , \mem[187][4] , \mem[187][3] ,
         \mem[187][2] , \mem[187][1] , \mem[187][0] , \mem[186][7] ,
         \mem[186][6] , \mem[186][5] , \mem[186][4] , \mem[186][3] ,
         \mem[186][2] , \mem[186][1] , \mem[186][0] , \mem[185][7] ,
         \mem[185][6] , \mem[185][5] , \mem[185][4] , \mem[185][3] ,
         \mem[185][2] , \mem[185][1] , \mem[185][0] , \mem[184][7] ,
         \mem[184][6] , \mem[184][5] , \mem[184][4] , \mem[184][3] ,
         \mem[184][2] , \mem[184][1] , \mem[184][0] , \mem[183][7] ,
         \mem[183][6] , \mem[183][5] , \mem[183][4] , \mem[183][3] ,
         \mem[183][2] , \mem[183][1] , \mem[183][0] , \mem[182][7] ,
         \mem[182][6] , \mem[182][5] , \mem[182][4] , \mem[182][3] ,
         \mem[182][2] , \mem[182][1] , \mem[182][0] , \mem[181][7] ,
         \mem[181][6] , \mem[181][5] , \mem[181][4] , \mem[181][3] ,
         \mem[181][2] , \mem[181][1] , \mem[181][0] , \mem[180][7] ,
         \mem[180][6] , \mem[180][5] , \mem[180][4] , \mem[180][3] ,
         \mem[180][2] , \mem[180][1] , \mem[180][0] , \mem[179][7] ,
         \mem[179][6] , \mem[179][5] , \mem[179][4] , \mem[179][3] ,
         \mem[179][2] , \mem[179][1] , \mem[179][0] , \mem[178][7] ,
         \mem[178][6] , \mem[178][5] , \mem[178][4] , \mem[178][3] ,
         \mem[178][2] , \mem[178][1] , \mem[178][0] , \mem[177][7] ,
         \mem[177][6] , \mem[177][5] , \mem[177][4] , \mem[177][3] ,
         \mem[177][2] , \mem[177][1] , \mem[177][0] , \mem[176][7] ,
         \mem[176][6] , \mem[176][5] , \mem[176][4] , \mem[176][3] ,
         \mem[176][2] , \mem[176][1] , \mem[176][0] , \mem[175][7] ,
         \mem[175][6] , \mem[175][5] , \mem[175][4] , \mem[175][3] ,
         \mem[175][2] , \mem[175][1] , \mem[175][0] , \mem[174][7] ,
         \mem[174][6] , \mem[174][5] , \mem[174][4] , \mem[174][3] ,
         \mem[174][2] , \mem[174][1] , \mem[174][0] , \mem[173][7] ,
         \mem[173][6] , \mem[173][5] , \mem[173][4] , \mem[173][3] ,
         \mem[173][2] , \mem[173][1] , \mem[173][0] , \mem[172][7] ,
         \mem[172][6] , \mem[172][5] , \mem[172][4] , \mem[172][3] ,
         \mem[172][2] , \mem[172][1] , \mem[172][0] , \mem[171][7] ,
         \mem[171][6] , \mem[171][5] , \mem[171][4] , \mem[171][3] ,
         \mem[171][2] , \mem[171][1] , \mem[171][0] , \mem[170][7] ,
         \mem[170][6] , \mem[170][5] , \mem[170][4] , \mem[170][3] ,
         \mem[170][2] , \mem[170][1] , \mem[170][0] , \mem[169][7] ,
         \mem[169][6] , \mem[169][5] , \mem[169][4] , \mem[169][3] ,
         \mem[169][2] , \mem[169][1] , \mem[169][0] , \mem[168][7] ,
         \mem[168][6] , \mem[168][5] , \mem[168][4] , \mem[168][3] ,
         \mem[168][2] , \mem[168][1] , \mem[168][0] , \mem[167][7] ,
         \mem[167][6] , \mem[167][5] , \mem[167][4] , \mem[167][3] ,
         \mem[167][2] , \mem[167][1] , \mem[167][0] , \mem[166][7] ,
         \mem[166][6] , \mem[166][5] , \mem[166][4] , \mem[166][3] ,
         \mem[166][2] , \mem[166][1] , \mem[166][0] , \mem[165][7] ,
         \mem[165][6] , \mem[165][5] , \mem[165][4] , \mem[165][3] ,
         \mem[165][2] , \mem[165][1] , \mem[165][0] , \mem[164][7] ,
         \mem[164][6] , \mem[164][5] , \mem[164][4] , \mem[164][3] ,
         \mem[164][2] , \mem[164][1] , \mem[164][0] , \mem[163][7] ,
         \mem[163][6] , \mem[163][5] , \mem[163][4] , \mem[163][3] ,
         \mem[163][2] , \mem[163][1] , \mem[163][0] , \mem[162][7] ,
         \mem[162][6] , \mem[162][5] , \mem[162][4] , \mem[162][3] ,
         \mem[162][2] , \mem[162][1] , \mem[162][0] , \mem[161][7] ,
         \mem[161][6] , \mem[161][5] , \mem[161][4] , \mem[161][3] ,
         \mem[161][2] , \mem[161][1] , \mem[161][0] , \mem[160][7] ,
         \mem[160][6] , \mem[160][5] , \mem[160][4] , \mem[160][3] ,
         \mem[160][2] , \mem[160][1] , \mem[160][0] , \mem[159][7] ,
         \mem[159][6] , \mem[159][5] , \mem[159][4] , \mem[159][3] ,
         \mem[159][2] , \mem[159][1] , \mem[159][0] , \mem[158][7] ,
         \mem[158][6] , \mem[158][5] , \mem[158][4] , \mem[158][3] ,
         \mem[158][2] , \mem[158][1] , \mem[158][0] , \mem[157][7] ,
         \mem[157][6] , \mem[157][5] , \mem[157][4] , \mem[157][3] ,
         \mem[157][2] , \mem[157][1] , \mem[157][0] , \mem[156][7] ,
         \mem[156][6] , \mem[156][5] , \mem[156][4] , \mem[156][3] ,
         \mem[156][2] , \mem[156][1] , \mem[156][0] , \mem[155][7] ,
         \mem[155][6] , \mem[155][5] , \mem[155][4] , \mem[155][3] ,
         \mem[155][2] , \mem[155][1] , \mem[155][0] , \mem[154][7] ,
         \mem[154][6] , \mem[154][5] , \mem[154][4] , \mem[154][3] ,
         \mem[154][2] , \mem[154][1] , \mem[154][0] , \mem[153][7] ,
         \mem[153][6] , \mem[153][5] , \mem[153][4] , \mem[153][3] ,
         \mem[153][2] , \mem[153][1] , \mem[153][0] , \mem[152][7] ,
         \mem[152][6] , \mem[152][5] , \mem[152][4] , \mem[152][3] ,
         \mem[152][2] , \mem[152][1] , \mem[152][0] , \mem[151][7] ,
         \mem[151][6] , \mem[151][5] , \mem[151][4] , \mem[151][3] ,
         \mem[151][2] , \mem[151][1] , \mem[151][0] , \mem[150][7] ,
         \mem[150][6] , \mem[150][5] , \mem[150][4] , \mem[150][3] ,
         \mem[150][2] , \mem[150][1] , \mem[150][0] , \mem[149][7] ,
         \mem[149][6] , \mem[149][5] , \mem[149][4] , \mem[149][3] ,
         \mem[149][2] , \mem[149][1] , \mem[149][0] , \mem[148][7] ,
         \mem[148][6] , \mem[148][5] , \mem[148][4] , \mem[148][3] ,
         \mem[148][2] , \mem[148][1] , \mem[148][0] , \mem[147][7] ,
         \mem[147][6] , \mem[147][5] , \mem[147][4] , \mem[147][3] ,
         \mem[147][2] , \mem[147][1] , \mem[147][0] , \mem[146][7] ,
         \mem[146][6] , \mem[146][5] , \mem[146][4] , \mem[146][3] ,
         \mem[146][2] , \mem[146][1] , \mem[146][0] , \mem[145][7] ,
         \mem[145][6] , \mem[145][5] , \mem[145][4] , \mem[145][3] ,
         \mem[145][2] , \mem[145][1] , \mem[145][0] , \mem[144][7] ,
         \mem[144][6] , \mem[144][5] , \mem[144][4] , \mem[144][3] ,
         \mem[144][2] , \mem[144][1] , \mem[144][0] , \mem[143][7] ,
         \mem[143][6] , \mem[143][5] , \mem[143][4] , \mem[143][3] ,
         \mem[143][2] , \mem[143][1] , \mem[143][0] , \mem[142][7] ,
         \mem[142][6] , \mem[142][5] , \mem[142][4] , \mem[142][3] ,
         \mem[142][2] , \mem[142][1] , \mem[142][0] , \mem[141][7] ,
         \mem[141][6] , \mem[141][5] , \mem[141][4] , \mem[141][3] ,
         \mem[141][2] , \mem[141][1] , \mem[141][0] , \mem[140][7] ,
         \mem[140][6] , \mem[140][5] , \mem[140][4] , \mem[140][3] ,
         \mem[140][2] , \mem[140][1] , \mem[140][0] , \mem[139][7] ,
         \mem[139][6] , \mem[139][5] , \mem[139][4] , \mem[139][3] ,
         \mem[139][2] , \mem[139][1] , \mem[139][0] , \mem[138][7] ,
         \mem[138][6] , \mem[138][5] , \mem[138][4] , \mem[138][3] ,
         \mem[138][2] , \mem[138][1] , \mem[138][0] , \mem[137][7] ,
         \mem[137][6] , \mem[137][5] , \mem[137][4] , \mem[137][3] ,
         \mem[137][2] , \mem[137][1] , \mem[137][0] , \mem[136][7] ,
         \mem[136][6] , \mem[136][5] , \mem[136][4] , \mem[136][3] ,
         \mem[136][2] , \mem[136][1] , \mem[136][0] , \mem[135][7] ,
         \mem[135][6] , \mem[135][5] , \mem[135][4] , \mem[135][3] ,
         \mem[135][2] , \mem[135][1] , \mem[135][0] , \mem[134][7] ,
         \mem[134][6] , \mem[134][5] , \mem[134][4] , \mem[134][3] ,
         \mem[134][2] , \mem[134][1] , \mem[134][0] , \mem[133][7] ,
         \mem[133][6] , \mem[133][5] , \mem[133][4] , \mem[133][3] ,
         \mem[133][2] , \mem[133][1] , \mem[133][0] , \mem[132][7] ,
         \mem[132][6] , \mem[132][5] , \mem[132][4] , \mem[132][3] ,
         \mem[132][2] , \mem[132][1] , \mem[132][0] , \mem[131][7] ,
         \mem[131][6] , \mem[131][5] , \mem[131][4] , \mem[131][3] ,
         \mem[131][2] , \mem[131][1] , \mem[131][0] , \mem[130][7] ,
         \mem[130][6] , \mem[130][5] , \mem[130][4] , \mem[130][3] ,
         \mem[130][2] , \mem[130][1] , \mem[130][0] , \mem[129][7] ,
         \mem[129][6] , \mem[129][5] , \mem[129][4] , \mem[129][3] ,
         \mem[129][2] , \mem[129][1] , \mem[129][0] , \mem[128][7] ,
         \mem[128][6] , \mem[128][5] , \mem[128][4] , \mem[128][3] ,
         \mem[128][2] , \mem[128][1] , \mem[128][0] , \mem[127][7] ,
         \mem[127][6] , \mem[127][5] , \mem[127][4] , \mem[127][3] ,
         \mem[127][2] , \mem[127][1] , \mem[127][0] , \mem[126][7] ,
         \mem[126][6] , \mem[126][5] , \mem[126][4] , \mem[126][3] ,
         \mem[126][2] , \mem[126][1] , \mem[126][0] , \mem[125][7] ,
         \mem[125][6] , \mem[125][5] , \mem[125][4] , \mem[125][3] ,
         \mem[125][2] , \mem[125][1] , \mem[125][0] , \mem[124][7] ,
         \mem[124][6] , \mem[124][5] , \mem[124][4] , \mem[124][3] ,
         \mem[124][2] , \mem[124][1] , \mem[124][0] , \mem[123][7] ,
         \mem[123][6] , \mem[123][5] , \mem[123][4] , \mem[123][3] ,
         \mem[123][2] , \mem[123][1] , \mem[123][0] , \mem[122][7] ,
         \mem[122][6] , \mem[122][5] , \mem[122][4] , \mem[122][3] ,
         \mem[122][2] , \mem[122][1] , \mem[122][0] , \mem[121][7] ,
         \mem[121][6] , \mem[121][5] , \mem[121][4] , \mem[121][3] ,
         \mem[121][2] , \mem[121][1] , \mem[121][0] , \mem[120][7] ,
         \mem[120][6] , \mem[120][5] , \mem[120][4] , \mem[120][3] ,
         \mem[120][2] , \mem[120][1] , \mem[120][0] , \mem[119][7] ,
         \mem[119][6] , \mem[119][5] , \mem[119][4] , \mem[119][3] ,
         \mem[119][2] , \mem[119][1] , \mem[119][0] , \mem[118][7] ,
         \mem[118][6] , \mem[118][5] , \mem[118][4] , \mem[118][3] ,
         \mem[118][2] , \mem[118][1] , \mem[118][0] , \mem[117][7] ,
         \mem[117][6] , \mem[117][5] , \mem[117][4] , \mem[117][3] ,
         \mem[117][2] , \mem[117][1] , \mem[117][0] , \mem[116][7] ,
         \mem[116][6] , \mem[116][5] , \mem[116][4] , \mem[116][3] ,
         \mem[116][2] , \mem[116][1] , \mem[116][0] , \mem[115][7] ,
         \mem[115][6] , \mem[115][5] , \mem[115][4] , \mem[115][3] ,
         \mem[115][2] , \mem[115][1] , \mem[115][0] , \mem[114][7] ,
         \mem[114][6] , \mem[114][5] , \mem[114][4] , \mem[114][3] ,
         \mem[114][2] , \mem[114][1] , \mem[114][0] , \mem[113][7] ,
         \mem[113][6] , \mem[113][5] , \mem[113][4] , \mem[113][3] ,
         \mem[113][2] , \mem[113][1] , \mem[113][0] , \mem[112][7] ,
         \mem[112][6] , \mem[112][5] , \mem[112][4] , \mem[112][3] ,
         \mem[112][2] , \mem[112][1] , \mem[112][0] , \mem[111][7] ,
         \mem[111][6] , \mem[111][5] , \mem[111][4] , \mem[111][3] ,
         \mem[111][2] , \mem[111][1] , \mem[111][0] , \mem[110][7] ,
         \mem[110][6] , \mem[110][5] , \mem[110][4] , \mem[110][3] ,
         \mem[110][2] , \mem[110][1] , \mem[110][0] , \mem[109][7] ,
         \mem[109][6] , \mem[109][5] , \mem[109][4] , \mem[109][3] ,
         \mem[109][2] , \mem[109][1] , \mem[109][0] , \mem[108][7] ,
         \mem[108][6] , \mem[108][5] , \mem[108][4] , \mem[108][3] ,
         \mem[108][2] , \mem[108][1] , \mem[108][0] , \mem[107][7] ,
         \mem[107][6] , \mem[107][5] , \mem[107][4] , \mem[107][3] ,
         \mem[107][2] , \mem[107][1] , \mem[107][0] , \mem[106][7] ,
         \mem[106][6] , \mem[106][5] , \mem[106][4] , \mem[106][3] ,
         \mem[106][2] , \mem[106][1] , \mem[106][0] , \mem[105][7] ,
         \mem[105][6] , \mem[105][5] , \mem[105][4] , \mem[105][3] ,
         \mem[105][2] , \mem[105][1] , \mem[105][0] , \mem[104][7] ,
         \mem[104][6] , \mem[104][5] , \mem[104][4] , \mem[104][3] ,
         \mem[104][2] , \mem[104][1] , \mem[104][0] , \mem[103][7] ,
         \mem[103][6] , \mem[103][5] , \mem[103][4] , \mem[103][3] ,
         \mem[103][2] , \mem[103][1] , \mem[103][0] , \mem[102][7] ,
         \mem[102][6] , \mem[102][5] , \mem[102][4] , \mem[102][3] ,
         \mem[102][2] , \mem[102][1] , \mem[102][0] , \mem[101][7] ,
         \mem[101][6] , \mem[101][5] , \mem[101][4] , \mem[101][3] ,
         \mem[101][2] , \mem[101][1] , \mem[101][0] , \mem[100][7] ,
         \mem[100][6] , \mem[100][5] , \mem[100][4] , \mem[100][3] ,
         \mem[100][2] , \mem[100][1] , \mem[100][0] , \mem[99][7] ,
         \mem[99][6] , \mem[99][5] , \mem[99][4] , \mem[99][3] , \mem[99][2] ,
         \mem[99][1] , \mem[99][0] , \mem[98][7] , \mem[98][6] , \mem[98][5] ,
         \mem[98][4] , \mem[98][3] , \mem[98][2] , \mem[98][1] , \mem[98][0] ,
         \mem[97][7] , \mem[97][6] , \mem[97][5] , \mem[97][4] , \mem[97][3] ,
         \mem[97][2] , \mem[97][1] , \mem[97][0] , \mem[96][7] , \mem[96][6] ,
         \mem[96][5] , \mem[96][4] , \mem[96][3] , \mem[96][2] , \mem[96][1] ,
         \mem[96][0] , \mem[95][7] , \mem[95][6] , \mem[95][5] , \mem[95][4] ,
         \mem[95][3] , \mem[95][2] , \mem[95][1] , \mem[95][0] , \mem[94][7] ,
         \mem[94][6] , \mem[94][5] , \mem[94][4] , \mem[94][3] , \mem[94][2] ,
         \mem[94][1] , \mem[94][0] , \mem[93][7] , \mem[93][6] , \mem[93][5] ,
         \mem[93][4] , \mem[93][3] , \mem[93][2] , \mem[93][1] , \mem[93][0] ,
         \mem[92][7] , \mem[92][6] , \mem[92][5] , \mem[92][4] , \mem[92][3] ,
         \mem[92][2] , \mem[92][1] , \mem[92][0] , \mem[91][7] , \mem[91][6] ,
         \mem[91][5] , \mem[91][4] , \mem[91][3] , \mem[91][2] , \mem[91][1] ,
         \mem[91][0] , \mem[90][7] , \mem[90][6] , \mem[90][5] , \mem[90][4] ,
         \mem[90][3] , \mem[90][2] , \mem[90][1] , \mem[90][0] , \mem[89][7] ,
         \mem[89][6] , \mem[89][5] , \mem[89][4] , \mem[89][3] , \mem[89][2] ,
         \mem[89][1] , \mem[89][0] , \mem[88][7] , \mem[88][6] , \mem[88][5] ,
         \mem[88][4] , \mem[88][3] , \mem[88][2] , \mem[88][1] , \mem[88][0] ,
         \mem[87][7] , \mem[87][6] , \mem[87][5] , \mem[87][4] , \mem[87][3] ,
         \mem[87][2] , \mem[87][1] , \mem[87][0] , \mem[86][7] , \mem[86][6] ,
         \mem[86][5] , \mem[86][4] , \mem[86][3] , \mem[86][2] , \mem[86][1] ,
         \mem[86][0] , \mem[85][7] , \mem[85][6] , \mem[85][5] , \mem[85][4] ,
         \mem[85][3] , \mem[85][2] , \mem[85][1] , \mem[85][0] , \mem[84][7] ,
         \mem[84][6] , \mem[84][5] , \mem[84][4] , \mem[84][3] , \mem[84][2] ,
         \mem[84][1] , \mem[84][0] , \mem[83][7] , \mem[83][6] , \mem[83][5] ,
         \mem[83][4] , \mem[83][3] , \mem[83][2] , \mem[83][1] , \mem[83][0] ,
         \mem[82][7] , \mem[82][6] , \mem[82][5] , \mem[82][4] , \mem[82][3] ,
         \mem[82][2] , \mem[82][1] , \mem[82][0] , \mem[81][7] , \mem[81][6] ,
         \mem[81][5] , \mem[81][4] , \mem[81][3] , \mem[81][2] , \mem[81][1] ,
         \mem[81][0] , \mem[80][7] , \mem[80][6] , \mem[80][5] , \mem[80][4] ,
         \mem[80][3] , \mem[80][2] , \mem[80][1] , \mem[80][0] , \mem[79][7] ,
         \mem[79][6] , \mem[79][5] , \mem[79][4] , \mem[79][3] , \mem[79][2] ,
         \mem[79][1] , \mem[79][0] , \mem[78][7] , \mem[78][6] , \mem[78][5] ,
         \mem[78][4] , \mem[78][3] , \mem[78][2] , \mem[78][1] , \mem[78][0] ,
         \mem[77][7] , \mem[77][6] , \mem[77][5] , \mem[77][4] , \mem[77][3] ,
         \mem[77][2] , \mem[77][1] , \mem[77][0] , \mem[76][7] , \mem[76][6] ,
         \mem[76][5] , \mem[76][4] , \mem[76][3] , \mem[76][2] , \mem[76][1] ,
         \mem[76][0] , \mem[75][7] , \mem[75][6] , \mem[75][5] , \mem[75][4] ,
         \mem[75][3] , \mem[75][2] , \mem[75][1] , \mem[75][0] , \mem[74][7] ,
         \mem[74][6] , \mem[74][5] , \mem[74][4] , \mem[74][3] , \mem[74][2] ,
         \mem[74][1] , \mem[74][0] , \mem[73][7] , \mem[73][6] , \mem[73][5] ,
         \mem[73][4] , \mem[73][3] , \mem[73][2] , \mem[73][1] , \mem[73][0] ,
         \mem[72][7] , \mem[72][6] , \mem[72][5] , \mem[72][4] , \mem[72][3] ,
         \mem[72][2] , \mem[72][1] , \mem[72][0] , \mem[71][7] , \mem[71][6] ,
         \mem[71][5] , \mem[71][4] , \mem[71][3] , \mem[71][2] , \mem[71][1] ,
         \mem[71][0] , \mem[70][7] , \mem[70][6] , \mem[70][5] , \mem[70][4] ,
         \mem[70][3] , \mem[70][2] , \mem[70][1] , \mem[70][0] , \mem[69][7] ,
         \mem[69][6] , \mem[69][5] , \mem[69][4] , \mem[69][3] , \mem[69][2] ,
         \mem[69][1] , \mem[69][0] , \mem[68][7] , \mem[68][6] , \mem[68][5] ,
         \mem[68][4] , \mem[68][3] , \mem[68][2] , \mem[68][1] , \mem[68][0] ,
         \mem[67][7] , \mem[67][6] , \mem[67][5] , \mem[67][4] , \mem[67][3] ,
         \mem[67][2] , \mem[67][1] , \mem[67][0] , \mem[66][7] , \mem[66][6] ,
         \mem[66][5] , \mem[66][4] , \mem[66][3] , \mem[66][2] , \mem[66][1] ,
         \mem[66][0] , \mem[65][7] , \mem[65][6] , \mem[65][5] , \mem[65][4] ,
         \mem[65][3] , \mem[65][2] , \mem[65][1] , \mem[65][0] , \mem[64][7] ,
         \mem[64][6] , \mem[64][5] , \mem[64][4] , \mem[64][3] , \mem[64][2] ,
         \mem[64][1] , \mem[64][0] , \mem[63][7] , \mem[63][6] , \mem[63][5] ,
         \mem[63][4] , \mem[63][3] , \mem[63][2] , \mem[63][1] , \mem[63][0] ,
         \mem[62][7] , \mem[62][6] , \mem[62][5] , \mem[62][4] , \mem[62][3] ,
         \mem[62][2] , \mem[62][1] , \mem[62][0] , \mem[61][7] , \mem[61][6] ,
         \mem[61][5] , \mem[61][4] , \mem[61][3] , \mem[61][2] , \mem[61][1] ,
         \mem[61][0] , \mem[60][7] , \mem[60][6] , \mem[60][5] , \mem[60][4] ,
         \mem[60][3] , \mem[60][2] , \mem[60][1] , \mem[60][0] , \mem[59][7] ,
         \mem[59][6] , \mem[59][5] , \mem[59][4] , \mem[59][3] , \mem[59][2] ,
         \mem[59][1] , \mem[59][0] , \mem[58][7] , \mem[58][6] , \mem[58][5] ,
         \mem[58][4] , \mem[58][3] , \mem[58][2] , \mem[58][1] , \mem[58][0] ,
         \mem[57][7] , \mem[57][6] , \mem[57][5] , \mem[57][4] , \mem[57][3] ,
         \mem[57][2] , \mem[57][1] , \mem[57][0] , \mem[56][7] , \mem[56][6] ,
         \mem[56][5] , \mem[56][4] , \mem[56][3] , \mem[56][2] , \mem[56][1] ,
         \mem[56][0] , \mem[55][7] , \mem[55][6] , \mem[55][5] , \mem[55][4] ,
         \mem[55][3] , \mem[55][2] , \mem[55][1] , \mem[55][0] , \mem[54][7] ,
         \mem[54][6] , \mem[54][5] , \mem[54][4] , \mem[54][3] , \mem[54][2] ,
         \mem[54][1] , \mem[54][0] , \mem[53][7] , \mem[53][6] , \mem[53][5] ,
         \mem[53][4] , \mem[53][3] , \mem[53][2] , \mem[53][1] , \mem[53][0] ,
         \mem[52][7] , \mem[52][6] , \mem[52][5] , \mem[52][4] , \mem[52][3] ,
         \mem[52][2] , \mem[52][1] , \mem[52][0] , \mem[51][7] , \mem[51][6] ,
         \mem[51][5] , \mem[51][4] , \mem[51][3] , \mem[51][2] , \mem[51][1] ,
         \mem[51][0] , \mem[50][7] , \mem[50][6] , \mem[50][5] , \mem[50][4] ,
         \mem[50][3] , \mem[50][2] , \mem[50][1] , \mem[50][0] , \mem[49][7] ,
         \mem[49][6] , \mem[49][5] , \mem[49][4] , \mem[49][3] , \mem[49][2] ,
         \mem[49][1] , \mem[49][0] , \mem[48][7] , \mem[48][6] , \mem[48][5] ,
         \mem[48][4] , \mem[48][3] , \mem[48][2] , \mem[48][1] , \mem[48][0] ,
         \mem[47][7] , \mem[47][6] , \mem[47][5] , \mem[47][4] , \mem[47][3] ,
         \mem[47][2] , \mem[47][1] , \mem[47][0] , \mem[46][7] , \mem[46][6] ,
         \mem[46][5] , \mem[46][4] , \mem[46][3] , \mem[46][2] , \mem[46][1] ,
         \mem[46][0] , \mem[45][7] , \mem[45][6] , \mem[45][5] , \mem[45][4] ,
         \mem[45][3] , \mem[45][2] , \mem[45][1] , \mem[45][0] , \mem[44][7] ,
         \mem[44][6] , \mem[44][5] , \mem[44][4] , \mem[44][3] , \mem[44][2] ,
         \mem[44][1] , \mem[44][0] , \mem[43][7] , \mem[43][6] , \mem[43][5] ,
         \mem[43][4] , \mem[43][3] , \mem[43][2] , \mem[43][1] , \mem[43][0] ,
         \mem[42][7] , \mem[42][6] , \mem[42][5] , \mem[42][4] , \mem[42][3] ,
         \mem[42][2] , \mem[42][1] , \mem[42][0] , \mem[41][7] , \mem[41][6] ,
         \mem[41][5] , \mem[41][4] , \mem[41][3] , \mem[41][2] , \mem[41][1] ,
         \mem[41][0] , \mem[40][7] , \mem[40][6] , \mem[40][5] , \mem[40][4] ,
         \mem[40][3] , \mem[40][2] , \mem[40][1] , \mem[40][0] , \mem[39][7] ,
         \mem[39][6] , \mem[39][5] , \mem[39][4] , \mem[39][3] , \mem[39][2] ,
         \mem[39][1] , \mem[39][0] , \mem[38][7] , \mem[38][6] , \mem[38][5] ,
         \mem[38][4] , \mem[38][3] , \mem[38][2] , \mem[38][1] , \mem[38][0] ,
         \mem[37][7] , \mem[37][6] , \mem[37][5] , \mem[37][4] , \mem[37][3] ,
         \mem[37][2] , \mem[37][1] , \mem[37][0] , \mem[36][7] , \mem[36][6] ,
         \mem[36][5] , \mem[36][4] , \mem[36][3] , \mem[36][2] , \mem[36][1] ,
         \mem[36][0] , \mem[35][7] , \mem[35][6] , \mem[35][5] , \mem[35][4] ,
         \mem[35][3] , \mem[35][2] , \mem[35][1] , \mem[35][0] , \mem[34][7] ,
         \mem[34][6] , \mem[34][5] , \mem[34][4] , \mem[34][3] , \mem[34][2] ,
         \mem[34][1] , \mem[34][0] , \mem[33][7] , \mem[33][6] , \mem[33][5] ,
         \mem[33][4] , \mem[33][3] , \mem[33][2] , \mem[33][1] , \mem[33][0] ,
         \mem[32][7] , \mem[32][6] , \mem[32][5] , \mem[32][4] , \mem[32][3] ,
         \mem[32][2] , \mem[32][1] , \mem[32][0] , \mem[31][7] , \mem[31][6] ,
         \mem[31][5] , \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] ,
         \mem[31][0] , \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] ,
         \mem[30][3] , \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] ,
         \mem[29][6] , \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] ,
         \mem[29][1] , \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] ,
         \mem[28][4] , \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] ,
         \mem[27][7] , \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] ,
         \mem[27][2] , \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] ,
         \mem[26][5] , \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] ,
         \mem[26][0] , \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] ,
         \mem[25][3] , \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] ,
         \mem[24][6] , \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] ,
         \mem[24][1] , \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] ,
         \mem[23][4] , \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] ,
         \mem[22][7] , \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] ,
         \mem[22][2] , \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] ,
         \mem[21][5] , \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] ,
         \mem[21][0] , \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] ,
         \mem[20][3] , \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] ,
         \mem[19][6] , \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] ,
         \mem[19][1] , \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] ,
         \mem[18][4] , \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] ,
         \mem[17][7] , \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] ,
         \mem[17][2] , \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] ,
         \mem[16][5] , \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] ,
         \mem[16][0] , \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] ,
         \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] ,
         \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] ,
         \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] ,
         \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] ,
         \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] ,
         \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] ,
         \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] ,
         \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] ,
         \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] ,
         \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] ,
         \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] ,
         \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] ,
         \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] ,
         \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] ,
         \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] ,
         \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] ,
         \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N28, N29, N30,
         N31, N32, N33, N34, N35, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
         n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,
         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,
         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
         n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,
         n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
         n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
         n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072,
         n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,
         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
         n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,
         n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
         n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
         n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144,
         n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
         n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,
         n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168,
         n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176,
         n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
         n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192,
         n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200,
         n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
         n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216,
         n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224,
         n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232,
         n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240,
         n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
         n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256,
         n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264,
         n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,
         n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,
         n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288,
         n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296,
         n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304,
         n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
         n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320,
         n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,
         n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336,
         n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344,
         n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
         n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360,
         n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368,
         n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
         n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,
         n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392,
         n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400,
         n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408,
         n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416,
         n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
         n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432,
         n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
         n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
         n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472,
         n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480,
         n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488,
         n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,
         n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504,
         n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512,
         n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520,
         n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528,
         n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536,
         n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544,
         n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552,
         n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560,
         n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,
         n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576,
         n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584,
         n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592,
         n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600,
         n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608,
         n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616,
         n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624,
         n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,
         n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
         n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648,
         n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656,
         n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664,
         n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672,
         n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680,
         n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688,
         n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696,
         n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704,
         n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712,
         n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720,
         n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728,
         n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736,
         n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744,
         n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752,
         n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760,
         n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768,
         n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776,
         n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,
         n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792,
         n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800,
         n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808,
         n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816,
         n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824,
         n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,
         n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840,
         n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848,
         n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,
         n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864,
         n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872,
         n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880,
         n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888,
         n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896,
         n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904,
         n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912,
         n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920,
         n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928,
         n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936,
         n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944,
         n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
         n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960,
         n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968,
         n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976,
         n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984,
         n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992,
         n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000,
         n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008,
         n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016,
         n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
         n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032,
         n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040,
         n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048,
         n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056,
         n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064,
         n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072,
         n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080,
         n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088,
         n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
         n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104,
         n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112,
         n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120,
         n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128,
         n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136,
         n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,
         n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152,
         n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160,
         n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
         n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176,
         n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184,
         n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192,
         n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200,
         n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208,
         n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,
         n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224,
         n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232,
         n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
         n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248,
         n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256,
         n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264,
         n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272,
         n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280,
         n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,
         n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296,
         n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304,
         n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,
         n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320,
         n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
         n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336,
         n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
         n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352,
         n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360,
         n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368,
         n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,
         n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384,
         n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392,
         n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400,
         n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408,
         n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416,
         n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424,
         n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432,
         n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440,
         n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448,
         n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456,
         n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464,
         n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472,
         n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480,
         n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488,
         n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496,
         n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504,
         n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512,
         n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520,
         n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528,
         n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536,
         n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544,
         n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552,
         n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560,
         n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568,
         n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576,
         n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584,
         n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592,
         n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600,
         n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608,
         n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616,
         n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624,
         n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632,
         n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640,
         n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648,
         n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656,
         n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664,
         n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672,
         n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680,
         n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688,
         n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696,
         n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704,
         n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712,
         n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720,
         n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728,
         n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736,
         n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744,
         n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752,
         n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760,
         n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768,
         n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776,
         n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784,
         n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792,
         n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800,
         n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808,
         n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816,
         n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824,
         n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832,
         n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840,
         n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848,
         n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856,
         n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864,
         n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872,
         n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880,
         n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888,
         n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896,
         n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904,
         n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912,
         n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920,
         n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928,
         n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936,
         n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944,
         n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952,
         n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960,
         n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968,
         n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976,
         n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984,
         n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992,
         n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000,
         n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008,
         n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016,
         n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024,
         n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032,
         n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040,
         n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048,
         n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056,
         n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064,
         n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072,
         n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080,
         n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088,
         n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096,
         n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104,
         n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112,
         n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120,
         n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128,
         n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136,
         n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144,
         n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152,
         n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160,
         n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168,
         n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176,
         n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184,
         n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192,
         n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200,
         n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208,
         n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216,
         n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224,
         n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232,
         n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240,
         n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248,
         n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256,
         n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264,
         n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272,
         n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280,
         n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288,
         n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296,
         n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304,
         n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312,
         n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320,
         n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328,
         n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336,
         n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344,
         n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352,
         n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360,
         n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368,
         n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376,
         n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384,
         n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392,
         n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400,
         n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408,
         n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416,
         n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424,
         n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432,
         n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440,
         n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448,
         n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456,
         n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464,
         n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472,
         n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480,
         n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488,
         n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496,
         n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504,
         n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512,
         n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520,
         n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528,
         n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536,
         n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544,
         n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552,
         n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560,
         n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568,
         n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576,
         n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584,
         n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592,
         n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600,
         n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608,
         n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616,
         n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624,
         n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632,
         n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640,
         n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648,
         n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656,
         n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664,
         n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672,
         n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680,
         n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688,
         n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696,
         n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704,
         n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712,
         n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720,
         n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728,
         n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736,
         n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744,
         n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752,
         n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760,
         n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768,
         n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776,
         n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784,
         n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792,
         n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800,
         n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808,
         n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816,
         n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824,
         n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832,
         n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840,
         n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848,
         n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856,
         n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864,
         n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872,
         n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880,
         n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888,
         n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896,
         n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904,
         n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912,
         n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920,
         n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928,
         n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936,
         n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944,
         n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952,
         n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960,
         n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968,
         n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976,
         n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984,
         n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992,
         n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000,
         n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008,
         n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016,
         n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024,
         n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032,
         n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040,
         n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048,
         n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056,
         n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064,
         n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072,
         n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080,
         n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088,
         n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096,
         n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104,
         n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112,
         n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120,
         n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128,
         n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136,
         n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144,
         n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152,
         n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160,
         n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168,
         n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176,
         n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184,
         n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192,
         n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200,
         n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208,
         n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216,
         n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224,
         n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232,
         n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240,
         n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248,
         n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256,
         n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264,
         n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272,
         n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280,
         n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288,
         n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296,
         n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304,
         n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312,
         n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320,
         n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328,
         n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336,
         n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344,
         n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352,
         n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360,
         n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368,
         n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376,
         n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384,
         n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392,
         n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400,
         n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408,
         n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416,
         n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424,
         n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432,
         n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440,
         n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448,
         n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456,
         n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464,
         n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472,
         n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480,
         n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488,
         n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496,
         n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504,
         n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512,
         n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520,
         n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528,
         n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536,
         n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544,
         n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552,
         n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560,
         n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568,
         n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576,
         n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584,
         n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592,
         n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600,
         n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608,
         n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616,
         n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624,
         n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632,
         n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640,
         n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648,
         n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656,
         n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664,
         n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672,
         n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680,
         n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688,
         n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696,
         n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704,
         n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712,
         n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720,
         n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728,
         n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736,
         n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744,
         n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752,
         n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760,
         n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768,
         n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776,
         n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784,
         n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792,
         n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800,
         n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808,
         n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816,
         n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824,
         n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832,
         n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840,
         n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848,
         n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856,
         n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864,
         n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872,
         n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880,
         n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888,
         n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896,
         n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904,
         n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912,
         n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920,
         n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928,
         n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936,
         n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944,
         n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952,
         n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960,
         n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968,
         n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976,
         n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984,
         n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992,
         n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000,
         n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008,
         n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016,
         n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024,
         n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032,
         n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040,
         n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048,
         n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056,
         n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064,
         n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072,
         n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080,
         n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088,
         n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,
         n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104,
         n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112,
         n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120,
         n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128,
         n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136,
         n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144,
         n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152,
         n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160,
         n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168,
         n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176,
         n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184,
         n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192,
         n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200,
         n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208,
         n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216,
         n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224,
         n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232,
         n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240,
         n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248,
         n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256,
         n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264,
         n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272,
         n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280,
         n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288,
         n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296,
         n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304,
         n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312,
         n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320,
         n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328,
         n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336,
         n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344,
         n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352,
         n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360,
         n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368,
         n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376,
         n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384,
         n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392,
         n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400,
         n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408,
         n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416,
         n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,
         n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432,
         n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440,
         n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448,
         n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456,
         n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464,
         n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472,
         n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480,
         n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488,
         n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496,
         n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504,
         n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512,
         n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520,
         n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528,
         n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536,
         n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544,
         n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552,
         n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560,
         n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568,
         n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576,
         n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584,
         n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592,
         n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600,
         n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608,
         n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616,
         n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624,
         n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632,
         n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640,
         n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648,
         n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656,
         n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664,
         n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672,
         n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680,
         n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688,
         n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696,
         n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704,
         n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712,
         n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720,
         n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728,
         n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736,
         n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744,
         n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752,
         n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760,
         n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768,
         n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776,
         n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784,
         n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792,
         n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800,
         n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808,
         n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816,
         n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824,
         n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832,
         n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840,
         n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848,
         n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856,
         n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864,
         n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872,
         n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880,
         n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888,
         n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896,
         n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904,
         n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912,
         n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920,
         n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928,
         n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936,
         n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944,
         n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952,
         n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960,
         n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968,
         n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976,
         n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984,
         n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992,
         n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000,
         n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008,
         n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016,
         n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024,
         n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032,
         n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040,
         n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048,
         n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056,
         n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064,
         n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072,
         n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080,
         n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088,
         n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096,
         n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104,
         n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112,
         n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120,
         n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128,
         n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136,
         n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144,
         n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152,
         n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160,
         n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168,
         n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176,
         n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184,
         n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192,
         n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200,
         n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208,
         n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,
         n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224,
         n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232,
         n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240,
         n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248,
         n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256,
         n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264,
         n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272,
         n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280,
         n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288,
         n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296,
         n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304,
         n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312,
         n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320,
         n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328,
         n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336,
         n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344,
         n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352,
         n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360,
         n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368,
         n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376,
         n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384,
         n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392,
         n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400,
         n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408,
         n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416,
         n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424,
         n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432,
         n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440,
         n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448,
         n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456,
         n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464,
         n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472,
         n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480,
         n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488,
         n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496,
         n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504,
         n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512,
         n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520,
         n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528,
         n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536,
         n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544,
         n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552,
         n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560,
         n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568,
         n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576,
         n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584,
         n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592,
         n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600,
         n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608,
         n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616,
         n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624,
         n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632,
         n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640,
         n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648,
         n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656,
         n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664,
         n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672,
         n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680,
         n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688,
         n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696,
         n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704,
         n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712,
         n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720,
         n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728,
         n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736,
         n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744,
         n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752,
         n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760,
         n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768,
         n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776,
         n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784,
         n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,
         n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800,
         n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808,
         n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816,
         n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824,
         n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832,
         n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840,
         n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848,
         n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856,
         n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864,
         n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872,
         n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880,
         n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888,
         n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896,
         n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904,
         n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912,
         n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920,
         n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928,
         n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936,
         n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944,
         n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952,
         n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960,
         n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968,
         n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976,
         n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984,
         n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992,
         n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000,
         n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008,
         n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016,
         n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024,
         n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032,
         n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040,
         n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048,
         n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056,
         n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064,
         n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072,
         n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080,
         n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088,
         n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096,
         n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104,
         n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112,
         n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120,
         n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128,
         n27129, n27130, n27131;
  assign N18 = addr[0];
  assign N19 = addr[1];
  assign N20 = addr[2];
  assign N21 = addr[3];
  assign N22 = addr[4];
  assign N23 = addr[5];
  assign N24 = addr[6];
  assign N25 = addr[7];
  assign N26 = addr[8];
  assign N27 = addr[9];

  DFF_X1 \data_out_reg[7]  ( .D(N28), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N29), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N30), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N31), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N32), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N33), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N34), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N35), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[1023][7]  ( .D(n8609), .CK(clk), .Q(\mem[1023][7] ) );
  DFF_X1 \mem_reg[1023][6]  ( .D(n8610), .CK(clk), .Q(\mem[1023][6] ) );
  DFF_X1 \mem_reg[1023][5]  ( .D(n8611), .CK(clk), .Q(\mem[1023][5] ) );
  DFF_X1 \mem_reg[1023][4]  ( .D(n8612), .CK(clk), .Q(\mem[1023][4] ) );
  DFF_X1 \mem_reg[1023][3]  ( .D(n8613), .CK(clk), .Q(\mem[1023][3] ) );
  DFF_X1 \mem_reg[1023][2]  ( .D(n8614), .CK(clk), .Q(\mem[1023][2] ) );
  DFF_X1 \mem_reg[1023][1]  ( .D(n8615), .CK(clk), .Q(\mem[1023][1] ) );
  DFF_X1 \mem_reg[1023][0]  ( .D(n8616), .CK(clk), .Q(\mem[1023][0] ) );
  DFF_X1 \mem_reg[1022][7]  ( .D(n8617), .CK(clk), .Q(\mem[1022][7] ) );
  DFF_X1 \mem_reg[1022][6]  ( .D(n8618), .CK(clk), .Q(\mem[1022][6] ) );
  DFF_X1 \mem_reg[1022][5]  ( .D(n8619), .CK(clk), .Q(\mem[1022][5] ) );
  DFF_X1 \mem_reg[1022][4]  ( .D(n8620), .CK(clk), .Q(\mem[1022][4] ) );
  DFF_X1 \mem_reg[1022][3]  ( .D(n8621), .CK(clk), .Q(\mem[1022][3] ) );
  DFF_X1 \mem_reg[1022][2]  ( .D(n8622), .CK(clk), .Q(\mem[1022][2] ) );
  DFF_X1 \mem_reg[1022][1]  ( .D(n8623), .CK(clk), .Q(\mem[1022][1] ) );
  DFF_X1 \mem_reg[1022][0]  ( .D(n8624), .CK(clk), .Q(\mem[1022][0] ) );
  DFF_X1 \mem_reg[1021][7]  ( .D(n8625), .CK(clk), .Q(\mem[1021][7] ) );
  DFF_X1 \mem_reg[1021][6]  ( .D(n8626), .CK(clk), .Q(\mem[1021][6] ) );
  DFF_X1 \mem_reg[1021][5]  ( .D(n8627), .CK(clk), .Q(\mem[1021][5] ) );
  DFF_X1 \mem_reg[1021][4]  ( .D(n8628), .CK(clk), .Q(\mem[1021][4] ) );
  DFF_X1 \mem_reg[1021][3]  ( .D(n8629), .CK(clk), .Q(\mem[1021][3] ) );
  DFF_X1 \mem_reg[1021][2]  ( .D(n8630), .CK(clk), .Q(\mem[1021][2] ) );
  DFF_X1 \mem_reg[1021][1]  ( .D(n8631), .CK(clk), .Q(\mem[1021][1] ) );
  DFF_X1 \mem_reg[1021][0]  ( .D(n8632), .CK(clk), .Q(\mem[1021][0] ) );
  DFF_X1 \mem_reg[1020][7]  ( .D(n8633), .CK(clk), .Q(\mem[1020][7] ) );
  DFF_X1 \mem_reg[1020][6]  ( .D(n8634), .CK(clk), .Q(\mem[1020][6] ) );
  DFF_X1 \mem_reg[1020][5]  ( .D(n8635), .CK(clk), .Q(\mem[1020][5] ) );
  DFF_X1 \mem_reg[1020][4]  ( .D(n8636), .CK(clk), .Q(\mem[1020][4] ) );
  DFF_X1 \mem_reg[1020][3]  ( .D(n8637), .CK(clk), .Q(\mem[1020][3] ) );
  DFF_X1 \mem_reg[1020][2]  ( .D(n8638), .CK(clk), .Q(\mem[1020][2] ) );
  DFF_X1 \mem_reg[1020][1]  ( .D(n8639), .CK(clk), .Q(\mem[1020][1] ) );
  DFF_X1 \mem_reg[1020][0]  ( .D(n8640), .CK(clk), .Q(\mem[1020][0] ) );
  DFF_X1 \mem_reg[1019][7]  ( .D(n8641), .CK(clk), .Q(\mem[1019][7] ) );
  DFF_X1 \mem_reg[1019][6]  ( .D(n8642), .CK(clk), .Q(\mem[1019][6] ) );
  DFF_X1 \mem_reg[1019][5]  ( .D(n8643), .CK(clk), .Q(\mem[1019][5] ) );
  DFF_X1 \mem_reg[1019][4]  ( .D(n8644), .CK(clk), .Q(\mem[1019][4] ) );
  DFF_X1 \mem_reg[1019][3]  ( .D(n8645), .CK(clk), .Q(\mem[1019][3] ) );
  DFF_X1 \mem_reg[1019][2]  ( .D(n8646), .CK(clk), .Q(\mem[1019][2] ) );
  DFF_X1 \mem_reg[1019][1]  ( .D(n8647), .CK(clk), .Q(\mem[1019][1] ) );
  DFF_X1 \mem_reg[1019][0]  ( .D(n8648), .CK(clk), .Q(\mem[1019][0] ) );
  DFF_X1 \mem_reg[1018][7]  ( .D(n8649), .CK(clk), .Q(\mem[1018][7] ) );
  DFF_X1 \mem_reg[1018][6]  ( .D(n8650), .CK(clk), .Q(\mem[1018][6] ) );
  DFF_X1 \mem_reg[1018][5]  ( .D(n8651), .CK(clk), .Q(\mem[1018][5] ) );
  DFF_X1 \mem_reg[1018][4]  ( .D(n8652), .CK(clk), .Q(\mem[1018][4] ) );
  DFF_X1 \mem_reg[1018][3]  ( .D(n8653), .CK(clk), .Q(\mem[1018][3] ) );
  DFF_X1 \mem_reg[1018][2]  ( .D(n8654), .CK(clk), .Q(\mem[1018][2] ) );
  DFF_X1 \mem_reg[1018][1]  ( .D(n8655), .CK(clk), .Q(\mem[1018][1] ) );
  DFF_X1 \mem_reg[1018][0]  ( .D(n8656), .CK(clk), .Q(\mem[1018][0] ) );
  DFF_X1 \mem_reg[1017][7]  ( .D(n8657), .CK(clk), .Q(\mem[1017][7] ) );
  DFF_X1 \mem_reg[1017][6]  ( .D(n8658), .CK(clk), .Q(\mem[1017][6] ) );
  DFF_X1 \mem_reg[1017][5]  ( .D(n8659), .CK(clk), .Q(\mem[1017][5] ) );
  DFF_X1 \mem_reg[1017][4]  ( .D(n8660), .CK(clk), .Q(\mem[1017][4] ) );
  DFF_X1 \mem_reg[1017][3]  ( .D(n8661), .CK(clk), .Q(\mem[1017][3] ) );
  DFF_X1 \mem_reg[1017][2]  ( .D(n8662), .CK(clk), .Q(\mem[1017][2] ) );
  DFF_X1 \mem_reg[1017][1]  ( .D(n8663), .CK(clk), .Q(\mem[1017][1] ) );
  DFF_X1 \mem_reg[1017][0]  ( .D(n8664), .CK(clk), .Q(\mem[1017][0] ) );
  DFF_X1 \mem_reg[1016][7]  ( .D(n8665), .CK(clk), .Q(\mem[1016][7] ) );
  DFF_X1 \mem_reg[1016][6]  ( .D(n8666), .CK(clk), .Q(\mem[1016][6] ) );
  DFF_X1 \mem_reg[1016][5]  ( .D(n8667), .CK(clk), .Q(\mem[1016][5] ) );
  DFF_X1 \mem_reg[1016][4]  ( .D(n8668), .CK(clk), .Q(\mem[1016][4] ) );
  DFF_X1 \mem_reg[1016][3]  ( .D(n8669), .CK(clk), .Q(\mem[1016][3] ) );
  DFF_X1 \mem_reg[1016][2]  ( .D(n8670), .CK(clk), .Q(\mem[1016][2] ) );
  DFF_X1 \mem_reg[1016][1]  ( .D(n8671), .CK(clk), .Q(\mem[1016][1] ) );
  DFF_X1 \mem_reg[1016][0]  ( .D(n8672), .CK(clk), .Q(\mem[1016][0] ) );
  DFF_X1 \mem_reg[1015][7]  ( .D(n8673), .CK(clk), .Q(\mem[1015][7] ) );
  DFF_X1 \mem_reg[1015][6]  ( .D(n8674), .CK(clk), .Q(\mem[1015][6] ) );
  DFF_X1 \mem_reg[1015][5]  ( .D(n8675), .CK(clk), .Q(\mem[1015][5] ) );
  DFF_X1 \mem_reg[1015][4]  ( .D(n8676), .CK(clk), .Q(\mem[1015][4] ) );
  DFF_X1 \mem_reg[1015][3]  ( .D(n8677), .CK(clk), .Q(\mem[1015][3] ) );
  DFF_X1 \mem_reg[1015][2]  ( .D(n8678), .CK(clk), .Q(\mem[1015][2] ) );
  DFF_X1 \mem_reg[1015][1]  ( .D(n8679), .CK(clk), .Q(\mem[1015][1] ) );
  DFF_X1 \mem_reg[1015][0]  ( .D(n8680), .CK(clk), .Q(\mem[1015][0] ) );
  DFF_X1 \mem_reg[1014][7]  ( .D(n8681), .CK(clk), .Q(\mem[1014][7] ) );
  DFF_X1 \mem_reg[1014][6]  ( .D(n8682), .CK(clk), .Q(\mem[1014][6] ) );
  DFF_X1 \mem_reg[1014][5]  ( .D(n8683), .CK(clk), .Q(\mem[1014][5] ) );
  DFF_X1 \mem_reg[1014][4]  ( .D(n8684), .CK(clk), .Q(\mem[1014][4] ) );
  DFF_X1 \mem_reg[1014][3]  ( .D(n8685), .CK(clk), .Q(\mem[1014][3] ) );
  DFF_X1 \mem_reg[1014][2]  ( .D(n8686), .CK(clk), .Q(\mem[1014][2] ) );
  DFF_X1 \mem_reg[1014][1]  ( .D(n8687), .CK(clk), .Q(\mem[1014][1] ) );
  DFF_X1 \mem_reg[1014][0]  ( .D(n8688), .CK(clk), .Q(\mem[1014][0] ) );
  DFF_X1 \mem_reg[1013][7]  ( .D(n8689), .CK(clk), .Q(\mem[1013][7] ) );
  DFF_X1 \mem_reg[1013][6]  ( .D(n8690), .CK(clk), .Q(\mem[1013][6] ) );
  DFF_X1 \mem_reg[1013][5]  ( .D(n8691), .CK(clk), .Q(\mem[1013][5] ) );
  DFF_X1 \mem_reg[1013][4]  ( .D(n8692), .CK(clk), .Q(\mem[1013][4] ) );
  DFF_X1 \mem_reg[1013][3]  ( .D(n8693), .CK(clk), .Q(\mem[1013][3] ) );
  DFF_X1 \mem_reg[1013][2]  ( .D(n8694), .CK(clk), .Q(\mem[1013][2] ) );
  DFF_X1 \mem_reg[1013][1]  ( .D(n8695), .CK(clk), .Q(\mem[1013][1] ) );
  DFF_X1 \mem_reg[1013][0]  ( .D(n8696), .CK(clk), .Q(\mem[1013][0] ) );
  DFF_X1 \mem_reg[1012][7]  ( .D(n8697), .CK(clk), .Q(\mem[1012][7] ) );
  DFF_X1 \mem_reg[1012][6]  ( .D(n8698), .CK(clk), .Q(\mem[1012][6] ) );
  DFF_X1 \mem_reg[1012][5]  ( .D(n8699), .CK(clk), .Q(\mem[1012][5] ) );
  DFF_X1 \mem_reg[1012][4]  ( .D(n8700), .CK(clk), .Q(\mem[1012][4] ) );
  DFF_X1 \mem_reg[1012][3]  ( .D(n8701), .CK(clk), .Q(\mem[1012][3] ) );
  DFF_X1 \mem_reg[1012][2]  ( .D(n8702), .CK(clk), .Q(\mem[1012][2] ) );
  DFF_X1 \mem_reg[1012][1]  ( .D(n8703), .CK(clk), .Q(\mem[1012][1] ) );
  DFF_X1 \mem_reg[1012][0]  ( .D(n8704), .CK(clk), .Q(\mem[1012][0] ) );
  DFF_X1 \mem_reg[1011][7]  ( .D(n8705), .CK(clk), .Q(\mem[1011][7] ) );
  DFF_X1 \mem_reg[1011][6]  ( .D(n8706), .CK(clk), .Q(\mem[1011][6] ) );
  DFF_X1 \mem_reg[1011][5]  ( .D(n8707), .CK(clk), .Q(\mem[1011][5] ) );
  DFF_X1 \mem_reg[1011][4]  ( .D(n8708), .CK(clk), .Q(\mem[1011][4] ) );
  DFF_X1 \mem_reg[1011][3]  ( .D(n8709), .CK(clk), .Q(\mem[1011][3] ) );
  DFF_X1 \mem_reg[1011][2]  ( .D(n8710), .CK(clk), .Q(\mem[1011][2] ) );
  DFF_X1 \mem_reg[1011][1]  ( .D(n8711), .CK(clk), .Q(\mem[1011][1] ) );
  DFF_X1 \mem_reg[1011][0]  ( .D(n8712), .CK(clk), .Q(\mem[1011][0] ) );
  DFF_X1 \mem_reg[1010][7]  ( .D(n8713), .CK(clk), .Q(\mem[1010][7] ) );
  DFF_X1 \mem_reg[1010][6]  ( .D(n8714), .CK(clk), .Q(\mem[1010][6] ) );
  DFF_X1 \mem_reg[1010][5]  ( .D(n8715), .CK(clk), .Q(\mem[1010][5] ) );
  DFF_X1 \mem_reg[1010][4]  ( .D(n8716), .CK(clk), .Q(\mem[1010][4] ) );
  DFF_X1 \mem_reg[1010][3]  ( .D(n8717), .CK(clk), .Q(\mem[1010][3] ) );
  DFF_X1 \mem_reg[1010][2]  ( .D(n8718), .CK(clk), .Q(\mem[1010][2] ) );
  DFF_X1 \mem_reg[1010][1]  ( .D(n8719), .CK(clk), .Q(\mem[1010][1] ) );
  DFF_X1 \mem_reg[1010][0]  ( .D(n8720), .CK(clk), .Q(\mem[1010][0] ) );
  DFF_X1 \mem_reg[1009][7]  ( .D(n8721), .CK(clk), .Q(\mem[1009][7] ) );
  DFF_X1 \mem_reg[1009][6]  ( .D(n8722), .CK(clk), .Q(\mem[1009][6] ) );
  DFF_X1 \mem_reg[1009][5]  ( .D(n8723), .CK(clk), .Q(\mem[1009][5] ) );
  DFF_X1 \mem_reg[1009][4]  ( .D(n8724), .CK(clk), .Q(\mem[1009][4] ) );
  DFF_X1 \mem_reg[1009][3]  ( .D(n8725), .CK(clk), .Q(\mem[1009][3] ) );
  DFF_X1 \mem_reg[1009][2]  ( .D(n8726), .CK(clk), .Q(\mem[1009][2] ) );
  DFF_X1 \mem_reg[1009][1]  ( .D(n8727), .CK(clk), .Q(\mem[1009][1] ) );
  DFF_X1 \mem_reg[1009][0]  ( .D(n8728), .CK(clk), .Q(\mem[1009][0] ) );
  DFF_X1 \mem_reg[1008][7]  ( .D(n8729), .CK(clk), .Q(\mem[1008][7] ) );
  DFF_X1 \mem_reg[1008][6]  ( .D(n8730), .CK(clk), .Q(\mem[1008][6] ) );
  DFF_X1 \mem_reg[1008][5]  ( .D(n8731), .CK(clk), .Q(\mem[1008][5] ) );
  DFF_X1 \mem_reg[1008][4]  ( .D(n8732), .CK(clk), .Q(\mem[1008][4] ) );
  DFF_X1 \mem_reg[1008][3]  ( .D(n8733), .CK(clk), .Q(\mem[1008][3] ) );
  DFF_X1 \mem_reg[1008][2]  ( .D(n8734), .CK(clk), .Q(\mem[1008][2] ) );
  DFF_X1 \mem_reg[1008][1]  ( .D(n8735), .CK(clk), .Q(\mem[1008][1] ) );
  DFF_X1 \mem_reg[1008][0]  ( .D(n8736), .CK(clk), .Q(\mem[1008][0] ) );
  DFF_X1 \mem_reg[1007][7]  ( .D(n8737), .CK(clk), .Q(\mem[1007][7] ) );
  DFF_X1 \mem_reg[1007][6]  ( .D(n8738), .CK(clk), .Q(\mem[1007][6] ) );
  DFF_X1 \mem_reg[1007][5]  ( .D(n8739), .CK(clk), .Q(\mem[1007][5] ) );
  DFF_X1 \mem_reg[1007][4]  ( .D(n8740), .CK(clk), .Q(\mem[1007][4] ) );
  DFF_X1 \mem_reg[1007][3]  ( .D(n8741), .CK(clk), .Q(\mem[1007][3] ) );
  DFF_X1 \mem_reg[1007][2]  ( .D(n8742), .CK(clk), .Q(\mem[1007][2] ) );
  DFF_X1 \mem_reg[1007][1]  ( .D(n8743), .CK(clk), .Q(\mem[1007][1] ) );
  DFF_X1 \mem_reg[1007][0]  ( .D(n8744), .CK(clk), .Q(\mem[1007][0] ) );
  DFF_X1 \mem_reg[1006][7]  ( .D(n8745), .CK(clk), .Q(\mem[1006][7] ) );
  DFF_X1 \mem_reg[1006][6]  ( .D(n8746), .CK(clk), .Q(\mem[1006][6] ) );
  DFF_X1 \mem_reg[1006][5]  ( .D(n8747), .CK(clk), .Q(\mem[1006][5] ) );
  DFF_X1 \mem_reg[1006][4]  ( .D(n8748), .CK(clk), .Q(\mem[1006][4] ) );
  DFF_X1 \mem_reg[1006][3]  ( .D(n8749), .CK(clk), .Q(\mem[1006][3] ) );
  DFF_X1 \mem_reg[1006][2]  ( .D(n8750), .CK(clk), .Q(\mem[1006][2] ) );
  DFF_X1 \mem_reg[1006][1]  ( .D(n8751), .CK(clk), .Q(\mem[1006][1] ) );
  DFF_X1 \mem_reg[1006][0]  ( .D(n8752), .CK(clk), .Q(\mem[1006][0] ) );
  DFF_X1 \mem_reg[1005][7]  ( .D(n8753), .CK(clk), .Q(\mem[1005][7] ) );
  DFF_X1 \mem_reg[1005][6]  ( .D(n8754), .CK(clk), .Q(\mem[1005][6] ) );
  DFF_X1 \mem_reg[1005][5]  ( .D(n8755), .CK(clk), .Q(\mem[1005][5] ) );
  DFF_X1 \mem_reg[1005][4]  ( .D(n8756), .CK(clk), .Q(\mem[1005][4] ) );
  DFF_X1 \mem_reg[1005][3]  ( .D(n8757), .CK(clk), .Q(\mem[1005][3] ) );
  DFF_X1 \mem_reg[1005][2]  ( .D(n8758), .CK(clk), .Q(\mem[1005][2] ) );
  DFF_X1 \mem_reg[1005][1]  ( .D(n8759), .CK(clk), .Q(\mem[1005][1] ) );
  DFF_X1 \mem_reg[1005][0]  ( .D(n8760), .CK(clk), .Q(\mem[1005][0] ) );
  DFF_X1 \mem_reg[1004][7]  ( .D(n8761), .CK(clk), .Q(\mem[1004][7] ) );
  DFF_X1 \mem_reg[1004][6]  ( .D(n8762), .CK(clk), .Q(\mem[1004][6] ) );
  DFF_X1 \mem_reg[1004][5]  ( .D(n8763), .CK(clk), .Q(\mem[1004][5] ) );
  DFF_X1 \mem_reg[1004][4]  ( .D(n8764), .CK(clk), .Q(\mem[1004][4] ) );
  DFF_X1 \mem_reg[1004][3]  ( .D(n8765), .CK(clk), .Q(\mem[1004][3] ) );
  DFF_X1 \mem_reg[1004][2]  ( .D(n8766), .CK(clk), .Q(\mem[1004][2] ) );
  DFF_X1 \mem_reg[1004][1]  ( .D(n8767), .CK(clk), .Q(\mem[1004][1] ) );
  DFF_X1 \mem_reg[1004][0]  ( .D(n8768), .CK(clk), .Q(\mem[1004][0] ) );
  DFF_X1 \mem_reg[1003][7]  ( .D(n8769), .CK(clk), .Q(\mem[1003][7] ) );
  DFF_X1 \mem_reg[1003][6]  ( .D(n8770), .CK(clk), .Q(\mem[1003][6] ) );
  DFF_X1 \mem_reg[1003][5]  ( .D(n8771), .CK(clk), .Q(\mem[1003][5] ) );
  DFF_X1 \mem_reg[1003][4]  ( .D(n8772), .CK(clk), .Q(\mem[1003][4] ) );
  DFF_X1 \mem_reg[1003][3]  ( .D(n8773), .CK(clk), .Q(\mem[1003][3] ) );
  DFF_X1 \mem_reg[1003][2]  ( .D(n8774), .CK(clk), .Q(\mem[1003][2] ) );
  DFF_X1 \mem_reg[1003][1]  ( .D(n8775), .CK(clk), .Q(\mem[1003][1] ) );
  DFF_X1 \mem_reg[1003][0]  ( .D(n8776), .CK(clk), .Q(\mem[1003][0] ) );
  DFF_X1 \mem_reg[1002][7]  ( .D(n8777), .CK(clk), .Q(\mem[1002][7] ) );
  DFF_X1 \mem_reg[1002][6]  ( .D(n8778), .CK(clk), .Q(\mem[1002][6] ) );
  DFF_X1 \mem_reg[1002][5]  ( .D(n8779), .CK(clk), .Q(\mem[1002][5] ) );
  DFF_X1 \mem_reg[1002][4]  ( .D(n8780), .CK(clk), .Q(\mem[1002][4] ) );
  DFF_X1 \mem_reg[1002][3]  ( .D(n8781), .CK(clk), .Q(\mem[1002][3] ) );
  DFF_X1 \mem_reg[1002][2]  ( .D(n8782), .CK(clk), .Q(\mem[1002][2] ) );
  DFF_X1 \mem_reg[1002][1]  ( .D(n8783), .CK(clk), .Q(\mem[1002][1] ) );
  DFF_X1 \mem_reg[1002][0]  ( .D(n8784), .CK(clk), .Q(\mem[1002][0] ) );
  DFF_X1 \mem_reg[1001][7]  ( .D(n8785), .CK(clk), .Q(\mem[1001][7] ) );
  DFF_X1 \mem_reg[1001][6]  ( .D(n8786), .CK(clk), .Q(\mem[1001][6] ) );
  DFF_X1 \mem_reg[1001][5]  ( .D(n8787), .CK(clk), .Q(\mem[1001][5] ) );
  DFF_X1 \mem_reg[1001][4]  ( .D(n8788), .CK(clk), .Q(\mem[1001][4] ) );
  DFF_X1 \mem_reg[1001][3]  ( .D(n8789), .CK(clk), .Q(\mem[1001][3] ) );
  DFF_X1 \mem_reg[1001][2]  ( .D(n8790), .CK(clk), .Q(\mem[1001][2] ) );
  DFF_X1 \mem_reg[1001][1]  ( .D(n8791), .CK(clk), .Q(\mem[1001][1] ) );
  DFF_X1 \mem_reg[1001][0]  ( .D(n8792), .CK(clk), .Q(\mem[1001][0] ) );
  DFF_X1 \mem_reg[1000][7]  ( .D(n8793), .CK(clk), .Q(\mem[1000][7] ) );
  DFF_X1 \mem_reg[1000][6]  ( .D(n8794), .CK(clk), .Q(\mem[1000][6] ) );
  DFF_X1 \mem_reg[1000][5]  ( .D(n8795), .CK(clk), .Q(\mem[1000][5] ) );
  DFF_X1 \mem_reg[1000][4]  ( .D(n8796), .CK(clk), .Q(\mem[1000][4] ) );
  DFF_X1 \mem_reg[1000][3]  ( .D(n8797), .CK(clk), .Q(\mem[1000][3] ) );
  DFF_X1 \mem_reg[1000][2]  ( .D(n8798), .CK(clk), .Q(\mem[1000][2] ) );
  DFF_X1 \mem_reg[1000][1]  ( .D(n8799), .CK(clk), .Q(\mem[1000][1] ) );
  DFF_X1 \mem_reg[1000][0]  ( .D(n8800), .CK(clk), .Q(\mem[1000][0] ) );
  DFF_X1 \mem_reg[999][7]  ( .D(n8801), .CK(clk), .Q(\mem[999][7] ) );
  DFF_X1 \mem_reg[999][6]  ( .D(n8802), .CK(clk), .Q(\mem[999][6] ) );
  DFF_X1 \mem_reg[999][5]  ( .D(n8803), .CK(clk), .Q(\mem[999][5] ) );
  DFF_X1 \mem_reg[999][4]  ( .D(n8804), .CK(clk), .Q(\mem[999][4] ) );
  DFF_X1 \mem_reg[999][3]  ( .D(n8805), .CK(clk), .Q(\mem[999][3] ) );
  DFF_X1 \mem_reg[999][2]  ( .D(n8806), .CK(clk), .Q(\mem[999][2] ) );
  DFF_X1 \mem_reg[999][1]  ( .D(n8807), .CK(clk), .Q(\mem[999][1] ) );
  DFF_X1 \mem_reg[999][0]  ( .D(n8808), .CK(clk), .Q(\mem[999][0] ) );
  DFF_X1 \mem_reg[998][7]  ( .D(n8809), .CK(clk), .Q(\mem[998][7] ) );
  DFF_X1 \mem_reg[998][6]  ( .D(n8810), .CK(clk), .Q(\mem[998][6] ) );
  DFF_X1 \mem_reg[998][5]  ( .D(n8811), .CK(clk), .Q(\mem[998][5] ) );
  DFF_X1 \mem_reg[998][4]  ( .D(n8812), .CK(clk), .Q(\mem[998][4] ) );
  DFF_X1 \mem_reg[998][3]  ( .D(n8813), .CK(clk), .Q(\mem[998][3] ) );
  DFF_X1 \mem_reg[998][2]  ( .D(n8814), .CK(clk), .Q(\mem[998][2] ) );
  DFF_X1 \mem_reg[998][1]  ( .D(n8815), .CK(clk), .Q(\mem[998][1] ) );
  DFF_X1 \mem_reg[998][0]  ( .D(n8816), .CK(clk), .Q(\mem[998][0] ) );
  DFF_X1 \mem_reg[997][7]  ( .D(n8817), .CK(clk), .Q(\mem[997][7] ) );
  DFF_X1 \mem_reg[997][6]  ( .D(n8818), .CK(clk), .Q(\mem[997][6] ) );
  DFF_X1 \mem_reg[997][5]  ( .D(n8819), .CK(clk), .Q(\mem[997][5] ) );
  DFF_X1 \mem_reg[997][4]  ( .D(n8820), .CK(clk), .Q(\mem[997][4] ) );
  DFF_X1 \mem_reg[997][3]  ( .D(n8821), .CK(clk), .Q(\mem[997][3] ) );
  DFF_X1 \mem_reg[997][2]  ( .D(n8822), .CK(clk), .Q(\mem[997][2] ) );
  DFF_X1 \mem_reg[997][1]  ( .D(n8823), .CK(clk), .Q(\mem[997][1] ) );
  DFF_X1 \mem_reg[997][0]  ( .D(n8824), .CK(clk), .Q(\mem[997][0] ) );
  DFF_X1 \mem_reg[996][7]  ( .D(n8825), .CK(clk), .Q(\mem[996][7] ) );
  DFF_X1 \mem_reg[996][6]  ( .D(n8826), .CK(clk), .Q(\mem[996][6] ) );
  DFF_X1 \mem_reg[996][5]  ( .D(n8827), .CK(clk), .Q(\mem[996][5] ) );
  DFF_X1 \mem_reg[996][4]  ( .D(n8828), .CK(clk), .Q(\mem[996][4] ) );
  DFF_X1 \mem_reg[996][3]  ( .D(n8829), .CK(clk), .Q(\mem[996][3] ) );
  DFF_X1 \mem_reg[996][2]  ( .D(n8830), .CK(clk), .Q(\mem[996][2] ) );
  DFF_X1 \mem_reg[996][1]  ( .D(n8831), .CK(clk), .Q(\mem[996][1] ) );
  DFF_X1 \mem_reg[996][0]  ( .D(n8832), .CK(clk), .Q(\mem[996][0] ) );
  DFF_X1 \mem_reg[995][7]  ( .D(n8833), .CK(clk), .Q(\mem[995][7] ) );
  DFF_X1 \mem_reg[995][6]  ( .D(n8834), .CK(clk), .Q(\mem[995][6] ) );
  DFF_X1 \mem_reg[995][5]  ( .D(n8835), .CK(clk), .Q(\mem[995][5] ) );
  DFF_X1 \mem_reg[995][4]  ( .D(n8836), .CK(clk), .Q(\mem[995][4] ) );
  DFF_X1 \mem_reg[995][3]  ( .D(n8837), .CK(clk), .Q(\mem[995][3] ) );
  DFF_X1 \mem_reg[995][2]  ( .D(n8838), .CK(clk), .Q(\mem[995][2] ) );
  DFF_X1 \mem_reg[995][1]  ( .D(n8839), .CK(clk), .Q(\mem[995][1] ) );
  DFF_X1 \mem_reg[995][0]  ( .D(n8840), .CK(clk), .Q(\mem[995][0] ) );
  DFF_X1 \mem_reg[994][7]  ( .D(n8841), .CK(clk), .Q(\mem[994][7] ) );
  DFF_X1 \mem_reg[994][6]  ( .D(n8842), .CK(clk), .Q(\mem[994][6] ) );
  DFF_X1 \mem_reg[994][5]  ( .D(n8843), .CK(clk), .Q(\mem[994][5] ) );
  DFF_X1 \mem_reg[994][4]  ( .D(n8844), .CK(clk), .Q(\mem[994][4] ) );
  DFF_X1 \mem_reg[994][3]  ( .D(n8845), .CK(clk), .Q(\mem[994][3] ) );
  DFF_X1 \mem_reg[994][2]  ( .D(n8846), .CK(clk), .Q(\mem[994][2] ) );
  DFF_X1 \mem_reg[994][1]  ( .D(n8847), .CK(clk), .Q(\mem[994][1] ) );
  DFF_X1 \mem_reg[994][0]  ( .D(n8848), .CK(clk), .Q(\mem[994][0] ) );
  DFF_X1 \mem_reg[993][7]  ( .D(n8849), .CK(clk), .Q(\mem[993][7] ) );
  DFF_X1 \mem_reg[993][6]  ( .D(n8850), .CK(clk), .Q(\mem[993][6] ) );
  DFF_X1 \mem_reg[993][5]  ( .D(n8851), .CK(clk), .Q(\mem[993][5] ) );
  DFF_X1 \mem_reg[993][4]  ( .D(n8852), .CK(clk), .Q(\mem[993][4] ) );
  DFF_X1 \mem_reg[993][3]  ( .D(n8853), .CK(clk), .Q(\mem[993][3] ) );
  DFF_X1 \mem_reg[993][2]  ( .D(n8854), .CK(clk), .Q(\mem[993][2] ) );
  DFF_X1 \mem_reg[993][1]  ( .D(n8855), .CK(clk), .Q(\mem[993][1] ) );
  DFF_X1 \mem_reg[993][0]  ( .D(n8856), .CK(clk), .Q(\mem[993][0] ) );
  DFF_X1 \mem_reg[992][7]  ( .D(n8857), .CK(clk), .Q(\mem[992][7] ) );
  DFF_X1 \mem_reg[992][6]  ( .D(n8858), .CK(clk), .Q(\mem[992][6] ) );
  DFF_X1 \mem_reg[992][5]  ( .D(n8859), .CK(clk), .Q(\mem[992][5] ) );
  DFF_X1 \mem_reg[992][4]  ( .D(n8860), .CK(clk), .Q(\mem[992][4] ) );
  DFF_X1 \mem_reg[992][3]  ( .D(n8861), .CK(clk), .Q(\mem[992][3] ) );
  DFF_X1 \mem_reg[992][2]  ( .D(n8862), .CK(clk), .Q(\mem[992][2] ) );
  DFF_X1 \mem_reg[992][1]  ( .D(n8863), .CK(clk), .Q(\mem[992][1] ) );
  DFF_X1 \mem_reg[992][0]  ( .D(n8864), .CK(clk), .Q(\mem[992][0] ) );
  DFF_X1 \mem_reg[991][7]  ( .D(n8865), .CK(clk), .Q(\mem[991][7] ) );
  DFF_X1 \mem_reg[991][6]  ( .D(n8866), .CK(clk), .Q(\mem[991][6] ) );
  DFF_X1 \mem_reg[991][5]  ( .D(n8867), .CK(clk), .Q(\mem[991][5] ) );
  DFF_X1 \mem_reg[991][4]  ( .D(n8868), .CK(clk), .Q(\mem[991][4] ) );
  DFF_X1 \mem_reg[991][3]  ( .D(n8869), .CK(clk), .Q(\mem[991][3] ) );
  DFF_X1 \mem_reg[991][2]  ( .D(n8870), .CK(clk), .Q(\mem[991][2] ) );
  DFF_X1 \mem_reg[991][1]  ( .D(n8871), .CK(clk), .Q(\mem[991][1] ) );
  DFF_X1 \mem_reg[991][0]  ( .D(n8872), .CK(clk), .Q(\mem[991][0] ) );
  DFF_X1 \mem_reg[990][7]  ( .D(n8873), .CK(clk), .Q(\mem[990][7] ) );
  DFF_X1 \mem_reg[990][6]  ( .D(n8874), .CK(clk), .Q(\mem[990][6] ) );
  DFF_X1 \mem_reg[990][5]  ( .D(n8875), .CK(clk), .Q(\mem[990][5] ) );
  DFF_X1 \mem_reg[990][4]  ( .D(n8876), .CK(clk), .Q(\mem[990][4] ) );
  DFF_X1 \mem_reg[990][3]  ( .D(n8877), .CK(clk), .Q(\mem[990][3] ) );
  DFF_X1 \mem_reg[990][2]  ( .D(n8878), .CK(clk), .Q(\mem[990][2] ) );
  DFF_X1 \mem_reg[990][1]  ( .D(n8879), .CK(clk), .Q(\mem[990][1] ) );
  DFF_X1 \mem_reg[990][0]  ( .D(n8880), .CK(clk), .Q(\mem[990][0] ) );
  DFF_X1 \mem_reg[989][7]  ( .D(n8881), .CK(clk), .Q(\mem[989][7] ) );
  DFF_X1 \mem_reg[989][6]  ( .D(n8882), .CK(clk), .Q(\mem[989][6] ) );
  DFF_X1 \mem_reg[989][5]  ( .D(n8883), .CK(clk), .Q(\mem[989][5] ) );
  DFF_X1 \mem_reg[989][4]  ( .D(n8884), .CK(clk), .Q(\mem[989][4] ) );
  DFF_X1 \mem_reg[989][3]  ( .D(n8885), .CK(clk), .Q(\mem[989][3] ) );
  DFF_X1 \mem_reg[989][2]  ( .D(n8886), .CK(clk), .Q(\mem[989][2] ) );
  DFF_X1 \mem_reg[989][1]  ( .D(n8887), .CK(clk), .Q(\mem[989][1] ) );
  DFF_X1 \mem_reg[989][0]  ( .D(n8888), .CK(clk), .Q(\mem[989][0] ) );
  DFF_X1 \mem_reg[988][7]  ( .D(n8889), .CK(clk), .Q(\mem[988][7] ) );
  DFF_X1 \mem_reg[988][6]  ( .D(n8890), .CK(clk), .Q(\mem[988][6] ) );
  DFF_X1 \mem_reg[988][5]  ( .D(n8891), .CK(clk), .Q(\mem[988][5] ) );
  DFF_X1 \mem_reg[988][4]  ( .D(n8892), .CK(clk), .Q(\mem[988][4] ) );
  DFF_X1 \mem_reg[988][3]  ( .D(n8893), .CK(clk), .Q(\mem[988][3] ) );
  DFF_X1 \mem_reg[988][2]  ( .D(n8894), .CK(clk), .Q(\mem[988][2] ) );
  DFF_X1 \mem_reg[988][1]  ( .D(n8895), .CK(clk), .Q(\mem[988][1] ) );
  DFF_X1 \mem_reg[988][0]  ( .D(n8896), .CK(clk), .Q(\mem[988][0] ) );
  DFF_X1 \mem_reg[987][7]  ( .D(n8897), .CK(clk), .Q(\mem[987][7] ) );
  DFF_X1 \mem_reg[987][6]  ( .D(n8898), .CK(clk), .Q(\mem[987][6] ) );
  DFF_X1 \mem_reg[987][5]  ( .D(n8899), .CK(clk), .Q(\mem[987][5] ) );
  DFF_X1 \mem_reg[987][4]  ( .D(n8900), .CK(clk), .Q(\mem[987][4] ) );
  DFF_X1 \mem_reg[987][3]  ( .D(n8901), .CK(clk), .Q(\mem[987][3] ) );
  DFF_X1 \mem_reg[987][2]  ( .D(n8902), .CK(clk), .Q(\mem[987][2] ) );
  DFF_X1 \mem_reg[987][1]  ( .D(n8903), .CK(clk), .Q(\mem[987][1] ) );
  DFF_X1 \mem_reg[987][0]  ( .D(n8904), .CK(clk), .Q(\mem[987][0] ) );
  DFF_X1 \mem_reg[986][7]  ( .D(n8905), .CK(clk), .Q(\mem[986][7] ) );
  DFF_X1 \mem_reg[986][6]  ( .D(n8906), .CK(clk), .Q(\mem[986][6] ) );
  DFF_X1 \mem_reg[986][5]  ( .D(n8907), .CK(clk), .Q(\mem[986][5] ) );
  DFF_X1 \mem_reg[986][4]  ( .D(n8908), .CK(clk), .Q(\mem[986][4] ) );
  DFF_X1 \mem_reg[986][3]  ( .D(n8909), .CK(clk), .Q(\mem[986][3] ) );
  DFF_X1 \mem_reg[986][2]  ( .D(n8910), .CK(clk), .Q(\mem[986][2] ) );
  DFF_X1 \mem_reg[986][1]  ( .D(n8911), .CK(clk), .Q(\mem[986][1] ) );
  DFF_X1 \mem_reg[986][0]  ( .D(n8912), .CK(clk), .Q(\mem[986][0] ) );
  DFF_X1 \mem_reg[985][7]  ( .D(n8913), .CK(clk), .Q(\mem[985][7] ) );
  DFF_X1 \mem_reg[985][6]  ( .D(n8914), .CK(clk), .Q(\mem[985][6] ) );
  DFF_X1 \mem_reg[985][5]  ( .D(n8915), .CK(clk), .Q(\mem[985][5] ) );
  DFF_X1 \mem_reg[985][4]  ( .D(n8916), .CK(clk), .Q(\mem[985][4] ) );
  DFF_X1 \mem_reg[985][3]  ( .D(n8917), .CK(clk), .Q(\mem[985][3] ) );
  DFF_X1 \mem_reg[985][2]  ( .D(n8918), .CK(clk), .Q(\mem[985][2] ) );
  DFF_X1 \mem_reg[985][1]  ( .D(n8919), .CK(clk), .Q(\mem[985][1] ) );
  DFF_X1 \mem_reg[985][0]  ( .D(n8920), .CK(clk), .Q(\mem[985][0] ) );
  DFF_X1 \mem_reg[984][7]  ( .D(n8921), .CK(clk), .Q(\mem[984][7] ) );
  DFF_X1 \mem_reg[984][6]  ( .D(n8922), .CK(clk), .Q(\mem[984][6] ) );
  DFF_X1 \mem_reg[984][5]  ( .D(n8923), .CK(clk), .Q(\mem[984][5] ) );
  DFF_X1 \mem_reg[984][4]  ( .D(n8924), .CK(clk), .Q(\mem[984][4] ) );
  DFF_X1 \mem_reg[984][3]  ( .D(n8925), .CK(clk), .Q(\mem[984][3] ) );
  DFF_X1 \mem_reg[984][2]  ( .D(n8926), .CK(clk), .Q(\mem[984][2] ) );
  DFF_X1 \mem_reg[984][1]  ( .D(n8927), .CK(clk), .Q(\mem[984][1] ) );
  DFF_X1 \mem_reg[984][0]  ( .D(n8928), .CK(clk), .Q(\mem[984][0] ) );
  DFF_X1 \mem_reg[983][7]  ( .D(n8929), .CK(clk), .Q(\mem[983][7] ) );
  DFF_X1 \mem_reg[983][6]  ( .D(n8930), .CK(clk), .Q(\mem[983][6] ) );
  DFF_X1 \mem_reg[983][5]  ( .D(n8931), .CK(clk), .Q(\mem[983][5] ) );
  DFF_X1 \mem_reg[983][4]  ( .D(n8932), .CK(clk), .Q(\mem[983][4] ) );
  DFF_X1 \mem_reg[983][3]  ( .D(n8933), .CK(clk), .Q(\mem[983][3] ) );
  DFF_X1 \mem_reg[983][2]  ( .D(n8934), .CK(clk), .Q(\mem[983][2] ) );
  DFF_X1 \mem_reg[983][1]  ( .D(n8935), .CK(clk), .Q(\mem[983][1] ) );
  DFF_X1 \mem_reg[983][0]  ( .D(n8936), .CK(clk), .Q(\mem[983][0] ) );
  DFF_X1 \mem_reg[982][7]  ( .D(n8937), .CK(clk), .Q(\mem[982][7] ) );
  DFF_X1 \mem_reg[982][6]  ( .D(n8938), .CK(clk), .Q(\mem[982][6] ) );
  DFF_X1 \mem_reg[982][5]  ( .D(n8939), .CK(clk), .Q(\mem[982][5] ) );
  DFF_X1 \mem_reg[982][4]  ( .D(n8940), .CK(clk), .Q(\mem[982][4] ) );
  DFF_X1 \mem_reg[982][3]  ( .D(n8941), .CK(clk), .Q(\mem[982][3] ) );
  DFF_X1 \mem_reg[982][2]  ( .D(n8942), .CK(clk), .Q(\mem[982][2] ) );
  DFF_X1 \mem_reg[982][1]  ( .D(n8943), .CK(clk), .Q(\mem[982][1] ) );
  DFF_X1 \mem_reg[982][0]  ( .D(n8944), .CK(clk), .Q(\mem[982][0] ) );
  DFF_X1 \mem_reg[981][7]  ( .D(n8945), .CK(clk), .Q(\mem[981][7] ) );
  DFF_X1 \mem_reg[981][6]  ( .D(n8946), .CK(clk), .Q(\mem[981][6] ) );
  DFF_X1 \mem_reg[981][5]  ( .D(n8947), .CK(clk), .Q(\mem[981][5] ) );
  DFF_X1 \mem_reg[981][4]  ( .D(n8948), .CK(clk), .Q(\mem[981][4] ) );
  DFF_X1 \mem_reg[981][3]  ( .D(n8949), .CK(clk), .Q(\mem[981][3] ) );
  DFF_X1 \mem_reg[981][2]  ( .D(n8950), .CK(clk), .Q(\mem[981][2] ) );
  DFF_X1 \mem_reg[981][1]  ( .D(n8951), .CK(clk), .Q(\mem[981][1] ) );
  DFF_X1 \mem_reg[981][0]  ( .D(n8952), .CK(clk), .Q(\mem[981][0] ) );
  DFF_X1 \mem_reg[980][7]  ( .D(n8953), .CK(clk), .Q(\mem[980][7] ) );
  DFF_X1 \mem_reg[980][6]  ( .D(n8954), .CK(clk), .Q(\mem[980][6] ) );
  DFF_X1 \mem_reg[980][5]  ( .D(n8955), .CK(clk), .Q(\mem[980][5] ) );
  DFF_X1 \mem_reg[980][4]  ( .D(n8956), .CK(clk), .Q(\mem[980][4] ) );
  DFF_X1 \mem_reg[980][3]  ( .D(n8957), .CK(clk), .Q(\mem[980][3] ) );
  DFF_X1 \mem_reg[980][2]  ( .D(n8958), .CK(clk), .Q(\mem[980][2] ) );
  DFF_X1 \mem_reg[980][1]  ( .D(n8959), .CK(clk), .Q(\mem[980][1] ) );
  DFF_X1 \mem_reg[980][0]  ( .D(n8960), .CK(clk), .Q(\mem[980][0] ) );
  DFF_X1 \mem_reg[979][7]  ( .D(n8961), .CK(clk), .Q(\mem[979][7] ) );
  DFF_X1 \mem_reg[979][6]  ( .D(n8962), .CK(clk), .Q(\mem[979][6] ) );
  DFF_X1 \mem_reg[979][5]  ( .D(n8963), .CK(clk), .Q(\mem[979][5] ) );
  DFF_X1 \mem_reg[979][4]  ( .D(n8964), .CK(clk), .Q(\mem[979][4] ) );
  DFF_X1 \mem_reg[979][3]  ( .D(n8965), .CK(clk), .Q(\mem[979][3] ) );
  DFF_X1 \mem_reg[979][2]  ( .D(n8966), .CK(clk), .Q(\mem[979][2] ) );
  DFF_X1 \mem_reg[979][1]  ( .D(n8967), .CK(clk), .Q(\mem[979][1] ) );
  DFF_X1 \mem_reg[979][0]  ( .D(n8968), .CK(clk), .Q(\mem[979][0] ) );
  DFF_X1 \mem_reg[978][7]  ( .D(n8969), .CK(clk), .Q(\mem[978][7] ) );
  DFF_X1 \mem_reg[978][6]  ( .D(n8970), .CK(clk), .Q(\mem[978][6] ) );
  DFF_X1 \mem_reg[978][5]  ( .D(n8971), .CK(clk), .Q(\mem[978][5] ) );
  DFF_X1 \mem_reg[978][4]  ( .D(n8972), .CK(clk), .Q(\mem[978][4] ) );
  DFF_X1 \mem_reg[978][3]  ( .D(n8973), .CK(clk), .Q(\mem[978][3] ) );
  DFF_X1 \mem_reg[978][2]  ( .D(n8974), .CK(clk), .Q(\mem[978][2] ) );
  DFF_X1 \mem_reg[978][1]  ( .D(n8975), .CK(clk), .Q(\mem[978][1] ) );
  DFF_X1 \mem_reg[978][0]  ( .D(n8976), .CK(clk), .Q(\mem[978][0] ) );
  DFF_X1 \mem_reg[977][7]  ( .D(n8977), .CK(clk), .Q(\mem[977][7] ) );
  DFF_X1 \mem_reg[977][6]  ( .D(n8978), .CK(clk), .Q(\mem[977][6] ) );
  DFF_X1 \mem_reg[977][5]  ( .D(n8979), .CK(clk), .Q(\mem[977][5] ) );
  DFF_X1 \mem_reg[977][4]  ( .D(n8980), .CK(clk), .Q(\mem[977][4] ) );
  DFF_X1 \mem_reg[977][3]  ( .D(n8981), .CK(clk), .Q(\mem[977][3] ) );
  DFF_X1 \mem_reg[977][2]  ( .D(n8982), .CK(clk), .Q(\mem[977][2] ) );
  DFF_X1 \mem_reg[977][1]  ( .D(n8983), .CK(clk), .Q(\mem[977][1] ) );
  DFF_X1 \mem_reg[977][0]  ( .D(n8984), .CK(clk), .Q(\mem[977][0] ) );
  DFF_X1 \mem_reg[976][7]  ( .D(n8985), .CK(clk), .Q(\mem[976][7] ) );
  DFF_X1 \mem_reg[976][6]  ( .D(n8986), .CK(clk), .Q(\mem[976][6] ) );
  DFF_X1 \mem_reg[976][5]  ( .D(n8987), .CK(clk), .Q(\mem[976][5] ) );
  DFF_X1 \mem_reg[976][4]  ( .D(n8988), .CK(clk), .Q(\mem[976][4] ) );
  DFF_X1 \mem_reg[976][3]  ( .D(n8989), .CK(clk), .Q(\mem[976][3] ) );
  DFF_X1 \mem_reg[976][2]  ( .D(n8990), .CK(clk), .Q(\mem[976][2] ) );
  DFF_X1 \mem_reg[976][1]  ( .D(n8991), .CK(clk), .Q(\mem[976][1] ) );
  DFF_X1 \mem_reg[976][0]  ( .D(n8992), .CK(clk), .Q(\mem[976][0] ) );
  DFF_X1 \mem_reg[975][7]  ( .D(n8993), .CK(clk), .Q(\mem[975][7] ) );
  DFF_X1 \mem_reg[975][6]  ( .D(n8994), .CK(clk), .Q(\mem[975][6] ) );
  DFF_X1 \mem_reg[975][5]  ( .D(n8995), .CK(clk), .Q(\mem[975][5] ) );
  DFF_X1 \mem_reg[975][4]  ( .D(n8996), .CK(clk), .Q(\mem[975][4] ) );
  DFF_X1 \mem_reg[975][3]  ( .D(n8997), .CK(clk), .Q(\mem[975][3] ) );
  DFF_X1 \mem_reg[975][2]  ( .D(n8998), .CK(clk), .Q(\mem[975][2] ) );
  DFF_X1 \mem_reg[975][1]  ( .D(n8999), .CK(clk), .Q(\mem[975][1] ) );
  DFF_X1 \mem_reg[975][0]  ( .D(n9000), .CK(clk), .Q(\mem[975][0] ) );
  DFF_X1 \mem_reg[974][7]  ( .D(n9001), .CK(clk), .Q(\mem[974][7] ) );
  DFF_X1 \mem_reg[974][6]  ( .D(n9002), .CK(clk), .Q(\mem[974][6] ) );
  DFF_X1 \mem_reg[974][5]  ( .D(n9003), .CK(clk), .Q(\mem[974][5] ) );
  DFF_X1 \mem_reg[974][4]  ( .D(n9004), .CK(clk), .Q(\mem[974][4] ) );
  DFF_X1 \mem_reg[974][3]  ( .D(n9005), .CK(clk), .Q(\mem[974][3] ) );
  DFF_X1 \mem_reg[974][2]  ( .D(n9006), .CK(clk), .Q(\mem[974][2] ) );
  DFF_X1 \mem_reg[974][1]  ( .D(n9007), .CK(clk), .Q(\mem[974][1] ) );
  DFF_X1 \mem_reg[974][0]  ( .D(n9008), .CK(clk), .Q(\mem[974][0] ) );
  DFF_X1 \mem_reg[973][7]  ( .D(n9009), .CK(clk), .Q(\mem[973][7] ) );
  DFF_X1 \mem_reg[973][6]  ( .D(n9010), .CK(clk), .Q(\mem[973][6] ) );
  DFF_X1 \mem_reg[973][5]  ( .D(n9011), .CK(clk), .Q(\mem[973][5] ) );
  DFF_X1 \mem_reg[973][4]  ( .D(n9012), .CK(clk), .Q(\mem[973][4] ) );
  DFF_X1 \mem_reg[973][3]  ( .D(n9013), .CK(clk), .Q(\mem[973][3] ) );
  DFF_X1 \mem_reg[973][2]  ( .D(n9014), .CK(clk), .Q(\mem[973][2] ) );
  DFF_X1 \mem_reg[973][1]  ( .D(n9015), .CK(clk), .Q(\mem[973][1] ) );
  DFF_X1 \mem_reg[973][0]  ( .D(n9016), .CK(clk), .Q(\mem[973][0] ) );
  DFF_X1 \mem_reg[972][7]  ( .D(n9017), .CK(clk), .Q(\mem[972][7] ) );
  DFF_X1 \mem_reg[972][6]  ( .D(n9018), .CK(clk), .Q(\mem[972][6] ) );
  DFF_X1 \mem_reg[972][5]  ( .D(n9019), .CK(clk), .Q(\mem[972][5] ) );
  DFF_X1 \mem_reg[972][4]  ( .D(n9020), .CK(clk), .Q(\mem[972][4] ) );
  DFF_X1 \mem_reg[972][3]  ( .D(n9021), .CK(clk), .Q(\mem[972][3] ) );
  DFF_X1 \mem_reg[972][2]  ( .D(n9022), .CK(clk), .Q(\mem[972][2] ) );
  DFF_X1 \mem_reg[972][1]  ( .D(n9023), .CK(clk), .Q(\mem[972][1] ) );
  DFF_X1 \mem_reg[972][0]  ( .D(n9024), .CK(clk), .Q(\mem[972][0] ) );
  DFF_X1 \mem_reg[971][7]  ( .D(n9025), .CK(clk), .Q(\mem[971][7] ) );
  DFF_X1 \mem_reg[971][6]  ( .D(n9026), .CK(clk), .Q(\mem[971][6] ) );
  DFF_X1 \mem_reg[971][5]  ( .D(n9027), .CK(clk), .Q(\mem[971][5] ) );
  DFF_X1 \mem_reg[971][4]  ( .D(n9028), .CK(clk), .Q(\mem[971][4] ) );
  DFF_X1 \mem_reg[971][3]  ( .D(n9029), .CK(clk), .Q(\mem[971][3] ) );
  DFF_X1 \mem_reg[971][2]  ( .D(n9030), .CK(clk), .Q(\mem[971][2] ) );
  DFF_X1 \mem_reg[971][1]  ( .D(n9031), .CK(clk), .Q(\mem[971][1] ) );
  DFF_X1 \mem_reg[971][0]  ( .D(n9032), .CK(clk), .Q(\mem[971][0] ) );
  DFF_X1 \mem_reg[970][7]  ( .D(n9033), .CK(clk), .Q(\mem[970][7] ) );
  DFF_X1 \mem_reg[970][6]  ( .D(n9034), .CK(clk), .Q(\mem[970][6] ) );
  DFF_X1 \mem_reg[970][5]  ( .D(n9035), .CK(clk), .Q(\mem[970][5] ) );
  DFF_X1 \mem_reg[970][4]  ( .D(n9036), .CK(clk), .Q(\mem[970][4] ) );
  DFF_X1 \mem_reg[970][3]  ( .D(n9037), .CK(clk), .Q(\mem[970][3] ) );
  DFF_X1 \mem_reg[970][2]  ( .D(n9038), .CK(clk), .Q(\mem[970][2] ) );
  DFF_X1 \mem_reg[970][1]  ( .D(n9039), .CK(clk), .Q(\mem[970][1] ) );
  DFF_X1 \mem_reg[970][0]  ( .D(n9040), .CK(clk), .Q(\mem[970][0] ) );
  DFF_X1 \mem_reg[969][7]  ( .D(n9041), .CK(clk), .Q(\mem[969][7] ) );
  DFF_X1 \mem_reg[969][6]  ( .D(n9042), .CK(clk), .Q(\mem[969][6] ) );
  DFF_X1 \mem_reg[969][5]  ( .D(n9043), .CK(clk), .Q(\mem[969][5] ) );
  DFF_X1 \mem_reg[969][4]  ( .D(n9044), .CK(clk), .Q(\mem[969][4] ) );
  DFF_X1 \mem_reg[969][3]  ( .D(n9045), .CK(clk), .Q(\mem[969][3] ) );
  DFF_X1 \mem_reg[969][2]  ( .D(n9046), .CK(clk), .Q(\mem[969][2] ) );
  DFF_X1 \mem_reg[969][1]  ( .D(n9047), .CK(clk), .Q(\mem[969][1] ) );
  DFF_X1 \mem_reg[969][0]  ( .D(n9048), .CK(clk), .Q(\mem[969][0] ) );
  DFF_X1 \mem_reg[968][7]  ( .D(n9049), .CK(clk), .Q(\mem[968][7] ) );
  DFF_X1 \mem_reg[968][6]  ( .D(n9050), .CK(clk), .Q(\mem[968][6] ) );
  DFF_X1 \mem_reg[968][5]  ( .D(n9051), .CK(clk), .Q(\mem[968][5] ) );
  DFF_X1 \mem_reg[968][4]  ( .D(n9052), .CK(clk), .Q(\mem[968][4] ) );
  DFF_X1 \mem_reg[968][3]  ( .D(n9053), .CK(clk), .Q(\mem[968][3] ) );
  DFF_X1 \mem_reg[968][2]  ( .D(n9054), .CK(clk), .Q(\mem[968][2] ) );
  DFF_X1 \mem_reg[968][1]  ( .D(n9055), .CK(clk), .Q(\mem[968][1] ) );
  DFF_X1 \mem_reg[968][0]  ( .D(n9056), .CK(clk), .Q(\mem[968][0] ) );
  DFF_X1 \mem_reg[967][7]  ( .D(n9057), .CK(clk), .Q(\mem[967][7] ) );
  DFF_X1 \mem_reg[967][6]  ( .D(n9058), .CK(clk), .Q(\mem[967][6] ) );
  DFF_X1 \mem_reg[967][5]  ( .D(n9059), .CK(clk), .Q(\mem[967][5] ) );
  DFF_X1 \mem_reg[967][4]  ( .D(n9060), .CK(clk), .Q(\mem[967][4] ) );
  DFF_X1 \mem_reg[967][3]  ( .D(n9061), .CK(clk), .Q(\mem[967][3] ) );
  DFF_X1 \mem_reg[967][2]  ( .D(n9062), .CK(clk), .Q(\mem[967][2] ) );
  DFF_X1 \mem_reg[967][1]  ( .D(n9063), .CK(clk), .Q(\mem[967][1] ) );
  DFF_X1 \mem_reg[967][0]  ( .D(n9064), .CK(clk), .Q(\mem[967][0] ) );
  DFF_X1 \mem_reg[966][7]  ( .D(n9065), .CK(clk), .Q(\mem[966][7] ) );
  DFF_X1 \mem_reg[966][6]  ( .D(n9066), .CK(clk), .Q(\mem[966][6] ) );
  DFF_X1 \mem_reg[966][5]  ( .D(n9067), .CK(clk), .Q(\mem[966][5] ) );
  DFF_X1 \mem_reg[966][4]  ( .D(n9068), .CK(clk), .Q(\mem[966][4] ) );
  DFF_X1 \mem_reg[966][3]  ( .D(n9069), .CK(clk), .Q(\mem[966][3] ) );
  DFF_X1 \mem_reg[966][2]  ( .D(n9070), .CK(clk), .Q(\mem[966][2] ) );
  DFF_X1 \mem_reg[966][1]  ( .D(n9071), .CK(clk), .Q(\mem[966][1] ) );
  DFF_X1 \mem_reg[966][0]  ( .D(n9072), .CK(clk), .Q(\mem[966][0] ) );
  DFF_X1 \mem_reg[965][7]  ( .D(n9073), .CK(clk), .Q(\mem[965][7] ) );
  DFF_X1 \mem_reg[965][6]  ( .D(n9074), .CK(clk), .Q(\mem[965][6] ) );
  DFF_X1 \mem_reg[965][5]  ( .D(n9075), .CK(clk), .Q(\mem[965][5] ) );
  DFF_X1 \mem_reg[965][4]  ( .D(n9076), .CK(clk), .Q(\mem[965][4] ) );
  DFF_X1 \mem_reg[965][3]  ( .D(n9077), .CK(clk), .Q(\mem[965][3] ) );
  DFF_X1 \mem_reg[965][2]  ( .D(n9078), .CK(clk), .Q(\mem[965][2] ) );
  DFF_X1 \mem_reg[965][1]  ( .D(n9079), .CK(clk), .Q(\mem[965][1] ) );
  DFF_X1 \mem_reg[965][0]  ( .D(n9080), .CK(clk), .Q(\mem[965][0] ) );
  DFF_X1 \mem_reg[964][7]  ( .D(n9081), .CK(clk), .Q(\mem[964][7] ) );
  DFF_X1 \mem_reg[964][6]  ( .D(n9082), .CK(clk), .Q(\mem[964][6] ) );
  DFF_X1 \mem_reg[964][5]  ( .D(n9083), .CK(clk), .Q(\mem[964][5] ) );
  DFF_X1 \mem_reg[964][4]  ( .D(n9084), .CK(clk), .Q(\mem[964][4] ) );
  DFF_X1 \mem_reg[964][3]  ( .D(n9085), .CK(clk), .Q(\mem[964][3] ) );
  DFF_X1 \mem_reg[964][2]  ( .D(n9086), .CK(clk), .Q(\mem[964][2] ) );
  DFF_X1 \mem_reg[964][1]  ( .D(n9087), .CK(clk), .Q(\mem[964][1] ) );
  DFF_X1 \mem_reg[964][0]  ( .D(n9088), .CK(clk), .Q(\mem[964][0] ) );
  DFF_X1 \mem_reg[963][7]  ( .D(n9089), .CK(clk), .Q(\mem[963][7] ) );
  DFF_X1 \mem_reg[963][6]  ( .D(n9090), .CK(clk), .Q(\mem[963][6] ) );
  DFF_X1 \mem_reg[963][5]  ( .D(n9091), .CK(clk), .Q(\mem[963][5] ) );
  DFF_X1 \mem_reg[963][4]  ( .D(n9092), .CK(clk), .Q(\mem[963][4] ) );
  DFF_X1 \mem_reg[963][3]  ( .D(n9093), .CK(clk), .Q(\mem[963][3] ) );
  DFF_X1 \mem_reg[963][2]  ( .D(n9094), .CK(clk), .Q(\mem[963][2] ) );
  DFF_X1 \mem_reg[963][1]  ( .D(n9095), .CK(clk), .Q(\mem[963][1] ) );
  DFF_X1 \mem_reg[963][0]  ( .D(n9096), .CK(clk), .Q(\mem[963][0] ) );
  DFF_X1 \mem_reg[962][7]  ( .D(n9097), .CK(clk), .Q(\mem[962][7] ) );
  DFF_X1 \mem_reg[962][6]  ( .D(n9098), .CK(clk), .Q(\mem[962][6] ) );
  DFF_X1 \mem_reg[962][5]  ( .D(n9099), .CK(clk), .Q(\mem[962][5] ) );
  DFF_X1 \mem_reg[962][4]  ( .D(n9100), .CK(clk), .Q(\mem[962][4] ) );
  DFF_X1 \mem_reg[962][3]  ( .D(n9101), .CK(clk), .Q(\mem[962][3] ) );
  DFF_X1 \mem_reg[962][2]  ( .D(n9102), .CK(clk), .Q(\mem[962][2] ) );
  DFF_X1 \mem_reg[962][1]  ( .D(n9103), .CK(clk), .Q(\mem[962][1] ) );
  DFF_X1 \mem_reg[962][0]  ( .D(n9104), .CK(clk), .Q(\mem[962][0] ) );
  DFF_X1 \mem_reg[961][7]  ( .D(n9105), .CK(clk), .Q(\mem[961][7] ) );
  DFF_X1 \mem_reg[961][6]  ( .D(n9106), .CK(clk), .Q(\mem[961][6] ) );
  DFF_X1 \mem_reg[961][5]  ( .D(n9107), .CK(clk), .Q(\mem[961][5] ) );
  DFF_X1 \mem_reg[961][4]  ( .D(n9108), .CK(clk), .Q(\mem[961][4] ) );
  DFF_X1 \mem_reg[961][3]  ( .D(n9109), .CK(clk), .Q(\mem[961][3] ) );
  DFF_X1 \mem_reg[961][2]  ( .D(n9110), .CK(clk), .Q(\mem[961][2] ) );
  DFF_X1 \mem_reg[961][1]  ( .D(n9111), .CK(clk), .Q(\mem[961][1] ) );
  DFF_X1 \mem_reg[961][0]  ( .D(n9112), .CK(clk), .Q(\mem[961][0] ) );
  DFF_X1 \mem_reg[960][7]  ( .D(n9113), .CK(clk), .Q(\mem[960][7] ) );
  DFF_X1 \mem_reg[960][6]  ( .D(n9114), .CK(clk), .Q(\mem[960][6] ) );
  DFF_X1 \mem_reg[960][5]  ( .D(n9115), .CK(clk), .Q(\mem[960][5] ) );
  DFF_X1 \mem_reg[960][4]  ( .D(n9116), .CK(clk), .Q(\mem[960][4] ) );
  DFF_X1 \mem_reg[960][3]  ( .D(n9117), .CK(clk), .Q(\mem[960][3] ) );
  DFF_X1 \mem_reg[960][2]  ( .D(n9118), .CK(clk), .Q(\mem[960][2] ) );
  DFF_X1 \mem_reg[960][1]  ( .D(n9119), .CK(clk), .Q(\mem[960][1] ) );
  DFF_X1 \mem_reg[960][0]  ( .D(n9120), .CK(clk), .Q(\mem[960][0] ) );
  DFF_X1 \mem_reg[959][7]  ( .D(n9121), .CK(clk), .Q(\mem[959][7] ) );
  DFF_X1 \mem_reg[959][6]  ( .D(n9122), .CK(clk), .Q(\mem[959][6] ) );
  DFF_X1 \mem_reg[959][5]  ( .D(n9123), .CK(clk), .Q(\mem[959][5] ) );
  DFF_X1 \mem_reg[959][4]  ( .D(n9124), .CK(clk), .Q(\mem[959][4] ) );
  DFF_X1 \mem_reg[959][3]  ( .D(n9125), .CK(clk), .Q(\mem[959][3] ) );
  DFF_X1 \mem_reg[959][2]  ( .D(n9126), .CK(clk), .Q(\mem[959][2] ) );
  DFF_X1 \mem_reg[959][1]  ( .D(n9127), .CK(clk), .Q(\mem[959][1] ) );
  DFF_X1 \mem_reg[959][0]  ( .D(n9128), .CK(clk), .Q(\mem[959][0] ) );
  DFF_X1 \mem_reg[958][7]  ( .D(n9129), .CK(clk), .Q(\mem[958][7] ) );
  DFF_X1 \mem_reg[958][6]  ( .D(n9130), .CK(clk), .Q(\mem[958][6] ) );
  DFF_X1 \mem_reg[958][5]  ( .D(n9131), .CK(clk), .Q(\mem[958][5] ) );
  DFF_X1 \mem_reg[958][4]  ( .D(n9132), .CK(clk), .Q(\mem[958][4] ) );
  DFF_X1 \mem_reg[958][3]  ( .D(n9133), .CK(clk), .Q(\mem[958][3] ) );
  DFF_X1 \mem_reg[958][2]  ( .D(n9134), .CK(clk), .Q(\mem[958][2] ) );
  DFF_X1 \mem_reg[958][1]  ( .D(n9135), .CK(clk), .Q(\mem[958][1] ) );
  DFF_X1 \mem_reg[958][0]  ( .D(n9136), .CK(clk), .Q(\mem[958][0] ) );
  DFF_X1 \mem_reg[957][7]  ( .D(n9137), .CK(clk), .Q(\mem[957][7] ) );
  DFF_X1 \mem_reg[957][6]  ( .D(n9138), .CK(clk), .Q(\mem[957][6] ) );
  DFF_X1 \mem_reg[957][5]  ( .D(n9139), .CK(clk), .Q(\mem[957][5] ) );
  DFF_X1 \mem_reg[957][4]  ( .D(n9140), .CK(clk), .Q(\mem[957][4] ) );
  DFF_X1 \mem_reg[957][3]  ( .D(n9141), .CK(clk), .Q(\mem[957][3] ) );
  DFF_X1 \mem_reg[957][2]  ( .D(n9142), .CK(clk), .Q(\mem[957][2] ) );
  DFF_X1 \mem_reg[957][1]  ( .D(n9143), .CK(clk), .Q(\mem[957][1] ) );
  DFF_X1 \mem_reg[957][0]  ( .D(n9144), .CK(clk), .Q(\mem[957][0] ) );
  DFF_X1 \mem_reg[956][7]  ( .D(n9145), .CK(clk), .Q(\mem[956][7] ) );
  DFF_X1 \mem_reg[956][6]  ( .D(n9146), .CK(clk), .Q(\mem[956][6] ) );
  DFF_X1 \mem_reg[956][5]  ( .D(n9147), .CK(clk), .Q(\mem[956][5] ) );
  DFF_X1 \mem_reg[956][4]  ( .D(n9148), .CK(clk), .Q(\mem[956][4] ) );
  DFF_X1 \mem_reg[956][3]  ( .D(n9149), .CK(clk), .Q(\mem[956][3] ) );
  DFF_X1 \mem_reg[956][2]  ( .D(n9150), .CK(clk), .Q(\mem[956][2] ) );
  DFF_X1 \mem_reg[956][1]  ( .D(n9151), .CK(clk), .Q(\mem[956][1] ) );
  DFF_X1 \mem_reg[956][0]  ( .D(n9152), .CK(clk), .Q(\mem[956][0] ) );
  DFF_X1 \mem_reg[955][7]  ( .D(n9153), .CK(clk), .Q(\mem[955][7] ) );
  DFF_X1 \mem_reg[955][6]  ( .D(n9154), .CK(clk), .Q(\mem[955][6] ) );
  DFF_X1 \mem_reg[955][5]  ( .D(n9155), .CK(clk), .Q(\mem[955][5] ) );
  DFF_X1 \mem_reg[955][4]  ( .D(n9156), .CK(clk), .Q(\mem[955][4] ) );
  DFF_X1 \mem_reg[955][3]  ( .D(n9157), .CK(clk), .Q(\mem[955][3] ) );
  DFF_X1 \mem_reg[955][2]  ( .D(n9158), .CK(clk), .Q(\mem[955][2] ) );
  DFF_X1 \mem_reg[955][1]  ( .D(n9159), .CK(clk), .Q(\mem[955][1] ) );
  DFF_X1 \mem_reg[955][0]  ( .D(n9160), .CK(clk), .Q(\mem[955][0] ) );
  DFF_X1 \mem_reg[954][7]  ( .D(n9161), .CK(clk), .Q(\mem[954][7] ) );
  DFF_X1 \mem_reg[954][6]  ( .D(n9162), .CK(clk), .Q(\mem[954][6] ) );
  DFF_X1 \mem_reg[954][5]  ( .D(n9163), .CK(clk), .Q(\mem[954][5] ) );
  DFF_X1 \mem_reg[954][4]  ( .D(n9164), .CK(clk), .Q(\mem[954][4] ) );
  DFF_X1 \mem_reg[954][3]  ( .D(n9165), .CK(clk), .Q(\mem[954][3] ) );
  DFF_X1 \mem_reg[954][2]  ( .D(n9166), .CK(clk), .Q(\mem[954][2] ) );
  DFF_X1 \mem_reg[954][1]  ( .D(n9167), .CK(clk), .Q(\mem[954][1] ) );
  DFF_X1 \mem_reg[954][0]  ( .D(n9168), .CK(clk), .Q(\mem[954][0] ) );
  DFF_X1 \mem_reg[953][7]  ( .D(n9169), .CK(clk), .Q(\mem[953][7] ) );
  DFF_X1 \mem_reg[953][6]  ( .D(n9170), .CK(clk), .Q(\mem[953][6] ) );
  DFF_X1 \mem_reg[953][5]  ( .D(n9171), .CK(clk), .Q(\mem[953][5] ) );
  DFF_X1 \mem_reg[953][4]  ( .D(n9172), .CK(clk), .Q(\mem[953][4] ) );
  DFF_X1 \mem_reg[953][3]  ( .D(n9173), .CK(clk), .Q(\mem[953][3] ) );
  DFF_X1 \mem_reg[953][2]  ( .D(n9174), .CK(clk), .Q(\mem[953][2] ) );
  DFF_X1 \mem_reg[953][1]  ( .D(n9175), .CK(clk), .Q(\mem[953][1] ) );
  DFF_X1 \mem_reg[953][0]  ( .D(n9176), .CK(clk), .Q(\mem[953][0] ) );
  DFF_X1 \mem_reg[952][7]  ( .D(n9177), .CK(clk), .Q(\mem[952][7] ) );
  DFF_X1 \mem_reg[952][6]  ( .D(n9178), .CK(clk), .Q(\mem[952][6] ) );
  DFF_X1 \mem_reg[952][5]  ( .D(n9179), .CK(clk), .Q(\mem[952][5] ) );
  DFF_X1 \mem_reg[952][4]  ( .D(n9180), .CK(clk), .Q(\mem[952][4] ) );
  DFF_X1 \mem_reg[952][3]  ( .D(n9181), .CK(clk), .Q(\mem[952][3] ) );
  DFF_X1 \mem_reg[952][2]  ( .D(n9182), .CK(clk), .Q(\mem[952][2] ) );
  DFF_X1 \mem_reg[952][1]  ( .D(n9183), .CK(clk), .Q(\mem[952][1] ) );
  DFF_X1 \mem_reg[952][0]  ( .D(n9184), .CK(clk), .Q(\mem[952][0] ) );
  DFF_X1 \mem_reg[951][7]  ( .D(n9185), .CK(clk), .Q(\mem[951][7] ) );
  DFF_X1 \mem_reg[951][6]  ( .D(n9186), .CK(clk), .Q(\mem[951][6] ) );
  DFF_X1 \mem_reg[951][5]  ( .D(n9187), .CK(clk), .Q(\mem[951][5] ) );
  DFF_X1 \mem_reg[951][4]  ( .D(n9188), .CK(clk), .Q(\mem[951][4] ) );
  DFF_X1 \mem_reg[951][3]  ( .D(n9189), .CK(clk), .Q(\mem[951][3] ) );
  DFF_X1 \mem_reg[951][2]  ( .D(n9190), .CK(clk), .Q(\mem[951][2] ) );
  DFF_X1 \mem_reg[951][1]  ( .D(n9191), .CK(clk), .Q(\mem[951][1] ) );
  DFF_X1 \mem_reg[951][0]  ( .D(n9192), .CK(clk), .Q(\mem[951][0] ) );
  DFF_X1 \mem_reg[950][7]  ( .D(n9193), .CK(clk), .Q(\mem[950][7] ) );
  DFF_X1 \mem_reg[950][6]  ( .D(n9194), .CK(clk), .Q(\mem[950][6] ) );
  DFF_X1 \mem_reg[950][5]  ( .D(n9195), .CK(clk), .Q(\mem[950][5] ) );
  DFF_X1 \mem_reg[950][4]  ( .D(n9196), .CK(clk), .Q(\mem[950][4] ) );
  DFF_X1 \mem_reg[950][3]  ( .D(n9197), .CK(clk), .Q(\mem[950][3] ) );
  DFF_X1 \mem_reg[950][2]  ( .D(n9198), .CK(clk), .Q(\mem[950][2] ) );
  DFF_X1 \mem_reg[950][1]  ( .D(n9199), .CK(clk), .Q(\mem[950][1] ) );
  DFF_X1 \mem_reg[950][0]  ( .D(n9200), .CK(clk), .Q(\mem[950][0] ) );
  DFF_X1 \mem_reg[949][7]  ( .D(n9201), .CK(clk), .Q(\mem[949][7] ) );
  DFF_X1 \mem_reg[949][6]  ( .D(n9202), .CK(clk), .Q(\mem[949][6] ) );
  DFF_X1 \mem_reg[949][5]  ( .D(n9203), .CK(clk), .Q(\mem[949][5] ) );
  DFF_X1 \mem_reg[949][4]  ( .D(n9204), .CK(clk), .Q(\mem[949][4] ) );
  DFF_X1 \mem_reg[949][3]  ( .D(n9205), .CK(clk), .Q(\mem[949][3] ) );
  DFF_X1 \mem_reg[949][2]  ( .D(n9206), .CK(clk), .Q(\mem[949][2] ) );
  DFF_X1 \mem_reg[949][1]  ( .D(n9207), .CK(clk), .Q(\mem[949][1] ) );
  DFF_X1 \mem_reg[949][0]  ( .D(n9208), .CK(clk), .Q(\mem[949][0] ) );
  DFF_X1 \mem_reg[948][7]  ( .D(n9209), .CK(clk), .Q(\mem[948][7] ) );
  DFF_X1 \mem_reg[948][6]  ( .D(n9210), .CK(clk), .Q(\mem[948][6] ) );
  DFF_X1 \mem_reg[948][5]  ( .D(n9211), .CK(clk), .Q(\mem[948][5] ) );
  DFF_X1 \mem_reg[948][4]  ( .D(n9212), .CK(clk), .Q(\mem[948][4] ) );
  DFF_X1 \mem_reg[948][3]  ( .D(n9213), .CK(clk), .Q(\mem[948][3] ) );
  DFF_X1 \mem_reg[948][2]  ( .D(n9214), .CK(clk), .Q(\mem[948][2] ) );
  DFF_X1 \mem_reg[948][1]  ( .D(n9215), .CK(clk), .Q(\mem[948][1] ) );
  DFF_X1 \mem_reg[948][0]  ( .D(n9216), .CK(clk), .Q(\mem[948][0] ) );
  DFF_X1 \mem_reg[947][7]  ( .D(n9217), .CK(clk), .Q(\mem[947][7] ) );
  DFF_X1 \mem_reg[947][6]  ( .D(n9218), .CK(clk), .Q(\mem[947][6] ) );
  DFF_X1 \mem_reg[947][5]  ( .D(n9219), .CK(clk), .Q(\mem[947][5] ) );
  DFF_X1 \mem_reg[947][4]  ( .D(n9220), .CK(clk), .Q(\mem[947][4] ) );
  DFF_X1 \mem_reg[947][3]  ( .D(n9221), .CK(clk), .Q(\mem[947][3] ) );
  DFF_X1 \mem_reg[947][2]  ( .D(n9222), .CK(clk), .Q(\mem[947][2] ) );
  DFF_X1 \mem_reg[947][1]  ( .D(n18529), .CK(clk), .Q(\mem[947][1] ) );
  DFF_X1 \mem_reg[947][0]  ( .D(n18530), .CK(clk), .Q(\mem[947][0] ) );
  DFF_X1 \mem_reg[946][7]  ( .D(n18531), .CK(clk), .Q(\mem[946][7] ) );
  DFF_X1 \mem_reg[946][6]  ( .D(n18532), .CK(clk), .Q(\mem[946][6] ) );
  DFF_X1 \mem_reg[946][5]  ( .D(n18533), .CK(clk), .Q(\mem[946][5] ) );
  DFF_X1 \mem_reg[946][4]  ( .D(n18534), .CK(clk), .Q(\mem[946][4] ) );
  DFF_X1 \mem_reg[946][3]  ( .D(n18535), .CK(clk), .Q(\mem[946][3] ) );
  DFF_X1 \mem_reg[946][2]  ( .D(n18536), .CK(clk), .Q(\mem[946][2] ) );
  DFF_X1 \mem_reg[946][1]  ( .D(n18537), .CK(clk), .Q(\mem[946][1] ) );
  DFF_X1 \mem_reg[946][0]  ( .D(n18538), .CK(clk), .Q(\mem[946][0] ) );
  DFF_X1 \mem_reg[945][7]  ( .D(n18539), .CK(clk), .Q(\mem[945][7] ) );
  DFF_X1 \mem_reg[945][6]  ( .D(n18540), .CK(clk), .Q(\mem[945][6] ) );
  DFF_X1 \mem_reg[945][5]  ( .D(n18541), .CK(clk), .Q(\mem[945][5] ) );
  DFF_X1 \mem_reg[945][4]  ( .D(n18542), .CK(clk), .Q(\mem[945][4] ) );
  DFF_X1 \mem_reg[945][3]  ( .D(n18543), .CK(clk), .Q(\mem[945][3] ) );
  DFF_X1 \mem_reg[945][2]  ( .D(n18544), .CK(clk), .Q(\mem[945][2] ) );
  DFF_X1 \mem_reg[945][1]  ( .D(n18545), .CK(clk), .Q(\mem[945][1] ) );
  DFF_X1 \mem_reg[945][0]  ( .D(n18546), .CK(clk), .Q(\mem[945][0] ) );
  DFF_X1 \mem_reg[944][7]  ( .D(n18547), .CK(clk), .Q(\mem[944][7] ) );
  DFF_X1 \mem_reg[944][6]  ( .D(n18548), .CK(clk), .Q(\mem[944][6] ) );
  DFF_X1 \mem_reg[944][5]  ( .D(n18549), .CK(clk), .Q(\mem[944][5] ) );
  DFF_X1 \mem_reg[944][4]  ( .D(n18550), .CK(clk), .Q(\mem[944][4] ) );
  DFF_X1 \mem_reg[944][3]  ( .D(n18551), .CK(clk), .Q(\mem[944][3] ) );
  DFF_X1 \mem_reg[944][2]  ( .D(n18552), .CK(clk), .Q(\mem[944][2] ) );
  DFF_X1 \mem_reg[944][1]  ( .D(n18553), .CK(clk), .Q(\mem[944][1] ) );
  DFF_X1 \mem_reg[944][0]  ( .D(n18554), .CK(clk), .Q(\mem[944][0] ) );
  DFF_X1 \mem_reg[943][7]  ( .D(n18555), .CK(clk), .Q(\mem[943][7] ) );
  DFF_X1 \mem_reg[943][6]  ( .D(n18556), .CK(clk), .Q(\mem[943][6] ) );
  DFF_X1 \mem_reg[943][5]  ( .D(n18557), .CK(clk), .Q(\mem[943][5] ) );
  DFF_X1 \mem_reg[943][4]  ( .D(n18558), .CK(clk), .Q(\mem[943][4] ) );
  DFF_X1 \mem_reg[943][3]  ( .D(n18559), .CK(clk), .Q(\mem[943][3] ) );
  DFF_X1 \mem_reg[943][2]  ( .D(n18560), .CK(clk), .Q(\mem[943][2] ) );
  DFF_X1 \mem_reg[943][1]  ( .D(n18561), .CK(clk), .Q(\mem[943][1] ) );
  DFF_X1 \mem_reg[943][0]  ( .D(n18562), .CK(clk), .Q(\mem[943][0] ) );
  DFF_X1 \mem_reg[942][7]  ( .D(n18563), .CK(clk), .Q(\mem[942][7] ) );
  DFF_X1 \mem_reg[942][6]  ( .D(n18564), .CK(clk), .Q(\mem[942][6] ) );
  DFF_X1 \mem_reg[942][5]  ( .D(n18565), .CK(clk), .Q(\mem[942][5] ) );
  DFF_X1 \mem_reg[942][4]  ( .D(n18566), .CK(clk), .Q(\mem[942][4] ) );
  DFF_X1 \mem_reg[942][3]  ( .D(n18567), .CK(clk), .Q(\mem[942][3] ) );
  DFF_X1 \mem_reg[942][2]  ( .D(n18568), .CK(clk), .Q(\mem[942][2] ) );
  DFF_X1 \mem_reg[942][1]  ( .D(n18569), .CK(clk), .Q(\mem[942][1] ) );
  DFF_X1 \mem_reg[942][0]  ( .D(n18570), .CK(clk), .Q(\mem[942][0] ) );
  DFF_X1 \mem_reg[941][7]  ( .D(n18571), .CK(clk), .Q(\mem[941][7] ) );
  DFF_X1 \mem_reg[941][6]  ( .D(n18572), .CK(clk), .Q(\mem[941][6] ) );
  DFF_X1 \mem_reg[941][5]  ( .D(n18573), .CK(clk), .Q(\mem[941][5] ) );
  DFF_X1 \mem_reg[941][4]  ( .D(n18574), .CK(clk), .Q(\mem[941][4] ) );
  DFF_X1 \mem_reg[941][3]  ( .D(n18575), .CK(clk), .Q(\mem[941][3] ) );
  DFF_X1 \mem_reg[941][2]  ( .D(n18576), .CK(clk), .Q(\mem[941][2] ) );
  DFF_X1 \mem_reg[941][1]  ( .D(n18577), .CK(clk), .Q(\mem[941][1] ) );
  DFF_X1 \mem_reg[941][0]  ( .D(n18578), .CK(clk), .Q(\mem[941][0] ) );
  DFF_X1 \mem_reg[940][7]  ( .D(n18579), .CK(clk), .Q(\mem[940][7] ) );
  DFF_X1 \mem_reg[940][6]  ( .D(n18580), .CK(clk), .Q(\mem[940][6] ) );
  DFF_X1 \mem_reg[940][5]  ( .D(n18581), .CK(clk), .Q(\mem[940][5] ) );
  DFF_X1 \mem_reg[940][4]  ( .D(n18582), .CK(clk), .Q(\mem[940][4] ) );
  DFF_X1 \mem_reg[940][3]  ( .D(n18583), .CK(clk), .Q(\mem[940][3] ) );
  DFF_X1 \mem_reg[940][2]  ( .D(n18584), .CK(clk), .Q(\mem[940][2] ) );
  DFF_X1 \mem_reg[940][1]  ( .D(n18585), .CK(clk), .Q(\mem[940][1] ) );
  DFF_X1 \mem_reg[940][0]  ( .D(n18586), .CK(clk), .Q(\mem[940][0] ) );
  DFF_X1 \mem_reg[939][7]  ( .D(n18587), .CK(clk), .Q(\mem[939][7] ) );
  DFF_X1 \mem_reg[939][6]  ( .D(n18588), .CK(clk), .Q(\mem[939][6] ) );
  DFF_X1 \mem_reg[939][5]  ( .D(n18589), .CK(clk), .Q(\mem[939][5] ) );
  DFF_X1 \mem_reg[939][4]  ( .D(n18590), .CK(clk), .Q(\mem[939][4] ) );
  DFF_X1 \mem_reg[939][3]  ( .D(n18591), .CK(clk), .Q(\mem[939][3] ) );
  DFF_X1 \mem_reg[939][2]  ( .D(n18592), .CK(clk), .Q(\mem[939][2] ) );
  DFF_X1 \mem_reg[939][1]  ( .D(n18593), .CK(clk), .Q(\mem[939][1] ) );
  DFF_X1 \mem_reg[939][0]  ( .D(n18594), .CK(clk), .Q(\mem[939][0] ) );
  DFF_X1 \mem_reg[938][7]  ( .D(n18595), .CK(clk), .Q(\mem[938][7] ) );
  DFF_X1 \mem_reg[938][6]  ( .D(n18596), .CK(clk), .Q(\mem[938][6] ) );
  DFF_X1 \mem_reg[938][5]  ( .D(n18597), .CK(clk), .Q(\mem[938][5] ) );
  DFF_X1 \mem_reg[938][4]  ( .D(n18598), .CK(clk), .Q(\mem[938][4] ) );
  DFF_X1 \mem_reg[938][3]  ( .D(n18599), .CK(clk), .Q(\mem[938][3] ) );
  DFF_X1 \mem_reg[938][2]  ( .D(n18600), .CK(clk), .Q(\mem[938][2] ) );
  DFF_X1 \mem_reg[938][1]  ( .D(n18601), .CK(clk), .Q(\mem[938][1] ) );
  DFF_X1 \mem_reg[938][0]  ( .D(n18602), .CK(clk), .Q(\mem[938][0] ) );
  DFF_X1 \mem_reg[937][7]  ( .D(n18603), .CK(clk), .Q(\mem[937][7] ) );
  DFF_X1 \mem_reg[937][6]  ( .D(n18604), .CK(clk), .Q(\mem[937][6] ) );
  DFF_X1 \mem_reg[937][5]  ( .D(n18605), .CK(clk), .Q(\mem[937][5] ) );
  DFF_X1 \mem_reg[937][4]  ( .D(n18606), .CK(clk), .Q(\mem[937][4] ) );
  DFF_X1 \mem_reg[937][3]  ( .D(n18607), .CK(clk), .Q(\mem[937][3] ) );
  DFF_X1 \mem_reg[937][2]  ( .D(n18608), .CK(clk), .Q(\mem[937][2] ) );
  DFF_X1 \mem_reg[937][1]  ( .D(n18609), .CK(clk), .Q(\mem[937][1] ) );
  DFF_X1 \mem_reg[937][0]  ( .D(n18610), .CK(clk), .Q(\mem[937][0] ) );
  DFF_X1 \mem_reg[936][7]  ( .D(n18611), .CK(clk), .Q(\mem[936][7] ) );
  DFF_X1 \mem_reg[936][6]  ( .D(n18612), .CK(clk), .Q(\mem[936][6] ) );
  DFF_X1 \mem_reg[936][5]  ( .D(n18613), .CK(clk), .Q(\mem[936][5] ) );
  DFF_X1 \mem_reg[936][4]  ( .D(n18614), .CK(clk), .Q(\mem[936][4] ) );
  DFF_X1 \mem_reg[936][3]  ( .D(n18615), .CK(clk), .Q(\mem[936][3] ) );
  DFF_X1 \mem_reg[936][2]  ( .D(n18616), .CK(clk), .Q(\mem[936][2] ) );
  DFF_X1 \mem_reg[936][1]  ( .D(n18617), .CK(clk), .Q(\mem[936][1] ) );
  DFF_X1 \mem_reg[936][0]  ( .D(n18618), .CK(clk), .Q(\mem[936][0] ) );
  DFF_X1 \mem_reg[935][7]  ( .D(n18619), .CK(clk), .Q(\mem[935][7] ) );
  DFF_X1 \mem_reg[935][6]  ( .D(n18620), .CK(clk), .Q(\mem[935][6] ) );
  DFF_X1 \mem_reg[935][5]  ( .D(n18621), .CK(clk), .Q(\mem[935][5] ) );
  DFF_X1 \mem_reg[935][4]  ( .D(n18622), .CK(clk), .Q(\mem[935][4] ) );
  DFF_X1 \mem_reg[935][3]  ( .D(n18623), .CK(clk), .Q(\mem[935][3] ) );
  DFF_X1 \mem_reg[935][2]  ( .D(n18624), .CK(clk), .Q(\mem[935][2] ) );
  DFF_X1 \mem_reg[935][1]  ( .D(n18625), .CK(clk), .Q(\mem[935][1] ) );
  DFF_X1 \mem_reg[935][0]  ( .D(n18626), .CK(clk), .Q(\mem[935][0] ) );
  DFF_X1 \mem_reg[934][7]  ( .D(n18627), .CK(clk), .Q(\mem[934][7] ) );
  DFF_X1 \mem_reg[934][6]  ( .D(n18628), .CK(clk), .Q(\mem[934][6] ) );
  DFF_X1 \mem_reg[934][5]  ( .D(n18629), .CK(clk), .Q(\mem[934][5] ) );
  DFF_X1 \mem_reg[934][4]  ( .D(n18630), .CK(clk), .Q(\mem[934][4] ) );
  DFF_X1 \mem_reg[934][3]  ( .D(n18631), .CK(clk), .Q(\mem[934][3] ) );
  DFF_X1 \mem_reg[934][2]  ( .D(n18632), .CK(clk), .Q(\mem[934][2] ) );
  DFF_X1 \mem_reg[934][1]  ( .D(n18633), .CK(clk), .Q(\mem[934][1] ) );
  DFF_X1 \mem_reg[934][0]  ( .D(n18634), .CK(clk), .Q(\mem[934][0] ) );
  DFF_X1 \mem_reg[933][7]  ( .D(n18635), .CK(clk), .Q(\mem[933][7] ) );
  DFF_X1 \mem_reg[933][6]  ( .D(n18636), .CK(clk), .Q(\mem[933][6] ) );
  DFF_X1 \mem_reg[933][5]  ( .D(n18637), .CK(clk), .Q(\mem[933][5] ) );
  DFF_X1 \mem_reg[933][4]  ( .D(n18638), .CK(clk), .Q(\mem[933][4] ) );
  DFF_X1 \mem_reg[933][3]  ( .D(n18639), .CK(clk), .Q(\mem[933][3] ) );
  DFF_X1 \mem_reg[933][2]  ( .D(n18640), .CK(clk), .Q(\mem[933][2] ) );
  DFF_X1 \mem_reg[933][1]  ( .D(n18641), .CK(clk), .Q(\mem[933][1] ) );
  DFF_X1 \mem_reg[933][0]  ( .D(n18642), .CK(clk), .Q(\mem[933][0] ) );
  DFF_X1 \mem_reg[932][7]  ( .D(n18643), .CK(clk), .Q(\mem[932][7] ) );
  DFF_X1 \mem_reg[932][6]  ( .D(n18644), .CK(clk), .Q(\mem[932][6] ) );
  DFF_X1 \mem_reg[932][5]  ( .D(n18645), .CK(clk), .Q(\mem[932][5] ) );
  DFF_X1 \mem_reg[932][4]  ( .D(n18646), .CK(clk), .Q(\mem[932][4] ) );
  DFF_X1 \mem_reg[932][3]  ( .D(n18647), .CK(clk), .Q(\mem[932][3] ) );
  DFF_X1 \mem_reg[932][2]  ( .D(n18648), .CK(clk), .Q(\mem[932][2] ) );
  DFF_X1 \mem_reg[932][1]  ( .D(n18649), .CK(clk), .Q(\mem[932][1] ) );
  DFF_X1 \mem_reg[932][0]  ( .D(n18650), .CK(clk), .Q(\mem[932][0] ) );
  DFF_X1 \mem_reg[931][7]  ( .D(n18651), .CK(clk), .Q(\mem[931][7] ) );
  DFF_X1 \mem_reg[931][6]  ( .D(n18652), .CK(clk), .Q(\mem[931][6] ) );
  DFF_X1 \mem_reg[931][5]  ( .D(n18653), .CK(clk), .Q(\mem[931][5] ) );
  DFF_X1 \mem_reg[931][4]  ( .D(n18654), .CK(clk), .Q(\mem[931][4] ) );
  DFF_X1 \mem_reg[931][3]  ( .D(n18655), .CK(clk), .Q(\mem[931][3] ) );
  DFF_X1 \mem_reg[931][2]  ( .D(n18656), .CK(clk), .Q(\mem[931][2] ) );
  DFF_X1 \mem_reg[931][1]  ( .D(n18657), .CK(clk), .Q(\mem[931][1] ) );
  DFF_X1 \mem_reg[931][0]  ( .D(n18658), .CK(clk), .Q(\mem[931][0] ) );
  DFF_X1 \mem_reg[930][7]  ( .D(n18659), .CK(clk), .Q(\mem[930][7] ) );
  DFF_X1 \mem_reg[930][6]  ( .D(n18660), .CK(clk), .Q(\mem[930][6] ) );
  DFF_X1 \mem_reg[930][5]  ( .D(n18661), .CK(clk), .Q(\mem[930][5] ) );
  DFF_X1 \mem_reg[930][4]  ( .D(n18662), .CK(clk), .Q(\mem[930][4] ) );
  DFF_X1 \mem_reg[930][3]  ( .D(n18663), .CK(clk), .Q(\mem[930][3] ) );
  DFF_X1 \mem_reg[930][2]  ( .D(n18664), .CK(clk), .Q(\mem[930][2] ) );
  DFF_X1 \mem_reg[930][1]  ( .D(n18665), .CK(clk), .Q(\mem[930][1] ) );
  DFF_X1 \mem_reg[930][0]  ( .D(n18666), .CK(clk), .Q(\mem[930][0] ) );
  DFF_X1 \mem_reg[929][7]  ( .D(n18667), .CK(clk), .Q(\mem[929][7] ) );
  DFF_X1 \mem_reg[929][6]  ( .D(n18668), .CK(clk), .Q(\mem[929][6] ) );
  DFF_X1 \mem_reg[929][5]  ( .D(n18669), .CK(clk), .Q(\mem[929][5] ) );
  DFF_X1 \mem_reg[929][4]  ( .D(n18670), .CK(clk), .Q(\mem[929][4] ) );
  DFF_X1 \mem_reg[929][3]  ( .D(n18671), .CK(clk), .Q(\mem[929][3] ) );
  DFF_X1 \mem_reg[929][2]  ( .D(n18672), .CK(clk), .Q(\mem[929][2] ) );
  DFF_X1 \mem_reg[929][1]  ( .D(n18673), .CK(clk), .Q(\mem[929][1] ) );
  DFF_X1 \mem_reg[929][0]  ( .D(n18674), .CK(clk), .Q(\mem[929][0] ) );
  DFF_X1 \mem_reg[928][7]  ( .D(n18675), .CK(clk), .Q(\mem[928][7] ) );
  DFF_X1 \mem_reg[928][6]  ( .D(n18676), .CK(clk), .Q(\mem[928][6] ) );
  DFF_X1 \mem_reg[928][5]  ( .D(n18677), .CK(clk), .Q(\mem[928][5] ) );
  DFF_X1 \mem_reg[928][4]  ( .D(n18678), .CK(clk), .Q(\mem[928][4] ) );
  DFF_X1 \mem_reg[928][3]  ( .D(n18679), .CK(clk), .Q(\mem[928][3] ) );
  DFF_X1 \mem_reg[928][2]  ( .D(n18680), .CK(clk), .Q(\mem[928][2] ) );
  DFF_X1 \mem_reg[928][1]  ( .D(n18681), .CK(clk), .Q(\mem[928][1] ) );
  DFF_X1 \mem_reg[928][0]  ( .D(n18682), .CK(clk), .Q(\mem[928][0] ) );
  DFF_X1 \mem_reg[927][7]  ( .D(n18683), .CK(clk), .Q(\mem[927][7] ) );
  DFF_X1 \mem_reg[927][6]  ( .D(n18684), .CK(clk), .Q(\mem[927][6] ) );
  DFF_X1 \mem_reg[927][5]  ( .D(n18685), .CK(clk), .Q(\mem[927][5] ) );
  DFF_X1 \mem_reg[927][4]  ( .D(n18686), .CK(clk), .Q(\mem[927][4] ) );
  DFF_X1 \mem_reg[927][3]  ( .D(n18687), .CK(clk), .Q(\mem[927][3] ) );
  DFF_X1 \mem_reg[927][2]  ( .D(n18688), .CK(clk), .Q(\mem[927][2] ) );
  DFF_X1 \mem_reg[927][1]  ( .D(n18689), .CK(clk), .Q(\mem[927][1] ) );
  DFF_X1 \mem_reg[927][0]  ( .D(n18690), .CK(clk), .Q(\mem[927][0] ) );
  DFF_X1 \mem_reg[926][7]  ( .D(n18691), .CK(clk), .Q(\mem[926][7] ) );
  DFF_X1 \mem_reg[926][6]  ( .D(n18692), .CK(clk), .Q(\mem[926][6] ) );
  DFF_X1 \mem_reg[926][5]  ( .D(n18693), .CK(clk), .Q(\mem[926][5] ) );
  DFF_X1 \mem_reg[926][4]  ( .D(n18694), .CK(clk), .Q(\mem[926][4] ) );
  DFF_X1 \mem_reg[926][3]  ( .D(n18695), .CK(clk), .Q(\mem[926][3] ) );
  DFF_X1 \mem_reg[926][2]  ( .D(n18696), .CK(clk), .Q(\mem[926][2] ) );
  DFF_X1 \mem_reg[926][1]  ( .D(n18697), .CK(clk), .Q(\mem[926][1] ) );
  DFF_X1 \mem_reg[926][0]  ( .D(n18698), .CK(clk), .Q(\mem[926][0] ) );
  DFF_X1 \mem_reg[925][7]  ( .D(n18699), .CK(clk), .Q(\mem[925][7] ) );
  DFF_X1 \mem_reg[925][6]  ( .D(n18700), .CK(clk), .Q(\mem[925][6] ) );
  DFF_X1 \mem_reg[925][5]  ( .D(n18701), .CK(clk), .Q(\mem[925][5] ) );
  DFF_X1 \mem_reg[925][4]  ( .D(n18702), .CK(clk), .Q(\mem[925][4] ) );
  DFF_X1 \mem_reg[925][3]  ( .D(n18703), .CK(clk), .Q(\mem[925][3] ) );
  DFF_X1 \mem_reg[925][2]  ( .D(n18704), .CK(clk), .Q(\mem[925][2] ) );
  DFF_X1 \mem_reg[925][1]  ( .D(n18705), .CK(clk), .Q(\mem[925][1] ) );
  DFF_X1 \mem_reg[925][0]  ( .D(n18706), .CK(clk), .Q(\mem[925][0] ) );
  DFF_X1 \mem_reg[924][7]  ( .D(n18707), .CK(clk), .Q(\mem[924][7] ) );
  DFF_X1 \mem_reg[924][6]  ( .D(n18708), .CK(clk), .Q(\mem[924][6] ) );
  DFF_X1 \mem_reg[924][5]  ( .D(n18709), .CK(clk), .Q(\mem[924][5] ) );
  DFF_X1 \mem_reg[924][4]  ( .D(n18710), .CK(clk), .Q(\mem[924][4] ) );
  DFF_X1 \mem_reg[924][3]  ( .D(n18711), .CK(clk), .Q(\mem[924][3] ) );
  DFF_X1 \mem_reg[924][2]  ( .D(n18712), .CK(clk), .Q(\mem[924][2] ) );
  DFF_X1 \mem_reg[924][1]  ( .D(n18713), .CK(clk), .Q(\mem[924][1] ) );
  DFF_X1 \mem_reg[924][0]  ( .D(n18714), .CK(clk), .Q(\mem[924][0] ) );
  DFF_X1 \mem_reg[923][7]  ( .D(n18715), .CK(clk), .Q(\mem[923][7] ) );
  DFF_X1 \mem_reg[923][6]  ( .D(n18716), .CK(clk), .Q(\mem[923][6] ) );
  DFF_X1 \mem_reg[923][5]  ( .D(n18717), .CK(clk), .Q(\mem[923][5] ) );
  DFF_X1 \mem_reg[923][4]  ( .D(n18718), .CK(clk), .Q(\mem[923][4] ) );
  DFF_X1 \mem_reg[923][3]  ( .D(n18719), .CK(clk), .Q(\mem[923][3] ) );
  DFF_X1 \mem_reg[923][2]  ( .D(n18720), .CK(clk), .Q(\mem[923][2] ) );
  DFF_X1 \mem_reg[923][1]  ( .D(n18721), .CK(clk), .Q(\mem[923][1] ) );
  DFF_X1 \mem_reg[923][0]  ( .D(n18722), .CK(clk), .Q(\mem[923][0] ) );
  DFF_X1 \mem_reg[922][7]  ( .D(n18723), .CK(clk), .Q(\mem[922][7] ) );
  DFF_X1 \mem_reg[922][6]  ( .D(n18724), .CK(clk), .Q(\mem[922][6] ) );
  DFF_X1 \mem_reg[922][5]  ( .D(n18725), .CK(clk), .Q(\mem[922][5] ) );
  DFF_X1 \mem_reg[922][4]  ( .D(n18726), .CK(clk), .Q(\mem[922][4] ) );
  DFF_X1 \mem_reg[922][3]  ( .D(n18727), .CK(clk), .Q(\mem[922][3] ) );
  DFF_X1 \mem_reg[922][2]  ( .D(n18728), .CK(clk), .Q(\mem[922][2] ) );
  DFF_X1 \mem_reg[922][1]  ( .D(n18729), .CK(clk), .Q(\mem[922][1] ) );
  DFF_X1 \mem_reg[922][0]  ( .D(n18730), .CK(clk), .Q(\mem[922][0] ) );
  DFF_X1 \mem_reg[921][7]  ( .D(n18731), .CK(clk), .Q(\mem[921][7] ) );
  DFF_X1 \mem_reg[921][6]  ( .D(n18732), .CK(clk), .Q(\mem[921][6] ) );
  DFF_X1 \mem_reg[921][5]  ( .D(n18733), .CK(clk), .Q(\mem[921][5] ) );
  DFF_X1 \mem_reg[921][4]  ( .D(n18734), .CK(clk), .Q(\mem[921][4] ) );
  DFF_X1 \mem_reg[921][3]  ( .D(n18735), .CK(clk), .Q(\mem[921][3] ) );
  DFF_X1 \mem_reg[921][2]  ( .D(n18736), .CK(clk), .Q(\mem[921][2] ) );
  DFF_X1 \mem_reg[921][1]  ( .D(n18737), .CK(clk), .Q(\mem[921][1] ) );
  DFF_X1 \mem_reg[921][0]  ( .D(n18738), .CK(clk), .Q(\mem[921][0] ) );
  DFF_X1 \mem_reg[920][7]  ( .D(n18739), .CK(clk), .Q(\mem[920][7] ) );
  DFF_X1 \mem_reg[920][6]  ( .D(n18740), .CK(clk), .Q(\mem[920][6] ) );
  DFF_X1 \mem_reg[920][5]  ( .D(n18741), .CK(clk), .Q(\mem[920][5] ) );
  DFF_X1 \mem_reg[920][4]  ( .D(n18742), .CK(clk), .Q(\mem[920][4] ) );
  DFF_X1 \mem_reg[920][3]  ( .D(n18743), .CK(clk), .Q(\mem[920][3] ) );
  DFF_X1 \mem_reg[920][2]  ( .D(n18744), .CK(clk), .Q(\mem[920][2] ) );
  DFF_X1 \mem_reg[920][1]  ( .D(n18745), .CK(clk), .Q(\mem[920][1] ) );
  DFF_X1 \mem_reg[920][0]  ( .D(n18746), .CK(clk), .Q(\mem[920][0] ) );
  DFF_X1 \mem_reg[919][7]  ( .D(n18747), .CK(clk), .Q(\mem[919][7] ) );
  DFF_X1 \mem_reg[919][6]  ( .D(n18748), .CK(clk), .Q(\mem[919][6] ) );
  DFF_X1 \mem_reg[919][5]  ( .D(n18749), .CK(clk), .Q(\mem[919][5] ) );
  DFF_X1 \mem_reg[919][4]  ( .D(n18750), .CK(clk), .Q(\mem[919][4] ) );
  DFF_X1 \mem_reg[919][3]  ( .D(n18751), .CK(clk), .Q(\mem[919][3] ) );
  DFF_X1 \mem_reg[919][2]  ( .D(n18752), .CK(clk), .Q(\mem[919][2] ) );
  DFF_X1 \mem_reg[919][1]  ( .D(n18753), .CK(clk), .Q(\mem[919][1] ) );
  DFF_X1 \mem_reg[919][0]  ( .D(n18754), .CK(clk), .Q(\mem[919][0] ) );
  DFF_X1 \mem_reg[918][7]  ( .D(n18755), .CK(clk), .Q(\mem[918][7] ) );
  DFF_X1 \mem_reg[918][6]  ( .D(n18756), .CK(clk), .Q(\mem[918][6] ) );
  DFF_X1 \mem_reg[918][5]  ( .D(n18757), .CK(clk), .Q(\mem[918][5] ) );
  DFF_X1 \mem_reg[918][4]  ( .D(n18758), .CK(clk), .Q(\mem[918][4] ) );
  DFF_X1 \mem_reg[918][3]  ( .D(n18759), .CK(clk), .Q(\mem[918][3] ) );
  DFF_X1 \mem_reg[918][2]  ( .D(n18760), .CK(clk), .Q(\mem[918][2] ) );
  DFF_X1 \mem_reg[918][1]  ( .D(n18761), .CK(clk), .Q(\mem[918][1] ) );
  DFF_X1 \mem_reg[918][0]  ( .D(n18762), .CK(clk), .Q(\mem[918][0] ) );
  DFF_X1 \mem_reg[917][7]  ( .D(n18763), .CK(clk), .Q(\mem[917][7] ) );
  DFF_X1 \mem_reg[917][6]  ( .D(n18764), .CK(clk), .Q(\mem[917][6] ) );
  DFF_X1 \mem_reg[917][5]  ( .D(n18765), .CK(clk), .Q(\mem[917][5] ) );
  DFF_X1 \mem_reg[917][4]  ( .D(n18766), .CK(clk), .Q(\mem[917][4] ) );
  DFF_X1 \mem_reg[917][3]  ( .D(n18767), .CK(clk), .Q(\mem[917][3] ) );
  DFF_X1 \mem_reg[917][2]  ( .D(n18768), .CK(clk), .Q(\mem[917][2] ) );
  DFF_X1 \mem_reg[917][1]  ( .D(n18769), .CK(clk), .Q(\mem[917][1] ) );
  DFF_X1 \mem_reg[917][0]  ( .D(n18770), .CK(clk), .Q(\mem[917][0] ) );
  DFF_X1 \mem_reg[916][7]  ( .D(n18771), .CK(clk), .Q(\mem[916][7] ) );
  DFF_X1 \mem_reg[916][6]  ( .D(n18772), .CK(clk), .Q(\mem[916][6] ) );
  DFF_X1 \mem_reg[916][5]  ( .D(n18773), .CK(clk), .Q(\mem[916][5] ) );
  DFF_X1 \mem_reg[916][4]  ( .D(n18774), .CK(clk), .Q(\mem[916][4] ) );
  DFF_X1 \mem_reg[916][3]  ( .D(n18775), .CK(clk), .Q(\mem[916][3] ) );
  DFF_X1 \mem_reg[916][2]  ( .D(n18776), .CK(clk), .Q(\mem[916][2] ) );
  DFF_X1 \mem_reg[916][1]  ( .D(n18777), .CK(clk), .Q(\mem[916][1] ) );
  DFF_X1 \mem_reg[916][0]  ( .D(n18778), .CK(clk), .Q(\mem[916][0] ) );
  DFF_X1 \mem_reg[915][7]  ( .D(n18779), .CK(clk), .Q(\mem[915][7] ) );
  DFF_X1 \mem_reg[915][6]  ( .D(n18780), .CK(clk), .Q(\mem[915][6] ) );
  DFF_X1 \mem_reg[915][5]  ( .D(n18781), .CK(clk), .Q(\mem[915][5] ) );
  DFF_X1 \mem_reg[915][4]  ( .D(n18782), .CK(clk), .Q(\mem[915][4] ) );
  DFF_X1 \mem_reg[915][3]  ( .D(n18783), .CK(clk), .Q(\mem[915][3] ) );
  DFF_X1 \mem_reg[915][2]  ( .D(n18784), .CK(clk), .Q(\mem[915][2] ) );
  DFF_X1 \mem_reg[915][1]  ( .D(n18785), .CK(clk), .Q(\mem[915][1] ) );
  DFF_X1 \mem_reg[915][0]  ( .D(n18786), .CK(clk), .Q(\mem[915][0] ) );
  DFF_X1 \mem_reg[914][7]  ( .D(n18787), .CK(clk), .Q(\mem[914][7] ) );
  DFF_X1 \mem_reg[914][6]  ( .D(n18788), .CK(clk), .Q(\mem[914][6] ) );
  DFF_X1 \mem_reg[914][5]  ( .D(n18789), .CK(clk), .Q(\mem[914][5] ) );
  DFF_X1 \mem_reg[914][4]  ( .D(n18790), .CK(clk), .Q(\mem[914][4] ) );
  DFF_X1 \mem_reg[914][3]  ( .D(n18791), .CK(clk), .Q(\mem[914][3] ) );
  DFF_X1 \mem_reg[914][2]  ( .D(n18792), .CK(clk), .Q(\mem[914][2] ) );
  DFF_X1 \mem_reg[914][1]  ( .D(n18793), .CK(clk), .Q(\mem[914][1] ) );
  DFF_X1 \mem_reg[914][0]  ( .D(n18794), .CK(clk), .Q(\mem[914][0] ) );
  DFF_X1 \mem_reg[913][7]  ( .D(n18795), .CK(clk), .Q(\mem[913][7] ) );
  DFF_X1 \mem_reg[913][6]  ( .D(n18796), .CK(clk), .Q(\mem[913][6] ) );
  DFF_X1 \mem_reg[913][5]  ( .D(n18797), .CK(clk), .Q(\mem[913][5] ) );
  DFF_X1 \mem_reg[913][4]  ( .D(n18798), .CK(clk), .Q(\mem[913][4] ) );
  DFF_X1 \mem_reg[913][3]  ( .D(n18799), .CK(clk), .Q(\mem[913][3] ) );
  DFF_X1 \mem_reg[913][2]  ( .D(n18800), .CK(clk), .Q(\mem[913][2] ) );
  DFF_X1 \mem_reg[913][1]  ( .D(n18801), .CK(clk), .Q(\mem[913][1] ) );
  DFF_X1 \mem_reg[913][0]  ( .D(n18802), .CK(clk), .Q(\mem[913][0] ) );
  DFF_X1 \mem_reg[912][7]  ( .D(n18803), .CK(clk), .Q(\mem[912][7] ) );
  DFF_X1 \mem_reg[912][6]  ( .D(n18804), .CK(clk), .Q(\mem[912][6] ) );
  DFF_X1 \mem_reg[912][5]  ( .D(n18805), .CK(clk), .Q(\mem[912][5] ) );
  DFF_X1 \mem_reg[912][4]  ( .D(n18806), .CK(clk), .Q(\mem[912][4] ) );
  DFF_X1 \mem_reg[912][3]  ( .D(n18807), .CK(clk), .Q(\mem[912][3] ) );
  DFF_X1 \mem_reg[912][2]  ( .D(n18808), .CK(clk), .Q(\mem[912][2] ) );
  DFF_X1 \mem_reg[912][1]  ( .D(n18809), .CK(clk), .Q(\mem[912][1] ) );
  DFF_X1 \mem_reg[912][0]  ( .D(n18810), .CK(clk), .Q(\mem[912][0] ) );
  DFF_X1 \mem_reg[911][7]  ( .D(n18811), .CK(clk), .Q(\mem[911][7] ) );
  DFF_X1 \mem_reg[911][6]  ( .D(n18812), .CK(clk), .Q(\mem[911][6] ) );
  DFF_X1 \mem_reg[911][5]  ( .D(n18813), .CK(clk), .Q(\mem[911][5] ) );
  DFF_X1 \mem_reg[911][4]  ( .D(n18814), .CK(clk), .Q(\mem[911][4] ) );
  DFF_X1 \mem_reg[911][3]  ( .D(n18815), .CK(clk), .Q(\mem[911][3] ) );
  DFF_X1 \mem_reg[911][2]  ( .D(n18816), .CK(clk), .Q(\mem[911][2] ) );
  DFF_X1 \mem_reg[911][1]  ( .D(n18817), .CK(clk), .Q(\mem[911][1] ) );
  DFF_X1 \mem_reg[911][0]  ( .D(n18818), .CK(clk), .Q(\mem[911][0] ) );
  DFF_X1 \mem_reg[910][7]  ( .D(n18819), .CK(clk), .Q(\mem[910][7] ) );
  DFF_X1 \mem_reg[910][6]  ( .D(n18820), .CK(clk), .Q(\mem[910][6] ) );
  DFF_X1 \mem_reg[910][5]  ( .D(n18821), .CK(clk), .Q(\mem[910][5] ) );
  DFF_X1 \mem_reg[910][4]  ( .D(n18822), .CK(clk), .Q(\mem[910][4] ) );
  DFF_X1 \mem_reg[910][3]  ( .D(n18823), .CK(clk), .Q(\mem[910][3] ) );
  DFF_X1 \mem_reg[910][2]  ( .D(n18824), .CK(clk), .Q(\mem[910][2] ) );
  DFF_X1 \mem_reg[910][1]  ( .D(n18825), .CK(clk), .Q(\mem[910][1] ) );
  DFF_X1 \mem_reg[910][0]  ( .D(n18826), .CK(clk), .Q(\mem[910][0] ) );
  DFF_X1 \mem_reg[909][7]  ( .D(n18827), .CK(clk), .Q(\mem[909][7] ) );
  DFF_X1 \mem_reg[909][6]  ( .D(n18828), .CK(clk), .Q(\mem[909][6] ) );
  DFF_X1 \mem_reg[909][5]  ( .D(n18829), .CK(clk), .Q(\mem[909][5] ) );
  DFF_X1 \mem_reg[909][4]  ( .D(n18830), .CK(clk), .Q(\mem[909][4] ) );
  DFF_X1 \mem_reg[909][3]  ( .D(n18831), .CK(clk), .Q(\mem[909][3] ) );
  DFF_X1 \mem_reg[909][2]  ( .D(n18832), .CK(clk), .Q(\mem[909][2] ) );
  DFF_X1 \mem_reg[909][1]  ( .D(n18833), .CK(clk), .Q(\mem[909][1] ) );
  DFF_X1 \mem_reg[909][0]  ( .D(n18834), .CK(clk), .Q(\mem[909][0] ) );
  DFF_X1 \mem_reg[908][7]  ( .D(n18835), .CK(clk), .Q(\mem[908][7] ) );
  DFF_X1 \mem_reg[908][6]  ( .D(n18836), .CK(clk), .Q(\mem[908][6] ) );
  DFF_X1 \mem_reg[908][5]  ( .D(n18837), .CK(clk), .Q(\mem[908][5] ) );
  DFF_X1 \mem_reg[908][4]  ( .D(n18838), .CK(clk), .Q(\mem[908][4] ) );
  DFF_X1 \mem_reg[908][3]  ( .D(n18839), .CK(clk), .Q(\mem[908][3] ) );
  DFF_X1 \mem_reg[908][2]  ( .D(n18840), .CK(clk), .Q(\mem[908][2] ) );
  DFF_X1 \mem_reg[908][1]  ( .D(n18841), .CK(clk), .Q(\mem[908][1] ) );
  DFF_X1 \mem_reg[908][0]  ( .D(n18842), .CK(clk), .Q(\mem[908][0] ) );
  DFF_X1 \mem_reg[907][7]  ( .D(n18843), .CK(clk), .Q(\mem[907][7] ) );
  DFF_X1 \mem_reg[907][6]  ( .D(n18844), .CK(clk), .Q(\mem[907][6] ) );
  DFF_X1 \mem_reg[907][5]  ( .D(n18845), .CK(clk), .Q(\mem[907][5] ) );
  DFF_X1 \mem_reg[907][4]  ( .D(n18846), .CK(clk), .Q(\mem[907][4] ) );
  DFF_X1 \mem_reg[907][3]  ( .D(n18847), .CK(clk), .Q(\mem[907][3] ) );
  DFF_X1 \mem_reg[907][2]  ( .D(n18848), .CK(clk), .Q(\mem[907][2] ) );
  DFF_X1 \mem_reg[907][1]  ( .D(n18849), .CK(clk), .Q(\mem[907][1] ) );
  DFF_X1 \mem_reg[907][0]  ( .D(n18850), .CK(clk), .Q(\mem[907][0] ) );
  DFF_X1 \mem_reg[906][7]  ( .D(n18851), .CK(clk), .Q(\mem[906][7] ) );
  DFF_X1 \mem_reg[906][6]  ( .D(n18852), .CK(clk), .Q(\mem[906][6] ) );
  DFF_X1 \mem_reg[906][5]  ( .D(n18853), .CK(clk), .Q(\mem[906][5] ) );
  DFF_X1 \mem_reg[906][4]  ( .D(n18854), .CK(clk), .Q(\mem[906][4] ) );
  DFF_X1 \mem_reg[906][3]  ( .D(n18855), .CK(clk), .Q(\mem[906][3] ) );
  DFF_X1 \mem_reg[906][2]  ( .D(n18856), .CK(clk), .Q(\mem[906][2] ) );
  DFF_X1 \mem_reg[906][1]  ( .D(n18857), .CK(clk), .Q(\mem[906][1] ) );
  DFF_X1 \mem_reg[906][0]  ( .D(n18858), .CK(clk), .Q(\mem[906][0] ) );
  DFF_X1 \mem_reg[905][7]  ( .D(n18859), .CK(clk), .Q(\mem[905][7] ) );
  DFF_X1 \mem_reg[905][6]  ( .D(n18860), .CK(clk), .Q(\mem[905][6] ) );
  DFF_X1 \mem_reg[905][5]  ( .D(n18861), .CK(clk), .Q(\mem[905][5] ) );
  DFF_X1 \mem_reg[905][4]  ( .D(n18862), .CK(clk), .Q(\mem[905][4] ) );
  DFF_X1 \mem_reg[905][3]  ( .D(n18863), .CK(clk), .Q(\mem[905][3] ) );
  DFF_X1 \mem_reg[905][2]  ( .D(n18864), .CK(clk), .Q(\mem[905][2] ) );
  DFF_X1 \mem_reg[905][1]  ( .D(n18865), .CK(clk), .Q(\mem[905][1] ) );
  DFF_X1 \mem_reg[905][0]  ( .D(n18866), .CK(clk), .Q(\mem[905][0] ) );
  DFF_X1 \mem_reg[904][7]  ( .D(n18867), .CK(clk), .Q(\mem[904][7] ) );
  DFF_X1 \mem_reg[904][6]  ( .D(n18868), .CK(clk), .Q(\mem[904][6] ) );
  DFF_X1 \mem_reg[904][5]  ( .D(n18869), .CK(clk), .Q(\mem[904][5] ) );
  DFF_X1 \mem_reg[904][4]  ( .D(n18870), .CK(clk), .Q(\mem[904][4] ) );
  DFF_X1 \mem_reg[904][3]  ( .D(n18871), .CK(clk), .Q(\mem[904][3] ) );
  DFF_X1 \mem_reg[904][2]  ( .D(n18872), .CK(clk), .Q(\mem[904][2] ) );
  DFF_X1 \mem_reg[904][1]  ( .D(n18873), .CK(clk), .Q(\mem[904][1] ) );
  DFF_X1 \mem_reg[904][0]  ( .D(n18874), .CK(clk), .Q(\mem[904][0] ) );
  DFF_X1 \mem_reg[903][7]  ( .D(n18875), .CK(clk), .Q(\mem[903][7] ) );
  DFF_X1 \mem_reg[903][6]  ( .D(n18876), .CK(clk), .Q(\mem[903][6] ) );
  DFF_X1 \mem_reg[903][5]  ( .D(n18877), .CK(clk), .Q(\mem[903][5] ) );
  DFF_X1 \mem_reg[903][4]  ( .D(n18878), .CK(clk), .Q(\mem[903][4] ) );
  DFF_X1 \mem_reg[903][3]  ( .D(n18879), .CK(clk), .Q(\mem[903][3] ) );
  DFF_X1 \mem_reg[903][2]  ( .D(n18880), .CK(clk), .Q(\mem[903][2] ) );
  DFF_X1 \mem_reg[903][1]  ( .D(n18881), .CK(clk), .Q(\mem[903][1] ) );
  DFF_X1 \mem_reg[903][0]  ( .D(n18882), .CK(clk), .Q(\mem[903][0] ) );
  DFF_X1 \mem_reg[902][7]  ( .D(n18883), .CK(clk), .Q(\mem[902][7] ) );
  DFF_X1 \mem_reg[902][6]  ( .D(n18884), .CK(clk), .Q(\mem[902][6] ) );
  DFF_X1 \mem_reg[902][5]  ( .D(n18885), .CK(clk), .Q(\mem[902][5] ) );
  DFF_X1 \mem_reg[902][4]  ( .D(n18886), .CK(clk), .Q(\mem[902][4] ) );
  DFF_X1 \mem_reg[902][3]  ( .D(n18887), .CK(clk), .Q(\mem[902][3] ) );
  DFF_X1 \mem_reg[902][2]  ( .D(n18888), .CK(clk), .Q(\mem[902][2] ) );
  DFF_X1 \mem_reg[902][1]  ( .D(n18889), .CK(clk), .Q(\mem[902][1] ) );
  DFF_X1 \mem_reg[902][0]  ( .D(n18890), .CK(clk), .Q(\mem[902][0] ) );
  DFF_X1 \mem_reg[901][7]  ( .D(n18891), .CK(clk), .Q(\mem[901][7] ) );
  DFF_X1 \mem_reg[901][6]  ( .D(n18892), .CK(clk), .Q(\mem[901][6] ) );
  DFF_X1 \mem_reg[901][5]  ( .D(n18893), .CK(clk), .Q(\mem[901][5] ) );
  DFF_X1 \mem_reg[901][4]  ( .D(n18894), .CK(clk), .Q(\mem[901][4] ) );
  DFF_X1 \mem_reg[901][3]  ( .D(n18895), .CK(clk), .Q(\mem[901][3] ) );
  DFF_X1 \mem_reg[901][2]  ( .D(n18896), .CK(clk), .Q(\mem[901][2] ) );
  DFF_X1 \mem_reg[901][1]  ( .D(n18897), .CK(clk), .Q(\mem[901][1] ) );
  DFF_X1 \mem_reg[901][0]  ( .D(n18898), .CK(clk), .Q(\mem[901][0] ) );
  DFF_X1 \mem_reg[900][7]  ( .D(n18899), .CK(clk), .Q(\mem[900][7] ) );
  DFF_X1 \mem_reg[900][6]  ( .D(n18900), .CK(clk), .Q(\mem[900][6] ) );
  DFF_X1 \mem_reg[900][5]  ( .D(n18901), .CK(clk), .Q(\mem[900][5] ) );
  DFF_X1 \mem_reg[900][4]  ( .D(n18902), .CK(clk), .Q(\mem[900][4] ) );
  DFF_X1 \mem_reg[900][3]  ( .D(n18903), .CK(clk), .Q(\mem[900][3] ) );
  DFF_X1 \mem_reg[900][2]  ( .D(n18904), .CK(clk), .Q(\mem[900][2] ) );
  DFF_X1 \mem_reg[900][1]  ( .D(n18905), .CK(clk), .Q(\mem[900][1] ) );
  DFF_X1 \mem_reg[900][0]  ( .D(n18906), .CK(clk), .Q(\mem[900][0] ) );
  DFF_X1 \mem_reg[899][7]  ( .D(n18907), .CK(clk), .Q(\mem[899][7] ) );
  DFF_X1 \mem_reg[899][6]  ( .D(n18908), .CK(clk), .Q(\mem[899][6] ) );
  DFF_X1 \mem_reg[899][5]  ( .D(n18909), .CK(clk), .Q(\mem[899][5] ) );
  DFF_X1 \mem_reg[899][4]  ( .D(n18910), .CK(clk), .Q(\mem[899][4] ) );
  DFF_X1 \mem_reg[899][3]  ( .D(n18911), .CK(clk), .Q(\mem[899][3] ) );
  DFF_X1 \mem_reg[899][2]  ( .D(n18912), .CK(clk), .Q(\mem[899][2] ) );
  DFF_X1 \mem_reg[899][1]  ( .D(n18913), .CK(clk), .Q(\mem[899][1] ) );
  DFF_X1 \mem_reg[899][0]  ( .D(n18914), .CK(clk), .Q(\mem[899][0] ) );
  DFF_X1 \mem_reg[898][7]  ( .D(n18915), .CK(clk), .Q(\mem[898][7] ) );
  DFF_X1 \mem_reg[898][6]  ( .D(n18916), .CK(clk), .Q(\mem[898][6] ) );
  DFF_X1 \mem_reg[898][5]  ( .D(n18917), .CK(clk), .Q(\mem[898][5] ) );
  DFF_X1 \mem_reg[898][4]  ( .D(n18918), .CK(clk), .Q(\mem[898][4] ) );
  DFF_X1 \mem_reg[898][3]  ( .D(n18919), .CK(clk), .Q(\mem[898][3] ) );
  DFF_X1 \mem_reg[898][2]  ( .D(n18920), .CK(clk), .Q(\mem[898][2] ) );
  DFF_X1 \mem_reg[898][1]  ( .D(n18921), .CK(clk), .Q(\mem[898][1] ) );
  DFF_X1 \mem_reg[898][0]  ( .D(n18922), .CK(clk), .Q(\mem[898][0] ) );
  DFF_X1 \mem_reg[897][7]  ( .D(n18923), .CK(clk), .Q(\mem[897][7] ) );
  DFF_X1 \mem_reg[897][6]  ( .D(n18924), .CK(clk), .Q(\mem[897][6] ) );
  DFF_X1 \mem_reg[897][5]  ( .D(n18925), .CK(clk), .Q(\mem[897][5] ) );
  DFF_X1 \mem_reg[897][4]  ( .D(n18926), .CK(clk), .Q(\mem[897][4] ) );
  DFF_X1 \mem_reg[897][3]  ( .D(n18927), .CK(clk), .Q(\mem[897][3] ) );
  DFF_X1 \mem_reg[897][2]  ( .D(n18928), .CK(clk), .Q(\mem[897][2] ) );
  DFF_X1 \mem_reg[897][1]  ( .D(n18929), .CK(clk), .Q(\mem[897][1] ) );
  DFF_X1 \mem_reg[897][0]  ( .D(n18930), .CK(clk), .Q(\mem[897][0] ) );
  DFF_X1 \mem_reg[896][7]  ( .D(n18931), .CK(clk), .Q(\mem[896][7] ) );
  DFF_X1 \mem_reg[896][6]  ( .D(n18932), .CK(clk), .Q(\mem[896][6] ) );
  DFF_X1 \mem_reg[896][5]  ( .D(n18933), .CK(clk), .Q(\mem[896][5] ) );
  DFF_X1 \mem_reg[896][4]  ( .D(n18934), .CK(clk), .Q(\mem[896][4] ) );
  DFF_X1 \mem_reg[896][3]  ( .D(n18935), .CK(clk), .Q(\mem[896][3] ) );
  DFF_X1 \mem_reg[896][2]  ( .D(n18936), .CK(clk), .Q(\mem[896][2] ) );
  DFF_X1 \mem_reg[896][1]  ( .D(n18937), .CK(clk), .Q(\mem[896][1] ) );
  DFF_X1 \mem_reg[896][0]  ( .D(n18938), .CK(clk), .Q(\mem[896][0] ) );
  DFF_X1 \mem_reg[895][7]  ( .D(n18939), .CK(clk), .Q(\mem[895][7] ) );
  DFF_X1 \mem_reg[895][6]  ( .D(n18940), .CK(clk), .Q(\mem[895][6] ) );
  DFF_X1 \mem_reg[895][5]  ( .D(n18941), .CK(clk), .Q(\mem[895][5] ) );
  DFF_X1 \mem_reg[895][4]  ( .D(n18942), .CK(clk), .Q(\mem[895][4] ) );
  DFF_X1 \mem_reg[895][3]  ( .D(n18943), .CK(clk), .Q(\mem[895][3] ) );
  DFF_X1 \mem_reg[895][2]  ( .D(n18944), .CK(clk), .Q(\mem[895][2] ) );
  DFF_X1 \mem_reg[895][1]  ( .D(n18945), .CK(clk), .Q(\mem[895][1] ) );
  DFF_X1 \mem_reg[895][0]  ( .D(n18946), .CK(clk), .Q(\mem[895][0] ) );
  DFF_X1 \mem_reg[894][7]  ( .D(n18947), .CK(clk), .Q(\mem[894][7] ) );
  DFF_X1 \mem_reg[894][6]  ( .D(n18948), .CK(clk), .Q(\mem[894][6] ) );
  DFF_X1 \mem_reg[894][5]  ( .D(n18949), .CK(clk), .Q(\mem[894][5] ) );
  DFF_X1 \mem_reg[894][4]  ( .D(n18950), .CK(clk), .Q(\mem[894][4] ) );
  DFF_X1 \mem_reg[894][3]  ( .D(n18951), .CK(clk), .Q(\mem[894][3] ) );
  DFF_X1 \mem_reg[894][2]  ( .D(n18952), .CK(clk), .Q(\mem[894][2] ) );
  DFF_X1 \mem_reg[894][1]  ( .D(n18953), .CK(clk), .Q(\mem[894][1] ) );
  DFF_X1 \mem_reg[894][0]  ( .D(n18954), .CK(clk), .Q(\mem[894][0] ) );
  DFF_X1 \mem_reg[893][7]  ( .D(n18955), .CK(clk), .Q(\mem[893][7] ) );
  DFF_X1 \mem_reg[893][6]  ( .D(n18956), .CK(clk), .Q(\mem[893][6] ) );
  DFF_X1 \mem_reg[893][5]  ( .D(n18957), .CK(clk), .Q(\mem[893][5] ) );
  DFF_X1 \mem_reg[893][4]  ( .D(n18958), .CK(clk), .Q(\mem[893][4] ) );
  DFF_X1 \mem_reg[893][3]  ( .D(n18959), .CK(clk), .Q(\mem[893][3] ) );
  DFF_X1 \mem_reg[893][2]  ( .D(n18960), .CK(clk), .Q(\mem[893][2] ) );
  DFF_X1 \mem_reg[893][1]  ( .D(n18961), .CK(clk), .Q(\mem[893][1] ) );
  DFF_X1 \mem_reg[893][0]  ( .D(n18962), .CK(clk), .Q(\mem[893][0] ) );
  DFF_X1 \mem_reg[892][7]  ( .D(n18963), .CK(clk), .Q(\mem[892][7] ) );
  DFF_X1 \mem_reg[892][6]  ( .D(n18964), .CK(clk), .Q(\mem[892][6] ) );
  DFF_X1 \mem_reg[892][5]  ( .D(n18965), .CK(clk), .Q(\mem[892][5] ) );
  DFF_X1 \mem_reg[892][4]  ( .D(n18966), .CK(clk), .Q(\mem[892][4] ) );
  DFF_X1 \mem_reg[892][3]  ( .D(n18967), .CK(clk), .Q(\mem[892][3] ) );
  DFF_X1 \mem_reg[892][2]  ( .D(n18968), .CK(clk), .Q(\mem[892][2] ) );
  DFF_X1 \mem_reg[892][1]  ( .D(n18969), .CK(clk), .Q(\mem[892][1] ) );
  DFF_X1 \mem_reg[892][0]  ( .D(n18970), .CK(clk), .Q(\mem[892][0] ) );
  DFF_X1 \mem_reg[891][7]  ( .D(n18971), .CK(clk), .Q(\mem[891][7] ) );
  DFF_X1 \mem_reg[891][6]  ( .D(n18972), .CK(clk), .Q(\mem[891][6] ) );
  DFF_X1 \mem_reg[891][5]  ( .D(n18973), .CK(clk), .Q(\mem[891][5] ) );
  DFF_X1 \mem_reg[891][4]  ( .D(n18974), .CK(clk), .Q(\mem[891][4] ) );
  DFF_X1 \mem_reg[891][3]  ( .D(n18975), .CK(clk), .Q(\mem[891][3] ) );
  DFF_X1 \mem_reg[891][2]  ( .D(n18976), .CK(clk), .Q(\mem[891][2] ) );
  DFF_X1 \mem_reg[891][1]  ( .D(n18977), .CK(clk), .Q(\mem[891][1] ) );
  DFF_X1 \mem_reg[891][0]  ( .D(n18978), .CK(clk), .Q(\mem[891][0] ) );
  DFF_X1 \mem_reg[890][7]  ( .D(n18979), .CK(clk), .Q(\mem[890][7] ) );
  DFF_X1 \mem_reg[890][6]  ( .D(n18980), .CK(clk), .Q(\mem[890][6] ) );
  DFF_X1 \mem_reg[890][5]  ( .D(n18981), .CK(clk), .Q(\mem[890][5] ) );
  DFF_X1 \mem_reg[890][4]  ( .D(n18982), .CK(clk), .Q(\mem[890][4] ) );
  DFF_X1 \mem_reg[890][3]  ( .D(n18983), .CK(clk), .Q(\mem[890][3] ) );
  DFF_X1 \mem_reg[890][2]  ( .D(n18984), .CK(clk), .Q(\mem[890][2] ) );
  DFF_X1 \mem_reg[890][1]  ( .D(n18985), .CK(clk), .Q(\mem[890][1] ) );
  DFF_X1 \mem_reg[890][0]  ( .D(n18986), .CK(clk), .Q(\mem[890][0] ) );
  DFF_X1 \mem_reg[889][7]  ( .D(n18987), .CK(clk), .Q(\mem[889][7] ) );
  DFF_X1 \mem_reg[889][6]  ( .D(n18988), .CK(clk), .Q(\mem[889][6] ) );
  DFF_X1 \mem_reg[889][5]  ( .D(n18989), .CK(clk), .Q(\mem[889][5] ) );
  DFF_X1 \mem_reg[889][4]  ( .D(n18990), .CK(clk), .Q(\mem[889][4] ) );
  DFF_X1 \mem_reg[889][3]  ( .D(n18991), .CK(clk), .Q(\mem[889][3] ) );
  DFF_X1 \mem_reg[889][2]  ( .D(n18992), .CK(clk), .Q(\mem[889][2] ) );
  DFF_X1 \mem_reg[889][1]  ( .D(n18993), .CK(clk), .Q(\mem[889][1] ) );
  DFF_X1 \mem_reg[889][0]  ( .D(n18994), .CK(clk), .Q(\mem[889][0] ) );
  DFF_X1 \mem_reg[888][7]  ( .D(n18995), .CK(clk), .Q(\mem[888][7] ) );
  DFF_X1 \mem_reg[888][6]  ( .D(n18996), .CK(clk), .Q(\mem[888][6] ) );
  DFF_X1 \mem_reg[888][5]  ( .D(n18997), .CK(clk), .Q(\mem[888][5] ) );
  DFF_X1 \mem_reg[888][4]  ( .D(n18998), .CK(clk), .Q(\mem[888][4] ) );
  DFF_X1 \mem_reg[888][3]  ( .D(n18999), .CK(clk), .Q(\mem[888][3] ) );
  DFF_X1 \mem_reg[888][2]  ( .D(n19000), .CK(clk), .Q(\mem[888][2] ) );
  DFF_X1 \mem_reg[888][1]  ( .D(n19001), .CK(clk), .Q(\mem[888][1] ) );
  DFF_X1 \mem_reg[888][0]  ( .D(n19002), .CK(clk), .Q(\mem[888][0] ) );
  DFF_X1 \mem_reg[887][7]  ( .D(n19003), .CK(clk), .Q(\mem[887][7] ) );
  DFF_X1 \mem_reg[887][6]  ( .D(n19004), .CK(clk), .Q(\mem[887][6] ) );
  DFF_X1 \mem_reg[887][5]  ( .D(n19005), .CK(clk), .Q(\mem[887][5] ) );
  DFF_X1 \mem_reg[887][4]  ( .D(n19006), .CK(clk), .Q(\mem[887][4] ) );
  DFF_X1 \mem_reg[887][3]  ( .D(n19007), .CK(clk), .Q(\mem[887][3] ) );
  DFF_X1 \mem_reg[887][2]  ( .D(n19008), .CK(clk), .Q(\mem[887][2] ) );
  DFF_X1 \mem_reg[887][1]  ( .D(n19009), .CK(clk), .Q(\mem[887][1] ) );
  DFF_X1 \mem_reg[887][0]  ( .D(n19010), .CK(clk), .Q(\mem[887][0] ) );
  DFF_X1 \mem_reg[886][7]  ( .D(n19011), .CK(clk), .Q(\mem[886][7] ) );
  DFF_X1 \mem_reg[886][6]  ( .D(n19012), .CK(clk), .Q(\mem[886][6] ) );
  DFF_X1 \mem_reg[886][5]  ( .D(n19013), .CK(clk), .Q(\mem[886][5] ) );
  DFF_X1 \mem_reg[886][4]  ( .D(n19014), .CK(clk), .Q(\mem[886][4] ) );
  DFF_X1 \mem_reg[886][3]  ( .D(n19015), .CK(clk), .Q(\mem[886][3] ) );
  DFF_X1 \mem_reg[886][2]  ( .D(n19016), .CK(clk), .Q(\mem[886][2] ) );
  DFF_X1 \mem_reg[886][1]  ( .D(n19017), .CK(clk), .Q(\mem[886][1] ) );
  DFF_X1 \mem_reg[886][0]  ( .D(n19018), .CK(clk), .Q(\mem[886][0] ) );
  DFF_X1 \mem_reg[885][7]  ( .D(n19019), .CK(clk), .Q(\mem[885][7] ) );
  DFF_X1 \mem_reg[885][6]  ( .D(n19020), .CK(clk), .Q(\mem[885][6] ) );
  DFF_X1 \mem_reg[885][5]  ( .D(n19021), .CK(clk), .Q(\mem[885][5] ) );
  DFF_X1 \mem_reg[885][4]  ( .D(n19022), .CK(clk), .Q(\mem[885][4] ) );
  DFF_X1 \mem_reg[885][3]  ( .D(n19023), .CK(clk), .Q(\mem[885][3] ) );
  DFF_X1 \mem_reg[885][2]  ( .D(n19024), .CK(clk), .Q(\mem[885][2] ) );
  DFF_X1 \mem_reg[885][1]  ( .D(n19025), .CK(clk), .Q(\mem[885][1] ) );
  DFF_X1 \mem_reg[885][0]  ( .D(n19026), .CK(clk), .Q(\mem[885][0] ) );
  DFF_X1 \mem_reg[884][7]  ( .D(n19027), .CK(clk), .Q(\mem[884][7] ) );
  DFF_X1 \mem_reg[884][6]  ( .D(n19028), .CK(clk), .Q(\mem[884][6] ) );
  DFF_X1 \mem_reg[884][5]  ( .D(n19029), .CK(clk), .Q(\mem[884][5] ) );
  DFF_X1 \mem_reg[884][4]  ( .D(n19030), .CK(clk), .Q(\mem[884][4] ) );
  DFF_X1 \mem_reg[884][3]  ( .D(n19031), .CK(clk), .Q(\mem[884][3] ) );
  DFF_X1 \mem_reg[884][2]  ( .D(n19032), .CK(clk), .Q(\mem[884][2] ) );
  DFF_X1 \mem_reg[884][1]  ( .D(n19033), .CK(clk), .Q(\mem[884][1] ) );
  DFF_X1 \mem_reg[884][0]  ( .D(n19034), .CK(clk), .Q(\mem[884][0] ) );
  DFF_X1 \mem_reg[883][7]  ( .D(n19035), .CK(clk), .Q(\mem[883][7] ) );
  DFF_X1 \mem_reg[883][6]  ( .D(n19036), .CK(clk), .Q(\mem[883][6] ) );
  DFF_X1 \mem_reg[883][5]  ( .D(n19037), .CK(clk), .Q(\mem[883][5] ) );
  DFF_X1 \mem_reg[883][4]  ( .D(n19038), .CK(clk), .Q(\mem[883][4] ) );
  DFF_X1 \mem_reg[883][3]  ( .D(n19039), .CK(clk), .Q(\mem[883][3] ) );
  DFF_X1 \mem_reg[883][2]  ( .D(n19040), .CK(clk), .Q(\mem[883][2] ) );
  DFF_X1 \mem_reg[883][1]  ( .D(n19041), .CK(clk), .Q(\mem[883][1] ) );
  DFF_X1 \mem_reg[883][0]  ( .D(n19042), .CK(clk), .Q(\mem[883][0] ) );
  DFF_X1 \mem_reg[882][7]  ( .D(n19043), .CK(clk), .Q(\mem[882][7] ) );
  DFF_X1 \mem_reg[882][6]  ( .D(n19044), .CK(clk), .Q(\mem[882][6] ) );
  DFF_X1 \mem_reg[882][5]  ( .D(n19045), .CK(clk), .Q(\mem[882][5] ) );
  DFF_X1 \mem_reg[882][4]  ( .D(n19046), .CK(clk), .Q(\mem[882][4] ) );
  DFF_X1 \mem_reg[882][3]  ( .D(n19047), .CK(clk), .Q(\mem[882][3] ) );
  DFF_X1 \mem_reg[882][2]  ( .D(n19048), .CK(clk), .Q(\mem[882][2] ) );
  DFF_X1 \mem_reg[882][1]  ( .D(n19049), .CK(clk), .Q(\mem[882][1] ) );
  DFF_X1 \mem_reg[882][0]  ( .D(n19050), .CK(clk), .Q(\mem[882][0] ) );
  DFF_X1 \mem_reg[881][7]  ( .D(n19051), .CK(clk), .Q(\mem[881][7] ) );
  DFF_X1 \mem_reg[881][6]  ( .D(n19052), .CK(clk), .Q(\mem[881][6] ) );
  DFF_X1 \mem_reg[881][5]  ( .D(n19053), .CK(clk), .Q(\mem[881][5] ) );
  DFF_X1 \mem_reg[881][4]  ( .D(n19054), .CK(clk), .Q(\mem[881][4] ) );
  DFF_X1 \mem_reg[881][3]  ( .D(n19055), .CK(clk), .Q(\mem[881][3] ) );
  DFF_X1 \mem_reg[881][2]  ( .D(n19056), .CK(clk), .Q(\mem[881][2] ) );
  DFF_X1 \mem_reg[881][1]  ( .D(n19057), .CK(clk), .Q(\mem[881][1] ) );
  DFF_X1 \mem_reg[881][0]  ( .D(n19058), .CK(clk), .Q(\mem[881][0] ) );
  DFF_X1 \mem_reg[880][7]  ( .D(n19059), .CK(clk), .Q(\mem[880][7] ) );
  DFF_X1 \mem_reg[880][6]  ( .D(n19060), .CK(clk), .Q(\mem[880][6] ) );
  DFF_X1 \mem_reg[880][5]  ( .D(n19061), .CK(clk), .Q(\mem[880][5] ) );
  DFF_X1 \mem_reg[880][4]  ( .D(n19062), .CK(clk), .Q(\mem[880][4] ) );
  DFF_X1 \mem_reg[880][3]  ( .D(n19063), .CK(clk), .Q(\mem[880][3] ) );
  DFF_X1 \mem_reg[880][2]  ( .D(n19064), .CK(clk), .Q(\mem[880][2] ) );
  DFF_X1 \mem_reg[880][1]  ( .D(n19065), .CK(clk), .Q(\mem[880][1] ) );
  DFF_X1 \mem_reg[880][0]  ( .D(n19066), .CK(clk), .Q(\mem[880][0] ) );
  DFF_X1 \mem_reg[879][7]  ( .D(n19067), .CK(clk), .Q(\mem[879][7] ) );
  DFF_X1 \mem_reg[879][6]  ( .D(n19068), .CK(clk), .Q(\mem[879][6] ) );
  DFF_X1 \mem_reg[879][5]  ( .D(n19069), .CK(clk), .Q(\mem[879][5] ) );
  DFF_X1 \mem_reg[879][4]  ( .D(n19070), .CK(clk), .Q(\mem[879][4] ) );
  DFF_X1 \mem_reg[879][3]  ( .D(n19071), .CK(clk), .Q(\mem[879][3] ) );
  DFF_X1 \mem_reg[879][2]  ( .D(n19072), .CK(clk), .Q(\mem[879][2] ) );
  DFF_X1 \mem_reg[879][1]  ( .D(n19073), .CK(clk), .Q(\mem[879][1] ) );
  DFF_X1 \mem_reg[879][0]  ( .D(n19074), .CK(clk), .Q(\mem[879][0] ) );
  DFF_X1 \mem_reg[878][7]  ( .D(n19075), .CK(clk), .Q(\mem[878][7] ) );
  DFF_X1 \mem_reg[878][6]  ( .D(n19076), .CK(clk), .Q(\mem[878][6] ) );
  DFF_X1 \mem_reg[878][5]  ( .D(n19077), .CK(clk), .Q(\mem[878][5] ) );
  DFF_X1 \mem_reg[878][4]  ( .D(n19078), .CK(clk), .Q(\mem[878][4] ) );
  DFF_X1 \mem_reg[878][3]  ( .D(n19079), .CK(clk), .Q(\mem[878][3] ) );
  DFF_X1 \mem_reg[878][2]  ( .D(n19080), .CK(clk), .Q(\mem[878][2] ) );
  DFF_X1 \mem_reg[878][1]  ( .D(n19081), .CK(clk), .Q(\mem[878][1] ) );
  DFF_X1 \mem_reg[878][0]  ( .D(n19082), .CK(clk), .Q(\mem[878][0] ) );
  DFF_X1 \mem_reg[877][7]  ( .D(n19083), .CK(clk), .Q(\mem[877][7] ) );
  DFF_X1 \mem_reg[877][6]  ( .D(n19084), .CK(clk), .Q(\mem[877][6] ) );
  DFF_X1 \mem_reg[877][5]  ( .D(n19085), .CK(clk), .Q(\mem[877][5] ) );
  DFF_X1 \mem_reg[877][4]  ( .D(n19086), .CK(clk), .Q(\mem[877][4] ) );
  DFF_X1 \mem_reg[877][3]  ( .D(n19087), .CK(clk), .Q(\mem[877][3] ) );
  DFF_X1 \mem_reg[877][2]  ( .D(n19088), .CK(clk), .Q(\mem[877][2] ) );
  DFF_X1 \mem_reg[877][1]  ( .D(n19089), .CK(clk), .Q(\mem[877][1] ) );
  DFF_X1 \mem_reg[877][0]  ( .D(n19090), .CK(clk), .Q(\mem[877][0] ) );
  DFF_X1 \mem_reg[876][7]  ( .D(n19091), .CK(clk), .Q(\mem[876][7] ) );
  DFF_X1 \mem_reg[876][6]  ( .D(n19092), .CK(clk), .Q(\mem[876][6] ) );
  DFF_X1 \mem_reg[876][5]  ( .D(n19093), .CK(clk), .Q(\mem[876][5] ) );
  DFF_X1 \mem_reg[876][4]  ( .D(n19094), .CK(clk), .Q(\mem[876][4] ) );
  DFF_X1 \mem_reg[876][3]  ( .D(n19095), .CK(clk), .Q(\mem[876][3] ) );
  DFF_X1 \mem_reg[876][2]  ( .D(n19096), .CK(clk), .Q(\mem[876][2] ) );
  DFF_X1 \mem_reg[876][1]  ( .D(n19097), .CK(clk), .Q(\mem[876][1] ) );
  DFF_X1 \mem_reg[876][0]  ( .D(n19098), .CK(clk), .Q(\mem[876][0] ) );
  DFF_X1 \mem_reg[875][7]  ( .D(n19099), .CK(clk), .Q(\mem[875][7] ) );
  DFF_X1 \mem_reg[875][6]  ( .D(n19100), .CK(clk), .Q(\mem[875][6] ) );
  DFF_X1 \mem_reg[875][5]  ( .D(n19101), .CK(clk), .Q(\mem[875][5] ) );
  DFF_X1 \mem_reg[875][4]  ( .D(n19102), .CK(clk), .Q(\mem[875][4] ) );
  DFF_X1 \mem_reg[875][3]  ( .D(n19103), .CK(clk), .Q(\mem[875][3] ) );
  DFF_X1 \mem_reg[875][2]  ( .D(n19104), .CK(clk), .Q(\mem[875][2] ) );
  DFF_X1 \mem_reg[875][1]  ( .D(n19105), .CK(clk), .Q(\mem[875][1] ) );
  DFF_X1 \mem_reg[875][0]  ( .D(n19106), .CK(clk), .Q(\mem[875][0] ) );
  DFF_X1 \mem_reg[874][7]  ( .D(n19107), .CK(clk), .Q(\mem[874][7] ) );
  DFF_X1 \mem_reg[874][6]  ( .D(n19108), .CK(clk), .Q(\mem[874][6] ) );
  DFF_X1 \mem_reg[874][5]  ( .D(n19109), .CK(clk), .Q(\mem[874][5] ) );
  DFF_X1 \mem_reg[874][4]  ( .D(n19110), .CK(clk), .Q(\mem[874][4] ) );
  DFF_X1 \mem_reg[874][3]  ( .D(n19111), .CK(clk), .Q(\mem[874][3] ) );
  DFF_X1 \mem_reg[874][2]  ( .D(n19112), .CK(clk), .Q(\mem[874][2] ) );
  DFF_X1 \mem_reg[874][1]  ( .D(n19113), .CK(clk), .Q(\mem[874][1] ) );
  DFF_X1 \mem_reg[874][0]  ( .D(n19114), .CK(clk), .Q(\mem[874][0] ) );
  DFF_X1 \mem_reg[873][7]  ( .D(n19115), .CK(clk), .Q(\mem[873][7] ) );
  DFF_X1 \mem_reg[873][6]  ( .D(n19116), .CK(clk), .Q(\mem[873][6] ) );
  DFF_X1 \mem_reg[873][5]  ( .D(n19117), .CK(clk), .Q(\mem[873][5] ) );
  DFF_X1 \mem_reg[873][4]  ( .D(n19118), .CK(clk), .Q(\mem[873][4] ) );
  DFF_X1 \mem_reg[873][3]  ( .D(n19119), .CK(clk), .Q(\mem[873][3] ) );
  DFF_X1 \mem_reg[873][2]  ( .D(n19120), .CK(clk), .Q(\mem[873][2] ) );
  DFF_X1 \mem_reg[873][1]  ( .D(n19121), .CK(clk), .Q(\mem[873][1] ) );
  DFF_X1 \mem_reg[873][0]  ( .D(n19122), .CK(clk), .Q(\mem[873][0] ) );
  DFF_X1 \mem_reg[872][7]  ( .D(n19123), .CK(clk), .Q(\mem[872][7] ) );
  DFF_X1 \mem_reg[872][6]  ( .D(n19124), .CK(clk), .Q(\mem[872][6] ) );
  DFF_X1 \mem_reg[872][5]  ( .D(n19125), .CK(clk), .Q(\mem[872][5] ) );
  DFF_X1 \mem_reg[872][4]  ( .D(n19126), .CK(clk), .Q(\mem[872][4] ) );
  DFF_X1 \mem_reg[872][3]  ( .D(n19127), .CK(clk), .Q(\mem[872][3] ) );
  DFF_X1 \mem_reg[872][2]  ( .D(n19128), .CK(clk), .Q(\mem[872][2] ) );
  DFF_X1 \mem_reg[872][1]  ( .D(n19129), .CK(clk), .Q(\mem[872][1] ) );
  DFF_X1 \mem_reg[872][0]  ( .D(n19130), .CK(clk), .Q(\mem[872][0] ) );
  DFF_X1 \mem_reg[871][7]  ( .D(n19131), .CK(clk), .Q(\mem[871][7] ) );
  DFF_X1 \mem_reg[871][6]  ( .D(n19132), .CK(clk), .Q(\mem[871][6] ) );
  DFF_X1 \mem_reg[871][5]  ( .D(n19133), .CK(clk), .Q(\mem[871][5] ) );
  DFF_X1 \mem_reg[871][4]  ( .D(n19134), .CK(clk), .Q(\mem[871][4] ) );
  DFF_X1 \mem_reg[871][3]  ( .D(n19135), .CK(clk), .Q(\mem[871][3] ) );
  DFF_X1 \mem_reg[871][2]  ( .D(n19136), .CK(clk), .Q(\mem[871][2] ) );
  DFF_X1 \mem_reg[871][1]  ( .D(n19137), .CK(clk), .Q(\mem[871][1] ) );
  DFF_X1 \mem_reg[871][0]  ( .D(n19138), .CK(clk), .Q(\mem[871][0] ) );
  DFF_X1 \mem_reg[870][7]  ( .D(n19139), .CK(clk), .Q(\mem[870][7] ) );
  DFF_X1 \mem_reg[870][6]  ( .D(n19140), .CK(clk), .Q(\mem[870][6] ) );
  DFF_X1 \mem_reg[870][5]  ( .D(n19141), .CK(clk), .Q(\mem[870][5] ) );
  DFF_X1 \mem_reg[870][4]  ( .D(n19142), .CK(clk), .Q(\mem[870][4] ) );
  DFF_X1 \mem_reg[870][3]  ( .D(n19143), .CK(clk), .Q(\mem[870][3] ) );
  DFF_X1 \mem_reg[870][2]  ( .D(n19144), .CK(clk), .Q(\mem[870][2] ) );
  DFF_X1 \mem_reg[870][1]  ( .D(n19145), .CK(clk), .Q(\mem[870][1] ) );
  DFF_X1 \mem_reg[870][0]  ( .D(n19146), .CK(clk), .Q(\mem[870][0] ) );
  DFF_X1 \mem_reg[869][7]  ( .D(n19147), .CK(clk), .Q(\mem[869][7] ) );
  DFF_X1 \mem_reg[869][6]  ( .D(n19148), .CK(clk), .Q(\mem[869][6] ) );
  DFF_X1 \mem_reg[869][5]  ( .D(n19149), .CK(clk), .Q(\mem[869][5] ) );
  DFF_X1 \mem_reg[869][4]  ( .D(n19150), .CK(clk), .Q(\mem[869][4] ) );
  DFF_X1 \mem_reg[869][3]  ( .D(n19151), .CK(clk), .Q(\mem[869][3] ) );
  DFF_X1 \mem_reg[869][2]  ( .D(n19152), .CK(clk), .Q(\mem[869][2] ) );
  DFF_X1 \mem_reg[869][1]  ( .D(n19153), .CK(clk), .Q(\mem[869][1] ) );
  DFF_X1 \mem_reg[869][0]  ( .D(n19154), .CK(clk), .Q(\mem[869][0] ) );
  DFF_X1 \mem_reg[868][7]  ( .D(n19155), .CK(clk), .Q(\mem[868][7] ) );
  DFF_X1 \mem_reg[868][6]  ( .D(n19156), .CK(clk), .Q(\mem[868][6] ) );
  DFF_X1 \mem_reg[868][5]  ( .D(n19157), .CK(clk), .Q(\mem[868][5] ) );
  DFF_X1 \mem_reg[868][4]  ( .D(n19158), .CK(clk), .Q(\mem[868][4] ) );
  DFF_X1 \mem_reg[868][3]  ( .D(n19159), .CK(clk), .Q(\mem[868][3] ) );
  DFF_X1 \mem_reg[868][2]  ( .D(n19160), .CK(clk), .Q(\mem[868][2] ) );
  DFF_X1 \mem_reg[868][1]  ( .D(n19161), .CK(clk), .Q(\mem[868][1] ) );
  DFF_X1 \mem_reg[868][0]  ( .D(n19162), .CK(clk), .Q(\mem[868][0] ) );
  DFF_X1 \mem_reg[867][7]  ( .D(n19163), .CK(clk), .Q(\mem[867][7] ) );
  DFF_X1 \mem_reg[867][6]  ( .D(n19164), .CK(clk), .Q(\mem[867][6] ) );
  DFF_X1 \mem_reg[867][5]  ( .D(n19165), .CK(clk), .Q(\mem[867][5] ) );
  DFF_X1 \mem_reg[867][4]  ( .D(n19166), .CK(clk), .Q(\mem[867][4] ) );
  DFF_X1 \mem_reg[867][3]  ( .D(n19167), .CK(clk), .Q(\mem[867][3] ) );
  DFF_X1 \mem_reg[867][2]  ( .D(n19168), .CK(clk), .Q(\mem[867][2] ) );
  DFF_X1 \mem_reg[867][1]  ( .D(n19169), .CK(clk), .Q(\mem[867][1] ) );
  DFF_X1 \mem_reg[867][0]  ( .D(n19170), .CK(clk), .Q(\mem[867][0] ) );
  DFF_X1 \mem_reg[866][7]  ( .D(n19171), .CK(clk), .Q(\mem[866][7] ) );
  DFF_X1 \mem_reg[866][6]  ( .D(n19172), .CK(clk), .Q(\mem[866][6] ) );
  DFF_X1 \mem_reg[866][5]  ( .D(n19173), .CK(clk), .Q(\mem[866][5] ) );
  DFF_X1 \mem_reg[866][4]  ( .D(n19174), .CK(clk), .Q(\mem[866][4] ) );
  DFF_X1 \mem_reg[866][3]  ( .D(n19175), .CK(clk), .Q(\mem[866][3] ) );
  DFF_X1 \mem_reg[866][2]  ( .D(n19176), .CK(clk), .Q(\mem[866][2] ) );
  DFF_X1 \mem_reg[866][1]  ( .D(n19177), .CK(clk), .Q(\mem[866][1] ) );
  DFF_X1 \mem_reg[866][0]  ( .D(n19178), .CK(clk), .Q(\mem[866][0] ) );
  DFF_X1 \mem_reg[865][7]  ( .D(n19179), .CK(clk), .Q(\mem[865][7] ) );
  DFF_X1 \mem_reg[865][6]  ( .D(n19180), .CK(clk), .Q(\mem[865][6] ) );
  DFF_X1 \mem_reg[865][5]  ( .D(n19181), .CK(clk), .Q(\mem[865][5] ) );
  DFF_X1 \mem_reg[865][4]  ( .D(n19182), .CK(clk), .Q(\mem[865][4] ) );
  DFF_X1 \mem_reg[865][3]  ( .D(n19183), .CK(clk), .Q(\mem[865][3] ) );
  DFF_X1 \mem_reg[865][2]  ( .D(n19184), .CK(clk), .Q(\mem[865][2] ) );
  DFF_X1 \mem_reg[865][1]  ( .D(n19185), .CK(clk), .Q(\mem[865][1] ) );
  DFF_X1 \mem_reg[865][0]  ( .D(n19186), .CK(clk), .Q(\mem[865][0] ) );
  DFF_X1 \mem_reg[864][7]  ( .D(n19187), .CK(clk), .Q(\mem[864][7] ) );
  DFF_X1 \mem_reg[864][6]  ( .D(n19188), .CK(clk), .Q(\mem[864][6] ) );
  DFF_X1 \mem_reg[864][5]  ( .D(n19189), .CK(clk), .Q(\mem[864][5] ) );
  DFF_X1 \mem_reg[864][4]  ( .D(n19190), .CK(clk), .Q(\mem[864][4] ) );
  DFF_X1 \mem_reg[864][3]  ( .D(n19191), .CK(clk), .Q(\mem[864][3] ) );
  DFF_X1 \mem_reg[864][2]  ( .D(n19192), .CK(clk), .Q(\mem[864][2] ) );
  DFF_X1 \mem_reg[864][1]  ( .D(n19193), .CK(clk), .Q(\mem[864][1] ) );
  DFF_X1 \mem_reg[864][0]  ( .D(n19194), .CK(clk), .Q(\mem[864][0] ) );
  DFF_X1 \mem_reg[863][7]  ( .D(n19195), .CK(clk), .Q(\mem[863][7] ) );
  DFF_X1 \mem_reg[863][6]  ( .D(n19196), .CK(clk), .Q(\mem[863][6] ) );
  DFF_X1 \mem_reg[863][5]  ( .D(n19197), .CK(clk), .Q(\mem[863][5] ) );
  DFF_X1 \mem_reg[863][4]  ( .D(n19198), .CK(clk), .Q(\mem[863][4] ) );
  DFF_X1 \mem_reg[863][3]  ( .D(n19199), .CK(clk), .Q(\mem[863][3] ) );
  DFF_X1 \mem_reg[863][2]  ( .D(n19200), .CK(clk), .Q(\mem[863][2] ) );
  DFF_X1 \mem_reg[863][1]  ( .D(n19201), .CK(clk), .Q(\mem[863][1] ) );
  DFF_X1 \mem_reg[863][0]  ( .D(n19202), .CK(clk), .Q(\mem[863][0] ) );
  DFF_X1 \mem_reg[862][7]  ( .D(n19203), .CK(clk), .Q(\mem[862][7] ) );
  DFF_X1 \mem_reg[862][6]  ( .D(n19204), .CK(clk), .Q(\mem[862][6] ) );
  DFF_X1 \mem_reg[862][5]  ( .D(n19205), .CK(clk), .Q(\mem[862][5] ) );
  DFF_X1 \mem_reg[862][4]  ( .D(n19206), .CK(clk), .Q(\mem[862][4] ) );
  DFF_X1 \mem_reg[862][3]  ( .D(n19207), .CK(clk), .Q(\mem[862][3] ) );
  DFF_X1 \mem_reg[862][2]  ( .D(n19208), .CK(clk), .Q(\mem[862][2] ) );
  DFF_X1 \mem_reg[862][1]  ( .D(n19209), .CK(clk), .Q(\mem[862][1] ) );
  DFF_X1 \mem_reg[862][0]  ( .D(n19210), .CK(clk), .Q(\mem[862][0] ) );
  DFF_X1 \mem_reg[861][7]  ( .D(n19211), .CK(clk), .Q(\mem[861][7] ) );
  DFF_X1 \mem_reg[861][6]  ( .D(n19212), .CK(clk), .Q(\mem[861][6] ) );
  DFF_X1 \mem_reg[861][5]  ( .D(n19213), .CK(clk), .Q(\mem[861][5] ) );
  DFF_X1 \mem_reg[861][4]  ( .D(n19214), .CK(clk), .Q(\mem[861][4] ) );
  DFF_X1 \mem_reg[861][3]  ( .D(n19215), .CK(clk), .Q(\mem[861][3] ) );
  DFF_X1 \mem_reg[861][2]  ( .D(n19216), .CK(clk), .Q(\mem[861][2] ) );
  DFF_X1 \mem_reg[861][1]  ( .D(n19217), .CK(clk), .Q(\mem[861][1] ) );
  DFF_X1 \mem_reg[861][0]  ( .D(n19218), .CK(clk), .Q(\mem[861][0] ) );
  DFF_X1 \mem_reg[860][7]  ( .D(n19219), .CK(clk), .Q(\mem[860][7] ) );
  DFF_X1 \mem_reg[860][6]  ( .D(n19220), .CK(clk), .Q(\mem[860][6] ) );
  DFF_X1 \mem_reg[860][5]  ( .D(n19221), .CK(clk), .Q(\mem[860][5] ) );
  DFF_X1 \mem_reg[860][4]  ( .D(n19222), .CK(clk), .Q(\mem[860][4] ) );
  DFF_X1 \mem_reg[860][3]  ( .D(n19223), .CK(clk), .Q(\mem[860][3] ) );
  DFF_X1 \mem_reg[860][2]  ( .D(n19224), .CK(clk), .Q(\mem[860][2] ) );
  DFF_X1 \mem_reg[860][1]  ( .D(n19225), .CK(clk), .Q(\mem[860][1] ) );
  DFF_X1 \mem_reg[860][0]  ( .D(n19226), .CK(clk), .Q(\mem[860][0] ) );
  DFF_X1 \mem_reg[859][7]  ( .D(n19227), .CK(clk), .Q(\mem[859][7] ) );
  DFF_X1 \mem_reg[859][6]  ( .D(n19228), .CK(clk), .Q(\mem[859][6] ) );
  DFF_X1 \mem_reg[859][5]  ( .D(n19229), .CK(clk), .Q(\mem[859][5] ) );
  DFF_X1 \mem_reg[859][4]  ( .D(n19230), .CK(clk), .Q(\mem[859][4] ) );
  DFF_X1 \mem_reg[859][3]  ( .D(n19231), .CK(clk), .Q(\mem[859][3] ) );
  DFF_X1 \mem_reg[859][2]  ( .D(n19232), .CK(clk), .Q(\mem[859][2] ) );
  DFF_X1 \mem_reg[859][1]  ( .D(n19233), .CK(clk), .Q(\mem[859][1] ) );
  DFF_X1 \mem_reg[859][0]  ( .D(n19234), .CK(clk), .Q(\mem[859][0] ) );
  DFF_X1 \mem_reg[858][7]  ( .D(n19235), .CK(clk), .Q(\mem[858][7] ) );
  DFF_X1 \mem_reg[858][6]  ( .D(n19236), .CK(clk), .Q(\mem[858][6] ) );
  DFF_X1 \mem_reg[858][5]  ( .D(n19237), .CK(clk), .Q(\mem[858][5] ) );
  DFF_X1 \mem_reg[858][4]  ( .D(n19238), .CK(clk), .Q(\mem[858][4] ) );
  DFF_X1 \mem_reg[858][3]  ( .D(n19239), .CK(clk), .Q(\mem[858][3] ) );
  DFF_X1 \mem_reg[858][2]  ( .D(n19240), .CK(clk), .Q(\mem[858][2] ) );
  DFF_X1 \mem_reg[858][1]  ( .D(n19241), .CK(clk), .Q(\mem[858][1] ) );
  DFF_X1 \mem_reg[858][0]  ( .D(n19242), .CK(clk), .Q(\mem[858][0] ) );
  DFF_X1 \mem_reg[857][7]  ( .D(n19243), .CK(clk), .Q(\mem[857][7] ) );
  DFF_X1 \mem_reg[857][6]  ( .D(n19244), .CK(clk), .Q(\mem[857][6] ) );
  DFF_X1 \mem_reg[857][5]  ( .D(n19245), .CK(clk), .Q(\mem[857][5] ) );
  DFF_X1 \mem_reg[857][4]  ( .D(n19246), .CK(clk), .Q(\mem[857][4] ) );
  DFF_X1 \mem_reg[857][3]  ( .D(n19247), .CK(clk), .Q(\mem[857][3] ) );
  DFF_X1 \mem_reg[857][2]  ( .D(n19248), .CK(clk), .Q(\mem[857][2] ) );
  DFF_X1 \mem_reg[857][1]  ( .D(n19249), .CK(clk), .Q(\mem[857][1] ) );
  DFF_X1 \mem_reg[857][0]  ( .D(n19250), .CK(clk), .Q(\mem[857][0] ) );
  DFF_X1 \mem_reg[856][7]  ( .D(n19251), .CK(clk), .Q(\mem[856][7] ) );
  DFF_X1 \mem_reg[856][6]  ( .D(n19252), .CK(clk), .Q(\mem[856][6] ) );
  DFF_X1 \mem_reg[856][5]  ( .D(n19253), .CK(clk), .Q(\mem[856][5] ) );
  DFF_X1 \mem_reg[856][4]  ( .D(n19254), .CK(clk), .Q(\mem[856][4] ) );
  DFF_X1 \mem_reg[856][3]  ( .D(n19255), .CK(clk), .Q(\mem[856][3] ) );
  DFF_X1 \mem_reg[856][2]  ( .D(n19256), .CK(clk), .Q(\mem[856][2] ) );
  DFF_X1 \mem_reg[856][1]  ( .D(n19257), .CK(clk), .Q(\mem[856][1] ) );
  DFF_X1 \mem_reg[856][0]  ( .D(n19258), .CK(clk), .Q(\mem[856][0] ) );
  DFF_X1 \mem_reg[855][7]  ( .D(n19259), .CK(clk), .Q(\mem[855][7] ) );
  DFF_X1 \mem_reg[855][6]  ( .D(n19260), .CK(clk), .Q(\mem[855][6] ) );
  DFF_X1 \mem_reg[855][5]  ( .D(n19261), .CK(clk), .Q(\mem[855][5] ) );
  DFF_X1 \mem_reg[855][4]  ( .D(n19262), .CK(clk), .Q(\mem[855][4] ) );
  DFF_X1 \mem_reg[855][3]  ( .D(n19263), .CK(clk), .Q(\mem[855][3] ) );
  DFF_X1 \mem_reg[855][2]  ( .D(n19264), .CK(clk), .Q(\mem[855][2] ) );
  DFF_X1 \mem_reg[855][1]  ( .D(n19265), .CK(clk), .Q(\mem[855][1] ) );
  DFF_X1 \mem_reg[855][0]  ( .D(n19266), .CK(clk), .Q(\mem[855][0] ) );
  DFF_X1 \mem_reg[854][7]  ( .D(n19267), .CK(clk), .Q(\mem[854][7] ) );
  DFF_X1 \mem_reg[854][6]  ( .D(n19268), .CK(clk), .Q(\mem[854][6] ) );
  DFF_X1 \mem_reg[854][5]  ( .D(n19269), .CK(clk), .Q(\mem[854][5] ) );
  DFF_X1 \mem_reg[854][4]  ( .D(n19270), .CK(clk), .Q(\mem[854][4] ) );
  DFF_X1 \mem_reg[854][3]  ( .D(n19271), .CK(clk), .Q(\mem[854][3] ) );
  DFF_X1 \mem_reg[854][2]  ( .D(n19272), .CK(clk), .Q(\mem[854][2] ) );
  DFF_X1 \mem_reg[854][1]  ( .D(n19273), .CK(clk), .Q(\mem[854][1] ) );
  DFF_X1 \mem_reg[854][0]  ( .D(n19274), .CK(clk), .Q(\mem[854][0] ) );
  DFF_X1 \mem_reg[853][7]  ( .D(n19275), .CK(clk), .Q(\mem[853][7] ) );
  DFF_X1 \mem_reg[853][6]  ( .D(n19276), .CK(clk), .Q(\mem[853][6] ) );
  DFF_X1 \mem_reg[853][5]  ( .D(n19277), .CK(clk), .Q(\mem[853][5] ) );
  DFF_X1 \mem_reg[853][4]  ( .D(n19278), .CK(clk), .Q(\mem[853][4] ) );
  DFF_X1 \mem_reg[853][3]  ( .D(n19279), .CK(clk), .Q(\mem[853][3] ) );
  DFF_X1 \mem_reg[853][2]  ( .D(n19280), .CK(clk), .Q(\mem[853][2] ) );
  DFF_X1 \mem_reg[853][1]  ( .D(n19281), .CK(clk), .Q(\mem[853][1] ) );
  DFF_X1 \mem_reg[853][0]  ( .D(n19282), .CK(clk), .Q(\mem[853][0] ) );
  DFF_X1 \mem_reg[852][7]  ( .D(n19283), .CK(clk), .Q(\mem[852][7] ) );
  DFF_X1 \mem_reg[852][6]  ( .D(n19284), .CK(clk), .Q(\mem[852][6] ) );
  DFF_X1 \mem_reg[852][5]  ( .D(n19285), .CK(clk), .Q(\mem[852][5] ) );
  DFF_X1 \mem_reg[852][4]  ( .D(n19286), .CK(clk), .Q(\mem[852][4] ) );
  DFF_X1 \mem_reg[852][3]  ( .D(n19287), .CK(clk), .Q(\mem[852][3] ) );
  DFF_X1 \mem_reg[852][2]  ( .D(n19288), .CK(clk), .Q(\mem[852][2] ) );
  DFF_X1 \mem_reg[852][1]  ( .D(n19289), .CK(clk), .Q(\mem[852][1] ) );
  DFF_X1 \mem_reg[852][0]  ( .D(n19290), .CK(clk), .Q(\mem[852][0] ) );
  DFF_X1 \mem_reg[851][7]  ( .D(n19291), .CK(clk), .Q(\mem[851][7] ) );
  DFF_X1 \mem_reg[851][6]  ( .D(n19292), .CK(clk), .Q(\mem[851][6] ) );
  DFF_X1 \mem_reg[851][5]  ( .D(n19293), .CK(clk), .Q(\mem[851][5] ) );
  DFF_X1 \mem_reg[851][4]  ( .D(n19294), .CK(clk), .Q(\mem[851][4] ) );
  DFF_X1 \mem_reg[851][3]  ( .D(n19295), .CK(clk), .Q(\mem[851][3] ) );
  DFF_X1 \mem_reg[851][2]  ( .D(n19296), .CK(clk), .Q(\mem[851][2] ) );
  DFF_X1 \mem_reg[851][1]  ( .D(n19297), .CK(clk), .Q(\mem[851][1] ) );
  DFF_X1 \mem_reg[851][0]  ( .D(n19298), .CK(clk), .Q(\mem[851][0] ) );
  DFF_X1 \mem_reg[850][7]  ( .D(n19299), .CK(clk), .Q(\mem[850][7] ) );
  DFF_X1 \mem_reg[850][6]  ( .D(n19300), .CK(clk), .Q(\mem[850][6] ) );
  DFF_X1 \mem_reg[850][5]  ( .D(n19301), .CK(clk), .Q(\mem[850][5] ) );
  DFF_X1 \mem_reg[850][4]  ( .D(n19302), .CK(clk), .Q(\mem[850][4] ) );
  DFF_X1 \mem_reg[850][3]  ( .D(n19303), .CK(clk), .Q(\mem[850][3] ) );
  DFF_X1 \mem_reg[850][2]  ( .D(n19304), .CK(clk), .Q(\mem[850][2] ) );
  DFF_X1 \mem_reg[850][1]  ( .D(n19305), .CK(clk), .Q(\mem[850][1] ) );
  DFF_X1 \mem_reg[850][0]  ( .D(n19306), .CK(clk), .Q(\mem[850][0] ) );
  DFF_X1 \mem_reg[849][7]  ( .D(n19307), .CK(clk), .Q(\mem[849][7] ) );
  DFF_X1 \mem_reg[849][6]  ( .D(n19308), .CK(clk), .Q(\mem[849][6] ) );
  DFF_X1 \mem_reg[849][5]  ( .D(n19309), .CK(clk), .Q(\mem[849][5] ) );
  DFF_X1 \mem_reg[849][4]  ( .D(n19310), .CK(clk), .Q(\mem[849][4] ) );
  DFF_X1 \mem_reg[849][3]  ( .D(n19311), .CK(clk), .Q(\mem[849][3] ) );
  DFF_X1 \mem_reg[849][2]  ( .D(n19312), .CK(clk), .Q(\mem[849][2] ) );
  DFF_X1 \mem_reg[849][1]  ( .D(n19313), .CK(clk), .Q(\mem[849][1] ) );
  DFF_X1 \mem_reg[849][0]  ( .D(n19314), .CK(clk), .Q(\mem[849][0] ) );
  DFF_X1 \mem_reg[848][7]  ( .D(n19315), .CK(clk), .Q(\mem[848][7] ) );
  DFF_X1 \mem_reg[848][6]  ( .D(n19316), .CK(clk), .Q(\mem[848][6] ) );
  DFF_X1 \mem_reg[848][5]  ( .D(n19317), .CK(clk), .Q(\mem[848][5] ) );
  DFF_X1 \mem_reg[848][4]  ( .D(n19318), .CK(clk), .Q(\mem[848][4] ) );
  DFF_X1 \mem_reg[848][3]  ( .D(n19319), .CK(clk), .Q(\mem[848][3] ) );
  DFF_X1 \mem_reg[848][2]  ( .D(n19320), .CK(clk), .Q(\mem[848][2] ) );
  DFF_X1 \mem_reg[848][1]  ( .D(n19321), .CK(clk), .Q(\mem[848][1] ) );
  DFF_X1 \mem_reg[848][0]  ( .D(n19322), .CK(clk), .Q(\mem[848][0] ) );
  DFF_X1 \mem_reg[847][7]  ( .D(n19323), .CK(clk), .Q(\mem[847][7] ) );
  DFF_X1 \mem_reg[847][6]  ( .D(n19324), .CK(clk), .Q(\mem[847][6] ) );
  DFF_X1 \mem_reg[847][5]  ( .D(n19325), .CK(clk), .Q(\mem[847][5] ) );
  DFF_X1 \mem_reg[847][4]  ( .D(n19326), .CK(clk), .Q(\mem[847][4] ) );
  DFF_X1 \mem_reg[847][3]  ( .D(n19327), .CK(clk), .Q(\mem[847][3] ) );
  DFF_X1 \mem_reg[847][2]  ( .D(n19328), .CK(clk), .Q(\mem[847][2] ) );
  DFF_X1 \mem_reg[847][1]  ( .D(n19329), .CK(clk), .Q(\mem[847][1] ) );
  DFF_X1 \mem_reg[847][0]  ( .D(n19330), .CK(clk), .Q(\mem[847][0] ) );
  DFF_X1 \mem_reg[846][7]  ( .D(n19331), .CK(clk), .Q(\mem[846][7] ) );
  DFF_X1 \mem_reg[846][6]  ( .D(n19332), .CK(clk), .Q(\mem[846][6] ) );
  DFF_X1 \mem_reg[846][5]  ( .D(n19333), .CK(clk), .Q(\mem[846][5] ) );
  DFF_X1 \mem_reg[846][4]  ( .D(n19334), .CK(clk), .Q(\mem[846][4] ) );
  DFF_X1 \mem_reg[846][3]  ( .D(n19335), .CK(clk), .Q(\mem[846][3] ) );
  DFF_X1 \mem_reg[846][2]  ( .D(n19336), .CK(clk), .Q(\mem[846][2] ) );
  DFF_X1 \mem_reg[846][1]  ( .D(n19337), .CK(clk), .Q(\mem[846][1] ) );
  DFF_X1 \mem_reg[846][0]  ( .D(n19338), .CK(clk), .Q(\mem[846][0] ) );
  DFF_X1 \mem_reg[845][7]  ( .D(n19339), .CK(clk), .Q(\mem[845][7] ) );
  DFF_X1 \mem_reg[845][6]  ( .D(n19340), .CK(clk), .Q(\mem[845][6] ) );
  DFF_X1 \mem_reg[845][5]  ( .D(n19341), .CK(clk), .Q(\mem[845][5] ) );
  DFF_X1 \mem_reg[845][4]  ( .D(n19342), .CK(clk), .Q(\mem[845][4] ) );
  DFF_X1 \mem_reg[845][3]  ( .D(n19343), .CK(clk), .Q(\mem[845][3] ) );
  DFF_X1 \mem_reg[845][2]  ( .D(n19344), .CK(clk), .Q(\mem[845][2] ) );
  DFF_X1 \mem_reg[845][1]  ( .D(n19345), .CK(clk), .Q(\mem[845][1] ) );
  DFF_X1 \mem_reg[845][0]  ( .D(n19346), .CK(clk), .Q(\mem[845][0] ) );
  DFF_X1 \mem_reg[844][7]  ( .D(n19347), .CK(clk), .Q(\mem[844][7] ) );
  DFF_X1 \mem_reg[844][6]  ( .D(n19348), .CK(clk), .Q(\mem[844][6] ) );
  DFF_X1 \mem_reg[844][5]  ( .D(n19349), .CK(clk), .Q(\mem[844][5] ) );
  DFF_X1 \mem_reg[844][4]  ( .D(n19350), .CK(clk), .Q(\mem[844][4] ) );
  DFF_X1 \mem_reg[844][3]  ( .D(n19351), .CK(clk), .Q(\mem[844][3] ) );
  DFF_X1 \mem_reg[844][2]  ( .D(n19352), .CK(clk), .Q(\mem[844][2] ) );
  DFF_X1 \mem_reg[844][1]  ( .D(n19353), .CK(clk), .Q(\mem[844][1] ) );
  DFF_X1 \mem_reg[844][0]  ( .D(n19354), .CK(clk), .Q(\mem[844][0] ) );
  DFF_X1 \mem_reg[843][7]  ( .D(n19355), .CK(clk), .Q(\mem[843][7] ) );
  DFF_X1 \mem_reg[843][6]  ( .D(n19356), .CK(clk), .Q(\mem[843][6] ) );
  DFF_X1 \mem_reg[843][5]  ( .D(n19357), .CK(clk), .Q(\mem[843][5] ) );
  DFF_X1 \mem_reg[843][4]  ( .D(n19358), .CK(clk), .Q(\mem[843][4] ) );
  DFF_X1 \mem_reg[843][3]  ( .D(n19359), .CK(clk), .Q(\mem[843][3] ) );
  DFF_X1 \mem_reg[843][2]  ( .D(n19360), .CK(clk), .Q(\mem[843][2] ) );
  DFF_X1 \mem_reg[843][1]  ( .D(n19361), .CK(clk), .Q(\mem[843][1] ) );
  DFF_X1 \mem_reg[843][0]  ( .D(n19362), .CK(clk), .Q(\mem[843][0] ) );
  DFF_X1 \mem_reg[842][7]  ( .D(n19363), .CK(clk), .Q(\mem[842][7] ) );
  DFF_X1 \mem_reg[842][6]  ( .D(n19364), .CK(clk), .Q(\mem[842][6] ) );
  DFF_X1 \mem_reg[842][5]  ( .D(n19365), .CK(clk), .Q(\mem[842][5] ) );
  DFF_X1 \mem_reg[842][4]  ( .D(n19366), .CK(clk), .Q(\mem[842][4] ) );
  DFF_X1 \mem_reg[842][3]  ( .D(n19367), .CK(clk), .Q(\mem[842][3] ) );
  DFF_X1 \mem_reg[842][2]  ( .D(n19368), .CK(clk), .Q(\mem[842][2] ) );
  DFF_X1 \mem_reg[842][1]  ( .D(n19369), .CK(clk), .Q(\mem[842][1] ) );
  DFF_X1 \mem_reg[842][0]  ( .D(n19370), .CK(clk), .Q(\mem[842][0] ) );
  DFF_X1 \mem_reg[841][7]  ( .D(n19371), .CK(clk), .Q(\mem[841][7] ) );
  DFF_X1 \mem_reg[841][6]  ( .D(n19372), .CK(clk), .Q(\mem[841][6] ) );
  DFF_X1 \mem_reg[841][5]  ( .D(n19373), .CK(clk), .Q(\mem[841][5] ) );
  DFF_X1 \mem_reg[841][4]  ( .D(n19374), .CK(clk), .Q(\mem[841][4] ) );
  DFF_X1 \mem_reg[841][3]  ( .D(n19375), .CK(clk), .Q(\mem[841][3] ) );
  DFF_X1 \mem_reg[841][2]  ( .D(n19376), .CK(clk), .Q(\mem[841][2] ) );
  DFF_X1 \mem_reg[841][1]  ( .D(n19377), .CK(clk), .Q(\mem[841][1] ) );
  DFF_X1 \mem_reg[841][0]  ( .D(n19378), .CK(clk), .Q(\mem[841][0] ) );
  DFF_X1 \mem_reg[840][7]  ( .D(n19379), .CK(clk), .Q(\mem[840][7] ) );
  DFF_X1 \mem_reg[840][6]  ( .D(n19380), .CK(clk), .Q(\mem[840][6] ) );
  DFF_X1 \mem_reg[840][5]  ( .D(n19381), .CK(clk), .Q(\mem[840][5] ) );
  DFF_X1 \mem_reg[840][4]  ( .D(n19382), .CK(clk), .Q(\mem[840][4] ) );
  DFF_X1 \mem_reg[840][3]  ( .D(n19383), .CK(clk), .Q(\mem[840][3] ) );
  DFF_X1 \mem_reg[840][2]  ( .D(n19384), .CK(clk), .Q(\mem[840][2] ) );
  DFF_X1 \mem_reg[840][1]  ( .D(n19385), .CK(clk), .Q(\mem[840][1] ) );
  DFF_X1 \mem_reg[840][0]  ( .D(n19386), .CK(clk), .Q(\mem[840][0] ) );
  DFF_X1 \mem_reg[839][7]  ( .D(n19387), .CK(clk), .Q(\mem[839][7] ) );
  DFF_X1 \mem_reg[839][6]  ( .D(n19388), .CK(clk), .Q(\mem[839][6] ) );
  DFF_X1 \mem_reg[839][5]  ( .D(n19389), .CK(clk), .Q(\mem[839][5] ) );
  DFF_X1 \mem_reg[839][4]  ( .D(n19390), .CK(clk), .Q(\mem[839][4] ) );
  DFF_X1 \mem_reg[839][3]  ( .D(n19391), .CK(clk), .Q(\mem[839][3] ) );
  DFF_X1 \mem_reg[839][2]  ( .D(n19392), .CK(clk), .Q(\mem[839][2] ) );
  DFF_X1 \mem_reg[839][1]  ( .D(n19393), .CK(clk), .Q(\mem[839][1] ) );
  DFF_X1 \mem_reg[839][0]  ( .D(n19394), .CK(clk), .Q(\mem[839][0] ) );
  DFF_X1 \mem_reg[838][7]  ( .D(n19395), .CK(clk), .Q(\mem[838][7] ) );
  DFF_X1 \mem_reg[838][6]  ( .D(n19396), .CK(clk), .Q(\mem[838][6] ) );
  DFF_X1 \mem_reg[838][5]  ( .D(n19397), .CK(clk), .Q(\mem[838][5] ) );
  DFF_X1 \mem_reg[838][4]  ( .D(n19398), .CK(clk), .Q(\mem[838][4] ) );
  DFF_X1 \mem_reg[838][3]  ( .D(n19399), .CK(clk), .Q(\mem[838][3] ) );
  DFF_X1 \mem_reg[838][2]  ( .D(n19400), .CK(clk), .Q(\mem[838][2] ) );
  DFF_X1 \mem_reg[838][1]  ( .D(n19401), .CK(clk), .Q(\mem[838][1] ) );
  DFF_X1 \mem_reg[838][0]  ( .D(n19402), .CK(clk), .Q(\mem[838][0] ) );
  DFF_X1 \mem_reg[837][7]  ( .D(n19403), .CK(clk), .Q(\mem[837][7] ) );
  DFF_X1 \mem_reg[837][6]  ( .D(n19404), .CK(clk), .Q(\mem[837][6] ) );
  DFF_X1 \mem_reg[837][5]  ( .D(n19405), .CK(clk), .Q(\mem[837][5] ) );
  DFF_X1 \mem_reg[837][4]  ( .D(n19406), .CK(clk), .Q(\mem[837][4] ) );
  DFF_X1 \mem_reg[837][3]  ( .D(n19407), .CK(clk), .Q(\mem[837][3] ) );
  DFF_X1 \mem_reg[837][2]  ( .D(n19408), .CK(clk), .Q(\mem[837][2] ) );
  DFF_X1 \mem_reg[837][1]  ( .D(n19409), .CK(clk), .Q(\mem[837][1] ) );
  DFF_X1 \mem_reg[837][0]  ( .D(n19410), .CK(clk), .Q(\mem[837][0] ) );
  DFF_X1 \mem_reg[836][7]  ( .D(n19411), .CK(clk), .Q(\mem[836][7] ) );
  DFF_X1 \mem_reg[836][6]  ( .D(n19412), .CK(clk), .Q(\mem[836][6] ) );
  DFF_X1 \mem_reg[836][5]  ( .D(n19413), .CK(clk), .Q(\mem[836][5] ) );
  DFF_X1 \mem_reg[836][4]  ( .D(n19414), .CK(clk), .Q(\mem[836][4] ) );
  DFF_X1 \mem_reg[836][3]  ( .D(n19415), .CK(clk), .Q(\mem[836][3] ) );
  DFF_X1 \mem_reg[836][2]  ( .D(n19416), .CK(clk), .Q(\mem[836][2] ) );
  DFF_X1 \mem_reg[836][1]  ( .D(n19417), .CK(clk), .Q(\mem[836][1] ) );
  DFF_X1 \mem_reg[836][0]  ( .D(n19418), .CK(clk), .Q(\mem[836][0] ) );
  DFF_X1 \mem_reg[835][7]  ( .D(n19419), .CK(clk), .Q(\mem[835][7] ) );
  DFF_X1 \mem_reg[835][6]  ( .D(n19420), .CK(clk), .Q(\mem[835][6] ) );
  DFF_X1 \mem_reg[835][5]  ( .D(n19421), .CK(clk), .Q(\mem[835][5] ) );
  DFF_X1 \mem_reg[835][4]  ( .D(n19422), .CK(clk), .Q(\mem[835][4] ) );
  DFF_X1 \mem_reg[835][3]  ( .D(n19423), .CK(clk), .Q(\mem[835][3] ) );
  DFF_X1 \mem_reg[835][2]  ( .D(n19424), .CK(clk), .Q(\mem[835][2] ) );
  DFF_X1 \mem_reg[835][1]  ( .D(n19425), .CK(clk), .Q(\mem[835][1] ) );
  DFF_X1 \mem_reg[835][0]  ( .D(n19426), .CK(clk), .Q(\mem[835][0] ) );
  DFF_X1 \mem_reg[834][7]  ( .D(n19427), .CK(clk), .Q(\mem[834][7] ) );
  DFF_X1 \mem_reg[834][6]  ( .D(n19428), .CK(clk), .Q(\mem[834][6] ) );
  DFF_X1 \mem_reg[834][5]  ( .D(n19429), .CK(clk), .Q(\mem[834][5] ) );
  DFF_X1 \mem_reg[834][4]  ( .D(n19430), .CK(clk), .Q(\mem[834][4] ) );
  DFF_X1 \mem_reg[834][3]  ( .D(n19431), .CK(clk), .Q(\mem[834][3] ) );
  DFF_X1 \mem_reg[834][2]  ( .D(n19432), .CK(clk), .Q(\mem[834][2] ) );
  DFF_X1 \mem_reg[834][1]  ( .D(n19433), .CK(clk), .Q(\mem[834][1] ) );
  DFF_X1 \mem_reg[834][0]  ( .D(n19434), .CK(clk), .Q(\mem[834][0] ) );
  DFF_X1 \mem_reg[833][7]  ( .D(n19435), .CK(clk), .Q(\mem[833][7] ) );
  DFF_X1 \mem_reg[833][6]  ( .D(n19436), .CK(clk), .Q(\mem[833][6] ) );
  DFF_X1 \mem_reg[833][5]  ( .D(n19437), .CK(clk), .Q(\mem[833][5] ) );
  DFF_X1 \mem_reg[833][4]  ( .D(n19438), .CK(clk), .Q(\mem[833][4] ) );
  DFF_X1 \mem_reg[833][3]  ( .D(n19439), .CK(clk), .Q(\mem[833][3] ) );
  DFF_X1 \mem_reg[833][2]  ( .D(n19440), .CK(clk), .Q(\mem[833][2] ) );
  DFF_X1 \mem_reg[833][1]  ( .D(n19441), .CK(clk), .Q(\mem[833][1] ) );
  DFF_X1 \mem_reg[833][0]  ( .D(n19442), .CK(clk), .Q(\mem[833][0] ) );
  DFF_X1 \mem_reg[832][7]  ( .D(n19443), .CK(clk), .Q(\mem[832][7] ) );
  DFF_X1 \mem_reg[832][6]  ( .D(n19444), .CK(clk), .Q(\mem[832][6] ) );
  DFF_X1 \mem_reg[832][5]  ( .D(n19445), .CK(clk), .Q(\mem[832][5] ) );
  DFF_X1 \mem_reg[832][4]  ( .D(n19446), .CK(clk), .Q(\mem[832][4] ) );
  DFF_X1 \mem_reg[832][3]  ( .D(n19447), .CK(clk), .Q(\mem[832][3] ) );
  DFF_X1 \mem_reg[832][2]  ( .D(n19448), .CK(clk), .Q(\mem[832][2] ) );
  DFF_X1 \mem_reg[832][1]  ( .D(n19449), .CK(clk), .Q(\mem[832][1] ) );
  DFF_X1 \mem_reg[832][0]  ( .D(n19450), .CK(clk), .Q(\mem[832][0] ) );
  DFF_X1 \mem_reg[831][7]  ( .D(n19451), .CK(clk), .Q(\mem[831][7] ) );
  DFF_X1 \mem_reg[831][6]  ( .D(n19452), .CK(clk), .Q(\mem[831][6] ) );
  DFF_X1 \mem_reg[831][5]  ( .D(n19453), .CK(clk), .Q(\mem[831][5] ) );
  DFF_X1 \mem_reg[831][4]  ( .D(n19454), .CK(clk), .Q(\mem[831][4] ) );
  DFF_X1 \mem_reg[831][3]  ( .D(n19455), .CK(clk), .Q(\mem[831][3] ) );
  DFF_X1 \mem_reg[831][2]  ( .D(n19456), .CK(clk), .Q(\mem[831][2] ) );
  DFF_X1 \mem_reg[831][1]  ( .D(n19457), .CK(clk), .Q(\mem[831][1] ) );
  DFF_X1 \mem_reg[831][0]  ( .D(n19458), .CK(clk), .Q(\mem[831][0] ) );
  DFF_X1 \mem_reg[830][7]  ( .D(n19459), .CK(clk), .Q(\mem[830][7] ) );
  DFF_X1 \mem_reg[830][6]  ( .D(n19460), .CK(clk), .Q(\mem[830][6] ) );
  DFF_X1 \mem_reg[830][5]  ( .D(n19461), .CK(clk), .Q(\mem[830][5] ) );
  DFF_X1 \mem_reg[830][4]  ( .D(n19462), .CK(clk), .Q(\mem[830][4] ) );
  DFF_X1 \mem_reg[830][3]  ( .D(n19463), .CK(clk), .Q(\mem[830][3] ) );
  DFF_X1 \mem_reg[830][2]  ( .D(n19464), .CK(clk), .Q(\mem[830][2] ) );
  DFF_X1 \mem_reg[830][1]  ( .D(n19465), .CK(clk), .Q(\mem[830][1] ) );
  DFF_X1 \mem_reg[830][0]  ( .D(n19466), .CK(clk), .Q(\mem[830][0] ) );
  DFF_X1 \mem_reg[829][7]  ( .D(n19467), .CK(clk), .Q(\mem[829][7] ) );
  DFF_X1 \mem_reg[829][6]  ( .D(n19468), .CK(clk), .Q(\mem[829][6] ) );
  DFF_X1 \mem_reg[829][5]  ( .D(n19469), .CK(clk), .Q(\mem[829][5] ) );
  DFF_X1 \mem_reg[829][4]  ( .D(n19470), .CK(clk), .Q(\mem[829][4] ) );
  DFF_X1 \mem_reg[829][3]  ( .D(n19471), .CK(clk), .Q(\mem[829][3] ) );
  DFF_X1 \mem_reg[829][2]  ( .D(n19472), .CK(clk), .Q(\mem[829][2] ) );
  DFF_X1 \mem_reg[829][1]  ( .D(n19473), .CK(clk), .Q(\mem[829][1] ) );
  DFF_X1 \mem_reg[829][0]  ( .D(n19474), .CK(clk), .Q(\mem[829][0] ) );
  DFF_X1 \mem_reg[828][7]  ( .D(n19475), .CK(clk), .Q(\mem[828][7] ) );
  DFF_X1 \mem_reg[828][6]  ( .D(n19476), .CK(clk), .Q(\mem[828][6] ) );
  DFF_X1 \mem_reg[828][5]  ( .D(n19477), .CK(clk), .Q(\mem[828][5] ) );
  DFF_X1 \mem_reg[828][4]  ( .D(n19478), .CK(clk), .Q(\mem[828][4] ) );
  DFF_X1 \mem_reg[828][3]  ( .D(n19479), .CK(clk), .Q(\mem[828][3] ) );
  DFF_X1 \mem_reg[828][2]  ( .D(n19480), .CK(clk), .Q(\mem[828][2] ) );
  DFF_X1 \mem_reg[828][1]  ( .D(n19481), .CK(clk), .Q(\mem[828][1] ) );
  DFF_X1 \mem_reg[828][0]  ( .D(n19482), .CK(clk), .Q(\mem[828][0] ) );
  DFF_X1 \mem_reg[827][7]  ( .D(n19483), .CK(clk), .Q(\mem[827][7] ) );
  DFF_X1 \mem_reg[827][6]  ( .D(n19484), .CK(clk), .Q(\mem[827][6] ) );
  DFF_X1 \mem_reg[827][5]  ( .D(n19485), .CK(clk), .Q(\mem[827][5] ) );
  DFF_X1 \mem_reg[827][4]  ( .D(n19486), .CK(clk), .Q(\mem[827][4] ) );
  DFF_X1 \mem_reg[827][3]  ( .D(n19487), .CK(clk), .Q(\mem[827][3] ) );
  DFF_X1 \mem_reg[827][2]  ( .D(n19488), .CK(clk), .Q(\mem[827][2] ) );
  DFF_X1 \mem_reg[827][1]  ( .D(n19489), .CK(clk), .Q(\mem[827][1] ) );
  DFF_X1 \mem_reg[827][0]  ( .D(n19490), .CK(clk), .Q(\mem[827][0] ) );
  DFF_X1 \mem_reg[826][7]  ( .D(n19491), .CK(clk), .Q(\mem[826][7] ) );
  DFF_X1 \mem_reg[826][6]  ( .D(n19492), .CK(clk), .Q(\mem[826][6] ) );
  DFF_X1 \mem_reg[826][5]  ( .D(n19493), .CK(clk), .Q(\mem[826][5] ) );
  DFF_X1 \mem_reg[826][4]  ( .D(n19494), .CK(clk), .Q(\mem[826][4] ) );
  DFF_X1 \mem_reg[826][3]  ( .D(n19495), .CK(clk), .Q(\mem[826][3] ) );
  DFF_X1 \mem_reg[826][2]  ( .D(n19496), .CK(clk), .Q(\mem[826][2] ) );
  DFF_X1 \mem_reg[826][1]  ( .D(n19497), .CK(clk), .Q(\mem[826][1] ) );
  DFF_X1 \mem_reg[826][0]  ( .D(n19498), .CK(clk), .Q(\mem[826][0] ) );
  DFF_X1 \mem_reg[825][7]  ( .D(n19499), .CK(clk), .Q(\mem[825][7] ) );
  DFF_X1 \mem_reg[825][6]  ( .D(n19500), .CK(clk), .Q(\mem[825][6] ) );
  DFF_X1 \mem_reg[825][5]  ( .D(n19501), .CK(clk), .Q(\mem[825][5] ) );
  DFF_X1 \mem_reg[825][4]  ( .D(n19502), .CK(clk), .Q(\mem[825][4] ) );
  DFF_X1 \mem_reg[825][3]  ( .D(n19503), .CK(clk), .Q(\mem[825][3] ) );
  DFF_X1 \mem_reg[825][2]  ( .D(n19504), .CK(clk), .Q(\mem[825][2] ) );
  DFF_X1 \mem_reg[825][1]  ( .D(n19505), .CK(clk), .Q(\mem[825][1] ) );
  DFF_X1 \mem_reg[825][0]  ( .D(n19506), .CK(clk), .Q(\mem[825][0] ) );
  DFF_X1 \mem_reg[824][7]  ( .D(n19507), .CK(clk), .Q(\mem[824][7] ) );
  DFF_X1 \mem_reg[824][6]  ( .D(n19508), .CK(clk), .Q(\mem[824][6] ) );
  DFF_X1 \mem_reg[824][5]  ( .D(n19509), .CK(clk), .Q(\mem[824][5] ) );
  DFF_X1 \mem_reg[824][4]  ( .D(n19510), .CK(clk), .Q(\mem[824][4] ) );
  DFF_X1 \mem_reg[824][3]  ( .D(n19511), .CK(clk), .Q(\mem[824][3] ) );
  DFF_X1 \mem_reg[824][2]  ( .D(n19512), .CK(clk), .Q(\mem[824][2] ) );
  DFF_X1 \mem_reg[824][1]  ( .D(n19513), .CK(clk), .Q(\mem[824][1] ) );
  DFF_X1 \mem_reg[824][0]  ( .D(n19514), .CK(clk), .Q(\mem[824][0] ) );
  DFF_X1 \mem_reg[823][7]  ( .D(n19515), .CK(clk), .Q(\mem[823][7] ) );
  DFF_X1 \mem_reg[823][6]  ( .D(n19516), .CK(clk), .Q(\mem[823][6] ) );
  DFF_X1 \mem_reg[823][5]  ( .D(n19517), .CK(clk), .Q(\mem[823][5] ) );
  DFF_X1 \mem_reg[823][4]  ( .D(n19518), .CK(clk), .Q(\mem[823][4] ) );
  DFF_X1 \mem_reg[823][3]  ( .D(n19519), .CK(clk), .Q(\mem[823][3] ) );
  DFF_X1 \mem_reg[823][2]  ( .D(n19520), .CK(clk), .Q(\mem[823][2] ) );
  DFF_X1 \mem_reg[823][1]  ( .D(n19521), .CK(clk), .Q(\mem[823][1] ) );
  DFF_X1 \mem_reg[823][0]  ( .D(n19522), .CK(clk), .Q(\mem[823][0] ) );
  DFF_X1 \mem_reg[822][7]  ( .D(n19523), .CK(clk), .Q(\mem[822][7] ) );
  DFF_X1 \mem_reg[822][6]  ( .D(n19524), .CK(clk), .Q(\mem[822][6] ) );
  DFF_X1 \mem_reg[822][5]  ( .D(n19525), .CK(clk), .Q(\mem[822][5] ) );
  DFF_X1 \mem_reg[822][4]  ( .D(n19526), .CK(clk), .Q(\mem[822][4] ) );
  DFF_X1 \mem_reg[822][3]  ( .D(n19527), .CK(clk), .Q(\mem[822][3] ) );
  DFF_X1 \mem_reg[822][2]  ( .D(n19528), .CK(clk), .Q(\mem[822][2] ) );
  DFF_X1 \mem_reg[822][1]  ( .D(n19529), .CK(clk), .Q(\mem[822][1] ) );
  DFF_X1 \mem_reg[822][0]  ( .D(n19530), .CK(clk), .Q(\mem[822][0] ) );
  DFF_X1 \mem_reg[821][7]  ( .D(n19531), .CK(clk), .Q(\mem[821][7] ) );
  DFF_X1 \mem_reg[821][6]  ( .D(n19532), .CK(clk), .Q(\mem[821][6] ) );
  DFF_X1 \mem_reg[821][5]  ( .D(n19533), .CK(clk), .Q(\mem[821][5] ) );
  DFF_X1 \mem_reg[821][4]  ( .D(n19534), .CK(clk), .Q(\mem[821][4] ) );
  DFF_X1 \mem_reg[821][3]  ( .D(n19535), .CK(clk), .Q(\mem[821][3] ) );
  DFF_X1 \mem_reg[821][2]  ( .D(n19536), .CK(clk), .Q(\mem[821][2] ) );
  DFF_X1 \mem_reg[821][1]  ( .D(n19537), .CK(clk), .Q(\mem[821][1] ) );
  DFF_X1 \mem_reg[821][0]  ( .D(n19538), .CK(clk), .Q(\mem[821][0] ) );
  DFF_X1 \mem_reg[820][7]  ( .D(n19539), .CK(clk), .Q(\mem[820][7] ) );
  DFF_X1 \mem_reg[820][6]  ( .D(n19540), .CK(clk), .Q(\mem[820][6] ) );
  DFF_X1 \mem_reg[820][5]  ( .D(n19541), .CK(clk), .Q(\mem[820][5] ) );
  DFF_X1 \mem_reg[820][4]  ( .D(n19542), .CK(clk), .Q(\mem[820][4] ) );
  DFF_X1 \mem_reg[820][3]  ( .D(n19543), .CK(clk), .Q(\mem[820][3] ) );
  DFF_X1 \mem_reg[820][2]  ( .D(n19544), .CK(clk), .Q(\mem[820][2] ) );
  DFF_X1 \mem_reg[820][1]  ( .D(n19545), .CK(clk), .Q(\mem[820][1] ) );
  DFF_X1 \mem_reg[820][0]  ( .D(n19546), .CK(clk), .Q(\mem[820][0] ) );
  DFF_X1 \mem_reg[819][7]  ( .D(n19547), .CK(clk), .Q(\mem[819][7] ) );
  DFF_X1 \mem_reg[819][6]  ( .D(n19548), .CK(clk), .Q(\mem[819][6] ) );
  DFF_X1 \mem_reg[819][5]  ( .D(n19549), .CK(clk), .Q(\mem[819][5] ) );
  DFF_X1 \mem_reg[819][4]  ( .D(n19550), .CK(clk), .Q(\mem[819][4] ) );
  DFF_X1 \mem_reg[819][3]  ( .D(n19551), .CK(clk), .Q(\mem[819][3] ) );
  DFF_X1 \mem_reg[819][2]  ( .D(n19552), .CK(clk), .Q(\mem[819][2] ) );
  DFF_X1 \mem_reg[819][1]  ( .D(n19553), .CK(clk), .Q(\mem[819][1] ) );
  DFF_X1 \mem_reg[819][0]  ( .D(n19554), .CK(clk), .Q(\mem[819][0] ) );
  DFF_X1 \mem_reg[818][7]  ( .D(n19555), .CK(clk), .Q(\mem[818][7] ) );
  DFF_X1 \mem_reg[818][6]  ( .D(n19556), .CK(clk), .Q(\mem[818][6] ) );
  DFF_X1 \mem_reg[818][5]  ( .D(n19557), .CK(clk), .Q(\mem[818][5] ) );
  DFF_X1 \mem_reg[818][4]  ( .D(n19558), .CK(clk), .Q(\mem[818][4] ) );
  DFF_X1 \mem_reg[818][3]  ( .D(n19559), .CK(clk), .Q(\mem[818][3] ) );
  DFF_X1 \mem_reg[818][2]  ( .D(n19560), .CK(clk), .Q(\mem[818][2] ) );
  DFF_X1 \mem_reg[818][1]  ( .D(n19561), .CK(clk), .Q(\mem[818][1] ) );
  DFF_X1 \mem_reg[818][0]  ( .D(n19562), .CK(clk), .Q(\mem[818][0] ) );
  DFF_X1 \mem_reg[817][7]  ( .D(n19563), .CK(clk), .Q(\mem[817][7] ) );
  DFF_X1 \mem_reg[817][6]  ( .D(n19564), .CK(clk), .Q(\mem[817][6] ) );
  DFF_X1 \mem_reg[817][5]  ( .D(n19565), .CK(clk), .Q(\mem[817][5] ) );
  DFF_X1 \mem_reg[817][4]  ( .D(n19566), .CK(clk), .Q(\mem[817][4] ) );
  DFF_X1 \mem_reg[817][3]  ( .D(n19567), .CK(clk), .Q(\mem[817][3] ) );
  DFF_X1 \mem_reg[817][2]  ( .D(n19568), .CK(clk), .Q(\mem[817][2] ) );
  DFF_X1 \mem_reg[817][1]  ( .D(n19569), .CK(clk), .Q(\mem[817][1] ) );
  DFF_X1 \mem_reg[817][0]  ( .D(n19570), .CK(clk), .Q(\mem[817][0] ) );
  DFF_X1 \mem_reg[816][7]  ( .D(n19571), .CK(clk), .Q(\mem[816][7] ) );
  DFF_X1 \mem_reg[816][6]  ( .D(n19572), .CK(clk), .Q(\mem[816][6] ) );
  DFF_X1 \mem_reg[816][5]  ( .D(n19573), .CK(clk), .Q(\mem[816][5] ) );
  DFF_X1 \mem_reg[816][4]  ( .D(n19574), .CK(clk), .Q(\mem[816][4] ) );
  DFF_X1 \mem_reg[816][3]  ( .D(n19575), .CK(clk), .Q(\mem[816][3] ) );
  DFF_X1 \mem_reg[816][2]  ( .D(n19576), .CK(clk), .Q(\mem[816][2] ) );
  DFF_X1 \mem_reg[816][1]  ( .D(n19577), .CK(clk), .Q(\mem[816][1] ) );
  DFF_X1 \mem_reg[816][0]  ( .D(n19578), .CK(clk), .Q(\mem[816][0] ) );
  DFF_X1 \mem_reg[815][7]  ( .D(n19579), .CK(clk), .Q(\mem[815][7] ) );
  DFF_X1 \mem_reg[815][6]  ( .D(n19580), .CK(clk), .Q(\mem[815][6] ) );
  DFF_X1 \mem_reg[815][5]  ( .D(n19581), .CK(clk), .Q(\mem[815][5] ) );
  DFF_X1 \mem_reg[815][4]  ( .D(n19582), .CK(clk), .Q(\mem[815][4] ) );
  DFF_X1 \mem_reg[815][3]  ( .D(n19583), .CK(clk), .Q(\mem[815][3] ) );
  DFF_X1 \mem_reg[815][2]  ( .D(n19584), .CK(clk), .Q(\mem[815][2] ) );
  DFF_X1 \mem_reg[815][1]  ( .D(n19585), .CK(clk), .Q(\mem[815][1] ) );
  DFF_X1 \mem_reg[815][0]  ( .D(n19586), .CK(clk), .Q(\mem[815][0] ) );
  DFF_X1 \mem_reg[814][7]  ( .D(n19587), .CK(clk), .Q(\mem[814][7] ) );
  DFF_X1 \mem_reg[814][6]  ( .D(n19588), .CK(clk), .Q(\mem[814][6] ) );
  DFF_X1 \mem_reg[814][5]  ( .D(n19589), .CK(clk), .Q(\mem[814][5] ) );
  DFF_X1 \mem_reg[814][4]  ( .D(n19590), .CK(clk), .Q(\mem[814][4] ) );
  DFF_X1 \mem_reg[814][3]  ( .D(n19591), .CK(clk), .Q(\mem[814][3] ) );
  DFF_X1 \mem_reg[814][2]  ( .D(n19592), .CK(clk), .Q(\mem[814][2] ) );
  DFF_X1 \mem_reg[814][1]  ( .D(n19593), .CK(clk), .Q(\mem[814][1] ) );
  DFF_X1 \mem_reg[814][0]  ( .D(n19594), .CK(clk), .Q(\mem[814][0] ) );
  DFF_X1 \mem_reg[813][7]  ( .D(n19595), .CK(clk), .Q(\mem[813][7] ) );
  DFF_X1 \mem_reg[813][6]  ( .D(n19596), .CK(clk), .Q(\mem[813][6] ) );
  DFF_X1 \mem_reg[813][5]  ( .D(n19597), .CK(clk), .Q(\mem[813][5] ) );
  DFF_X1 \mem_reg[813][4]  ( .D(n19598), .CK(clk), .Q(\mem[813][4] ) );
  DFF_X1 \mem_reg[813][3]  ( .D(n19599), .CK(clk), .Q(\mem[813][3] ) );
  DFF_X1 \mem_reg[813][2]  ( .D(n19600), .CK(clk), .Q(\mem[813][2] ) );
  DFF_X1 \mem_reg[813][1]  ( .D(n19601), .CK(clk), .Q(\mem[813][1] ) );
  DFF_X1 \mem_reg[813][0]  ( .D(n19602), .CK(clk), .Q(\mem[813][0] ) );
  DFF_X1 \mem_reg[812][7]  ( .D(n19603), .CK(clk), .Q(\mem[812][7] ) );
  DFF_X1 \mem_reg[812][6]  ( .D(n19604), .CK(clk), .Q(\mem[812][6] ) );
  DFF_X1 \mem_reg[812][5]  ( .D(n19605), .CK(clk), .Q(\mem[812][5] ) );
  DFF_X1 \mem_reg[812][4]  ( .D(n19606), .CK(clk), .Q(\mem[812][4] ) );
  DFF_X1 \mem_reg[812][3]  ( .D(n19607), .CK(clk), .Q(\mem[812][3] ) );
  DFF_X1 \mem_reg[812][2]  ( .D(n19608), .CK(clk), .Q(\mem[812][2] ) );
  DFF_X1 \mem_reg[812][1]  ( .D(n19609), .CK(clk), .Q(\mem[812][1] ) );
  DFF_X1 \mem_reg[812][0]  ( .D(n19610), .CK(clk), .Q(\mem[812][0] ) );
  DFF_X1 \mem_reg[811][7]  ( .D(n19611), .CK(clk), .Q(\mem[811][7] ) );
  DFF_X1 \mem_reg[811][6]  ( .D(n19612), .CK(clk), .Q(\mem[811][6] ) );
  DFF_X1 \mem_reg[811][5]  ( .D(n19613), .CK(clk), .Q(\mem[811][5] ) );
  DFF_X1 \mem_reg[811][4]  ( .D(n19614), .CK(clk), .Q(\mem[811][4] ) );
  DFF_X1 \mem_reg[811][3]  ( .D(n19615), .CK(clk), .Q(\mem[811][3] ) );
  DFF_X1 \mem_reg[811][2]  ( .D(n19616), .CK(clk), .Q(\mem[811][2] ) );
  DFF_X1 \mem_reg[811][1]  ( .D(n19617), .CK(clk), .Q(\mem[811][1] ) );
  DFF_X1 \mem_reg[811][0]  ( .D(n19618), .CK(clk), .Q(\mem[811][0] ) );
  DFF_X1 \mem_reg[810][7]  ( .D(n19619), .CK(clk), .Q(\mem[810][7] ) );
  DFF_X1 \mem_reg[810][6]  ( .D(n19620), .CK(clk), .Q(\mem[810][6] ) );
  DFF_X1 \mem_reg[810][5]  ( .D(n19621), .CK(clk), .Q(\mem[810][5] ) );
  DFF_X1 \mem_reg[810][4]  ( .D(n19622), .CK(clk), .Q(\mem[810][4] ) );
  DFF_X1 \mem_reg[810][3]  ( .D(n19623), .CK(clk), .Q(\mem[810][3] ) );
  DFF_X1 \mem_reg[810][2]  ( .D(n19624), .CK(clk), .Q(\mem[810][2] ) );
  DFF_X1 \mem_reg[810][1]  ( .D(n19625), .CK(clk), .Q(\mem[810][1] ) );
  DFF_X1 \mem_reg[810][0]  ( .D(n19626), .CK(clk), .Q(\mem[810][0] ) );
  DFF_X1 \mem_reg[809][7]  ( .D(n19627), .CK(clk), .Q(\mem[809][7] ) );
  DFF_X1 \mem_reg[809][6]  ( .D(n19628), .CK(clk), .Q(\mem[809][6] ) );
  DFF_X1 \mem_reg[809][5]  ( .D(n19629), .CK(clk), .Q(\mem[809][5] ) );
  DFF_X1 \mem_reg[809][4]  ( .D(n19630), .CK(clk), .Q(\mem[809][4] ) );
  DFF_X1 \mem_reg[809][3]  ( .D(n19631), .CK(clk), .Q(\mem[809][3] ) );
  DFF_X1 \mem_reg[809][2]  ( .D(n19632), .CK(clk), .Q(\mem[809][2] ) );
  DFF_X1 \mem_reg[809][1]  ( .D(n19633), .CK(clk), .Q(\mem[809][1] ) );
  DFF_X1 \mem_reg[809][0]  ( .D(n19634), .CK(clk), .Q(\mem[809][0] ) );
  DFF_X1 \mem_reg[808][7]  ( .D(n19635), .CK(clk), .Q(\mem[808][7] ) );
  DFF_X1 \mem_reg[808][6]  ( .D(n19636), .CK(clk), .Q(\mem[808][6] ) );
  DFF_X1 \mem_reg[808][5]  ( .D(n19637), .CK(clk), .Q(\mem[808][5] ) );
  DFF_X1 \mem_reg[808][4]  ( .D(n19638), .CK(clk), .Q(\mem[808][4] ) );
  DFF_X1 \mem_reg[808][3]  ( .D(n19639), .CK(clk), .Q(\mem[808][3] ) );
  DFF_X1 \mem_reg[808][2]  ( .D(n19640), .CK(clk), .Q(\mem[808][2] ) );
  DFF_X1 \mem_reg[808][1]  ( .D(n19641), .CK(clk), .Q(\mem[808][1] ) );
  DFF_X1 \mem_reg[808][0]  ( .D(n19642), .CK(clk), .Q(\mem[808][0] ) );
  DFF_X1 \mem_reg[807][7]  ( .D(n19643), .CK(clk), .Q(\mem[807][7] ) );
  DFF_X1 \mem_reg[807][6]  ( .D(n19644), .CK(clk), .Q(\mem[807][6] ) );
  DFF_X1 \mem_reg[807][5]  ( .D(n19645), .CK(clk), .Q(\mem[807][5] ) );
  DFF_X1 \mem_reg[807][4]  ( .D(n19646), .CK(clk), .Q(\mem[807][4] ) );
  DFF_X1 \mem_reg[807][3]  ( .D(n19647), .CK(clk), .Q(\mem[807][3] ) );
  DFF_X1 \mem_reg[807][2]  ( .D(n19648), .CK(clk), .Q(\mem[807][2] ) );
  DFF_X1 \mem_reg[807][1]  ( .D(n19649), .CK(clk), .Q(\mem[807][1] ) );
  DFF_X1 \mem_reg[807][0]  ( .D(n19650), .CK(clk), .Q(\mem[807][0] ) );
  DFF_X1 \mem_reg[806][7]  ( .D(n19651), .CK(clk), .Q(\mem[806][7] ) );
  DFF_X1 \mem_reg[806][6]  ( .D(n19652), .CK(clk), .Q(\mem[806][6] ) );
  DFF_X1 \mem_reg[806][5]  ( .D(n19653), .CK(clk), .Q(\mem[806][5] ) );
  DFF_X1 \mem_reg[806][4]  ( .D(n19654), .CK(clk), .Q(\mem[806][4] ) );
  DFF_X1 \mem_reg[806][3]  ( .D(n19655), .CK(clk), .Q(\mem[806][3] ) );
  DFF_X1 \mem_reg[806][2]  ( .D(n19656), .CK(clk), .Q(\mem[806][2] ) );
  DFF_X1 \mem_reg[806][1]  ( .D(n19657), .CK(clk), .Q(\mem[806][1] ) );
  DFF_X1 \mem_reg[806][0]  ( .D(n19658), .CK(clk), .Q(\mem[806][0] ) );
  DFF_X1 \mem_reg[805][7]  ( .D(n19659), .CK(clk), .Q(\mem[805][7] ) );
  DFF_X1 \mem_reg[805][6]  ( .D(n19660), .CK(clk), .Q(\mem[805][6] ) );
  DFF_X1 \mem_reg[805][5]  ( .D(n19661), .CK(clk), .Q(\mem[805][5] ) );
  DFF_X1 \mem_reg[805][4]  ( .D(n19662), .CK(clk), .Q(\mem[805][4] ) );
  DFF_X1 \mem_reg[805][3]  ( .D(n19663), .CK(clk), .Q(\mem[805][3] ) );
  DFF_X1 \mem_reg[805][2]  ( .D(n19664), .CK(clk), .Q(\mem[805][2] ) );
  DFF_X1 \mem_reg[805][1]  ( .D(n19665), .CK(clk), .Q(\mem[805][1] ) );
  DFF_X1 \mem_reg[805][0]  ( .D(n19666), .CK(clk), .Q(\mem[805][0] ) );
  DFF_X1 \mem_reg[804][7]  ( .D(n19667), .CK(clk), .Q(\mem[804][7] ) );
  DFF_X1 \mem_reg[804][6]  ( .D(n19668), .CK(clk), .Q(\mem[804][6] ) );
  DFF_X1 \mem_reg[804][5]  ( .D(n19669), .CK(clk), .Q(\mem[804][5] ) );
  DFF_X1 \mem_reg[804][4]  ( .D(n19670), .CK(clk), .Q(\mem[804][4] ) );
  DFF_X1 \mem_reg[804][3]  ( .D(n19671), .CK(clk), .Q(\mem[804][3] ) );
  DFF_X1 \mem_reg[804][2]  ( .D(n19672), .CK(clk), .Q(\mem[804][2] ) );
  DFF_X1 \mem_reg[804][1]  ( .D(n19673), .CK(clk), .Q(\mem[804][1] ) );
  DFF_X1 \mem_reg[804][0]  ( .D(n19674), .CK(clk), .Q(\mem[804][0] ) );
  DFF_X1 \mem_reg[803][7]  ( .D(n19675), .CK(clk), .Q(\mem[803][7] ) );
  DFF_X1 \mem_reg[803][6]  ( .D(n19676), .CK(clk), .Q(\mem[803][6] ) );
  DFF_X1 \mem_reg[803][5]  ( .D(n19677), .CK(clk), .Q(\mem[803][5] ) );
  DFF_X1 \mem_reg[803][4]  ( .D(n19678), .CK(clk), .Q(\mem[803][4] ) );
  DFF_X1 \mem_reg[803][3]  ( .D(n19679), .CK(clk), .Q(\mem[803][3] ) );
  DFF_X1 \mem_reg[803][2]  ( .D(n19680), .CK(clk), .Q(\mem[803][2] ) );
  DFF_X1 \mem_reg[803][1]  ( .D(n19681), .CK(clk), .Q(\mem[803][1] ) );
  DFF_X1 \mem_reg[803][0]  ( .D(n19682), .CK(clk), .Q(\mem[803][0] ) );
  DFF_X1 \mem_reg[802][7]  ( .D(n19683), .CK(clk), .Q(\mem[802][7] ) );
  DFF_X1 \mem_reg[802][6]  ( .D(n19684), .CK(clk), .Q(\mem[802][6] ) );
  DFF_X1 \mem_reg[802][5]  ( .D(n19685), .CK(clk), .Q(\mem[802][5] ) );
  DFF_X1 \mem_reg[802][4]  ( .D(n19686), .CK(clk), .Q(\mem[802][4] ) );
  DFF_X1 \mem_reg[802][3]  ( .D(n19687), .CK(clk), .Q(\mem[802][3] ) );
  DFF_X1 \mem_reg[802][2]  ( .D(n19688), .CK(clk), .Q(\mem[802][2] ) );
  DFF_X1 \mem_reg[802][1]  ( .D(n19689), .CK(clk), .Q(\mem[802][1] ) );
  DFF_X1 \mem_reg[802][0]  ( .D(n19690), .CK(clk), .Q(\mem[802][0] ) );
  DFF_X1 \mem_reg[801][7]  ( .D(n19691), .CK(clk), .Q(\mem[801][7] ) );
  DFF_X1 \mem_reg[801][6]  ( .D(n19692), .CK(clk), .Q(\mem[801][6] ) );
  DFF_X1 \mem_reg[801][5]  ( .D(n19693), .CK(clk), .Q(\mem[801][5] ) );
  DFF_X1 \mem_reg[801][4]  ( .D(n19694), .CK(clk), .Q(\mem[801][4] ) );
  DFF_X1 \mem_reg[801][3]  ( .D(n19695), .CK(clk), .Q(\mem[801][3] ) );
  DFF_X1 \mem_reg[801][2]  ( .D(n19696), .CK(clk), .Q(\mem[801][2] ) );
  DFF_X1 \mem_reg[801][1]  ( .D(n19697), .CK(clk), .Q(\mem[801][1] ) );
  DFF_X1 \mem_reg[801][0]  ( .D(n19698), .CK(clk), .Q(\mem[801][0] ) );
  DFF_X1 \mem_reg[800][7]  ( .D(n19699), .CK(clk), .Q(\mem[800][7] ) );
  DFF_X1 \mem_reg[800][6]  ( .D(n19700), .CK(clk), .Q(\mem[800][6] ) );
  DFF_X1 \mem_reg[800][5]  ( .D(n19701), .CK(clk), .Q(\mem[800][5] ) );
  DFF_X1 \mem_reg[800][4]  ( .D(n19702), .CK(clk), .Q(\mem[800][4] ) );
  DFF_X1 \mem_reg[800][3]  ( .D(n19703), .CK(clk), .Q(\mem[800][3] ) );
  DFF_X1 \mem_reg[800][2]  ( .D(n19704), .CK(clk), .Q(\mem[800][2] ) );
  DFF_X1 \mem_reg[800][1]  ( .D(n19705), .CK(clk), .Q(\mem[800][1] ) );
  DFF_X1 \mem_reg[800][0]  ( .D(n19706), .CK(clk), .Q(\mem[800][0] ) );
  DFF_X1 \mem_reg[799][7]  ( .D(n19707), .CK(clk), .Q(\mem[799][7] ) );
  DFF_X1 \mem_reg[799][6]  ( .D(n19708), .CK(clk), .Q(\mem[799][6] ) );
  DFF_X1 \mem_reg[799][5]  ( .D(n19709), .CK(clk), .Q(\mem[799][5] ) );
  DFF_X1 \mem_reg[799][4]  ( .D(n19710), .CK(clk), .Q(\mem[799][4] ) );
  DFF_X1 \mem_reg[799][3]  ( .D(n19711), .CK(clk), .Q(\mem[799][3] ) );
  DFF_X1 \mem_reg[799][2]  ( .D(n19712), .CK(clk), .Q(\mem[799][2] ) );
  DFF_X1 \mem_reg[799][1]  ( .D(n19713), .CK(clk), .Q(\mem[799][1] ) );
  DFF_X1 \mem_reg[799][0]  ( .D(n19714), .CK(clk), .Q(\mem[799][0] ) );
  DFF_X1 \mem_reg[798][7]  ( .D(n19715), .CK(clk), .Q(\mem[798][7] ) );
  DFF_X1 \mem_reg[798][6]  ( .D(n19716), .CK(clk), .Q(\mem[798][6] ) );
  DFF_X1 \mem_reg[798][5]  ( .D(n19717), .CK(clk), .Q(\mem[798][5] ) );
  DFF_X1 \mem_reg[798][4]  ( .D(n19718), .CK(clk), .Q(\mem[798][4] ) );
  DFF_X1 \mem_reg[798][3]  ( .D(n19719), .CK(clk), .Q(\mem[798][3] ) );
  DFF_X1 \mem_reg[798][2]  ( .D(n19720), .CK(clk), .Q(\mem[798][2] ) );
  DFF_X1 \mem_reg[798][1]  ( .D(n19721), .CK(clk), .Q(\mem[798][1] ) );
  DFF_X1 \mem_reg[798][0]  ( .D(n19722), .CK(clk), .Q(\mem[798][0] ) );
  DFF_X1 \mem_reg[797][7]  ( .D(n19723), .CK(clk), .Q(\mem[797][7] ) );
  DFF_X1 \mem_reg[797][6]  ( .D(n19724), .CK(clk), .Q(\mem[797][6] ) );
  DFF_X1 \mem_reg[797][5]  ( .D(n19725), .CK(clk), .Q(\mem[797][5] ) );
  DFF_X1 \mem_reg[797][4]  ( .D(n19726), .CK(clk), .Q(\mem[797][4] ) );
  DFF_X1 \mem_reg[797][3]  ( .D(n19727), .CK(clk), .Q(\mem[797][3] ) );
  DFF_X1 \mem_reg[797][2]  ( .D(n19728), .CK(clk), .Q(\mem[797][2] ) );
  DFF_X1 \mem_reg[797][1]  ( .D(n19729), .CK(clk), .Q(\mem[797][1] ) );
  DFF_X1 \mem_reg[797][0]  ( .D(n19730), .CK(clk), .Q(\mem[797][0] ) );
  DFF_X1 \mem_reg[796][7]  ( .D(n19731), .CK(clk), .Q(\mem[796][7] ) );
  DFF_X1 \mem_reg[796][6]  ( .D(n19732), .CK(clk), .Q(\mem[796][6] ) );
  DFF_X1 \mem_reg[796][5]  ( .D(n19733), .CK(clk), .Q(\mem[796][5] ) );
  DFF_X1 \mem_reg[796][4]  ( .D(n19734), .CK(clk), .Q(\mem[796][4] ) );
  DFF_X1 \mem_reg[796][3]  ( .D(n19735), .CK(clk), .Q(\mem[796][3] ) );
  DFF_X1 \mem_reg[796][2]  ( .D(n19736), .CK(clk), .Q(\mem[796][2] ) );
  DFF_X1 \mem_reg[796][1]  ( .D(n19737), .CK(clk), .Q(\mem[796][1] ) );
  DFF_X1 \mem_reg[796][0]  ( .D(n19738), .CK(clk), .Q(\mem[796][0] ) );
  DFF_X1 \mem_reg[795][7]  ( .D(n19739), .CK(clk), .Q(\mem[795][7] ) );
  DFF_X1 \mem_reg[795][6]  ( .D(n19740), .CK(clk), .Q(\mem[795][6] ) );
  DFF_X1 \mem_reg[795][5]  ( .D(n19741), .CK(clk), .Q(\mem[795][5] ) );
  DFF_X1 \mem_reg[795][4]  ( .D(n19742), .CK(clk), .Q(\mem[795][4] ) );
  DFF_X1 \mem_reg[795][3]  ( .D(n19743), .CK(clk), .Q(\mem[795][3] ) );
  DFF_X1 \mem_reg[795][2]  ( .D(n19744), .CK(clk), .Q(\mem[795][2] ) );
  DFF_X1 \mem_reg[795][1]  ( .D(n19745), .CK(clk), .Q(\mem[795][1] ) );
  DFF_X1 \mem_reg[795][0]  ( .D(n19746), .CK(clk), .Q(\mem[795][0] ) );
  DFF_X1 \mem_reg[794][7]  ( .D(n19747), .CK(clk), .Q(\mem[794][7] ) );
  DFF_X1 \mem_reg[794][6]  ( .D(n19748), .CK(clk), .Q(\mem[794][6] ) );
  DFF_X1 \mem_reg[794][5]  ( .D(n19749), .CK(clk), .Q(\mem[794][5] ) );
  DFF_X1 \mem_reg[794][4]  ( .D(n19750), .CK(clk), .Q(\mem[794][4] ) );
  DFF_X1 \mem_reg[794][3]  ( .D(n19751), .CK(clk), .Q(\mem[794][3] ) );
  DFF_X1 \mem_reg[794][2]  ( .D(n19752), .CK(clk), .Q(\mem[794][2] ) );
  DFF_X1 \mem_reg[794][1]  ( .D(n19753), .CK(clk), .Q(\mem[794][1] ) );
  DFF_X1 \mem_reg[794][0]  ( .D(n19754), .CK(clk), .Q(\mem[794][0] ) );
  DFF_X1 \mem_reg[793][7]  ( .D(n19755), .CK(clk), .Q(\mem[793][7] ) );
  DFF_X1 \mem_reg[793][6]  ( .D(n19756), .CK(clk), .Q(\mem[793][6] ) );
  DFF_X1 \mem_reg[793][5]  ( .D(n19757), .CK(clk), .Q(\mem[793][5] ) );
  DFF_X1 \mem_reg[793][4]  ( .D(n19758), .CK(clk), .Q(\mem[793][4] ) );
  DFF_X1 \mem_reg[793][3]  ( .D(n19759), .CK(clk), .Q(\mem[793][3] ) );
  DFF_X1 \mem_reg[793][2]  ( .D(n19760), .CK(clk), .Q(\mem[793][2] ) );
  DFF_X1 \mem_reg[793][1]  ( .D(n19761), .CK(clk), .Q(\mem[793][1] ) );
  DFF_X1 \mem_reg[793][0]  ( .D(n19762), .CK(clk), .Q(\mem[793][0] ) );
  DFF_X1 \mem_reg[792][7]  ( .D(n19763), .CK(clk), .Q(\mem[792][7] ) );
  DFF_X1 \mem_reg[792][6]  ( .D(n19764), .CK(clk), .Q(\mem[792][6] ) );
  DFF_X1 \mem_reg[792][5]  ( .D(n19765), .CK(clk), .Q(\mem[792][5] ) );
  DFF_X1 \mem_reg[792][4]  ( .D(n19766), .CK(clk), .Q(\mem[792][4] ) );
  DFF_X1 \mem_reg[792][3]  ( .D(n19767), .CK(clk), .Q(\mem[792][3] ) );
  DFF_X1 \mem_reg[792][2]  ( .D(n19768), .CK(clk), .Q(\mem[792][2] ) );
  DFF_X1 \mem_reg[792][1]  ( .D(n19769), .CK(clk), .Q(\mem[792][1] ) );
  DFF_X1 \mem_reg[792][0]  ( .D(n19770), .CK(clk), .Q(\mem[792][0] ) );
  DFF_X1 \mem_reg[791][7]  ( .D(n19771), .CK(clk), .Q(\mem[791][7] ) );
  DFF_X1 \mem_reg[791][6]  ( .D(n19772), .CK(clk), .Q(\mem[791][6] ) );
  DFF_X1 \mem_reg[791][5]  ( .D(n19773), .CK(clk), .Q(\mem[791][5] ) );
  DFF_X1 \mem_reg[791][4]  ( .D(n19774), .CK(clk), .Q(\mem[791][4] ) );
  DFF_X1 \mem_reg[791][3]  ( .D(n19775), .CK(clk), .Q(\mem[791][3] ) );
  DFF_X1 \mem_reg[791][2]  ( .D(n19776), .CK(clk), .Q(\mem[791][2] ) );
  DFF_X1 \mem_reg[791][1]  ( .D(n19777), .CK(clk), .Q(\mem[791][1] ) );
  DFF_X1 \mem_reg[791][0]  ( .D(n19778), .CK(clk), .Q(\mem[791][0] ) );
  DFF_X1 \mem_reg[790][7]  ( .D(n19779), .CK(clk), .Q(\mem[790][7] ) );
  DFF_X1 \mem_reg[790][6]  ( .D(n19780), .CK(clk), .Q(\mem[790][6] ) );
  DFF_X1 \mem_reg[790][5]  ( .D(n19781), .CK(clk), .Q(\mem[790][5] ) );
  DFF_X1 \mem_reg[790][4]  ( .D(n19782), .CK(clk), .Q(\mem[790][4] ) );
  DFF_X1 \mem_reg[790][3]  ( .D(n19783), .CK(clk), .Q(\mem[790][3] ) );
  DFF_X1 \mem_reg[790][2]  ( .D(n19784), .CK(clk), .Q(\mem[790][2] ) );
  DFF_X1 \mem_reg[790][1]  ( .D(n19785), .CK(clk), .Q(\mem[790][1] ) );
  DFF_X1 \mem_reg[790][0]  ( .D(n19786), .CK(clk), .Q(\mem[790][0] ) );
  DFF_X1 \mem_reg[789][7]  ( .D(n19787), .CK(clk), .Q(\mem[789][7] ) );
  DFF_X1 \mem_reg[789][6]  ( .D(n19788), .CK(clk), .Q(\mem[789][6] ) );
  DFF_X1 \mem_reg[789][5]  ( .D(n19789), .CK(clk), .Q(\mem[789][5] ) );
  DFF_X1 \mem_reg[789][4]  ( .D(n19790), .CK(clk), .Q(\mem[789][4] ) );
  DFF_X1 \mem_reg[789][3]  ( .D(n19791), .CK(clk), .Q(\mem[789][3] ) );
  DFF_X1 \mem_reg[789][2]  ( .D(n19792), .CK(clk), .Q(\mem[789][2] ) );
  DFF_X1 \mem_reg[789][1]  ( .D(n19793), .CK(clk), .Q(\mem[789][1] ) );
  DFF_X1 \mem_reg[789][0]  ( .D(n19794), .CK(clk), .Q(\mem[789][0] ) );
  DFF_X1 \mem_reg[788][7]  ( .D(n19795), .CK(clk), .Q(\mem[788][7] ) );
  DFF_X1 \mem_reg[788][6]  ( .D(n19796), .CK(clk), .Q(\mem[788][6] ) );
  DFF_X1 \mem_reg[788][5]  ( .D(n19797), .CK(clk), .Q(\mem[788][5] ) );
  DFF_X1 \mem_reg[788][4]  ( .D(n19798), .CK(clk), .Q(\mem[788][4] ) );
  DFF_X1 \mem_reg[788][3]  ( .D(n19799), .CK(clk), .Q(\mem[788][3] ) );
  DFF_X1 \mem_reg[788][2]  ( .D(n19800), .CK(clk), .Q(\mem[788][2] ) );
  DFF_X1 \mem_reg[788][1]  ( .D(n19801), .CK(clk), .Q(\mem[788][1] ) );
  DFF_X1 \mem_reg[788][0]  ( .D(n19802), .CK(clk), .Q(\mem[788][0] ) );
  DFF_X1 \mem_reg[787][7]  ( .D(n19803), .CK(clk), .Q(\mem[787][7] ) );
  DFF_X1 \mem_reg[787][6]  ( .D(n19804), .CK(clk), .Q(\mem[787][6] ) );
  DFF_X1 \mem_reg[787][5]  ( .D(n19805), .CK(clk), .Q(\mem[787][5] ) );
  DFF_X1 \mem_reg[787][4]  ( .D(n19806), .CK(clk), .Q(\mem[787][4] ) );
  DFF_X1 \mem_reg[787][3]  ( .D(n19807), .CK(clk), .Q(\mem[787][3] ) );
  DFF_X1 \mem_reg[787][2]  ( .D(n19808), .CK(clk), .Q(\mem[787][2] ) );
  DFF_X1 \mem_reg[787][1]  ( .D(n19809), .CK(clk), .Q(\mem[787][1] ) );
  DFF_X1 \mem_reg[787][0]  ( .D(n19810), .CK(clk), .Q(\mem[787][0] ) );
  DFF_X1 \mem_reg[786][7]  ( .D(n19811), .CK(clk), .Q(\mem[786][7] ) );
  DFF_X1 \mem_reg[786][6]  ( .D(n19812), .CK(clk), .Q(\mem[786][6] ) );
  DFF_X1 \mem_reg[786][5]  ( .D(n19813), .CK(clk), .Q(\mem[786][5] ) );
  DFF_X1 \mem_reg[786][4]  ( .D(n19814), .CK(clk), .Q(\mem[786][4] ) );
  DFF_X1 \mem_reg[786][3]  ( .D(n19815), .CK(clk), .Q(\mem[786][3] ) );
  DFF_X1 \mem_reg[786][2]  ( .D(n19816), .CK(clk), .Q(\mem[786][2] ) );
  DFF_X1 \mem_reg[786][1]  ( .D(n19817), .CK(clk), .Q(\mem[786][1] ) );
  DFF_X1 \mem_reg[786][0]  ( .D(n19818), .CK(clk), .Q(\mem[786][0] ) );
  DFF_X1 \mem_reg[785][7]  ( .D(n19819), .CK(clk), .Q(\mem[785][7] ) );
  DFF_X1 \mem_reg[785][6]  ( .D(n19820), .CK(clk), .Q(\mem[785][6] ) );
  DFF_X1 \mem_reg[785][5]  ( .D(n19821), .CK(clk), .Q(\mem[785][5] ) );
  DFF_X1 \mem_reg[785][4]  ( .D(n19822), .CK(clk), .Q(\mem[785][4] ) );
  DFF_X1 \mem_reg[785][3]  ( .D(n19823), .CK(clk), .Q(\mem[785][3] ) );
  DFF_X1 \mem_reg[785][2]  ( .D(n19824), .CK(clk), .Q(\mem[785][2] ) );
  DFF_X1 \mem_reg[785][1]  ( .D(n19825), .CK(clk), .Q(\mem[785][1] ) );
  DFF_X1 \mem_reg[785][0]  ( .D(n19826), .CK(clk), .Q(\mem[785][0] ) );
  DFF_X1 \mem_reg[784][7]  ( .D(n19827), .CK(clk), .Q(\mem[784][7] ) );
  DFF_X1 \mem_reg[784][6]  ( .D(n19828), .CK(clk), .Q(\mem[784][6] ) );
  DFF_X1 \mem_reg[784][5]  ( .D(n19829), .CK(clk), .Q(\mem[784][5] ) );
  DFF_X1 \mem_reg[784][4]  ( .D(n19830), .CK(clk), .Q(\mem[784][4] ) );
  DFF_X1 \mem_reg[784][3]  ( .D(n19831), .CK(clk), .Q(\mem[784][3] ) );
  DFF_X1 \mem_reg[784][2]  ( .D(n19832), .CK(clk), .Q(\mem[784][2] ) );
  DFF_X1 \mem_reg[784][1]  ( .D(n19833), .CK(clk), .Q(\mem[784][1] ) );
  DFF_X1 \mem_reg[784][0]  ( .D(n19834), .CK(clk), .Q(\mem[784][0] ) );
  DFF_X1 \mem_reg[783][7]  ( .D(n19835), .CK(clk), .Q(\mem[783][7] ) );
  DFF_X1 \mem_reg[783][6]  ( .D(n19836), .CK(clk), .Q(\mem[783][6] ) );
  DFF_X1 \mem_reg[783][5]  ( .D(n19837), .CK(clk), .Q(\mem[783][5] ) );
  DFF_X1 \mem_reg[783][4]  ( .D(n19838), .CK(clk), .Q(\mem[783][4] ) );
  DFF_X1 \mem_reg[783][3]  ( .D(n19839), .CK(clk), .Q(\mem[783][3] ) );
  DFF_X1 \mem_reg[783][2]  ( .D(n19840), .CK(clk), .Q(\mem[783][2] ) );
  DFF_X1 \mem_reg[783][1]  ( .D(n19841), .CK(clk), .Q(\mem[783][1] ) );
  DFF_X1 \mem_reg[783][0]  ( .D(n19842), .CK(clk), .Q(\mem[783][0] ) );
  DFF_X1 \mem_reg[782][7]  ( .D(n19843), .CK(clk), .Q(\mem[782][7] ) );
  DFF_X1 \mem_reg[782][6]  ( .D(n19844), .CK(clk), .Q(\mem[782][6] ) );
  DFF_X1 \mem_reg[782][5]  ( .D(n19845), .CK(clk), .Q(\mem[782][5] ) );
  DFF_X1 \mem_reg[782][4]  ( .D(n19846), .CK(clk), .Q(\mem[782][4] ) );
  DFF_X1 \mem_reg[782][3]  ( .D(n19847), .CK(clk), .Q(\mem[782][3] ) );
  DFF_X1 \mem_reg[782][2]  ( .D(n19848), .CK(clk), .Q(\mem[782][2] ) );
  DFF_X1 \mem_reg[782][1]  ( .D(n19849), .CK(clk), .Q(\mem[782][1] ) );
  DFF_X1 \mem_reg[782][0]  ( .D(n19850), .CK(clk), .Q(\mem[782][0] ) );
  DFF_X1 \mem_reg[781][7]  ( .D(n19851), .CK(clk), .Q(\mem[781][7] ) );
  DFF_X1 \mem_reg[781][6]  ( .D(n19852), .CK(clk), .Q(\mem[781][6] ) );
  DFF_X1 \mem_reg[781][5]  ( .D(n19853), .CK(clk), .Q(\mem[781][5] ) );
  DFF_X1 \mem_reg[781][4]  ( .D(n19854), .CK(clk), .Q(\mem[781][4] ) );
  DFF_X1 \mem_reg[781][3]  ( .D(n19855), .CK(clk), .Q(\mem[781][3] ) );
  DFF_X1 \mem_reg[781][2]  ( .D(n19856), .CK(clk), .Q(\mem[781][2] ) );
  DFF_X1 \mem_reg[781][1]  ( .D(n19857), .CK(clk), .Q(\mem[781][1] ) );
  DFF_X1 \mem_reg[781][0]  ( .D(n19858), .CK(clk), .Q(\mem[781][0] ) );
  DFF_X1 \mem_reg[780][7]  ( .D(n19859), .CK(clk), .Q(\mem[780][7] ) );
  DFF_X1 \mem_reg[780][6]  ( .D(n19860), .CK(clk), .Q(\mem[780][6] ) );
  DFF_X1 \mem_reg[780][5]  ( .D(n19861), .CK(clk), .Q(\mem[780][5] ) );
  DFF_X1 \mem_reg[780][4]  ( .D(n19862), .CK(clk), .Q(\mem[780][4] ) );
  DFF_X1 \mem_reg[780][3]  ( .D(n19863), .CK(clk), .Q(\mem[780][3] ) );
  DFF_X1 \mem_reg[780][2]  ( .D(n19864), .CK(clk), .Q(\mem[780][2] ) );
  DFF_X1 \mem_reg[780][1]  ( .D(n19865), .CK(clk), .Q(\mem[780][1] ) );
  DFF_X1 \mem_reg[780][0]  ( .D(n19866), .CK(clk), .Q(\mem[780][0] ) );
  DFF_X1 \mem_reg[779][7]  ( .D(n19867), .CK(clk), .Q(\mem[779][7] ) );
  DFF_X1 \mem_reg[779][6]  ( .D(n19868), .CK(clk), .Q(\mem[779][6] ) );
  DFF_X1 \mem_reg[779][5]  ( .D(n19869), .CK(clk), .Q(\mem[779][5] ) );
  DFF_X1 \mem_reg[779][4]  ( .D(n19870), .CK(clk), .Q(\mem[779][4] ) );
  DFF_X1 \mem_reg[779][3]  ( .D(n19871), .CK(clk), .Q(\mem[779][3] ) );
  DFF_X1 \mem_reg[779][2]  ( .D(n19872), .CK(clk), .Q(\mem[779][2] ) );
  DFF_X1 \mem_reg[779][1]  ( .D(n19873), .CK(clk), .Q(\mem[779][1] ) );
  DFF_X1 \mem_reg[779][0]  ( .D(n19874), .CK(clk), .Q(\mem[779][0] ) );
  DFF_X1 \mem_reg[778][7]  ( .D(n19875), .CK(clk), .Q(\mem[778][7] ) );
  DFF_X1 \mem_reg[778][6]  ( .D(n19876), .CK(clk), .Q(\mem[778][6] ) );
  DFF_X1 \mem_reg[778][5]  ( .D(n19877), .CK(clk), .Q(\mem[778][5] ) );
  DFF_X1 \mem_reg[778][4]  ( .D(n19878), .CK(clk), .Q(\mem[778][4] ) );
  DFF_X1 \mem_reg[778][3]  ( .D(n19879), .CK(clk), .Q(\mem[778][3] ) );
  DFF_X1 \mem_reg[778][2]  ( .D(n19880), .CK(clk), .Q(\mem[778][2] ) );
  DFF_X1 \mem_reg[778][1]  ( .D(n19881), .CK(clk), .Q(\mem[778][1] ) );
  DFF_X1 \mem_reg[778][0]  ( .D(n19882), .CK(clk), .Q(\mem[778][0] ) );
  DFF_X1 \mem_reg[777][7]  ( .D(n19883), .CK(clk), .Q(\mem[777][7] ) );
  DFF_X1 \mem_reg[777][6]  ( .D(n19884), .CK(clk), .Q(\mem[777][6] ) );
  DFF_X1 \mem_reg[777][5]  ( .D(n19885), .CK(clk), .Q(\mem[777][5] ) );
  DFF_X1 \mem_reg[777][4]  ( .D(n19886), .CK(clk), .Q(\mem[777][4] ) );
  DFF_X1 \mem_reg[777][3]  ( .D(n19887), .CK(clk), .Q(\mem[777][3] ) );
  DFF_X1 \mem_reg[777][2]  ( .D(n19888), .CK(clk), .Q(\mem[777][2] ) );
  DFF_X1 \mem_reg[777][1]  ( .D(n19889), .CK(clk), .Q(\mem[777][1] ) );
  DFF_X1 \mem_reg[777][0]  ( .D(n19890), .CK(clk), .Q(\mem[777][0] ) );
  DFF_X1 \mem_reg[776][7]  ( .D(n19891), .CK(clk), .Q(\mem[776][7] ) );
  DFF_X1 \mem_reg[776][6]  ( .D(n19892), .CK(clk), .Q(\mem[776][6] ) );
  DFF_X1 \mem_reg[776][5]  ( .D(n19893), .CK(clk), .Q(\mem[776][5] ) );
  DFF_X1 \mem_reg[776][4]  ( .D(n19894), .CK(clk), .Q(\mem[776][4] ) );
  DFF_X1 \mem_reg[776][3]  ( .D(n19895), .CK(clk), .Q(\mem[776][3] ) );
  DFF_X1 \mem_reg[776][2]  ( .D(n19896), .CK(clk), .Q(\mem[776][2] ) );
  DFF_X1 \mem_reg[776][1]  ( .D(n19897), .CK(clk), .Q(\mem[776][1] ) );
  DFF_X1 \mem_reg[776][0]  ( .D(n19898), .CK(clk), .Q(\mem[776][0] ) );
  DFF_X1 \mem_reg[775][7]  ( .D(n19899), .CK(clk), .Q(\mem[775][7] ) );
  DFF_X1 \mem_reg[775][6]  ( .D(n19900), .CK(clk), .Q(\mem[775][6] ) );
  DFF_X1 \mem_reg[775][5]  ( .D(n19901), .CK(clk), .Q(\mem[775][5] ) );
  DFF_X1 \mem_reg[775][4]  ( .D(n19902), .CK(clk), .Q(\mem[775][4] ) );
  DFF_X1 \mem_reg[775][3]  ( .D(n19903), .CK(clk), .Q(\mem[775][3] ) );
  DFF_X1 \mem_reg[775][2]  ( .D(n19904), .CK(clk), .Q(\mem[775][2] ) );
  DFF_X1 \mem_reg[775][1]  ( .D(n19905), .CK(clk), .Q(\mem[775][1] ) );
  DFF_X1 \mem_reg[775][0]  ( .D(n19906), .CK(clk), .Q(\mem[775][0] ) );
  DFF_X1 \mem_reg[774][7]  ( .D(n19907), .CK(clk), .Q(\mem[774][7] ) );
  DFF_X1 \mem_reg[774][6]  ( .D(n19908), .CK(clk), .Q(\mem[774][6] ) );
  DFF_X1 \mem_reg[774][5]  ( .D(n19909), .CK(clk), .Q(\mem[774][5] ) );
  DFF_X1 \mem_reg[774][4]  ( .D(n19910), .CK(clk), .Q(\mem[774][4] ) );
  DFF_X1 \mem_reg[774][3]  ( .D(n19911), .CK(clk), .Q(\mem[774][3] ) );
  DFF_X1 \mem_reg[774][2]  ( .D(n19912), .CK(clk), .Q(\mem[774][2] ) );
  DFF_X1 \mem_reg[774][1]  ( .D(n19913), .CK(clk), .Q(\mem[774][1] ) );
  DFF_X1 \mem_reg[774][0]  ( .D(n19914), .CK(clk), .Q(\mem[774][0] ) );
  DFF_X1 \mem_reg[773][7]  ( .D(n19915), .CK(clk), .Q(\mem[773][7] ) );
  DFF_X1 \mem_reg[773][6]  ( .D(n19916), .CK(clk), .Q(\mem[773][6] ) );
  DFF_X1 \mem_reg[773][5]  ( .D(n19917), .CK(clk), .Q(\mem[773][5] ) );
  DFF_X1 \mem_reg[773][4]  ( .D(n19918), .CK(clk), .Q(\mem[773][4] ) );
  DFF_X1 \mem_reg[773][3]  ( .D(n19919), .CK(clk), .Q(\mem[773][3] ) );
  DFF_X1 \mem_reg[773][2]  ( .D(n19920), .CK(clk), .Q(\mem[773][2] ) );
  DFF_X1 \mem_reg[773][1]  ( .D(n19921), .CK(clk), .Q(\mem[773][1] ) );
  DFF_X1 \mem_reg[773][0]  ( .D(n19922), .CK(clk), .Q(\mem[773][0] ) );
  DFF_X1 \mem_reg[772][7]  ( .D(n19923), .CK(clk), .Q(\mem[772][7] ) );
  DFF_X1 \mem_reg[772][6]  ( .D(n19924), .CK(clk), .Q(\mem[772][6] ) );
  DFF_X1 \mem_reg[772][5]  ( .D(n19925), .CK(clk), .Q(\mem[772][5] ) );
  DFF_X1 \mem_reg[772][4]  ( .D(n19926), .CK(clk), .Q(\mem[772][4] ) );
  DFF_X1 \mem_reg[772][3]  ( .D(n19927), .CK(clk), .Q(\mem[772][3] ) );
  DFF_X1 \mem_reg[772][2]  ( .D(n19928), .CK(clk), .Q(\mem[772][2] ) );
  DFF_X1 \mem_reg[772][1]  ( .D(n19929), .CK(clk), .Q(\mem[772][1] ) );
  DFF_X1 \mem_reg[772][0]  ( .D(n19930), .CK(clk), .Q(\mem[772][0] ) );
  DFF_X1 \mem_reg[771][7]  ( .D(n19931), .CK(clk), .Q(\mem[771][7] ) );
  DFF_X1 \mem_reg[771][6]  ( .D(n19932), .CK(clk), .Q(\mem[771][6] ) );
  DFF_X1 \mem_reg[771][5]  ( .D(n19933), .CK(clk), .Q(\mem[771][5] ) );
  DFF_X1 \mem_reg[771][4]  ( .D(n19934), .CK(clk), .Q(\mem[771][4] ) );
  DFF_X1 \mem_reg[771][3]  ( .D(n19935), .CK(clk), .Q(\mem[771][3] ) );
  DFF_X1 \mem_reg[771][2]  ( .D(n19936), .CK(clk), .Q(\mem[771][2] ) );
  DFF_X1 \mem_reg[771][1]  ( .D(n19937), .CK(clk), .Q(\mem[771][1] ) );
  DFF_X1 \mem_reg[771][0]  ( .D(n19938), .CK(clk), .Q(\mem[771][0] ) );
  DFF_X1 \mem_reg[770][7]  ( .D(n19939), .CK(clk), .Q(\mem[770][7] ) );
  DFF_X1 \mem_reg[770][6]  ( .D(n19940), .CK(clk), .Q(\mem[770][6] ) );
  DFF_X1 \mem_reg[770][5]  ( .D(n19941), .CK(clk), .Q(\mem[770][5] ) );
  DFF_X1 \mem_reg[770][4]  ( .D(n19942), .CK(clk), .Q(\mem[770][4] ) );
  DFF_X1 \mem_reg[770][3]  ( .D(n19943), .CK(clk), .Q(\mem[770][3] ) );
  DFF_X1 \mem_reg[770][2]  ( .D(n19944), .CK(clk), .Q(\mem[770][2] ) );
  DFF_X1 \mem_reg[770][1]  ( .D(n19945), .CK(clk), .Q(\mem[770][1] ) );
  DFF_X1 \mem_reg[770][0]  ( .D(n19946), .CK(clk), .Q(\mem[770][0] ) );
  DFF_X1 \mem_reg[769][7]  ( .D(n19947), .CK(clk), .Q(\mem[769][7] ) );
  DFF_X1 \mem_reg[769][6]  ( .D(n19948), .CK(clk), .Q(\mem[769][6] ) );
  DFF_X1 \mem_reg[769][5]  ( .D(n19949), .CK(clk), .Q(\mem[769][5] ) );
  DFF_X1 \mem_reg[769][4]  ( .D(n19950), .CK(clk), .Q(\mem[769][4] ) );
  DFF_X1 \mem_reg[769][3]  ( .D(n19951), .CK(clk), .Q(\mem[769][3] ) );
  DFF_X1 \mem_reg[769][2]  ( .D(n19952), .CK(clk), .Q(\mem[769][2] ) );
  DFF_X1 \mem_reg[769][1]  ( .D(n19953), .CK(clk), .Q(\mem[769][1] ) );
  DFF_X1 \mem_reg[769][0]  ( .D(n19954), .CK(clk), .Q(\mem[769][0] ) );
  DFF_X1 \mem_reg[768][7]  ( .D(n19955), .CK(clk), .Q(\mem[768][7] ) );
  DFF_X1 \mem_reg[768][6]  ( .D(n19956), .CK(clk), .Q(\mem[768][6] ) );
  DFF_X1 \mem_reg[768][5]  ( .D(n19957), .CK(clk), .Q(\mem[768][5] ) );
  DFF_X1 \mem_reg[768][4]  ( .D(n19958), .CK(clk), .Q(\mem[768][4] ) );
  DFF_X1 \mem_reg[768][3]  ( .D(n19959), .CK(clk), .Q(\mem[768][3] ) );
  DFF_X1 \mem_reg[768][2]  ( .D(n19960), .CK(clk), .Q(\mem[768][2] ) );
  DFF_X1 \mem_reg[768][1]  ( .D(n19961), .CK(clk), .Q(\mem[768][1] ) );
  DFF_X1 \mem_reg[768][0]  ( .D(n19962), .CK(clk), .Q(\mem[768][0] ) );
  DFF_X1 \mem_reg[767][7]  ( .D(n19963), .CK(clk), .Q(\mem[767][7] ) );
  DFF_X1 \mem_reg[767][6]  ( .D(n19964), .CK(clk), .Q(\mem[767][6] ) );
  DFF_X1 \mem_reg[767][5]  ( .D(n19965), .CK(clk), .Q(\mem[767][5] ) );
  DFF_X1 \mem_reg[767][4]  ( .D(n19966), .CK(clk), .Q(\mem[767][4] ) );
  DFF_X1 \mem_reg[767][3]  ( .D(n19967), .CK(clk), .Q(\mem[767][3] ) );
  DFF_X1 \mem_reg[767][2]  ( .D(n19968), .CK(clk), .Q(\mem[767][2] ) );
  DFF_X1 \mem_reg[767][1]  ( .D(n19969), .CK(clk), .Q(\mem[767][1] ) );
  DFF_X1 \mem_reg[767][0]  ( .D(n19970), .CK(clk), .Q(\mem[767][0] ) );
  DFF_X1 \mem_reg[766][7]  ( .D(n19971), .CK(clk), .Q(\mem[766][7] ) );
  DFF_X1 \mem_reg[766][6]  ( .D(n19972), .CK(clk), .Q(\mem[766][6] ) );
  DFF_X1 \mem_reg[766][5]  ( .D(n19973), .CK(clk), .Q(\mem[766][5] ) );
  DFF_X1 \mem_reg[766][4]  ( .D(n19974), .CK(clk), .Q(\mem[766][4] ) );
  DFF_X1 \mem_reg[766][3]  ( .D(n19975), .CK(clk), .Q(\mem[766][3] ) );
  DFF_X1 \mem_reg[766][2]  ( .D(n19976), .CK(clk), .Q(\mem[766][2] ) );
  DFF_X1 \mem_reg[766][1]  ( .D(n19977), .CK(clk), .Q(\mem[766][1] ) );
  DFF_X1 \mem_reg[766][0]  ( .D(n19978), .CK(clk), .Q(\mem[766][0] ) );
  DFF_X1 \mem_reg[765][7]  ( .D(n19979), .CK(clk), .Q(\mem[765][7] ) );
  DFF_X1 \mem_reg[765][6]  ( .D(n19980), .CK(clk), .Q(\mem[765][6] ) );
  DFF_X1 \mem_reg[765][5]  ( .D(n19981), .CK(clk), .Q(\mem[765][5] ) );
  DFF_X1 \mem_reg[765][4]  ( .D(n19982), .CK(clk), .Q(\mem[765][4] ) );
  DFF_X1 \mem_reg[765][3]  ( .D(n19983), .CK(clk), .Q(\mem[765][3] ) );
  DFF_X1 \mem_reg[765][2]  ( .D(n19984), .CK(clk), .Q(\mem[765][2] ) );
  DFF_X1 \mem_reg[765][1]  ( .D(n19985), .CK(clk), .Q(\mem[765][1] ) );
  DFF_X1 \mem_reg[765][0]  ( .D(n19986), .CK(clk), .Q(\mem[765][0] ) );
  DFF_X1 \mem_reg[764][7]  ( .D(n19987), .CK(clk), .Q(\mem[764][7] ) );
  DFF_X1 \mem_reg[764][6]  ( .D(n19988), .CK(clk), .Q(\mem[764][6] ) );
  DFF_X1 \mem_reg[764][5]  ( .D(n19989), .CK(clk), .Q(\mem[764][5] ) );
  DFF_X1 \mem_reg[764][4]  ( .D(n19990), .CK(clk), .Q(\mem[764][4] ) );
  DFF_X1 \mem_reg[764][3]  ( .D(n19991), .CK(clk), .Q(\mem[764][3] ) );
  DFF_X1 \mem_reg[764][2]  ( .D(n19992), .CK(clk), .Q(\mem[764][2] ) );
  DFF_X1 \mem_reg[764][1]  ( .D(n19993), .CK(clk), .Q(\mem[764][1] ) );
  DFF_X1 \mem_reg[764][0]  ( .D(n19994), .CK(clk), .Q(\mem[764][0] ) );
  DFF_X1 \mem_reg[763][7]  ( .D(n19995), .CK(clk), .Q(\mem[763][7] ) );
  DFF_X1 \mem_reg[763][6]  ( .D(n19996), .CK(clk), .Q(\mem[763][6] ) );
  DFF_X1 \mem_reg[763][5]  ( .D(n19997), .CK(clk), .Q(\mem[763][5] ) );
  DFF_X1 \mem_reg[763][4]  ( .D(n19998), .CK(clk), .Q(\mem[763][4] ) );
  DFF_X1 \mem_reg[763][3]  ( .D(n19999), .CK(clk), .Q(\mem[763][3] ) );
  DFF_X1 \mem_reg[763][2]  ( .D(n20000), .CK(clk), .Q(\mem[763][2] ) );
  DFF_X1 \mem_reg[763][1]  ( .D(n20001), .CK(clk), .Q(\mem[763][1] ) );
  DFF_X1 \mem_reg[763][0]  ( .D(n20002), .CK(clk), .Q(\mem[763][0] ) );
  DFF_X1 \mem_reg[762][7]  ( .D(n20003), .CK(clk), .Q(\mem[762][7] ) );
  DFF_X1 \mem_reg[762][6]  ( .D(n20004), .CK(clk), .Q(\mem[762][6] ) );
  DFF_X1 \mem_reg[762][5]  ( .D(n20005), .CK(clk), .Q(\mem[762][5] ) );
  DFF_X1 \mem_reg[762][4]  ( .D(n20006), .CK(clk), .Q(\mem[762][4] ) );
  DFF_X1 \mem_reg[762][3]  ( .D(n20007), .CK(clk), .Q(\mem[762][3] ) );
  DFF_X1 \mem_reg[762][2]  ( .D(n20008), .CK(clk), .Q(\mem[762][2] ) );
  DFF_X1 \mem_reg[762][1]  ( .D(n20009), .CK(clk), .Q(\mem[762][1] ) );
  DFF_X1 \mem_reg[762][0]  ( .D(n20010), .CK(clk), .Q(\mem[762][0] ) );
  DFF_X1 \mem_reg[761][7]  ( .D(n20011), .CK(clk), .Q(\mem[761][7] ) );
  DFF_X1 \mem_reg[761][6]  ( .D(n20012), .CK(clk), .Q(\mem[761][6] ) );
  DFF_X1 \mem_reg[761][5]  ( .D(n20013), .CK(clk), .Q(\mem[761][5] ) );
  DFF_X1 \mem_reg[761][4]  ( .D(n20014), .CK(clk), .Q(\mem[761][4] ) );
  DFF_X1 \mem_reg[761][3]  ( .D(n20015), .CK(clk), .Q(\mem[761][3] ) );
  DFF_X1 \mem_reg[761][2]  ( .D(n20016), .CK(clk), .Q(\mem[761][2] ) );
  DFF_X1 \mem_reg[761][1]  ( .D(n20017), .CK(clk), .Q(\mem[761][1] ) );
  DFF_X1 \mem_reg[761][0]  ( .D(n20018), .CK(clk), .Q(\mem[761][0] ) );
  DFF_X1 \mem_reg[760][7]  ( .D(n20019), .CK(clk), .Q(\mem[760][7] ) );
  DFF_X1 \mem_reg[760][6]  ( .D(n20020), .CK(clk), .Q(\mem[760][6] ) );
  DFF_X1 \mem_reg[760][5]  ( .D(n20021), .CK(clk), .Q(\mem[760][5] ) );
  DFF_X1 \mem_reg[760][4]  ( .D(n20022), .CK(clk), .Q(\mem[760][4] ) );
  DFF_X1 \mem_reg[760][3]  ( .D(n20023), .CK(clk), .Q(\mem[760][3] ) );
  DFF_X1 \mem_reg[760][2]  ( .D(n20024), .CK(clk), .Q(\mem[760][2] ) );
  DFF_X1 \mem_reg[760][1]  ( .D(n20025), .CK(clk), .Q(\mem[760][1] ) );
  DFF_X1 \mem_reg[760][0]  ( .D(n20026), .CK(clk), .Q(\mem[760][0] ) );
  DFF_X1 \mem_reg[759][7]  ( .D(n20027), .CK(clk), .Q(\mem[759][7] ) );
  DFF_X1 \mem_reg[759][6]  ( .D(n20028), .CK(clk), .Q(\mem[759][6] ) );
  DFF_X1 \mem_reg[759][5]  ( .D(n20029), .CK(clk), .Q(\mem[759][5] ) );
  DFF_X1 \mem_reg[759][4]  ( .D(n20030), .CK(clk), .Q(\mem[759][4] ) );
  DFF_X1 \mem_reg[759][3]  ( .D(n20031), .CK(clk), .Q(\mem[759][3] ) );
  DFF_X1 \mem_reg[759][2]  ( .D(n20032), .CK(clk), .Q(\mem[759][2] ) );
  DFF_X1 \mem_reg[759][1]  ( .D(n20033), .CK(clk), .Q(\mem[759][1] ) );
  DFF_X1 \mem_reg[759][0]  ( .D(n20034), .CK(clk), .Q(\mem[759][0] ) );
  DFF_X1 \mem_reg[758][7]  ( .D(n20035), .CK(clk), .Q(\mem[758][7] ) );
  DFF_X1 \mem_reg[758][6]  ( .D(n20036), .CK(clk), .Q(\mem[758][6] ) );
  DFF_X1 \mem_reg[758][5]  ( .D(n20037), .CK(clk), .Q(\mem[758][5] ) );
  DFF_X1 \mem_reg[758][4]  ( .D(n20038), .CK(clk), .Q(\mem[758][4] ) );
  DFF_X1 \mem_reg[758][3]  ( .D(n20039), .CK(clk), .Q(\mem[758][3] ) );
  DFF_X1 \mem_reg[758][2]  ( .D(n20040), .CK(clk), .Q(\mem[758][2] ) );
  DFF_X1 \mem_reg[758][1]  ( .D(n20041), .CK(clk), .Q(\mem[758][1] ) );
  DFF_X1 \mem_reg[758][0]  ( .D(n20042), .CK(clk), .Q(\mem[758][0] ) );
  DFF_X1 \mem_reg[757][7]  ( .D(n20043), .CK(clk), .Q(\mem[757][7] ) );
  DFF_X1 \mem_reg[757][6]  ( .D(n20044), .CK(clk), .Q(\mem[757][6] ) );
  DFF_X1 \mem_reg[757][5]  ( .D(n20045), .CK(clk), .Q(\mem[757][5] ) );
  DFF_X1 \mem_reg[757][4]  ( .D(n20046), .CK(clk), .Q(\mem[757][4] ) );
  DFF_X1 \mem_reg[757][3]  ( .D(n20047), .CK(clk), .Q(\mem[757][3] ) );
  DFF_X1 \mem_reg[757][2]  ( .D(n20048), .CK(clk), .Q(\mem[757][2] ) );
  DFF_X1 \mem_reg[757][1]  ( .D(n20049), .CK(clk), .Q(\mem[757][1] ) );
  DFF_X1 \mem_reg[757][0]  ( .D(n20050), .CK(clk), .Q(\mem[757][0] ) );
  DFF_X1 \mem_reg[756][7]  ( .D(n20051), .CK(clk), .Q(\mem[756][7] ) );
  DFF_X1 \mem_reg[756][6]  ( .D(n20052), .CK(clk), .Q(\mem[756][6] ) );
  DFF_X1 \mem_reg[756][5]  ( .D(n20053), .CK(clk), .Q(\mem[756][5] ) );
  DFF_X1 \mem_reg[756][4]  ( .D(n20054), .CK(clk), .Q(\mem[756][4] ) );
  DFF_X1 \mem_reg[756][3]  ( .D(n20055), .CK(clk), .Q(\mem[756][3] ) );
  DFF_X1 \mem_reg[756][2]  ( .D(n20056), .CK(clk), .Q(\mem[756][2] ) );
  DFF_X1 \mem_reg[756][1]  ( .D(n20057), .CK(clk), .Q(\mem[756][1] ) );
  DFF_X1 \mem_reg[756][0]  ( .D(n20058), .CK(clk), .Q(\mem[756][0] ) );
  DFF_X1 \mem_reg[755][7]  ( .D(n20059), .CK(clk), .Q(\mem[755][7] ) );
  DFF_X1 \mem_reg[755][6]  ( .D(n20060), .CK(clk), .Q(\mem[755][6] ) );
  DFF_X1 \mem_reg[755][5]  ( .D(n20061), .CK(clk), .Q(\mem[755][5] ) );
  DFF_X1 \mem_reg[755][4]  ( .D(n20062), .CK(clk), .Q(\mem[755][4] ) );
  DFF_X1 \mem_reg[755][3]  ( .D(n20063), .CK(clk), .Q(\mem[755][3] ) );
  DFF_X1 \mem_reg[755][2]  ( .D(n20064), .CK(clk), .Q(\mem[755][2] ) );
  DFF_X1 \mem_reg[755][1]  ( .D(n20065), .CK(clk), .Q(\mem[755][1] ) );
  DFF_X1 \mem_reg[755][0]  ( .D(n20066), .CK(clk), .Q(\mem[755][0] ) );
  DFF_X1 \mem_reg[754][7]  ( .D(n20067), .CK(clk), .Q(\mem[754][7] ) );
  DFF_X1 \mem_reg[754][6]  ( .D(n20068), .CK(clk), .Q(\mem[754][6] ) );
  DFF_X1 \mem_reg[754][5]  ( .D(n20069), .CK(clk), .Q(\mem[754][5] ) );
  DFF_X1 \mem_reg[754][4]  ( .D(n20070), .CK(clk), .Q(\mem[754][4] ) );
  DFF_X1 \mem_reg[754][3]  ( .D(n20071), .CK(clk), .Q(\mem[754][3] ) );
  DFF_X1 \mem_reg[754][2]  ( .D(n20072), .CK(clk), .Q(\mem[754][2] ) );
  DFF_X1 \mem_reg[754][1]  ( .D(n20073), .CK(clk), .Q(\mem[754][1] ) );
  DFF_X1 \mem_reg[754][0]  ( .D(n20074), .CK(clk), .Q(\mem[754][0] ) );
  DFF_X1 \mem_reg[753][7]  ( .D(n20075), .CK(clk), .Q(\mem[753][7] ) );
  DFF_X1 \mem_reg[753][6]  ( .D(n20076), .CK(clk), .Q(\mem[753][6] ) );
  DFF_X1 \mem_reg[753][5]  ( .D(n20077), .CK(clk), .Q(\mem[753][5] ) );
  DFF_X1 \mem_reg[753][4]  ( .D(n20078), .CK(clk), .Q(\mem[753][4] ) );
  DFF_X1 \mem_reg[753][3]  ( .D(n20079), .CK(clk), .Q(\mem[753][3] ) );
  DFF_X1 \mem_reg[753][2]  ( .D(n20080), .CK(clk), .Q(\mem[753][2] ) );
  DFF_X1 \mem_reg[753][1]  ( .D(n20081), .CK(clk), .Q(\mem[753][1] ) );
  DFF_X1 \mem_reg[753][0]  ( .D(n20082), .CK(clk), .Q(\mem[753][0] ) );
  DFF_X1 \mem_reg[752][7]  ( .D(n20083), .CK(clk), .Q(\mem[752][7] ) );
  DFF_X1 \mem_reg[752][6]  ( .D(n20084), .CK(clk), .Q(\mem[752][6] ) );
  DFF_X1 \mem_reg[752][5]  ( .D(n20085), .CK(clk), .Q(\mem[752][5] ) );
  DFF_X1 \mem_reg[752][4]  ( .D(n20086), .CK(clk), .Q(\mem[752][4] ) );
  DFF_X1 \mem_reg[752][3]  ( .D(n20087), .CK(clk), .Q(\mem[752][3] ) );
  DFF_X1 \mem_reg[752][2]  ( .D(n20088), .CK(clk), .Q(\mem[752][2] ) );
  DFF_X1 \mem_reg[752][1]  ( .D(n20089), .CK(clk), .Q(\mem[752][1] ) );
  DFF_X1 \mem_reg[752][0]  ( .D(n20090), .CK(clk), .Q(\mem[752][0] ) );
  DFF_X1 \mem_reg[751][7]  ( .D(n20091), .CK(clk), .Q(\mem[751][7] ) );
  DFF_X1 \mem_reg[751][6]  ( .D(n20092), .CK(clk), .Q(\mem[751][6] ) );
  DFF_X1 \mem_reg[751][5]  ( .D(n20093), .CK(clk), .Q(\mem[751][5] ) );
  DFF_X1 \mem_reg[751][4]  ( .D(n20094), .CK(clk), .Q(\mem[751][4] ) );
  DFF_X1 \mem_reg[751][3]  ( .D(n20095), .CK(clk), .Q(\mem[751][3] ) );
  DFF_X1 \mem_reg[751][2]  ( .D(n20096), .CK(clk), .Q(\mem[751][2] ) );
  DFF_X1 \mem_reg[751][1]  ( .D(n20097), .CK(clk), .Q(\mem[751][1] ) );
  DFF_X1 \mem_reg[751][0]  ( .D(n20098), .CK(clk), .Q(\mem[751][0] ) );
  DFF_X1 \mem_reg[750][7]  ( .D(n20099), .CK(clk), .Q(\mem[750][7] ) );
  DFF_X1 \mem_reg[750][6]  ( .D(n20100), .CK(clk), .Q(\mem[750][6] ) );
  DFF_X1 \mem_reg[750][5]  ( .D(n20101), .CK(clk), .Q(\mem[750][5] ) );
  DFF_X1 \mem_reg[750][4]  ( .D(n20102), .CK(clk), .Q(\mem[750][4] ) );
  DFF_X1 \mem_reg[750][3]  ( .D(n20103), .CK(clk), .Q(\mem[750][3] ) );
  DFF_X1 \mem_reg[750][2]  ( .D(n20104), .CK(clk), .Q(\mem[750][2] ) );
  DFF_X1 \mem_reg[750][1]  ( .D(n20105), .CK(clk), .Q(\mem[750][1] ) );
  DFF_X1 \mem_reg[750][0]  ( .D(n20106), .CK(clk), .Q(\mem[750][0] ) );
  DFF_X1 \mem_reg[749][7]  ( .D(n20107), .CK(clk), .Q(\mem[749][7] ) );
  DFF_X1 \mem_reg[749][6]  ( .D(n20108), .CK(clk), .Q(\mem[749][6] ) );
  DFF_X1 \mem_reg[749][5]  ( .D(n20109), .CK(clk), .Q(\mem[749][5] ) );
  DFF_X1 \mem_reg[749][4]  ( .D(n20110), .CK(clk), .Q(\mem[749][4] ) );
  DFF_X1 \mem_reg[749][3]  ( .D(n20111), .CK(clk), .Q(\mem[749][3] ) );
  DFF_X1 \mem_reg[749][2]  ( .D(n20112), .CK(clk), .Q(\mem[749][2] ) );
  DFF_X1 \mem_reg[749][1]  ( .D(n20113), .CK(clk), .Q(\mem[749][1] ) );
  DFF_X1 \mem_reg[749][0]  ( .D(n20114), .CK(clk), .Q(\mem[749][0] ) );
  DFF_X1 \mem_reg[748][7]  ( .D(n20115), .CK(clk), .Q(\mem[748][7] ) );
  DFF_X1 \mem_reg[748][6]  ( .D(n20116), .CK(clk), .Q(\mem[748][6] ) );
  DFF_X1 \mem_reg[748][5]  ( .D(n20117), .CK(clk), .Q(\mem[748][5] ) );
  DFF_X1 \mem_reg[748][4]  ( .D(n20118), .CK(clk), .Q(\mem[748][4] ) );
  DFF_X1 \mem_reg[748][3]  ( .D(n20119), .CK(clk), .Q(\mem[748][3] ) );
  DFF_X1 \mem_reg[748][2]  ( .D(n20120), .CK(clk), .Q(\mem[748][2] ) );
  DFF_X1 \mem_reg[748][1]  ( .D(n20121), .CK(clk), .Q(\mem[748][1] ) );
  DFF_X1 \mem_reg[748][0]  ( .D(n20122), .CK(clk), .Q(\mem[748][0] ) );
  DFF_X1 \mem_reg[747][7]  ( .D(n20123), .CK(clk), .Q(\mem[747][7] ) );
  DFF_X1 \mem_reg[747][6]  ( .D(n20124), .CK(clk), .Q(\mem[747][6] ) );
  DFF_X1 \mem_reg[747][5]  ( .D(n20125), .CK(clk), .Q(\mem[747][5] ) );
  DFF_X1 \mem_reg[747][4]  ( .D(n20126), .CK(clk), .Q(\mem[747][4] ) );
  DFF_X1 \mem_reg[747][3]  ( .D(n20127), .CK(clk), .Q(\mem[747][3] ) );
  DFF_X1 \mem_reg[747][2]  ( .D(n20128), .CK(clk), .Q(\mem[747][2] ) );
  DFF_X1 \mem_reg[747][1]  ( .D(n20129), .CK(clk), .Q(\mem[747][1] ) );
  DFF_X1 \mem_reg[747][0]  ( .D(n20130), .CK(clk), .Q(\mem[747][0] ) );
  DFF_X1 \mem_reg[746][7]  ( .D(n20131), .CK(clk), .Q(\mem[746][7] ) );
  DFF_X1 \mem_reg[746][6]  ( .D(n20132), .CK(clk), .Q(\mem[746][6] ) );
  DFF_X1 \mem_reg[746][5]  ( .D(n20133), .CK(clk), .Q(\mem[746][5] ) );
  DFF_X1 \mem_reg[746][4]  ( .D(n20134), .CK(clk), .Q(\mem[746][4] ) );
  DFF_X1 \mem_reg[746][3]  ( .D(n20135), .CK(clk), .Q(\mem[746][3] ) );
  DFF_X1 \mem_reg[746][2]  ( .D(n20136), .CK(clk), .Q(\mem[746][2] ) );
  DFF_X1 \mem_reg[746][1]  ( .D(n20137), .CK(clk), .Q(\mem[746][1] ) );
  DFF_X1 \mem_reg[746][0]  ( .D(n20138), .CK(clk), .Q(\mem[746][0] ) );
  DFF_X1 \mem_reg[745][7]  ( .D(n20139), .CK(clk), .Q(\mem[745][7] ) );
  DFF_X1 \mem_reg[745][6]  ( .D(n20140), .CK(clk), .Q(\mem[745][6] ) );
  DFF_X1 \mem_reg[745][5]  ( .D(n20141), .CK(clk), .Q(\mem[745][5] ) );
  DFF_X1 \mem_reg[745][4]  ( .D(n20142), .CK(clk), .Q(\mem[745][4] ) );
  DFF_X1 \mem_reg[745][3]  ( .D(n20143), .CK(clk), .Q(\mem[745][3] ) );
  DFF_X1 \mem_reg[745][2]  ( .D(n20144), .CK(clk), .Q(\mem[745][2] ) );
  DFF_X1 \mem_reg[745][1]  ( .D(n20145), .CK(clk), .Q(\mem[745][1] ) );
  DFF_X1 \mem_reg[745][0]  ( .D(n20146), .CK(clk), .Q(\mem[745][0] ) );
  DFF_X1 \mem_reg[744][7]  ( .D(n20147), .CK(clk), .Q(\mem[744][7] ) );
  DFF_X1 \mem_reg[744][6]  ( .D(n20148), .CK(clk), .Q(\mem[744][6] ) );
  DFF_X1 \mem_reg[744][5]  ( .D(n20149), .CK(clk), .Q(\mem[744][5] ) );
  DFF_X1 \mem_reg[744][4]  ( .D(n20150), .CK(clk), .Q(\mem[744][4] ) );
  DFF_X1 \mem_reg[744][3]  ( .D(n20151), .CK(clk), .Q(\mem[744][3] ) );
  DFF_X1 \mem_reg[744][2]  ( .D(n20152), .CK(clk), .Q(\mem[744][2] ) );
  DFF_X1 \mem_reg[744][1]  ( .D(n20153), .CK(clk), .Q(\mem[744][1] ) );
  DFF_X1 \mem_reg[744][0]  ( .D(n20154), .CK(clk), .Q(\mem[744][0] ) );
  DFF_X1 \mem_reg[743][7]  ( .D(n20155), .CK(clk), .Q(\mem[743][7] ) );
  DFF_X1 \mem_reg[743][6]  ( .D(n20156), .CK(clk), .Q(\mem[743][6] ) );
  DFF_X1 \mem_reg[743][5]  ( .D(n20157), .CK(clk), .Q(\mem[743][5] ) );
  DFF_X1 \mem_reg[743][4]  ( .D(n20158), .CK(clk), .Q(\mem[743][4] ) );
  DFF_X1 \mem_reg[743][3]  ( .D(n20159), .CK(clk), .Q(\mem[743][3] ) );
  DFF_X1 \mem_reg[743][2]  ( .D(n20160), .CK(clk), .Q(\mem[743][2] ) );
  DFF_X1 \mem_reg[743][1]  ( .D(n20161), .CK(clk), .Q(\mem[743][1] ) );
  DFF_X1 \mem_reg[743][0]  ( .D(n20162), .CK(clk), .Q(\mem[743][0] ) );
  DFF_X1 \mem_reg[742][7]  ( .D(n20163), .CK(clk), .Q(\mem[742][7] ) );
  DFF_X1 \mem_reg[742][6]  ( .D(n20164), .CK(clk), .Q(\mem[742][6] ) );
  DFF_X1 \mem_reg[742][5]  ( .D(n20165), .CK(clk), .Q(\mem[742][5] ) );
  DFF_X1 \mem_reg[742][4]  ( .D(n20166), .CK(clk), .Q(\mem[742][4] ) );
  DFF_X1 \mem_reg[742][3]  ( .D(n20167), .CK(clk), .Q(\mem[742][3] ) );
  DFF_X1 \mem_reg[742][2]  ( .D(n20168), .CK(clk), .Q(\mem[742][2] ) );
  DFF_X1 \mem_reg[742][1]  ( .D(n20169), .CK(clk), .Q(\mem[742][1] ) );
  DFF_X1 \mem_reg[742][0]  ( .D(n20170), .CK(clk), .Q(\mem[742][0] ) );
  DFF_X1 \mem_reg[741][7]  ( .D(n20171), .CK(clk), .Q(\mem[741][7] ) );
  DFF_X1 \mem_reg[741][6]  ( .D(n20172), .CK(clk), .Q(\mem[741][6] ) );
  DFF_X1 \mem_reg[741][5]  ( .D(n20173), .CK(clk), .Q(\mem[741][5] ) );
  DFF_X1 \mem_reg[741][4]  ( .D(n20174), .CK(clk), .Q(\mem[741][4] ) );
  DFF_X1 \mem_reg[741][3]  ( .D(n20175), .CK(clk), .Q(\mem[741][3] ) );
  DFF_X1 \mem_reg[741][2]  ( .D(n20176), .CK(clk), .Q(\mem[741][2] ) );
  DFF_X1 \mem_reg[741][1]  ( .D(n20177), .CK(clk), .Q(\mem[741][1] ) );
  DFF_X1 \mem_reg[741][0]  ( .D(n20178), .CK(clk), .Q(\mem[741][0] ) );
  DFF_X1 \mem_reg[740][7]  ( .D(n20179), .CK(clk), .Q(\mem[740][7] ) );
  DFF_X1 \mem_reg[740][6]  ( .D(n20180), .CK(clk), .Q(\mem[740][6] ) );
  DFF_X1 \mem_reg[740][5]  ( .D(n20181), .CK(clk), .Q(\mem[740][5] ) );
  DFF_X1 \mem_reg[740][4]  ( .D(n20182), .CK(clk), .Q(\mem[740][4] ) );
  DFF_X1 \mem_reg[740][3]  ( .D(n20183), .CK(clk), .Q(\mem[740][3] ) );
  DFF_X1 \mem_reg[740][2]  ( .D(n20184), .CK(clk), .Q(\mem[740][2] ) );
  DFF_X1 \mem_reg[740][1]  ( .D(n20185), .CK(clk), .Q(\mem[740][1] ) );
  DFF_X1 \mem_reg[740][0]  ( .D(n20186), .CK(clk), .Q(\mem[740][0] ) );
  DFF_X1 \mem_reg[739][7]  ( .D(n20187), .CK(clk), .Q(\mem[739][7] ) );
  DFF_X1 \mem_reg[739][6]  ( .D(n20188), .CK(clk), .Q(\mem[739][6] ) );
  DFF_X1 \mem_reg[739][5]  ( .D(n20189), .CK(clk), .Q(\mem[739][5] ) );
  DFF_X1 \mem_reg[739][4]  ( .D(n20190), .CK(clk), .Q(\mem[739][4] ) );
  DFF_X1 \mem_reg[739][3]  ( .D(n20191), .CK(clk), .Q(\mem[739][3] ) );
  DFF_X1 \mem_reg[739][2]  ( .D(n20192), .CK(clk), .Q(\mem[739][2] ) );
  DFF_X1 \mem_reg[739][1]  ( .D(n20193), .CK(clk), .Q(\mem[739][1] ) );
  DFF_X1 \mem_reg[739][0]  ( .D(n20194), .CK(clk), .Q(\mem[739][0] ) );
  DFF_X1 \mem_reg[738][7]  ( .D(n20195), .CK(clk), .Q(\mem[738][7] ) );
  DFF_X1 \mem_reg[738][6]  ( .D(n20196), .CK(clk), .Q(\mem[738][6] ) );
  DFF_X1 \mem_reg[738][5]  ( .D(n20197), .CK(clk), .Q(\mem[738][5] ) );
  DFF_X1 \mem_reg[738][4]  ( .D(n20198), .CK(clk), .Q(\mem[738][4] ) );
  DFF_X1 \mem_reg[738][3]  ( .D(n20199), .CK(clk), .Q(\mem[738][3] ) );
  DFF_X1 \mem_reg[738][2]  ( .D(n20200), .CK(clk), .Q(\mem[738][2] ) );
  DFF_X1 \mem_reg[738][1]  ( .D(n20201), .CK(clk), .Q(\mem[738][1] ) );
  DFF_X1 \mem_reg[738][0]  ( .D(n20202), .CK(clk), .Q(\mem[738][0] ) );
  DFF_X1 \mem_reg[737][7]  ( .D(n20203), .CK(clk), .Q(\mem[737][7] ) );
  DFF_X1 \mem_reg[737][6]  ( .D(n20204), .CK(clk), .Q(\mem[737][6] ) );
  DFF_X1 \mem_reg[737][5]  ( .D(n20205), .CK(clk), .Q(\mem[737][5] ) );
  DFF_X1 \mem_reg[737][4]  ( .D(n20206), .CK(clk), .Q(\mem[737][4] ) );
  DFF_X1 \mem_reg[737][3]  ( .D(n20207), .CK(clk), .Q(\mem[737][3] ) );
  DFF_X1 \mem_reg[737][2]  ( .D(n20208), .CK(clk), .Q(\mem[737][2] ) );
  DFF_X1 \mem_reg[737][1]  ( .D(n20209), .CK(clk), .Q(\mem[737][1] ) );
  DFF_X1 \mem_reg[737][0]  ( .D(n20210), .CK(clk), .Q(\mem[737][0] ) );
  DFF_X1 \mem_reg[736][7]  ( .D(n20211), .CK(clk), .Q(\mem[736][7] ) );
  DFF_X1 \mem_reg[736][6]  ( .D(n20212), .CK(clk), .Q(\mem[736][6] ) );
  DFF_X1 \mem_reg[736][5]  ( .D(n20213), .CK(clk), .Q(\mem[736][5] ) );
  DFF_X1 \mem_reg[736][4]  ( .D(n20214), .CK(clk), .Q(\mem[736][4] ) );
  DFF_X1 \mem_reg[736][3]  ( .D(n20215), .CK(clk), .Q(\mem[736][3] ) );
  DFF_X1 \mem_reg[736][2]  ( .D(n20216), .CK(clk), .Q(\mem[736][2] ) );
  DFF_X1 \mem_reg[736][1]  ( .D(n20217), .CK(clk), .Q(\mem[736][1] ) );
  DFF_X1 \mem_reg[736][0]  ( .D(n20218), .CK(clk), .Q(\mem[736][0] ) );
  DFF_X1 \mem_reg[735][7]  ( .D(n20219), .CK(clk), .Q(\mem[735][7] ) );
  DFF_X1 \mem_reg[735][6]  ( .D(n20220), .CK(clk), .Q(\mem[735][6] ) );
  DFF_X1 \mem_reg[735][5]  ( .D(n20221), .CK(clk), .Q(\mem[735][5] ) );
  DFF_X1 \mem_reg[735][4]  ( .D(n20222), .CK(clk), .Q(\mem[735][4] ) );
  DFF_X1 \mem_reg[735][3]  ( .D(n20223), .CK(clk), .Q(\mem[735][3] ) );
  DFF_X1 \mem_reg[735][2]  ( .D(n20224), .CK(clk), .Q(\mem[735][2] ) );
  DFF_X1 \mem_reg[735][1]  ( .D(n20225), .CK(clk), .Q(\mem[735][1] ) );
  DFF_X1 \mem_reg[735][0]  ( .D(n20226), .CK(clk), .Q(\mem[735][0] ) );
  DFF_X1 \mem_reg[734][7]  ( .D(n20227), .CK(clk), .Q(\mem[734][7] ) );
  DFF_X1 \mem_reg[734][6]  ( .D(n20228), .CK(clk), .Q(\mem[734][6] ) );
  DFF_X1 \mem_reg[734][5]  ( .D(n20229), .CK(clk), .Q(\mem[734][5] ) );
  DFF_X1 \mem_reg[734][4]  ( .D(n20230), .CK(clk), .Q(\mem[734][4] ) );
  DFF_X1 \mem_reg[734][3]  ( .D(n20231), .CK(clk), .Q(\mem[734][3] ) );
  DFF_X1 \mem_reg[734][2]  ( .D(n20232), .CK(clk), .Q(\mem[734][2] ) );
  DFF_X1 \mem_reg[734][1]  ( .D(n20233), .CK(clk), .Q(\mem[734][1] ) );
  DFF_X1 \mem_reg[734][0]  ( .D(n20234), .CK(clk), .Q(\mem[734][0] ) );
  DFF_X1 \mem_reg[733][7]  ( .D(n20235), .CK(clk), .Q(\mem[733][7] ) );
  DFF_X1 \mem_reg[733][6]  ( .D(n20236), .CK(clk), .Q(\mem[733][6] ) );
  DFF_X1 \mem_reg[733][5]  ( .D(n20237), .CK(clk), .Q(\mem[733][5] ) );
  DFF_X1 \mem_reg[733][4]  ( .D(n20238), .CK(clk), .Q(\mem[733][4] ) );
  DFF_X1 \mem_reg[733][3]  ( .D(n20239), .CK(clk), .Q(\mem[733][3] ) );
  DFF_X1 \mem_reg[733][2]  ( .D(n20240), .CK(clk), .Q(\mem[733][2] ) );
  DFF_X1 \mem_reg[733][1]  ( .D(n20241), .CK(clk), .Q(\mem[733][1] ) );
  DFF_X1 \mem_reg[733][0]  ( .D(n20242), .CK(clk), .Q(\mem[733][0] ) );
  DFF_X1 \mem_reg[732][7]  ( .D(n20243), .CK(clk), .Q(\mem[732][7] ) );
  DFF_X1 \mem_reg[732][6]  ( .D(n20244), .CK(clk), .Q(\mem[732][6] ) );
  DFF_X1 \mem_reg[732][5]  ( .D(n20245), .CK(clk), .Q(\mem[732][5] ) );
  DFF_X1 \mem_reg[732][4]  ( .D(n20246), .CK(clk), .Q(\mem[732][4] ) );
  DFF_X1 \mem_reg[732][3]  ( .D(n20247), .CK(clk), .Q(\mem[732][3] ) );
  DFF_X1 \mem_reg[732][2]  ( .D(n20248), .CK(clk), .Q(\mem[732][2] ) );
  DFF_X1 \mem_reg[732][1]  ( .D(n20249), .CK(clk), .Q(\mem[732][1] ) );
  DFF_X1 \mem_reg[732][0]  ( .D(n20250), .CK(clk), .Q(\mem[732][0] ) );
  DFF_X1 \mem_reg[731][7]  ( .D(n20251), .CK(clk), .Q(\mem[731][7] ) );
  DFF_X1 \mem_reg[731][6]  ( .D(n20252), .CK(clk), .Q(\mem[731][6] ) );
  DFF_X1 \mem_reg[731][5]  ( .D(n20253), .CK(clk), .Q(\mem[731][5] ) );
  DFF_X1 \mem_reg[731][4]  ( .D(n20254), .CK(clk), .Q(\mem[731][4] ) );
  DFF_X1 \mem_reg[731][3]  ( .D(n20255), .CK(clk), .Q(\mem[731][3] ) );
  DFF_X1 \mem_reg[731][2]  ( .D(n20256), .CK(clk), .Q(\mem[731][2] ) );
  DFF_X1 \mem_reg[731][1]  ( .D(n20257), .CK(clk), .Q(\mem[731][1] ) );
  DFF_X1 \mem_reg[731][0]  ( .D(n20258), .CK(clk), .Q(\mem[731][0] ) );
  DFF_X1 \mem_reg[730][7]  ( .D(n20259), .CK(clk), .Q(\mem[730][7] ) );
  DFF_X1 \mem_reg[730][6]  ( .D(n20260), .CK(clk), .Q(\mem[730][6] ) );
  DFF_X1 \mem_reg[730][5]  ( .D(n20261), .CK(clk), .Q(\mem[730][5] ) );
  DFF_X1 \mem_reg[730][4]  ( .D(n20262), .CK(clk), .Q(\mem[730][4] ) );
  DFF_X1 \mem_reg[730][3]  ( .D(n20263), .CK(clk), .Q(\mem[730][3] ) );
  DFF_X1 \mem_reg[730][2]  ( .D(n20264), .CK(clk), .Q(\mem[730][2] ) );
  DFF_X1 \mem_reg[730][1]  ( .D(n20265), .CK(clk), .Q(\mem[730][1] ) );
  DFF_X1 \mem_reg[730][0]  ( .D(n20266), .CK(clk), .Q(\mem[730][0] ) );
  DFF_X1 \mem_reg[729][7]  ( .D(n20267), .CK(clk), .Q(\mem[729][7] ) );
  DFF_X1 \mem_reg[729][6]  ( .D(n20268), .CK(clk), .Q(\mem[729][6] ) );
  DFF_X1 \mem_reg[729][5]  ( .D(n20269), .CK(clk), .Q(\mem[729][5] ) );
  DFF_X1 \mem_reg[729][4]  ( .D(n20270), .CK(clk), .Q(\mem[729][4] ) );
  DFF_X1 \mem_reg[729][3]  ( .D(n20271), .CK(clk), .Q(\mem[729][3] ) );
  DFF_X1 \mem_reg[729][2]  ( .D(n20272), .CK(clk), .Q(\mem[729][2] ) );
  DFF_X1 \mem_reg[729][1]  ( .D(n20273), .CK(clk), .Q(\mem[729][1] ) );
  DFF_X1 \mem_reg[729][0]  ( .D(n20274), .CK(clk), .Q(\mem[729][0] ) );
  DFF_X1 \mem_reg[728][7]  ( .D(n20275), .CK(clk), .Q(\mem[728][7] ) );
  DFF_X1 \mem_reg[728][6]  ( .D(n20276), .CK(clk), .Q(\mem[728][6] ) );
  DFF_X1 \mem_reg[728][5]  ( .D(n20277), .CK(clk), .Q(\mem[728][5] ) );
  DFF_X1 \mem_reg[728][4]  ( .D(n20278), .CK(clk), .Q(\mem[728][4] ) );
  DFF_X1 \mem_reg[728][3]  ( .D(n20279), .CK(clk), .Q(\mem[728][3] ) );
  DFF_X1 \mem_reg[728][2]  ( .D(n20280), .CK(clk), .Q(\mem[728][2] ) );
  DFF_X1 \mem_reg[728][1]  ( .D(n20281), .CK(clk), .Q(\mem[728][1] ) );
  DFF_X1 \mem_reg[728][0]  ( .D(n20282), .CK(clk), .Q(\mem[728][0] ) );
  DFF_X1 \mem_reg[727][7]  ( .D(n20283), .CK(clk), .Q(\mem[727][7] ) );
  DFF_X1 \mem_reg[727][6]  ( .D(n20284), .CK(clk), .Q(\mem[727][6] ) );
  DFF_X1 \mem_reg[727][5]  ( .D(n20285), .CK(clk), .Q(\mem[727][5] ) );
  DFF_X1 \mem_reg[727][4]  ( .D(n20286), .CK(clk), .Q(\mem[727][4] ) );
  DFF_X1 \mem_reg[727][3]  ( .D(n20287), .CK(clk), .Q(\mem[727][3] ) );
  DFF_X1 \mem_reg[727][2]  ( .D(n20288), .CK(clk), .Q(\mem[727][2] ) );
  DFF_X1 \mem_reg[727][1]  ( .D(n20289), .CK(clk), .Q(\mem[727][1] ) );
  DFF_X1 \mem_reg[727][0]  ( .D(n20290), .CK(clk), .Q(\mem[727][0] ) );
  DFF_X1 \mem_reg[726][7]  ( .D(n20291), .CK(clk), .Q(\mem[726][7] ) );
  DFF_X1 \mem_reg[726][6]  ( .D(n20292), .CK(clk), .Q(\mem[726][6] ) );
  DFF_X1 \mem_reg[726][5]  ( .D(n20293), .CK(clk), .Q(\mem[726][5] ) );
  DFF_X1 \mem_reg[726][4]  ( .D(n20294), .CK(clk), .Q(\mem[726][4] ) );
  DFF_X1 \mem_reg[726][3]  ( .D(n20295), .CK(clk), .Q(\mem[726][3] ) );
  DFF_X1 \mem_reg[726][2]  ( .D(n20296), .CK(clk), .Q(\mem[726][2] ) );
  DFF_X1 \mem_reg[726][1]  ( .D(n20297), .CK(clk), .Q(\mem[726][1] ) );
  DFF_X1 \mem_reg[726][0]  ( .D(n20298), .CK(clk), .Q(\mem[726][0] ) );
  DFF_X1 \mem_reg[725][7]  ( .D(n20299), .CK(clk), .Q(\mem[725][7] ) );
  DFF_X1 \mem_reg[725][6]  ( .D(n20300), .CK(clk), .Q(\mem[725][6] ) );
  DFF_X1 \mem_reg[725][5]  ( .D(n20301), .CK(clk), .Q(\mem[725][5] ) );
  DFF_X1 \mem_reg[725][4]  ( .D(n20302), .CK(clk), .Q(\mem[725][4] ) );
  DFF_X1 \mem_reg[725][3]  ( .D(n20303), .CK(clk), .Q(\mem[725][3] ) );
  DFF_X1 \mem_reg[725][2]  ( .D(n20304), .CK(clk), .Q(\mem[725][2] ) );
  DFF_X1 \mem_reg[725][1]  ( .D(n20305), .CK(clk), .Q(\mem[725][1] ) );
  DFF_X1 \mem_reg[725][0]  ( .D(n20306), .CK(clk), .Q(\mem[725][0] ) );
  DFF_X1 \mem_reg[724][7]  ( .D(n20307), .CK(clk), .Q(\mem[724][7] ) );
  DFF_X1 \mem_reg[724][6]  ( .D(n20308), .CK(clk), .Q(\mem[724][6] ) );
  DFF_X1 \mem_reg[724][5]  ( .D(n20309), .CK(clk), .Q(\mem[724][5] ) );
  DFF_X1 \mem_reg[724][4]  ( .D(n20310), .CK(clk), .Q(\mem[724][4] ) );
  DFF_X1 \mem_reg[724][3]  ( .D(n20311), .CK(clk), .Q(\mem[724][3] ) );
  DFF_X1 \mem_reg[724][2]  ( .D(n20312), .CK(clk), .Q(\mem[724][2] ) );
  DFF_X1 \mem_reg[724][1]  ( .D(n20313), .CK(clk), .Q(\mem[724][1] ) );
  DFF_X1 \mem_reg[724][0]  ( .D(n20314), .CK(clk), .Q(\mem[724][0] ) );
  DFF_X1 \mem_reg[723][7]  ( .D(n20315), .CK(clk), .Q(\mem[723][7] ) );
  DFF_X1 \mem_reg[723][6]  ( .D(n20316), .CK(clk), .Q(\mem[723][6] ) );
  DFF_X1 \mem_reg[723][5]  ( .D(n20317), .CK(clk), .Q(\mem[723][5] ) );
  DFF_X1 \mem_reg[723][4]  ( .D(n20318), .CK(clk), .Q(\mem[723][4] ) );
  DFF_X1 \mem_reg[723][3]  ( .D(n20319), .CK(clk), .Q(\mem[723][3] ) );
  DFF_X1 \mem_reg[723][2]  ( .D(n20320), .CK(clk), .Q(\mem[723][2] ) );
  DFF_X1 \mem_reg[723][1]  ( .D(n20321), .CK(clk), .Q(\mem[723][1] ) );
  DFF_X1 \mem_reg[723][0]  ( .D(n20322), .CK(clk), .Q(\mem[723][0] ) );
  DFF_X1 \mem_reg[722][7]  ( .D(n20323), .CK(clk), .Q(\mem[722][7] ) );
  DFF_X1 \mem_reg[722][6]  ( .D(n20324), .CK(clk), .Q(\mem[722][6] ) );
  DFF_X1 \mem_reg[722][5]  ( .D(n20325), .CK(clk), .Q(\mem[722][5] ) );
  DFF_X1 \mem_reg[722][4]  ( .D(n20326), .CK(clk), .Q(\mem[722][4] ) );
  DFF_X1 \mem_reg[722][3]  ( .D(n20327), .CK(clk), .Q(\mem[722][3] ) );
  DFF_X1 \mem_reg[722][2]  ( .D(n20328), .CK(clk), .Q(\mem[722][2] ) );
  DFF_X1 \mem_reg[722][1]  ( .D(n20329), .CK(clk), .Q(\mem[722][1] ) );
  DFF_X1 \mem_reg[722][0]  ( .D(n20330), .CK(clk), .Q(\mem[722][0] ) );
  DFF_X1 \mem_reg[721][7]  ( .D(n20331), .CK(clk), .Q(\mem[721][7] ) );
  DFF_X1 \mem_reg[721][6]  ( .D(n20332), .CK(clk), .Q(\mem[721][6] ) );
  DFF_X1 \mem_reg[721][5]  ( .D(n20333), .CK(clk), .Q(\mem[721][5] ) );
  DFF_X1 \mem_reg[721][4]  ( .D(n20334), .CK(clk), .Q(\mem[721][4] ) );
  DFF_X1 \mem_reg[721][3]  ( .D(n20335), .CK(clk), .Q(\mem[721][3] ) );
  DFF_X1 \mem_reg[721][2]  ( .D(n20336), .CK(clk), .Q(\mem[721][2] ) );
  DFF_X1 \mem_reg[721][1]  ( .D(n20337), .CK(clk), .Q(\mem[721][1] ) );
  DFF_X1 \mem_reg[721][0]  ( .D(n20338), .CK(clk), .Q(\mem[721][0] ) );
  DFF_X1 \mem_reg[720][7]  ( .D(n20339), .CK(clk), .Q(\mem[720][7] ) );
  DFF_X1 \mem_reg[720][6]  ( .D(n20340), .CK(clk), .Q(\mem[720][6] ) );
  DFF_X1 \mem_reg[720][5]  ( .D(n20341), .CK(clk), .Q(\mem[720][5] ) );
  DFF_X1 \mem_reg[720][4]  ( .D(n20342), .CK(clk), .Q(\mem[720][4] ) );
  DFF_X1 \mem_reg[720][3]  ( .D(n20343), .CK(clk), .Q(\mem[720][3] ) );
  DFF_X1 \mem_reg[720][2]  ( .D(n20344), .CK(clk), .Q(\mem[720][2] ) );
  DFF_X1 \mem_reg[720][1]  ( .D(n20345), .CK(clk), .Q(\mem[720][1] ) );
  DFF_X1 \mem_reg[720][0]  ( .D(n20346), .CK(clk), .Q(\mem[720][0] ) );
  DFF_X1 \mem_reg[719][7]  ( .D(n20347), .CK(clk), .Q(\mem[719][7] ) );
  DFF_X1 \mem_reg[719][6]  ( .D(n20348), .CK(clk), .Q(\mem[719][6] ) );
  DFF_X1 \mem_reg[719][5]  ( .D(n20349), .CK(clk), .Q(\mem[719][5] ) );
  DFF_X1 \mem_reg[719][4]  ( .D(n20350), .CK(clk), .Q(\mem[719][4] ) );
  DFF_X1 \mem_reg[719][3]  ( .D(n20351), .CK(clk), .Q(\mem[719][3] ) );
  DFF_X1 \mem_reg[719][2]  ( .D(n20352), .CK(clk), .Q(\mem[719][2] ) );
  DFF_X1 \mem_reg[719][1]  ( .D(n20353), .CK(clk), .Q(\mem[719][1] ) );
  DFF_X1 \mem_reg[719][0]  ( .D(n20354), .CK(clk), .Q(\mem[719][0] ) );
  DFF_X1 \mem_reg[718][7]  ( .D(n20355), .CK(clk), .Q(\mem[718][7] ) );
  DFF_X1 \mem_reg[718][6]  ( .D(n20356), .CK(clk), .Q(\mem[718][6] ) );
  DFF_X1 \mem_reg[718][5]  ( .D(n20357), .CK(clk), .Q(\mem[718][5] ) );
  DFF_X1 \mem_reg[718][4]  ( .D(n20358), .CK(clk), .Q(\mem[718][4] ) );
  DFF_X1 \mem_reg[718][3]  ( .D(n20359), .CK(clk), .Q(\mem[718][3] ) );
  DFF_X1 \mem_reg[718][2]  ( .D(n20360), .CK(clk), .Q(\mem[718][2] ) );
  DFF_X1 \mem_reg[718][1]  ( .D(n20361), .CK(clk), .Q(\mem[718][1] ) );
  DFF_X1 \mem_reg[718][0]  ( .D(n20362), .CK(clk), .Q(\mem[718][0] ) );
  DFF_X1 \mem_reg[717][7]  ( .D(n20363), .CK(clk), .Q(\mem[717][7] ) );
  DFF_X1 \mem_reg[717][6]  ( .D(n20364), .CK(clk), .Q(\mem[717][6] ) );
  DFF_X1 \mem_reg[717][5]  ( .D(n20365), .CK(clk), .Q(\mem[717][5] ) );
  DFF_X1 \mem_reg[717][4]  ( .D(n20366), .CK(clk), .Q(\mem[717][4] ) );
  DFF_X1 \mem_reg[717][3]  ( .D(n20367), .CK(clk), .Q(\mem[717][3] ) );
  DFF_X1 \mem_reg[717][2]  ( .D(n20368), .CK(clk), .Q(\mem[717][2] ) );
  DFF_X1 \mem_reg[717][1]  ( .D(n20369), .CK(clk), .Q(\mem[717][1] ) );
  DFF_X1 \mem_reg[717][0]  ( .D(n20370), .CK(clk), .Q(\mem[717][0] ) );
  DFF_X1 \mem_reg[716][7]  ( .D(n20371), .CK(clk), .Q(\mem[716][7] ) );
  DFF_X1 \mem_reg[716][6]  ( .D(n20372), .CK(clk), .Q(\mem[716][6] ) );
  DFF_X1 \mem_reg[716][5]  ( .D(n20373), .CK(clk), .Q(\mem[716][5] ) );
  DFF_X1 \mem_reg[716][4]  ( .D(n20374), .CK(clk), .Q(\mem[716][4] ) );
  DFF_X1 \mem_reg[716][3]  ( .D(n20375), .CK(clk), .Q(\mem[716][3] ) );
  DFF_X1 \mem_reg[716][2]  ( .D(n20376), .CK(clk), .Q(\mem[716][2] ) );
  DFF_X1 \mem_reg[716][1]  ( .D(n20377), .CK(clk), .Q(\mem[716][1] ) );
  DFF_X1 \mem_reg[716][0]  ( .D(n20378), .CK(clk), .Q(\mem[716][0] ) );
  DFF_X1 \mem_reg[715][7]  ( .D(n20379), .CK(clk), .Q(\mem[715][7] ) );
  DFF_X1 \mem_reg[715][6]  ( .D(n20380), .CK(clk), .Q(\mem[715][6] ) );
  DFF_X1 \mem_reg[715][5]  ( .D(n20381), .CK(clk), .Q(\mem[715][5] ) );
  DFF_X1 \mem_reg[715][4]  ( .D(n20382), .CK(clk), .Q(\mem[715][4] ) );
  DFF_X1 \mem_reg[715][3]  ( .D(n20383), .CK(clk), .Q(\mem[715][3] ) );
  DFF_X1 \mem_reg[715][2]  ( .D(n20384), .CK(clk), .Q(\mem[715][2] ) );
  DFF_X1 \mem_reg[715][1]  ( .D(n20385), .CK(clk), .Q(\mem[715][1] ) );
  DFF_X1 \mem_reg[715][0]  ( .D(n20386), .CK(clk), .Q(\mem[715][0] ) );
  DFF_X1 \mem_reg[714][7]  ( .D(n20387), .CK(clk), .Q(\mem[714][7] ) );
  DFF_X1 \mem_reg[714][6]  ( .D(n20388), .CK(clk), .Q(\mem[714][6] ) );
  DFF_X1 \mem_reg[714][5]  ( .D(n20389), .CK(clk), .Q(\mem[714][5] ) );
  DFF_X1 \mem_reg[714][4]  ( .D(n20390), .CK(clk), .Q(\mem[714][4] ) );
  DFF_X1 \mem_reg[714][3]  ( .D(n20391), .CK(clk), .Q(\mem[714][3] ) );
  DFF_X1 \mem_reg[714][2]  ( .D(n20392), .CK(clk), .Q(\mem[714][2] ) );
  DFF_X1 \mem_reg[714][1]  ( .D(n20393), .CK(clk), .Q(\mem[714][1] ) );
  DFF_X1 \mem_reg[714][0]  ( .D(n20394), .CK(clk), .Q(\mem[714][0] ) );
  DFF_X1 \mem_reg[713][7]  ( .D(n20395), .CK(clk), .Q(\mem[713][7] ) );
  DFF_X1 \mem_reg[713][6]  ( .D(n20396), .CK(clk), .Q(\mem[713][6] ) );
  DFF_X1 \mem_reg[713][5]  ( .D(n20397), .CK(clk), .Q(\mem[713][5] ) );
  DFF_X1 \mem_reg[713][4]  ( .D(n20398), .CK(clk), .Q(\mem[713][4] ) );
  DFF_X1 \mem_reg[713][3]  ( .D(n20399), .CK(clk), .Q(\mem[713][3] ) );
  DFF_X1 \mem_reg[713][2]  ( .D(n20400), .CK(clk), .Q(\mem[713][2] ) );
  DFF_X1 \mem_reg[713][1]  ( .D(n20401), .CK(clk), .Q(\mem[713][1] ) );
  DFF_X1 \mem_reg[713][0]  ( .D(n20402), .CK(clk), .Q(\mem[713][0] ) );
  DFF_X1 \mem_reg[712][7]  ( .D(n20403), .CK(clk), .Q(\mem[712][7] ) );
  DFF_X1 \mem_reg[712][6]  ( .D(n20404), .CK(clk), .Q(\mem[712][6] ) );
  DFF_X1 \mem_reg[712][5]  ( .D(n20405), .CK(clk), .Q(\mem[712][5] ) );
  DFF_X1 \mem_reg[712][4]  ( .D(n20406), .CK(clk), .Q(\mem[712][4] ) );
  DFF_X1 \mem_reg[712][3]  ( .D(n20407), .CK(clk), .Q(\mem[712][3] ) );
  DFF_X1 \mem_reg[712][2]  ( .D(n20408), .CK(clk), .Q(\mem[712][2] ) );
  DFF_X1 \mem_reg[712][1]  ( .D(n20409), .CK(clk), .Q(\mem[712][1] ) );
  DFF_X1 \mem_reg[712][0]  ( .D(n20410), .CK(clk), .Q(\mem[712][0] ) );
  DFF_X1 \mem_reg[711][7]  ( .D(n20411), .CK(clk), .Q(\mem[711][7] ) );
  DFF_X1 \mem_reg[711][6]  ( .D(n20412), .CK(clk), .Q(\mem[711][6] ) );
  DFF_X1 \mem_reg[711][5]  ( .D(n20413), .CK(clk), .Q(\mem[711][5] ) );
  DFF_X1 \mem_reg[711][4]  ( .D(n20414), .CK(clk), .Q(\mem[711][4] ) );
  DFF_X1 \mem_reg[711][3]  ( .D(n20415), .CK(clk), .Q(\mem[711][3] ) );
  DFF_X1 \mem_reg[711][2]  ( .D(n20416), .CK(clk), .Q(\mem[711][2] ) );
  DFF_X1 \mem_reg[711][1]  ( .D(n20417), .CK(clk), .Q(\mem[711][1] ) );
  DFF_X1 \mem_reg[711][0]  ( .D(n20418), .CK(clk), .Q(\mem[711][0] ) );
  DFF_X1 \mem_reg[710][7]  ( .D(n20419), .CK(clk), .Q(\mem[710][7] ) );
  DFF_X1 \mem_reg[710][6]  ( .D(n20420), .CK(clk), .Q(\mem[710][6] ) );
  DFF_X1 \mem_reg[710][5]  ( .D(n20421), .CK(clk), .Q(\mem[710][5] ) );
  DFF_X1 \mem_reg[710][4]  ( .D(n20422), .CK(clk), .Q(\mem[710][4] ) );
  DFF_X1 \mem_reg[710][3]  ( .D(n20423), .CK(clk), .Q(\mem[710][3] ) );
  DFF_X1 \mem_reg[710][2]  ( .D(n20424), .CK(clk), .Q(\mem[710][2] ) );
  DFF_X1 \mem_reg[710][1]  ( .D(n20425), .CK(clk), .Q(\mem[710][1] ) );
  DFF_X1 \mem_reg[710][0]  ( .D(n20426), .CK(clk), .Q(\mem[710][0] ) );
  DFF_X1 \mem_reg[709][7]  ( .D(n20427), .CK(clk), .Q(\mem[709][7] ) );
  DFF_X1 \mem_reg[709][6]  ( .D(n20428), .CK(clk), .Q(\mem[709][6] ) );
  DFF_X1 \mem_reg[709][5]  ( .D(n20429), .CK(clk), .Q(\mem[709][5] ) );
  DFF_X1 \mem_reg[709][4]  ( .D(n20430), .CK(clk), .Q(\mem[709][4] ) );
  DFF_X1 \mem_reg[709][3]  ( .D(n20431), .CK(clk), .Q(\mem[709][3] ) );
  DFF_X1 \mem_reg[709][2]  ( .D(n20432), .CK(clk), .Q(\mem[709][2] ) );
  DFF_X1 \mem_reg[709][1]  ( .D(n20433), .CK(clk), .Q(\mem[709][1] ) );
  DFF_X1 \mem_reg[709][0]  ( .D(n20434), .CK(clk), .Q(\mem[709][0] ) );
  DFF_X1 \mem_reg[708][7]  ( .D(n20435), .CK(clk), .Q(\mem[708][7] ) );
  DFF_X1 \mem_reg[708][6]  ( .D(n20436), .CK(clk), .Q(\mem[708][6] ) );
  DFF_X1 \mem_reg[708][5]  ( .D(n20437), .CK(clk), .Q(\mem[708][5] ) );
  DFF_X1 \mem_reg[708][4]  ( .D(n20438), .CK(clk), .Q(\mem[708][4] ) );
  DFF_X1 \mem_reg[708][3]  ( .D(n20439), .CK(clk), .Q(\mem[708][3] ) );
  DFF_X1 \mem_reg[708][2]  ( .D(n20440), .CK(clk), .Q(\mem[708][2] ) );
  DFF_X1 \mem_reg[708][1]  ( .D(n20441), .CK(clk), .Q(\mem[708][1] ) );
  DFF_X1 \mem_reg[708][0]  ( .D(n20442), .CK(clk), .Q(\mem[708][0] ) );
  DFF_X1 \mem_reg[707][7]  ( .D(n20443), .CK(clk), .Q(\mem[707][7] ) );
  DFF_X1 \mem_reg[707][6]  ( .D(n20444), .CK(clk), .Q(\mem[707][6] ) );
  DFF_X1 \mem_reg[707][5]  ( .D(n20445), .CK(clk), .Q(\mem[707][5] ) );
  DFF_X1 \mem_reg[707][4]  ( .D(n20446), .CK(clk), .Q(\mem[707][4] ) );
  DFF_X1 \mem_reg[707][3]  ( .D(n20447), .CK(clk), .Q(\mem[707][3] ) );
  DFF_X1 \mem_reg[707][2]  ( .D(n20448), .CK(clk), .Q(\mem[707][2] ) );
  DFF_X1 \mem_reg[707][1]  ( .D(n20449), .CK(clk), .Q(\mem[707][1] ) );
  DFF_X1 \mem_reg[707][0]  ( .D(n20450), .CK(clk), .Q(\mem[707][0] ) );
  DFF_X1 \mem_reg[706][7]  ( .D(n20451), .CK(clk), .Q(\mem[706][7] ) );
  DFF_X1 \mem_reg[706][6]  ( .D(n20452), .CK(clk), .Q(\mem[706][6] ) );
  DFF_X1 \mem_reg[706][5]  ( .D(n20453), .CK(clk), .Q(\mem[706][5] ) );
  DFF_X1 \mem_reg[706][4]  ( .D(n20454), .CK(clk), .Q(\mem[706][4] ) );
  DFF_X1 \mem_reg[706][3]  ( .D(n20455), .CK(clk), .Q(\mem[706][3] ) );
  DFF_X1 \mem_reg[706][2]  ( .D(n20456), .CK(clk), .Q(\mem[706][2] ) );
  DFF_X1 \mem_reg[706][1]  ( .D(n20457), .CK(clk), .Q(\mem[706][1] ) );
  DFF_X1 \mem_reg[706][0]  ( .D(n20458), .CK(clk), .Q(\mem[706][0] ) );
  DFF_X1 \mem_reg[705][7]  ( .D(n20459), .CK(clk), .Q(\mem[705][7] ) );
  DFF_X1 \mem_reg[705][6]  ( .D(n20460), .CK(clk), .Q(\mem[705][6] ) );
  DFF_X1 \mem_reg[705][5]  ( .D(n20461), .CK(clk), .Q(\mem[705][5] ) );
  DFF_X1 \mem_reg[705][4]  ( .D(n20462), .CK(clk), .Q(\mem[705][4] ) );
  DFF_X1 \mem_reg[705][3]  ( .D(n20463), .CK(clk), .Q(\mem[705][3] ) );
  DFF_X1 \mem_reg[705][2]  ( .D(n20464), .CK(clk), .Q(\mem[705][2] ) );
  DFF_X1 \mem_reg[705][1]  ( .D(n20465), .CK(clk), .Q(\mem[705][1] ) );
  DFF_X1 \mem_reg[705][0]  ( .D(n20466), .CK(clk), .Q(\mem[705][0] ) );
  DFF_X1 \mem_reg[704][7]  ( .D(n20467), .CK(clk), .Q(\mem[704][7] ) );
  DFF_X1 \mem_reg[704][6]  ( .D(n20468), .CK(clk), .Q(\mem[704][6] ) );
  DFF_X1 \mem_reg[704][5]  ( .D(n20469), .CK(clk), .Q(\mem[704][5] ) );
  DFF_X1 \mem_reg[704][4]  ( .D(n20470), .CK(clk), .Q(\mem[704][4] ) );
  DFF_X1 \mem_reg[704][3]  ( .D(n20471), .CK(clk), .Q(\mem[704][3] ) );
  DFF_X1 \mem_reg[704][2]  ( .D(n20472), .CK(clk), .Q(\mem[704][2] ) );
  DFF_X1 \mem_reg[704][1]  ( .D(n20473), .CK(clk), .Q(\mem[704][1] ) );
  DFF_X1 \mem_reg[704][0]  ( .D(n20474), .CK(clk), .Q(\mem[704][0] ) );
  DFF_X1 \mem_reg[703][7]  ( .D(n20475), .CK(clk), .Q(\mem[703][7] ) );
  DFF_X1 \mem_reg[703][6]  ( .D(n20476), .CK(clk), .Q(\mem[703][6] ) );
  DFF_X1 \mem_reg[703][5]  ( .D(n20477), .CK(clk), .Q(\mem[703][5] ) );
  DFF_X1 \mem_reg[703][4]  ( .D(n20478), .CK(clk), .Q(\mem[703][4] ) );
  DFF_X1 \mem_reg[703][3]  ( .D(n20479), .CK(clk), .Q(\mem[703][3] ) );
  DFF_X1 \mem_reg[703][2]  ( .D(n20480), .CK(clk), .Q(\mem[703][2] ) );
  DFF_X1 \mem_reg[703][1]  ( .D(n20481), .CK(clk), .Q(\mem[703][1] ) );
  DFF_X1 \mem_reg[703][0]  ( .D(n20482), .CK(clk), .Q(\mem[703][0] ) );
  DFF_X1 \mem_reg[702][7]  ( .D(n20483), .CK(clk), .Q(\mem[702][7] ) );
  DFF_X1 \mem_reg[702][6]  ( .D(n20484), .CK(clk), .Q(\mem[702][6] ) );
  DFF_X1 \mem_reg[702][5]  ( .D(n20485), .CK(clk), .Q(\mem[702][5] ) );
  DFF_X1 \mem_reg[702][4]  ( .D(n20486), .CK(clk), .Q(\mem[702][4] ) );
  DFF_X1 \mem_reg[702][3]  ( .D(n20487), .CK(clk), .Q(\mem[702][3] ) );
  DFF_X1 \mem_reg[702][2]  ( .D(n20488), .CK(clk), .Q(\mem[702][2] ) );
  DFF_X1 \mem_reg[702][1]  ( .D(n20489), .CK(clk), .Q(\mem[702][1] ) );
  DFF_X1 \mem_reg[702][0]  ( .D(n20490), .CK(clk), .Q(\mem[702][0] ) );
  DFF_X1 \mem_reg[701][7]  ( .D(n20491), .CK(clk), .Q(\mem[701][7] ) );
  DFF_X1 \mem_reg[701][6]  ( .D(n20492), .CK(clk), .Q(\mem[701][6] ) );
  DFF_X1 \mem_reg[701][5]  ( .D(n20493), .CK(clk), .Q(\mem[701][5] ) );
  DFF_X1 \mem_reg[701][4]  ( .D(n20494), .CK(clk), .Q(\mem[701][4] ) );
  DFF_X1 \mem_reg[701][3]  ( .D(n20495), .CK(clk), .Q(\mem[701][3] ) );
  DFF_X1 \mem_reg[701][2]  ( .D(n20496), .CK(clk), .Q(\mem[701][2] ) );
  DFF_X1 \mem_reg[701][1]  ( .D(n20497), .CK(clk), .Q(\mem[701][1] ) );
  DFF_X1 \mem_reg[701][0]  ( .D(n20498), .CK(clk), .Q(\mem[701][0] ) );
  DFF_X1 \mem_reg[700][7]  ( .D(n20499), .CK(clk), .Q(\mem[700][7] ) );
  DFF_X1 \mem_reg[700][6]  ( .D(n20500), .CK(clk), .Q(\mem[700][6] ) );
  DFF_X1 \mem_reg[700][5]  ( .D(n20501), .CK(clk), .Q(\mem[700][5] ) );
  DFF_X1 \mem_reg[700][4]  ( .D(n20502), .CK(clk), .Q(\mem[700][4] ) );
  DFF_X1 \mem_reg[700][3]  ( .D(n20503), .CK(clk), .Q(\mem[700][3] ) );
  DFF_X1 \mem_reg[700][2]  ( .D(n20504), .CK(clk), .Q(\mem[700][2] ) );
  DFF_X1 \mem_reg[700][1]  ( .D(n20505), .CK(clk), .Q(\mem[700][1] ) );
  DFF_X1 \mem_reg[700][0]  ( .D(n20506), .CK(clk), .Q(\mem[700][0] ) );
  DFF_X1 \mem_reg[699][7]  ( .D(n20507), .CK(clk), .Q(\mem[699][7] ) );
  DFF_X1 \mem_reg[699][6]  ( .D(n20508), .CK(clk), .Q(\mem[699][6] ) );
  DFF_X1 \mem_reg[699][5]  ( .D(n20509), .CK(clk), .Q(\mem[699][5] ) );
  DFF_X1 \mem_reg[699][4]  ( .D(n20510), .CK(clk), .Q(\mem[699][4] ) );
  DFF_X1 \mem_reg[699][3]  ( .D(n20511), .CK(clk), .Q(\mem[699][3] ) );
  DFF_X1 \mem_reg[699][2]  ( .D(n20512), .CK(clk), .Q(\mem[699][2] ) );
  DFF_X1 \mem_reg[699][1]  ( .D(n20513), .CK(clk), .Q(\mem[699][1] ) );
  DFF_X1 \mem_reg[699][0]  ( .D(n20514), .CK(clk), .Q(\mem[699][0] ) );
  DFF_X1 \mem_reg[698][7]  ( .D(n20515), .CK(clk), .Q(\mem[698][7] ) );
  DFF_X1 \mem_reg[698][6]  ( .D(n20516), .CK(clk), .Q(\mem[698][6] ) );
  DFF_X1 \mem_reg[698][5]  ( .D(n20517), .CK(clk), .Q(\mem[698][5] ) );
  DFF_X1 \mem_reg[698][4]  ( .D(n20518), .CK(clk), .Q(\mem[698][4] ) );
  DFF_X1 \mem_reg[698][3]  ( .D(n20519), .CK(clk), .Q(\mem[698][3] ) );
  DFF_X1 \mem_reg[698][2]  ( .D(n20520), .CK(clk), .Q(\mem[698][2] ) );
  DFF_X1 \mem_reg[698][1]  ( .D(n20521), .CK(clk), .Q(\mem[698][1] ) );
  DFF_X1 \mem_reg[698][0]  ( .D(n20522), .CK(clk), .Q(\mem[698][0] ) );
  DFF_X1 \mem_reg[697][7]  ( .D(n20523), .CK(clk), .Q(\mem[697][7] ) );
  DFF_X1 \mem_reg[697][6]  ( .D(n20524), .CK(clk), .Q(\mem[697][6] ) );
  DFF_X1 \mem_reg[697][5]  ( .D(n20525), .CK(clk), .Q(\mem[697][5] ) );
  DFF_X1 \mem_reg[697][4]  ( .D(n20526), .CK(clk), .Q(\mem[697][4] ) );
  DFF_X1 \mem_reg[697][3]  ( .D(n20527), .CK(clk), .Q(\mem[697][3] ) );
  DFF_X1 \mem_reg[697][2]  ( .D(n20528), .CK(clk), .Q(\mem[697][2] ) );
  DFF_X1 \mem_reg[697][1]  ( .D(n20529), .CK(clk), .Q(\mem[697][1] ) );
  DFF_X1 \mem_reg[697][0]  ( .D(n20530), .CK(clk), .Q(\mem[697][0] ) );
  DFF_X1 \mem_reg[696][7]  ( .D(n20531), .CK(clk), .Q(\mem[696][7] ) );
  DFF_X1 \mem_reg[696][6]  ( .D(n20532), .CK(clk), .Q(\mem[696][6] ) );
  DFF_X1 \mem_reg[696][5]  ( .D(n20533), .CK(clk), .Q(\mem[696][5] ) );
  DFF_X1 \mem_reg[696][4]  ( .D(n20534), .CK(clk), .Q(\mem[696][4] ) );
  DFF_X1 \mem_reg[696][3]  ( .D(n20535), .CK(clk), .Q(\mem[696][3] ) );
  DFF_X1 \mem_reg[696][2]  ( .D(n20536), .CK(clk), .Q(\mem[696][2] ) );
  DFF_X1 \mem_reg[696][1]  ( .D(n20537), .CK(clk), .Q(\mem[696][1] ) );
  DFF_X1 \mem_reg[696][0]  ( .D(n20538), .CK(clk), .Q(\mem[696][0] ) );
  DFF_X1 \mem_reg[695][7]  ( .D(n20539), .CK(clk), .Q(\mem[695][7] ) );
  DFF_X1 \mem_reg[695][6]  ( .D(n20540), .CK(clk), .Q(\mem[695][6] ) );
  DFF_X1 \mem_reg[695][5]  ( .D(n20541), .CK(clk), .Q(\mem[695][5] ) );
  DFF_X1 \mem_reg[695][4]  ( .D(n20542), .CK(clk), .Q(\mem[695][4] ) );
  DFF_X1 \mem_reg[695][3]  ( .D(n20543), .CK(clk), .Q(\mem[695][3] ) );
  DFF_X1 \mem_reg[695][2]  ( .D(n20544), .CK(clk), .Q(\mem[695][2] ) );
  DFF_X1 \mem_reg[695][1]  ( .D(n20545), .CK(clk), .Q(\mem[695][1] ) );
  DFF_X1 \mem_reg[695][0]  ( .D(n20546), .CK(clk), .Q(\mem[695][0] ) );
  DFF_X1 \mem_reg[694][7]  ( .D(n20547), .CK(clk), .Q(\mem[694][7] ) );
  DFF_X1 \mem_reg[694][6]  ( .D(n20548), .CK(clk), .Q(\mem[694][6] ) );
  DFF_X1 \mem_reg[694][5]  ( .D(n20549), .CK(clk), .Q(\mem[694][5] ) );
  DFF_X1 \mem_reg[694][4]  ( .D(n20550), .CK(clk), .Q(\mem[694][4] ) );
  DFF_X1 \mem_reg[694][3]  ( .D(n20551), .CK(clk), .Q(\mem[694][3] ) );
  DFF_X1 \mem_reg[694][2]  ( .D(n20552), .CK(clk), .Q(\mem[694][2] ) );
  DFF_X1 \mem_reg[694][1]  ( .D(n20553), .CK(clk), .Q(\mem[694][1] ) );
  DFF_X1 \mem_reg[694][0]  ( .D(n20554), .CK(clk), .Q(\mem[694][0] ) );
  DFF_X1 \mem_reg[693][7]  ( .D(n20555), .CK(clk), .Q(\mem[693][7] ) );
  DFF_X1 \mem_reg[693][6]  ( .D(n20556), .CK(clk), .Q(\mem[693][6] ) );
  DFF_X1 \mem_reg[693][5]  ( .D(n20557), .CK(clk), .Q(\mem[693][5] ) );
  DFF_X1 \mem_reg[693][4]  ( .D(n20558), .CK(clk), .Q(\mem[693][4] ) );
  DFF_X1 \mem_reg[693][3]  ( .D(n20559), .CK(clk), .Q(\mem[693][3] ) );
  DFF_X1 \mem_reg[693][2]  ( .D(n20560), .CK(clk), .Q(\mem[693][2] ) );
  DFF_X1 \mem_reg[693][1]  ( .D(n20561), .CK(clk), .Q(\mem[693][1] ) );
  DFF_X1 \mem_reg[693][0]  ( .D(n20562), .CK(clk), .Q(\mem[693][0] ) );
  DFF_X1 \mem_reg[692][7]  ( .D(n20563), .CK(clk), .Q(\mem[692][7] ) );
  DFF_X1 \mem_reg[692][6]  ( .D(n20564), .CK(clk), .Q(\mem[692][6] ) );
  DFF_X1 \mem_reg[692][5]  ( .D(n20565), .CK(clk), .Q(\mem[692][5] ) );
  DFF_X1 \mem_reg[692][4]  ( .D(n20566), .CK(clk), .Q(\mem[692][4] ) );
  DFF_X1 \mem_reg[692][3]  ( .D(n20567), .CK(clk), .Q(\mem[692][3] ) );
  DFF_X1 \mem_reg[692][2]  ( .D(n20568), .CK(clk), .Q(\mem[692][2] ) );
  DFF_X1 \mem_reg[692][1]  ( .D(n20569), .CK(clk), .Q(\mem[692][1] ) );
  DFF_X1 \mem_reg[692][0]  ( .D(n20570), .CK(clk), .Q(\mem[692][0] ) );
  DFF_X1 \mem_reg[691][7]  ( .D(n20571), .CK(clk), .Q(\mem[691][7] ) );
  DFF_X1 \mem_reg[691][6]  ( .D(n20572), .CK(clk), .Q(\mem[691][6] ) );
  DFF_X1 \mem_reg[691][5]  ( .D(n20573), .CK(clk), .Q(\mem[691][5] ) );
  DFF_X1 \mem_reg[691][4]  ( .D(n20574), .CK(clk), .Q(\mem[691][4] ) );
  DFF_X1 \mem_reg[691][3]  ( .D(n20575), .CK(clk), .Q(\mem[691][3] ) );
  DFF_X1 \mem_reg[691][2]  ( .D(n20576), .CK(clk), .Q(\mem[691][2] ) );
  DFF_X1 \mem_reg[691][1]  ( .D(n20577), .CK(clk), .Q(\mem[691][1] ) );
  DFF_X1 \mem_reg[691][0]  ( .D(n20578), .CK(clk), .Q(\mem[691][0] ) );
  DFF_X1 \mem_reg[690][7]  ( .D(n20579), .CK(clk), .Q(\mem[690][7] ) );
  DFF_X1 \mem_reg[690][6]  ( .D(n20580), .CK(clk), .Q(\mem[690][6] ) );
  DFF_X1 \mem_reg[690][5]  ( .D(n20581), .CK(clk), .Q(\mem[690][5] ) );
  DFF_X1 \mem_reg[690][4]  ( .D(n20582), .CK(clk), .Q(\mem[690][4] ) );
  DFF_X1 \mem_reg[690][3]  ( .D(n20583), .CK(clk), .Q(\mem[690][3] ) );
  DFF_X1 \mem_reg[690][2]  ( .D(n20584), .CK(clk), .Q(\mem[690][2] ) );
  DFF_X1 \mem_reg[690][1]  ( .D(n20585), .CK(clk), .Q(\mem[690][1] ) );
  DFF_X1 \mem_reg[690][0]  ( .D(n20586), .CK(clk), .Q(\mem[690][0] ) );
  DFF_X1 \mem_reg[689][7]  ( .D(n20587), .CK(clk), .Q(\mem[689][7] ) );
  DFF_X1 \mem_reg[689][6]  ( .D(n20588), .CK(clk), .Q(\mem[689][6] ) );
  DFF_X1 \mem_reg[689][5]  ( .D(n20589), .CK(clk), .Q(\mem[689][5] ) );
  DFF_X1 \mem_reg[689][4]  ( .D(n20590), .CK(clk), .Q(\mem[689][4] ) );
  DFF_X1 \mem_reg[689][3]  ( .D(n20591), .CK(clk), .Q(\mem[689][3] ) );
  DFF_X1 \mem_reg[689][2]  ( .D(n20592), .CK(clk), .Q(\mem[689][2] ) );
  DFF_X1 \mem_reg[689][1]  ( .D(n20593), .CK(clk), .Q(\mem[689][1] ) );
  DFF_X1 \mem_reg[689][0]  ( .D(n20594), .CK(clk), .Q(\mem[689][0] ) );
  DFF_X1 \mem_reg[688][7]  ( .D(n20595), .CK(clk), .Q(\mem[688][7] ) );
  DFF_X1 \mem_reg[688][6]  ( .D(n20596), .CK(clk), .Q(\mem[688][6] ) );
  DFF_X1 \mem_reg[688][5]  ( .D(n20597), .CK(clk), .Q(\mem[688][5] ) );
  DFF_X1 \mem_reg[688][4]  ( .D(n20598), .CK(clk), .Q(\mem[688][4] ) );
  DFF_X1 \mem_reg[688][3]  ( .D(n20599), .CK(clk), .Q(\mem[688][3] ) );
  DFF_X1 \mem_reg[688][2]  ( .D(n20600), .CK(clk), .Q(\mem[688][2] ) );
  DFF_X1 \mem_reg[688][1]  ( .D(n20601), .CK(clk), .Q(\mem[688][1] ) );
  DFF_X1 \mem_reg[688][0]  ( .D(n20602), .CK(clk), .Q(\mem[688][0] ) );
  DFF_X1 \mem_reg[687][7]  ( .D(n20603), .CK(clk), .Q(\mem[687][7] ) );
  DFF_X1 \mem_reg[687][6]  ( .D(n20604), .CK(clk), .Q(\mem[687][6] ) );
  DFF_X1 \mem_reg[687][5]  ( .D(n20605), .CK(clk), .Q(\mem[687][5] ) );
  DFF_X1 \mem_reg[687][4]  ( .D(n20606), .CK(clk), .Q(\mem[687][4] ) );
  DFF_X1 \mem_reg[687][3]  ( .D(n20607), .CK(clk), .Q(\mem[687][3] ) );
  DFF_X1 \mem_reg[687][2]  ( .D(n20608), .CK(clk), .Q(\mem[687][2] ) );
  DFF_X1 \mem_reg[687][1]  ( .D(n20609), .CK(clk), .Q(\mem[687][1] ) );
  DFF_X1 \mem_reg[687][0]  ( .D(n20610), .CK(clk), .Q(\mem[687][0] ) );
  DFF_X1 \mem_reg[686][7]  ( .D(n20611), .CK(clk), .Q(\mem[686][7] ) );
  DFF_X1 \mem_reg[686][6]  ( .D(n20612), .CK(clk), .Q(\mem[686][6] ) );
  DFF_X1 \mem_reg[686][5]  ( .D(n20613), .CK(clk), .Q(\mem[686][5] ) );
  DFF_X1 \mem_reg[686][4]  ( .D(n20614), .CK(clk), .Q(\mem[686][4] ) );
  DFF_X1 \mem_reg[686][3]  ( .D(n20615), .CK(clk), .Q(\mem[686][3] ) );
  DFF_X1 \mem_reg[686][2]  ( .D(n20616), .CK(clk), .Q(\mem[686][2] ) );
  DFF_X1 \mem_reg[686][1]  ( .D(n20617), .CK(clk), .Q(\mem[686][1] ) );
  DFF_X1 \mem_reg[686][0]  ( .D(n20618), .CK(clk), .Q(\mem[686][0] ) );
  DFF_X1 \mem_reg[685][7]  ( .D(n20619), .CK(clk), .Q(\mem[685][7] ) );
  DFF_X1 \mem_reg[685][6]  ( .D(n20620), .CK(clk), .Q(\mem[685][6] ) );
  DFF_X1 \mem_reg[685][5]  ( .D(n20621), .CK(clk), .Q(\mem[685][5] ) );
  DFF_X1 \mem_reg[685][4]  ( .D(n20622), .CK(clk), .Q(\mem[685][4] ) );
  DFF_X1 \mem_reg[685][3]  ( .D(n20623), .CK(clk), .Q(\mem[685][3] ) );
  DFF_X1 \mem_reg[685][2]  ( .D(n20624), .CK(clk), .Q(\mem[685][2] ) );
  DFF_X1 \mem_reg[685][1]  ( .D(n20625), .CK(clk), .Q(\mem[685][1] ) );
  DFF_X1 \mem_reg[685][0]  ( .D(n20626), .CK(clk), .Q(\mem[685][0] ) );
  DFF_X1 \mem_reg[684][7]  ( .D(n20627), .CK(clk), .Q(\mem[684][7] ) );
  DFF_X1 \mem_reg[684][6]  ( .D(n20628), .CK(clk), .Q(\mem[684][6] ) );
  DFF_X1 \mem_reg[684][5]  ( .D(n20629), .CK(clk), .Q(\mem[684][5] ) );
  DFF_X1 \mem_reg[684][4]  ( .D(n20630), .CK(clk), .Q(\mem[684][4] ) );
  DFF_X1 \mem_reg[684][3]  ( .D(n20631), .CK(clk), .Q(\mem[684][3] ) );
  DFF_X1 \mem_reg[684][2]  ( .D(n20632), .CK(clk), .Q(\mem[684][2] ) );
  DFF_X1 \mem_reg[684][1]  ( .D(n20633), .CK(clk), .Q(\mem[684][1] ) );
  DFF_X1 \mem_reg[684][0]  ( .D(n20634), .CK(clk), .Q(\mem[684][0] ) );
  DFF_X1 \mem_reg[683][7]  ( .D(n20635), .CK(clk), .Q(\mem[683][7] ) );
  DFF_X1 \mem_reg[683][6]  ( .D(n20636), .CK(clk), .Q(\mem[683][6] ) );
  DFF_X1 \mem_reg[683][5]  ( .D(n20637), .CK(clk), .Q(\mem[683][5] ) );
  DFF_X1 \mem_reg[683][4]  ( .D(n20638), .CK(clk), .Q(\mem[683][4] ) );
  DFF_X1 \mem_reg[683][3]  ( .D(n20639), .CK(clk), .Q(\mem[683][3] ) );
  DFF_X1 \mem_reg[683][2]  ( .D(n20640), .CK(clk), .Q(\mem[683][2] ) );
  DFF_X1 \mem_reg[683][1]  ( .D(n20641), .CK(clk), .Q(\mem[683][1] ) );
  DFF_X1 \mem_reg[683][0]  ( .D(n20642), .CK(clk), .Q(\mem[683][0] ) );
  DFF_X1 \mem_reg[682][7]  ( .D(n20643), .CK(clk), .Q(\mem[682][7] ) );
  DFF_X1 \mem_reg[682][6]  ( .D(n20644), .CK(clk), .Q(\mem[682][6] ) );
  DFF_X1 \mem_reg[682][5]  ( .D(n20645), .CK(clk), .Q(\mem[682][5] ) );
  DFF_X1 \mem_reg[682][4]  ( .D(n20646), .CK(clk), .Q(\mem[682][4] ) );
  DFF_X1 \mem_reg[682][3]  ( .D(n20647), .CK(clk), .Q(\mem[682][3] ) );
  DFF_X1 \mem_reg[682][2]  ( .D(n20648), .CK(clk), .Q(\mem[682][2] ) );
  DFF_X1 \mem_reg[682][1]  ( .D(n20649), .CK(clk), .Q(\mem[682][1] ) );
  DFF_X1 \mem_reg[682][0]  ( .D(n20650), .CK(clk), .Q(\mem[682][0] ) );
  DFF_X1 \mem_reg[681][7]  ( .D(n20651), .CK(clk), .Q(\mem[681][7] ) );
  DFF_X1 \mem_reg[681][6]  ( .D(n20652), .CK(clk), .Q(\mem[681][6] ) );
  DFF_X1 \mem_reg[681][5]  ( .D(n20653), .CK(clk), .Q(\mem[681][5] ) );
  DFF_X1 \mem_reg[681][4]  ( .D(n20654), .CK(clk), .Q(\mem[681][4] ) );
  DFF_X1 \mem_reg[681][3]  ( .D(n20655), .CK(clk), .Q(\mem[681][3] ) );
  DFF_X1 \mem_reg[681][2]  ( .D(n20656), .CK(clk), .Q(\mem[681][2] ) );
  DFF_X1 \mem_reg[681][1]  ( .D(n20657), .CK(clk), .Q(\mem[681][1] ) );
  DFF_X1 \mem_reg[681][0]  ( .D(n20658), .CK(clk), .Q(\mem[681][0] ) );
  DFF_X1 \mem_reg[680][7]  ( .D(n20659), .CK(clk), .Q(\mem[680][7] ) );
  DFF_X1 \mem_reg[680][6]  ( .D(n20660), .CK(clk), .Q(\mem[680][6] ) );
  DFF_X1 \mem_reg[680][5]  ( .D(n20661), .CK(clk), .Q(\mem[680][5] ) );
  DFF_X1 \mem_reg[680][4]  ( .D(n20662), .CK(clk), .Q(\mem[680][4] ) );
  DFF_X1 \mem_reg[680][3]  ( .D(n20663), .CK(clk), .Q(\mem[680][3] ) );
  DFF_X1 \mem_reg[680][2]  ( .D(n20664), .CK(clk), .Q(\mem[680][2] ) );
  DFF_X1 \mem_reg[680][1]  ( .D(n20665), .CK(clk), .Q(\mem[680][1] ) );
  DFF_X1 \mem_reg[680][0]  ( .D(n20666), .CK(clk), .Q(\mem[680][0] ) );
  DFF_X1 \mem_reg[679][7]  ( .D(n20667), .CK(clk), .Q(\mem[679][7] ) );
  DFF_X1 \mem_reg[679][6]  ( .D(n20668), .CK(clk), .Q(\mem[679][6] ) );
  DFF_X1 \mem_reg[679][5]  ( .D(n20669), .CK(clk), .Q(\mem[679][5] ) );
  DFF_X1 \mem_reg[679][4]  ( .D(n20670), .CK(clk), .Q(\mem[679][4] ) );
  DFF_X1 \mem_reg[679][3]  ( .D(n20671), .CK(clk), .Q(\mem[679][3] ) );
  DFF_X1 \mem_reg[679][2]  ( .D(n20672), .CK(clk), .Q(\mem[679][2] ) );
  DFF_X1 \mem_reg[679][1]  ( .D(n20673), .CK(clk), .Q(\mem[679][1] ) );
  DFF_X1 \mem_reg[679][0]  ( .D(n20674), .CK(clk), .Q(\mem[679][0] ) );
  DFF_X1 \mem_reg[678][7]  ( .D(n20675), .CK(clk), .Q(\mem[678][7] ) );
  DFF_X1 \mem_reg[678][6]  ( .D(n20676), .CK(clk), .Q(\mem[678][6] ) );
  DFF_X1 \mem_reg[678][5]  ( .D(n20677), .CK(clk), .Q(\mem[678][5] ) );
  DFF_X1 \mem_reg[678][4]  ( .D(n20678), .CK(clk), .Q(\mem[678][4] ) );
  DFF_X1 \mem_reg[678][3]  ( .D(n20679), .CK(clk), .Q(\mem[678][3] ) );
  DFF_X1 \mem_reg[678][2]  ( .D(n20680), .CK(clk), .Q(\mem[678][2] ) );
  DFF_X1 \mem_reg[678][1]  ( .D(n20681), .CK(clk), .Q(\mem[678][1] ) );
  DFF_X1 \mem_reg[678][0]  ( .D(n20682), .CK(clk), .Q(\mem[678][0] ) );
  DFF_X1 \mem_reg[677][7]  ( .D(n20683), .CK(clk), .Q(\mem[677][7] ) );
  DFF_X1 \mem_reg[677][6]  ( .D(n20684), .CK(clk), .Q(\mem[677][6] ) );
  DFF_X1 \mem_reg[677][5]  ( .D(n20685), .CK(clk), .Q(\mem[677][5] ) );
  DFF_X1 \mem_reg[677][4]  ( .D(n20686), .CK(clk), .Q(\mem[677][4] ) );
  DFF_X1 \mem_reg[677][3]  ( .D(n20687), .CK(clk), .Q(\mem[677][3] ) );
  DFF_X1 \mem_reg[677][2]  ( .D(n20688), .CK(clk), .Q(\mem[677][2] ) );
  DFF_X1 \mem_reg[677][1]  ( .D(n20689), .CK(clk), .Q(\mem[677][1] ) );
  DFF_X1 \mem_reg[677][0]  ( .D(n20690), .CK(clk), .Q(\mem[677][0] ) );
  DFF_X1 \mem_reg[676][7]  ( .D(n20691), .CK(clk), .Q(\mem[676][7] ) );
  DFF_X1 \mem_reg[676][6]  ( .D(n20692), .CK(clk), .Q(\mem[676][6] ) );
  DFF_X1 \mem_reg[676][5]  ( .D(n20693), .CK(clk), .Q(\mem[676][5] ) );
  DFF_X1 \mem_reg[676][4]  ( .D(n20694), .CK(clk), .Q(\mem[676][4] ) );
  DFF_X1 \mem_reg[676][3]  ( .D(n20695), .CK(clk), .Q(\mem[676][3] ) );
  DFF_X1 \mem_reg[676][2]  ( .D(n20696), .CK(clk), .Q(\mem[676][2] ) );
  DFF_X1 \mem_reg[676][1]  ( .D(n20697), .CK(clk), .Q(\mem[676][1] ) );
  DFF_X1 \mem_reg[676][0]  ( .D(n20698), .CK(clk), .Q(\mem[676][0] ) );
  DFF_X1 \mem_reg[675][7]  ( .D(n20699), .CK(clk), .Q(\mem[675][7] ) );
  DFF_X1 \mem_reg[675][6]  ( .D(n20700), .CK(clk), .Q(\mem[675][6] ) );
  DFF_X1 \mem_reg[675][5]  ( .D(n20701), .CK(clk), .Q(\mem[675][5] ) );
  DFF_X1 \mem_reg[675][4]  ( .D(n20702), .CK(clk), .Q(\mem[675][4] ) );
  DFF_X1 \mem_reg[675][3]  ( .D(n20703), .CK(clk), .Q(\mem[675][3] ) );
  DFF_X1 \mem_reg[675][2]  ( .D(n20704), .CK(clk), .Q(\mem[675][2] ) );
  DFF_X1 \mem_reg[675][1]  ( .D(n20705), .CK(clk), .Q(\mem[675][1] ) );
  DFF_X1 \mem_reg[675][0]  ( .D(n20706), .CK(clk), .Q(\mem[675][0] ) );
  DFF_X1 \mem_reg[674][7]  ( .D(n20707), .CK(clk), .Q(\mem[674][7] ) );
  DFF_X1 \mem_reg[674][6]  ( .D(n20708), .CK(clk), .Q(\mem[674][6] ) );
  DFF_X1 \mem_reg[674][5]  ( .D(n20709), .CK(clk), .Q(\mem[674][5] ) );
  DFF_X1 \mem_reg[674][4]  ( .D(n20710), .CK(clk), .Q(\mem[674][4] ) );
  DFF_X1 \mem_reg[674][3]  ( .D(n20711), .CK(clk), .Q(\mem[674][3] ) );
  DFF_X1 \mem_reg[674][2]  ( .D(n20712), .CK(clk), .Q(\mem[674][2] ) );
  DFF_X1 \mem_reg[674][1]  ( .D(n20713), .CK(clk), .Q(\mem[674][1] ) );
  DFF_X1 \mem_reg[674][0]  ( .D(n20714), .CK(clk), .Q(\mem[674][0] ) );
  DFF_X1 \mem_reg[673][7]  ( .D(n20715), .CK(clk), .Q(\mem[673][7] ) );
  DFF_X1 \mem_reg[673][6]  ( .D(n20716), .CK(clk), .Q(\mem[673][6] ) );
  DFF_X1 \mem_reg[673][5]  ( .D(n20717), .CK(clk), .Q(\mem[673][5] ) );
  DFF_X1 \mem_reg[673][4]  ( .D(n20718), .CK(clk), .Q(\mem[673][4] ) );
  DFF_X1 \mem_reg[673][3]  ( .D(n20719), .CK(clk), .Q(\mem[673][3] ) );
  DFF_X1 \mem_reg[673][2]  ( .D(n20720), .CK(clk), .Q(\mem[673][2] ) );
  DFF_X1 \mem_reg[673][1]  ( .D(n20721), .CK(clk), .Q(\mem[673][1] ) );
  DFF_X1 \mem_reg[673][0]  ( .D(n20722), .CK(clk), .Q(\mem[673][0] ) );
  DFF_X1 \mem_reg[672][7]  ( .D(n20723), .CK(clk), .Q(\mem[672][7] ) );
  DFF_X1 \mem_reg[672][6]  ( .D(n20724), .CK(clk), .Q(\mem[672][6] ) );
  DFF_X1 \mem_reg[672][5]  ( .D(n20725), .CK(clk), .Q(\mem[672][5] ) );
  DFF_X1 \mem_reg[672][4]  ( .D(n20726), .CK(clk), .Q(\mem[672][4] ) );
  DFF_X1 \mem_reg[672][3]  ( .D(n20727), .CK(clk), .Q(\mem[672][3] ) );
  DFF_X1 \mem_reg[672][2]  ( .D(n20728), .CK(clk), .Q(\mem[672][2] ) );
  DFF_X1 \mem_reg[672][1]  ( .D(n20729), .CK(clk), .Q(\mem[672][1] ) );
  DFF_X1 \mem_reg[672][0]  ( .D(n20730), .CK(clk), .Q(\mem[672][0] ) );
  DFF_X1 \mem_reg[671][7]  ( .D(n20731), .CK(clk), .Q(\mem[671][7] ) );
  DFF_X1 \mem_reg[671][6]  ( .D(n20732), .CK(clk), .Q(\mem[671][6] ) );
  DFF_X1 \mem_reg[671][5]  ( .D(n20733), .CK(clk), .Q(\mem[671][5] ) );
  DFF_X1 \mem_reg[671][4]  ( .D(n20734), .CK(clk), .Q(\mem[671][4] ) );
  DFF_X1 \mem_reg[671][3]  ( .D(n20735), .CK(clk), .Q(\mem[671][3] ) );
  DFF_X1 \mem_reg[671][2]  ( .D(n20736), .CK(clk), .Q(\mem[671][2] ) );
  DFF_X1 \mem_reg[671][1]  ( .D(n20737), .CK(clk), .Q(\mem[671][1] ) );
  DFF_X1 \mem_reg[671][0]  ( .D(n20738), .CK(clk), .Q(\mem[671][0] ) );
  DFF_X1 \mem_reg[670][7]  ( .D(n20739), .CK(clk), .Q(\mem[670][7] ) );
  DFF_X1 \mem_reg[670][6]  ( .D(n20740), .CK(clk), .Q(\mem[670][6] ) );
  DFF_X1 \mem_reg[670][5]  ( .D(n20741), .CK(clk), .Q(\mem[670][5] ) );
  DFF_X1 \mem_reg[670][4]  ( .D(n20742), .CK(clk), .Q(\mem[670][4] ) );
  DFF_X1 \mem_reg[670][3]  ( .D(n20743), .CK(clk), .Q(\mem[670][3] ) );
  DFF_X1 \mem_reg[670][2]  ( .D(n20744), .CK(clk), .Q(\mem[670][2] ) );
  DFF_X1 \mem_reg[670][1]  ( .D(n20745), .CK(clk), .Q(\mem[670][1] ) );
  DFF_X1 \mem_reg[670][0]  ( .D(n20746), .CK(clk), .Q(\mem[670][0] ) );
  DFF_X1 \mem_reg[669][7]  ( .D(n20747), .CK(clk), .Q(\mem[669][7] ) );
  DFF_X1 \mem_reg[669][6]  ( .D(n20748), .CK(clk), .Q(\mem[669][6] ) );
  DFF_X1 \mem_reg[669][5]  ( .D(n20749), .CK(clk), .Q(\mem[669][5] ) );
  DFF_X1 \mem_reg[669][4]  ( .D(n20750), .CK(clk), .Q(\mem[669][4] ) );
  DFF_X1 \mem_reg[669][3]  ( .D(n20751), .CK(clk), .Q(\mem[669][3] ) );
  DFF_X1 \mem_reg[669][2]  ( .D(n20752), .CK(clk), .Q(\mem[669][2] ) );
  DFF_X1 \mem_reg[669][1]  ( .D(n20753), .CK(clk), .Q(\mem[669][1] ) );
  DFF_X1 \mem_reg[669][0]  ( .D(n20754), .CK(clk), .Q(\mem[669][0] ) );
  DFF_X1 \mem_reg[668][7]  ( .D(n20755), .CK(clk), .Q(\mem[668][7] ) );
  DFF_X1 \mem_reg[668][6]  ( .D(n20756), .CK(clk), .Q(\mem[668][6] ) );
  DFF_X1 \mem_reg[668][5]  ( .D(n20757), .CK(clk), .Q(\mem[668][5] ) );
  DFF_X1 \mem_reg[668][4]  ( .D(n20758), .CK(clk), .Q(\mem[668][4] ) );
  DFF_X1 \mem_reg[668][3]  ( .D(n20759), .CK(clk), .Q(\mem[668][3] ) );
  DFF_X1 \mem_reg[668][2]  ( .D(n20760), .CK(clk), .Q(\mem[668][2] ) );
  DFF_X1 \mem_reg[668][1]  ( .D(n20761), .CK(clk), .Q(\mem[668][1] ) );
  DFF_X1 \mem_reg[668][0]  ( .D(n20762), .CK(clk), .Q(\mem[668][0] ) );
  DFF_X1 \mem_reg[667][7]  ( .D(n20763), .CK(clk), .Q(\mem[667][7] ) );
  DFF_X1 \mem_reg[667][6]  ( .D(n20764), .CK(clk), .Q(\mem[667][6] ) );
  DFF_X1 \mem_reg[667][5]  ( .D(n20765), .CK(clk), .Q(\mem[667][5] ) );
  DFF_X1 \mem_reg[667][4]  ( .D(n20766), .CK(clk), .Q(\mem[667][4] ) );
  DFF_X1 \mem_reg[667][3]  ( .D(n20767), .CK(clk), .Q(\mem[667][3] ) );
  DFF_X1 \mem_reg[667][2]  ( .D(n20768), .CK(clk), .Q(\mem[667][2] ) );
  DFF_X1 \mem_reg[667][1]  ( .D(n20769), .CK(clk), .Q(\mem[667][1] ) );
  DFF_X1 \mem_reg[667][0]  ( .D(n20770), .CK(clk), .Q(\mem[667][0] ) );
  DFF_X1 \mem_reg[666][7]  ( .D(n20771), .CK(clk), .Q(\mem[666][7] ) );
  DFF_X1 \mem_reg[666][6]  ( .D(n20772), .CK(clk), .Q(\mem[666][6] ) );
  DFF_X1 \mem_reg[666][5]  ( .D(n20773), .CK(clk), .Q(\mem[666][5] ) );
  DFF_X1 \mem_reg[666][4]  ( .D(n20774), .CK(clk), .Q(\mem[666][4] ) );
  DFF_X1 \mem_reg[666][3]  ( .D(n20775), .CK(clk), .Q(\mem[666][3] ) );
  DFF_X1 \mem_reg[666][2]  ( .D(n20776), .CK(clk), .Q(\mem[666][2] ) );
  DFF_X1 \mem_reg[666][1]  ( .D(n20777), .CK(clk), .Q(\mem[666][1] ) );
  DFF_X1 \mem_reg[666][0]  ( .D(n20778), .CK(clk), .Q(\mem[666][0] ) );
  DFF_X1 \mem_reg[665][7]  ( .D(n20779), .CK(clk), .Q(\mem[665][7] ) );
  DFF_X1 \mem_reg[665][6]  ( .D(n20780), .CK(clk), .Q(\mem[665][6] ) );
  DFF_X1 \mem_reg[665][5]  ( .D(n20781), .CK(clk), .Q(\mem[665][5] ) );
  DFF_X1 \mem_reg[665][4]  ( .D(n20782), .CK(clk), .Q(\mem[665][4] ) );
  DFF_X1 \mem_reg[665][3]  ( .D(n20783), .CK(clk), .Q(\mem[665][3] ) );
  DFF_X1 \mem_reg[665][2]  ( .D(n20784), .CK(clk), .Q(\mem[665][2] ) );
  DFF_X1 \mem_reg[665][1]  ( .D(n20785), .CK(clk), .Q(\mem[665][1] ) );
  DFF_X1 \mem_reg[665][0]  ( .D(n20786), .CK(clk), .Q(\mem[665][0] ) );
  DFF_X1 \mem_reg[664][7]  ( .D(n20787), .CK(clk), .Q(\mem[664][7] ) );
  DFF_X1 \mem_reg[664][6]  ( .D(n20788), .CK(clk), .Q(\mem[664][6] ) );
  DFF_X1 \mem_reg[664][5]  ( .D(n20789), .CK(clk), .Q(\mem[664][5] ) );
  DFF_X1 \mem_reg[664][4]  ( .D(n20790), .CK(clk), .Q(\mem[664][4] ) );
  DFF_X1 \mem_reg[664][3]  ( .D(n20791), .CK(clk), .Q(\mem[664][3] ) );
  DFF_X1 \mem_reg[664][2]  ( .D(n20792), .CK(clk), .Q(\mem[664][2] ) );
  DFF_X1 \mem_reg[664][1]  ( .D(n20793), .CK(clk), .Q(\mem[664][1] ) );
  DFF_X1 \mem_reg[664][0]  ( .D(n20794), .CK(clk), .Q(\mem[664][0] ) );
  DFF_X1 \mem_reg[663][7]  ( .D(n20795), .CK(clk), .Q(\mem[663][7] ) );
  DFF_X1 \mem_reg[663][6]  ( .D(n20796), .CK(clk), .Q(\mem[663][6] ) );
  DFF_X1 \mem_reg[663][5]  ( .D(n20797), .CK(clk), .Q(\mem[663][5] ) );
  DFF_X1 \mem_reg[663][4]  ( .D(n20798), .CK(clk), .Q(\mem[663][4] ) );
  DFF_X1 \mem_reg[663][3]  ( .D(n20799), .CK(clk), .Q(\mem[663][3] ) );
  DFF_X1 \mem_reg[663][2]  ( .D(n20800), .CK(clk), .Q(\mem[663][2] ) );
  DFF_X1 \mem_reg[663][1]  ( .D(n20801), .CK(clk), .Q(\mem[663][1] ) );
  DFF_X1 \mem_reg[663][0]  ( .D(n20802), .CK(clk), .Q(\mem[663][0] ) );
  DFF_X1 \mem_reg[662][7]  ( .D(n20803), .CK(clk), .Q(\mem[662][7] ) );
  DFF_X1 \mem_reg[662][6]  ( .D(n20804), .CK(clk), .Q(\mem[662][6] ) );
  DFF_X1 \mem_reg[662][5]  ( .D(n20805), .CK(clk), .Q(\mem[662][5] ) );
  DFF_X1 \mem_reg[662][4]  ( .D(n20806), .CK(clk), .Q(\mem[662][4] ) );
  DFF_X1 \mem_reg[662][3]  ( .D(n20807), .CK(clk), .Q(\mem[662][3] ) );
  DFF_X1 \mem_reg[662][2]  ( .D(n20808), .CK(clk), .Q(\mem[662][2] ) );
  DFF_X1 \mem_reg[662][1]  ( .D(n20809), .CK(clk), .Q(\mem[662][1] ) );
  DFF_X1 \mem_reg[662][0]  ( .D(n20810), .CK(clk), .Q(\mem[662][0] ) );
  DFF_X1 \mem_reg[661][7]  ( .D(n20811), .CK(clk), .Q(\mem[661][7] ) );
  DFF_X1 \mem_reg[661][6]  ( .D(n20812), .CK(clk), .Q(\mem[661][6] ) );
  DFF_X1 \mem_reg[661][5]  ( .D(n20813), .CK(clk), .Q(\mem[661][5] ) );
  DFF_X1 \mem_reg[661][4]  ( .D(n20814), .CK(clk), .Q(\mem[661][4] ) );
  DFF_X1 \mem_reg[661][3]  ( .D(n20815), .CK(clk), .Q(\mem[661][3] ) );
  DFF_X1 \mem_reg[661][2]  ( .D(n20816), .CK(clk), .Q(\mem[661][2] ) );
  DFF_X1 \mem_reg[661][1]  ( .D(n20817), .CK(clk), .Q(\mem[661][1] ) );
  DFF_X1 \mem_reg[661][0]  ( .D(n20818), .CK(clk), .Q(\mem[661][0] ) );
  DFF_X1 \mem_reg[660][7]  ( .D(n20819), .CK(clk), .Q(\mem[660][7] ) );
  DFF_X1 \mem_reg[660][6]  ( .D(n20820), .CK(clk), .Q(\mem[660][6] ) );
  DFF_X1 \mem_reg[660][5]  ( .D(n20821), .CK(clk), .Q(\mem[660][5] ) );
  DFF_X1 \mem_reg[660][4]  ( .D(n20822), .CK(clk), .Q(\mem[660][4] ) );
  DFF_X1 \mem_reg[660][3]  ( .D(n20823), .CK(clk), .Q(\mem[660][3] ) );
  DFF_X1 \mem_reg[660][2]  ( .D(n20824), .CK(clk), .Q(\mem[660][2] ) );
  DFF_X1 \mem_reg[660][1]  ( .D(n20825), .CK(clk), .Q(\mem[660][1] ) );
  DFF_X1 \mem_reg[660][0]  ( .D(n20826), .CK(clk), .Q(\mem[660][0] ) );
  DFF_X1 \mem_reg[659][7]  ( .D(n20827), .CK(clk), .Q(\mem[659][7] ) );
  DFF_X1 \mem_reg[659][6]  ( .D(n20828), .CK(clk), .Q(\mem[659][6] ) );
  DFF_X1 \mem_reg[659][5]  ( .D(n20829), .CK(clk), .Q(\mem[659][5] ) );
  DFF_X1 \mem_reg[659][4]  ( .D(n20830), .CK(clk), .Q(\mem[659][4] ) );
  DFF_X1 \mem_reg[659][3]  ( .D(n20831), .CK(clk), .Q(\mem[659][3] ) );
  DFF_X1 \mem_reg[659][2]  ( .D(n20832), .CK(clk), .Q(\mem[659][2] ) );
  DFF_X1 \mem_reg[659][1]  ( .D(n20833), .CK(clk), .Q(\mem[659][1] ) );
  DFF_X1 \mem_reg[659][0]  ( .D(n20834), .CK(clk), .Q(\mem[659][0] ) );
  DFF_X1 \mem_reg[658][7]  ( .D(n20835), .CK(clk), .Q(\mem[658][7] ) );
  DFF_X1 \mem_reg[658][6]  ( .D(n20836), .CK(clk), .Q(\mem[658][6] ) );
  DFF_X1 \mem_reg[658][5]  ( .D(n20837), .CK(clk), .Q(\mem[658][5] ) );
  DFF_X1 \mem_reg[658][4]  ( .D(n20838), .CK(clk), .Q(\mem[658][4] ) );
  DFF_X1 \mem_reg[658][3]  ( .D(n20839), .CK(clk), .Q(\mem[658][3] ) );
  DFF_X1 \mem_reg[658][2]  ( .D(n20840), .CK(clk), .Q(\mem[658][2] ) );
  DFF_X1 \mem_reg[658][1]  ( .D(n20841), .CK(clk), .Q(\mem[658][1] ) );
  DFF_X1 \mem_reg[658][0]  ( .D(n20842), .CK(clk), .Q(\mem[658][0] ) );
  DFF_X1 \mem_reg[657][7]  ( .D(n20843), .CK(clk), .Q(\mem[657][7] ) );
  DFF_X1 \mem_reg[657][6]  ( .D(n20844), .CK(clk), .Q(\mem[657][6] ) );
  DFF_X1 \mem_reg[657][5]  ( .D(n20845), .CK(clk), .Q(\mem[657][5] ) );
  DFF_X1 \mem_reg[657][4]  ( .D(n20846), .CK(clk), .Q(\mem[657][4] ) );
  DFF_X1 \mem_reg[657][3]  ( .D(n20847), .CK(clk), .Q(\mem[657][3] ) );
  DFF_X1 \mem_reg[657][2]  ( .D(n20848), .CK(clk), .Q(\mem[657][2] ) );
  DFF_X1 \mem_reg[657][1]  ( .D(n20849), .CK(clk), .Q(\mem[657][1] ) );
  DFF_X1 \mem_reg[657][0]  ( .D(n20850), .CK(clk), .Q(\mem[657][0] ) );
  DFF_X1 \mem_reg[656][7]  ( .D(n20851), .CK(clk), .Q(\mem[656][7] ) );
  DFF_X1 \mem_reg[656][6]  ( .D(n20852), .CK(clk), .Q(\mem[656][6] ) );
  DFF_X1 \mem_reg[656][5]  ( .D(n20853), .CK(clk), .Q(\mem[656][5] ) );
  DFF_X1 \mem_reg[656][4]  ( .D(n20854), .CK(clk), .Q(\mem[656][4] ) );
  DFF_X1 \mem_reg[656][3]  ( .D(n20855), .CK(clk), .Q(\mem[656][3] ) );
  DFF_X1 \mem_reg[656][2]  ( .D(n20856), .CK(clk), .Q(\mem[656][2] ) );
  DFF_X1 \mem_reg[656][1]  ( .D(n20857), .CK(clk), .Q(\mem[656][1] ) );
  DFF_X1 \mem_reg[656][0]  ( .D(n20858), .CK(clk), .Q(\mem[656][0] ) );
  DFF_X1 \mem_reg[655][7]  ( .D(n20859), .CK(clk), .Q(\mem[655][7] ) );
  DFF_X1 \mem_reg[655][6]  ( .D(n20860), .CK(clk), .Q(\mem[655][6] ) );
  DFF_X1 \mem_reg[655][5]  ( .D(n20861), .CK(clk), .Q(\mem[655][5] ) );
  DFF_X1 \mem_reg[655][4]  ( .D(n20862), .CK(clk), .Q(\mem[655][4] ) );
  DFF_X1 \mem_reg[655][3]  ( .D(n20863), .CK(clk), .Q(\mem[655][3] ) );
  DFF_X1 \mem_reg[655][2]  ( .D(n20864), .CK(clk), .Q(\mem[655][2] ) );
  DFF_X1 \mem_reg[655][1]  ( .D(n20865), .CK(clk), .Q(\mem[655][1] ) );
  DFF_X1 \mem_reg[655][0]  ( .D(n20866), .CK(clk), .Q(\mem[655][0] ) );
  DFF_X1 \mem_reg[654][7]  ( .D(n20867), .CK(clk), .Q(\mem[654][7] ) );
  DFF_X1 \mem_reg[654][6]  ( .D(n20868), .CK(clk), .Q(\mem[654][6] ) );
  DFF_X1 \mem_reg[654][5]  ( .D(n20869), .CK(clk), .Q(\mem[654][5] ) );
  DFF_X1 \mem_reg[654][4]  ( .D(n20870), .CK(clk), .Q(\mem[654][4] ) );
  DFF_X1 \mem_reg[654][3]  ( .D(n20871), .CK(clk), .Q(\mem[654][3] ) );
  DFF_X1 \mem_reg[654][2]  ( .D(n20872), .CK(clk), .Q(\mem[654][2] ) );
  DFF_X1 \mem_reg[654][1]  ( .D(n20873), .CK(clk), .Q(\mem[654][1] ) );
  DFF_X1 \mem_reg[654][0]  ( .D(n20874), .CK(clk), .Q(\mem[654][0] ) );
  DFF_X1 \mem_reg[653][7]  ( .D(n20875), .CK(clk), .Q(\mem[653][7] ) );
  DFF_X1 \mem_reg[653][6]  ( .D(n20876), .CK(clk), .Q(\mem[653][6] ) );
  DFF_X1 \mem_reg[653][5]  ( .D(n20877), .CK(clk), .Q(\mem[653][5] ) );
  DFF_X1 \mem_reg[653][4]  ( .D(n20878), .CK(clk), .Q(\mem[653][4] ) );
  DFF_X1 \mem_reg[653][3]  ( .D(n20879), .CK(clk), .Q(\mem[653][3] ) );
  DFF_X1 \mem_reg[653][2]  ( .D(n20880), .CK(clk), .Q(\mem[653][2] ) );
  DFF_X1 \mem_reg[653][1]  ( .D(n20881), .CK(clk), .Q(\mem[653][1] ) );
  DFF_X1 \mem_reg[653][0]  ( .D(n20882), .CK(clk), .Q(\mem[653][0] ) );
  DFF_X1 \mem_reg[652][7]  ( .D(n20883), .CK(clk), .Q(\mem[652][7] ) );
  DFF_X1 \mem_reg[652][6]  ( .D(n20884), .CK(clk), .Q(\mem[652][6] ) );
  DFF_X1 \mem_reg[652][5]  ( .D(n20885), .CK(clk), .Q(\mem[652][5] ) );
  DFF_X1 \mem_reg[652][4]  ( .D(n20886), .CK(clk), .Q(\mem[652][4] ) );
  DFF_X1 \mem_reg[652][3]  ( .D(n20887), .CK(clk), .Q(\mem[652][3] ) );
  DFF_X1 \mem_reg[652][2]  ( .D(n20888), .CK(clk), .Q(\mem[652][2] ) );
  DFF_X1 \mem_reg[652][1]  ( .D(n20889), .CK(clk), .Q(\mem[652][1] ) );
  DFF_X1 \mem_reg[652][0]  ( .D(n20890), .CK(clk), .Q(\mem[652][0] ) );
  DFF_X1 \mem_reg[651][7]  ( .D(n20891), .CK(clk), .Q(\mem[651][7] ) );
  DFF_X1 \mem_reg[651][6]  ( .D(n20892), .CK(clk), .Q(\mem[651][6] ) );
  DFF_X1 \mem_reg[651][5]  ( .D(n20893), .CK(clk), .Q(\mem[651][5] ) );
  DFF_X1 \mem_reg[651][4]  ( .D(n20894), .CK(clk), .Q(\mem[651][4] ) );
  DFF_X1 \mem_reg[651][3]  ( .D(n20895), .CK(clk), .Q(\mem[651][3] ) );
  DFF_X1 \mem_reg[651][2]  ( .D(n20896), .CK(clk), .Q(\mem[651][2] ) );
  DFF_X1 \mem_reg[651][1]  ( .D(n20897), .CK(clk), .Q(\mem[651][1] ) );
  DFF_X1 \mem_reg[651][0]  ( .D(n20898), .CK(clk), .Q(\mem[651][0] ) );
  DFF_X1 \mem_reg[650][7]  ( .D(n20899), .CK(clk), .Q(\mem[650][7] ) );
  DFF_X1 \mem_reg[650][6]  ( .D(n20900), .CK(clk), .Q(\mem[650][6] ) );
  DFF_X1 \mem_reg[650][5]  ( .D(n20901), .CK(clk), .Q(\mem[650][5] ) );
  DFF_X1 \mem_reg[650][4]  ( .D(n20902), .CK(clk), .Q(\mem[650][4] ) );
  DFF_X1 \mem_reg[650][3]  ( .D(n20903), .CK(clk), .Q(\mem[650][3] ) );
  DFF_X1 \mem_reg[650][2]  ( .D(n20904), .CK(clk), .Q(\mem[650][2] ) );
  DFF_X1 \mem_reg[650][1]  ( .D(n20905), .CK(clk), .Q(\mem[650][1] ) );
  DFF_X1 \mem_reg[650][0]  ( .D(n20906), .CK(clk), .Q(\mem[650][0] ) );
  DFF_X1 \mem_reg[649][7]  ( .D(n20907), .CK(clk), .Q(\mem[649][7] ) );
  DFF_X1 \mem_reg[649][6]  ( .D(n20908), .CK(clk), .Q(\mem[649][6] ) );
  DFF_X1 \mem_reg[649][5]  ( .D(n20909), .CK(clk), .Q(\mem[649][5] ) );
  DFF_X1 \mem_reg[649][4]  ( .D(n20910), .CK(clk), .Q(\mem[649][4] ) );
  DFF_X1 \mem_reg[649][3]  ( .D(n20911), .CK(clk), .Q(\mem[649][3] ) );
  DFF_X1 \mem_reg[649][2]  ( .D(n20912), .CK(clk), .Q(\mem[649][2] ) );
  DFF_X1 \mem_reg[649][1]  ( .D(n20913), .CK(clk), .Q(\mem[649][1] ) );
  DFF_X1 \mem_reg[649][0]  ( .D(n20914), .CK(clk), .Q(\mem[649][0] ) );
  DFF_X1 \mem_reg[648][7]  ( .D(n20915), .CK(clk), .Q(\mem[648][7] ) );
  DFF_X1 \mem_reg[648][6]  ( .D(n20916), .CK(clk), .Q(\mem[648][6] ) );
  DFF_X1 \mem_reg[648][5]  ( .D(n20917), .CK(clk), .Q(\mem[648][5] ) );
  DFF_X1 \mem_reg[648][4]  ( .D(n20918), .CK(clk), .Q(\mem[648][4] ) );
  DFF_X1 \mem_reg[648][3]  ( .D(n20919), .CK(clk), .Q(\mem[648][3] ) );
  DFF_X1 \mem_reg[648][2]  ( .D(n20920), .CK(clk), .Q(\mem[648][2] ) );
  DFF_X1 \mem_reg[648][1]  ( .D(n20921), .CK(clk), .Q(\mem[648][1] ) );
  DFF_X1 \mem_reg[648][0]  ( .D(n20922), .CK(clk), .Q(\mem[648][0] ) );
  DFF_X1 \mem_reg[647][7]  ( .D(n20923), .CK(clk), .Q(\mem[647][7] ) );
  DFF_X1 \mem_reg[647][6]  ( .D(n20924), .CK(clk), .Q(\mem[647][6] ) );
  DFF_X1 \mem_reg[647][5]  ( .D(n20925), .CK(clk), .Q(\mem[647][5] ) );
  DFF_X1 \mem_reg[647][4]  ( .D(n20926), .CK(clk), .Q(\mem[647][4] ) );
  DFF_X1 \mem_reg[647][3]  ( .D(n20927), .CK(clk), .Q(\mem[647][3] ) );
  DFF_X1 \mem_reg[647][2]  ( .D(n20928), .CK(clk), .Q(\mem[647][2] ) );
  DFF_X1 \mem_reg[647][1]  ( .D(n20929), .CK(clk), .Q(\mem[647][1] ) );
  DFF_X1 \mem_reg[647][0]  ( .D(n20930), .CK(clk), .Q(\mem[647][0] ) );
  DFF_X1 \mem_reg[646][7]  ( .D(n20931), .CK(clk), .Q(\mem[646][7] ) );
  DFF_X1 \mem_reg[646][6]  ( .D(n20932), .CK(clk), .Q(\mem[646][6] ) );
  DFF_X1 \mem_reg[646][5]  ( .D(n20933), .CK(clk), .Q(\mem[646][5] ) );
  DFF_X1 \mem_reg[646][4]  ( .D(n20934), .CK(clk), .Q(\mem[646][4] ) );
  DFF_X1 \mem_reg[646][3]  ( .D(n20935), .CK(clk), .Q(\mem[646][3] ) );
  DFF_X1 \mem_reg[646][2]  ( .D(n20936), .CK(clk), .Q(\mem[646][2] ) );
  DFF_X1 \mem_reg[646][1]  ( .D(n20937), .CK(clk), .Q(\mem[646][1] ) );
  DFF_X1 \mem_reg[646][0]  ( .D(n20938), .CK(clk), .Q(\mem[646][0] ) );
  DFF_X1 \mem_reg[645][7]  ( .D(n20939), .CK(clk), .Q(\mem[645][7] ) );
  DFF_X1 \mem_reg[645][6]  ( .D(n20940), .CK(clk), .Q(\mem[645][6] ) );
  DFF_X1 \mem_reg[645][5]  ( .D(n20941), .CK(clk), .Q(\mem[645][5] ) );
  DFF_X1 \mem_reg[645][4]  ( .D(n20942), .CK(clk), .Q(\mem[645][4] ) );
  DFF_X1 \mem_reg[645][3]  ( .D(n20943), .CK(clk), .Q(\mem[645][3] ) );
  DFF_X1 \mem_reg[645][2]  ( .D(n20944), .CK(clk), .Q(\mem[645][2] ) );
  DFF_X1 \mem_reg[645][1]  ( .D(n20945), .CK(clk), .Q(\mem[645][1] ) );
  DFF_X1 \mem_reg[645][0]  ( .D(n20946), .CK(clk), .Q(\mem[645][0] ) );
  DFF_X1 \mem_reg[644][7]  ( .D(n20947), .CK(clk), .Q(\mem[644][7] ) );
  DFF_X1 \mem_reg[644][6]  ( .D(n20948), .CK(clk), .Q(\mem[644][6] ) );
  DFF_X1 \mem_reg[644][5]  ( .D(n20949), .CK(clk), .Q(\mem[644][5] ) );
  DFF_X1 \mem_reg[644][4]  ( .D(n20950), .CK(clk), .Q(\mem[644][4] ) );
  DFF_X1 \mem_reg[644][3]  ( .D(n20951), .CK(clk), .Q(\mem[644][3] ) );
  DFF_X1 \mem_reg[644][2]  ( .D(n20952), .CK(clk), .Q(\mem[644][2] ) );
  DFF_X1 \mem_reg[644][1]  ( .D(n20953), .CK(clk), .Q(\mem[644][1] ) );
  DFF_X1 \mem_reg[644][0]  ( .D(n20954), .CK(clk), .Q(\mem[644][0] ) );
  DFF_X1 \mem_reg[643][7]  ( .D(n20955), .CK(clk), .Q(\mem[643][7] ) );
  DFF_X1 \mem_reg[643][6]  ( .D(n20956), .CK(clk), .Q(\mem[643][6] ) );
  DFF_X1 \mem_reg[643][5]  ( .D(n20957), .CK(clk), .Q(\mem[643][5] ) );
  DFF_X1 \mem_reg[643][4]  ( .D(n20958), .CK(clk), .Q(\mem[643][4] ) );
  DFF_X1 \mem_reg[643][3]  ( .D(n20959), .CK(clk), .Q(\mem[643][3] ) );
  DFF_X1 \mem_reg[643][2]  ( .D(n20960), .CK(clk), .Q(\mem[643][2] ) );
  DFF_X1 \mem_reg[643][1]  ( .D(n20961), .CK(clk), .Q(\mem[643][1] ) );
  DFF_X1 \mem_reg[643][0]  ( .D(n20962), .CK(clk), .Q(\mem[643][0] ) );
  DFF_X1 \mem_reg[642][7]  ( .D(n20963), .CK(clk), .Q(\mem[642][7] ) );
  DFF_X1 \mem_reg[642][6]  ( .D(n20964), .CK(clk), .Q(\mem[642][6] ) );
  DFF_X1 \mem_reg[642][5]  ( .D(n20965), .CK(clk), .Q(\mem[642][5] ) );
  DFF_X1 \mem_reg[642][4]  ( .D(n20966), .CK(clk), .Q(\mem[642][4] ) );
  DFF_X1 \mem_reg[642][3]  ( .D(n20967), .CK(clk), .Q(\mem[642][3] ) );
  DFF_X1 \mem_reg[642][2]  ( .D(n20968), .CK(clk), .Q(\mem[642][2] ) );
  DFF_X1 \mem_reg[642][1]  ( .D(n20969), .CK(clk), .Q(\mem[642][1] ) );
  DFF_X1 \mem_reg[642][0]  ( .D(n20970), .CK(clk), .Q(\mem[642][0] ) );
  DFF_X1 \mem_reg[641][7]  ( .D(n20971), .CK(clk), .Q(\mem[641][7] ) );
  DFF_X1 \mem_reg[641][6]  ( .D(n20972), .CK(clk), .Q(\mem[641][6] ) );
  DFF_X1 \mem_reg[641][5]  ( .D(n20973), .CK(clk), .Q(\mem[641][5] ) );
  DFF_X1 \mem_reg[641][4]  ( .D(n20974), .CK(clk), .Q(\mem[641][4] ) );
  DFF_X1 \mem_reg[641][3]  ( .D(n20975), .CK(clk), .Q(\mem[641][3] ) );
  DFF_X1 \mem_reg[641][2]  ( .D(n20976), .CK(clk), .Q(\mem[641][2] ) );
  DFF_X1 \mem_reg[641][1]  ( .D(n20977), .CK(clk), .Q(\mem[641][1] ) );
  DFF_X1 \mem_reg[641][0]  ( .D(n20978), .CK(clk), .Q(\mem[641][0] ) );
  DFF_X1 \mem_reg[640][7]  ( .D(n20979), .CK(clk), .Q(\mem[640][7] ) );
  DFF_X1 \mem_reg[640][6]  ( .D(n20980), .CK(clk), .Q(\mem[640][6] ) );
  DFF_X1 \mem_reg[640][5]  ( .D(n20981), .CK(clk), .Q(\mem[640][5] ) );
  DFF_X1 \mem_reg[640][4]  ( .D(n20982), .CK(clk), .Q(\mem[640][4] ) );
  DFF_X1 \mem_reg[640][3]  ( .D(n20983), .CK(clk), .Q(\mem[640][3] ) );
  DFF_X1 \mem_reg[640][2]  ( .D(n20984), .CK(clk), .Q(\mem[640][2] ) );
  DFF_X1 \mem_reg[640][1]  ( .D(n20985), .CK(clk), .Q(\mem[640][1] ) );
  DFF_X1 \mem_reg[640][0]  ( .D(n20986), .CK(clk), .Q(\mem[640][0] ) );
  DFF_X1 \mem_reg[639][7]  ( .D(n20987), .CK(clk), .Q(\mem[639][7] ) );
  DFF_X1 \mem_reg[639][6]  ( .D(n20988), .CK(clk), .Q(\mem[639][6] ) );
  DFF_X1 \mem_reg[639][5]  ( .D(n20989), .CK(clk), .Q(\mem[639][5] ) );
  DFF_X1 \mem_reg[639][4]  ( .D(n20990), .CK(clk), .Q(\mem[639][4] ) );
  DFF_X1 \mem_reg[639][3]  ( .D(n20991), .CK(clk), .Q(\mem[639][3] ) );
  DFF_X1 \mem_reg[639][2]  ( .D(n20992), .CK(clk), .Q(\mem[639][2] ) );
  DFF_X1 \mem_reg[639][1]  ( .D(n20993), .CK(clk), .Q(\mem[639][1] ) );
  DFF_X1 \mem_reg[639][0]  ( .D(n20994), .CK(clk), .Q(\mem[639][0] ) );
  DFF_X1 \mem_reg[638][7]  ( .D(n20995), .CK(clk), .Q(\mem[638][7] ) );
  DFF_X1 \mem_reg[638][6]  ( .D(n20996), .CK(clk), .Q(\mem[638][6] ) );
  DFF_X1 \mem_reg[638][5]  ( .D(n20997), .CK(clk), .Q(\mem[638][5] ) );
  DFF_X1 \mem_reg[638][4]  ( .D(n20998), .CK(clk), .Q(\mem[638][4] ) );
  DFF_X1 \mem_reg[638][3]  ( .D(n20999), .CK(clk), .Q(\mem[638][3] ) );
  DFF_X1 \mem_reg[638][2]  ( .D(n21000), .CK(clk), .Q(\mem[638][2] ) );
  DFF_X1 \mem_reg[638][1]  ( .D(n21001), .CK(clk), .Q(\mem[638][1] ) );
  DFF_X1 \mem_reg[638][0]  ( .D(n21002), .CK(clk), .Q(\mem[638][0] ) );
  DFF_X1 \mem_reg[637][7]  ( .D(n21003), .CK(clk), .Q(\mem[637][7] ) );
  DFF_X1 \mem_reg[637][6]  ( .D(n21004), .CK(clk), .Q(\mem[637][6] ) );
  DFF_X1 \mem_reg[637][5]  ( .D(n21005), .CK(clk), .Q(\mem[637][5] ) );
  DFF_X1 \mem_reg[637][4]  ( .D(n21006), .CK(clk), .Q(\mem[637][4] ) );
  DFF_X1 \mem_reg[637][3]  ( .D(n21007), .CK(clk), .Q(\mem[637][3] ) );
  DFF_X1 \mem_reg[637][2]  ( .D(n21008), .CK(clk), .Q(\mem[637][2] ) );
  DFF_X1 \mem_reg[637][1]  ( .D(n21009), .CK(clk), .Q(\mem[637][1] ) );
  DFF_X1 \mem_reg[637][0]  ( .D(n21010), .CK(clk), .Q(\mem[637][0] ) );
  DFF_X1 \mem_reg[636][7]  ( .D(n21011), .CK(clk), .Q(\mem[636][7] ) );
  DFF_X1 \mem_reg[636][6]  ( .D(n21012), .CK(clk), .Q(\mem[636][6] ) );
  DFF_X1 \mem_reg[636][5]  ( .D(n21013), .CK(clk), .Q(\mem[636][5] ) );
  DFF_X1 \mem_reg[636][4]  ( .D(n21014), .CK(clk), .Q(\mem[636][4] ) );
  DFF_X1 \mem_reg[636][3]  ( .D(n21015), .CK(clk), .Q(\mem[636][3] ) );
  DFF_X1 \mem_reg[636][2]  ( .D(n21016), .CK(clk), .Q(\mem[636][2] ) );
  DFF_X1 \mem_reg[636][1]  ( .D(n21017), .CK(clk), .Q(\mem[636][1] ) );
  DFF_X1 \mem_reg[636][0]  ( .D(n21018), .CK(clk), .Q(\mem[636][0] ) );
  DFF_X1 \mem_reg[635][7]  ( .D(n21019), .CK(clk), .Q(\mem[635][7] ) );
  DFF_X1 \mem_reg[635][6]  ( .D(n21020), .CK(clk), .Q(\mem[635][6] ) );
  DFF_X1 \mem_reg[635][5]  ( .D(n21021), .CK(clk), .Q(\mem[635][5] ) );
  DFF_X1 \mem_reg[635][4]  ( .D(n21022), .CK(clk), .Q(\mem[635][4] ) );
  DFF_X1 \mem_reg[635][3]  ( .D(n21023), .CK(clk), .Q(\mem[635][3] ) );
  DFF_X1 \mem_reg[635][2]  ( .D(n21024), .CK(clk), .Q(\mem[635][2] ) );
  DFF_X1 \mem_reg[635][1]  ( .D(n21025), .CK(clk), .Q(\mem[635][1] ) );
  DFF_X1 \mem_reg[635][0]  ( .D(n21026), .CK(clk), .Q(\mem[635][0] ) );
  DFF_X1 \mem_reg[634][7]  ( .D(n21027), .CK(clk), .Q(\mem[634][7] ) );
  DFF_X1 \mem_reg[634][6]  ( .D(n21028), .CK(clk), .Q(\mem[634][6] ) );
  DFF_X1 \mem_reg[634][5]  ( .D(n21029), .CK(clk), .Q(\mem[634][5] ) );
  DFF_X1 \mem_reg[634][4]  ( .D(n21030), .CK(clk), .Q(\mem[634][4] ) );
  DFF_X1 \mem_reg[634][3]  ( .D(n21031), .CK(clk), .Q(\mem[634][3] ) );
  DFF_X1 \mem_reg[634][2]  ( .D(n21032), .CK(clk), .Q(\mem[634][2] ) );
  DFF_X1 \mem_reg[634][1]  ( .D(n21033), .CK(clk), .Q(\mem[634][1] ) );
  DFF_X1 \mem_reg[634][0]  ( .D(n21034), .CK(clk), .Q(\mem[634][0] ) );
  DFF_X1 \mem_reg[633][7]  ( .D(n21035), .CK(clk), .Q(\mem[633][7] ) );
  DFF_X1 \mem_reg[633][6]  ( .D(n21036), .CK(clk), .Q(\mem[633][6] ) );
  DFF_X1 \mem_reg[633][5]  ( .D(n21037), .CK(clk), .Q(\mem[633][5] ) );
  DFF_X1 \mem_reg[633][4]  ( .D(n21038), .CK(clk), .Q(\mem[633][4] ) );
  DFF_X1 \mem_reg[633][3]  ( .D(n21039), .CK(clk), .Q(\mem[633][3] ) );
  DFF_X1 \mem_reg[633][2]  ( .D(n21040), .CK(clk), .Q(\mem[633][2] ) );
  DFF_X1 \mem_reg[633][1]  ( .D(n21041), .CK(clk), .Q(\mem[633][1] ) );
  DFF_X1 \mem_reg[633][0]  ( .D(n21042), .CK(clk), .Q(\mem[633][0] ) );
  DFF_X1 \mem_reg[632][7]  ( .D(n21043), .CK(clk), .Q(\mem[632][7] ) );
  DFF_X1 \mem_reg[632][6]  ( .D(n21044), .CK(clk), .Q(\mem[632][6] ) );
  DFF_X1 \mem_reg[632][5]  ( .D(n21045), .CK(clk), .Q(\mem[632][5] ) );
  DFF_X1 \mem_reg[632][4]  ( .D(n21046), .CK(clk), .Q(\mem[632][4] ) );
  DFF_X1 \mem_reg[632][3]  ( .D(n21047), .CK(clk), .Q(\mem[632][3] ) );
  DFF_X1 \mem_reg[632][2]  ( .D(n21048), .CK(clk), .Q(\mem[632][2] ) );
  DFF_X1 \mem_reg[632][1]  ( .D(n21049), .CK(clk), .Q(\mem[632][1] ) );
  DFF_X1 \mem_reg[632][0]  ( .D(n21050), .CK(clk), .Q(\mem[632][0] ) );
  DFF_X1 \mem_reg[631][7]  ( .D(n21051), .CK(clk), .Q(\mem[631][7] ) );
  DFF_X1 \mem_reg[631][6]  ( .D(n21052), .CK(clk), .Q(\mem[631][6] ) );
  DFF_X1 \mem_reg[631][5]  ( .D(n21053), .CK(clk), .Q(\mem[631][5] ) );
  DFF_X1 \mem_reg[631][4]  ( .D(n21054), .CK(clk), .Q(\mem[631][4] ) );
  DFF_X1 \mem_reg[631][3]  ( .D(n21055), .CK(clk), .Q(\mem[631][3] ) );
  DFF_X1 \mem_reg[631][2]  ( .D(n21056), .CK(clk), .Q(\mem[631][2] ) );
  DFF_X1 \mem_reg[631][1]  ( .D(n21057), .CK(clk), .Q(\mem[631][1] ) );
  DFF_X1 \mem_reg[631][0]  ( .D(n21058), .CK(clk), .Q(\mem[631][0] ) );
  DFF_X1 \mem_reg[630][7]  ( .D(n21059), .CK(clk), .Q(\mem[630][7] ) );
  DFF_X1 \mem_reg[630][6]  ( .D(n21060), .CK(clk), .Q(\mem[630][6] ) );
  DFF_X1 \mem_reg[630][5]  ( .D(n21061), .CK(clk), .Q(\mem[630][5] ) );
  DFF_X1 \mem_reg[630][4]  ( .D(n21062), .CK(clk), .Q(\mem[630][4] ) );
  DFF_X1 \mem_reg[630][3]  ( .D(n21063), .CK(clk), .Q(\mem[630][3] ) );
  DFF_X1 \mem_reg[630][2]  ( .D(n21064), .CK(clk), .Q(\mem[630][2] ) );
  DFF_X1 \mem_reg[630][1]  ( .D(n21065), .CK(clk), .Q(\mem[630][1] ) );
  DFF_X1 \mem_reg[630][0]  ( .D(n21066), .CK(clk), .Q(\mem[630][0] ) );
  DFF_X1 \mem_reg[629][7]  ( .D(n21067), .CK(clk), .Q(\mem[629][7] ) );
  DFF_X1 \mem_reg[629][6]  ( .D(n21068), .CK(clk), .Q(\mem[629][6] ) );
  DFF_X1 \mem_reg[629][5]  ( .D(n21069), .CK(clk), .Q(\mem[629][5] ) );
  DFF_X1 \mem_reg[629][4]  ( .D(n21070), .CK(clk), .Q(\mem[629][4] ) );
  DFF_X1 \mem_reg[629][3]  ( .D(n21071), .CK(clk), .Q(\mem[629][3] ) );
  DFF_X1 \mem_reg[629][2]  ( .D(n21072), .CK(clk), .Q(\mem[629][2] ) );
  DFF_X1 \mem_reg[629][1]  ( .D(n21073), .CK(clk), .Q(\mem[629][1] ) );
  DFF_X1 \mem_reg[629][0]  ( .D(n21074), .CK(clk), .Q(\mem[629][0] ) );
  DFF_X1 \mem_reg[628][7]  ( .D(n21075), .CK(clk), .Q(\mem[628][7] ) );
  DFF_X1 \mem_reg[628][6]  ( .D(n21076), .CK(clk), .Q(\mem[628][6] ) );
  DFF_X1 \mem_reg[628][5]  ( .D(n21077), .CK(clk), .Q(\mem[628][5] ) );
  DFF_X1 \mem_reg[628][4]  ( .D(n21078), .CK(clk), .Q(\mem[628][4] ) );
  DFF_X1 \mem_reg[628][3]  ( .D(n21079), .CK(clk), .Q(\mem[628][3] ) );
  DFF_X1 \mem_reg[628][2]  ( .D(n21080), .CK(clk), .Q(\mem[628][2] ) );
  DFF_X1 \mem_reg[628][1]  ( .D(n21081), .CK(clk), .Q(\mem[628][1] ) );
  DFF_X1 \mem_reg[628][0]  ( .D(n21082), .CK(clk), .Q(\mem[628][0] ) );
  DFF_X1 \mem_reg[627][7]  ( .D(n21083), .CK(clk), .Q(\mem[627][7] ) );
  DFF_X1 \mem_reg[627][6]  ( .D(n21084), .CK(clk), .Q(\mem[627][6] ) );
  DFF_X1 \mem_reg[627][5]  ( .D(n21085), .CK(clk), .Q(\mem[627][5] ) );
  DFF_X1 \mem_reg[627][4]  ( .D(n21086), .CK(clk), .Q(\mem[627][4] ) );
  DFF_X1 \mem_reg[627][3]  ( .D(n21087), .CK(clk), .Q(\mem[627][3] ) );
  DFF_X1 \mem_reg[627][2]  ( .D(n21088), .CK(clk), .Q(\mem[627][2] ) );
  DFF_X1 \mem_reg[627][1]  ( .D(n21089), .CK(clk), .Q(\mem[627][1] ) );
  DFF_X1 \mem_reg[627][0]  ( .D(n21090), .CK(clk), .Q(\mem[627][0] ) );
  DFF_X1 \mem_reg[626][7]  ( .D(n21091), .CK(clk), .Q(\mem[626][7] ) );
  DFF_X1 \mem_reg[626][6]  ( .D(n21092), .CK(clk), .Q(\mem[626][6] ) );
  DFF_X1 \mem_reg[626][5]  ( .D(n21093), .CK(clk), .Q(\mem[626][5] ) );
  DFF_X1 \mem_reg[626][4]  ( .D(n21094), .CK(clk), .Q(\mem[626][4] ) );
  DFF_X1 \mem_reg[626][3]  ( .D(n21095), .CK(clk), .Q(\mem[626][3] ) );
  DFF_X1 \mem_reg[626][2]  ( .D(n21096), .CK(clk), .Q(\mem[626][2] ) );
  DFF_X1 \mem_reg[626][1]  ( .D(n21097), .CK(clk), .Q(\mem[626][1] ) );
  DFF_X1 \mem_reg[626][0]  ( .D(n21098), .CK(clk), .Q(\mem[626][0] ) );
  DFF_X1 \mem_reg[625][7]  ( .D(n21099), .CK(clk), .Q(\mem[625][7] ) );
  DFF_X1 \mem_reg[625][6]  ( .D(n21100), .CK(clk), .Q(\mem[625][6] ) );
  DFF_X1 \mem_reg[625][5]  ( .D(n21101), .CK(clk), .Q(\mem[625][5] ) );
  DFF_X1 \mem_reg[625][4]  ( .D(n21102), .CK(clk), .Q(\mem[625][4] ) );
  DFF_X1 \mem_reg[625][3]  ( .D(n21103), .CK(clk), .Q(\mem[625][3] ) );
  DFF_X1 \mem_reg[625][2]  ( .D(n21104), .CK(clk), .Q(\mem[625][2] ) );
  DFF_X1 \mem_reg[625][1]  ( .D(n21105), .CK(clk), .Q(\mem[625][1] ) );
  DFF_X1 \mem_reg[625][0]  ( .D(n21106), .CK(clk), .Q(\mem[625][0] ) );
  DFF_X1 \mem_reg[624][7]  ( .D(n21107), .CK(clk), .Q(\mem[624][7] ) );
  DFF_X1 \mem_reg[624][6]  ( .D(n21108), .CK(clk), .Q(\mem[624][6] ) );
  DFF_X1 \mem_reg[624][5]  ( .D(n21109), .CK(clk), .Q(\mem[624][5] ) );
  DFF_X1 \mem_reg[624][4]  ( .D(n21110), .CK(clk), .Q(\mem[624][4] ) );
  DFF_X1 \mem_reg[624][3]  ( .D(n21111), .CK(clk), .Q(\mem[624][3] ) );
  DFF_X1 \mem_reg[624][2]  ( .D(n21112), .CK(clk), .Q(\mem[624][2] ) );
  DFF_X1 \mem_reg[624][1]  ( .D(n21113), .CK(clk), .Q(\mem[624][1] ) );
  DFF_X1 \mem_reg[624][0]  ( .D(n21114), .CK(clk), .Q(\mem[624][0] ) );
  DFF_X1 \mem_reg[623][7]  ( .D(n21115), .CK(clk), .Q(\mem[623][7] ) );
  DFF_X1 \mem_reg[623][6]  ( .D(n21116), .CK(clk), .Q(\mem[623][6] ) );
  DFF_X1 \mem_reg[623][5]  ( .D(n21117), .CK(clk), .Q(\mem[623][5] ) );
  DFF_X1 \mem_reg[623][4]  ( .D(n21118), .CK(clk), .Q(\mem[623][4] ) );
  DFF_X1 \mem_reg[623][3]  ( .D(n21119), .CK(clk), .Q(\mem[623][3] ) );
  DFF_X1 \mem_reg[623][2]  ( .D(n21120), .CK(clk), .Q(\mem[623][2] ) );
  DFF_X1 \mem_reg[623][1]  ( .D(n21121), .CK(clk), .Q(\mem[623][1] ) );
  DFF_X1 \mem_reg[623][0]  ( .D(n21122), .CK(clk), .Q(\mem[623][0] ) );
  DFF_X1 \mem_reg[622][7]  ( .D(n21123), .CK(clk), .Q(\mem[622][7] ) );
  DFF_X1 \mem_reg[622][6]  ( .D(n21124), .CK(clk), .Q(\mem[622][6] ) );
  DFF_X1 \mem_reg[622][5]  ( .D(n21125), .CK(clk), .Q(\mem[622][5] ) );
  DFF_X1 \mem_reg[622][4]  ( .D(n21126), .CK(clk), .Q(\mem[622][4] ) );
  DFF_X1 \mem_reg[622][3]  ( .D(n21127), .CK(clk), .Q(\mem[622][3] ) );
  DFF_X1 \mem_reg[622][2]  ( .D(n21128), .CK(clk), .Q(\mem[622][2] ) );
  DFF_X1 \mem_reg[622][1]  ( .D(n21129), .CK(clk), .Q(\mem[622][1] ) );
  DFF_X1 \mem_reg[622][0]  ( .D(n21130), .CK(clk), .Q(\mem[622][0] ) );
  DFF_X1 \mem_reg[621][7]  ( .D(n21131), .CK(clk), .Q(\mem[621][7] ) );
  DFF_X1 \mem_reg[621][6]  ( .D(n21132), .CK(clk), .Q(\mem[621][6] ) );
  DFF_X1 \mem_reg[621][5]  ( .D(n21133), .CK(clk), .Q(\mem[621][5] ) );
  DFF_X1 \mem_reg[621][4]  ( .D(n21134), .CK(clk), .Q(\mem[621][4] ) );
  DFF_X1 \mem_reg[621][3]  ( .D(n21135), .CK(clk), .Q(\mem[621][3] ) );
  DFF_X1 \mem_reg[621][2]  ( .D(n21136), .CK(clk), .Q(\mem[621][2] ) );
  DFF_X1 \mem_reg[621][1]  ( .D(n21137), .CK(clk), .Q(\mem[621][1] ) );
  DFF_X1 \mem_reg[621][0]  ( .D(n21138), .CK(clk), .Q(\mem[621][0] ) );
  DFF_X1 \mem_reg[620][7]  ( .D(n21139), .CK(clk), .Q(\mem[620][7] ) );
  DFF_X1 \mem_reg[620][6]  ( .D(n21140), .CK(clk), .Q(\mem[620][6] ) );
  DFF_X1 \mem_reg[620][5]  ( .D(n21141), .CK(clk), .Q(\mem[620][5] ) );
  DFF_X1 \mem_reg[620][4]  ( .D(n21142), .CK(clk), .Q(\mem[620][4] ) );
  DFF_X1 \mem_reg[620][3]  ( .D(n21143), .CK(clk), .Q(\mem[620][3] ) );
  DFF_X1 \mem_reg[620][2]  ( .D(n21144), .CK(clk), .Q(\mem[620][2] ) );
  DFF_X1 \mem_reg[620][1]  ( .D(n21145), .CK(clk), .Q(\mem[620][1] ) );
  DFF_X1 \mem_reg[620][0]  ( .D(n21146), .CK(clk), .Q(\mem[620][0] ) );
  DFF_X1 \mem_reg[619][7]  ( .D(n21147), .CK(clk), .Q(\mem[619][7] ) );
  DFF_X1 \mem_reg[619][6]  ( .D(n21148), .CK(clk), .Q(\mem[619][6] ) );
  DFF_X1 \mem_reg[619][5]  ( .D(n21149), .CK(clk), .Q(\mem[619][5] ) );
  DFF_X1 \mem_reg[619][4]  ( .D(n21150), .CK(clk), .Q(\mem[619][4] ) );
  DFF_X1 \mem_reg[619][3]  ( .D(n21151), .CK(clk), .Q(\mem[619][3] ) );
  DFF_X1 \mem_reg[619][2]  ( .D(n21152), .CK(clk), .Q(\mem[619][2] ) );
  DFF_X1 \mem_reg[619][1]  ( .D(n21153), .CK(clk), .Q(\mem[619][1] ) );
  DFF_X1 \mem_reg[619][0]  ( .D(n21154), .CK(clk), .Q(\mem[619][0] ) );
  DFF_X1 \mem_reg[618][7]  ( .D(n21155), .CK(clk), .Q(\mem[618][7] ) );
  DFF_X1 \mem_reg[618][6]  ( .D(n21156), .CK(clk), .Q(\mem[618][6] ) );
  DFF_X1 \mem_reg[618][5]  ( .D(n21157), .CK(clk), .Q(\mem[618][5] ) );
  DFF_X1 \mem_reg[618][4]  ( .D(n21158), .CK(clk), .Q(\mem[618][4] ) );
  DFF_X1 \mem_reg[618][3]  ( .D(n21159), .CK(clk), .Q(\mem[618][3] ) );
  DFF_X1 \mem_reg[618][2]  ( .D(n21160), .CK(clk), .Q(\mem[618][2] ) );
  DFF_X1 \mem_reg[618][1]  ( .D(n21161), .CK(clk), .Q(\mem[618][1] ) );
  DFF_X1 \mem_reg[618][0]  ( .D(n21162), .CK(clk), .Q(\mem[618][0] ) );
  DFF_X1 \mem_reg[617][7]  ( .D(n21163), .CK(clk), .Q(\mem[617][7] ) );
  DFF_X1 \mem_reg[617][6]  ( .D(n21164), .CK(clk), .Q(\mem[617][6] ) );
  DFF_X1 \mem_reg[617][5]  ( .D(n21165), .CK(clk), .Q(\mem[617][5] ) );
  DFF_X1 \mem_reg[617][4]  ( .D(n21166), .CK(clk), .Q(\mem[617][4] ) );
  DFF_X1 \mem_reg[617][3]  ( .D(n21167), .CK(clk), .Q(\mem[617][3] ) );
  DFF_X1 \mem_reg[617][2]  ( .D(n21168), .CK(clk), .Q(\mem[617][2] ) );
  DFF_X1 \mem_reg[617][1]  ( .D(n21169), .CK(clk), .Q(\mem[617][1] ) );
  DFF_X1 \mem_reg[617][0]  ( .D(n21170), .CK(clk), .Q(\mem[617][0] ) );
  DFF_X1 \mem_reg[616][7]  ( .D(n21171), .CK(clk), .Q(\mem[616][7] ) );
  DFF_X1 \mem_reg[616][6]  ( .D(n21172), .CK(clk), .Q(\mem[616][6] ) );
  DFF_X1 \mem_reg[616][5]  ( .D(n21173), .CK(clk), .Q(\mem[616][5] ) );
  DFF_X1 \mem_reg[616][4]  ( .D(n21174), .CK(clk), .Q(\mem[616][4] ) );
  DFF_X1 \mem_reg[616][3]  ( .D(n21175), .CK(clk), .Q(\mem[616][3] ) );
  DFF_X1 \mem_reg[616][2]  ( .D(n21176), .CK(clk), .Q(\mem[616][2] ) );
  DFF_X1 \mem_reg[616][1]  ( .D(n21177), .CK(clk), .Q(\mem[616][1] ) );
  DFF_X1 \mem_reg[616][0]  ( .D(n21178), .CK(clk), .Q(\mem[616][0] ) );
  DFF_X1 \mem_reg[615][7]  ( .D(n21179), .CK(clk), .Q(\mem[615][7] ) );
  DFF_X1 \mem_reg[615][6]  ( .D(n21180), .CK(clk), .Q(\mem[615][6] ) );
  DFF_X1 \mem_reg[615][5]  ( .D(n21181), .CK(clk), .Q(\mem[615][5] ) );
  DFF_X1 \mem_reg[615][4]  ( .D(n21182), .CK(clk), .Q(\mem[615][4] ) );
  DFF_X1 \mem_reg[615][3]  ( .D(n21183), .CK(clk), .Q(\mem[615][3] ) );
  DFF_X1 \mem_reg[615][2]  ( .D(n21184), .CK(clk), .Q(\mem[615][2] ) );
  DFF_X1 \mem_reg[615][1]  ( .D(n21185), .CK(clk), .Q(\mem[615][1] ) );
  DFF_X1 \mem_reg[615][0]  ( .D(n21186), .CK(clk), .Q(\mem[615][0] ) );
  DFF_X1 \mem_reg[614][7]  ( .D(n21187), .CK(clk), .Q(\mem[614][7] ) );
  DFF_X1 \mem_reg[614][6]  ( .D(n21188), .CK(clk), .Q(\mem[614][6] ) );
  DFF_X1 \mem_reg[614][5]  ( .D(n21189), .CK(clk), .Q(\mem[614][5] ) );
  DFF_X1 \mem_reg[614][4]  ( .D(n21190), .CK(clk), .Q(\mem[614][4] ) );
  DFF_X1 \mem_reg[614][3]  ( .D(n21191), .CK(clk), .Q(\mem[614][3] ) );
  DFF_X1 \mem_reg[614][2]  ( .D(n21192), .CK(clk), .Q(\mem[614][2] ) );
  DFF_X1 \mem_reg[614][1]  ( .D(n21193), .CK(clk), .Q(\mem[614][1] ) );
  DFF_X1 \mem_reg[614][0]  ( .D(n21194), .CK(clk), .Q(\mem[614][0] ) );
  DFF_X1 \mem_reg[613][7]  ( .D(n21195), .CK(clk), .Q(\mem[613][7] ) );
  DFF_X1 \mem_reg[613][6]  ( .D(n21196), .CK(clk), .Q(\mem[613][6] ) );
  DFF_X1 \mem_reg[613][5]  ( .D(n21197), .CK(clk), .Q(\mem[613][5] ) );
  DFF_X1 \mem_reg[613][4]  ( .D(n21198), .CK(clk), .Q(\mem[613][4] ) );
  DFF_X1 \mem_reg[613][3]  ( .D(n21199), .CK(clk), .Q(\mem[613][3] ) );
  DFF_X1 \mem_reg[613][2]  ( .D(n21200), .CK(clk), .Q(\mem[613][2] ) );
  DFF_X1 \mem_reg[613][1]  ( .D(n21201), .CK(clk), .Q(\mem[613][1] ) );
  DFF_X1 \mem_reg[613][0]  ( .D(n21202), .CK(clk), .Q(\mem[613][0] ) );
  DFF_X1 \mem_reg[612][7]  ( .D(n21203), .CK(clk), .Q(\mem[612][7] ) );
  DFF_X1 \mem_reg[612][6]  ( .D(n21204), .CK(clk), .Q(\mem[612][6] ) );
  DFF_X1 \mem_reg[612][5]  ( .D(n21205), .CK(clk), .Q(\mem[612][5] ) );
  DFF_X1 \mem_reg[612][4]  ( .D(n21206), .CK(clk), .Q(\mem[612][4] ) );
  DFF_X1 \mem_reg[612][3]  ( .D(n21207), .CK(clk), .Q(\mem[612][3] ) );
  DFF_X1 \mem_reg[612][2]  ( .D(n21208), .CK(clk), .Q(\mem[612][2] ) );
  DFF_X1 \mem_reg[612][1]  ( .D(n21209), .CK(clk), .Q(\mem[612][1] ) );
  DFF_X1 \mem_reg[612][0]  ( .D(n21210), .CK(clk), .Q(\mem[612][0] ) );
  DFF_X1 \mem_reg[611][7]  ( .D(n21211), .CK(clk), .Q(\mem[611][7] ) );
  DFF_X1 \mem_reg[611][6]  ( .D(n21212), .CK(clk), .Q(\mem[611][6] ) );
  DFF_X1 \mem_reg[611][5]  ( .D(n21213), .CK(clk), .Q(\mem[611][5] ) );
  DFF_X1 \mem_reg[611][4]  ( .D(n21214), .CK(clk), .Q(\mem[611][4] ) );
  DFF_X1 \mem_reg[611][3]  ( .D(n21215), .CK(clk), .Q(\mem[611][3] ) );
  DFF_X1 \mem_reg[611][2]  ( .D(n21216), .CK(clk), .Q(\mem[611][2] ) );
  DFF_X1 \mem_reg[611][1]  ( .D(n21217), .CK(clk), .Q(\mem[611][1] ) );
  DFF_X1 \mem_reg[611][0]  ( .D(n21218), .CK(clk), .Q(\mem[611][0] ) );
  DFF_X1 \mem_reg[610][7]  ( .D(n21219), .CK(clk), .Q(\mem[610][7] ) );
  DFF_X1 \mem_reg[610][6]  ( .D(n21220), .CK(clk), .Q(\mem[610][6] ) );
  DFF_X1 \mem_reg[610][5]  ( .D(n21221), .CK(clk), .Q(\mem[610][5] ) );
  DFF_X1 \mem_reg[610][4]  ( .D(n21222), .CK(clk), .Q(\mem[610][4] ) );
  DFF_X1 \mem_reg[610][3]  ( .D(n21223), .CK(clk), .Q(\mem[610][3] ) );
  DFF_X1 \mem_reg[610][2]  ( .D(n21224), .CK(clk), .Q(\mem[610][2] ) );
  DFF_X1 \mem_reg[610][1]  ( .D(n21225), .CK(clk), .Q(\mem[610][1] ) );
  DFF_X1 \mem_reg[610][0]  ( .D(n21226), .CK(clk), .Q(\mem[610][0] ) );
  DFF_X1 \mem_reg[609][7]  ( .D(n21227), .CK(clk), .Q(\mem[609][7] ) );
  DFF_X1 \mem_reg[609][6]  ( .D(n21228), .CK(clk), .Q(\mem[609][6] ) );
  DFF_X1 \mem_reg[609][5]  ( .D(n21229), .CK(clk), .Q(\mem[609][5] ) );
  DFF_X1 \mem_reg[609][4]  ( .D(n21230), .CK(clk), .Q(\mem[609][4] ) );
  DFF_X1 \mem_reg[609][3]  ( .D(n21231), .CK(clk), .Q(\mem[609][3] ) );
  DFF_X1 \mem_reg[609][2]  ( .D(n21232), .CK(clk), .Q(\mem[609][2] ) );
  DFF_X1 \mem_reg[609][1]  ( .D(n21233), .CK(clk), .Q(\mem[609][1] ) );
  DFF_X1 \mem_reg[609][0]  ( .D(n21234), .CK(clk), .Q(\mem[609][0] ) );
  DFF_X1 \mem_reg[608][7]  ( .D(n21235), .CK(clk), .Q(\mem[608][7] ) );
  DFF_X1 \mem_reg[608][6]  ( .D(n21236), .CK(clk), .Q(\mem[608][6] ) );
  DFF_X1 \mem_reg[608][5]  ( .D(n21237), .CK(clk), .Q(\mem[608][5] ) );
  DFF_X1 \mem_reg[608][4]  ( .D(n21238), .CK(clk), .Q(\mem[608][4] ) );
  DFF_X1 \mem_reg[608][3]  ( .D(n21239), .CK(clk), .Q(\mem[608][3] ) );
  DFF_X1 \mem_reg[608][2]  ( .D(n21240), .CK(clk), .Q(\mem[608][2] ) );
  DFF_X1 \mem_reg[608][1]  ( .D(n21241), .CK(clk), .Q(\mem[608][1] ) );
  DFF_X1 \mem_reg[608][0]  ( .D(n21242), .CK(clk), .Q(\mem[608][0] ) );
  DFF_X1 \mem_reg[607][7]  ( .D(n21243), .CK(clk), .Q(\mem[607][7] ) );
  DFF_X1 \mem_reg[607][6]  ( .D(n21244), .CK(clk), .Q(\mem[607][6] ) );
  DFF_X1 \mem_reg[607][5]  ( .D(n21245), .CK(clk), .Q(\mem[607][5] ) );
  DFF_X1 \mem_reg[607][4]  ( .D(n21246), .CK(clk), .Q(\mem[607][4] ) );
  DFF_X1 \mem_reg[607][3]  ( .D(n21247), .CK(clk), .Q(\mem[607][3] ) );
  DFF_X1 \mem_reg[607][2]  ( .D(n21248), .CK(clk), .Q(\mem[607][2] ) );
  DFF_X1 \mem_reg[607][1]  ( .D(n21249), .CK(clk), .Q(\mem[607][1] ) );
  DFF_X1 \mem_reg[607][0]  ( .D(n21250), .CK(clk), .Q(\mem[607][0] ) );
  DFF_X1 \mem_reg[606][7]  ( .D(n21251), .CK(clk), .Q(\mem[606][7] ) );
  DFF_X1 \mem_reg[606][6]  ( .D(n21252), .CK(clk), .Q(\mem[606][6] ) );
  DFF_X1 \mem_reg[606][5]  ( .D(n21253), .CK(clk), .Q(\mem[606][5] ) );
  DFF_X1 \mem_reg[606][4]  ( .D(n21254), .CK(clk), .Q(\mem[606][4] ) );
  DFF_X1 \mem_reg[606][3]  ( .D(n21255), .CK(clk), .Q(\mem[606][3] ) );
  DFF_X1 \mem_reg[606][2]  ( .D(n21256), .CK(clk), .Q(\mem[606][2] ) );
  DFF_X1 \mem_reg[606][1]  ( .D(n21257), .CK(clk), .Q(\mem[606][1] ) );
  DFF_X1 \mem_reg[606][0]  ( .D(n21258), .CK(clk), .Q(\mem[606][0] ) );
  DFF_X1 \mem_reg[605][7]  ( .D(n21259), .CK(clk), .Q(\mem[605][7] ) );
  DFF_X1 \mem_reg[605][6]  ( .D(n21260), .CK(clk), .Q(\mem[605][6] ) );
  DFF_X1 \mem_reg[605][5]  ( .D(n21261), .CK(clk), .Q(\mem[605][5] ) );
  DFF_X1 \mem_reg[605][4]  ( .D(n21262), .CK(clk), .Q(\mem[605][4] ) );
  DFF_X1 \mem_reg[605][3]  ( .D(n21263), .CK(clk), .Q(\mem[605][3] ) );
  DFF_X1 \mem_reg[605][2]  ( .D(n21264), .CK(clk), .Q(\mem[605][2] ) );
  DFF_X1 \mem_reg[605][1]  ( .D(n21265), .CK(clk), .Q(\mem[605][1] ) );
  DFF_X1 \mem_reg[605][0]  ( .D(n21266), .CK(clk), .Q(\mem[605][0] ) );
  DFF_X1 \mem_reg[604][7]  ( .D(n21267), .CK(clk), .Q(\mem[604][7] ) );
  DFF_X1 \mem_reg[604][6]  ( .D(n21268), .CK(clk), .Q(\mem[604][6] ) );
  DFF_X1 \mem_reg[604][5]  ( .D(n21269), .CK(clk), .Q(\mem[604][5] ) );
  DFF_X1 \mem_reg[604][4]  ( .D(n21270), .CK(clk), .Q(\mem[604][4] ) );
  DFF_X1 \mem_reg[604][3]  ( .D(n21271), .CK(clk), .Q(\mem[604][3] ) );
  DFF_X1 \mem_reg[604][2]  ( .D(n21272), .CK(clk), .Q(\mem[604][2] ) );
  DFF_X1 \mem_reg[604][1]  ( .D(n21273), .CK(clk), .Q(\mem[604][1] ) );
  DFF_X1 \mem_reg[604][0]  ( .D(n21274), .CK(clk), .Q(\mem[604][0] ) );
  DFF_X1 \mem_reg[603][7]  ( .D(n21275), .CK(clk), .Q(\mem[603][7] ) );
  DFF_X1 \mem_reg[603][6]  ( .D(n21276), .CK(clk), .Q(\mem[603][6] ) );
  DFF_X1 \mem_reg[603][5]  ( .D(n21277), .CK(clk), .Q(\mem[603][5] ) );
  DFF_X1 \mem_reg[603][4]  ( .D(n21278), .CK(clk), .Q(\mem[603][4] ) );
  DFF_X1 \mem_reg[603][3]  ( .D(n21279), .CK(clk), .Q(\mem[603][3] ) );
  DFF_X1 \mem_reg[603][2]  ( .D(n21280), .CK(clk), .Q(\mem[603][2] ) );
  DFF_X1 \mem_reg[603][1]  ( .D(n21281), .CK(clk), .Q(\mem[603][1] ) );
  DFF_X1 \mem_reg[603][0]  ( .D(n21282), .CK(clk), .Q(\mem[603][0] ) );
  DFF_X1 \mem_reg[602][7]  ( .D(n21283), .CK(clk), .Q(\mem[602][7] ) );
  DFF_X1 \mem_reg[602][6]  ( .D(n21284), .CK(clk), .Q(\mem[602][6] ) );
  DFF_X1 \mem_reg[602][5]  ( .D(n21285), .CK(clk), .Q(\mem[602][5] ) );
  DFF_X1 \mem_reg[602][4]  ( .D(n21286), .CK(clk), .Q(\mem[602][4] ) );
  DFF_X1 \mem_reg[602][3]  ( .D(n21287), .CK(clk), .Q(\mem[602][3] ) );
  DFF_X1 \mem_reg[602][2]  ( .D(n21288), .CK(clk), .Q(\mem[602][2] ) );
  DFF_X1 \mem_reg[602][1]  ( .D(n21289), .CK(clk), .Q(\mem[602][1] ) );
  DFF_X1 \mem_reg[602][0]  ( .D(n21290), .CK(clk), .Q(\mem[602][0] ) );
  DFF_X1 \mem_reg[601][7]  ( .D(n21291), .CK(clk), .Q(\mem[601][7] ) );
  DFF_X1 \mem_reg[601][6]  ( .D(n21292), .CK(clk), .Q(\mem[601][6] ) );
  DFF_X1 \mem_reg[601][5]  ( .D(n21293), .CK(clk), .Q(\mem[601][5] ) );
  DFF_X1 \mem_reg[601][4]  ( .D(n21294), .CK(clk), .Q(\mem[601][4] ) );
  DFF_X1 \mem_reg[601][3]  ( .D(n21295), .CK(clk), .Q(\mem[601][3] ) );
  DFF_X1 \mem_reg[601][2]  ( .D(n21296), .CK(clk), .Q(\mem[601][2] ) );
  DFF_X1 \mem_reg[601][1]  ( .D(n21297), .CK(clk), .Q(\mem[601][1] ) );
  DFF_X1 \mem_reg[601][0]  ( .D(n21298), .CK(clk), .Q(\mem[601][0] ) );
  DFF_X1 \mem_reg[600][7]  ( .D(n21299), .CK(clk), .Q(\mem[600][7] ) );
  DFF_X1 \mem_reg[600][6]  ( .D(n21300), .CK(clk), .Q(\mem[600][6] ) );
  DFF_X1 \mem_reg[600][5]  ( .D(n21301), .CK(clk), .Q(\mem[600][5] ) );
  DFF_X1 \mem_reg[600][4]  ( .D(n21302), .CK(clk), .Q(\mem[600][4] ) );
  DFF_X1 \mem_reg[600][3]  ( .D(n21303), .CK(clk), .Q(\mem[600][3] ) );
  DFF_X1 \mem_reg[600][2]  ( .D(n21304), .CK(clk), .Q(\mem[600][2] ) );
  DFF_X1 \mem_reg[600][1]  ( .D(n21305), .CK(clk), .Q(\mem[600][1] ) );
  DFF_X1 \mem_reg[600][0]  ( .D(n21306), .CK(clk), .Q(\mem[600][0] ) );
  DFF_X1 \mem_reg[599][7]  ( .D(n21307), .CK(clk), .Q(\mem[599][7] ) );
  DFF_X1 \mem_reg[599][6]  ( .D(n21308), .CK(clk), .Q(\mem[599][6] ) );
  DFF_X1 \mem_reg[599][5]  ( .D(n21309), .CK(clk), .Q(\mem[599][5] ) );
  DFF_X1 \mem_reg[599][4]  ( .D(n21310), .CK(clk), .Q(\mem[599][4] ) );
  DFF_X1 \mem_reg[599][3]  ( .D(n21311), .CK(clk), .Q(\mem[599][3] ) );
  DFF_X1 \mem_reg[599][2]  ( .D(n21312), .CK(clk), .Q(\mem[599][2] ) );
  DFF_X1 \mem_reg[599][1]  ( .D(n21313), .CK(clk), .Q(\mem[599][1] ) );
  DFF_X1 \mem_reg[599][0]  ( .D(n21314), .CK(clk), .Q(\mem[599][0] ) );
  DFF_X1 \mem_reg[598][7]  ( .D(n21315), .CK(clk), .Q(\mem[598][7] ) );
  DFF_X1 \mem_reg[598][6]  ( .D(n21316), .CK(clk), .Q(\mem[598][6] ) );
  DFF_X1 \mem_reg[598][5]  ( .D(n21317), .CK(clk), .Q(\mem[598][5] ) );
  DFF_X1 \mem_reg[598][4]  ( .D(n21318), .CK(clk), .Q(\mem[598][4] ) );
  DFF_X1 \mem_reg[598][3]  ( .D(n21319), .CK(clk), .Q(\mem[598][3] ) );
  DFF_X1 \mem_reg[598][2]  ( .D(n21320), .CK(clk), .Q(\mem[598][2] ) );
  DFF_X1 \mem_reg[598][1]  ( .D(n21321), .CK(clk), .Q(\mem[598][1] ) );
  DFF_X1 \mem_reg[598][0]  ( .D(n21322), .CK(clk), .Q(\mem[598][0] ) );
  DFF_X1 \mem_reg[597][7]  ( .D(n21323), .CK(clk), .Q(\mem[597][7] ) );
  DFF_X1 \mem_reg[597][6]  ( .D(n21324), .CK(clk), .Q(\mem[597][6] ) );
  DFF_X1 \mem_reg[597][5]  ( .D(n21325), .CK(clk), .Q(\mem[597][5] ) );
  DFF_X1 \mem_reg[597][4]  ( .D(n21326), .CK(clk), .Q(\mem[597][4] ) );
  DFF_X1 \mem_reg[597][3]  ( .D(n21327), .CK(clk), .Q(\mem[597][3] ) );
  DFF_X1 \mem_reg[597][2]  ( .D(n21328), .CK(clk), .Q(\mem[597][2] ) );
  DFF_X1 \mem_reg[597][1]  ( .D(n21329), .CK(clk), .Q(\mem[597][1] ) );
  DFF_X1 \mem_reg[597][0]  ( .D(n21330), .CK(clk), .Q(\mem[597][0] ) );
  DFF_X1 \mem_reg[596][7]  ( .D(n21331), .CK(clk), .Q(\mem[596][7] ) );
  DFF_X1 \mem_reg[596][6]  ( .D(n21332), .CK(clk), .Q(\mem[596][6] ) );
  DFF_X1 \mem_reg[596][5]  ( .D(n21333), .CK(clk), .Q(\mem[596][5] ) );
  DFF_X1 \mem_reg[596][4]  ( .D(n21334), .CK(clk), .Q(\mem[596][4] ) );
  DFF_X1 \mem_reg[596][3]  ( .D(n21335), .CK(clk), .Q(\mem[596][3] ) );
  DFF_X1 \mem_reg[596][2]  ( .D(n21336), .CK(clk), .Q(\mem[596][2] ) );
  DFF_X1 \mem_reg[596][1]  ( .D(n21337), .CK(clk), .Q(\mem[596][1] ) );
  DFF_X1 \mem_reg[596][0]  ( .D(n21338), .CK(clk), .Q(\mem[596][0] ) );
  DFF_X1 \mem_reg[595][7]  ( .D(n21339), .CK(clk), .Q(\mem[595][7] ) );
  DFF_X1 \mem_reg[595][6]  ( .D(n21340), .CK(clk), .Q(\mem[595][6] ) );
  DFF_X1 \mem_reg[595][5]  ( .D(n21341), .CK(clk), .Q(\mem[595][5] ) );
  DFF_X1 \mem_reg[595][4]  ( .D(n21342), .CK(clk), .Q(\mem[595][4] ) );
  DFF_X1 \mem_reg[595][3]  ( .D(n21343), .CK(clk), .Q(\mem[595][3] ) );
  DFF_X1 \mem_reg[595][2]  ( .D(n21344), .CK(clk), .Q(\mem[595][2] ) );
  DFF_X1 \mem_reg[595][1]  ( .D(n21345), .CK(clk), .Q(\mem[595][1] ) );
  DFF_X1 \mem_reg[595][0]  ( .D(n21346), .CK(clk), .Q(\mem[595][0] ) );
  DFF_X1 \mem_reg[594][7]  ( .D(n21347), .CK(clk), .Q(\mem[594][7] ) );
  DFF_X1 \mem_reg[594][6]  ( .D(n21348), .CK(clk), .Q(\mem[594][6] ) );
  DFF_X1 \mem_reg[594][5]  ( .D(n21349), .CK(clk), .Q(\mem[594][5] ) );
  DFF_X1 \mem_reg[594][4]  ( .D(n21350), .CK(clk), .Q(\mem[594][4] ) );
  DFF_X1 \mem_reg[594][3]  ( .D(n21351), .CK(clk), .Q(\mem[594][3] ) );
  DFF_X1 \mem_reg[594][2]  ( .D(n21352), .CK(clk), .Q(\mem[594][2] ) );
  DFF_X1 \mem_reg[594][1]  ( .D(n21353), .CK(clk), .Q(\mem[594][1] ) );
  DFF_X1 \mem_reg[594][0]  ( .D(n21354), .CK(clk), .Q(\mem[594][0] ) );
  DFF_X1 \mem_reg[593][7]  ( .D(n21355), .CK(clk), .Q(\mem[593][7] ) );
  DFF_X1 \mem_reg[593][6]  ( .D(n21356), .CK(clk), .Q(\mem[593][6] ) );
  DFF_X1 \mem_reg[593][5]  ( .D(n21357), .CK(clk), .Q(\mem[593][5] ) );
  DFF_X1 \mem_reg[593][4]  ( .D(n21358), .CK(clk), .Q(\mem[593][4] ) );
  DFF_X1 \mem_reg[593][3]  ( .D(n21359), .CK(clk), .Q(\mem[593][3] ) );
  DFF_X1 \mem_reg[593][2]  ( .D(n21360), .CK(clk), .Q(\mem[593][2] ) );
  DFF_X1 \mem_reg[593][1]  ( .D(n21361), .CK(clk), .Q(\mem[593][1] ) );
  DFF_X1 \mem_reg[593][0]  ( .D(n21362), .CK(clk), .Q(\mem[593][0] ) );
  DFF_X1 \mem_reg[592][7]  ( .D(n21363), .CK(clk), .Q(\mem[592][7] ) );
  DFF_X1 \mem_reg[592][6]  ( .D(n21364), .CK(clk), .Q(\mem[592][6] ) );
  DFF_X1 \mem_reg[592][5]  ( .D(n21365), .CK(clk), .Q(\mem[592][5] ) );
  DFF_X1 \mem_reg[592][4]  ( .D(n21366), .CK(clk), .Q(\mem[592][4] ) );
  DFF_X1 \mem_reg[592][3]  ( .D(n21367), .CK(clk), .Q(\mem[592][3] ) );
  DFF_X1 \mem_reg[592][2]  ( .D(n21368), .CK(clk), .Q(\mem[592][2] ) );
  DFF_X1 \mem_reg[592][1]  ( .D(n21369), .CK(clk), .Q(\mem[592][1] ) );
  DFF_X1 \mem_reg[592][0]  ( .D(n21370), .CK(clk), .Q(\mem[592][0] ) );
  DFF_X1 \mem_reg[591][7]  ( .D(n21371), .CK(clk), .Q(\mem[591][7] ) );
  DFF_X1 \mem_reg[591][6]  ( .D(n21372), .CK(clk), .Q(\mem[591][6] ) );
  DFF_X1 \mem_reg[591][5]  ( .D(n21373), .CK(clk), .Q(\mem[591][5] ) );
  DFF_X1 \mem_reg[591][4]  ( .D(n21374), .CK(clk), .Q(\mem[591][4] ) );
  DFF_X1 \mem_reg[591][3]  ( .D(n21375), .CK(clk), .Q(\mem[591][3] ) );
  DFF_X1 \mem_reg[591][2]  ( .D(n21376), .CK(clk), .Q(\mem[591][2] ) );
  DFF_X1 \mem_reg[591][1]  ( .D(n21377), .CK(clk), .Q(\mem[591][1] ) );
  DFF_X1 \mem_reg[591][0]  ( .D(n21378), .CK(clk), .Q(\mem[591][0] ) );
  DFF_X1 \mem_reg[590][7]  ( .D(n21379), .CK(clk), .Q(\mem[590][7] ) );
  DFF_X1 \mem_reg[590][6]  ( .D(n21380), .CK(clk), .Q(\mem[590][6] ) );
  DFF_X1 \mem_reg[590][5]  ( .D(n21381), .CK(clk), .Q(\mem[590][5] ) );
  DFF_X1 \mem_reg[590][4]  ( .D(n21382), .CK(clk), .Q(\mem[590][4] ) );
  DFF_X1 \mem_reg[590][3]  ( .D(n21383), .CK(clk), .Q(\mem[590][3] ) );
  DFF_X1 \mem_reg[590][2]  ( .D(n21384), .CK(clk), .Q(\mem[590][2] ) );
  DFF_X1 \mem_reg[590][1]  ( .D(n21385), .CK(clk), .Q(\mem[590][1] ) );
  DFF_X1 \mem_reg[590][0]  ( .D(n21386), .CK(clk), .Q(\mem[590][0] ) );
  DFF_X1 \mem_reg[589][7]  ( .D(n21387), .CK(clk), .Q(\mem[589][7] ) );
  DFF_X1 \mem_reg[589][6]  ( .D(n21388), .CK(clk), .Q(\mem[589][6] ) );
  DFF_X1 \mem_reg[589][5]  ( .D(n21389), .CK(clk), .Q(\mem[589][5] ) );
  DFF_X1 \mem_reg[589][4]  ( .D(n21390), .CK(clk), .Q(\mem[589][4] ) );
  DFF_X1 \mem_reg[589][3]  ( .D(n21391), .CK(clk), .Q(\mem[589][3] ) );
  DFF_X1 \mem_reg[589][2]  ( .D(n21392), .CK(clk), .Q(\mem[589][2] ) );
  DFF_X1 \mem_reg[589][1]  ( .D(n21393), .CK(clk), .Q(\mem[589][1] ) );
  DFF_X1 \mem_reg[589][0]  ( .D(n21394), .CK(clk), .Q(\mem[589][0] ) );
  DFF_X1 \mem_reg[588][7]  ( .D(n21395), .CK(clk), .Q(\mem[588][7] ) );
  DFF_X1 \mem_reg[588][6]  ( .D(n21396), .CK(clk), .Q(\mem[588][6] ) );
  DFF_X1 \mem_reg[588][5]  ( .D(n21397), .CK(clk), .Q(\mem[588][5] ) );
  DFF_X1 \mem_reg[588][4]  ( .D(n21398), .CK(clk), .Q(\mem[588][4] ) );
  DFF_X1 \mem_reg[588][3]  ( .D(n21399), .CK(clk), .Q(\mem[588][3] ) );
  DFF_X1 \mem_reg[588][2]  ( .D(n21400), .CK(clk), .Q(\mem[588][2] ) );
  DFF_X1 \mem_reg[588][1]  ( .D(n21401), .CK(clk), .Q(\mem[588][1] ) );
  DFF_X1 \mem_reg[588][0]  ( .D(n21402), .CK(clk), .Q(\mem[588][0] ) );
  DFF_X1 \mem_reg[587][7]  ( .D(n21403), .CK(clk), .Q(\mem[587][7] ) );
  DFF_X1 \mem_reg[587][6]  ( .D(n21404), .CK(clk), .Q(\mem[587][6] ) );
  DFF_X1 \mem_reg[587][5]  ( .D(n21405), .CK(clk), .Q(\mem[587][5] ) );
  DFF_X1 \mem_reg[587][4]  ( .D(n21406), .CK(clk), .Q(\mem[587][4] ) );
  DFF_X1 \mem_reg[587][3]  ( .D(n21407), .CK(clk), .Q(\mem[587][3] ) );
  DFF_X1 \mem_reg[587][2]  ( .D(n21408), .CK(clk), .Q(\mem[587][2] ) );
  DFF_X1 \mem_reg[587][1]  ( .D(n21409), .CK(clk), .Q(\mem[587][1] ) );
  DFF_X1 \mem_reg[587][0]  ( .D(n21410), .CK(clk), .Q(\mem[587][0] ) );
  DFF_X1 \mem_reg[586][7]  ( .D(n21411), .CK(clk), .Q(\mem[586][7] ) );
  DFF_X1 \mem_reg[586][6]  ( .D(n21412), .CK(clk), .Q(\mem[586][6] ) );
  DFF_X1 \mem_reg[586][5]  ( .D(n21413), .CK(clk), .Q(\mem[586][5] ) );
  DFF_X1 \mem_reg[586][4]  ( .D(n21414), .CK(clk), .Q(\mem[586][4] ) );
  DFF_X1 \mem_reg[586][3]  ( .D(n21415), .CK(clk), .Q(\mem[586][3] ) );
  DFF_X1 \mem_reg[586][2]  ( .D(n21416), .CK(clk), .Q(\mem[586][2] ) );
  DFF_X1 \mem_reg[586][1]  ( .D(n21417), .CK(clk), .Q(\mem[586][1] ) );
  DFF_X1 \mem_reg[586][0]  ( .D(n21418), .CK(clk), .Q(\mem[586][0] ) );
  DFF_X1 \mem_reg[585][7]  ( .D(n21419), .CK(clk), .Q(\mem[585][7] ) );
  DFF_X1 \mem_reg[585][6]  ( .D(n21420), .CK(clk), .Q(\mem[585][6] ) );
  DFF_X1 \mem_reg[585][5]  ( .D(n21421), .CK(clk), .Q(\mem[585][5] ) );
  DFF_X1 \mem_reg[585][4]  ( .D(n21422), .CK(clk), .Q(\mem[585][4] ) );
  DFF_X1 \mem_reg[585][3]  ( .D(n21423), .CK(clk), .Q(\mem[585][3] ) );
  DFF_X1 \mem_reg[585][2]  ( .D(n21424), .CK(clk), .Q(\mem[585][2] ) );
  DFF_X1 \mem_reg[585][1]  ( .D(n21425), .CK(clk), .Q(\mem[585][1] ) );
  DFF_X1 \mem_reg[585][0]  ( .D(n21426), .CK(clk), .Q(\mem[585][0] ) );
  DFF_X1 \mem_reg[584][7]  ( .D(n21427), .CK(clk), .Q(\mem[584][7] ) );
  DFF_X1 \mem_reg[584][6]  ( .D(n21428), .CK(clk), .Q(\mem[584][6] ) );
  DFF_X1 \mem_reg[584][5]  ( .D(n21429), .CK(clk), .Q(\mem[584][5] ) );
  DFF_X1 \mem_reg[584][4]  ( .D(n21430), .CK(clk), .Q(\mem[584][4] ) );
  DFF_X1 \mem_reg[584][3]  ( .D(n21431), .CK(clk), .Q(\mem[584][3] ) );
  DFF_X1 \mem_reg[584][2]  ( .D(n21432), .CK(clk), .Q(\mem[584][2] ) );
  DFF_X1 \mem_reg[584][1]  ( .D(n21433), .CK(clk), .Q(\mem[584][1] ) );
  DFF_X1 \mem_reg[584][0]  ( .D(n21434), .CK(clk), .Q(\mem[584][0] ) );
  DFF_X1 \mem_reg[583][7]  ( .D(n21435), .CK(clk), .Q(\mem[583][7] ) );
  DFF_X1 \mem_reg[583][6]  ( .D(n21436), .CK(clk), .Q(\mem[583][6] ) );
  DFF_X1 \mem_reg[583][5]  ( .D(n21437), .CK(clk), .Q(\mem[583][5] ) );
  DFF_X1 \mem_reg[583][4]  ( .D(n21438), .CK(clk), .Q(\mem[583][4] ) );
  DFF_X1 \mem_reg[583][3]  ( .D(n21439), .CK(clk), .Q(\mem[583][3] ) );
  DFF_X1 \mem_reg[583][2]  ( .D(n21440), .CK(clk), .Q(\mem[583][2] ) );
  DFF_X1 \mem_reg[583][1]  ( .D(n21441), .CK(clk), .Q(\mem[583][1] ) );
  DFF_X1 \mem_reg[583][0]  ( .D(n21442), .CK(clk), .Q(\mem[583][0] ) );
  DFF_X1 \mem_reg[582][7]  ( .D(n21443), .CK(clk), .Q(\mem[582][7] ) );
  DFF_X1 \mem_reg[582][6]  ( .D(n21444), .CK(clk), .Q(\mem[582][6] ) );
  DFF_X1 \mem_reg[582][5]  ( .D(n21445), .CK(clk), .Q(\mem[582][5] ) );
  DFF_X1 \mem_reg[582][4]  ( .D(n21446), .CK(clk), .Q(\mem[582][4] ) );
  DFF_X1 \mem_reg[582][3]  ( .D(n21447), .CK(clk), .Q(\mem[582][3] ) );
  DFF_X1 \mem_reg[582][2]  ( .D(n21448), .CK(clk), .Q(\mem[582][2] ) );
  DFF_X1 \mem_reg[582][1]  ( .D(n21449), .CK(clk), .Q(\mem[582][1] ) );
  DFF_X1 \mem_reg[582][0]  ( .D(n21450), .CK(clk), .Q(\mem[582][0] ) );
  DFF_X1 \mem_reg[581][7]  ( .D(n21451), .CK(clk), .Q(\mem[581][7] ) );
  DFF_X1 \mem_reg[581][6]  ( .D(n21452), .CK(clk), .Q(\mem[581][6] ) );
  DFF_X1 \mem_reg[581][5]  ( .D(n21453), .CK(clk), .Q(\mem[581][5] ) );
  DFF_X1 \mem_reg[581][4]  ( .D(n21454), .CK(clk), .Q(\mem[581][4] ) );
  DFF_X1 \mem_reg[581][3]  ( .D(n21455), .CK(clk), .Q(\mem[581][3] ) );
  DFF_X1 \mem_reg[581][2]  ( .D(n21456), .CK(clk), .Q(\mem[581][2] ) );
  DFF_X1 \mem_reg[581][1]  ( .D(n21457), .CK(clk), .Q(\mem[581][1] ) );
  DFF_X1 \mem_reg[581][0]  ( .D(n21458), .CK(clk), .Q(\mem[581][0] ) );
  DFF_X1 \mem_reg[580][7]  ( .D(n21459), .CK(clk), .Q(\mem[580][7] ) );
  DFF_X1 \mem_reg[580][6]  ( .D(n21460), .CK(clk), .Q(\mem[580][6] ) );
  DFF_X1 \mem_reg[580][5]  ( .D(n21461), .CK(clk), .Q(\mem[580][5] ) );
  DFF_X1 \mem_reg[580][4]  ( .D(n21462), .CK(clk), .Q(\mem[580][4] ) );
  DFF_X1 \mem_reg[580][3]  ( .D(n21463), .CK(clk), .Q(\mem[580][3] ) );
  DFF_X1 \mem_reg[580][2]  ( .D(n21464), .CK(clk), .Q(\mem[580][2] ) );
  DFF_X1 \mem_reg[580][1]  ( .D(n21465), .CK(clk), .Q(\mem[580][1] ) );
  DFF_X1 \mem_reg[580][0]  ( .D(n21466), .CK(clk), .Q(\mem[580][0] ) );
  DFF_X1 \mem_reg[579][7]  ( .D(n21467), .CK(clk), .Q(\mem[579][7] ) );
  DFF_X1 \mem_reg[579][6]  ( .D(n21468), .CK(clk), .Q(\mem[579][6] ) );
  DFF_X1 \mem_reg[579][5]  ( .D(n21469), .CK(clk), .Q(\mem[579][5] ) );
  DFF_X1 \mem_reg[579][4]  ( .D(n21470), .CK(clk), .Q(\mem[579][4] ) );
  DFF_X1 \mem_reg[579][3]  ( .D(n21471), .CK(clk), .Q(\mem[579][3] ) );
  DFF_X1 \mem_reg[579][2]  ( .D(n21472), .CK(clk), .Q(\mem[579][2] ) );
  DFF_X1 \mem_reg[579][1]  ( .D(n21473), .CK(clk), .Q(\mem[579][1] ) );
  DFF_X1 \mem_reg[579][0]  ( .D(n21474), .CK(clk), .Q(\mem[579][0] ) );
  DFF_X1 \mem_reg[578][7]  ( .D(n21475), .CK(clk), .Q(\mem[578][7] ) );
  DFF_X1 \mem_reg[578][6]  ( .D(n21476), .CK(clk), .Q(\mem[578][6] ) );
  DFF_X1 \mem_reg[578][5]  ( .D(n21477), .CK(clk), .Q(\mem[578][5] ) );
  DFF_X1 \mem_reg[578][4]  ( .D(n21478), .CK(clk), .Q(\mem[578][4] ) );
  DFF_X1 \mem_reg[578][3]  ( .D(n21479), .CK(clk), .Q(\mem[578][3] ) );
  DFF_X1 \mem_reg[578][2]  ( .D(n21480), .CK(clk), .Q(\mem[578][2] ) );
  DFF_X1 \mem_reg[578][1]  ( .D(n21481), .CK(clk), .Q(\mem[578][1] ) );
  DFF_X1 \mem_reg[578][0]  ( .D(n21482), .CK(clk), .Q(\mem[578][0] ) );
  DFF_X1 \mem_reg[577][7]  ( .D(n21483), .CK(clk), .Q(\mem[577][7] ) );
  DFF_X1 \mem_reg[577][6]  ( .D(n21484), .CK(clk), .Q(\mem[577][6] ) );
  DFF_X1 \mem_reg[577][5]  ( .D(n21485), .CK(clk), .Q(\mem[577][5] ) );
  DFF_X1 \mem_reg[577][4]  ( .D(n21486), .CK(clk), .Q(\mem[577][4] ) );
  DFF_X1 \mem_reg[577][3]  ( .D(n21487), .CK(clk), .Q(\mem[577][3] ) );
  DFF_X1 \mem_reg[577][2]  ( .D(n21488), .CK(clk), .Q(\mem[577][2] ) );
  DFF_X1 \mem_reg[577][1]  ( .D(n21489), .CK(clk), .Q(\mem[577][1] ) );
  DFF_X1 \mem_reg[577][0]  ( .D(n21490), .CK(clk), .Q(\mem[577][0] ) );
  DFF_X1 \mem_reg[576][7]  ( .D(n21491), .CK(clk), .Q(\mem[576][7] ) );
  DFF_X1 \mem_reg[576][6]  ( .D(n21492), .CK(clk), .Q(\mem[576][6] ) );
  DFF_X1 \mem_reg[576][5]  ( .D(n21493), .CK(clk), .Q(\mem[576][5] ) );
  DFF_X1 \mem_reg[576][4]  ( .D(n21494), .CK(clk), .Q(\mem[576][4] ) );
  DFF_X1 \mem_reg[576][3]  ( .D(n21495), .CK(clk), .Q(\mem[576][3] ) );
  DFF_X1 \mem_reg[576][2]  ( .D(n21496), .CK(clk), .Q(\mem[576][2] ) );
  DFF_X1 \mem_reg[576][1]  ( .D(n21497), .CK(clk), .Q(\mem[576][1] ) );
  DFF_X1 \mem_reg[576][0]  ( .D(n21498), .CK(clk), .Q(\mem[576][0] ) );
  DFF_X1 \mem_reg[575][7]  ( .D(n21499), .CK(clk), .Q(\mem[575][7] ) );
  DFF_X1 \mem_reg[575][6]  ( .D(n21500), .CK(clk), .Q(\mem[575][6] ) );
  DFF_X1 \mem_reg[575][5]  ( .D(n21501), .CK(clk), .Q(\mem[575][5] ) );
  DFF_X1 \mem_reg[575][4]  ( .D(n21502), .CK(clk), .Q(\mem[575][4] ) );
  DFF_X1 \mem_reg[575][3]  ( .D(n21503), .CK(clk), .Q(\mem[575][3] ) );
  DFF_X1 \mem_reg[575][2]  ( .D(n21504), .CK(clk), .Q(\mem[575][2] ) );
  DFF_X1 \mem_reg[575][1]  ( .D(n21505), .CK(clk), .Q(\mem[575][1] ) );
  DFF_X1 \mem_reg[575][0]  ( .D(n21506), .CK(clk), .Q(\mem[575][0] ) );
  DFF_X1 \mem_reg[574][7]  ( .D(n21507), .CK(clk), .Q(\mem[574][7] ) );
  DFF_X1 \mem_reg[574][6]  ( .D(n21508), .CK(clk), .Q(\mem[574][6] ) );
  DFF_X1 \mem_reg[574][5]  ( .D(n21509), .CK(clk), .Q(\mem[574][5] ) );
  DFF_X1 \mem_reg[574][4]  ( .D(n21510), .CK(clk), .Q(\mem[574][4] ) );
  DFF_X1 \mem_reg[574][3]  ( .D(n21511), .CK(clk), .Q(\mem[574][3] ) );
  DFF_X1 \mem_reg[574][2]  ( .D(n21512), .CK(clk), .Q(\mem[574][2] ) );
  DFF_X1 \mem_reg[574][1]  ( .D(n21513), .CK(clk), .Q(\mem[574][1] ) );
  DFF_X1 \mem_reg[574][0]  ( .D(n21514), .CK(clk), .Q(\mem[574][0] ) );
  DFF_X1 \mem_reg[573][7]  ( .D(n21515), .CK(clk), .Q(\mem[573][7] ) );
  DFF_X1 \mem_reg[573][6]  ( .D(n21516), .CK(clk), .Q(\mem[573][6] ) );
  DFF_X1 \mem_reg[573][5]  ( .D(n21517), .CK(clk), .Q(\mem[573][5] ) );
  DFF_X1 \mem_reg[573][4]  ( .D(n21518), .CK(clk), .Q(\mem[573][4] ) );
  DFF_X1 \mem_reg[573][3]  ( .D(n21519), .CK(clk), .Q(\mem[573][3] ) );
  DFF_X1 \mem_reg[573][2]  ( .D(n21520), .CK(clk), .Q(\mem[573][2] ) );
  DFF_X1 \mem_reg[573][1]  ( .D(n21521), .CK(clk), .Q(\mem[573][1] ) );
  DFF_X1 \mem_reg[573][0]  ( .D(n21522), .CK(clk), .Q(\mem[573][0] ) );
  DFF_X1 \mem_reg[572][7]  ( .D(n21523), .CK(clk), .Q(\mem[572][7] ) );
  DFF_X1 \mem_reg[572][6]  ( .D(n21524), .CK(clk), .Q(\mem[572][6] ) );
  DFF_X1 \mem_reg[572][5]  ( .D(n21525), .CK(clk), .Q(\mem[572][5] ) );
  DFF_X1 \mem_reg[572][4]  ( .D(n21526), .CK(clk), .Q(\mem[572][4] ) );
  DFF_X1 \mem_reg[572][3]  ( .D(n21527), .CK(clk), .Q(\mem[572][3] ) );
  DFF_X1 \mem_reg[572][2]  ( .D(n21528), .CK(clk), .Q(\mem[572][2] ) );
  DFF_X1 \mem_reg[572][1]  ( .D(n21529), .CK(clk), .Q(\mem[572][1] ) );
  DFF_X1 \mem_reg[572][0]  ( .D(n21530), .CK(clk), .Q(\mem[572][0] ) );
  DFF_X1 \mem_reg[571][7]  ( .D(n21531), .CK(clk), .Q(\mem[571][7] ) );
  DFF_X1 \mem_reg[571][6]  ( .D(n21532), .CK(clk), .Q(\mem[571][6] ) );
  DFF_X1 \mem_reg[571][5]  ( .D(n21533), .CK(clk), .Q(\mem[571][5] ) );
  DFF_X1 \mem_reg[571][4]  ( .D(n21534), .CK(clk), .Q(\mem[571][4] ) );
  DFF_X1 \mem_reg[571][3]  ( .D(n21535), .CK(clk), .Q(\mem[571][3] ) );
  DFF_X1 \mem_reg[571][2]  ( .D(n21536), .CK(clk), .Q(\mem[571][2] ) );
  DFF_X1 \mem_reg[571][1]  ( .D(n21537), .CK(clk), .Q(\mem[571][1] ) );
  DFF_X1 \mem_reg[571][0]  ( .D(n21538), .CK(clk), .Q(\mem[571][0] ) );
  DFF_X1 \mem_reg[570][7]  ( .D(n21539), .CK(clk), .Q(\mem[570][7] ) );
  DFF_X1 \mem_reg[570][6]  ( .D(n21540), .CK(clk), .Q(\mem[570][6] ) );
  DFF_X1 \mem_reg[570][5]  ( .D(n21541), .CK(clk), .Q(\mem[570][5] ) );
  DFF_X1 \mem_reg[570][4]  ( .D(n21542), .CK(clk), .Q(\mem[570][4] ) );
  DFF_X1 \mem_reg[570][3]  ( .D(n21543), .CK(clk), .Q(\mem[570][3] ) );
  DFF_X1 \mem_reg[570][2]  ( .D(n21544), .CK(clk), .Q(\mem[570][2] ) );
  DFF_X1 \mem_reg[570][1]  ( .D(n21545), .CK(clk), .Q(\mem[570][1] ) );
  DFF_X1 \mem_reg[570][0]  ( .D(n21546), .CK(clk), .Q(\mem[570][0] ) );
  DFF_X1 \mem_reg[569][7]  ( .D(n21547), .CK(clk), .Q(\mem[569][7] ) );
  DFF_X1 \mem_reg[569][6]  ( .D(n21548), .CK(clk), .Q(\mem[569][6] ) );
  DFF_X1 \mem_reg[569][5]  ( .D(n21549), .CK(clk), .Q(\mem[569][5] ) );
  DFF_X1 \mem_reg[569][4]  ( .D(n21550), .CK(clk), .Q(\mem[569][4] ) );
  DFF_X1 \mem_reg[569][3]  ( .D(n21551), .CK(clk), .Q(\mem[569][3] ) );
  DFF_X1 \mem_reg[569][2]  ( .D(n21552), .CK(clk), .Q(\mem[569][2] ) );
  DFF_X1 \mem_reg[569][1]  ( .D(n21553), .CK(clk), .Q(\mem[569][1] ) );
  DFF_X1 \mem_reg[569][0]  ( .D(n21554), .CK(clk), .Q(\mem[569][0] ) );
  DFF_X1 \mem_reg[568][7]  ( .D(n21555), .CK(clk), .Q(\mem[568][7] ) );
  DFF_X1 \mem_reg[568][6]  ( .D(n21556), .CK(clk), .Q(\mem[568][6] ) );
  DFF_X1 \mem_reg[568][5]  ( .D(n21557), .CK(clk), .Q(\mem[568][5] ) );
  DFF_X1 \mem_reg[568][4]  ( .D(n21558), .CK(clk), .Q(\mem[568][4] ) );
  DFF_X1 \mem_reg[568][3]  ( .D(n21559), .CK(clk), .Q(\mem[568][3] ) );
  DFF_X1 \mem_reg[568][2]  ( .D(n21560), .CK(clk), .Q(\mem[568][2] ) );
  DFF_X1 \mem_reg[568][1]  ( .D(n21561), .CK(clk), .Q(\mem[568][1] ) );
  DFF_X1 \mem_reg[568][0]  ( .D(n21562), .CK(clk), .Q(\mem[568][0] ) );
  DFF_X1 \mem_reg[567][7]  ( .D(n21563), .CK(clk), .Q(\mem[567][7] ) );
  DFF_X1 \mem_reg[567][6]  ( .D(n21564), .CK(clk), .Q(\mem[567][6] ) );
  DFF_X1 \mem_reg[567][5]  ( .D(n21565), .CK(clk), .Q(\mem[567][5] ) );
  DFF_X1 \mem_reg[567][4]  ( .D(n21566), .CK(clk), .Q(\mem[567][4] ) );
  DFF_X1 \mem_reg[567][3]  ( .D(n21567), .CK(clk), .Q(\mem[567][3] ) );
  DFF_X1 \mem_reg[567][2]  ( .D(n21568), .CK(clk), .Q(\mem[567][2] ) );
  DFF_X1 \mem_reg[567][1]  ( .D(n21569), .CK(clk), .Q(\mem[567][1] ) );
  DFF_X1 \mem_reg[567][0]  ( .D(n21570), .CK(clk), .Q(\mem[567][0] ) );
  DFF_X1 \mem_reg[566][7]  ( .D(n21571), .CK(clk), .Q(\mem[566][7] ) );
  DFF_X1 \mem_reg[566][6]  ( .D(n21572), .CK(clk), .Q(\mem[566][6] ) );
  DFF_X1 \mem_reg[566][5]  ( .D(n21573), .CK(clk), .Q(\mem[566][5] ) );
  DFF_X1 \mem_reg[566][4]  ( .D(n21574), .CK(clk), .Q(\mem[566][4] ) );
  DFF_X1 \mem_reg[566][3]  ( .D(n21575), .CK(clk), .Q(\mem[566][3] ) );
  DFF_X1 \mem_reg[566][2]  ( .D(n21576), .CK(clk), .Q(\mem[566][2] ) );
  DFF_X1 \mem_reg[566][1]  ( .D(n21577), .CK(clk), .Q(\mem[566][1] ) );
  DFF_X1 \mem_reg[566][0]  ( .D(n21578), .CK(clk), .Q(\mem[566][0] ) );
  DFF_X1 \mem_reg[565][7]  ( .D(n21579), .CK(clk), .Q(\mem[565][7] ) );
  DFF_X1 \mem_reg[565][6]  ( .D(n21580), .CK(clk), .Q(\mem[565][6] ) );
  DFF_X1 \mem_reg[565][5]  ( .D(n21581), .CK(clk), .Q(\mem[565][5] ) );
  DFF_X1 \mem_reg[565][4]  ( .D(n21582), .CK(clk), .Q(\mem[565][4] ) );
  DFF_X1 \mem_reg[565][3]  ( .D(n21583), .CK(clk), .Q(\mem[565][3] ) );
  DFF_X1 \mem_reg[565][2]  ( .D(n21584), .CK(clk), .Q(\mem[565][2] ) );
  DFF_X1 \mem_reg[565][1]  ( .D(n21585), .CK(clk), .Q(\mem[565][1] ) );
  DFF_X1 \mem_reg[565][0]  ( .D(n21586), .CK(clk), .Q(\mem[565][0] ) );
  DFF_X1 \mem_reg[564][7]  ( .D(n21587), .CK(clk), .Q(\mem[564][7] ) );
  DFF_X1 \mem_reg[564][6]  ( .D(n21588), .CK(clk), .Q(\mem[564][6] ) );
  DFF_X1 \mem_reg[564][5]  ( .D(n21589), .CK(clk), .Q(\mem[564][5] ) );
  DFF_X1 \mem_reg[564][4]  ( .D(n21590), .CK(clk), .Q(\mem[564][4] ) );
  DFF_X1 \mem_reg[564][3]  ( .D(n21591), .CK(clk), .Q(\mem[564][3] ) );
  DFF_X1 \mem_reg[564][2]  ( .D(n21592), .CK(clk), .Q(\mem[564][2] ) );
  DFF_X1 \mem_reg[564][1]  ( .D(n21593), .CK(clk), .Q(\mem[564][1] ) );
  DFF_X1 \mem_reg[564][0]  ( .D(n21594), .CK(clk), .Q(\mem[564][0] ) );
  DFF_X1 \mem_reg[563][7]  ( .D(n21595), .CK(clk), .Q(\mem[563][7] ) );
  DFF_X1 \mem_reg[563][6]  ( .D(n21596), .CK(clk), .Q(\mem[563][6] ) );
  DFF_X1 \mem_reg[563][5]  ( .D(n21597), .CK(clk), .Q(\mem[563][5] ) );
  DFF_X1 \mem_reg[563][4]  ( .D(n21598), .CK(clk), .Q(\mem[563][4] ) );
  DFF_X1 \mem_reg[563][3]  ( .D(n21599), .CK(clk), .Q(\mem[563][3] ) );
  DFF_X1 \mem_reg[563][2]  ( .D(n21600), .CK(clk), .Q(\mem[563][2] ) );
  DFF_X1 \mem_reg[563][1]  ( .D(n21601), .CK(clk), .Q(\mem[563][1] ) );
  DFF_X1 \mem_reg[563][0]  ( .D(n21602), .CK(clk), .Q(\mem[563][0] ) );
  DFF_X1 \mem_reg[562][7]  ( .D(n21603), .CK(clk), .Q(\mem[562][7] ) );
  DFF_X1 \mem_reg[562][6]  ( .D(n21604), .CK(clk), .Q(\mem[562][6] ) );
  DFF_X1 \mem_reg[562][5]  ( .D(n21605), .CK(clk), .Q(\mem[562][5] ) );
  DFF_X1 \mem_reg[562][4]  ( .D(n21606), .CK(clk), .Q(\mem[562][4] ) );
  DFF_X1 \mem_reg[562][3]  ( .D(n21607), .CK(clk), .Q(\mem[562][3] ) );
  DFF_X1 \mem_reg[562][2]  ( .D(n21608), .CK(clk), .Q(\mem[562][2] ) );
  DFF_X1 \mem_reg[562][1]  ( .D(n21609), .CK(clk), .Q(\mem[562][1] ) );
  DFF_X1 \mem_reg[562][0]  ( .D(n21610), .CK(clk), .Q(\mem[562][0] ) );
  DFF_X1 \mem_reg[561][7]  ( .D(n21611), .CK(clk), .Q(\mem[561][7] ) );
  DFF_X1 \mem_reg[561][6]  ( .D(n21612), .CK(clk), .Q(\mem[561][6] ) );
  DFF_X1 \mem_reg[561][5]  ( .D(n21613), .CK(clk), .Q(\mem[561][5] ) );
  DFF_X1 \mem_reg[561][4]  ( .D(n21614), .CK(clk), .Q(\mem[561][4] ) );
  DFF_X1 \mem_reg[561][3]  ( .D(n21615), .CK(clk), .Q(\mem[561][3] ) );
  DFF_X1 \mem_reg[561][2]  ( .D(n21616), .CK(clk), .Q(\mem[561][2] ) );
  DFF_X1 \mem_reg[561][1]  ( .D(n21617), .CK(clk), .Q(\mem[561][1] ) );
  DFF_X1 \mem_reg[561][0]  ( .D(n21618), .CK(clk), .Q(\mem[561][0] ) );
  DFF_X1 \mem_reg[560][7]  ( .D(n21619), .CK(clk), .Q(\mem[560][7] ) );
  DFF_X1 \mem_reg[560][6]  ( .D(n21620), .CK(clk), .Q(\mem[560][6] ) );
  DFF_X1 \mem_reg[560][5]  ( .D(n21621), .CK(clk), .Q(\mem[560][5] ) );
  DFF_X1 \mem_reg[560][4]  ( .D(n21622), .CK(clk), .Q(\mem[560][4] ) );
  DFF_X1 \mem_reg[560][3]  ( .D(n21623), .CK(clk), .Q(\mem[560][3] ) );
  DFF_X1 \mem_reg[560][2]  ( .D(n21624), .CK(clk), .Q(\mem[560][2] ) );
  DFF_X1 \mem_reg[560][1]  ( .D(n21625), .CK(clk), .Q(\mem[560][1] ) );
  DFF_X1 \mem_reg[560][0]  ( .D(n21626), .CK(clk), .Q(\mem[560][0] ) );
  DFF_X1 \mem_reg[559][7]  ( .D(n21627), .CK(clk), .Q(\mem[559][7] ) );
  DFF_X1 \mem_reg[559][6]  ( .D(n21628), .CK(clk), .Q(\mem[559][6] ) );
  DFF_X1 \mem_reg[559][5]  ( .D(n21629), .CK(clk), .Q(\mem[559][5] ) );
  DFF_X1 \mem_reg[559][4]  ( .D(n21630), .CK(clk), .Q(\mem[559][4] ) );
  DFF_X1 \mem_reg[559][3]  ( .D(n21631), .CK(clk), .Q(\mem[559][3] ) );
  DFF_X1 \mem_reg[559][2]  ( .D(n21632), .CK(clk), .Q(\mem[559][2] ) );
  DFF_X1 \mem_reg[559][1]  ( .D(n21633), .CK(clk), .Q(\mem[559][1] ) );
  DFF_X1 \mem_reg[559][0]  ( .D(n21634), .CK(clk), .Q(\mem[559][0] ) );
  DFF_X1 \mem_reg[558][7]  ( .D(n21635), .CK(clk), .Q(\mem[558][7] ) );
  DFF_X1 \mem_reg[558][6]  ( .D(n21636), .CK(clk), .Q(\mem[558][6] ) );
  DFF_X1 \mem_reg[558][5]  ( .D(n21637), .CK(clk), .Q(\mem[558][5] ) );
  DFF_X1 \mem_reg[558][4]  ( .D(n21638), .CK(clk), .Q(\mem[558][4] ) );
  DFF_X1 \mem_reg[558][3]  ( .D(n21639), .CK(clk), .Q(\mem[558][3] ) );
  DFF_X1 \mem_reg[558][2]  ( .D(n21640), .CK(clk), .Q(\mem[558][2] ) );
  DFF_X1 \mem_reg[558][1]  ( .D(n21641), .CK(clk), .Q(\mem[558][1] ) );
  DFF_X1 \mem_reg[558][0]  ( .D(n21642), .CK(clk), .Q(\mem[558][0] ) );
  DFF_X1 \mem_reg[557][7]  ( .D(n21643), .CK(clk), .Q(\mem[557][7] ) );
  DFF_X1 \mem_reg[557][6]  ( .D(n21644), .CK(clk), .Q(\mem[557][6] ) );
  DFF_X1 \mem_reg[557][5]  ( .D(n21645), .CK(clk), .Q(\mem[557][5] ) );
  DFF_X1 \mem_reg[557][4]  ( .D(n21646), .CK(clk), .Q(\mem[557][4] ) );
  DFF_X1 \mem_reg[557][3]  ( .D(n21647), .CK(clk), .Q(\mem[557][3] ) );
  DFF_X1 \mem_reg[557][2]  ( .D(n21648), .CK(clk), .Q(\mem[557][2] ) );
  DFF_X1 \mem_reg[557][1]  ( .D(n21649), .CK(clk), .Q(\mem[557][1] ) );
  DFF_X1 \mem_reg[557][0]  ( .D(n21650), .CK(clk), .Q(\mem[557][0] ) );
  DFF_X1 \mem_reg[556][7]  ( .D(n21651), .CK(clk), .Q(\mem[556][7] ) );
  DFF_X1 \mem_reg[556][6]  ( .D(n21652), .CK(clk), .Q(\mem[556][6] ) );
  DFF_X1 \mem_reg[556][5]  ( .D(n21653), .CK(clk), .Q(\mem[556][5] ) );
  DFF_X1 \mem_reg[556][4]  ( .D(n21654), .CK(clk), .Q(\mem[556][4] ) );
  DFF_X1 \mem_reg[556][3]  ( .D(n21655), .CK(clk), .Q(\mem[556][3] ) );
  DFF_X1 \mem_reg[556][2]  ( .D(n21656), .CK(clk), .Q(\mem[556][2] ) );
  DFF_X1 \mem_reg[556][1]  ( .D(n21657), .CK(clk), .Q(\mem[556][1] ) );
  DFF_X1 \mem_reg[556][0]  ( .D(n21658), .CK(clk), .Q(\mem[556][0] ) );
  DFF_X1 \mem_reg[555][7]  ( .D(n21659), .CK(clk), .Q(\mem[555][7] ) );
  DFF_X1 \mem_reg[555][6]  ( .D(n21660), .CK(clk), .Q(\mem[555][6] ) );
  DFF_X1 \mem_reg[555][5]  ( .D(n21661), .CK(clk), .Q(\mem[555][5] ) );
  DFF_X1 \mem_reg[555][4]  ( .D(n21662), .CK(clk), .Q(\mem[555][4] ) );
  DFF_X1 \mem_reg[555][3]  ( .D(n21663), .CK(clk), .Q(\mem[555][3] ) );
  DFF_X1 \mem_reg[555][2]  ( .D(n21664), .CK(clk), .Q(\mem[555][2] ) );
  DFF_X1 \mem_reg[555][1]  ( .D(n21665), .CK(clk), .Q(\mem[555][1] ) );
  DFF_X1 \mem_reg[555][0]  ( .D(n21666), .CK(clk), .Q(\mem[555][0] ) );
  DFF_X1 \mem_reg[554][7]  ( .D(n21667), .CK(clk), .Q(\mem[554][7] ) );
  DFF_X1 \mem_reg[554][6]  ( .D(n21668), .CK(clk), .Q(\mem[554][6] ) );
  DFF_X1 \mem_reg[554][5]  ( .D(n21669), .CK(clk), .Q(\mem[554][5] ) );
  DFF_X1 \mem_reg[554][4]  ( .D(n21670), .CK(clk), .Q(\mem[554][4] ) );
  DFF_X1 \mem_reg[554][3]  ( .D(n21671), .CK(clk), .Q(\mem[554][3] ) );
  DFF_X1 \mem_reg[554][2]  ( .D(n21672), .CK(clk), .Q(\mem[554][2] ) );
  DFF_X1 \mem_reg[554][1]  ( .D(n21673), .CK(clk), .Q(\mem[554][1] ) );
  DFF_X1 \mem_reg[554][0]  ( .D(n21674), .CK(clk), .Q(\mem[554][0] ) );
  DFF_X1 \mem_reg[553][7]  ( .D(n21675), .CK(clk), .Q(\mem[553][7] ) );
  DFF_X1 \mem_reg[553][6]  ( .D(n21676), .CK(clk), .Q(\mem[553][6] ) );
  DFF_X1 \mem_reg[553][5]  ( .D(n21677), .CK(clk), .Q(\mem[553][5] ) );
  DFF_X1 \mem_reg[553][4]  ( .D(n21678), .CK(clk), .Q(\mem[553][4] ) );
  DFF_X1 \mem_reg[553][3]  ( .D(n21679), .CK(clk), .Q(\mem[553][3] ) );
  DFF_X1 \mem_reg[553][2]  ( .D(n21680), .CK(clk), .Q(\mem[553][2] ) );
  DFF_X1 \mem_reg[553][1]  ( .D(n21681), .CK(clk), .Q(\mem[553][1] ) );
  DFF_X1 \mem_reg[553][0]  ( .D(n21682), .CK(clk), .Q(\mem[553][0] ) );
  DFF_X1 \mem_reg[552][7]  ( .D(n21683), .CK(clk), .Q(\mem[552][7] ) );
  DFF_X1 \mem_reg[552][6]  ( .D(n21684), .CK(clk), .Q(\mem[552][6] ) );
  DFF_X1 \mem_reg[552][5]  ( .D(n21685), .CK(clk), .Q(\mem[552][5] ) );
  DFF_X1 \mem_reg[552][4]  ( .D(n21686), .CK(clk), .Q(\mem[552][4] ) );
  DFF_X1 \mem_reg[552][3]  ( .D(n21687), .CK(clk), .Q(\mem[552][3] ) );
  DFF_X1 \mem_reg[552][2]  ( .D(n21688), .CK(clk), .Q(\mem[552][2] ) );
  DFF_X1 \mem_reg[552][1]  ( .D(n21689), .CK(clk), .Q(\mem[552][1] ) );
  DFF_X1 \mem_reg[552][0]  ( .D(n21690), .CK(clk), .Q(\mem[552][0] ) );
  DFF_X1 \mem_reg[551][7]  ( .D(n21691), .CK(clk), .Q(\mem[551][7] ) );
  DFF_X1 \mem_reg[551][6]  ( .D(n21692), .CK(clk), .Q(\mem[551][6] ) );
  DFF_X1 \mem_reg[551][5]  ( .D(n21693), .CK(clk), .Q(\mem[551][5] ) );
  DFF_X1 \mem_reg[551][4]  ( .D(n21694), .CK(clk), .Q(\mem[551][4] ) );
  DFF_X1 \mem_reg[551][3]  ( .D(n21695), .CK(clk), .Q(\mem[551][3] ) );
  DFF_X1 \mem_reg[551][2]  ( .D(n21696), .CK(clk), .Q(\mem[551][2] ) );
  DFF_X1 \mem_reg[551][1]  ( .D(n21697), .CK(clk), .Q(\mem[551][1] ) );
  DFF_X1 \mem_reg[551][0]  ( .D(n21698), .CK(clk), .Q(\mem[551][0] ) );
  DFF_X1 \mem_reg[550][7]  ( .D(n21699), .CK(clk), .Q(\mem[550][7] ) );
  DFF_X1 \mem_reg[550][6]  ( .D(n21700), .CK(clk), .Q(\mem[550][6] ) );
  DFF_X1 \mem_reg[550][5]  ( .D(n21701), .CK(clk), .Q(\mem[550][5] ) );
  DFF_X1 \mem_reg[550][4]  ( .D(n21702), .CK(clk), .Q(\mem[550][4] ) );
  DFF_X1 \mem_reg[550][3]  ( .D(n21703), .CK(clk), .Q(\mem[550][3] ) );
  DFF_X1 \mem_reg[550][2]  ( .D(n21704), .CK(clk), .Q(\mem[550][2] ) );
  DFF_X1 \mem_reg[550][1]  ( .D(n21705), .CK(clk), .Q(\mem[550][1] ) );
  DFF_X1 \mem_reg[550][0]  ( .D(n21706), .CK(clk), .Q(\mem[550][0] ) );
  DFF_X1 \mem_reg[549][7]  ( .D(n21707), .CK(clk), .Q(\mem[549][7] ) );
  DFF_X1 \mem_reg[549][6]  ( .D(n21708), .CK(clk), .Q(\mem[549][6] ) );
  DFF_X1 \mem_reg[549][5]  ( .D(n21709), .CK(clk), .Q(\mem[549][5] ) );
  DFF_X1 \mem_reg[549][4]  ( .D(n21710), .CK(clk), .Q(\mem[549][4] ) );
  DFF_X1 \mem_reg[549][3]  ( .D(n21711), .CK(clk), .Q(\mem[549][3] ) );
  DFF_X1 \mem_reg[549][2]  ( .D(n21712), .CK(clk), .Q(\mem[549][2] ) );
  DFF_X1 \mem_reg[549][1]  ( .D(n21713), .CK(clk), .Q(\mem[549][1] ) );
  DFF_X1 \mem_reg[549][0]  ( .D(n21714), .CK(clk), .Q(\mem[549][0] ) );
  DFF_X1 \mem_reg[548][7]  ( .D(n21715), .CK(clk), .Q(\mem[548][7] ) );
  DFF_X1 \mem_reg[548][6]  ( .D(n21716), .CK(clk), .Q(\mem[548][6] ) );
  DFF_X1 \mem_reg[548][5]  ( .D(n21717), .CK(clk), .Q(\mem[548][5] ) );
  DFF_X1 \mem_reg[548][4]  ( .D(n21718), .CK(clk), .Q(\mem[548][4] ) );
  DFF_X1 \mem_reg[548][3]  ( .D(n21719), .CK(clk), .Q(\mem[548][3] ) );
  DFF_X1 \mem_reg[548][2]  ( .D(n21720), .CK(clk), .Q(\mem[548][2] ) );
  DFF_X1 \mem_reg[548][1]  ( .D(n21721), .CK(clk), .Q(\mem[548][1] ) );
  DFF_X1 \mem_reg[548][0]  ( .D(n21722), .CK(clk), .Q(\mem[548][0] ) );
  DFF_X1 \mem_reg[547][7]  ( .D(n21723), .CK(clk), .Q(\mem[547][7] ) );
  DFF_X1 \mem_reg[547][6]  ( .D(n21724), .CK(clk), .Q(\mem[547][6] ) );
  DFF_X1 \mem_reg[547][5]  ( .D(n21725), .CK(clk), .Q(\mem[547][5] ) );
  DFF_X1 \mem_reg[547][4]  ( .D(n21726), .CK(clk), .Q(\mem[547][4] ) );
  DFF_X1 \mem_reg[547][3]  ( .D(n21727), .CK(clk), .Q(\mem[547][3] ) );
  DFF_X1 \mem_reg[547][2]  ( .D(n21728), .CK(clk), .Q(\mem[547][2] ) );
  DFF_X1 \mem_reg[547][1]  ( .D(n21729), .CK(clk), .Q(\mem[547][1] ) );
  DFF_X1 \mem_reg[547][0]  ( .D(n21730), .CK(clk), .Q(\mem[547][0] ) );
  DFF_X1 \mem_reg[546][7]  ( .D(n21731), .CK(clk), .Q(\mem[546][7] ) );
  DFF_X1 \mem_reg[546][6]  ( .D(n21732), .CK(clk), .Q(\mem[546][6] ) );
  DFF_X1 \mem_reg[546][5]  ( .D(n21733), .CK(clk), .Q(\mem[546][5] ) );
  DFF_X1 \mem_reg[546][4]  ( .D(n21734), .CK(clk), .Q(\mem[546][4] ) );
  DFF_X1 \mem_reg[546][3]  ( .D(n21735), .CK(clk), .Q(\mem[546][3] ) );
  DFF_X1 \mem_reg[546][2]  ( .D(n21736), .CK(clk), .Q(\mem[546][2] ) );
  DFF_X1 \mem_reg[546][1]  ( .D(n21737), .CK(clk), .Q(\mem[546][1] ) );
  DFF_X1 \mem_reg[546][0]  ( .D(n21738), .CK(clk), .Q(\mem[546][0] ) );
  DFF_X1 \mem_reg[545][7]  ( .D(n21739), .CK(clk), .Q(\mem[545][7] ) );
  DFF_X1 \mem_reg[545][6]  ( .D(n21740), .CK(clk), .Q(\mem[545][6] ) );
  DFF_X1 \mem_reg[545][5]  ( .D(n21741), .CK(clk), .Q(\mem[545][5] ) );
  DFF_X1 \mem_reg[545][4]  ( .D(n21742), .CK(clk), .Q(\mem[545][4] ) );
  DFF_X1 \mem_reg[545][3]  ( .D(n21743), .CK(clk), .Q(\mem[545][3] ) );
  DFF_X1 \mem_reg[545][2]  ( .D(n21744), .CK(clk), .Q(\mem[545][2] ) );
  DFF_X1 \mem_reg[545][1]  ( .D(n21745), .CK(clk), .Q(\mem[545][1] ) );
  DFF_X1 \mem_reg[545][0]  ( .D(n21746), .CK(clk), .Q(\mem[545][0] ) );
  DFF_X1 \mem_reg[544][7]  ( .D(n21747), .CK(clk), .Q(\mem[544][7] ) );
  DFF_X1 \mem_reg[544][6]  ( .D(n21748), .CK(clk), .Q(\mem[544][6] ) );
  DFF_X1 \mem_reg[544][5]  ( .D(n21749), .CK(clk), .Q(\mem[544][5] ) );
  DFF_X1 \mem_reg[544][4]  ( .D(n21750), .CK(clk), .Q(\mem[544][4] ) );
  DFF_X1 \mem_reg[544][3]  ( .D(n21751), .CK(clk), .Q(\mem[544][3] ) );
  DFF_X1 \mem_reg[544][2]  ( .D(n21752), .CK(clk), .Q(\mem[544][2] ) );
  DFF_X1 \mem_reg[544][1]  ( .D(n21753), .CK(clk), .Q(\mem[544][1] ) );
  DFF_X1 \mem_reg[544][0]  ( .D(n21754), .CK(clk), .Q(\mem[544][0] ) );
  DFF_X1 \mem_reg[543][7]  ( .D(n21755), .CK(clk), .Q(\mem[543][7] ) );
  DFF_X1 \mem_reg[543][6]  ( .D(n21756), .CK(clk), .Q(\mem[543][6] ) );
  DFF_X1 \mem_reg[543][5]  ( .D(n21757), .CK(clk), .Q(\mem[543][5] ) );
  DFF_X1 \mem_reg[543][4]  ( .D(n21758), .CK(clk), .Q(\mem[543][4] ) );
  DFF_X1 \mem_reg[543][3]  ( .D(n21759), .CK(clk), .Q(\mem[543][3] ) );
  DFF_X1 \mem_reg[543][2]  ( .D(n21760), .CK(clk), .Q(\mem[543][2] ) );
  DFF_X1 \mem_reg[543][1]  ( .D(n21761), .CK(clk), .Q(\mem[543][1] ) );
  DFF_X1 \mem_reg[543][0]  ( .D(n21762), .CK(clk), .Q(\mem[543][0] ) );
  DFF_X1 \mem_reg[542][7]  ( .D(n21763), .CK(clk), .Q(\mem[542][7] ) );
  DFF_X1 \mem_reg[542][6]  ( .D(n21764), .CK(clk), .Q(\mem[542][6] ) );
  DFF_X1 \mem_reg[542][5]  ( .D(n21765), .CK(clk), .Q(\mem[542][5] ) );
  DFF_X1 \mem_reg[542][4]  ( .D(n21766), .CK(clk), .Q(\mem[542][4] ) );
  DFF_X1 \mem_reg[542][3]  ( .D(n21767), .CK(clk), .Q(\mem[542][3] ) );
  DFF_X1 \mem_reg[542][2]  ( .D(n21768), .CK(clk), .Q(\mem[542][2] ) );
  DFF_X1 \mem_reg[542][1]  ( .D(n21769), .CK(clk), .Q(\mem[542][1] ) );
  DFF_X1 \mem_reg[542][0]  ( .D(n21770), .CK(clk), .Q(\mem[542][0] ) );
  DFF_X1 \mem_reg[541][7]  ( .D(n21771), .CK(clk), .Q(\mem[541][7] ) );
  DFF_X1 \mem_reg[541][6]  ( .D(n21772), .CK(clk), .Q(\mem[541][6] ) );
  DFF_X1 \mem_reg[541][5]  ( .D(n21773), .CK(clk), .Q(\mem[541][5] ) );
  DFF_X1 \mem_reg[541][4]  ( .D(n21774), .CK(clk), .Q(\mem[541][4] ) );
  DFF_X1 \mem_reg[541][3]  ( .D(n21775), .CK(clk), .Q(\mem[541][3] ) );
  DFF_X1 \mem_reg[541][2]  ( .D(n21776), .CK(clk), .Q(\mem[541][2] ) );
  DFF_X1 \mem_reg[541][1]  ( .D(n21777), .CK(clk), .Q(\mem[541][1] ) );
  DFF_X1 \mem_reg[541][0]  ( .D(n21778), .CK(clk), .Q(\mem[541][0] ) );
  DFF_X1 \mem_reg[540][7]  ( .D(n21779), .CK(clk), .Q(\mem[540][7] ) );
  DFF_X1 \mem_reg[540][6]  ( .D(n21780), .CK(clk), .Q(\mem[540][6] ) );
  DFF_X1 \mem_reg[540][5]  ( .D(n21781), .CK(clk), .Q(\mem[540][5] ) );
  DFF_X1 \mem_reg[540][4]  ( .D(n21782), .CK(clk), .Q(\mem[540][4] ) );
  DFF_X1 \mem_reg[540][3]  ( .D(n21783), .CK(clk), .Q(\mem[540][3] ) );
  DFF_X1 \mem_reg[540][2]  ( .D(n21784), .CK(clk), .Q(\mem[540][2] ) );
  DFF_X1 \mem_reg[540][1]  ( .D(n21785), .CK(clk), .Q(\mem[540][1] ) );
  DFF_X1 \mem_reg[540][0]  ( .D(n21786), .CK(clk), .Q(\mem[540][0] ) );
  DFF_X1 \mem_reg[539][7]  ( .D(n21787), .CK(clk), .Q(\mem[539][7] ) );
  DFF_X1 \mem_reg[539][6]  ( .D(n21788), .CK(clk), .Q(\mem[539][6] ) );
  DFF_X1 \mem_reg[539][5]  ( .D(n21789), .CK(clk), .Q(\mem[539][5] ) );
  DFF_X1 \mem_reg[539][4]  ( .D(n21790), .CK(clk), .Q(\mem[539][4] ) );
  DFF_X1 \mem_reg[539][3]  ( .D(n21791), .CK(clk), .Q(\mem[539][3] ) );
  DFF_X1 \mem_reg[539][2]  ( .D(n21792), .CK(clk), .Q(\mem[539][2] ) );
  DFF_X1 \mem_reg[539][1]  ( .D(n21793), .CK(clk), .Q(\mem[539][1] ) );
  DFF_X1 \mem_reg[539][0]  ( .D(n21794), .CK(clk), .Q(\mem[539][0] ) );
  DFF_X1 \mem_reg[538][7]  ( .D(n21795), .CK(clk), .Q(\mem[538][7] ) );
  DFF_X1 \mem_reg[538][6]  ( .D(n21796), .CK(clk), .Q(\mem[538][6] ) );
  DFF_X1 \mem_reg[538][5]  ( .D(n21797), .CK(clk), .Q(\mem[538][5] ) );
  DFF_X1 \mem_reg[538][4]  ( .D(n21798), .CK(clk), .Q(\mem[538][4] ) );
  DFF_X1 \mem_reg[538][3]  ( .D(n21799), .CK(clk), .Q(\mem[538][3] ) );
  DFF_X1 \mem_reg[538][2]  ( .D(n21800), .CK(clk), .Q(\mem[538][2] ) );
  DFF_X1 \mem_reg[538][1]  ( .D(n21801), .CK(clk), .Q(\mem[538][1] ) );
  DFF_X1 \mem_reg[538][0]  ( .D(n21802), .CK(clk), .Q(\mem[538][0] ) );
  DFF_X1 \mem_reg[537][7]  ( .D(n21803), .CK(clk), .Q(\mem[537][7] ) );
  DFF_X1 \mem_reg[537][6]  ( .D(n21804), .CK(clk), .Q(\mem[537][6] ) );
  DFF_X1 \mem_reg[537][5]  ( .D(n21805), .CK(clk), .Q(\mem[537][5] ) );
  DFF_X1 \mem_reg[537][4]  ( .D(n21806), .CK(clk), .Q(\mem[537][4] ) );
  DFF_X1 \mem_reg[537][3]  ( .D(n21807), .CK(clk), .Q(\mem[537][3] ) );
  DFF_X1 \mem_reg[537][2]  ( .D(n21808), .CK(clk), .Q(\mem[537][2] ) );
  DFF_X1 \mem_reg[537][1]  ( .D(n21809), .CK(clk), .Q(\mem[537][1] ) );
  DFF_X1 \mem_reg[537][0]  ( .D(n21810), .CK(clk), .Q(\mem[537][0] ) );
  DFF_X1 \mem_reg[536][7]  ( .D(n21811), .CK(clk), .Q(\mem[536][7] ) );
  DFF_X1 \mem_reg[536][6]  ( .D(n21812), .CK(clk), .Q(\mem[536][6] ) );
  DFF_X1 \mem_reg[536][5]  ( .D(n21813), .CK(clk), .Q(\mem[536][5] ) );
  DFF_X1 \mem_reg[536][4]  ( .D(n21814), .CK(clk), .Q(\mem[536][4] ) );
  DFF_X1 \mem_reg[536][3]  ( .D(n21815), .CK(clk), .Q(\mem[536][3] ) );
  DFF_X1 \mem_reg[536][2]  ( .D(n21816), .CK(clk), .Q(\mem[536][2] ) );
  DFF_X1 \mem_reg[536][1]  ( .D(n21817), .CK(clk), .Q(\mem[536][1] ) );
  DFF_X1 \mem_reg[536][0]  ( .D(n21818), .CK(clk), .Q(\mem[536][0] ) );
  DFF_X1 \mem_reg[535][7]  ( .D(n21819), .CK(clk), .Q(\mem[535][7] ) );
  DFF_X1 \mem_reg[535][6]  ( .D(n21820), .CK(clk), .Q(\mem[535][6] ) );
  DFF_X1 \mem_reg[535][5]  ( .D(n21821), .CK(clk), .Q(\mem[535][5] ) );
  DFF_X1 \mem_reg[535][4]  ( .D(n21822), .CK(clk), .Q(\mem[535][4] ) );
  DFF_X1 \mem_reg[535][3]  ( .D(n21823), .CK(clk), .Q(\mem[535][3] ) );
  DFF_X1 \mem_reg[535][2]  ( .D(n21824), .CK(clk), .Q(\mem[535][2] ) );
  DFF_X1 \mem_reg[535][1]  ( .D(n21825), .CK(clk), .Q(\mem[535][1] ) );
  DFF_X1 \mem_reg[535][0]  ( .D(n21826), .CK(clk), .Q(\mem[535][0] ) );
  DFF_X1 \mem_reg[534][7]  ( .D(n21827), .CK(clk), .Q(\mem[534][7] ) );
  DFF_X1 \mem_reg[534][6]  ( .D(n21828), .CK(clk), .Q(\mem[534][6] ) );
  DFF_X1 \mem_reg[534][5]  ( .D(n21829), .CK(clk), .Q(\mem[534][5] ) );
  DFF_X1 \mem_reg[534][4]  ( .D(n21830), .CK(clk), .Q(\mem[534][4] ) );
  DFF_X1 \mem_reg[534][3]  ( .D(n21831), .CK(clk), .Q(\mem[534][3] ) );
  DFF_X1 \mem_reg[534][2]  ( .D(n21832), .CK(clk), .Q(\mem[534][2] ) );
  DFF_X1 \mem_reg[534][1]  ( .D(n21833), .CK(clk), .Q(\mem[534][1] ) );
  DFF_X1 \mem_reg[534][0]  ( .D(n21834), .CK(clk), .Q(\mem[534][0] ) );
  DFF_X1 \mem_reg[533][7]  ( .D(n21835), .CK(clk), .Q(\mem[533][7] ) );
  DFF_X1 \mem_reg[533][6]  ( .D(n21836), .CK(clk), .Q(\mem[533][6] ) );
  DFF_X1 \mem_reg[533][5]  ( .D(n21837), .CK(clk), .Q(\mem[533][5] ) );
  DFF_X1 \mem_reg[533][4]  ( .D(n21838), .CK(clk), .Q(\mem[533][4] ) );
  DFF_X1 \mem_reg[533][3]  ( .D(n21839), .CK(clk), .Q(\mem[533][3] ) );
  DFF_X1 \mem_reg[533][2]  ( .D(n21840), .CK(clk), .Q(\mem[533][2] ) );
  DFF_X1 \mem_reg[533][1]  ( .D(n21841), .CK(clk), .Q(\mem[533][1] ) );
  DFF_X1 \mem_reg[533][0]  ( .D(n21842), .CK(clk), .Q(\mem[533][0] ) );
  DFF_X1 \mem_reg[532][7]  ( .D(n21843), .CK(clk), .Q(\mem[532][7] ) );
  DFF_X1 \mem_reg[532][6]  ( .D(n21844), .CK(clk), .Q(\mem[532][6] ) );
  DFF_X1 \mem_reg[532][5]  ( .D(n21845), .CK(clk), .Q(\mem[532][5] ) );
  DFF_X1 \mem_reg[532][4]  ( .D(n21846), .CK(clk), .Q(\mem[532][4] ) );
  DFF_X1 \mem_reg[532][3]  ( .D(n21847), .CK(clk), .Q(\mem[532][3] ) );
  DFF_X1 \mem_reg[532][2]  ( .D(n21848), .CK(clk), .Q(\mem[532][2] ) );
  DFF_X1 \mem_reg[532][1]  ( .D(n21849), .CK(clk), .Q(\mem[532][1] ) );
  DFF_X1 \mem_reg[532][0]  ( .D(n21850), .CK(clk), .Q(\mem[532][0] ) );
  DFF_X1 \mem_reg[531][7]  ( .D(n21851), .CK(clk), .Q(\mem[531][7] ) );
  DFF_X1 \mem_reg[531][6]  ( .D(n21852), .CK(clk), .Q(\mem[531][6] ) );
  DFF_X1 \mem_reg[531][5]  ( .D(n21853), .CK(clk), .Q(\mem[531][5] ) );
  DFF_X1 \mem_reg[531][4]  ( .D(n21854), .CK(clk), .Q(\mem[531][4] ) );
  DFF_X1 \mem_reg[531][3]  ( .D(n21855), .CK(clk), .Q(\mem[531][3] ) );
  DFF_X1 \mem_reg[531][2]  ( .D(n21856), .CK(clk), .Q(\mem[531][2] ) );
  DFF_X1 \mem_reg[531][1]  ( .D(n21857), .CK(clk), .Q(\mem[531][1] ) );
  DFF_X1 \mem_reg[531][0]  ( .D(n21858), .CK(clk), .Q(\mem[531][0] ) );
  DFF_X1 \mem_reg[530][7]  ( .D(n21859), .CK(clk), .Q(\mem[530][7] ) );
  DFF_X1 \mem_reg[530][6]  ( .D(n21860), .CK(clk), .Q(\mem[530][6] ) );
  DFF_X1 \mem_reg[530][5]  ( .D(n21861), .CK(clk), .Q(\mem[530][5] ) );
  DFF_X1 \mem_reg[530][4]  ( .D(n21862), .CK(clk), .Q(\mem[530][4] ) );
  DFF_X1 \mem_reg[530][3]  ( .D(n21863), .CK(clk), .Q(\mem[530][3] ) );
  DFF_X1 \mem_reg[530][2]  ( .D(n21864), .CK(clk), .Q(\mem[530][2] ) );
  DFF_X1 \mem_reg[530][1]  ( .D(n21865), .CK(clk), .Q(\mem[530][1] ) );
  DFF_X1 \mem_reg[530][0]  ( .D(n21866), .CK(clk), .Q(\mem[530][0] ) );
  DFF_X1 \mem_reg[529][7]  ( .D(n21867), .CK(clk), .Q(\mem[529][7] ) );
  DFF_X1 \mem_reg[529][6]  ( .D(n21868), .CK(clk), .Q(\mem[529][6] ) );
  DFF_X1 \mem_reg[529][5]  ( .D(n21869), .CK(clk), .Q(\mem[529][5] ) );
  DFF_X1 \mem_reg[529][4]  ( .D(n21870), .CK(clk), .Q(\mem[529][4] ) );
  DFF_X1 \mem_reg[529][3]  ( .D(n21871), .CK(clk), .Q(\mem[529][3] ) );
  DFF_X1 \mem_reg[529][2]  ( .D(n21872), .CK(clk), .Q(\mem[529][2] ) );
  DFF_X1 \mem_reg[529][1]  ( .D(n21873), .CK(clk), .Q(\mem[529][1] ) );
  DFF_X1 \mem_reg[529][0]  ( .D(n21874), .CK(clk), .Q(\mem[529][0] ) );
  DFF_X1 \mem_reg[528][7]  ( .D(n21875), .CK(clk), .Q(\mem[528][7] ) );
  DFF_X1 \mem_reg[528][6]  ( .D(n21876), .CK(clk), .Q(\mem[528][6] ) );
  DFF_X1 \mem_reg[528][5]  ( .D(n21877), .CK(clk), .Q(\mem[528][5] ) );
  DFF_X1 \mem_reg[528][4]  ( .D(n21878), .CK(clk), .Q(\mem[528][4] ) );
  DFF_X1 \mem_reg[528][3]  ( .D(n21879), .CK(clk), .Q(\mem[528][3] ) );
  DFF_X1 \mem_reg[528][2]  ( .D(n21880), .CK(clk), .Q(\mem[528][2] ) );
  DFF_X1 \mem_reg[528][1]  ( .D(n21881), .CK(clk), .Q(\mem[528][1] ) );
  DFF_X1 \mem_reg[528][0]  ( .D(n21882), .CK(clk), .Q(\mem[528][0] ) );
  DFF_X1 \mem_reg[527][7]  ( .D(n21883), .CK(clk), .Q(\mem[527][7] ) );
  DFF_X1 \mem_reg[527][6]  ( .D(n21884), .CK(clk), .Q(\mem[527][6] ) );
  DFF_X1 \mem_reg[527][5]  ( .D(n21885), .CK(clk), .Q(\mem[527][5] ) );
  DFF_X1 \mem_reg[527][4]  ( .D(n21886), .CK(clk), .Q(\mem[527][4] ) );
  DFF_X1 \mem_reg[527][3]  ( .D(n21887), .CK(clk), .Q(\mem[527][3] ) );
  DFF_X1 \mem_reg[527][2]  ( .D(n21888), .CK(clk), .Q(\mem[527][2] ) );
  DFF_X1 \mem_reg[527][1]  ( .D(n21889), .CK(clk), .Q(\mem[527][1] ) );
  DFF_X1 \mem_reg[527][0]  ( .D(n21890), .CK(clk), .Q(\mem[527][0] ) );
  DFF_X1 \mem_reg[526][7]  ( .D(n21891), .CK(clk), .Q(\mem[526][7] ) );
  DFF_X1 \mem_reg[526][6]  ( .D(n21892), .CK(clk), .Q(\mem[526][6] ) );
  DFF_X1 \mem_reg[526][5]  ( .D(n21893), .CK(clk), .Q(\mem[526][5] ) );
  DFF_X1 \mem_reg[526][4]  ( .D(n21894), .CK(clk), .Q(\mem[526][4] ) );
  DFF_X1 \mem_reg[526][3]  ( .D(n21895), .CK(clk), .Q(\mem[526][3] ) );
  DFF_X1 \mem_reg[526][2]  ( .D(n21896), .CK(clk), .Q(\mem[526][2] ) );
  DFF_X1 \mem_reg[526][1]  ( .D(n21897), .CK(clk), .Q(\mem[526][1] ) );
  DFF_X1 \mem_reg[526][0]  ( .D(n21898), .CK(clk), .Q(\mem[526][0] ) );
  DFF_X1 \mem_reg[525][7]  ( .D(n21899), .CK(clk), .Q(\mem[525][7] ) );
  DFF_X1 \mem_reg[525][6]  ( .D(n21900), .CK(clk), .Q(\mem[525][6] ) );
  DFF_X1 \mem_reg[525][5]  ( .D(n21901), .CK(clk), .Q(\mem[525][5] ) );
  DFF_X1 \mem_reg[525][4]  ( .D(n21902), .CK(clk), .Q(\mem[525][4] ) );
  DFF_X1 \mem_reg[525][3]  ( .D(n21903), .CK(clk), .Q(\mem[525][3] ) );
  DFF_X1 \mem_reg[525][2]  ( .D(n21904), .CK(clk), .Q(\mem[525][2] ) );
  DFF_X1 \mem_reg[525][1]  ( .D(n21905), .CK(clk), .Q(\mem[525][1] ) );
  DFF_X1 \mem_reg[525][0]  ( .D(n21906), .CK(clk), .Q(\mem[525][0] ) );
  DFF_X1 \mem_reg[524][7]  ( .D(n21907), .CK(clk), .Q(\mem[524][7] ) );
  DFF_X1 \mem_reg[524][6]  ( .D(n21908), .CK(clk), .Q(\mem[524][6] ) );
  DFF_X1 \mem_reg[524][5]  ( .D(n21909), .CK(clk), .Q(\mem[524][5] ) );
  DFF_X1 \mem_reg[524][4]  ( .D(n21910), .CK(clk), .Q(\mem[524][4] ) );
  DFF_X1 \mem_reg[524][3]  ( .D(n21911), .CK(clk), .Q(\mem[524][3] ) );
  DFF_X1 \mem_reg[524][2]  ( .D(n21912), .CK(clk), .Q(\mem[524][2] ) );
  DFF_X1 \mem_reg[524][1]  ( .D(n21913), .CK(clk), .Q(\mem[524][1] ) );
  DFF_X1 \mem_reg[524][0]  ( .D(n21914), .CK(clk), .Q(\mem[524][0] ) );
  DFF_X1 \mem_reg[523][7]  ( .D(n21915), .CK(clk), .Q(\mem[523][7] ) );
  DFF_X1 \mem_reg[523][6]  ( .D(n21916), .CK(clk), .Q(\mem[523][6] ) );
  DFF_X1 \mem_reg[523][5]  ( .D(n21917), .CK(clk), .Q(\mem[523][5] ) );
  DFF_X1 \mem_reg[523][4]  ( .D(n21918), .CK(clk), .Q(\mem[523][4] ) );
  DFF_X1 \mem_reg[523][3]  ( .D(n21919), .CK(clk), .Q(\mem[523][3] ) );
  DFF_X1 \mem_reg[523][2]  ( .D(n21920), .CK(clk), .Q(\mem[523][2] ) );
  DFF_X1 \mem_reg[523][1]  ( .D(n21921), .CK(clk), .Q(\mem[523][1] ) );
  DFF_X1 \mem_reg[523][0]  ( .D(n21922), .CK(clk), .Q(\mem[523][0] ) );
  DFF_X1 \mem_reg[522][7]  ( .D(n21923), .CK(clk), .Q(\mem[522][7] ) );
  DFF_X1 \mem_reg[522][6]  ( .D(n21924), .CK(clk), .Q(\mem[522][6] ) );
  DFF_X1 \mem_reg[522][5]  ( .D(n21925), .CK(clk), .Q(\mem[522][5] ) );
  DFF_X1 \mem_reg[522][4]  ( .D(n21926), .CK(clk), .Q(\mem[522][4] ) );
  DFF_X1 \mem_reg[522][3]  ( .D(n21927), .CK(clk), .Q(\mem[522][3] ) );
  DFF_X1 \mem_reg[522][2]  ( .D(n21928), .CK(clk), .Q(\mem[522][2] ) );
  DFF_X1 \mem_reg[522][1]  ( .D(n21929), .CK(clk), .Q(\mem[522][1] ) );
  DFF_X1 \mem_reg[522][0]  ( .D(n21930), .CK(clk), .Q(\mem[522][0] ) );
  DFF_X1 \mem_reg[521][7]  ( .D(n21931), .CK(clk), .Q(\mem[521][7] ) );
  DFF_X1 \mem_reg[521][6]  ( .D(n21932), .CK(clk), .Q(\mem[521][6] ) );
  DFF_X1 \mem_reg[521][5]  ( .D(n21933), .CK(clk), .Q(\mem[521][5] ) );
  DFF_X1 \mem_reg[521][4]  ( .D(n21934), .CK(clk), .Q(\mem[521][4] ) );
  DFF_X1 \mem_reg[521][3]  ( .D(n21935), .CK(clk), .Q(\mem[521][3] ) );
  DFF_X1 \mem_reg[521][2]  ( .D(n21936), .CK(clk), .Q(\mem[521][2] ) );
  DFF_X1 \mem_reg[521][1]  ( .D(n21937), .CK(clk), .Q(\mem[521][1] ) );
  DFF_X1 \mem_reg[521][0]  ( .D(n21938), .CK(clk), .Q(\mem[521][0] ) );
  DFF_X1 \mem_reg[520][7]  ( .D(n21939), .CK(clk), .Q(\mem[520][7] ) );
  DFF_X1 \mem_reg[520][6]  ( .D(n21940), .CK(clk), .Q(\mem[520][6] ) );
  DFF_X1 \mem_reg[520][5]  ( .D(n21941), .CK(clk), .Q(\mem[520][5] ) );
  DFF_X1 \mem_reg[520][4]  ( .D(n21942), .CK(clk), .Q(\mem[520][4] ) );
  DFF_X1 \mem_reg[520][3]  ( .D(n21943), .CK(clk), .Q(\mem[520][3] ) );
  DFF_X1 \mem_reg[520][2]  ( .D(n21944), .CK(clk), .Q(\mem[520][2] ) );
  DFF_X1 \mem_reg[520][1]  ( .D(n21945), .CK(clk), .Q(\mem[520][1] ) );
  DFF_X1 \mem_reg[520][0]  ( .D(n21946), .CK(clk), .Q(\mem[520][0] ) );
  DFF_X1 \mem_reg[519][7]  ( .D(n21947), .CK(clk), .Q(\mem[519][7] ) );
  DFF_X1 \mem_reg[519][6]  ( .D(n21948), .CK(clk), .Q(\mem[519][6] ) );
  DFF_X1 \mem_reg[519][5]  ( .D(n21949), .CK(clk), .Q(\mem[519][5] ) );
  DFF_X1 \mem_reg[519][4]  ( .D(n21950), .CK(clk), .Q(\mem[519][4] ) );
  DFF_X1 \mem_reg[519][3]  ( .D(n21951), .CK(clk), .Q(\mem[519][3] ) );
  DFF_X1 \mem_reg[519][2]  ( .D(n21952), .CK(clk), .Q(\mem[519][2] ) );
  DFF_X1 \mem_reg[519][1]  ( .D(n21953), .CK(clk), .Q(\mem[519][1] ) );
  DFF_X1 \mem_reg[519][0]  ( .D(n21954), .CK(clk), .Q(\mem[519][0] ) );
  DFF_X1 \mem_reg[518][7]  ( .D(n21955), .CK(clk), .Q(\mem[518][7] ) );
  DFF_X1 \mem_reg[518][6]  ( .D(n21956), .CK(clk), .Q(\mem[518][6] ) );
  DFF_X1 \mem_reg[518][5]  ( .D(n21957), .CK(clk), .Q(\mem[518][5] ) );
  DFF_X1 \mem_reg[518][4]  ( .D(n21958), .CK(clk), .Q(\mem[518][4] ) );
  DFF_X1 \mem_reg[518][3]  ( .D(n21959), .CK(clk), .Q(\mem[518][3] ) );
  DFF_X1 \mem_reg[518][2]  ( .D(n21960), .CK(clk), .Q(\mem[518][2] ) );
  DFF_X1 \mem_reg[518][1]  ( .D(n21961), .CK(clk), .Q(\mem[518][1] ) );
  DFF_X1 \mem_reg[518][0]  ( .D(n21962), .CK(clk), .Q(\mem[518][0] ) );
  DFF_X1 \mem_reg[517][7]  ( .D(n21963), .CK(clk), .Q(\mem[517][7] ) );
  DFF_X1 \mem_reg[517][6]  ( .D(n21964), .CK(clk), .Q(\mem[517][6] ) );
  DFF_X1 \mem_reg[517][5]  ( .D(n21965), .CK(clk), .Q(\mem[517][5] ) );
  DFF_X1 \mem_reg[517][4]  ( .D(n21966), .CK(clk), .Q(\mem[517][4] ) );
  DFF_X1 \mem_reg[517][3]  ( .D(n21967), .CK(clk), .Q(\mem[517][3] ) );
  DFF_X1 \mem_reg[517][2]  ( .D(n21968), .CK(clk), .Q(\mem[517][2] ) );
  DFF_X1 \mem_reg[517][1]  ( .D(n21969), .CK(clk), .Q(\mem[517][1] ) );
  DFF_X1 \mem_reg[517][0]  ( .D(n21970), .CK(clk), .Q(\mem[517][0] ) );
  DFF_X1 \mem_reg[516][7]  ( .D(n21971), .CK(clk), .Q(\mem[516][7] ) );
  DFF_X1 \mem_reg[516][6]  ( .D(n21972), .CK(clk), .Q(\mem[516][6] ) );
  DFF_X1 \mem_reg[516][5]  ( .D(n21973), .CK(clk), .Q(\mem[516][5] ) );
  DFF_X1 \mem_reg[516][4]  ( .D(n21974), .CK(clk), .Q(\mem[516][4] ) );
  DFF_X1 \mem_reg[516][3]  ( .D(n21975), .CK(clk), .Q(\mem[516][3] ) );
  DFF_X1 \mem_reg[516][2]  ( .D(n21976), .CK(clk), .Q(\mem[516][2] ) );
  DFF_X1 \mem_reg[516][1]  ( .D(n21977), .CK(clk), .Q(\mem[516][1] ) );
  DFF_X1 \mem_reg[516][0]  ( .D(n21978), .CK(clk), .Q(\mem[516][0] ) );
  DFF_X1 \mem_reg[515][7]  ( .D(n21979), .CK(clk), .Q(\mem[515][7] ) );
  DFF_X1 \mem_reg[515][6]  ( .D(n21980), .CK(clk), .Q(\mem[515][6] ) );
  DFF_X1 \mem_reg[515][5]  ( .D(n21981), .CK(clk), .Q(\mem[515][5] ) );
  DFF_X1 \mem_reg[515][4]  ( .D(n21982), .CK(clk), .Q(\mem[515][4] ) );
  DFF_X1 \mem_reg[515][3]  ( .D(n21983), .CK(clk), .Q(\mem[515][3] ) );
  DFF_X1 \mem_reg[515][2]  ( .D(n21984), .CK(clk), .Q(\mem[515][2] ) );
  DFF_X1 \mem_reg[515][1]  ( .D(n21985), .CK(clk), .Q(\mem[515][1] ) );
  DFF_X1 \mem_reg[515][0]  ( .D(n21986), .CK(clk), .Q(\mem[515][0] ) );
  DFF_X1 \mem_reg[514][7]  ( .D(n21987), .CK(clk), .Q(\mem[514][7] ) );
  DFF_X1 \mem_reg[514][6]  ( .D(n21988), .CK(clk), .Q(\mem[514][6] ) );
  DFF_X1 \mem_reg[514][5]  ( .D(n21989), .CK(clk), .Q(\mem[514][5] ) );
  DFF_X1 \mem_reg[514][4]  ( .D(n21990), .CK(clk), .Q(\mem[514][4] ) );
  DFF_X1 \mem_reg[514][3]  ( .D(n21991), .CK(clk), .Q(\mem[514][3] ) );
  DFF_X1 \mem_reg[514][2]  ( .D(n21992), .CK(clk), .Q(\mem[514][2] ) );
  DFF_X1 \mem_reg[514][1]  ( .D(n21993), .CK(clk), .Q(\mem[514][1] ) );
  DFF_X1 \mem_reg[514][0]  ( .D(n21994), .CK(clk), .Q(\mem[514][0] ) );
  DFF_X1 \mem_reg[513][7]  ( .D(n21995), .CK(clk), .Q(\mem[513][7] ) );
  DFF_X1 \mem_reg[513][6]  ( .D(n21996), .CK(clk), .Q(\mem[513][6] ) );
  DFF_X1 \mem_reg[513][5]  ( .D(n21997), .CK(clk), .Q(\mem[513][5] ) );
  DFF_X1 \mem_reg[513][4]  ( .D(n21998), .CK(clk), .Q(\mem[513][4] ) );
  DFF_X1 \mem_reg[513][3]  ( .D(n21999), .CK(clk), .Q(\mem[513][3] ) );
  DFF_X1 \mem_reg[513][2]  ( .D(n22000), .CK(clk), .Q(\mem[513][2] ) );
  DFF_X1 \mem_reg[513][1]  ( .D(n22001), .CK(clk), .Q(\mem[513][1] ) );
  DFF_X1 \mem_reg[513][0]  ( .D(n22002), .CK(clk), .Q(\mem[513][0] ) );
  DFF_X1 \mem_reg[512][7]  ( .D(n22003), .CK(clk), .Q(\mem[512][7] ) );
  DFF_X1 \mem_reg[512][6]  ( .D(n22004), .CK(clk), .Q(\mem[512][6] ) );
  DFF_X1 \mem_reg[512][5]  ( .D(n22005), .CK(clk), .Q(\mem[512][5] ) );
  DFF_X1 \mem_reg[512][4]  ( .D(n22006), .CK(clk), .Q(\mem[512][4] ) );
  DFF_X1 \mem_reg[512][3]  ( .D(n22007), .CK(clk), .Q(\mem[512][3] ) );
  DFF_X1 \mem_reg[512][2]  ( .D(n22008), .CK(clk), .Q(\mem[512][2] ) );
  DFF_X1 \mem_reg[512][1]  ( .D(n22009), .CK(clk), .Q(\mem[512][1] ) );
  DFF_X1 \mem_reg[512][0]  ( .D(n22010), .CK(clk), .Q(\mem[512][0] ) );
  DFF_X1 \mem_reg[511][7]  ( .D(n22011), .CK(clk), .Q(\mem[511][7] ) );
  DFF_X1 \mem_reg[511][6]  ( .D(n22012), .CK(clk), .Q(\mem[511][6] ) );
  DFF_X1 \mem_reg[511][5]  ( .D(n22013), .CK(clk), .Q(\mem[511][5] ) );
  DFF_X1 \mem_reg[511][4]  ( .D(n22014), .CK(clk), .Q(\mem[511][4] ) );
  DFF_X1 \mem_reg[511][3]  ( .D(n22015), .CK(clk), .Q(\mem[511][3] ) );
  DFF_X1 \mem_reg[511][2]  ( .D(n22016), .CK(clk), .Q(\mem[511][2] ) );
  DFF_X1 \mem_reg[511][1]  ( .D(n22017), .CK(clk), .Q(\mem[511][1] ) );
  DFF_X1 \mem_reg[511][0]  ( .D(n22018), .CK(clk), .Q(\mem[511][0] ) );
  DFF_X1 \mem_reg[510][7]  ( .D(n22019), .CK(clk), .Q(\mem[510][7] ) );
  DFF_X1 \mem_reg[510][6]  ( .D(n22020), .CK(clk), .Q(\mem[510][6] ) );
  DFF_X1 \mem_reg[510][5]  ( .D(n22021), .CK(clk), .Q(\mem[510][5] ) );
  DFF_X1 \mem_reg[510][4]  ( .D(n22022), .CK(clk), .Q(\mem[510][4] ) );
  DFF_X1 \mem_reg[510][3]  ( .D(n22023), .CK(clk), .Q(\mem[510][3] ) );
  DFF_X1 \mem_reg[510][2]  ( .D(n22024), .CK(clk), .Q(\mem[510][2] ) );
  DFF_X1 \mem_reg[510][1]  ( .D(n22025), .CK(clk), .Q(\mem[510][1] ) );
  DFF_X1 \mem_reg[510][0]  ( .D(n22026), .CK(clk), .Q(\mem[510][0] ) );
  DFF_X1 \mem_reg[509][7]  ( .D(n22027), .CK(clk), .Q(\mem[509][7] ) );
  DFF_X1 \mem_reg[509][6]  ( .D(n22028), .CK(clk), .Q(\mem[509][6] ) );
  DFF_X1 \mem_reg[509][5]  ( .D(n22029), .CK(clk), .Q(\mem[509][5] ) );
  DFF_X1 \mem_reg[509][4]  ( .D(n22030), .CK(clk), .Q(\mem[509][4] ) );
  DFF_X1 \mem_reg[509][3]  ( .D(n22031), .CK(clk), .Q(\mem[509][3] ) );
  DFF_X1 \mem_reg[509][2]  ( .D(n22032), .CK(clk), .Q(\mem[509][2] ) );
  DFF_X1 \mem_reg[509][1]  ( .D(n22033), .CK(clk), .Q(\mem[509][1] ) );
  DFF_X1 \mem_reg[509][0]  ( .D(n22034), .CK(clk), .Q(\mem[509][0] ) );
  DFF_X1 \mem_reg[508][7]  ( .D(n22035), .CK(clk), .Q(\mem[508][7] ) );
  DFF_X1 \mem_reg[508][6]  ( .D(n22036), .CK(clk), .Q(\mem[508][6] ) );
  DFF_X1 \mem_reg[508][5]  ( .D(n22037), .CK(clk), .Q(\mem[508][5] ) );
  DFF_X1 \mem_reg[508][4]  ( .D(n22038), .CK(clk), .Q(\mem[508][4] ) );
  DFF_X1 \mem_reg[508][3]  ( .D(n22039), .CK(clk), .Q(\mem[508][3] ) );
  DFF_X1 \mem_reg[508][2]  ( .D(n22040), .CK(clk), .Q(\mem[508][2] ) );
  DFF_X1 \mem_reg[508][1]  ( .D(n22041), .CK(clk), .Q(\mem[508][1] ) );
  DFF_X1 \mem_reg[508][0]  ( .D(n22042), .CK(clk), .Q(\mem[508][0] ) );
  DFF_X1 \mem_reg[507][7]  ( .D(n22043), .CK(clk), .Q(\mem[507][7] ) );
  DFF_X1 \mem_reg[507][6]  ( .D(n22044), .CK(clk), .Q(\mem[507][6] ) );
  DFF_X1 \mem_reg[507][5]  ( .D(n22045), .CK(clk), .Q(\mem[507][5] ) );
  DFF_X1 \mem_reg[507][4]  ( .D(n22046), .CK(clk), .Q(\mem[507][4] ) );
  DFF_X1 \mem_reg[507][3]  ( .D(n22047), .CK(clk), .Q(\mem[507][3] ) );
  DFF_X1 \mem_reg[507][2]  ( .D(n22048), .CK(clk), .Q(\mem[507][2] ) );
  DFF_X1 \mem_reg[507][1]  ( .D(n22049), .CK(clk), .Q(\mem[507][1] ) );
  DFF_X1 \mem_reg[507][0]  ( .D(n22050), .CK(clk), .Q(\mem[507][0] ) );
  DFF_X1 \mem_reg[506][7]  ( .D(n22051), .CK(clk), .Q(\mem[506][7] ) );
  DFF_X1 \mem_reg[506][6]  ( .D(n22052), .CK(clk), .Q(\mem[506][6] ) );
  DFF_X1 \mem_reg[506][5]  ( .D(n22053), .CK(clk), .Q(\mem[506][5] ) );
  DFF_X1 \mem_reg[506][4]  ( .D(n22054), .CK(clk), .Q(\mem[506][4] ) );
  DFF_X1 \mem_reg[506][3]  ( .D(n22055), .CK(clk), .Q(\mem[506][3] ) );
  DFF_X1 \mem_reg[506][2]  ( .D(n22056), .CK(clk), .Q(\mem[506][2] ) );
  DFF_X1 \mem_reg[506][1]  ( .D(n22057), .CK(clk), .Q(\mem[506][1] ) );
  DFF_X1 \mem_reg[506][0]  ( .D(n22058), .CK(clk), .Q(\mem[506][0] ) );
  DFF_X1 \mem_reg[505][7]  ( .D(n22059), .CK(clk), .Q(\mem[505][7] ) );
  DFF_X1 \mem_reg[505][6]  ( .D(n22060), .CK(clk), .Q(\mem[505][6] ) );
  DFF_X1 \mem_reg[505][5]  ( .D(n22061), .CK(clk), .Q(\mem[505][5] ) );
  DFF_X1 \mem_reg[505][4]  ( .D(n22062), .CK(clk), .Q(\mem[505][4] ) );
  DFF_X1 \mem_reg[505][3]  ( .D(n22063), .CK(clk), .Q(\mem[505][3] ) );
  DFF_X1 \mem_reg[505][2]  ( .D(n22064), .CK(clk), .Q(\mem[505][2] ) );
  DFF_X1 \mem_reg[505][1]  ( .D(n22065), .CK(clk), .Q(\mem[505][1] ) );
  DFF_X1 \mem_reg[505][0]  ( .D(n22066), .CK(clk), .Q(\mem[505][0] ) );
  DFF_X1 \mem_reg[504][7]  ( .D(n22067), .CK(clk), .Q(\mem[504][7] ) );
  DFF_X1 \mem_reg[504][6]  ( .D(n22068), .CK(clk), .Q(\mem[504][6] ) );
  DFF_X1 \mem_reg[504][5]  ( .D(n22069), .CK(clk), .Q(\mem[504][5] ) );
  DFF_X1 \mem_reg[504][4]  ( .D(n22070), .CK(clk), .Q(\mem[504][4] ) );
  DFF_X1 \mem_reg[504][3]  ( .D(n22071), .CK(clk), .Q(\mem[504][3] ) );
  DFF_X1 \mem_reg[504][2]  ( .D(n22072), .CK(clk), .Q(\mem[504][2] ) );
  DFF_X1 \mem_reg[504][1]  ( .D(n22073), .CK(clk), .Q(\mem[504][1] ) );
  DFF_X1 \mem_reg[504][0]  ( .D(n22074), .CK(clk), .Q(\mem[504][0] ) );
  DFF_X1 \mem_reg[503][7]  ( .D(n22075), .CK(clk), .Q(\mem[503][7] ) );
  DFF_X1 \mem_reg[503][6]  ( .D(n22076), .CK(clk), .Q(\mem[503][6] ) );
  DFF_X1 \mem_reg[503][5]  ( .D(n22077), .CK(clk), .Q(\mem[503][5] ) );
  DFF_X1 \mem_reg[503][4]  ( .D(n22078), .CK(clk), .Q(\mem[503][4] ) );
  DFF_X1 \mem_reg[503][3]  ( .D(n22079), .CK(clk), .Q(\mem[503][3] ) );
  DFF_X1 \mem_reg[503][2]  ( .D(n22080), .CK(clk), .Q(\mem[503][2] ) );
  DFF_X1 \mem_reg[503][1]  ( .D(n22081), .CK(clk), .Q(\mem[503][1] ) );
  DFF_X1 \mem_reg[503][0]  ( .D(n22082), .CK(clk), .Q(\mem[503][0] ) );
  DFF_X1 \mem_reg[502][7]  ( .D(n22083), .CK(clk), .Q(\mem[502][7] ) );
  DFF_X1 \mem_reg[502][6]  ( .D(n22084), .CK(clk), .Q(\mem[502][6] ) );
  DFF_X1 \mem_reg[502][5]  ( .D(n22085), .CK(clk), .Q(\mem[502][5] ) );
  DFF_X1 \mem_reg[502][4]  ( .D(n22086), .CK(clk), .Q(\mem[502][4] ) );
  DFF_X1 \mem_reg[502][3]  ( .D(n22087), .CK(clk), .Q(\mem[502][3] ) );
  DFF_X1 \mem_reg[502][2]  ( .D(n22088), .CK(clk), .Q(\mem[502][2] ) );
  DFF_X1 \mem_reg[502][1]  ( .D(n22089), .CK(clk), .Q(\mem[502][1] ) );
  DFF_X1 \mem_reg[502][0]  ( .D(n22090), .CK(clk), .Q(\mem[502][0] ) );
  DFF_X1 \mem_reg[501][7]  ( .D(n22091), .CK(clk), .Q(\mem[501][7] ) );
  DFF_X1 \mem_reg[501][6]  ( .D(n22092), .CK(clk), .Q(\mem[501][6] ) );
  DFF_X1 \mem_reg[501][5]  ( .D(n22093), .CK(clk), .Q(\mem[501][5] ) );
  DFF_X1 \mem_reg[501][4]  ( .D(n22094), .CK(clk), .Q(\mem[501][4] ) );
  DFF_X1 \mem_reg[501][3]  ( .D(n22095), .CK(clk), .Q(\mem[501][3] ) );
  DFF_X1 \mem_reg[501][2]  ( .D(n22096), .CK(clk), .Q(\mem[501][2] ) );
  DFF_X1 \mem_reg[501][1]  ( .D(n22097), .CK(clk), .Q(\mem[501][1] ) );
  DFF_X1 \mem_reg[501][0]  ( .D(n22098), .CK(clk), .Q(\mem[501][0] ) );
  DFF_X1 \mem_reg[500][7]  ( .D(n22099), .CK(clk), .Q(\mem[500][7] ) );
  DFF_X1 \mem_reg[500][6]  ( .D(n22100), .CK(clk), .Q(\mem[500][6] ) );
  DFF_X1 \mem_reg[500][5]  ( .D(n22101), .CK(clk), .Q(\mem[500][5] ) );
  DFF_X1 \mem_reg[500][4]  ( .D(n22102), .CK(clk), .Q(\mem[500][4] ) );
  DFF_X1 \mem_reg[500][3]  ( .D(n22103), .CK(clk), .Q(\mem[500][3] ) );
  DFF_X1 \mem_reg[500][2]  ( .D(n22104), .CK(clk), .Q(\mem[500][2] ) );
  DFF_X1 \mem_reg[500][1]  ( .D(n22105), .CK(clk), .Q(\mem[500][1] ) );
  DFF_X1 \mem_reg[500][0]  ( .D(n22106), .CK(clk), .Q(\mem[500][0] ) );
  DFF_X1 \mem_reg[499][7]  ( .D(n22107), .CK(clk), .Q(\mem[499][7] ) );
  DFF_X1 \mem_reg[499][6]  ( .D(n22108), .CK(clk), .Q(\mem[499][6] ) );
  DFF_X1 \mem_reg[499][5]  ( .D(n22109), .CK(clk), .Q(\mem[499][5] ) );
  DFF_X1 \mem_reg[499][4]  ( .D(n22110), .CK(clk), .Q(\mem[499][4] ) );
  DFF_X1 \mem_reg[499][3]  ( .D(n22111), .CK(clk), .Q(\mem[499][3] ) );
  DFF_X1 \mem_reg[499][2]  ( .D(n22112), .CK(clk), .Q(\mem[499][2] ) );
  DFF_X1 \mem_reg[499][1]  ( .D(n22113), .CK(clk), .Q(\mem[499][1] ) );
  DFF_X1 \mem_reg[499][0]  ( .D(n22114), .CK(clk), .Q(\mem[499][0] ) );
  DFF_X1 \mem_reg[498][7]  ( .D(n22115), .CK(clk), .Q(\mem[498][7] ) );
  DFF_X1 \mem_reg[498][6]  ( .D(n22116), .CK(clk), .Q(\mem[498][6] ) );
  DFF_X1 \mem_reg[498][5]  ( .D(n22117), .CK(clk), .Q(\mem[498][5] ) );
  DFF_X1 \mem_reg[498][4]  ( .D(n22118), .CK(clk), .Q(\mem[498][4] ) );
  DFF_X1 \mem_reg[498][3]  ( .D(n22119), .CK(clk), .Q(\mem[498][3] ) );
  DFF_X1 \mem_reg[498][2]  ( .D(n22120), .CK(clk), .Q(\mem[498][2] ) );
  DFF_X1 \mem_reg[498][1]  ( .D(n22121), .CK(clk), .Q(\mem[498][1] ) );
  DFF_X1 \mem_reg[498][0]  ( .D(n22122), .CK(clk), .Q(\mem[498][0] ) );
  DFF_X1 \mem_reg[497][7]  ( .D(n22123), .CK(clk), .Q(\mem[497][7] ) );
  DFF_X1 \mem_reg[497][6]  ( .D(n22124), .CK(clk), .Q(\mem[497][6] ) );
  DFF_X1 \mem_reg[497][5]  ( .D(n22125), .CK(clk), .Q(\mem[497][5] ) );
  DFF_X1 \mem_reg[497][4]  ( .D(n22126), .CK(clk), .Q(\mem[497][4] ) );
  DFF_X1 \mem_reg[497][3]  ( .D(n22127), .CK(clk), .Q(\mem[497][3] ) );
  DFF_X1 \mem_reg[497][2]  ( .D(n22128), .CK(clk), .Q(\mem[497][2] ) );
  DFF_X1 \mem_reg[497][1]  ( .D(n22129), .CK(clk), .Q(\mem[497][1] ) );
  DFF_X1 \mem_reg[497][0]  ( .D(n22130), .CK(clk), .Q(\mem[497][0] ) );
  DFF_X1 \mem_reg[496][7]  ( .D(n22131), .CK(clk), .Q(\mem[496][7] ) );
  DFF_X1 \mem_reg[496][6]  ( .D(n22132), .CK(clk), .Q(\mem[496][6] ) );
  DFF_X1 \mem_reg[496][5]  ( .D(n22133), .CK(clk), .Q(\mem[496][5] ) );
  DFF_X1 \mem_reg[496][4]  ( .D(n22134), .CK(clk), .Q(\mem[496][4] ) );
  DFF_X1 \mem_reg[496][3]  ( .D(n22135), .CK(clk), .Q(\mem[496][3] ) );
  DFF_X1 \mem_reg[496][2]  ( .D(n22136), .CK(clk), .Q(\mem[496][2] ) );
  DFF_X1 \mem_reg[496][1]  ( .D(n22137), .CK(clk), .Q(\mem[496][1] ) );
  DFF_X1 \mem_reg[496][0]  ( .D(n22138), .CK(clk), .Q(\mem[496][0] ) );
  DFF_X1 \mem_reg[495][7]  ( .D(n22139), .CK(clk), .Q(\mem[495][7] ) );
  DFF_X1 \mem_reg[495][6]  ( .D(n22140), .CK(clk), .Q(\mem[495][6] ) );
  DFF_X1 \mem_reg[495][5]  ( .D(n22141), .CK(clk), .Q(\mem[495][5] ) );
  DFF_X1 \mem_reg[495][4]  ( .D(n22142), .CK(clk), .Q(\mem[495][4] ) );
  DFF_X1 \mem_reg[495][3]  ( .D(n22143), .CK(clk), .Q(\mem[495][3] ) );
  DFF_X1 \mem_reg[495][2]  ( .D(n22144), .CK(clk), .Q(\mem[495][2] ) );
  DFF_X1 \mem_reg[495][1]  ( .D(n22145), .CK(clk), .Q(\mem[495][1] ) );
  DFF_X1 \mem_reg[495][0]  ( .D(n22146), .CK(clk), .Q(\mem[495][0] ) );
  DFF_X1 \mem_reg[494][7]  ( .D(n22147), .CK(clk), .Q(\mem[494][7] ) );
  DFF_X1 \mem_reg[494][6]  ( .D(n22148), .CK(clk), .Q(\mem[494][6] ) );
  DFF_X1 \mem_reg[494][5]  ( .D(n22149), .CK(clk), .Q(\mem[494][5] ) );
  DFF_X1 \mem_reg[494][4]  ( .D(n22150), .CK(clk), .Q(\mem[494][4] ) );
  DFF_X1 \mem_reg[494][3]  ( .D(n22151), .CK(clk), .Q(\mem[494][3] ) );
  DFF_X1 \mem_reg[494][2]  ( .D(n22152), .CK(clk), .Q(\mem[494][2] ) );
  DFF_X1 \mem_reg[494][1]  ( .D(n22153), .CK(clk), .Q(\mem[494][1] ) );
  DFF_X1 \mem_reg[494][0]  ( .D(n22154), .CK(clk), .Q(\mem[494][0] ) );
  DFF_X1 \mem_reg[493][7]  ( .D(n22155), .CK(clk), .Q(\mem[493][7] ) );
  DFF_X1 \mem_reg[493][6]  ( .D(n22156), .CK(clk), .Q(\mem[493][6] ) );
  DFF_X1 \mem_reg[493][5]  ( .D(n22157), .CK(clk), .Q(\mem[493][5] ) );
  DFF_X1 \mem_reg[493][4]  ( .D(n22158), .CK(clk), .Q(\mem[493][4] ) );
  DFF_X1 \mem_reg[493][3]  ( .D(n22159), .CK(clk), .Q(\mem[493][3] ) );
  DFF_X1 \mem_reg[493][2]  ( .D(n22160), .CK(clk), .Q(\mem[493][2] ) );
  DFF_X1 \mem_reg[493][1]  ( .D(n22161), .CK(clk), .Q(\mem[493][1] ) );
  DFF_X1 \mem_reg[493][0]  ( .D(n22162), .CK(clk), .Q(\mem[493][0] ) );
  DFF_X1 \mem_reg[492][7]  ( .D(n22163), .CK(clk), .Q(\mem[492][7] ) );
  DFF_X1 \mem_reg[492][6]  ( .D(n22164), .CK(clk), .Q(\mem[492][6] ) );
  DFF_X1 \mem_reg[492][5]  ( .D(n22165), .CK(clk), .Q(\mem[492][5] ) );
  DFF_X1 \mem_reg[492][4]  ( .D(n22166), .CK(clk), .Q(\mem[492][4] ) );
  DFF_X1 \mem_reg[492][3]  ( .D(n22167), .CK(clk), .Q(\mem[492][3] ) );
  DFF_X1 \mem_reg[492][2]  ( .D(n22168), .CK(clk), .Q(\mem[492][2] ) );
  DFF_X1 \mem_reg[492][1]  ( .D(n22169), .CK(clk), .Q(\mem[492][1] ) );
  DFF_X1 \mem_reg[492][0]  ( .D(n22170), .CK(clk), .Q(\mem[492][0] ) );
  DFF_X1 \mem_reg[491][7]  ( .D(n22171), .CK(clk), .Q(\mem[491][7] ) );
  DFF_X1 \mem_reg[491][6]  ( .D(n22172), .CK(clk), .Q(\mem[491][6] ) );
  DFF_X1 \mem_reg[491][5]  ( .D(n22173), .CK(clk), .Q(\mem[491][5] ) );
  DFF_X1 \mem_reg[491][4]  ( .D(n22174), .CK(clk), .Q(\mem[491][4] ) );
  DFF_X1 \mem_reg[491][3]  ( .D(n22175), .CK(clk), .Q(\mem[491][3] ) );
  DFF_X1 \mem_reg[491][2]  ( .D(n22176), .CK(clk), .Q(\mem[491][2] ) );
  DFF_X1 \mem_reg[491][1]  ( .D(n22177), .CK(clk), .Q(\mem[491][1] ) );
  DFF_X1 \mem_reg[491][0]  ( .D(n22178), .CK(clk), .Q(\mem[491][0] ) );
  DFF_X1 \mem_reg[490][7]  ( .D(n22179), .CK(clk), .Q(\mem[490][7] ) );
  DFF_X1 \mem_reg[490][6]  ( .D(n22180), .CK(clk), .Q(\mem[490][6] ) );
  DFF_X1 \mem_reg[490][5]  ( .D(n22181), .CK(clk), .Q(\mem[490][5] ) );
  DFF_X1 \mem_reg[490][4]  ( .D(n22182), .CK(clk), .Q(\mem[490][4] ) );
  DFF_X1 \mem_reg[490][3]  ( .D(n22183), .CK(clk), .Q(\mem[490][3] ) );
  DFF_X1 \mem_reg[490][2]  ( .D(n22184), .CK(clk), .Q(\mem[490][2] ) );
  DFF_X1 \mem_reg[490][1]  ( .D(n22185), .CK(clk), .Q(\mem[490][1] ) );
  DFF_X1 \mem_reg[490][0]  ( .D(n22186), .CK(clk), .Q(\mem[490][0] ) );
  DFF_X1 \mem_reg[489][7]  ( .D(n22187), .CK(clk), .Q(\mem[489][7] ) );
  DFF_X1 \mem_reg[489][6]  ( .D(n22188), .CK(clk), .Q(\mem[489][6] ) );
  DFF_X1 \mem_reg[489][5]  ( .D(n22189), .CK(clk), .Q(\mem[489][5] ) );
  DFF_X1 \mem_reg[489][4]  ( .D(n22190), .CK(clk), .Q(\mem[489][4] ) );
  DFF_X1 \mem_reg[489][3]  ( .D(n22191), .CK(clk), .Q(\mem[489][3] ) );
  DFF_X1 \mem_reg[489][2]  ( .D(n22192), .CK(clk), .Q(\mem[489][2] ) );
  DFF_X1 \mem_reg[489][1]  ( .D(n22193), .CK(clk), .Q(\mem[489][1] ) );
  DFF_X1 \mem_reg[489][0]  ( .D(n22194), .CK(clk), .Q(\mem[489][0] ) );
  DFF_X1 \mem_reg[488][7]  ( .D(n22195), .CK(clk), .Q(\mem[488][7] ) );
  DFF_X1 \mem_reg[488][6]  ( .D(n22196), .CK(clk), .Q(\mem[488][6] ) );
  DFF_X1 \mem_reg[488][5]  ( .D(n22197), .CK(clk), .Q(\mem[488][5] ) );
  DFF_X1 \mem_reg[488][4]  ( .D(n22198), .CK(clk), .Q(\mem[488][4] ) );
  DFF_X1 \mem_reg[488][3]  ( .D(n22199), .CK(clk), .Q(\mem[488][3] ) );
  DFF_X1 \mem_reg[488][2]  ( .D(n22200), .CK(clk), .Q(\mem[488][2] ) );
  DFF_X1 \mem_reg[488][1]  ( .D(n22201), .CK(clk), .Q(\mem[488][1] ) );
  DFF_X1 \mem_reg[488][0]  ( .D(n22202), .CK(clk), .Q(\mem[488][0] ) );
  DFF_X1 \mem_reg[487][7]  ( .D(n22203), .CK(clk), .Q(\mem[487][7] ) );
  DFF_X1 \mem_reg[487][6]  ( .D(n22204), .CK(clk), .Q(\mem[487][6] ) );
  DFF_X1 \mem_reg[487][5]  ( .D(n22205), .CK(clk), .Q(\mem[487][5] ) );
  DFF_X1 \mem_reg[487][4]  ( .D(n22206), .CK(clk), .Q(\mem[487][4] ) );
  DFF_X1 \mem_reg[487][3]  ( .D(n22207), .CK(clk), .Q(\mem[487][3] ) );
  DFF_X1 \mem_reg[487][2]  ( .D(n22208), .CK(clk), .Q(\mem[487][2] ) );
  DFF_X1 \mem_reg[487][1]  ( .D(n22209), .CK(clk), .Q(\mem[487][1] ) );
  DFF_X1 \mem_reg[487][0]  ( .D(n22210), .CK(clk), .Q(\mem[487][0] ) );
  DFF_X1 \mem_reg[486][7]  ( .D(n22211), .CK(clk), .Q(\mem[486][7] ) );
  DFF_X1 \mem_reg[486][6]  ( .D(n22212), .CK(clk), .Q(\mem[486][6] ) );
  DFF_X1 \mem_reg[486][5]  ( .D(n22213), .CK(clk), .Q(\mem[486][5] ) );
  DFF_X1 \mem_reg[486][4]  ( .D(n22214), .CK(clk), .Q(\mem[486][4] ) );
  DFF_X1 \mem_reg[486][3]  ( .D(n22215), .CK(clk), .Q(\mem[486][3] ) );
  DFF_X1 \mem_reg[486][2]  ( .D(n22216), .CK(clk), .Q(\mem[486][2] ) );
  DFF_X1 \mem_reg[486][1]  ( .D(n22217), .CK(clk), .Q(\mem[486][1] ) );
  DFF_X1 \mem_reg[486][0]  ( .D(n22218), .CK(clk), .Q(\mem[486][0] ) );
  DFF_X1 \mem_reg[485][7]  ( .D(n22219), .CK(clk), .Q(\mem[485][7] ) );
  DFF_X1 \mem_reg[485][6]  ( .D(n22220), .CK(clk), .Q(\mem[485][6] ) );
  DFF_X1 \mem_reg[485][5]  ( .D(n22221), .CK(clk), .Q(\mem[485][5] ) );
  DFF_X1 \mem_reg[485][4]  ( .D(n22222), .CK(clk), .Q(\mem[485][4] ) );
  DFF_X1 \mem_reg[485][3]  ( .D(n22223), .CK(clk), .Q(\mem[485][3] ) );
  DFF_X1 \mem_reg[485][2]  ( .D(n22224), .CK(clk), .Q(\mem[485][2] ) );
  DFF_X1 \mem_reg[485][1]  ( .D(n22225), .CK(clk), .Q(\mem[485][1] ) );
  DFF_X1 \mem_reg[485][0]  ( .D(n22226), .CK(clk), .Q(\mem[485][0] ) );
  DFF_X1 \mem_reg[484][7]  ( .D(n22227), .CK(clk), .Q(\mem[484][7] ) );
  DFF_X1 \mem_reg[484][6]  ( .D(n22228), .CK(clk), .Q(\mem[484][6] ) );
  DFF_X1 \mem_reg[484][5]  ( .D(n22229), .CK(clk), .Q(\mem[484][5] ) );
  DFF_X1 \mem_reg[484][4]  ( .D(n22230), .CK(clk), .Q(\mem[484][4] ) );
  DFF_X1 \mem_reg[484][3]  ( .D(n22231), .CK(clk), .Q(\mem[484][3] ) );
  DFF_X1 \mem_reg[484][2]  ( .D(n22232), .CK(clk), .Q(\mem[484][2] ) );
  DFF_X1 \mem_reg[484][1]  ( .D(n22233), .CK(clk), .Q(\mem[484][1] ) );
  DFF_X1 \mem_reg[484][0]  ( .D(n22234), .CK(clk), .Q(\mem[484][0] ) );
  DFF_X1 \mem_reg[483][7]  ( .D(n22235), .CK(clk), .Q(\mem[483][7] ) );
  DFF_X1 \mem_reg[483][6]  ( .D(n22236), .CK(clk), .Q(\mem[483][6] ) );
  DFF_X1 \mem_reg[483][5]  ( .D(n22237), .CK(clk), .Q(\mem[483][5] ) );
  DFF_X1 \mem_reg[483][4]  ( .D(n22238), .CK(clk), .Q(\mem[483][4] ) );
  DFF_X1 \mem_reg[483][3]  ( .D(n22239), .CK(clk), .Q(\mem[483][3] ) );
  DFF_X1 \mem_reg[483][2]  ( .D(n22240), .CK(clk), .Q(\mem[483][2] ) );
  DFF_X1 \mem_reg[483][1]  ( .D(n22241), .CK(clk), .Q(\mem[483][1] ) );
  DFF_X1 \mem_reg[483][0]  ( .D(n22242), .CK(clk), .Q(\mem[483][0] ) );
  DFF_X1 \mem_reg[482][7]  ( .D(n22243), .CK(clk), .Q(\mem[482][7] ) );
  DFF_X1 \mem_reg[482][6]  ( .D(n22244), .CK(clk), .Q(\mem[482][6] ) );
  DFF_X1 \mem_reg[482][5]  ( .D(n22245), .CK(clk), .Q(\mem[482][5] ) );
  DFF_X1 \mem_reg[482][4]  ( .D(n22246), .CK(clk), .Q(\mem[482][4] ) );
  DFF_X1 \mem_reg[482][3]  ( .D(n22247), .CK(clk), .Q(\mem[482][3] ) );
  DFF_X1 \mem_reg[482][2]  ( .D(n22248), .CK(clk), .Q(\mem[482][2] ) );
  DFF_X1 \mem_reg[482][1]  ( .D(n22249), .CK(clk), .Q(\mem[482][1] ) );
  DFF_X1 \mem_reg[482][0]  ( .D(n22250), .CK(clk), .Q(\mem[482][0] ) );
  DFF_X1 \mem_reg[481][7]  ( .D(n22251), .CK(clk), .Q(\mem[481][7] ) );
  DFF_X1 \mem_reg[481][6]  ( .D(n22252), .CK(clk), .Q(\mem[481][6] ) );
  DFF_X1 \mem_reg[481][5]  ( .D(n22253), .CK(clk), .Q(\mem[481][5] ) );
  DFF_X1 \mem_reg[481][4]  ( .D(n22254), .CK(clk), .Q(\mem[481][4] ) );
  DFF_X1 \mem_reg[481][3]  ( .D(n22255), .CK(clk), .Q(\mem[481][3] ) );
  DFF_X1 \mem_reg[481][2]  ( .D(n22256), .CK(clk), .Q(\mem[481][2] ) );
  DFF_X1 \mem_reg[481][1]  ( .D(n22257), .CK(clk), .Q(\mem[481][1] ) );
  DFF_X1 \mem_reg[481][0]  ( .D(n22258), .CK(clk), .Q(\mem[481][0] ) );
  DFF_X1 \mem_reg[480][7]  ( .D(n22259), .CK(clk), .Q(\mem[480][7] ) );
  DFF_X1 \mem_reg[480][6]  ( .D(n22260), .CK(clk), .Q(\mem[480][6] ) );
  DFF_X1 \mem_reg[480][5]  ( .D(n22261), .CK(clk), .Q(\mem[480][5] ) );
  DFF_X1 \mem_reg[480][4]  ( .D(n22262), .CK(clk), .Q(\mem[480][4] ) );
  DFF_X1 \mem_reg[480][3]  ( .D(n22263), .CK(clk), .Q(\mem[480][3] ) );
  DFF_X1 \mem_reg[480][2]  ( .D(n22264), .CK(clk), .Q(\mem[480][2] ) );
  DFF_X1 \mem_reg[480][1]  ( .D(n22265), .CK(clk), .Q(\mem[480][1] ) );
  DFF_X1 \mem_reg[480][0]  ( .D(n22266), .CK(clk), .Q(\mem[480][0] ) );
  DFF_X1 \mem_reg[479][7]  ( .D(n22267), .CK(clk), .Q(\mem[479][7] ) );
  DFF_X1 \mem_reg[479][6]  ( .D(n22268), .CK(clk), .Q(\mem[479][6] ) );
  DFF_X1 \mem_reg[479][5]  ( .D(n22269), .CK(clk), .Q(\mem[479][5] ) );
  DFF_X1 \mem_reg[479][4]  ( .D(n22270), .CK(clk), .Q(\mem[479][4] ) );
  DFF_X1 \mem_reg[479][3]  ( .D(n22271), .CK(clk), .Q(\mem[479][3] ) );
  DFF_X1 \mem_reg[479][2]  ( .D(n22272), .CK(clk), .Q(\mem[479][2] ) );
  DFF_X1 \mem_reg[479][1]  ( .D(n22273), .CK(clk), .Q(\mem[479][1] ) );
  DFF_X1 \mem_reg[479][0]  ( .D(n22274), .CK(clk), .Q(\mem[479][0] ) );
  DFF_X1 \mem_reg[478][7]  ( .D(n22275), .CK(clk), .Q(\mem[478][7] ) );
  DFF_X1 \mem_reg[478][6]  ( .D(n22276), .CK(clk), .Q(\mem[478][6] ) );
  DFF_X1 \mem_reg[478][5]  ( .D(n22277), .CK(clk), .Q(\mem[478][5] ) );
  DFF_X1 \mem_reg[478][4]  ( .D(n22278), .CK(clk), .Q(\mem[478][4] ) );
  DFF_X1 \mem_reg[478][3]  ( .D(n22279), .CK(clk), .Q(\mem[478][3] ) );
  DFF_X1 \mem_reg[478][2]  ( .D(n22280), .CK(clk), .Q(\mem[478][2] ) );
  DFF_X1 \mem_reg[478][1]  ( .D(n22281), .CK(clk), .Q(\mem[478][1] ) );
  DFF_X1 \mem_reg[478][0]  ( .D(n22282), .CK(clk), .Q(\mem[478][0] ) );
  DFF_X1 \mem_reg[477][7]  ( .D(n22283), .CK(clk), .Q(\mem[477][7] ) );
  DFF_X1 \mem_reg[477][6]  ( .D(n22284), .CK(clk), .Q(\mem[477][6] ) );
  DFF_X1 \mem_reg[477][5]  ( .D(n22285), .CK(clk), .Q(\mem[477][5] ) );
  DFF_X1 \mem_reg[477][4]  ( .D(n22286), .CK(clk), .Q(\mem[477][4] ) );
  DFF_X1 \mem_reg[477][3]  ( .D(n22287), .CK(clk), .Q(\mem[477][3] ) );
  DFF_X1 \mem_reg[477][2]  ( .D(n22288), .CK(clk), .Q(\mem[477][2] ) );
  DFF_X1 \mem_reg[477][1]  ( .D(n22289), .CK(clk), .Q(\mem[477][1] ) );
  DFF_X1 \mem_reg[477][0]  ( .D(n22290), .CK(clk), .Q(\mem[477][0] ) );
  DFF_X1 \mem_reg[476][7]  ( .D(n22291), .CK(clk), .Q(\mem[476][7] ) );
  DFF_X1 \mem_reg[476][6]  ( .D(n22292), .CK(clk), .Q(\mem[476][6] ) );
  DFF_X1 \mem_reg[476][5]  ( .D(n22293), .CK(clk), .Q(\mem[476][5] ) );
  DFF_X1 \mem_reg[476][4]  ( .D(n22294), .CK(clk), .Q(\mem[476][4] ) );
  DFF_X1 \mem_reg[476][3]  ( .D(n22295), .CK(clk), .Q(\mem[476][3] ) );
  DFF_X1 \mem_reg[476][2]  ( .D(n22296), .CK(clk), .Q(\mem[476][2] ) );
  DFF_X1 \mem_reg[476][1]  ( .D(n22297), .CK(clk), .Q(\mem[476][1] ) );
  DFF_X1 \mem_reg[476][0]  ( .D(n22298), .CK(clk), .Q(\mem[476][0] ) );
  DFF_X1 \mem_reg[475][7]  ( .D(n22299), .CK(clk), .Q(\mem[475][7] ) );
  DFF_X1 \mem_reg[475][6]  ( .D(n22300), .CK(clk), .Q(\mem[475][6] ) );
  DFF_X1 \mem_reg[475][5]  ( .D(n22301), .CK(clk), .Q(\mem[475][5] ) );
  DFF_X1 \mem_reg[475][4]  ( .D(n22302), .CK(clk), .Q(\mem[475][4] ) );
  DFF_X1 \mem_reg[475][3]  ( .D(n22303), .CK(clk), .Q(\mem[475][3] ) );
  DFF_X1 \mem_reg[475][2]  ( .D(n22304), .CK(clk), .Q(\mem[475][2] ) );
  DFF_X1 \mem_reg[475][1]  ( .D(n22305), .CK(clk), .Q(\mem[475][1] ) );
  DFF_X1 \mem_reg[475][0]  ( .D(n22306), .CK(clk), .Q(\mem[475][0] ) );
  DFF_X1 \mem_reg[474][7]  ( .D(n22307), .CK(clk), .Q(\mem[474][7] ) );
  DFF_X1 \mem_reg[474][6]  ( .D(n22308), .CK(clk), .Q(\mem[474][6] ) );
  DFF_X1 \mem_reg[474][5]  ( .D(n22309), .CK(clk), .Q(\mem[474][5] ) );
  DFF_X1 \mem_reg[474][4]  ( .D(n22310), .CK(clk), .Q(\mem[474][4] ) );
  DFF_X1 \mem_reg[474][3]  ( .D(n22311), .CK(clk), .Q(\mem[474][3] ) );
  DFF_X1 \mem_reg[474][2]  ( .D(n22312), .CK(clk), .Q(\mem[474][2] ) );
  DFF_X1 \mem_reg[474][1]  ( .D(n22313), .CK(clk), .Q(\mem[474][1] ) );
  DFF_X1 \mem_reg[474][0]  ( .D(n22314), .CK(clk), .Q(\mem[474][0] ) );
  DFF_X1 \mem_reg[473][7]  ( .D(n22315), .CK(clk), .Q(\mem[473][7] ) );
  DFF_X1 \mem_reg[473][6]  ( .D(n22316), .CK(clk), .Q(\mem[473][6] ) );
  DFF_X1 \mem_reg[473][5]  ( .D(n22317), .CK(clk), .Q(\mem[473][5] ) );
  DFF_X1 \mem_reg[473][4]  ( .D(n22318), .CK(clk), .Q(\mem[473][4] ) );
  DFF_X1 \mem_reg[473][3]  ( .D(n22319), .CK(clk), .Q(\mem[473][3] ) );
  DFF_X1 \mem_reg[473][2]  ( .D(n22320), .CK(clk), .Q(\mem[473][2] ) );
  DFF_X1 \mem_reg[473][1]  ( .D(n22321), .CK(clk), .Q(\mem[473][1] ) );
  DFF_X1 \mem_reg[473][0]  ( .D(n22322), .CK(clk), .Q(\mem[473][0] ) );
  DFF_X1 \mem_reg[472][7]  ( .D(n22323), .CK(clk), .Q(\mem[472][7] ) );
  DFF_X1 \mem_reg[472][6]  ( .D(n22324), .CK(clk), .Q(\mem[472][6] ) );
  DFF_X1 \mem_reg[472][5]  ( .D(n22325), .CK(clk), .Q(\mem[472][5] ) );
  DFF_X1 \mem_reg[472][4]  ( .D(n22326), .CK(clk), .Q(\mem[472][4] ) );
  DFF_X1 \mem_reg[472][3]  ( .D(n22327), .CK(clk), .Q(\mem[472][3] ) );
  DFF_X1 \mem_reg[472][2]  ( .D(n22328), .CK(clk), .Q(\mem[472][2] ) );
  DFF_X1 \mem_reg[472][1]  ( .D(n22329), .CK(clk), .Q(\mem[472][1] ) );
  DFF_X1 \mem_reg[472][0]  ( .D(n22330), .CK(clk), .Q(\mem[472][0] ) );
  DFF_X1 \mem_reg[471][7]  ( .D(n22331), .CK(clk), .Q(\mem[471][7] ) );
  DFF_X1 \mem_reg[471][6]  ( .D(n22332), .CK(clk), .Q(\mem[471][6] ) );
  DFF_X1 \mem_reg[471][5]  ( .D(n22333), .CK(clk), .Q(\mem[471][5] ) );
  DFF_X1 \mem_reg[471][4]  ( .D(n22334), .CK(clk), .Q(\mem[471][4] ) );
  DFF_X1 \mem_reg[471][3]  ( .D(n22335), .CK(clk), .Q(\mem[471][3] ) );
  DFF_X1 \mem_reg[471][2]  ( .D(n22336), .CK(clk), .Q(\mem[471][2] ) );
  DFF_X1 \mem_reg[471][1]  ( .D(n22337), .CK(clk), .Q(\mem[471][1] ) );
  DFF_X1 \mem_reg[471][0]  ( .D(n22338), .CK(clk), .Q(\mem[471][0] ) );
  DFF_X1 \mem_reg[470][7]  ( .D(n22339), .CK(clk), .Q(\mem[470][7] ) );
  DFF_X1 \mem_reg[470][6]  ( .D(n22340), .CK(clk), .Q(\mem[470][6] ) );
  DFF_X1 \mem_reg[470][5]  ( .D(n22341), .CK(clk), .Q(\mem[470][5] ) );
  DFF_X1 \mem_reg[470][4]  ( .D(n22342), .CK(clk), .Q(\mem[470][4] ) );
  DFF_X1 \mem_reg[470][3]  ( .D(n22343), .CK(clk), .Q(\mem[470][3] ) );
  DFF_X1 \mem_reg[470][2]  ( .D(n22344), .CK(clk), .Q(\mem[470][2] ) );
  DFF_X1 \mem_reg[470][1]  ( .D(n22345), .CK(clk), .Q(\mem[470][1] ) );
  DFF_X1 \mem_reg[470][0]  ( .D(n22346), .CK(clk), .Q(\mem[470][0] ) );
  DFF_X1 \mem_reg[469][7]  ( .D(n22347), .CK(clk), .Q(\mem[469][7] ) );
  DFF_X1 \mem_reg[469][6]  ( .D(n22348), .CK(clk), .Q(\mem[469][6] ) );
  DFF_X1 \mem_reg[469][5]  ( .D(n22349), .CK(clk), .Q(\mem[469][5] ) );
  DFF_X1 \mem_reg[469][4]  ( .D(n22350), .CK(clk), .Q(\mem[469][4] ) );
  DFF_X1 \mem_reg[469][3]  ( .D(n22351), .CK(clk), .Q(\mem[469][3] ) );
  DFF_X1 \mem_reg[469][2]  ( .D(n22352), .CK(clk), .Q(\mem[469][2] ) );
  DFF_X1 \mem_reg[469][1]  ( .D(n22353), .CK(clk), .Q(\mem[469][1] ) );
  DFF_X1 \mem_reg[469][0]  ( .D(n22354), .CK(clk), .Q(\mem[469][0] ) );
  DFF_X1 \mem_reg[468][7]  ( .D(n22355), .CK(clk), .Q(\mem[468][7] ) );
  DFF_X1 \mem_reg[468][6]  ( .D(n22356), .CK(clk), .Q(\mem[468][6] ) );
  DFF_X1 \mem_reg[468][5]  ( .D(n22357), .CK(clk), .Q(\mem[468][5] ) );
  DFF_X1 \mem_reg[468][4]  ( .D(n22358), .CK(clk), .Q(\mem[468][4] ) );
  DFF_X1 \mem_reg[468][3]  ( .D(n22359), .CK(clk), .Q(\mem[468][3] ) );
  DFF_X1 \mem_reg[468][2]  ( .D(n22360), .CK(clk), .Q(\mem[468][2] ) );
  DFF_X1 \mem_reg[468][1]  ( .D(n22361), .CK(clk), .Q(\mem[468][1] ) );
  DFF_X1 \mem_reg[468][0]  ( .D(n22362), .CK(clk), .Q(\mem[468][0] ) );
  DFF_X1 \mem_reg[467][7]  ( .D(n22363), .CK(clk), .Q(\mem[467][7] ) );
  DFF_X1 \mem_reg[467][6]  ( .D(n22364), .CK(clk), .Q(\mem[467][6] ) );
  DFF_X1 \mem_reg[467][5]  ( .D(n22365), .CK(clk), .Q(\mem[467][5] ) );
  DFF_X1 \mem_reg[467][4]  ( .D(n22366), .CK(clk), .Q(\mem[467][4] ) );
  DFF_X1 \mem_reg[467][3]  ( .D(n22367), .CK(clk), .Q(\mem[467][3] ) );
  DFF_X1 \mem_reg[467][2]  ( .D(n22368), .CK(clk), .Q(\mem[467][2] ) );
  DFF_X1 \mem_reg[467][1]  ( .D(n22369), .CK(clk), .Q(\mem[467][1] ) );
  DFF_X1 \mem_reg[467][0]  ( .D(n22370), .CK(clk), .Q(\mem[467][0] ) );
  DFF_X1 \mem_reg[466][7]  ( .D(n22371), .CK(clk), .Q(\mem[466][7] ) );
  DFF_X1 \mem_reg[466][6]  ( .D(n22372), .CK(clk), .Q(\mem[466][6] ) );
  DFF_X1 \mem_reg[466][5]  ( .D(n22373), .CK(clk), .Q(\mem[466][5] ) );
  DFF_X1 \mem_reg[466][4]  ( .D(n22374), .CK(clk), .Q(\mem[466][4] ) );
  DFF_X1 \mem_reg[466][3]  ( .D(n22375), .CK(clk), .Q(\mem[466][3] ) );
  DFF_X1 \mem_reg[466][2]  ( .D(n22376), .CK(clk), .Q(\mem[466][2] ) );
  DFF_X1 \mem_reg[466][1]  ( .D(n22377), .CK(clk), .Q(\mem[466][1] ) );
  DFF_X1 \mem_reg[466][0]  ( .D(n22378), .CK(clk), .Q(\mem[466][0] ) );
  DFF_X1 \mem_reg[465][7]  ( .D(n22379), .CK(clk), .Q(\mem[465][7] ) );
  DFF_X1 \mem_reg[465][6]  ( .D(n22380), .CK(clk), .Q(\mem[465][6] ) );
  DFF_X1 \mem_reg[465][5]  ( .D(n22381), .CK(clk), .Q(\mem[465][5] ) );
  DFF_X1 \mem_reg[465][4]  ( .D(n22382), .CK(clk), .Q(\mem[465][4] ) );
  DFF_X1 \mem_reg[465][3]  ( .D(n22383), .CK(clk), .Q(\mem[465][3] ) );
  DFF_X1 \mem_reg[465][2]  ( .D(n22384), .CK(clk), .Q(\mem[465][2] ) );
  DFF_X1 \mem_reg[465][1]  ( .D(n22385), .CK(clk), .Q(\mem[465][1] ) );
  DFF_X1 \mem_reg[465][0]  ( .D(n22386), .CK(clk), .Q(\mem[465][0] ) );
  DFF_X1 \mem_reg[464][7]  ( .D(n22387), .CK(clk), .Q(\mem[464][7] ) );
  DFF_X1 \mem_reg[464][6]  ( .D(n22388), .CK(clk), .Q(\mem[464][6] ) );
  DFF_X1 \mem_reg[464][5]  ( .D(n22389), .CK(clk), .Q(\mem[464][5] ) );
  DFF_X1 \mem_reg[464][4]  ( .D(n22390), .CK(clk), .Q(\mem[464][4] ) );
  DFF_X1 \mem_reg[464][3]  ( .D(n22391), .CK(clk), .Q(\mem[464][3] ) );
  DFF_X1 \mem_reg[464][2]  ( .D(n22392), .CK(clk), .Q(\mem[464][2] ) );
  DFF_X1 \mem_reg[464][1]  ( .D(n22393), .CK(clk), .Q(\mem[464][1] ) );
  DFF_X1 \mem_reg[464][0]  ( .D(n22394), .CK(clk), .Q(\mem[464][0] ) );
  DFF_X1 \mem_reg[463][7]  ( .D(n22395), .CK(clk), .Q(\mem[463][7] ) );
  DFF_X1 \mem_reg[463][6]  ( .D(n22396), .CK(clk), .Q(\mem[463][6] ) );
  DFF_X1 \mem_reg[463][5]  ( .D(n22397), .CK(clk), .Q(\mem[463][5] ) );
  DFF_X1 \mem_reg[463][4]  ( .D(n22398), .CK(clk), .Q(\mem[463][4] ) );
  DFF_X1 \mem_reg[463][3]  ( .D(n22399), .CK(clk), .Q(\mem[463][3] ) );
  DFF_X1 \mem_reg[463][2]  ( .D(n22400), .CK(clk), .Q(\mem[463][2] ) );
  DFF_X1 \mem_reg[463][1]  ( .D(n22401), .CK(clk), .Q(\mem[463][1] ) );
  DFF_X1 \mem_reg[463][0]  ( .D(n22402), .CK(clk), .Q(\mem[463][0] ) );
  DFF_X1 \mem_reg[462][7]  ( .D(n22403), .CK(clk), .Q(\mem[462][7] ) );
  DFF_X1 \mem_reg[462][6]  ( .D(n22404), .CK(clk), .Q(\mem[462][6] ) );
  DFF_X1 \mem_reg[462][5]  ( .D(n22405), .CK(clk), .Q(\mem[462][5] ) );
  DFF_X1 \mem_reg[462][4]  ( .D(n22406), .CK(clk), .Q(\mem[462][4] ) );
  DFF_X1 \mem_reg[462][3]  ( .D(n22407), .CK(clk), .Q(\mem[462][3] ) );
  DFF_X1 \mem_reg[462][2]  ( .D(n22408), .CK(clk), .Q(\mem[462][2] ) );
  DFF_X1 \mem_reg[462][1]  ( .D(n22409), .CK(clk), .Q(\mem[462][1] ) );
  DFF_X1 \mem_reg[462][0]  ( .D(n22410), .CK(clk), .Q(\mem[462][0] ) );
  DFF_X1 \mem_reg[461][7]  ( .D(n22411), .CK(clk), .Q(\mem[461][7] ) );
  DFF_X1 \mem_reg[461][6]  ( .D(n22412), .CK(clk), .Q(\mem[461][6] ) );
  DFF_X1 \mem_reg[461][5]  ( .D(n22413), .CK(clk), .Q(\mem[461][5] ) );
  DFF_X1 \mem_reg[461][4]  ( .D(n22414), .CK(clk), .Q(\mem[461][4] ) );
  DFF_X1 \mem_reg[461][3]  ( .D(n22415), .CK(clk), .Q(\mem[461][3] ) );
  DFF_X1 \mem_reg[461][2]  ( .D(n22416), .CK(clk), .Q(\mem[461][2] ) );
  DFF_X1 \mem_reg[461][1]  ( .D(n22417), .CK(clk), .Q(\mem[461][1] ) );
  DFF_X1 \mem_reg[461][0]  ( .D(n22418), .CK(clk), .Q(\mem[461][0] ) );
  DFF_X1 \mem_reg[460][7]  ( .D(n22419), .CK(clk), .Q(\mem[460][7] ) );
  DFF_X1 \mem_reg[460][6]  ( .D(n22420), .CK(clk), .Q(\mem[460][6] ) );
  DFF_X1 \mem_reg[460][5]  ( .D(n22421), .CK(clk), .Q(\mem[460][5] ) );
  DFF_X1 \mem_reg[460][4]  ( .D(n22422), .CK(clk), .Q(\mem[460][4] ) );
  DFF_X1 \mem_reg[460][3]  ( .D(n22423), .CK(clk), .Q(\mem[460][3] ) );
  DFF_X1 \mem_reg[460][2]  ( .D(n22424), .CK(clk), .Q(\mem[460][2] ) );
  DFF_X1 \mem_reg[460][1]  ( .D(n22425), .CK(clk), .Q(\mem[460][1] ) );
  DFF_X1 \mem_reg[460][0]  ( .D(n22426), .CK(clk), .Q(\mem[460][0] ) );
  DFF_X1 \mem_reg[459][7]  ( .D(n22427), .CK(clk), .Q(\mem[459][7] ) );
  DFF_X1 \mem_reg[459][6]  ( .D(n22428), .CK(clk), .Q(\mem[459][6] ) );
  DFF_X1 \mem_reg[459][5]  ( .D(n22429), .CK(clk), .Q(\mem[459][5] ) );
  DFF_X1 \mem_reg[459][4]  ( .D(n22430), .CK(clk), .Q(\mem[459][4] ) );
  DFF_X1 \mem_reg[459][3]  ( .D(n22431), .CK(clk), .Q(\mem[459][3] ) );
  DFF_X1 \mem_reg[459][2]  ( .D(n22432), .CK(clk), .Q(\mem[459][2] ) );
  DFF_X1 \mem_reg[459][1]  ( .D(n22433), .CK(clk), .Q(\mem[459][1] ) );
  DFF_X1 \mem_reg[459][0]  ( .D(n22434), .CK(clk), .Q(\mem[459][0] ) );
  DFF_X1 \mem_reg[458][7]  ( .D(n22435), .CK(clk), .Q(\mem[458][7] ) );
  DFF_X1 \mem_reg[458][6]  ( .D(n22436), .CK(clk), .Q(\mem[458][6] ) );
  DFF_X1 \mem_reg[458][5]  ( .D(n22437), .CK(clk), .Q(\mem[458][5] ) );
  DFF_X1 \mem_reg[458][4]  ( .D(n22438), .CK(clk), .Q(\mem[458][4] ) );
  DFF_X1 \mem_reg[458][3]  ( .D(n22439), .CK(clk), .Q(\mem[458][3] ) );
  DFF_X1 \mem_reg[458][2]  ( .D(n22440), .CK(clk), .Q(\mem[458][2] ) );
  DFF_X1 \mem_reg[458][1]  ( .D(n22441), .CK(clk), .Q(\mem[458][1] ) );
  DFF_X1 \mem_reg[458][0]  ( .D(n22442), .CK(clk), .Q(\mem[458][0] ) );
  DFF_X1 \mem_reg[457][7]  ( .D(n22443), .CK(clk), .Q(\mem[457][7] ) );
  DFF_X1 \mem_reg[457][6]  ( .D(n22444), .CK(clk), .Q(\mem[457][6] ) );
  DFF_X1 \mem_reg[457][5]  ( .D(n22445), .CK(clk), .Q(\mem[457][5] ) );
  DFF_X1 \mem_reg[457][4]  ( .D(n22446), .CK(clk), .Q(\mem[457][4] ) );
  DFF_X1 \mem_reg[457][3]  ( .D(n22447), .CK(clk), .Q(\mem[457][3] ) );
  DFF_X1 \mem_reg[457][2]  ( .D(n22448), .CK(clk), .Q(\mem[457][2] ) );
  DFF_X1 \mem_reg[457][1]  ( .D(n22449), .CK(clk), .Q(\mem[457][1] ) );
  DFF_X1 \mem_reg[457][0]  ( .D(n22450), .CK(clk), .Q(\mem[457][0] ) );
  DFF_X1 \mem_reg[456][7]  ( .D(n22451), .CK(clk), .Q(\mem[456][7] ) );
  DFF_X1 \mem_reg[456][6]  ( .D(n22452), .CK(clk), .Q(\mem[456][6] ) );
  DFF_X1 \mem_reg[456][5]  ( .D(n22453), .CK(clk), .Q(\mem[456][5] ) );
  DFF_X1 \mem_reg[456][4]  ( .D(n22454), .CK(clk), .Q(\mem[456][4] ) );
  DFF_X1 \mem_reg[456][3]  ( .D(n22455), .CK(clk), .Q(\mem[456][3] ) );
  DFF_X1 \mem_reg[456][2]  ( .D(n22456), .CK(clk), .Q(\mem[456][2] ) );
  DFF_X1 \mem_reg[456][1]  ( .D(n22457), .CK(clk), .Q(\mem[456][1] ) );
  DFF_X1 \mem_reg[456][0]  ( .D(n22458), .CK(clk), .Q(\mem[456][0] ) );
  DFF_X1 \mem_reg[455][7]  ( .D(n22459), .CK(clk), .Q(\mem[455][7] ) );
  DFF_X1 \mem_reg[455][6]  ( .D(n22460), .CK(clk), .Q(\mem[455][6] ) );
  DFF_X1 \mem_reg[455][5]  ( .D(n22461), .CK(clk), .Q(\mem[455][5] ) );
  DFF_X1 \mem_reg[455][4]  ( .D(n22462), .CK(clk), .Q(\mem[455][4] ) );
  DFF_X1 \mem_reg[455][3]  ( .D(n22463), .CK(clk), .Q(\mem[455][3] ) );
  DFF_X1 \mem_reg[455][2]  ( .D(n22464), .CK(clk), .Q(\mem[455][2] ) );
  DFF_X1 \mem_reg[455][1]  ( .D(n22465), .CK(clk), .Q(\mem[455][1] ) );
  DFF_X1 \mem_reg[455][0]  ( .D(n22466), .CK(clk), .Q(\mem[455][0] ) );
  DFF_X1 \mem_reg[454][7]  ( .D(n22467), .CK(clk), .Q(\mem[454][7] ) );
  DFF_X1 \mem_reg[454][6]  ( .D(n22468), .CK(clk), .Q(\mem[454][6] ) );
  DFF_X1 \mem_reg[454][5]  ( .D(n22469), .CK(clk), .Q(\mem[454][5] ) );
  DFF_X1 \mem_reg[454][4]  ( .D(n22470), .CK(clk), .Q(\mem[454][4] ) );
  DFF_X1 \mem_reg[454][3]  ( .D(n22471), .CK(clk), .Q(\mem[454][3] ) );
  DFF_X1 \mem_reg[454][2]  ( .D(n22472), .CK(clk), .Q(\mem[454][2] ) );
  DFF_X1 \mem_reg[454][1]  ( .D(n22473), .CK(clk), .Q(\mem[454][1] ) );
  DFF_X1 \mem_reg[454][0]  ( .D(n22474), .CK(clk), .Q(\mem[454][0] ) );
  DFF_X1 \mem_reg[453][7]  ( .D(n22475), .CK(clk), .Q(\mem[453][7] ) );
  DFF_X1 \mem_reg[453][6]  ( .D(n22476), .CK(clk), .Q(\mem[453][6] ) );
  DFF_X1 \mem_reg[453][5]  ( .D(n22477), .CK(clk), .Q(\mem[453][5] ) );
  DFF_X1 \mem_reg[453][4]  ( .D(n22478), .CK(clk), .Q(\mem[453][4] ) );
  DFF_X1 \mem_reg[453][3]  ( .D(n22479), .CK(clk), .Q(\mem[453][3] ) );
  DFF_X1 \mem_reg[453][2]  ( .D(n22480), .CK(clk), .Q(\mem[453][2] ) );
  DFF_X1 \mem_reg[453][1]  ( .D(n22481), .CK(clk), .Q(\mem[453][1] ) );
  DFF_X1 \mem_reg[453][0]  ( .D(n22482), .CK(clk), .Q(\mem[453][0] ) );
  DFF_X1 \mem_reg[452][7]  ( .D(n22483), .CK(clk), .Q(\mem[452][7] ) );
  DFF_X1 \mem_reg[452][6]  ( .D(n22484), .CK(clk), .Q(\mem[452][6] ) );
  DFF_X1 \mem_reg[452][5]  ( .D(n22485), .CK(clk), .Q(\mem[452][5] ) );
  DFF_X1 \mem_reg[452][4]  ( .D(n22486), .CK(clk), .Q(\mem[452][4] ) );
  DFF_X1 \mem_reg[452][3]  ( .D(n22487), .CK(clk), .Q(\mem[452][3] ) );
  DFF_X1 \mem_reg[452][2]  ( .D(n22488), .CK(clk), .Q(\mem[452][2] ) );
  DFF_X1 \mem_reg[452][1]  ( .D(n22489), .CK(clk), .Q(\mem[452][1] ) );
  DFF_X1 \mem_reg[452][0]  ( .D(n22490), .CK(clk), .Q(\mem[452][0] ) );
  DFF_X1 \mem_reg[451][7]  ( .D(n22491), .CK(clk), .Q(\mem[451][7] ) );
  DFF_X1 \mem_reg[451][6]  ( .D(n22492), .CK(clk), .Q(\mem[451][6] ) );
  DFF_X1 \mem_reg[451][5]  ( .D(n22493), .CK(clk), .Q(\mem[451][5] ) );
  DFF_X1 \mem_reg[451][4]  ( .D(n22494), .CK(clk), .Q(\mem[451][4] ) );
  DFF_X1 \mem_reg[451][3]  ( .D(n22495), .CK(clk), .Q(\mem[451][3] ) );
  DFF_X1 \mem_reg[451][2]  ( .D(n22496), .CK(clk), .Q(\mem[451][2] ) );
  DFF_X1 \mem_reg[451][1]  ( .D(n22497), .CK(clk), .Q(\mem[451][1] ) );
  DFF_X1 \mem_reg[451][0]  ( .D(n22498), .CK(clk), .Q(\mem[451][0] ) );
  DFF_X1 \mem_reg[450][7]  ( .D(n22499), .CK(clk), .Q(\mem[450][7] ) );
  DFF_X1 \mem_reg[450][6]  ( .D(n22500), .CK(clk), .Q(\mem[450][6] ) );
  DFF_X1 \mem_reg[450][5]  ( .D(n22501), .CK(clk), .Q(\mem[450][5] ) );
  DFF_X1 \mem_reg[450][4]  ( .D(n22502), .CK(clk), .Q(\mem[450][4] ) );
  DFF_X1 \mem_reg[450][3]  ( .D(n22503), .CK(clk), .Q(\mem[450][3] ) );
  DFF_X1 \mem_reg[450][2]  ( .D(n22504), .CK(clk), .Q(\mem[450][2] ) );
  DFF_X1 \mem_reg[450][1]  ( .D(n22505), .CK(clk), .Q(\mem[450][1] ) );
  DFF_X1 \mem_reg[450][0]  ( .D(n22506), .CK(clk), .Q(\mem[450][0] ) );
  DFF_X1 \mem_reg[449][7]  ( .D(n22507), .CK(clk), .Q(\mem[449][7] ) );
  DFF_X1 \mem_reg[449][6]  ( .D(n22508), .CK(clk), .Q(\mem[449][6] ) );
  DFF_X1 \mem_reg[449][5]  ( .D(n22509), .CK(clk), .Q(\mem[449][5] ) );
  DFF_X1 \mem_reg[449][4]  ( .D(n22510), .CK(clk), .Q(\mem[449][4] ) );
  DFF_X1 \mem_reg[449][3]  ( .D(n22511), .CK(clk), .Q(\mem[449][3] ) );
  DFF_X1 \mem_reg[449][2]  ( .D(n22512), .CK(clk), .Q(\mem[449][2] ) );
  DFF_X1 \mem_reg[449][1]  ( .D(n22513), .CK(clk), .Q(\mem[449][1] ) );
  DFF_X1 \mem_reg[449][0]  ( .D(n22514), .CK(clk), .Q(\mem[449][0] ) );
  DFF_X1 \mem_reg[448][7]  ( .D(n22515), .CK(clk), .Q(\mem[448][7] ) );
  DFF_X1 \mem_reg[448][6]  ( .D(n22516), .CK(clk), .Q(\mem[448][6] ) );
  DFF_X1 \mem_reg[448][5]  ( .D(n22517), .CK(clk), .Q(\mem[448][5] ) );
  DFF_X1 \mem_reg[448][4]  ( .D(n22518), .CK(clk), .Q(\mem[448][4] ) );
  DFF_X1 \mem_reg[448][3]  ( .D(n22519), .CK(clk), .Q(\mem[448][3] ) );
  DFF_X1 \mem_reg[448][2]  ( .D(n22520), .CK(clk), .Q(\mem[448][2] ) );
  DFF_X1 \mem_reg[448][1]  ( .D(n22521), .CK(clk), .Q(\mem[448][1] ) );
  DFF_X1 \mem_reg[448][0]  ( .D(n22522), .CK(clk), .Q(\mem[448][0] ) );
  DFF_X1 \mem_reg[447][7]  ( .D(n22523), .CK(clk), .Q(\mem[447][7] ) );
  DFF_X1 \mem_reg[447][6]  ( .D(n22524), .CK(clk), .Q(\mem[447][6] ) );
  DFF_X1 \mem_reg[447][5]  ( .D(n22525), .CK(clk), .Q(\mem[447][5] ) );
  DFF_X1 \mem_reg[447][4]  ( .D(n22526), .CK(clk), .Q(\mem[447][4] ) );
  DFF_X1 \mem_reg[447][3]  ( .D(n22527), .CK(clk), .Q(\mem[447][3] ) );
  DFF_X1 \mem_reg[447][2]  ( .D(n22528), .CK(clk), .Q(\mem[447][2] ) );
  DFF_X1 \mem_reg[447][1]  ( .D(n22529), .CK(clk), .Q(\mem[447][1] ) );
  DFF_X1 \mem_reg[447][0]  ( .D(n22530), .CK(clk), .Q(\mem[447][0] ) );
  DFF_X1 \mem_reg[446][7]  ( .D(n22531), .CK(clk), .Q(\mem[446][7] ) );
  DFF_X1 \mem_reg[446][6]  ( .D(n22532), .CK(clk), .Q(\mem[446][6] ) );
  DFF_X1 \mem_reg[446][5]  ( .D(n22533), .CK(clk), .Q(\mem[446][5] ) );
  DFF_X1 \mem_reg[446][4]  ( .D(n22534), .CK(clk), .Q(\mem[446][4] ) );
  DFF_X1 \mem_reg[446][3]  ( .D(n22535), .CK(clk), .Q(\mem[446][3] ) );
  DFF_X1 \mem_reg[446][2]  ( .D(n22536), .CK(clk), .Q(\mem[446][2] ) );
  DFF_X1 \mem_reg[446][1]  ( .D(n22537), .CK(clk), .Q(\mem[446][1] ) );
  DFF_X1 \mem_reg[446][0]  ( .D(n22538), .CK(clk), .Q(\mem[446][0] ) );
  DFF_X1 \mem_reg[445][7]  ( .D(n22539), .CK(clk), .Q(\mem[445][7] ) );
  DFF_X1 \mem_reg[445][6]  ( .D(n22540), .CK(clk), .Q(\mem[445][6] ) );
  DFF_X1 \mem_reg[445][5]  ( .D(n22541), .CK(clk), .Q(\mem[445][5] ) );
  DFF_X1 \mem_reg[445][4]  ( .D(n22542), .CK(clk), .Q(\mem[445][4] ) );
  DFF_X1 \mem_reg[445][3]  ( .D(n22543), .CK(clk), .Q(\mem[445][3] ) );
  DFF_X1 \mem_reg[445][2]  ( .D(n22544), .CK(clk), .Q(\mem[445][2] ) );
  DFF_X1 \mem_reg[445][1]  ( .D(n22545), .CK(clk), .Q(\mem[445][1] ) );
  DFF_X1 \mem_reg[445][0]  ( .D(n22546), .CK(clk), .Q(\mem[445][0] ) );
  DFF_X1 \mem_reg[444][7]  ( .D(n22547), .CK(clk), .Q(\mem[444][7] ) );
  DFF_X1 \mem_reg[444][6]  ( .D(n22548), .CK(clk), .Q(\mem[444][6] ) );
  DFF_X1 \mem_reg[444][5]  ( .D(n22549), .CK(clk), .Q(\mem[444][5] ) );
  DFF_X1 \mem_reg[444][4]  ( .D(n22550), .CK(clk), .Q(\mem[444][4] ) );
  DFF_X1 \mem_reg[444][3]  ( .D(n22551), .CK(clk), .Q(\mem[444][3] ) );
  DFF_X1 \mem_reg[444][2]  ( .D(n22552), .CK(clk), .Q(\mem[444][2] ) );
  DFF_X1 \mem_reg[444][1]  ( .D(n22553), .CK(clk), .Q(\mem[444][1] ) );
  DFF_X1 \mem_reg[444][0]  ( .D(n22554), .CK(clk), .Q(\mem[444][0] ) );
  DFF_X1 \mem_reg[443][7]  ( .D(n22555), .CK(clk), .Q(\mem[443][7] ) );
  DFF_X1 \mem_reg[443][6]  ( .D(n22556), .CK(clk), .Q(\mem[443][6] ) );
  DFF_X1 \mem_reg[443][5]  ( .D(n22557), .CK(clk), .Q(\mem[443][5] ) );
  DFF_X1 \mem_reg[443][4]  ( .D(n22558), .CK(clk), .Q(\mem[443][4] ) );
  DFF_X1 \mem_reg[443][3]  ( .D(n22559), .CK(clk), .Q(\mem[443][3] ) );
  DFF_X1 \mem_reg[443][2]  ( .D(n22560), .CK(clk), .Q(\mem[443][2] ) );
  DFF_X1 \mem_reg[443][1]  ( .D(n22561), .CK(clk), .Q(\mem[443][1] ) );
  DFF_X1 \mem_reg[443][0]  ( .D(n22562), .CK(clk), .Q(\mem[443][0] ) );
  DFF_X1 \mem_reg[442][7]  ( .D(n22563), .CK(clk), .Q(\mem[442][7] ) );
  DFF_X1 \mem_reg[442][6]  ( .D(n22564), .CK(clk), .Q(\mem[442][6] ) );
  DFF_X1 \mem_reg[442][5]  ( .D(n22565), .CK(clk), .Q(\mem[442][5] ) );
  DFF_X1 \mem_reg[442][4]  ( .D(n22566), .CK(clk), .Q(\mem[442][4] ) );
  DFF_X1 \mem_reg[442][3]  ( .D(n22567), .CK(clk), .Q(\mem[442][3] ) );
  DFF_X1 \mem_reg[442][2]  ( .D(n22568), .CK(clk), .Q(\mem[442][2] ) );
  DFF_X1 \mem_reg[442][1]  ( .D(n22569), .CK(clk), .Q(\mem[442][1] ) );
  DFF_X1 \mem_reg[442][0]  ( .D(n22570), .CK(clk), .Q(\mem[442][0] ) );
  DFF_X1 \mem_reg[441][7]  ( .D(n22571), .CK(clk), .Q(\mem[441][7] ) );
  DFF_X1 \mem_reg[441][6]  ( .D(n22572), .CK(clk), .Q(\mem[441][6] ) );
  DFF_X1 \mem_reg[441][5]  ( .D(n22573), .CK(clk), .Q(\mem[441][5] ) );
  DFF_X1 \mem_reg[441][4]  ( .D(n22574), .CK(clk), .Q(\mem[441][4] ) );
  DFF_X1 \mem_reg[441][3]  ( .D(n22575), .CK(clk), .Q(\mem[441][3] ) );
  DFF_X1 \mem_reg[441][2]  ( .D(n22576), .CK(clk), .Q(\mem[441][2] ) );
  DFF_X1 \mem_reg[441][1]  ( .D(n22577), .CK(clk), .Q(\mem[441][1] ) );
  DFF_X1 \mem_reg[441][0]  ( .D(n22578), .CK(clk), .Q(\mem[441][0] ) );
  DFF_X1 \mem_reg[440][7]  ( .D(n22579), .CK(clk), .Q(\mem[440][7] ) );
  DFF_X1 \mem_reg[440][6]  ( .D(n22580), .CK(clk), .Q(\mem[440][6] ) );
  DFF_X1 \mem_reg[440][5]  ( .D(n22581), .CK(clk), .Q(\mem[440][5] ) );
  DFF_X1 \mem_reg[440][4]  ( .D(n22582), .CK(clk), .Q(\mem[440][4] ) );
  DFF_X1 \mem_reg[440][3]  ( .D(n22583), .CK(clk), .Q(\mem[440][3] ) );
  DFF_X1 \mem_reg[440][2]  ( .D(n22584), .CK(clk), .Q(\mem[440][2] ) );
  DFF_X1 \mem_reg[440][1]  ( .D(n22585), .CK(clk), .Q(\mem[440][1] ) );
  DFF_X1 \mem_reg[440][0]  ( .D(n22586), .CK(clk), .Q(\mem[440][0] ) );
  DFF_X1 \mem_reg[439][7]  ( .D(n22587), .CK(clk), .Q(\mem[439][7] ) );
  DFF_X1 \mem_reg[439][6]  ( .D(n22588), .CK(clk), .Q(\mem[439][6] ) );
  DFF_X1 \mem_reg[439][5]  ( .D(n22589), .CK(clk), .Q(\mem[439][5] ) );
  DFF_X1 \mem_reg[439][4]  ( .D(n22590), .CK(clk), .Q(\mem[439][4] ) );
  DFF_X1 \mem_reg[439][3]  ( .D(n22591), .CK(clk), .Q(\mem[439][3] ) );
  DFF_X1 \mem_reg[439][2]  ( .D(n22592), .CK(clk), .Q(\mem[439][2] ) );
  DFF_X1 \mem_reg[439][1]  ( .D(n22593), .CK(clk), .Q(\mem[439][1] ) );
  DFF_X1 \mem_reg[439][0]  ( .D(n22594), .CK(clk), .Q(\mem[439][0] ) );
  DFF_X1 \mem_reg[438][7]  ( .D(n22595), .CK(clk), .Q(\mem[438][7] ) );
  DFF_X1 \mem_reg[438][6]  ( .D(n22596), .CK(clk), .Q(\mem[438][6] ) );
  DFF_X1 \mem_reg[438][5]  ( .D(n22597), .CK(clk), .Q(\mem[438][5] ) );
  DFF_X1 \mem_reg[438][4]  ( .D(n22598), .CK(clk), .Q(\mem[438][4] ) );
  DFF_X1 \mem_reg[438][3]  ( .D(n22599), .CK(clk), .Q(\mem[438][3] ) );
  DFF_X1 \mem_reg[438][2]  ( .D(n22600), .CK(clk), .Q(\mem[438][2] ) );
  DFF_X1 \mem_reg[438][1]  ( .D(n22601), .CK(clk), .Q(\mem[438][1] ) );
  DFF_X1 \mem_reg[438][0]  ( .D(n22602), .CK(clk), .Q(\mem[438][0] ) );
  DFF_X1 \mem_reg[437][7]  ( .D(n22603), .CK(clk), .Q(\mem[437][7] ) );
  DFF_X1 \mem_reg[437][6]  ( .D(n22604), .CK(clk), .Q(\mem[437][6] ) );
  DFF_X1 \mem_reg[437][5]  ( .D(n22605), .CK(clk), .Q(\mem[437][5] ) );
  DFF_X1 \mem_reg[437][4]  ( .D(n22606), .CK(clk), .Q(\mem[437][4] ) );
  DFF_X1 \mem_reg[437][3]  ( .D(n22607), .CK(clk), .Q(\mem[437][3] ) );
  DFF_X1 \mem_reg[437][2]  ( .D(n22608), .CK(clk), .Q(\mem[437][2] ) );
  DFF_X1 \mem_reg[437][1]  ( .D(n22609), .CK(clk), .Q(\mem[437][1] ) );
  DFF_X1 \mem_reg[437][0]  ( .D(n22610), .CK(clk), .Q(\mem[437][0] ) );
  DFF_X1 \mem_reg[436][7]  ( .D(n22611), .CK(clk), .Q(\mem[436][7] ) );
  DFF_X1 \mem_reg[436][6]  ( .D(n22612), .CK(clk), .Q(\mem[436][6] ) );
  DFF_X1 \mem_reg[436][5]  ( .D(n22613), .CK(clk), .Q(\mem[436][5] ) );
  DFF_X1 \mem_reg[436][4]  ( .D(n22614), .CK(clk), .Q(\mem[436][4] ) );
  DFF_X1 \mem_reg[436][3]  ( .D(n22615), .CK(clk), .Q(\mem[436][3] ) );
  DFF_X1 \mem_reg[436][2]  ( .D(n22616), .CK(clk), .Q(\mem[436][2] ) );
  DFF_X1 \mem_reg[436][1]  ( .D(n22617), .CK(clk), .Q(\mem[436][1] ) );
  DFF_X1 \mem_reg[436][0]  ( .D(n22618), .CK(clk), .Q(\mem[436][0] ) );
  DFF_X1 \mem_reg[435][7]  ( .D(n22619), .CK(clk), .Q(\mem[435][7] ) );
  DFF_X1 \mem_reg[435][6]  ( .D(n22620), .CK(clk), .Q(\mem[435][6] ) );
  DFF_X1 \mem_reg[435][5]  ( .D(n22621), .CK(clk), .Q(\mem[435][5] ) );
  DFF_X1 \mem_reg[435][4]  ( .D(n22622), .CK(clk), .Q(\mem[435][4] ) );
  DFF_X1 \mem_reg[435][3]  ( .D(n22623), .CK(clk), .Q(\mem[435][3] ) );
  DFF_X1 \mem_reg[435][2]  ( .D(n22624), .CK(clk), .Q(\mem[435][2] ) );
  DFF_X1 \mem_reg[435][1]  ( .D(n22625), .CK(clk), .Q(\mem[435][1] ) );
  DFF_X1 \mem_reg[435][0]  ( .D(n22626), .CK(clk), .Q(\mem[435][0] ) );
  DFF_X1 \mem_reg[434][7]  ( .D(n22627), .CK(clk), .Q(\mem[434][7] ) );
  DFF_X1 \mem_reg[434][6]  ( .D(n22628), .CK(clk), .Q(\mem[434][6] ) );
  DFF_X1 \mem_reg[434][5]  ( .D(n22629), .CK(clk), .Q(\mem[434][5] ) );
  DFF_X1 \mem_reg[434][4]  ( .D(n22630), .CK(clk), .Q(\mem[434][4] ) );
  DFF_X1 \mem_reg[434][3]  ( .D(n22631), .CK(clk), .Q(\mem[434][3] ) );
  DFF_X1 \mem_reg[434][2]  ( .D(n22632), .CK(clk), .Q(\mem[434][2] ) );
  DFF_X1 \mem_reg[434][1]  ( .D(n22633), .CK(clk), .Q(\mem[434][1] ) );
  DFF_X1 \mem_reg[434][0]  ( .D(n22634), .CK(clk), .Q(\mem[434][0] ) );
  DFF_X1 \mem_reg[433][7]  ( .D(n22635), .CK(clk), .Q(\mem[433][7] ) );
  DFF_X1 \mem_reg[433][6]  ( .D(n22636), .CK(clk), .Q(\mem[433][6] ) );
  DFF_X1 \mem_reg[433][5]  ( .D(n22637), .CK(clk), .Q(\mem[433][5] ) );
  DFF_X1 \mem_reg[433][4]  ( .D(n22638), .CK(clk), .Q(\mem[433][4] ) );
  DFF_X1 \mem_reg[433][3]  ( .D(n22639), .CK(clk), .Q(\mem[433][3] ) );
  DFF_X1 \mem_reg[433][2]  ( .D(n22640), .CK(clk), .Q(\mem[433][2] ) );
  DFF_X1 \mem_reg[433][1]  ( .D(n22641), .CK(clk), .Q(\mem[433][1] ) );
  DFF_X1 \mem_reg[433][0]  ( .D(n22642), .CK(clk), .Q(\mem[433][0] ) );
  DFF_X1 \mem_reg[432][7]  ( .D(n22643), .CK(clk), .Q(\mem[432][7] ) );
  DFF_X1 \mem_reg[432][6]  ( .D(n22644), .CK(clk), .Q(\mem[432][6] ) );
  DFF_X1 \mem_reg[432][5]  ( .D(n22645), .CK(clk), .Q(\mem[432][5] ) );
  DFF_X1 \mem_reg[432][4]  ( .D(n22646), .CK(clk), .Q(\mem[432][4] ) );
  DFF_X1 \mem_reg[432][3]  ( .D(n22647), .CK(clk), .Q(\mem[432][3] ) );
  DFF_X1 \mem_reg[432][2]  ( .D(n22648), .CK(clk), .Q(\mem[432][2] ) );
  DFF_X1 \mem_reg[432][1]  ( .D(n22649), .CK(clk), .Q(\mem[432][1] ) );
  DFF_X1 \mem_reg[432][0]  ( .D(n22650), .CK(clk), .Q(\mem[432][0] ) );
  DFF_X1 \mem_reg[431][7]  ( .D(n22651), .CK(clk), .Q(\mem[431][7] ) );
  DFF_X1 \mem_reg[431][6]  ( .D(n22652), .CK(clk), .Q(\mem[431][6] ) );
  DFF_X1 \mem_reg[431][5]  ( .D(n22653), .CK(clk), .Q(\mem[431][5] ) );
  DFF_X1 \mem_reg[431][4]  ( .D(n22654), .CK(clk), .Q(\mem[431][4] ) );
  DFF_X1 \mem_reg[431][3]  ( .D(n22655), .CK(clk), .Q(\mem[431][3] ) );
  DFF_X1 \mem_reg[431][2]  ( .D(n22656), .CK(clk), .Q(\mem[431][2] ) );
  DFF_X1 \mem_reg[431][1]  ( .D(n22657), .CK(clk), .Q(\mem[431][1] ) );
  DFF_X1 \mem_reg[431][0]  ( .D(n22658), .CK(clk), .Q(\mem[431][0] ) );
  DFF_X1 \mem_reg[430][7]  ( .D(n22659), .CK(clk), .Q(\mem[430][7] ) );
  DFF_X1 \mem_reg[430][6]  ( .D(n22660), .CK(clk), .Q(\mem[430][6] ) );
  DFF_X1 \mem_reg[430][5]  ( .D(n22661), .CK(clk), .Q(\mem[430][5] ) );
  DFF_X1 \mem_reg[430][4]  ( .D(n22662), .CK(clk), .Q(\mem[430][4] ) );
  DFF_X1 \mem_reg[430][3]  ( .D(n22663), .CK(clk), .Q(\mem[430][3] ) );
  DFF_X1 \mem_reg[430][2]  ( .D(n22664), .CK(clk), .Q(\mem[430][2] ) );
  DFF_X1 \mem_reg[430][1]  ( .D(n22665), .CK(clk), .Q(\mem[430][1] ) );
  DFF_X1 \mem_reg[430][0]  ( .D(n22666), .CK(clk), .Q(\mem[430][0] ) );
  DFF_X1 \mem_reg[429][7]  ( .D(n22667), .CK(clk), .Q(\mem[429][7] ) );
  DFF_X1 \mem_reg[429][6]  ( .D(n22668), .CK(clk), .Q(\mem[429][6] ) );
  DFF_X1 \mem_reg[429][5]  ( .D(n22669), .CK(clk), .Q(\mem[429][5] ) );
  DFF_X1 \mem_reg[429][4]  ( .D(n22670), .CK(clk), .Q(\mem[429][4] ) );
  DFF_X1 \mem_reg[429][3]  ( .D(n22671), .CK(clk), .Q(\mem[429][3] ) );
  DFF_X1 \mem_reg[429][2]  ( .D(n22672), .CK(clk), .Q(\mem[429][2] ) );
  DFF_X1 \mem_reg[429][1]  ( .D(n22673), .CK(clk), .Q(\mem[429][1] ) );
  DFF_X1 \mem_reg[429][0]  ( .D(n22674), .CK(clk), .Q(\mem[429][0] ) );
  DFF_X1 \mem_reg[428][7]  ( .D(n22675), .CK(clk), .Q(\mem[428][7] ) );
  DFF_X1 \mem_reg[428][6]  ( .D(n22676), .CK(clk), .Q(\mem[428][6] ) );
  DFF_X1 \mem_reg[428][5]  ( .D(n22677), .CK(clk), .Q(\mem[428][5] ) );
  DFF_X1 \mem_reg[428][4]  ( .D(n22678), .CK(clk), .Q(\mem[428][4] ) );
  DFF_X1 \mem_reg[428][3]  ( .D(n22679), .CK(clk), .Q(\mem[428][3] ) );
  DFF_X1 \mem_reg[428][2]  ( .D(n22680), .CK(clk), .Q(\mem[428][2] ) );
  DFF_X1 \mem_reg[428][1]  ( .D(n22681), .CK(clk), .Q(\mem[428][1] ) );
  DFF_X1 \mem_reg[428][0]  ( .D(n22682), .CK(clk), .Q(\mem[428][0] ) );
  DFF_X1 \mem_reg[427][7]  ( .D(n22683), .CK(clk), .Q(\mem[427][7] ) );
  DFF_X1 \mem_reg[427][6]  ( .D(n22684), .CK(clk), .Q(\mem[427][6] ) );
  DFF_X1 \mem_reg[427][5]  ( .D(n22685), .CK(clk), .Q(\mem[427][5] ) );
  DFF_X1 \mem_reg[427][4]  ( .D(n22686), .CK(clk), .Q(\mem[427][4] ) );
  DFF_X1 \mem_reg[427][3]  ( .D(n22687), .CK(clk), .Q(\mem[427][3] ) );
  DFF_X1 \mem_reg[427][2]  ( .D(n22688), .CK(clk), .Q(\mem[427][2] ) );
  DFF_X1 \mem_reg[427][1]  ( .D(n22689), .CK(clk), .Q(\mem[427][1] ) );
  DFF_X1 \mem_reg[427][0]  ( .D(n22690), .CK(clk), .Q(\mem[427][0] ) );
  DFF_X1 \mem_reg[426][7]  ( .D(n22691), .CK(clk), .Q(\mem[426][7] ) );
  DFF_X1 \mem_reg[426][6]  ( .D(n22692), .CK(clk), .Q(\mem[426][6] ) );
  DFF_X1 \mem_reg[426][5]  ( .D(n22693), .CK(clk), .Q(\mem[426][5] ) );
  DFF_X1 \mem_reg[426][4]  ( .D(n22694), .CK(clk), .Q(\mem[426][4] ) );
  DFF_X1 \mem_reg[426][3]  ( .D(n22695), .CK(clk), .Q(\mem[426][3] ) );
  DFF_X1 \mem_reg[426][2]  ( .D(n22696), .CK(clk), .Q(\mem[426][2] ) );
  DFF_X1 \mem_reg[426][1]  ( .D(n22697), .CK(clk), .Q(\mem[426][1] ) );
  DFF_X1 \mem_reg[426][0]  ( .D(n22698), .CK(clk), .Q(\mem[426][0] ) );
  DFF_X1 \mem_reg[425][7]  ( .D(n22699), .CK(clk), .Q(\mem[425][7] ) );
  DFF_X1 \mem_reg[425][6]  ( .D(n22700), .CK(clk), .Q(\mem[425][6] ) );
  DFF_X1 \mem_reg[425][5]  ( .D(n22701), .CK(clk), .Q(\mem[425][5] ) );
  DFF_X1 \mem_reg[425][4]  ( .D(n22702), .CK(clk), .Q(\mem[425][4] ) );
  DFF_X1 \mem_reg[425][3]  ( .D(n22703), .CK(clk), .Q(\mem[425][3] ) );
  DFF_X1 \mem_reg[425][2]  ( .D(n22704), .CK(clk), .Q(\mem[425][2] ) );
  DFF_X1 \mem_reg[425][1]  ( .D(n22705), .CK(clk), .Q(\mem[425][1] ) );
  DFF_X1 \mem_reg[425][0]  ( .D(n22706), .CK(clk), .Q(\mem[425][0] ) );
  DFF_X1 \mem_reg[424][7]  ( .D(n22707), .CK(clk), .Q(\mem[424][7] ) );
  DFF_X1 \mem_reg[424][6]  ( .D(n22708), .CK(clk), .Q(\mem[424][6] ) );
  DFF_X1 \mem_reg[424][5]  ( .D(n22709), .CK(clk), .Q(\mem[424][5] ) );
  DFF_X1 \mem_reg[424][4]  ( .D(n22710), .CK(clk), .Q(\mem[424][4] ) );
  DFF_X1 \mem_reg[424][3]  ( .D(n22711), .CK(clk), .Q(\mem[424][3] ) );
  DFF_X1 \mem_reg[424][2]  ( .D(n22712), .CK(clk), .Q(\mem[424][2] ) );
  DFF_X1 \mem_reg[424][1]  ( .D(n22713), .CK(clk), .Q(\mem[424][1] ) );
  DFF_X1 \mem_reg[424][0]  ( .D(n22714), .CK(clk), .Q(\mem[424][0] ) );
  DFF_X1 \mem_reg[423][7]  ( .D(n22715), .CK(clk), .Q(\mem[423][7] ) );
  DFF_X1 \mem_reg[423][6]  ( .D(n22716), .CK(clk), .Q(\mem[423][6] ) );
  DFF_X1 \mem_reg[423][5]  ( .D(n22717), .CK(clk), .Q(\mem[423][5] ) );
  DFF_X1 \mem_reg[423][4]  ( .D(n22718), .CK(clk), .Q(\mem[423][4] ) );
  DFF_X1 \mem_reg[423][3]  ( .D(n22719), .CK(clk), .Q(\mem[423][3] ) );
  DFF_X1 \mem_reg[423][2]  ( .D(n22720), .CK(clk), .Q(\mem[423][2] ) );
  DFF_X1 \mem_reg[423][1]  ( .D(n22721), .CK(clk), .Q(\mem[423][1] ) );
  DFF_X1 \mem_reg[423][0]  ( .D(n22722), .CK(clk), .Q(\mem[423][0] ) );
  DFF_X1 \mem_reg[422][7]  ( .D(n22723), .CK(clk), .Q(\mem[422][7] ) );
  DFF_X1 \mem_reg[422][6]  ( .D(n22724), .CK(clk), .Q(\mem[422][6] ) );
  DFF_X1 \mem_reg[422][5]  ( .D(n22725), .CK(clk), .Q(\mem[422][5] ) );
  DFF_X1 \mem_reg[422][4]  ( .D(n22726), .CK(clk), .Q(\mem[422][4] ) );
  DFF_X1 \mem_reg[422][3]  ( .D(n22727), .CK(clk), .Q(\mem[422][3] ) );
  DFF_X1 \mem_reg[422][2]  ( .D(n22728), .CK(clk), .Q(\mem[422][2] ) );
  DFF_X1 \mem_reg[422][1]  ( .D(n22729), .CK(clk), .Q(\mem[422][1] ) );
  DFF_X1 \mem_reg[422][0]  ( .D(n22730), .CK(clk), .Q(\mem[422][0] ) );
  DFF_X1 \mem_reg[421][7]  ( .D(n22731), .CK(clk), .Q(\mem[421][7] ) );
  DFF_X1 \mem_reg[421][6]  ( .D(n22732), .CK(clk), .Q(\mem[421][6] ) );
  DFF_X1 \mem_reg[421][5]  ( .D(n22733), .CK(clk), .Q(\mem[421][5] ) );
  DFF_X1 \mem_reg[421][4]  ( .D(n22734), .CK(clk), .Q(\mem[421][4] ) );
  DFF_X1 \mem_reg[421][3]  ( .D(n22735), .CK(clk), .Q(\mem[421][3] ) );
  DFF_X1 \mem_reg[421][2]  ( .D(n22736), .CK(clk), .Q(\mem[421][2] ) );
  DFF_X1 \mem_reg[421][1]  ( .D(n22737), .CK(clk), .Q(\mem[421][1] ) );
  DFF_X1 \mem_reg[421][0]  ( .D(n22738), .CK(clk), .Q(\mem[421][0] ) );
  DFF_X1 \mem_reg[420][7]  ( .D(n22739), .CK(clk), .Q(\mem[420][7] ) );
  DFF_X1 \mem_reg[420][6]  ( .D(n22740), .CK(clk), .Q(\mem[420][6] ) );
  DFF_X1 \mem_reg[420][5]  ( .D(n22741), .CK(clk), .Q(\mem[420][5] ) );
  DFF_X1 \mem_reg[420][4]  ( .D(n22742), .CK(clk), .Q(\mem[420][4] ) );
  DFF_X1 \mem_reg[420][3]  ( .D(n22743), .CK(clk), .Q(\mem[420][3] ) );
  DFF_X1 \mem_reg[420][2]  ( .D(n22744), .CK(clk), .Q(\mem[420][2] ) );
  DFF_X1 \mem_reg[420][1]  ( .D(n22745), .CK(clk), .Q(\mem[420][1] ) );
  DFF_X1 \mem_reg[420][0]  ( .D(n22746), .CK(clk), .Q(\mem[420][0] ) );
  DFF_X1 \mem_reg[419][7]  ( .D(n22747), .CK(clk), .Q(\mem[419][7] ) );
  DFF_X1 \mem_reg[419][6]  ( .D(n22748), .CK(clk), .Q(\mem[419][6] ) );
  DFF_X1 \mem_reg[419][5]  ( .D(n22749), .CK(clk), .Q(\mem[419][5] ) );
  DFF_X1 \mem_reg[419][4]  ( .D(n22750), .CK(clk), .Q(\mem[419][4] ) );
  DFF_X1 \mem_reg[419][3]  ( .D(n22751), .CK(clk), .Q(\mem[419][3] ) );
  DFF_X1 \mem_reg[419][2]  ( .D(n22752), .CK(clk), .Q(\mem[419][2] ) );
  DFF_X1 \mem_reg[419][1]  ( .D(n22753), .CK(clk), .Q(\mem[419][1] ) );
  DFF_X1 \mem_reg[419][0]  ( .D(n22754), .CK(clk), .Q(\mem[419][0] ) );
  DFF_X1 \mem_reg[418][7]  ( .D(n22755), .CK(clk), .Q(\mem[418][7] ) );
  DFF_X1 \mem_reg[418][6]  ( .D(n22756), .CK(clk), .Q(\mem[418][6] ) );
  DFF_X1 \mem_reg[418][5]  ( .D(n22757), .CK(clk), .Q(\mem[418][5] ) );
  DFF_X1 \mem_reg[418][4]  ( .D(n22758), .CK(clk), .Q(\mem[418][4] ) );
  DFF_X1 \mem_reg[418][3]  ( .D(n22759), .CK(clk), .Q(\mem[418][3] ) );
  DFF_X1 \mem_reg[418][2]  ( .D(n22760), .CK(clk), .Q(\mem[418][2] ) );
  DFF_X1 \mem_reg[418][1]  ( .D(n22761), .CK(clk), .Q(\mem[418][1] ) );
  DFF_X1 \mem_reg[418][0]  ( .D(n22762), .CK(clk), .Q(\mem[418][0] ) );
  DFF_X1 \mem_reg[417][7]  ( .D(n22763), .CK(clk), .Q(\mem[417][7] ) );
  DFF_X1 \mem_reg[417][6]  ( .D(n22764), .CK(clk), .Q(\mem[417][6] ) );
  DFF_X1 \mem_reg[417][5]  ( .D(n22765), .CK(clk), .Q(\mem[417][5] ) );
  DFF_X1 \mem_reg[417][4]  ( .D(n22766), .CK(clk), .Q(\mem[417][4] ) );
  DFF_X1 \mem_reg[417][3]  ( .D(n22767), .CK(clk), .Q(\mem[417][3] ) );
  DFF_X1 \mem_reg[417][2]  ( .D(n22768), .CK(clk), .Q(\mem[417][2] ) );
  DFF_X1 \mem_reg[417][1]  ( .D(n22769), .CK(clk), .Q(\mem[417][1] ) );
  DFF_X1 \mem_reg[417][0]  ( .D(n22770), .CK(clk), .Q(\mem[417][0] ) );
  DFF_X1 \mem_reg[416][7]  ( .D(n22771), .CK(clk), .Q(\mem[416][7] ) );
  DFF_X1 \mem_reg[416][6]  ( .D(n22772), .CK(clk), .Q(\mem[416][6] ) );
  DFF_X1 \mem_reg[416][5]  ( .D(n22773), .CK(clk), .Q(\mem[416][5] ) );
  DFF_X1 \mem_reg[416][4]  ( .D(n22774), .CK(clk), .Q(\mem[416][4] ) );
  DFF_X1 \mem_reg[416][3]  ( .D(n22775), .CK(clk), .Q(\mem[416][3] ) );
  DFF_X1 \mem_reg[416][2]  ( .D(n22776), .CK(clk), .Q(\mem[416][2] ) );
  DFF_X1 \mem_reg[416][1]  ( .D(n22777), .CK(clk), .Q(\mem[416][1] ) );
  DFF_X1 \mem_reg[416][0]  ( .D(n22778), .CK(clk), .Q(\mem[416][0] ) );
  DFF_X1 \mem_reg[415][7]  ( .D(n22779), .CK(clk), .Q(\mem[415][7] ) );
  DFF_X1 \mem_reg[415][6]  ( .D(n22780), .CK(clk), .Q(\mem[415][6] ) );
  DFF_X1 \mem_reg[415][5]  ( .D(n22781), .CK(clk), .Q(\mem[415][5] ) );
  DFF_X1 \mem_reg[415][4]  ( .D(n22782), .CK(clk), .Q(\mem[415][4] ) );
  DFF_X1 \mem_reg[415][3]  ( .D(n22783), .CK(clk), .Q(\mem[415][3] ) );
  DFF_X1 \mem_reg[415][2]  ( .D(n22784), .CK(clk), .Q(\mem[415][2] ) );
  DFF_X1 \mem_reg[415][1]  ( .D(n22785), .CK(clk), .Q(\mem[415][1] ) );
  DFF_X1 \mem_reg[415][0]  ( .D(n22786), .CK(clk), .Q(\mem[415][0] ) );
  DFF_X1 \mem_reg[414][7]  ( .D(n22787), .CK(clk), .Q(\mem[414][7] ) );
  DFF_X1 \mem_reg[414][6]  ( .D(n22788), .CK(clk), .Q(\mem[414][6] ) );
  DFF_X1 \mem_reg[414][5]  ( .D(n22789), .CK(clk), .Q(\mem[414][5] ) );
  DFF_X1 \mem_reg[414][4]  ( .D(n22790), .CK(clk), .Q(\mem[414][4] ) );
  DFF_X1 \mem_reg[414][3]  ( .D(n22791), .CK(clk), .Q(\mem[414][3] ) );
  DFF_X1 \mem_reg[414][2]  ( .D(n22792), .CK(clk), .Q(\mem[414][2] ) );
  DFF_X1 \mem_reg[414][1]  ( .D(n22793), .CK(clk), .Q(\mem[414][1] ) );
  DFF_X1 \mem_reg[414][0]  ( .D(n22794), .CK(clk), .Q(\mem[414][0] ) );
  DFF_X1 \mem_reg[413][7]  ( .D(n22795), .CK(clk), .Q(\mem[413][7] ) );
  DFF_X1 \mem_reg[413][6]  ( .D(n22796), .CK(clk), .Q(\mem[413][6] ) );
  DFF_X1 \mem_reg[413][5]  ( .D(n22797), .CK(clk), .Q(\mem[413][5] ) );
  DFF_X1 \mem_reg[413][4]  ( .D(n22798), .CK(clk), .Q(\mem[413][4] ) );
  DFF_X1 \mem_reg[413][3]  ( .D(n22799), .CK(clk), .Q(\mem[413][3] ) );
  DFF_X1 \mem_reg[413][2]  ( .D(n22800), .CK(clk), .Q(\mem[413][2] ) );
  DFF_X1 \mem_reg[413][1]  ( .D(n22801), .CK(clk), .Q(\mem[413][1] ) );
  DFF_X1 \mem_reg[413][0]  ( .D(n22802), .CK(clk), .Q(\mem[413][0] ) );
  DFF_X1 \mem_reg[412][7]  ( .D(n22803), .CK(clk), .Q(\mem[412][7] ) );
  DFF_X1 \mem_reg[412][6]  ( .D(n22804), .CK(clk), .Q(\mem[412][6] ) );
  DFF_X1 \mem_reg[412][5]  ( .D(n22805), .CK(clk), .Q(\mem[412][5] ) );
  DFF_X1 \mem_reg[412][4]  ( .D(n22806), .CK(clk), .Q(\mem[412][4] ) );
  DFF_X1 \mem_reg[412][3]  ( .D(n22807), .CK(clk), .Q(\mem[412][3] ) );
  DFF_X1 \mem_reg[412][2]  ( .D(n22808), .CK(clk), .Q(\mem[412][2] ) );
  DFF_X1 \mem_reg[412][1]  ( .D(n22809), .CK(clk), .Q(\mem[412][1] ) );
  DFF_X1 \mem_reg[412][0]  ( .D(n22810), .CK(clk), .Q(\mem[412][0] ) );
  DFF_X1 \mem_reg[411][7]  ( .D(n22811), .CK(clk), .Q(\mem[411][7] ) );
  DFF_X1 \mem_reg[411][6]  ( .D(n22812), .CK(clk), .Q(\mem[411][6] ) );
  DFF_X1 \mem_reg[411][5]  ( .D(n22813), .CK(clk), .Q(\mem[411][5] ) );
  DFF_X1 \mem_reg[411][4]  ( .D(n22814), .CK(clk), .Q(\mem[411][4] ) );
  DFF_X1 \mem_reg[411][3]  ( .D(n22815), .CK(clk), .Q(\mem[411][3] ) );
  DFF_X1 \mem_reg[411][2]  ( .D(n22816), .CK(clk), .Q(\mem[411][2] ) );
  DFF_X1 \mem_reg[411][1]  ( .D(n22817), .CK(clk), .Q(\mem[411][1] ) );
  DFF_X1 \mem_reg[411][0]  ( .D(n22818), .CK(clk), .Q(\mem[411][0] ) );
  DFF_X1 \mem_reg[410][7]  ( .D(n22819), .CK(clk), .Q(\mem[410][7] ) );
  DFF_X1 \mem_reg[410][6]  ( .D(n22820), .CK(clk), .Q(\mem[410][6] ) );
  DFF_X1 \mem_reg[410][5]  ( .D(n22821), .CK(clk), .Q(\mem[410][5] ) );
  DFF_X1 \mem_reg[410][4]  ( .D(n22822), .CK(clk), .Q(\mem[410][4] ) );
  DFF_X1 \mem_reg[410][3]  ( .D(n22823), .CK(clk), .Q(\mem[410][3] ) );
  DFF_X1 \mem_reg[410][2]  ( .D(n22824), .CK(clk), .Q(\mem[410][2] ) );
  DFF_X1 \mem_reg[410][1]  ( .D(n22825), .CK(clk), .Q(\mem[410][1] ) );
  DFF_X1 \mem_reg[410][0]  ( .D(n22826), .CK(clk), .Q(\mem[410][0] ) );
  DFF_X1 \mem_reg[409][7]  ( .D(n22827), .CK(clk), .Q(\mem[409][7] ) );
  DFF_X1 \mem_reg[409][6]  ( .D(n22828), .CK(clk), .Q(\mem[409][6] ) );
  DFF_X1 \mem_reg[409][5]  ( .D(n22829), .CK(clk), .Q(\mem[409][5] ) );
  DFF_X1 \mem_reg[409][4]  ( .D(n22830), .CK(clk), .Q(\mem[409][4] ) );
  DFF_X1 \mem_reg[409][3]  ( .D(n22831), .CK(clk), .Q(\mem[409][3] ) );
  DFF_X1 \mem_reg[409][2]  ( .D(n22832), .CK(clk), .Q(\mem[409][2] ) );
  DFF_X1 \mem_reg[409][1]  ( .D(n22833), .CK(clk), .Q(\mem[409][1] ) );
  DFF_X1 \mem_reg[409][0]  ( .D(n22834), .CK(clk), .Q(\mem[409][0] ) );
  DFF_X1 \mem_reg[408][7]  ( .D(n22835), .CK(clk), .Q(\mem[408][7] ) );
  DFF_X1 \mem_reg[408][6]  ( .D(n22836), .CK(clk), .Q(\mem[408][6] ) );
  DFF_X1 \mem_reg[408][5]  ( .D(n22837), .CK(clk), .Q(\mem[408][5] ) );
  DFF_X1 \mem_reg[408][4]  ( .D(n22838), .CK(clk), .Q(\mem[408][4] ) );
  DFF_X1 \mem_reg[408][3]  ( .D(n22839), .CK(clk), .Q(\mem[408][3] ) );
  DFF_X1 \mem_reg[408][2]  ( .D(n22840), .CK(clk), .Q(\mem[408][2] ) );
  DFF_X1 \mem_reg[408][1]  ( .D(n22841), .CK(clk), .Q(\mem[408][1] ) );
  DFF_X1 \mem_reg[408][0]  ( .D(n22842), .CK(clk), .Q(\mem[408][0] ) );
  DFF_X1 \mem_reg[407][7]  ( .D(n22843), .CK(clk), .Q(\mem[407][7] ) );
  DFF_X1 \mem_reg[407][6]  ( .D(n22844), .CK(clk), .Q(\mem[407][6] ) );
  DFF_X1 \mem_reg[407][5]  ( .D(n22845), .CK(clk), .Q(\mem[407][5] ) );
  DFF_X1 \mem_reg[407][4]  ( .D(n22846), .CK(clk), .Q(\mem[407][4] ) );
  DFF_X1 \mem_reg[407][3]  ( .D(n22847), .CK(clk), .Q(\mem[407][3] ) );
  DFF_X1 \mem_reg[407][2]  ( .D(n22848), .CK(clk), .Q(\mem[407][2] ) );
  DFF_X1 \mem_reg[407][1]  ( .D(n22849), .CK(clk), .Q(\mem[407][1] ) );
  DFF_X1 \mem_reg[407][0]  ( .D(n22850), .CK(clk), .Q(\mem[407][0] ) );
  DFF_X1 \mem_reg[406][7]  ( .D(n22851), .CK(clk), .Q(\mem[406][7] ) );
  DFF_X1 \mem_reg[406][6]  ( .D(n22852), .CK(clk), .Q(\mem[406][6] ) );
  DFF_X1 \mem_reg[406][5]  ( .D(n22853), .CK(clk), .Q(\mem[406][5] ) );
  DFF_X1 \mem_reg[406][4]  ( .D(n22854), .CK(clk), .Q(\mem[406][4] ) );
  DFF_X1 \mem_reg[406][3]  ( .D(n22855), .CK(clk), .Q(\mem[406][3] ) );
  DFF_X1 \mem_reg[406][2]  ( .D(n22856), .CK(clk), .Q(\mem[406][2] ) );
  DFF_X1 \mem_reg[406][1]  ( .D(n22857), .CK(clk), .Q(\mem[406][1] ) );
  DFF_X1 \mem_reg[406][0]  ( .D(n22858), .CK(clk), .Q(\mem[406][0] ) );
  DFF_X1 \mem_reg[405][7]  ( .D(n22859), .CK(clk), .Q(\mem[405][7] ) );
  DFF_X1 \mem_reg[405][6]  ( .D(n22860), .CK(clk), .Q(\mem[405][6] ) );
  DFF_X1 \mem_reg[405][5]  ( .D(n22861), .CK(clk), .Q(\mem[405][5] ) );
  DFF_X1 \mem_reg[405][4]  ( .D(n22862), .CK(clk), .Q(\mem[405][4] ) );
  DFF_X1 \mem_reg[405][3]  ( .D(n22863), .CK(clk), .Q(\mem[405][3] ) );
  DFF_X1 \mem_reg[405][2]  ( .D(n22864), .CK(clk), .Q(\mem[405][2] ) );
  DFF_X1 \mem_reg[405][1]  ( .D(n22865), .CK(clk), .Q(\mem[405][1] ) );
  DFF_X1 \mem_reg[405][0]  ( .D(n22866), .CK(clk), .Q(\mem[405][0] ) );
  DFF_X1 \mem_reg[404][7]  ( .D(n22867), .CK(clk), .Q(\mem[404][7] ) );
  DFF_X1 \mem_reg[404][6]  ( .D(n22868), .CK(clk), .Q(\mem[404][6] ) );
  DFF_X1 \mem_reg[404][5]  ( .D(n22869), .CK(clk), .Q(\mem[404][5] ) );
  DFF_X1 \mem_reg[404][4]  ( .D(n22870), .CK(clk), .Q(\mem[404][4] ) );
  DFF_X1 \mem_reg[404][3]  ( .D(n22871), .CK(clk), .Q(\mem[404][3] ) );
  DFF_X1 \mem_reg[404][2]  ( .D(n22872), .CK(clk), .Q(\mem[404][2] ) );
  DFF_X1 \mem_reg[404][1]  ( .D(n22873), .CK(clk), .Q(\mem[404][1] ) );
  DFF_X1 \mem_reg[404][0]  ( .D(n22874), .CK(clk), .Q(\mem[404][0] ) );
  DFF_X1 \mem_reg[403][7]  ( .D(n22875), .CK(clk), .Q(\mem[403][7] ) );
  DFF_X1 \mem_reg[403][6]  ( .D(n22876), .CK(clk), .Q(\mem[403][6] ) );
  DFF_X1 \mem_reg[403][5]  ( .D(n22877), .CK(clk), .Q(\mem[403][5] ) );
  DFF_X1 \mem_reg[403][4]  ( .D(n22878), .CK(clk), .Q(\mem[403][4] ) );
  DFF_X1 \mem_reg[403][3]  ( .D(n22879), .CK(clk), .Q(\mem[403][3] ) );
  DFF_X1 \mem_reg[403][2]  ( .D(n22880), .CK(clk), .Q(\mem[403][2] ) );
  DFF_X1 \mem_reg[403][1]  ( .D(n22881), .CK(clk), .Q(\mem[403][1] ) );
  DFF_X1 \mem_reg[403][0]  ( .D(n22882), .CK(clk), .Q(\mem[403][0] ) );
  DFF_X1 \mem_reg[402][7]  ( .D(n22883), .CK(clk), .Q(\mem[402][7] ) );
  DFF_X1 \mem_reg[402][6]  ( .D(n22884), .CK(clk), .Q(\mem[402][6] ) );
  DFF_X1 \mem_reg[402][5]  ( .D(n22885), .CK(clk), .Q(\mem[402][5] ) );
  DFF_X1 \mem_reg[402][4]  ( .D(n22886), .CK(clk), .Q(\mem[402][4] ) );
  DFF_X1 \mem_reg[402][3]  ( .D(n22887), .CK(clk), .Q(\mem[402][3] ) );
  DFF_X1 \mem_reg[402][2]  ( .D(n22888), .CK(clk), .Q(\mem[402][2] ) );
  DFF_X1 \mem_reg[402][1]  ( .D(n22889), .CK(clk), .Q(\mem[402][1] ) );
  DFF_X1 \mem_reg[402][0]  ( .D(n22890), .CK(clk), .Q(\mem[402][0] ) );
  DFF_X1 \mem_reg[401][7]  ( .D(n22891), .CK(clk), .Q(\mem[401][7] ) );
  DFF_X1 \mem_reg[401][6]  ( .D(n22892), .CK(clk), .Q(\mem[401][6] ) );
  DFF_X1 \mem_reg[401][5]  ( .D(n22893), .CK(clk), .Q(\mem[401][5] ) );
  DFF_X1 \mem_reg[401][4]  ( .D(n22894), .CK(clk), .Q(\mem[401][4] ) );
  DFF_X1 \mem_reg[401][3]  ( .D(n22895), .CK(clk), .Q(\mem[401][3] ) );
  DFF_X1 \mem_reg[401][2]  ( .D(n22896), .CK(clk), .Q(\mem[401][2] ) );
  DFF_X1 \mem_reg[401][1]  ( .D(n22897), .CK(clk), .Q(\mem[401][1] ) );
  DFF_X1 \mem_reg[401][0]  ( .D(n22898), .CK(clk), .Q(\mem[401][0] ) );
  DFF_X1 \mem_reg[400][7]  ( .D(n22899), .CK(clk), .Q(\mem[400][7] ) );
  DFF_X1 \mem_reg[400][6]  ( .D(n22900), .CK(clk), .Q(\mem[400][6] ) );
  DFF_X1 \mem_reg[400][5]  ( .D(n22901), .CK(clk), .Q(\mem[400][5] ) );
  DFF_X1 \mem_reg[400][4]  ( .D(n22902), .CK(clk), .Q(\mem[400][4] ) );
  DFF_X1 \mem_reg[400][3]  ( .D(n22903), .CK(clk), .Q(\mem[400][3] ) );
  DFF_X1 \mem_reg[400][2]  ( .D(n22904), .CK(clk), .Q(\mem[400][2] ) );
  DFF_X1 \mem_reg[400][1]  ( .D(n22905), .CK(clk), .Q(\mem[400][1] ) );
  DFF_X1 \mem_reg[400][0]  ( .D(n22906), .CK(clk), .Q(\mem[400][0] ) );
  DFF_X1 \mem_reg[399][7]  ( .D(n22907), .CK(clk), .Q(\mem[399][7] ) );
  DFF_X1 \mem_reg[399][6]  ( .D(n22908), .CK(clk), .Q(\mem[399][6] ) );
  DFF_X1 \mem_reg[399][5]  ( .D(n22909), .CK(clk), .Q(\mem[399][5] ) );
  DFF_X1 \mem_reg[399][4]  ( .D(n22910), .CK(clk), .Q(\mem[399][4] ) );
  DFF_X1 \mem_reg[399][3]  ( .D(n22911), .CK(clk), .Q(\mem[399][3] ) );
  DFF_X1 \mem_reg[399][2]  ( .D(n22912), .CK(clk), .Q(\mem[399][2] ) );
  DFF_X1 \mem_reg[399][1]  ( .D(n22913), .CK(clk), .Q(\mem[399][1] ) );
  DFF_X1 \mem_reg[399][0]  ( .D(n22914), .CK(clk), .Q(\mem[399][0] ) );
  DFF_X1 \mem_reg[398][7]  ( .D(n22915), .CK(clk), .Q(\mem[398][7] ) );
  DFF_X1 \mem_reg[398][6]  ( .D(n22916), .CK(clk), .Q(\mem[398][6] ) );
  DFF_X1 \mem_reg[398][5]  ( .D(n22917), .CK(clk), .Q(\mem[398][5] ) );
  DFF_X1 \mem_reg[398][4]  ( .D(n22918), .CK(clk), .Q(\mem[398][4] ) );
  DFF_X1 \mem_reg[398][3]  ( .D(n22919), .CK(clk), .Q(\mem[398][3] ) );
  DFF_X1 \mem_reg[398][2]  ( .D(n22920), .CK(clk), .Q(\mem[398][2] ) );
  DFF_X1 \mem_reg[398][1]  ( .D(n22921), .CK(clk), .Q(\mem[398][1] ) );
  DFF_X1 \mem_reg[398][0]  ( .D(n22922), .CK(clk), .Q(\mem[398][0] ) );
  DFF_X1 \mem_reg[397][7]  ( .D(n22923), .CK(clk), .Q(\mem[397][7] ) );
  DFF_X1 \mem_reg[397][6]  ( .D(n22924), .CK(clk), .Q(\mem[397][6] ) );
  DFF_X1 \mem_reg[397][5]  ( .D(n22925), .CK(clk), .Q(\mem[397][5] ) );
  DFF_X1 \mem_reg[397][4]  ( .D(n22926), .CK(clk), .Q(\mem[397][4] ) );
  DFF_X1 \mem_reg[397][3]  ( .D(n22927), .CK(clk), .Q(\mem[397][3] ) );
  DFF_X1 \mem_reg[397][2]  ( .D(n22928), .CK(clk), .Q(\mem[397][2] ) );
  DFF_X1 \mem_reg[397][1]  ( .D(n22929), .CK(clk), .Q(\mem[397][1] ) );
  DFF_X1 \mem_reg[397][0]  ( .D(n22930), .CK(clk), .Q(\mem[397][0] ) );
  DFF_X1 \mem_reg[396][7]  ( .D(n22931), .CK(clk), .Q(\mem[396][7] ) );
  DFF_X1 \mem_reg[396][6]  ( .D(n22932), .CK(clk), .Q(\mem[396][6] ) );
  DFF_X1 \mem_reg[396][5]  ( .D(n22933), .CK(clk), .Q(\mem[396][5] ) );
  DFF_X1 \mem_reg[396][4]  ( .D(n22934), .CK(clk), .Q(\mem[396][4] ) );
  DFF_X1 \mem_reg[396][3]  ( .D(n22935), .CK(clk), .Q(\mem[396][3] ) );
  DFF_X1 \mem_reg[396][2]  ( .D(n22936), .CK(clk), .Q(\mem[396][2] ) );
  DFF_X1 \mem_reg[396][1]  ( .D(n22937), .CK(clk), .Q(\mem[396][1] ) );
  DFF_X1 \mem_reg[396][0]  ( .D(n22938), .CK(clk), .Q(\mem[396][0] ) );
  DFF_X1 \mem_reg[395][7]  ( .D(n22939), .CK(clk), .Q(\mem[395][7] ) );
  DFF_X1 \mem_reg[395][6]  ( .D(n22940), .CK(clk), .Q(\mem[395][6] ) );
  DFF_X1 \mem_reg[395][5]  ( .D(n22941), .CK(clk), .Q(\mem[395][5] ) );
  DFF_X1 \mem_reg[395][4]  ( .D(n22942), .CK(clk), .Q(\mem[395][4] ) );
  DFF_X1 \mem_reg[395][3]  ( .D(n22943), .CK(clk), .Q(\mem[395][3] ) );
  DFF_X1 \mem_reg[395][2]  ( .D(n22944), .CK(clk), .Q(\mem[395][2] ) );
  DFF_X1 \mem_reg[395][1]  ( .D(n22945), .CK(clk), .Q(\mem[395][1] ) );
  DFF_X1 \mem_reg[395][0]  ( .D(n22946), .CK(clk), .Q(\mem[395][0] ) );
  DFF_X1 \mem_reg[394][7]  ( .D(n22947), .CK(clk), .Q(\mem[394][7] ) );
  DFF_X1 \mem_reg[394][6]  ( .D(n22948), .CK(clk), .Q(\mem[394][6] ) );
  DFF_X1 \mem_reg[394][5]  ( .D(n22949), .CK(clk), .Q(\mem[394][5] ) );
  DFF_X1 \mem_reg[394][4]  ( .D(n22950), .CK(clk), .Q(\mem[394][4] ) );
  DFF_X1 \mem_reg[394][3]  ( .D(n22951), .CK(clk), .Q(\mem[394][3] ) );
  DFF_X1 \mem_reg[394][2]  ( .D(n22952), .CK(clk), .Q(\mem[394][2] ) );
  DFF_X1 \mem_reg[394][1]  ( .D(n22953), .CK(clk), .Q(\mem[394][1] ) );
  DFF_X1 \mem_reg[394][0]  ( .D(n22954), .CK(clk), .Q(\mem[394][0] ) );
  DFF_X1 \mem_reg[393][7]  ( .D(n22955), .CK(clk), .Q(\mem[393][7] ) );
  DFF_X1 \mem_reg[393][6]  ( .D(n22956), .CK(clk), .Q(\mem[393][6] ) );
  DFF_X1 \mem_reg[393][5]  ( .D(n22957), .CK(clk), .Q(\mem[393][5] ) );
  DFF_X1 \mem_reg[393][4]  ( .D(n22958), .CK(clk), .Q(\mem[393][4] ) );
  DFF_X1 \mem_reg[393][3]  ( .D(n22959), .CK(clk), .Q(\mem[393][3] ) );
  DFF_X1 \mem_reg[393][2]  ( .D(n22960), .CK(clk), .Q(\mem[393][2] ) );
  DFF_X1 \mem_reg[393][1]  ( .D(n22961), .CK(clk), .Q(\mem[393][1] ) );
  DFF_X1 \mem_reg[393][0]  ( .D(n22962), .CK(clk), .Q(\mem[393][0] ) );
  DFF_X1 \mem_reg[392][7]  ( .D(n22963), .CK(clk), .Q(\mem[392][7] ) );
  DFF_X1 \mem_reg[392][6]  ( .D(n22964), .CK(clk), .Q(\mem[392][6] ) );
  DFF_X1 \mem_reg[392][5]  ( .D(n22965), .CK(clk), .Q(\mem[392][5] ) );
  DFF_X1 \mem_reg[392][4]  ( .D(n22966), .CK(clk), .Q(\mem[392][4] ) );
  DFF_X1 \mem_reg[392][3]  ( .D(n22967), .CK(clk), .Q(\mem[392][3] ) );
  DFF_X1 \mem_reg[392][2]  ( .D(n22968), .CK(clk), .Q(\mem[392][2] ) );
  DFF_X1 \mem_reg[392][1]  ( .D(n22969), .CK(clk), .Q(\mem[392][1] ) );
  DFF_X1 \mem_reg[392][0]  ( .D(n22970), .CK(clk), .Q(\mem[392][0] ) );
  DFF_X1 \mem_reg[391][7]  ( .D(n22971), .CK(clk), .Q(\mem[391][7] ) );
  DFF_X1 \mem_reg[391][6]  ( .D(n22972), .CK(clk), .Q(\mem[391][6] ) );
  DFF_X1 \mem_reg[391][5]  ( .D(n22973), .CK(clk), .Q(\mem[391][5] ) );
  DFF_X1 \mem_reg[391][4]  ( .D(n22974), .CK(clk), .Q(\mem[391][4] ) );
  DFF_X1 \mem_reg[391][3]  ( .D(n22975), .CK(clk), .Q(\mem[391][3] ) );
  DFF_X1 \mem_reg[391][2]  ( .D(n22976), .CK(clk), .Q(\mem[391][2] ) );
  DFF_X1 \mem_reg[391][1]  ( .D(n22977), .CK(clk), .Q(\mem[391][1] ) );
  DFF_X1 \mem_reg[391][0]  ( .D(n22978), .CK(clk), .Q(\mem[391][0] ) );
  DFF_X1 \mem_reg[390][7]  ( .D(n22979), .CK(clk), .Q(\mem[390][7] ) );
  DFF_X1 \mem_reg[390][6]  ( .D(n22980), .CK(clk), .Q(\mem[390][6] ) );
  DFF_X1 \mem_reg[390][5]  ( .D(n22981), .CK(clk), .Q(\mem[390][5] ) );
  DFF_X1 \mem_reg[390][4]  ( .D(n22982), .CK(clk), .Q(\mem[390][4] ) );
  DFF_X1 \mem_reg[390][3]  ( .D(n22983), .CK(clk), .Q(\mem[390][3] ) );
  DFF_X1 \mem_reg[390][2]  ( .D(n22984), .CK(clk), .Q(\mem[390][2] ) );
  DFF_X1 \mem_reg[390][1]  ( .D(n22985), .CK(clk), .Q(\mem[390][1] ) );
  DFF_X1 \mem_reg[390][0]  ( .D(n22986), .CK(clk), .Q(\mem[390][0] ) );
  DFF_X1 \mem_reg[389][7]  ( .D(n22987), .CK(clk), .Q(\mem[389][7] ) );
  DFF_X1 \mem_reg[389][6]  ( .D(n22988), .CK(clk), .Q(\mem[389][6] ) );
  DFF_X1 \mem_reg[389][5]  ( .D(n22989), .CK(clk), .Q(\mem[389][5] ) );
  DFF_X1 \mem_reg[389][4]  ( .D(n22990), .CK(clk), .Q(\mem[389][4] ) );
  DFF_X1 \mem_reg[389][3]  ( .D(n22991), .CK(clk), .Q(\mem[389][3] ) );
  DFF_X1 \mem_reg[389][2]  ( .D(n22992), .CK(clk), .Q(\mem[389][2] ) );
  DFF_X1 \mem_reg[389][1]  ( .D(n22993), .CK(clk), .Q(\mem[389][1] ) );
  DFF_X1 \mem_reg[389][0]  ( .D(n22994), .CK(clk), .Q(\mem[389][0] ) );
  DFF_X1 \mem_reg[388][7]  ( .D(n22995), .CK(clk), .Q(\mem[388][7] ) );
  DFF_X1 \mem_reg[388][6]  ( .D(n22996), .CK(clk), .Q(\mem[388][6] ) );
  DFF_X1 \mem_reg[388][5]  ( .D(n22997), .CK(clk), .Q(\mem[388][5] ) );
  DFF_X1 \mem_reg[388][4]  ( .D(n22998), .CK(clk), .Q(\mem[388][4] ) );
  DFF_X1 \mem_reg[388][3]  ( .D(n22999), .CK(clk), .Q(\mem[388][3] ) );
  DFF_X1 \mem_reg[388][2]  ( .D(n23000), .CK(clk), .Q(\mem[388][2] ) );
  DFF_X1 \mem_reg[388][1]  ( .D(n23001), .CK(clk), .Q(\mem[388][1] ) );
  DFF_X1 \mem_reg[388][0]  ( .D(n23002), .CK(clk), .Q(\mem[388][0] ) );
  DFF_X1 \mem_reg[387][7]  ( .D(n23003), .CK(clk), .Q(\mem[387][7] ) );
  DFF_X1 \mem_reg[387][6]  ( .D(n23004), .CK(clk), .Q(\mem[387][6] ) );
  DFF_X1 \mem_reg[387][5]  ( .D(n23005), .CK(clk), .Q(\mem[387][5] ) );
  DFF_X1 \mem_reg[387][4]  ( .D(n23006), .CK(clk), .Q(\mem[387][4] ) );
  DFF_X1 \mem_reg[387][3]  ( .D(n23007), .CK(clk), .Q(\mem[387][3] ) );
  DFF_X1 \mem_reg[387][2]  ( .D(n23008), .CK(clk), .Q(\mem[387][2] ) );
  DFF_X1 \mem_reg[387][1]  ( .D(n23009), .CK(clk), .Q(\mem[387][1] ) );
  DFF_X1 \mem_reg[387][0]  ( .D(n23010), .CK(clk), .Q(\mem[387][0] ) );
  DFF_X1 \mem_reg[386][7]  ( .D(n23011), .CK(clk), .Q(\mem[386][7] ) );
  DFF_X1 \mem_reg[386][6]  ( .D(n23012), .CK(clk), .Q(\mem[386][6] ) );
  DFF_X1 \mem_reg[386][5]  ( .D(n23013), .CK(clk), .Q(\mem[386][5] ) );
  DFF_X1 \mem_reg[386][4]  ( .D(n23014), .CK(clk), .Q(\mem[386][4] ) );
  DFF_X1 \mem_reg[386][3]  ( .D(n23015), .CK(clk), .Q(\mem[386][3] ) );
  DFF_X1 \mem_reg[386][2]  ( .D(n23016), .CK(clk), .Q(\mem[386][2] ) );
  DFF_X1 \mem_reg[386][1]  ( .D(n23017), .CK(clk), .Q(\mem[386][1] ) );
  DFF_X1 \mem_reg[386][0]  ( .D(n23018), .CK(clk), .Q(\mem[386][0] ) );
  DFF_X1 \mem_reg[385][7]  ( .D(n23019), .CK(clk), .Q(\mem[385][7] ) );
  DFF_X1 \mem_reg[385][6]  ( .D(n23020), .CK(clk), .Q(\mem[385][6] ) );
  DFF_X1 \mem_reg[385][5]  ( .D(n23021), .CK(clk), .Q(\mem[385][5] ) );
  DFF_X1 \mem_reg[385][4]  ( .D(n23022), .CK(clk), .Q(\mem[385][4] ) );
  DFF_X1 \mem_reg[385][3]  ( .D(n23023), .CK(clk), .Q(\mem[385][3] ) );
  DFF_X1 \mem_reg[385][2]  ( .D(n23024), .CK(clk), .Q(\mem[385][2] ) );
  DFF_X1 \mem_reg[385][1]  ( .D(n23025), .CK(clk), .Q(\mem[385][1] ) );
  DFF_X1 \mem_reg[385][0]  ( .D(n23026), .CK(clk), .Q(\mem[385][0] ) );
  DFF_X1 \mem_reg[384][7]  ( .D(n23027), .CK(clk), .Q(\mem[384][7] ) );
  DFF_X1 \mem_reg[384][6]  ( .D(n23028), .CK(clk), .Q(\mem[384][6] ) );
  DFF_X1 \mem_reg[384][5]  ( .D(n23029), .CK(clk), .Q(\mem[384][5] ) );
  DFF_X1 \mem_reg[384][4]  ( .D(n23030), .CK(clk), .Q(\mem[384][4] ) );
  DFF_X1 \mem_reg[384][3]  ( .D(n23031), .CK(clk), .Q(\mem[384][3] ) );
  DFF_X1 \mem_reg[384][2]  ( .D(n23032), .CK(clk), .Q(\mem[384][2] ) );
  DFF_X1 \mem_reg[384][1]  ( .D(n23033), .CK(clk), .Q(\mem[384][1] ) );
  DFF_X1 \mem_reg[384][0]  ( .D(n23034), .CK(clk), .Q(\mem[384][0] ) );
  DFF_X1 \mem_reg[383][7]  ( .D(n23035), .CK(clk), .Q(\mem[383][7] ) );
  DFF_X1 \mem_reg[383][6]  ( .D(n23036), .CK(clk), .Q(\mem[383][6] ) );
  DFF_X1 \mem_reg[383][5]  ( .D(n23037), .CK(clk), .Q(\mem[383][5] ) );
  DFF_X1 \mem_reg[383][4]  ( .D(n23038), .CK(clk), .Q(\mem[383][4] ) );
  DFF_X1 \mem_reg[383][3]  ( .D(n23039), .CK(clk), .Q(\mem[383][3] ) );
  DFF_X1 \mem_reg[383][2]  ( .D(n23040), .CK(clk), .Q(\mem[383][2] ) );
  DFF_X1 \mem_reg[383][1]  ( .D(n23041), .CK(clk), .Q(\mem[383][1] ) );
  DFF_X1 \mem_reg[383][0]  ( .D(n23042), .CK(clk), .Q(\mem[383][0] ) );
  DFF_X1 \mem_reg[382][7]  ( .D(n23043), .CK(clk), .Q(\mem[382][7] ) );
  DFF_X1 \mem_reg[382][6]  ( .D(n23044), .CK(clk), .Q(\mem[382][6] ) );
  DFF_X1 \mem_reg[382][5]  ( .D(n23045), .CK(clk), .Q(\mem[382][5] ) );
  DFF_X1 \mem_reg[382][4]  ( .D(n23046), .CK(clk), .Q(\mem[382][4] ) );
  DFF_X1 \mem_reg[382][3]  ( .D(n23047), .CK(clk), .Q(\mem[382][3] ) );
  DFF_X1 \mem_reg[382][2]  ( .D(n23048), .CK(clk), .Q(\mem[382][2] ) );
  DFF_X1 \mem_reg[382][1]  ( .D(n23049), .CK(clk), .Q(\mem[382][1] ) );
  DFF_X1 \mem_reg[382][0]  ( .D(n23050), .CK(clk), .Q(\mem[382][0] ) );
  DFF_X1 \mem_reg[381][7]  ( .D(n23051), .CK(clk), .Q(\mem[381][7] ) );
  DFF_X1 \mem_reg[381][6]  ( .D(n23052), .CK(clk), .Q(\mem[381][6] ) );
  DFF_X1 \mem_reg[381][5]  ( .D(n23053), .CK(clk), .Q(\mem[381][5] ) );
  DFF_X1 \mem_reg[381][4]  ( .D(n23054), .CK(clk), .Q(\mem[381][4] ) );
  DFF_X1 \mem_reg[381][3]  ( .D(n23055), .CK(clk), .Q(\mem[381][3] ) );
  DFF_X1 \mem_reg[381][2]  ( .D(n23056), .CK(clk), .Q(\mem[381][2] ) );
  DFF_X1 \mem_reg[381][1]  ( .D(n23057), .CK(clk), .Q(\mem[381][1] ) );
  DFF_X1 \mem_reg[381][0]  ( .D(n23058), .CK(clk), .Q(\mem[381][0] ) );
  DFF_X1 \mem_reg[380][7]  ( .D(n23059), .CK(clk), .Q(\mem[380][7] ) );
  DFF_X1 \mem_reg[380][6]  ( .D(n23060), .CK(clk), .Q(\mem[380][6] ) );
  DFF_X1 \mem_reg[380][5]  ( .D(n23061), .CK(clk), .Q(\mem[380][5] ) );
  DFF_X1 \mem_reg[380][4]  ( .D(n23062), .CK(clk), .Q(\mem[380][4] ) );
  DFF_X1 \mem_reg[380][3]  ( .D(n23063), .CK(clk), .Q(\mem[380][3] ) );
  DFF_X1 \mem_reg[380][2]  ( .D(n23064), .CK(clk), .Q(\mem[380][2] ) );
  DFF_X1 \mem_reg[380][1]  ( .D(n23065), .CK(clk), .Q(\mem[380][1] ) );
  DFF_X1 \mem_reg[380][0]  ( .D(n23066), .CK(clk), .Q(\mem[380][0] ) );
  DFF_X1 \mem_reg[379][7]  ( .D(n23067), .CK(clk), .Q(\mem[379][7] ) );
  DFF_X1 \mem_reg[379][6]  ( .D(n23068), .CK(clk), .Q(\mem[379][6] ) );
  DFF_X1 \mem_reg[379][5]  ( .D(n23069), .CK(clk), .Q(\mem[379][5] ) );
  DFF_X1 \mem_reg[379][4]  ( .D(n23070), .CK(clk), .Q(\mem[379][4] ) );
  DFF_X1 \mem_reg[379][3]  ( .D(n23071), .CK(clk), .Q(\mem[379][3] ) );
  DFF_X1 \mem_reg[379][2]  ( .D(n23072), .CK(clk), .Q(\mem[379][2] ) );
  DFF_X1 \mem_reg[379][1]  ( .D(n23073), .CK(clk), .Q(\mem[379][1] ) );
  DFF_X1 \mem_reg[379][0]  ( .D(n23074), .CK(clk), .Q(\mem[379][0] ) );
  DFF_X1 \mem_reg[378][7]  ( .D(n23075), .CK(clk), .Q(\mem[378][7] ) );
  DFF_X1 \mem_reg[378][6]  ( .D(n23076), .CK(clk), .Q(\mem[378][6] ) );
  DFF_X1 \mem_reg[378][5]  ( .D(n23077), .CK(clk), .Q(\mem[378][5] ) );
  DFF_X1 \mem_reg[378][4]  ( .D(n23078), .CK(clk), .Q(\mem[378][4] ) );
  DFF_X1 \mem_reg[378][3]  ( .D(n23079), .CK(clk), .Q(\mem[378][3] ) );
  DFF_X1 \mem_reg[378][2]  ( .D(n23080), .CK(clk), .Q(\mem[378][2] ) );
  DFF_X1 \mem_reg[378][1]  ( .D(n23081), .CK(clk), .Q(\mem[378][1] ) );
  DFF_X1 \mem_reg[378][0]  ( .D(n23082), .CK(clk), .Q(\mem[378][0] ) );
  DFF_X1 \mem_reg[377][7]  ( .D(n23083), .CK(clk), .Q(\mem[377][7] ) );
  DFF_X1 \mem_reg[377][6]  ( .D(n23084), .CK(clk), .Q(\mem[377][6] ) );
  DFF_X1 \mem_reg[377][5]  ( .D(n23085), .CK(clk), .Q(\mem[377][5] ) );
  DFF_X1 \mem_reg[377][4]  ( .D(n23086), .CK(clk), .Q(\mem[377][4] ) );
  DFF_X1 \mem_reg[377][3]  ( .D(n23087), .CK(clk), .Q(\mem[377][3] ) );
  DFF_X1 \mem_reg[377][2]  ( .D(n23088), .CK(clk), .Q(\mem[377][2] ) );
  DFF_X1 \mem_reg[377][1]  ( .D(n23089), .CK(clk), .Q(\mem[377][1] ) );
  DFF_X1 \mem_reg[377][0]  ( .D(n23090), .CK(clk), .Q(\mem[377][0] ) );
  DFF_X1 \mem_reg[376][7]  ( .D(n23091), .CK(clk), .Q(\mem[376][7] ) );
  DFF_X1 \mem_reg[376][6]  ( .D(n23092), .CK(clk), .Q(\mem[376][6] ) );
  DFF_X1 \mem_reg[376][5]  ( .D(n23093), .CK(clk), .Q(\mem[376][5] ) );
  DFF_X1 \mem_reg[376][4]  ( .D(n23094), .CK(clk), .Q(\mem[376][4] ) );
  DFF_X1 \mem_reg[376][3]  ( .D(n23095), .CK(clk), .Q(\mem[376][3] ) );
  DFF_X1 \mem_reg[376][2]  ( .D(n23096), .CK(clk), .Q(\mem[376][2] ) );
  DFF_X1 \mem_reg[376][1]  ( .D(n23097), .CK(clk), .Q(\mem[376][1] ) );
  DFF_X1 \mem_reg[376][0]  ( .D(n23098), .CK(clk), .Q(\mem[376][0] ) );
  DFF_X1 \mem_reg[375][7]  ( .D(n23099), .CK(clk), .Q(\mem[375][7] ) );
  DFF_X1 \mem_reg[375][6]  ( .D(n23100), .CK(clk), .Q(\mem[375][6] ) );
  DFF_X1 \mem_reg[375][5]  ( .D(n23101), .CK(clk), .Q(\mem[375][5] ) );
  DFF_X1 \mem_reg[375][4]  ( .D(n23102), .CK(clk), .Q(\mem[375][4] ) );
  DFF_X1 \mem_reg[375][3]  ( .D(n23103), .CK(clk), .Q(\mem[375][3] ) );
  DFF_X1 \mem_reg[375][2]  ( .D(n23104), .CK(clk), .Q(\mem[375][2] ) );
  DFF_X1 \mem_reg[375][1]  ( .D(n23105), .CK(clk), .Q(\mem[375][1] ) );
  DFF_X1 \mem_reg[375][0]  ( .D(n23106), .CK(clk), .Q(\mem[375][0] ) );
  DFF_X1 \mem_reg[374][7]  ( .D(n23107), .CK(clk), .Q(\mem[374][7] ) );
  DFF_X1 \mem_reg[374][6]  ( .D(n23108), .CK(clk), .Q(\mem[374][6] ) );
  DFF_X1 \mem_reg[374][5]  ( .D(n23109), .CK(clk), .Q(\mem[374][5] ) );
  DFF_X1 \mem_reg[374][4]  ( .D(n23110), .CK(clk), .Q(\mem[374][4] ) );
  DFF_X1 \mem_reg[374][3]  ( .D(n23111), .CK(clk), .Q(\mem[374][3] ) );
  DFF_X1 \mem_reg[374][2]  ( .D(n23112), .CK(clk), .Q(\mem[374][2] ) );
  DFF_X1 \mem_reg[374][1]  ( .D(n23113), .CK(clk), .Q(\mem[374][1] ) );
  DFF_X1 \mem_reg[374][0]  ( .D(n23114), .CK(clk), .Q(\mem[374][0] ) );
  DFF_X1 \mem_reg[373][7]  ( .D(n23115), .CK(clk), .Q(\mem[373][7] ) );
  DFF_X1 \mem_reg[373][6]  ( .D(n23116), .CK(clk), .Q(\mem[373][6] ) );
  DFF_X1 \mem_reg[373][5]  ( .D(n23117), .CK(clk), .Q(\mem[373][5] ) );
  DFF_X1 \mem_reg[373][4]  ( .D(n23118), .CK(clk), .Q(\mem[373][4] ) );
  DFF_X1 \mem_reg[373][3]  ( .D(n23119), .CK(clk), .Q(\mem[373][3] ) );
  DFF_X1 \mem_reg[373][2]  ( .D(n23120), .CK(clk), .Q(\mem[373][2] ) );
  DFF_X1 \mem_reg[373][1]  ( .D(n23121), .CK(clk), .Q(\mem[373][1] ) );
  DFF_X1 \mem_reg[373][0]  ( .D(n23122), .CK(clk), .Q(\mem[373][0] ) );
  DFF_X1 \mem_reg[372][7]  ( .D(n23123), .CK(clk), .Q(\mem[372][7] ) );
  DFF_X1 \mem_reg[372][6]  ( .D(n23124), .CK(clk), .Q(\mem[372][6] ) );
  DFF_X1 \mem_reg[372][5]  ( .D(n23125), .CK(clk), .Q(\mem[372][5] ) );
  DFF_X1 \mem_reg[372][4]  ( .D(n23126), .CK(clk), .Q(\mem[372][4] ) );
  DFF_X1 \mem_reg[372][3]  ( .D(n23127), .CK(clk), .Q(\mem[372][3] ) );
  DFF_X1 \mem_reg[372][2]  ( .D(n23128), .CK(clk), .Q(\mem[372][2] ) );
  DFF_X1 \mem_reg[372][1]  ( .D(n23129), .CK(clk), .Q(\mem[372][1] ) );
  DFF_X1 \mem_reg[372][0]  ( .D(n23130), .CK(clk), .Q(\mem[372][0] ) );
  DFF_X1 \mem_reg[371][7]  ( .D(n23131), .CK(clk), .Q(\mem[371][7] ) );
  DFF_X1 \mem_reg[371][6]  ( .D(n23132), .CK(clk), .Q(\mem[371][6] ) );
  DFF_X1 \mem_reg[371][5]  ( .D(n23133), .CK(clk), .Q(\mem[371][5] ) );
  DFF_X1 \mem_reg[371][4]  ( .D(n23134), .CK(clk), .Q(\mem[371][4] ) );
  DFF_X1 \mem_reg[371][3]  ( .D(n23135), .CK(clk), .Q(\mem[371][3] ) );
  DFF_X1 \mem_reg[371][2]  ( .D(n23136), .CK(clk), .Q(\mem[371][2] ) );
  DFF_X1 \mem_reg[371][1]  ( .D(n23137), .CK(clk), .Q(\mem[371][1] ) );
  DFF_X1 \mem_reg[371][0]  ( .D(n23138), .CK(clk), .Q(\mem[371][0] ) );
  DFF_X1 \mem_reg[370][7]  ( .D(n23139), .CK(clk), .Q(\mem[370][7] ) );
  DFF_X1 \mem_reg[370][6]  ( .D(n23140), .CK(clk), .Q(\mem[370][6] ) );
  DFF_X1 \mem_reg[370][5]  ( .D(n23141), .CK(clk), .Q(\mem[370][5] ) );
  DFF_X1 \mem_reg[370][4]  ( .D(n23142), .CK(clk), .Q(\mem[370][4] ) );
  DFF_X1 \mem_reg[370][3]  ( .D(n23143), .CK(clk), .Q(\mem[370][3] ) );
  DFF_X1 \mem_reg[370][2]  ( .D(n23144), .CK(clk), .Q(\mem[370][2] ) );
  DFF_X1 \mem_reg[370][1]  ( .D(n23145), .CK(clk), .Q(\mem[370][1] ) );
  DFF_X1 \mem_reg[370][0]  ( .D(n23146), .CK(clk), .Q(\mem[370][0] ) );
  DFF_X1 \mem_reg[369][7]  ( .D(n23147), .CK(clk), .Q(\mem[369][7] ) );
  DFF_X1 \mem_reg[369][6]  ( .D(n23148), .CK(clk), .Q(\mem[369][6] ) );
  DFF_X1 \mem_reg[369][5]  ( .D(n23149), .CK(clk), .Q(\mem[369][5] ) );
  DFF_X1 \mem_reg[369][4]  ( .D(n23150), .CK(clk), .Q(\mem[369][4] ) );
  DFF_X1 \mem_reg[369][3]  ( .D(n23151), .CK(clk), .Q(\mem[369][3] ) );
  DFF_X1 \mem_reg[369][2]  ( .D(n23152), .CK(clk), .Q(\mem[369][2] ) );
  DFF_X1 \mem_reg[369][1]  ( .D(n23153), .CK(clk), .Q(\mem[369][1] ) );
  DFF_X1 \mem_reg[369][0]  ( .D(n23154), .CK(clk), .Q(\mem[369][0] ) );
  DFF_X1 \mem_reg[368][7]  ( .D(n23155), .CK(clk), .Q(\mem[368][7] ) );
  DFF_X1 \mem_reg[368][6]  ( .D(n23156), .CK(clk), .Q(\mem[368][6] ) );
  DFF_X1 \mem_reg[368][5]  ( .D(n23157), .CK(clk), .Q(\mem[368][5] ) );
  DFF_X1 \mem_reg[368][4]  ( .D(n23158), .CK(clk), .Q(\mem[368][4] ) );
  DFF_X1 \mem_reg[368][3]  ( .D(n23159), .CK(clk), .Q(\mem[368][3] ) );
  DFF_X1 \mem_reg[368][2]  ( .D(n23160), .CK(clk), .Q(\mem[368][2] ) );
  DFF_X1 \mem_reg[368][1]  ( .D(n23161), .CK(clk), .Q(\mem[368][1] ) );
  DFF_X1 \mem_reg[368][0]  ( .D(n23162), .CK(clk), .Q(\mem[368][0] ) );
  DFF_X1 \mem_reg[367][7]  ( .D(n23163), .CK(clk), .Q(\mem[367][7] ) );
  DFF_X1 \mem_reg[367][6]  ( .D(n23164), .CK(clk), .Q(\mem[367][6] ) );
  DFF_X1 \mem_reg[367][5]  ( .D(n23165), .CK(clk), .Q(\mem[367][5] ) );
  DFF_X1 \mem_reg[367][4]  ( .D(n23166), .CK(clk), .Q(\mem[367][4] ) );
  DFF_X1 \mem_reg[367][3]  ( .D(n23167), .CK(clk), .Q(\mem[367][3] ) );
  DFF_X1 \mem_reg[367][2]  ( .D(n23168), .CK(clk), .Q(\mem[367][2] ) );
  DFF_X1 \mem_reg[367][1]  ( .D(n23169), .CK(clk), .Q(\mem[367][1] ) );
  DFF_X1 \mem_reg[367][0]  ( .D(n23170), .CK(clk), .Q(\mem[367][0] ) );
  DFF_X1 \mem_reg[366][7]  ( .D(n23171), .CK(clk), .Q(\mem[366][7] ) );
  DFF_X1 \mem_reg[366][6]  ( .D(n23172), .CK(clk), .Q(\mem[366][6] ) );
  DFF_X1 \mem_reg[366][5]  ( .D(n23173), .CK(clk), .Q(\mem[366][5] ) );
  DFF_X1 \mem_reg[366][4]  ( .D(n23174), .CK(clk), .Q(\mem[366][4] ) );
  DFF_X1 \mem_reg[366][3]  ( .D(n23175), .CK(clk), .Q(\mem[366][3] ) );
  DFF_X1 \mem_reg[366][2]  ( .D(n23176), .CK(clk), .Q(\mem[366][2] ) );
  DFF_X1 \mem_reg[366][1]  ( .D(n23177), .CK(clk), .Q(\mem[366][1] ) );
  DFF_X1 \mem_reg[366][0]  ( .D(n23178), .CK(clk), .Q(\mem[366][0] ) );
  DFF_X1 \mem_reg[365][7]  ( .D(n23179), .CK(clk), .Q(\mem[365][7] ) );
  DFF_X1 \mem_reg[365][6]  ( .D(n23180), .CK(clk), .Q(\mem[365][6] ) );
  DFF_X1 \mem_reg[365][5]  ( .D(n23181), .CK(clk), .Q(\mem[365][5] ) );
  DFF_X1 \mem_reg[365][4]  ( .D(n23182), .CK(clk), .Q(\mem[365][4] ) );
  DFF_X1 \mem_reg[365][3]  ( .D(n23183), .CK(clk), .Q(\mem[365][3] ) );
  DFF_X1 \mem_reg[365][2]  ( .D(n23184), .CK(clk), .Q(\mem[365][2] ) );
  DFF_X1 \mem_reg[365][1]  ( .D(n23185), .CK(clk), .Q(\mem[365][1] ) );
  DFF_X1 \mem_reg[365][0]  ( .D(n23186), .CK(clk), .Q(\mem[365][0] ) );
  DFF_X1 \mem_reg[364][7]  ( .D(n23187), .CK(clk), .Q(\mem[364][7] ) );
  DFF_X1 \mem_reg[364][6]  ( .D(n23188), .CK(clk), .Q(\mem[364][6] ) );
  DFF_X1 \mem_reg[364][5]  ( .D(n23189), .CK(clk), .Q(\mem[364][5] ) );
  DFF_X1 \mem_reg[364][4]  ( .D(n23190), .CK(clk), .Q(\mem[364][4] ) );
  DFF_X1 \mem_reg[364][3]  ( .D(n23191), .CK(clk), .Q(\mem[364][3] ) );
  DFF_X1 \mem_reg[364][2]  ( .D(n23192), .CK(clk), .Q(\mem[364][2] ) );
  DFF_X1 \mem_reg[364][1]  ( .D(n23193), .CK(clk), .Q(\mem[364][1] ) );
  DFF_X1 \mem_reg[364][0]  ( .D(n23194), .CK(clk), .Q(\mem[364][0] ) );
  DFF_X1 \mem_reg[363][7]  ( .D(n23195), .CK(clk), .Q(\mem[363][7] ) );
  DFF_X1 \mem_reg[363][6]  ( .D(n23196), .CK(clk), .Q(\mem[363][6] ) );
  DFF_X1 \mem_reg[363][5]  ( .D(n23197), .CK(clk), .Q(\mem[363][5] ) );
  DFF_X1 \mem_reg[363][4]  ( .D(n23198), .CK(clk), .Q(\mem[363][4] ) );
  DFF_X1 \mem_reg[363][3]  ( .D(n23199), .CK(clk), .Q(\mem[363][3] ) );
  DFF_X1 \mem_reg[363][2]  ( .D(n23200), .CK(clk), .Q(\mem[363][2] ) );
  DFF_X1 \mem_reg[363][1]  ( .D(n23201), .CK(clk), .Q(\mem[363][1] ) );
  DFF_X1 \mem_reg[363][0]  ( .D(n23202), .CK(clk), .Q(\mem[363][0] ) );
  DFF_X1 \mem_reg[362][7]  ( .D(n23203), .CK(clk), .Q(\mem[362][7] ) );
  DFF_X1 \mem_reg[362][6]  ( .D(n23204), .CK(clk), .Q(\mem[362][6] ) );
  DFF_X1 \mem_reg[362][5]  ( .D(n23205), .CK(clk), .Q(\mem[362][5] ) );
  DFF_X1 \mem_reg[362][4]  ( .D(n23206), .CK(clk), .Q(\mem[362][4] ) );
  DFF_X1 \mem_reg[362][3]  ( .D(n23207), .CK(clk), .Q(\mem[362][3] ) );
  DFF_X1 \mem_reg[362][2]  ( .D(n23208), .CK(clk), .Q(\mem[362][2] ) );
  DFF_X1 \mem_reg[362][1]  ( .D(n23209), .CK(clk), .Q(\mem[362][1] ) );
  DFF_X1 \mem_reg[362][0]  ( .D(n23210), .CK(clk), .Q(\mem[362][0] ) );
  DFF_X1 \mem_reg[361][7]  ( .D(n23211), .CK(clk), .Q(\mem[361][7] ) );
  DFF_X1 \mem_reg[361][6]  ( .D(n23212), .CK(clk), .Q(\mem[361][6] ) );
  DFF_X1 \mem_reg[361][5]  ( .D(n23213), .CK(clk), .Q(\mem[361][5] ) );
  DFF_X1 \mem_reg[361][4]  ( .D(n23214), .CK(clk), .Q(\mem[361][4] ) );
  DFF_X1 \mem_reg[361][3]  ( .D(n23215), .CK(clk), .Q(\mem[361][3] ) );
  DFF_X1 \mem_reg[361][2]  ( .D(n23216), .CK(clk), .Q(\mem[361][2] ) );
  DFF_X1 \mem_reg[361][1]  ( .D(n23217), .CK(clk), .Q(\mem[361][1] ) );
  DFF_X1 \mem_reg[361][0]  ( .D(n23218), .CK(clk), .Q(\mem[361][0] ) );
  DFF_X1 \mem_reg[360][7]  ( .D(n23219), .CK(clk), .Q(\mem[360][7] ) );
  DFF_X1 \mem_reg[360][6]  ( .D(n23220), .CK(clk), .Q(\mem[360][6] ) );
  DFF_X1 \mem_reg[360][5]  ( .D(n23221), .CK(clk), .Q(\mem[360][5] ) );
  DFF_X1 \mem_reg[360][4]  ( .D(n23222), .CK(clk), .Q(\mem[360][4] ) );
  DFF_X1 \mem_reg[360][3]  ( .D(n23223), .CK(clk), .Q(\mem[360][3] ) );
  DFF_X1 \mem_reg[360][2]  ( .D(n23224), .CK(clk), .Q(\mem[360][2] ) );
  DFF_X1 \mem_reg[360][1]  ( .D(n23225), .CK(clk), .Q(\mem[360][1] ) );
  DFF_X1 \mem_reg[360][0]  ( .D(n23226), .CK(clk), .Q(\mem[360][0] ) );
  DFF_X1 \mem_reg[359][7]  ( .D(n23227), .CK(clk), .Q(\mem[359][7] ) );
  DFF_X1 \mem_reg[359][6]  ( .D(n23228), .CK(clk), .Q(\mem[359][6] ) );
  DFF_X1 \mem_reg[359][5]  ( .D(n23229), .CK(clk), .Q(\mem[359][5] ) );
  DFF_X1 \mem_reg[359][4]  ( .D(n23230), .CK(clk), .Q(\mem[359][4] ) );
  DFF_X1 \mem_reg[359][3]  ( .D(n23231), .CK(clk), .Q(\mem[359][3] ) );
  DFF_X1 \mem_reg[359][2]  ( .D(n23232), .CK(clk), .Q(\mem[359][2] ) );
  DFF_X1 \mem_reg[359][1]  ( .D(n23233), .CK(clk), .Q(\mem[359][1] ) );
  DFF_X1 \mem_reg[359][0]  ( .D(n23234), .CK(clk), .Q(\mem[359][0] ) );
  DFF_X1 \mem_reg[358][7]  ( .D(n23235), .CK(clk), .Q(\mem[358][7] ) );
  DFF_X1 \mem_reg[358][6]  ( .D(n23236), .CK(clk), .Q(\mem[358][6] ) );
  DFF_X1 \mem_reg[358][5]  ( .D(n23237), .CK(clk), .Q(\mem[358][5] ) );
  DFF_X1 \mem_reg[358][4]  ( .D(n23238), .CK(clk), .Q(\mem[358][4] ) );
  DFF_X1 \mem_reg[358][3]  ( .D(n23239), .CK(clk), .Q(\mem[358][3] ) );
  DFF_X1 \mem_reg[358][2]  ( .D(n23240), .CK(clk), .Q(\mem[358][2] ) );
  DFF_X1 \mem_reg[358][1]  ( .D(n23241), .CK(clk), .Q(\mem[358][1] ) );
  DFF_X1 \mem_reg[358][0]  ( .D(n23242), .CK(clk), .Q(\mem[358][0] ) );
  DFF_X1 \mem_reg[357][7]  ( .D(n23243), .CK(clk), .Q(\mem[357][7] ) );
  DFF_X1 \mem_reg[357][6]  ( .D(n23244), .CK(clk), .Q(\mem[357][6] ) );
  DFF_X1 \mem_reg[357][5]  ( .D(n23245), .CK(clk), .Q(\mem[357][5] ) );
  DFF_X1 \mem_reg[357][4]  ( .D(n23246), .CK(clk), .Q(\mem[357][4] ) );
  DFF_X1 \mem_reg[357][3]  ( .D(n23247), .CK(clk), .Q(\mem[357][3] ) );
  DFF_X1 \mem_reg[357][2]  ( .D(n23248), .CK(clk), .Q(\mem[357][2] ) );
  DFF_X1 \mem_reg[357][1]  ( .D(n23249), .CK(clk), .Q(\mem[357][1] ) );
  DFF_X1 \mem_reg[357][0]  ( .D(n23250), .CK(clk), .Q(\mem[357][0] ) );
  DFF_X1 \mem_reg[356][7]  ( .D(n23251), .CK(clk), .Q(\mem[356][7] ) );
  DFF_X1 \mem_reg[356][6]  ( .D(n23252), .CK(clk), .Q(\mem[356][6] ) );
  DFF_X1 \mem_reg[356][5]  ( .D(n23253), .CK(clk), .Q(\mem[356][5] ) );
  DFF_X1 \mem_reg[356][4]  ( .D(n23254), .CK(clk), .Q(\mem[356][4] ) );
  DFF_X1 \mem_reg[356][3]  ( .D(n23255), .CK(clk), .Q(\mem[356][3] ) );
  DFF_X1 \mem_reg[356][2]  ( .D(n23256), .CK(clk), .Q(\mem[356][2] ) );
  DFF_X1 \mem_reg[356][1]  ( .D(n23257), .CK(clk), .Q(\mem[356][1] ) );
  DFF_X1 \mem_reg[356][0]  ( .D(n23258), .CK(clk), .Q(\mem[356][0] ) );
  DFF_X1 \mem_reg[355][7]  ( .D(n23259), .CK(clk), .Q(\mem[355][7] ) );
  DFF_X1 \mem_reg[355][6]  ( .D(n23260), .CK(clk), .Q(\mem[355][6] ) );
  DFF_X1 \mem_reg[355][5]  ( .D(n23261), .CK(clk), .Q(\mem[355][5] ) );
  DFF_X1 \mem_reg[355][4]  ( .D(n23262), .CK(clk), .Q(\mem[355][4] ) );
  DFF_X1 \mem_reg[355][3]  ( .D(n23263), .CK(clk), .Q(\mem[355][3] ) );
  DFF_X1 \mem_reg[355][2]  ( .D(n23264), .CK(clk), .Q(\mem[355][2] ) );
  DFF_X1 \mem_reg[355][1]  ( .D(n23265), .CK(clk), .Q(\mem[355][1] ) );
  DFF_X1 \mem_reg[355][0]  ( .D(n23266), .CK(clk), .Q(\mem[355][0] ) );
  DFF_X1 \mem_reg[354][7]  ( .D(n23267), .CK(clk), .Q(\mem[354][7] ) );
  DFF_X1 \mem_reg[354][6]  ( .D(n23268), .CK(clk), .Q(\mem[354][6] ) );
  DFF_X1 \mem_reg[354][5]  ( .D(n23269), .CK(clk), .Q(\mem[354][5] ) );
  DFF_X1 \mem_reg[354][4]  ( .D(n23270), .CK(clk), .Q(\mem[354][4] ) );
  DFF_X1 \mem_reg[354][3]  ( .D(n23271), .CK(clk), .Q(\mem[354][3] ) );
  DFF_X1 \mem_reg[354][2]  ( .D(n23272), .CK(clk), .Q(\mem[354][2] ) );
  DFF_X1 \mem_reg[354][1]  ( .D(n23273), .CK(clk), .Q(\mem[354][1] ) );
  DFF_X1 \mem_reg[354][0]  ( .D(n23274), .CK(clk), .Q(\mem[354][0] ) );
  DFF_X1 \mem_reg[353][7]  ( .D(n23275), .CK(clk), .Q(\mem[353][7] ) );
  DFF_X1 \mem_reg[353][6]  ( .D(n23276), .CK(clk), .Q(\mem[353][6] ) );
  DFF_X1 \mem_reg[353][5]  ( .D(n23277), .CK(clk), .Q(\mem[353][5] ) );
  DFF_X1 \mem_reg[353][4]  ( .D(n23278), .CK(clk), .Q(\mem[353][4] ) );
  DFF_X1 \mem_reg[353][3]  ( .D(n23279), .CK(clk), .Q(\mem[353][3] ) );
  DFF_X1 \mem_reg[353][2]  ( .D(n23280), .CK(clk), .Q(\mem[353][2] ) );
  DFF_X1 \mem_reg[353][1]  ( .D(n23281), .CK(clk), .Q(\mem[353][1] ) );
  DFF_X1 \mem_reg[353][0]  ( .D(n23282), .CK(clk), .Q(\mem[353][0] ) );
  DFF_X1 \mem_reg[352][7]  ( .D(n23283), .CK(clk), .Q(\mem[352][7] ) );
  DFF_X1 \mem_reg[352][6]  ( .D(n23284), .CK(clk), .Q(\mem[352][6] ) );
  DFF_X1 \mem_reg[352][5]  ( .D(n23285), .CK(clk), .Q(\mem[352][5] ) );
  DFF_X1 \mem_reg[352][4]  ( .D(n23286), .CK(clk), .Q(\mem[352][4] ) );
  DFF_X1 \mem_reg[352][3]  ( .D(n23287), .CK(clk), .Q(\mem[352][3] ) );
  DFF_X1 \mem_reg[352][2]  ( .D(n23288), .CK(clk), .Q(\mem[352][2] ) );
  DFF_X1 \mem_reg[352][1]  ( .D(n23289), .CK(clk), .Q(\mem[352][1] ) );
  DFF_X1 \mem_reg[352][0]  ( .D(n23290), .CK(clk), .Q(\mem[352][0] ) );
  DFF_X1 \mem_reg[351][7]  ( .D(n23291), .CK(clk), .Q(\mem[351][7] ) );
  DFF_X1 \mem_reg[351][6]  ( .D(n23292), .CK(clk), .Q(\mem[351][6] ) );
  DFF_X1 \mem_reg[351][5]  ( .D(n23293), .CK(clk), .Q(\mem[351][5] ) );
  DFF_X1 \mem_reg[351][4]  ( .D(n23294), .CK(clk), .Q(\mem[351][4] ) );
  DFF_X1 \mem_reg[351][3]  ( .D(n23295), .CK(clk), .Q(\mem[351][3] ) );
  DFF_X1 \mem_reg[351][2]  ( .D(n23296), .CK(clk), .Q(\mem[351][2] ) );
  DFF_X1 \mem_reg[351][1]  ( .D(n23297), .CK(clk), .Q(\mem[351][1] ) );
  DFF_X1 \mem_reg[351][0]  ( .D(n23298), .CK(clk), .Q(\mem[351][0] ) );
  DFF_X1 \mem_reg[350][7]  ( .D(n23299), .CK(clk), .Q(\mem[350][7] ) );
  DFF_X1 \mem_reg[350][6]  ( .D(n23300), .CK(clk), .Q(\mem[350][6] ) );
  DFF_X1 \mem_reg[350][5]  ( .D(n23301), .CK(clk), .Q(\mem[350][5] ) );
  DFF_X1 \mem_reg[350][4]  ( .D(n23302), .CK(clk), .Q(\mem[350][4] ) );
  DFF_X1 \mem_reg[350][3]  ( .D(n23303), .CK(clk), .Q(\mem[350][3] ) );
  DFF_X1 \mem_reg[350][2]  ( .D(n23304), .CK(clk), .Q(\mem[350][2] ) );
  DFF_X1 \mem_reg[350][1]  ( .D(n23305), .CK(clk), .Q(\mem[350][1] ) );
  DFF_X1 \mem_reg[350][0]  ( .D(n23306), .CK(clk), .Q(\mem[350][0] ) );
  DFF_X1 \mem_reg[349][7]  ( .D(n23307), .CK(clk), .Q(\mem[349][7] ) );
  DFF_X1 \mem_reg[349][6]  ( .D(n23308), .CK(clk), .Q(\mem[349][6] ) );
  DFF_X1 \mem_reg[349][5]  ( .D(n23309), .CK(clk), .Q(\mem[349][5] ) );
  DFF_X1 \mem_reg[349][4]  ( .D(n23310), .CK(clk), .Q(\mem[349][4] ) );
  DFF_X1 \mem_reg[349][3]  ( .D(n23311), .CK(clk), .Q(\mem[349][3] ) );
  DFF_X1 \mem_reg[349][2]  ( .D(n23312), .CK(clk), .Q(\mem[349][2] ) );
  DFF_X1 \mem_reg[349][1]  ( .D(n23313), .CK(clk), .Q(\mem[349][1] ) );
  DFF_X1 \mem_reg[349][0]  ( .D(n23314), .CK(clk), .Q(\mem[349][0] ) );
  DFF_X1 \mem_reg[348][7]  ( .D(n23315), .CK(clk), .Q(\mem[348][7] ) );
  DFF_X1 \mem_reg[348][6]  ( .D(n23316), .CK(clk), .Q(\mem[348][6] ) );
  DFF_X1 \mem_reg[348][5]  ( .D(n23317), .CK(clk), .Q(\mem[348][5] ) );
  DFF_X1 \mem_reg[348][4]  ( .D(n23318), .CK(clk), .Q(\mem[348][4] ) );
  DFF_X1 \mem_reg[348][3]  ( .D(n23319), .CK(clk), .Q(\mem[348][3] ) );
  DFF_X1 \mem_reg[348][2]  ( .D(n23320), .CK(clk), .Q(\mem[348][2] ) );
  DFF_X1 \mem_reg[348][1]  ( .D(n23321), .CK(clk), .Q(\mem[348][1] ) );
  DFF_X1 \mem_reg[348][0]  ( .D(n23322), .CK(clk), .Q(\mem[348][0] ) );
  DFF_X1 \mem_reg[347][7]  ( .D(n23323), .CK(clk), .Q(\mem[347][7] ) );
  DFF_X1 \mem_reg[347][6]  ( .D(n23324), .CK(clk), .Q(\mem[347][6] ) );
  DFF_X1 \mem_reg[347][5]  ( .D(n23325), .CK(clk), .Q(\mem[347][5] ) );
  DFF_X1 \mem_reg[347][4]  ( .D(n23326), .CK(clk), .Q(\mem[347][4] ) );
  DFF_X1 \mem_reg[347][3]  ( .D(n23327), .CK(clk), .Q(\mem[347][3] ) );
  DFF_X1 \mem_reg[347][2]  ( .D(n23328), .CK(clk), .Q(\mem[347][2] ) );
  DFF_X1 \mem_reg[347][1]  ( .D(n23329), .CK(clk), .Q(\mem[347][1] ) );
  DFF_X1 \mem_reg[347][0]  ( .D(n23330), .CK(clk), .Q(\mem[347][0] ) );
  DFF_X1 \mem_reg[346][7]  ( .D(n23331), .CK(clk), .Q(\mem[346][7] ) );
  DFF_X1 \mem_reg[346][6]  ( .D(n23332), .CK(clk), .Q(\mem[346][6] ) );
  DFF_X1 \mem_reg[346][5]  ( .D(n23333), .CK(clk), .Q(\mem[346][5] ) );
  DFF_X1 \mem_reg[346][4]  ( .D(n23334), .CK(clk), .Q(\mem[346][4] ) );
  DFF_X1 \mem_reg[346][3]  ( .D(n23335), .CK(clk), .Q(\mem[346][3] ) );
  DFF_X1 \mem_reg[346][2]  ( .D(n23336), .CK(clk), .Q(\mem[346][2] ) );
  DFF_X1 \mem_reg[346][1]  ( .D(n23337), .CK(clk), .Q(\mem[346][1] ) );
  DFF_X1 \mem_reg[346][0]  ( .D(n23338), .CK(clk), .Q(\mem[346][0] ) );
  DFF_X1 \mem_reg[345][7]  ( .D(n23339), .CK(clk), .Q(\mem[345][7] ) );
  DFF_X1 \mem_reg[345][6]  ( .D(n23340), .CK(clk), .Q(\mem[345][6] ) );
  DFF_X1 \mem_reg[345][5]  ( .D(n23341), .CK(clk), .Q(\mem[345][5] ) );
  DFF_X1 \mem_reg[345][4]  ( .D(n23342), .CK(clk), .Q(\mem[345][4] ) );
  DFF_X1 \mem_reg[345][3]  ( .D(n23343), .CK(clk), .Q(\mem[345][3] ) );
  DFF_X1 \mem_reg[345][2]  ( .D(n23344), .CK(clk), .Q(\mem[345][2] ) );
  DFF_X1 \mem_reg[345][1]  ( .D(n23345), .CK(clk), .Q(\mem[345][1] ) );
  DFF_X1 \mem_reg[345][0]  ( .D(n23346), .CK(clk), .Q(\mem[345][0] ) );
  DFF_X1 \mem_reg[344][7]  ( .D(n23347), .CK(clk), .Q(\mem[344][7] ) );
  DFF_X1 \mem_reg[344][6]  ( .D(n23348), .CK(clk), .Q(\mem[344][6] ) );
  DFF_X1 \mem_reg[344][5]  ( .D(n23349), .CK(clk), .Q(\mem[344][5] ) );
  DFF_X1 \mem_reg[344][4]  ( .D(n23350), .CK(clk), .Q(\mem[344][4] ) );
  DFF_X1 \mem_reg[344][3]  ( .D(n23351), .CK(clk), .Q(\mem[344][3] ) );
  DFF_X1 \mem_reg[344][2]  ( .D(n23352), .CK(clk), .Q(\mem[344][2] ) );
  DFF_X1 \mem_reg[344][1]  ( .D(n23353), .CK(clk), .Q(\mem[344][1] ) );
  DFF_X1 \mem_reg[344][0]  ( .D(n23354), .CK(clk), .Q(\mem[344][0] ) );
  DFF_X1 \mem_reg[343][7]  ( .D(n23355), .CK(clk), .Q(\mem[343][7] ) );
  DFF_X1 \mem_reg[343][6]  ( .D(n23356), .CK(clk), .Q(\mem[343][6] ) );
  DFF_X1 \mem_reg[343][5]  ( .D(n23357), .CK(clk), .Q(\mem[343][5] ) );
  DFF_X1 \mem_reg[343][4]  ( .D(n23358), .CK(clk), .Q(\mem[343][4] ) );
  DFF_X1 \mem_reg[343][3]  ( .D(n23359), .CK(clk), .Q(\mem[343][3] ) );
  DFF_X1 \mem_reg[343][2]  ( .D(n23360), .CK(clk), .Q(\mem[343][2] ) );
  DFF_X1 \mem_reg[343][1]  ( .D(n23361), .CK(clk), .Q(\mem[343][1] ) );
  DFF_X1 \mem_reg[343][0]  ( .D(n23362), .CK(clk), .Q(\mem[343][0] ) );
  DFF_X1 \mem_reg[342][7]  ( .D(n23363), .CK(clk), .Q(\mem[342][7] ) );
  DFF_X1 \mem_reg[342][6]  ( .D(n23364), .CK(clk), .Q(\mem[342][6] ) );
  DFF_X1 \mem_reg[342][5]  ( .D(n23365), .CK(clk), .Q(\mem[342][5] ) );
  DFF_X1 \mem_reg[342][4]  ( .D(n23366), .CK(clk), .Q(\mem[342][4] ) );
  DFF_X1 \mem_reg[342][3]  ( .D(n23367), .CK(clk), .Q(\mem[342][3] ) );
  DFF_X1 \mem_reg[342][2]  ( .D(n23368), .CK(clk), .Q(\mem[342][2] ) );
  DFF_X1 \mem_reg[342][1]  ( .D(n23369), .CK(clk), .Q(\mem[342][1] ) );
  DFF_X1 \mem_reg[342][0]  ( .D(n23370), .CK(clk), .Q(\mem[342][0] ) );
  DFF_X1 \mem_reg[341][7]  ( .D(n23371), .CK(clk), .Q(\mem[341][7] ) );
  DFF_X1 \mem_reg[341][6]  ( .D(n23372), .CK(clk), .Q(\mem[341][6] ) );
  DFF_X1 \mem_reg[341][5]  ( .D(n23373), .CK(clk), .Q(\mem[341][5] ) );
  DFF_X1 \mem_reg[341][4]  ( .D(n23374), .CK(clk), .Q(\mem[341][4] ) );
  DFF_X1 \mem_reg[341][3]  ( .D(n23375), .CK(clk), .Q(\mem[341][3] ) );
  DFF_X1 \mem_reg[341][2]  ( .D(n23376), .CK(clk), .Q(\mem[341][2] ) );
  DFF_X1 \mem_reg[341][1]  ( .D(n23377), .CK(clk), .Q(\mem[341][1] ) );
  DFF_X1 \mem_reg[341][0]  ( .D(n23378), .CK(clk), .Q(\mem[341][0] ) );
  DFF_X1 \mem_reg[340][7]  ( .D(n23379), .CK(clk), .Q(\mem[340][7] ) );
  DFF_X1 \mem_reg[340][6]  ( .D(n23380), .CK(clk), .Q(\mem[340][6] ) );
  DFF_X1 \mem_reg[340][5]  ( .D(n23381), .CK(clk), .Q(\mem[340][5] ) );
  DFF_X1 \mem_reg[340][4]  ( .D(n23382), .CK(clk), .Q(\mem[340][4] ) );
  DFF_X1 \mem_reg[340][3]  ( .D(n23383), .CK(clk), .Q(\mem[340][3] ) );
  DFF_X1 \mem_reg[340][2]  ( .D(n23384), .CK(clk), .Q(\mem[340][2] ) );
  DFF_X1 \mem_reg[340][1]  ( .D(n23385), .CK(clk), .Q(\mem[340][1] ) );
  DFF_X1 \mem_reg[340][0]  ( .D(n23386), .CK(clk), .Q(\mem[340][0] ) );
  DFF_X1 \mem_reg[339][7]  ( .D(n23387), .CK(clk), .Q(\mem[339][7] ) );
  DFF_X1 \mem_reg[339][6]  ( .D(n23388), .CK(clk), .Q(\mem[339][6] ) );
  DFF_X1 \mem_reg[339][5]  ( .D(n23389), .CK(clk), .Q(\mem[339][5] ) );
  DFF_X1 \mem_reg[339][4]  ( .D(n23390), .CK(clk), .Q(\mem[339][4] ) );
  DFF_X1 \mem_reg[339][3]  ( .D(n23391), .CK(clk), .Q(\mem[339][3] ) );
  DFF_X1 \mem_reg[339][2]  ( .D(n23392), .CK(clk), .Q(\mem[339][2] ) );
  DFF_X1 \mem_reg[339][1]  ( .D(n23393), .CK(clk), .Q(\mem[339][1] ) );
  DFF_X1 \mem_reg[339][0]  ( .D(n23394), .CK(clk), .Q(\mem[339][0] ) );
  DFF_X1 \mem_reg[338][7]  ( .D(n23395), .CK(clk), .Q(\mem[338][7] ) );
  DFF_X1 \mem_reg[338][6]  ( .D(n23396), .CK(clk), .Q(\mem[338][6] ) );
  DFF_X1 \mem_reg[338][5]  ( .D(n23397), .CK(clk), .Q(\mem[338][5] ) );
  DFF_X1 \mem_reg[338][4]  ( .D(n23398), .CK(clk), .Q(\mem[338][4] ) );
  DFF_X1 \mem_reg[338][3]  ( .D(n23399), .CK(clk), .Q(\mem[338][3] ) );
  DFF_X1 \mem_reg[338][2]  ( .D(n23400), .CK(clk), .Q(\mem[338][2] ) );
  DFF_X1 \mem_reg[338][1]  ( .D(n23401), .CK(clk), .Q(\mem[338][1] ) );
  DFF_X1 \mem_reg[338][0]  ( .D(n23402), .CK(clk), .Q(\mem[338][0] ) );
  DFF_X1 \mem_reg[337][7]  ( .D(n23403), .CK(clk), .Q(\mem[337][7] ) );
  DFF_X1 \mem_reg[337][6]  ( .D(n23404), .CK(clk), .Q(\mem[337][6] ) );
  DFF_X1 \mem_reg[337][5]  ( .D(n23405), .CK(clk), .Q(\mem[337][5] ) );
  DFF_X1 \mem_reg[337][4]  ( .D(n23406), .CK(clk), .Q(\mem[337][4] ) );
  DFF_X1 \mem_reg[337][3]  ( .D(n23407), .CK(clk), .Q(\mem[337][3] ) );
  DFF_X1 \mem_reg[337][2]  ( .D(n23408), .CK(clk), .Q(\mem[337][2] ) );
  DFF_X1 \mem_reg[337][1]  ( .D(n23409), .CK(clk), .Q(\mem[337][1] ) );
  DFF_X1 \mem_reg[337][0]  ( .D(n23410), .CK(clk), .Q(\mem[337][0] ) );
  DFF_X1 \mem_reg[336][7]  ( .D(n23411), .CK(clk), .Q(\mem[336][7] ) );
  DFF_X1 \mem_reg[336][6]  ( .D(n23412), .CK(clk), .Q(\mem[336][6] ) );
  DFF_X1 \mem_reg[336][5]  ( .D(n23413), .CK(clk), .Q(\mem[336][5] ) );
  DFF_X1 \mem_reg[336][4]  ( .D(n23414), .CK(clk), .Q(\mem[336][4] ) );
  DFF_X1 \mem_reg[336][3]  ( .D(n23415), .CK(clk), .Q(\mem[336][3] ) );
  DFF_X1 \mem_reg[336][2]  ( .D(n23416), .CK(clk), .Q(\mem[336][2] ) );
  DFF_X1 \mem_reg[336][1]  ( .D(n23417), .CK(clk), .Q(\mem[336][1] ) );
  DFF_X1 \mem_reg[336][0]  ( .D(n23418), .CK(clk), .Q(\mem[336][0] ) );
  DFF_X1 \mem_reg[335][7]  ( .D(n23419), .CK(clk), .Q(\mem[335][7] ) );
  DFF_X1 \mem_reg[335][6]  ( .D(n23420), .CK(clk), .Q(\mem[335][6] ) );
  DFF_X1 \mem_reg[335][5]  ( .D(n23421), .CK(clk), .Q(\mem[335][5] ) );
  DFF_X1 \mem_reg[335][4]  ( .D(n23422), .CK(clk), .Q(\mem[335][4] ) );
  DFF_X1 \mem_reg[335][3]  ( .D(n23423), .CK(clk), .Q(\mem[335][3] ) );
  DFF_X1 \mem_reg[335][2]  ( .D(n23424), .CK(clk), .Q(\mem[335][2] ) );
  DFF_X1 \mem_reg[335][1]  ( .D(n23425), .CK(clk), .Q(\mem[335][1] ) );
  DFF_X1 \mem_reg[335][0]  ( .D(n23426), .CK(clk), .Q(\mem[335][0] ) );
  DFF_X1 \mem_reg[334][7]  ( .D(n23427), .CK(clk), .Q(\mem[334][7] ) );
  DFF_X1 \mem_reg[334][6]  ( .D(n23428), .CK(clk), .Q(\mem[334][6] ) );
  DFF_X1 \mem_reg[334][5]  ( .D(n23429), .CK(clk), .Q(\mem[334][5] ) );
  DFF_X1 \mem_reg[334][4]  ( .D(n23430), .CK(clk), .Q(\mem[334][4] ) );
  DFF_X1 \mem_reg[334][3]  ( .D(n23431), .CK(clk), .Q(\mem[334][3] ) );
  DFF_X1 \mem_reg[334][2]  ( .D(n23432), .CK(clk), .Q(\mem[334][2] ) );
  DFF_X1 \mem_reg[334][1]  ( .D(n23433), .CK(clk), .Q(\mem[334][1] ) );
  DFF_X1 \mem_reg[334][0]  ( .D(n23434), .CK(clk), .Q(\mem[334][0] ) );
  DFF_X1 \mem_reg[333][7]  ( .D(n23435), .CK(clk), .Q(\mem[333][7] ) );
  DFF_X1 \mem_reg[333][6]  ( .D(n23436), .CK(clk), .Q(\mem[333][6] ) );
  DFF_X1 \mem_reg[333][5]  ( .D(n23437), .CK(clk), .Q(\mem[333][5] ) );
  DFF_X1 \mem_reg[333][4]  ( .D(n23438), .CK(clk), .Q(\mem[333][4] ) );
  DFF_X1 \mem_reg[333][3]  ( .D(n23439), .CK(clk), .Q(\mem[333][3] ) );
  DFF_X1 \mem_reg[333][2]  ( .D(n23440), .CK(clk), .Q(\mem[333][2] ) );
  DFF_X1 \mem_reg[333][1]  ( .D(n23441), .CK(clk), .Q(\mem[333][1] ) );
  DFF_X1 \mem_reg[333][0]  ( .D(n23442), .CK(clk), .Q(\mem[333][0] ) );
  DFF_X1 \mem_reg[332][7]  ( .D(n23443), .CK(clk), .Q(\mem[332][7] ) );
  DFF_X1 \mem_reg[332][6]  ( .D(n23444), .CK(clk), .Q(\mem[332][6] ) );
  DFF_X1 \mem_reg[332][5]  ( .D(n23445), .CK(clk), .Q(\mem[332][5] ) );
  DFF_X1 \mem_reg[332][4]  ( .D(n23446), .CK(clk), .Q(\mem[332][4] ) );
  DFF_X1 \mem_reg[332][3]  ( .D(n23447), .CK(clk), .Q(\mem[332][3] ) );
  DFF_X1 \mem_reg[332][2]  ( .D(n23448), .CK(clk), .Q(\mem[332][2] ) );
  DFF_X1 \mem_reg[332][1]  ( .D(n23449), .CK(clk), .Q(\mem[332][1] ) );
  DFF_X1 \mem_reg[332][0]  ( .D(n23450), .CK(clk), .Q(\mem[332][0] ) );
  DFF_X1 \mem_reg[331][7]  ( .D(n23451), .CK(clk), .Q(\mem[331][7] ) );
  DFF_X1 \mem_reg[331][6]  ( .D(n23452), .CK(clk), .Q(\mem[331][6] ) );
  DFF_X1 \mem_reg[331][5]  ( .D(n23453), .CK(clk), .Q(\mem[331][5] ) );
  DFF_X1 \mem_reg[331][4]  ( .D(n23454), .CK(clk), .Q(\mem[331][4] ) );
  DFF_X1 \mem_reg[331][3]  ( .D(n23455), .CK(clk), .Q(\mem[331][3] ) );
  DFF_X1 \mem_reg[331][2]  ( .D(n23456), .CK(clk), .Q(\mem[331][2] ) );
  DFF_X1 \mem_reg[331][1]  ( .D(n23457), .CK(clk), .Q(\mem[331][1] ) );
  DFF_X1 \mem_reg[331][0]  ( .D(n23458), .CK(clk), .Q(\mem[331][0] ) );
  DFF_X1 \mem_reg[330][7]  ( .D(n23459), .CK(clk), .Q(\mem[330][7] ) );
  DFF_X1 \mem_reg[330][6]  ( .D(n23460), .CK(clk), .Q(\mem[330][6] ) );
  DFF_X1 \mem_reg[330][5]  ( .D(n23461), .CK(clk), .Q(\mem[330][5] ) );
  DFF_X1 \mem_reg[330][4]  ( .D(n23462), .CK(clk), .Q(\mem[330][4] ) );
  DFF_X1 \mem_reg[330][3]  ( .D(n23463), .CK(clk), .Q(\mem[330][3] ) );
  DFF_X1 \mem_reg[330][2]  ( .D(n23464), .CK(clk), .Q(\mem[330][2] ) );
  DFF_X1 \mem_reg[330][1]  ( .D(n23465), .CK(clk), .Q(\mem[330][1] ) );
  DFF_X1 \mem_reg[330][0]  ( .D(n23466), .CK(clk), .Q(\mem[330][0] ) );
  DFF_X1 \mem_reg[329][7]  ( .D(n23467), .CK(clk), .Q(\mem[329][7] ) );
  DFF_X1 \mem_reg[329][6]  ( .D(n23468), .CK(clk), .Q(\mem[329][6] ) );
  DFF_X1 \mem_reg[329][5]  ( .D(n23469), .CK(clk), .Q(\mem[329][5] ) );
  DFF_X1 \mem_reg[329][4]  ( .D(n23470), .CK(clk), .Q(\mem[329][4] ) );
  DFF_X1 \mem_reg[329][3]  ( .D(n23471), .CK(clk), .Q(\mem[329][3] ) );
  DFF_X1 \mem_reg[329][2]  ( .D(n23472), .CK(clk), .Q(\mem[329][2] ) );
  DFF_X1 \mem_reg[329][1]  ( .D(n23473), .CK(clk), .Q(\mem[329][1] ) );
  DFF_X1 \mem_reg[329][0]  ( .D(n23474), .CK(clk), .Q(\mem[329][0] ) );
  DFF_X1 \mem_reg[328][7]  ( .D(n23475), .CK(clk), .Q(\mem[328][7] ) );
  DFF_X1 \mem_reg[328][6]  ( .D(n23476), .CK(clk), .Q(\mem[328][6] ) );
  DFF_X1 \mem_reg[328][5]  ( .D(n23477), .CK(clk), .Q(\mem[328][5] ) );
  DFF_X1 \mem_reg[328][4]  ( .D(n23478), .CK(clk), .Q(\mem[328][4] ) );
  DFF_X1 \mem_reg[328][3]  ( .D(n23479), .CK(clk), .Q(\mem[328][3] ) );
  DFF_X1 \mem_reg[328][2]  ( .D(n23480), .CK(clk), .Q(\mem[328][2] ) );
  DFF_X1 \mem_reg[328][1]  ( .D(n23481), .CK(clk), .Q(\mem[328][1] ) );
  DFF_X1 \mem_reg[328][0]  ( .D(n23482), .CK(clk), .Q(\mem[328][0] ) );
  DFF_X1 \mem_reg[327][7]  ( .D(n23483), .CK(clk), .Q(\mem[327][7] ) );
  DFF_X1 \mem_reg[327][6]  ( .D(n23484), .CK(clk), .Q(\mem[327][6] ) );
  DFF_X1 \mem_reg[327][5]  ( .D(n23485), .CK(clk), .Q(\mem[327][5] ) );
  DFF_X1 \mem_reg[327][4]  ( .D(n23486), .CK(clk), .Q(\mem[327][4] ) );
  DFF_X1 \mem_reg[327][3]  ( .D(n23487), .CK(clk), .Q(\mem[327][3] ) );
  DFF_X1 \mem_reg[327][2]  ( .D(n23488), .CK(clk), .Q(\mem[327][2] ) );
  DFF_X1 \mem_reg[327][1]  ( .D(n23489), .CK(clk), .Q(\mem[327][1] ) );
  DFF_X1 \mem_reg[327][0]  ( .D(n23490), .CK(clk), .Q(\mem[327][0] ) );
  DFF_X1 \mem_reg[326][7]  ( .D(n23491), .CK(clk), .Q(\mem[326][7] ) );
  DFF_X1 \mem_reg[326][6]  ( .D(n23492), .CK(clk), .Q(\mem[326][6] ) );
  DFF_X1 \mem_reg[326][5]  ( .D(n23493), .CK(clk), .Q(\mem[326][5] ) );
  DFF_X1 \mem_reg[326][4]  ( .D(n23494), .CK(clk), .Q(\mem[326][4] ) );
  DFF_X1 \mem_reg[326][3]  ( .D(n23495), .CK(clk), .Q(\mem[326][3] ) );
  DFF_X1 \mem_reg[326][2]  ( .D(n23496), .CK(clk), .Q(\mem[326][2] ) );
  DFF_X1 \mem_reg[326][1]  ( .D(n23497), .CK(clk), .Q(\mem[326][1] ) );
  DFF_X1 \mem_reg[326][0]  ( .D(n23498), .CK(clk), .Q(\mem[326][0] ) );
  DFF_X1 \mem_reg[325][7]  ( .D(n23499), .CK(clk), .Q(\mem[325][7] ) );
  DFF_X1 \mem_reg[325][6]  ( .D(n23500), .CK(clk), .Q(\mem[325][6] ) );
  DFF_X1 \mem_reg[325][5]  ( .D(n23501), .CK(clk), .Q(\mem[325][5] ) );
  DFF_X1 \mem_reg[325][4]  ( .D(n23502), .CK(clk), .Q(\mem[325][4] ) );
  DFF_X1 \mem_reg[325][3]  ( .D(n23503), .CK(clk), .Q(\mem[325][3] ) );
  DFF_X1 \mem_reg[325][2]  ( .D(n23504), .CK(clk), .Q(\mem[325][2] ) );
  DFF_X1 \mem_reg[325][1]  ( .D(n23505), .CK(clk), .Q(\mem[325][1] ) );
  DFF_X1 \mem_reg[325][0]  ( .D(n23506), .CK(clk), .Q(\mem[325][0] ) );
  DFF_X1 \mem_reg[324][7]  ( .D(n23507), .CK(clk), .Q(\mem[324][7] ) );
  DFF_X1 \mem_reg[324][6]  ( .D(n23508), .CK(clk), .Q(\mem[324][6] ) );
  DFF_X1 \mem_reg[324][5]  ( .D(n23509), .CK(clk), .Q(\mem[324][5] ) );
  DFF_X1 \mem_reg[324][4]  ( .D(n23510), .CK(clk), .Q(\mem[324][4] ) );
  DFF_X1 \mem_reg[324][3]  ( .D(n23511), .CK(clk), .Q(\mem[324][3] ) );
  DFF_X1 \mem_reg[324][2]  ( .D(n23512), .CK(clk), .Q(\mem[324][2] ) );
  DFF_X1 \mem_reg[324][1]  ( .D(n23513), .CK(clk), .Q(\mem[324][1] ) );
  DFF_X1 \mem_reg[324][0]  ( .D(n23514), .CK(clk), .Q(\mem[324][0] ) );
  DFF_X1 \mem_reg[323][7]  ( .D(n23515), .CK(clk), .Q(\mem[323][7] ) );
  DFF_X1 \mem_reg[323][6]  ( .D(n23516), .CK(clk), .Q(\mem[323][6] ) );
  DFF_X1 \mem_reg[323][5]  ( .D(n23517), .CK(clk), .Q(\mem[323][5] ) );
  DFF_X1 \mem_reg[323][4]  ( .D(n23518), .CK(clk), .Q(\mem[323][4] ) );
  DFF_X1 \mem_reg[323][3]  ( .D(n23519), .CK(clk), .Q(\mem[323][3] ) );
  DFF_X1 \mem_reg[323][2]  ( .D(n23520), .CK(clk), .Q(\mem[323][2] ) );
  DFF_X1 \mem_reg[323][1]  ( .D(n23521), .CK(clk), .Q(\mem[323][1] ) );
  DFF_X1 \mem_reg[323][0]  ( .D(n23522), .CK(clk), .Q(\mem[323][0] ) );
  DFF_X1 \mem_reg[322][7]  ( .D(n23523), .CK(clk), .Q(\mem[322][7] ) );
  DFF_X1 \mem_reg[322][6]  ( .D(n23524), .CK(clk), .Q(\mem[322][6] ) );
  DFF_X1 \mem_reg[322][5]  ( .D(n23525), .CK(clk), .Q(\mem[322][5] ) );
  DFF_X1 \mem_reg[322][4]  ( .D(n23526), .CK(clk), .Q(\mem[322][4] ) );
  DFF_X1 \mem_reg[322][3]  ( .D(n23527), .CK(clk), .Q(\mem[322][3] ) );
  DFF_X1 \mem_reg[322][2]  ( .D(n23528), .CK(clk), .Q(\mem[322][2] ) );
  DFF_X1 \mem_reg[322][1]  ( .D(n23529), .CK(clk), .Q(\mem[322][1] ) );
  DFF_X1 \mem_reg[322][0]  ( .D(n23530), .CK(clk), .Q(\mem[322][0] ) );
  DFF_X1 \mem_reg[321][7]  ( .D(n23531), .CK(clk), .Q(\mem[321][7] ) );
  DFF_X1 \mem_reg[321][6]  ( .D(n23532), .CK(clk), .Q(\mem[321][6] ) );
  DFF_X1 \mem_reg[321][5]  ( .D(n23533), .CK(clk), .Q(\mem[321][5] ) );
  DFF_X1 \mem_reg[321][4]  ( .D(n23534), .CK(clk), .Q(\mem[321][4] ) );
  DFF_X1 \mem_reg[321][3]  ( .D(n23535), .CK(clk), .Q(\mem[321][3] ) );
  DFF_X1 \mem_reg[321][2]  ( .D(n23536), .CK(clk), .Q(\mem[321][2] ) );
  DFF_X1 \mem_reg[321][1]  ( .D(n23537), .CK(clk), .Q(\mem[321][1] ) );
  DFF_X1 \mem_reg[321][0]  ( .D(n23538), .CK(clk), .Q(\mem[321][0] ) );
  DFF_X1 \mem_reg[320][7]  ( .D(n23539), .CK(clk), .Q(\mem[320][7] ) );
  DFF_X1 \mem_reg[320][6]  ( .D(n23540), .CK(clk), .Q(\mem[320][6] ) );
  DFF_X1 \mem_reg[320][5]  ( .D(n23541), .CK(clk), .Q(\mem[320][5] ) );
  DFF_X1 \mem_reg[320][4]  ( .D(n23542), .CK(clk), .Q(\mem[320][4] ) );
  DFF_X1 \mem_reg[320][3]  ( .D(n23543), .CK(clk), .Q(\mem[320][3] ) );
  DFF_X1 \mem_reg[320][2]  ( .D(n23544), .CK(clk), .Q(\mem[320][2] ) );
  DFF_X1 \mem_reg[320][1]  ( .D(n23545), .CK(clk), .Q(\mem[320][1] ) );
  DFF_X1 \mem_reg[320][0]  ( .D(n23546), .CK(clk), .Q(\mem[320][0] ) );
  DFF_X1 \mem_reg[319][7]  ( .D(n23547), .CK(clk), .Q(\mem[319][7] ) );
  DFF_X1 \mem_reg[319][6]  ( .D(n23548), .CK(clk), .Q(\mem[319][6] ) );
  DFF_X1 \mem_reg[319][5]  ( .D(n23549), .CK(clk), .Q(\mem[319][5] ) );
  DFF_X1 \mem_reg[319][4]  ( .D(n23550), .CK(clk), .Q(\mem[319][4] ) );
  DFF_X1 \mem_reg[319][3]  ( .D(n23551), .CK(clk), .Q(\mem[319][3] ) );
  DFF_X1 \mem_reg[319][2]  ( .D(n23552), .CK(clk), .Q(\mem[319][2] ) );
  DFF_X1 \mem_reg[319][1]  ( .D(n23553), .CK(clk), .Q(\mem[319][1] ) );
  DFF_X1 \mem_reg[319][0]  ( .D(n23554), .CK(clk), .Q(\mem[319][0] ) );
  DFF_X1 \mem_reg[318][7]  ( .D(n23555), .CK(clk), .Q(\mem[318][7] ) );
  DFF_X1 \mem_reg[318][6]  ( .D(n23556), .CK(clk), .Q(\mem[318][6] ) );
  DFF_X1 \mem_reg[318][5]  ( .D(n23557), .CK(clk), .Q(\mem[318][5] ) );
  DFF_X1 \mem_reg[318][4]  ( .D(n23558), .CK(clk), .Q(\mem[318][4] ) );
  DFF_X1 \mem_reg[318][3]  ( .D(n23559), .CK(clk), .Q(\mem[318][3] ) );
  DFF_X1 \mem_reg[318][2]  ( .D(n23560), .CK(clk), .Q(\mem[318][2] ) );
  DFF_X1 \mem_reg[318][1]  ( .D(n23561), .CK(clk), .Q(\mem[318][1] ) );
  DFF_X1 \mem_reg[318][0]  ( .D(n23562), .CK(clk), .Q(\mem[318][0] ) );
  DFF_X1 \mem_reg[317][7]  ( .D(n23563), .CK(clk), .Q(\mem[317][7] ) );
  DFF_X1 \mem_reg[317][6]  ( .D(n23564), .CK(clk), .Q(\mem[317][6] ) );
  DFF_X1 \mem_reg[317][5]  ( .D(n23565), .CK(clk), .Q(\mem[317][5] ) );
  DFF_X1 \mem_reg[317][4]  ( .D(n23566), .CK(clk), .Q(\mem[317][4] ) );
  DFF_X1 \mem_reg[317][3]  ( .D(n23567), .CK(clk), .Q(\mem[317][3] ) );
  DFF_X1 \mem_reg[317][2]  ( .D(n23568), .CK(clk), .Q(\mem[317][2] ) );
  DFF_X1 \mem_reg[317][1]  ( .D(n23569), .CK(clk), .Q(\mem[317][1] ) );
  DFF_X1 \mem_reg[317][0]  ( .D(n23570), .CK(clk), .Q(\mem[317][0] ) );
  DFF_X1 \mem_reg[316][7]  ( .D(n23571), .CK(clk), .Q(\mem[316][7] ) );
  DFF_X1 \mem_reg[316][6]  ( .D(n23572), .CK(clk), .Q(\mem[316][6] ) );
  DFF_X1 \mem_reg[316][5]  ( .D(n23573), .CK(clk), .Q(\mem[316][5] ) );
  DFF_X1 \mem_reg[316][4]  ( .D(n23574), .CK(clk), .Q(\mem[316][4] ) );
  DFF_X1 \mem_reg[316][3]  ( .D(n23575), .CK(clk), .Q(\mem[316][3] ) );
  DFF_X1 \mem_reg[316][2]  ( .D(n23576), .CK(clk), .Q(\mem[316][2] ) );
  DFF_X1 \mem_reg[316][1]  ( .D(n23577), .CK(clk), .Q(\mem[316][1] ) );
  DFF_X1 \mem_reg[316][0]  ( .D(n23578), .CK(clk), .Q(\mem[316][0] ) );
  DFF_X1 \mem_reg[315][7]  ( .D(n23579), .CK(clk), .Q(\mem[315][7] ) );
  DFF_X1 \mem_reg[315][6]  ( .D(n23580), .CK(clk), .Q(\mem[315][6] ) );
  DFF_X1 \mem_reg[315][5]  ( .D(n23581), .CK(clk), .Q(\mem[315][5] ) );
  DFF_X1 \mem_reg[315][4]  ( .D(n23582), .CK(clk), .Q(\mem[315][4] ) );
  DFF_X1 \mem_reg[315][3]  ( .D(n23583), .CK(clk), .Q(\mem[315][3] ) );
  DFF_X1 \mem_reg[315][2]  ( .D(n23584), .CK(clk), .Q(\mem[315][2] ) );
  DFF_X1 \mem_reg[315][1]  ( .D(n23585), .CK(clk), .Q(\mem[315][1] ) );
  DFF_X1 \mem_reg[315][0]  ( .D(n23586), .CK(clk), .Q(\mem[315][0] ) );
  DFF_X1 \mem_reg[314][7]  ( .D(n23587), .CK(clk), .Q(\mem[314][7] ) );
  DFF_X1 \mem_reg[314][6]  ( .D(n23588), .CK(clk), .Q(\mem[314][6] ) );
  DFF_X1 \mem_reg[314][5]  ( .D(n23589), .CK(clk), .Q(\mem[314][5] ) );
  DFF_X1 \mem_reg[314][4]  ( .D(n23590), .CK(clk), .Q(\mem[314][4] ) );
  DFF_X1 \mem_reg[314][3]  ( .D(n23591), .CK(clk), .Q(\mem[314][3] ) );
  DFF_X1 \mem_reg[314][2]  ( .D(n23592), .CK(clk), .Q(\mem[314][2] ) );
  DFF_X1 \mem_reg[314][1]  ( .D(n23593), .CK(clk), .Q(\mem[314][1] ) );
  DFF_X1 \mem_reg[314][0]  ( .D(n23594), .CK(clk), .Q(\mem[314][0] ) );
  DFF_X1 \mem_reg[313][7]  ( .D(n23595), .CK(clk), .Q(\mem[313][7] ) );
  DFF_X1 \mem_reg[313][6]  ( .D(n23596), .CK(clk), .Q(\mem[313][6] ) );
  DFF_X1 \mem_reg[313][5]  ( .D(n23597), .CK(clk), .Q(\mem[313][5] ) );
  DFF_X1 \mem_reg[313][4]  ( .D(n23598), .CK(clk), .Q(\mem[313][4] ) );
  DFF_X1 \mem_reg[313][3]  ( .D(n23599), .CK(clk), .Q(\mem[313][3] ) );
  DFF_X1 \mem_reg[313][2]  ( .D(n23600), .CK(clk), .Q(\mem[313][2] ) );
  DFF_X1 \mem_reg[313][1]  ( .D(n23601), .CK(clk), .Q(\mem[313][1] ) );
  DFF_X1 \mem_reg[313][0]  ( .D(n23602), .CK(clk), .Q(\mem[313][0] ) );
  DFF_X1 \mem_reg[312][7]  ( .D(n23603), .CK(clk), .Q(\mem[312][7] ) );
  DFF_X1 \mem_reg[312][6]  ( .D(n23604), .CK(clk), .Q(\mem[312][6] ) );
  DFF_X1 \mem_reg[312][5]  ( .D(n23605), .CK(clk), .Q(\mem[312][5] ) );
  DFF_X1 \mem_reg[312][4]  ( .D(n23606), .CK(clk), .Q(\mem[312][4] ) );
  DFF_X1 \mem_reg[312][3]  ( .D(n23607), .CK(clk), .Q(\mem[312][3] ) );
  DFF_X1 \mem_reg[312][2]  ( .D(n23608), .CK(clk), .Q(\mem[312][2] ) );
  DFF_X1 \mem_reg[312][1]  ( .D(n23609), .CK(clk), .Q(\mem[312][1] ) );
  DFF_X1 \mem_reg[312][0]  ( .D(n23610), .CK(clk), .Q(\mem[312][0] ) );
  DFF_X1 \mem_reg[311][7]  ( .D(n23611), .CK(clk), .Q(\mem[311][7] ) );
  DFF_X1 \mem_reg[311][6]  ( .D(n23612), .CK(clk), .Q(\mem[311][6] ) );
  DFF_X1 \mem_reg[311][5]  ( .D(n23613), .CK(clk), .Q(\mem[311][5] ) );
  DFF_X1 \mem_reg[311][4]  ( .D(n23614), .CK(clk), .Q(\mem[311][4] ) );
  DFF_X1 \mem_reg[311][3]  ( .D(n23615), .CK(clk), .Q(\mem[311][3] ) );
  DFF_X1 \mem_reg[311][2]  ( .D(n23616), .CK(clk), .Q(\mem[311][2] ) );
  DFF_X1 \mem_reg[311][1]  ( .D(n23617), .CK(clk), .Q(\mem[311][1] ) );
  DFF_X1 \mem_reg[311][0]  ( .D(n23618), .CK(clk), .Q(\mem[311][0] ) );
  DFF_X1 \mem_reg[310][7]  ( .D(n23619), .CK(clk), .Q(\mem[310][7] ) );
  DFF_X1 \mem_reg[310][6]  ( .D(n23620), .CK(clk), .Q(\mem[310][6] ) );
  DFF_X1 \mem_reg[310][5]  ( .D(n23621), .CK(clk), .Q(\mem[310][5] ) );
  DFF_X1 \mem_reg[310][4]  ( .D(n23622), .CK(clk), .Q(\mem[310][4] ) );
  DFF_X1 \mem_reg[310][3]  ( .D(n23623), .CK(clk), .Q(\mem[310][3] ) );
  DFF_X1 \mem_reg[310][2]  ( .D(n23624), .CK(clk), .Q(\mem[310][2] ) );
  DFF_X1 \mem_reg[310][1]  ( .D(n23625), .CK(clk), .Q(\mem[310][1] ) );
  DFF_X1 \mem_reg[310][0]  ( .D(n23626), .CK(clk), .Q(\mem[310][0] ) );
  DFF_X1 \mem_reg[309][7]  ( .D(n23627), .CK(clk), .Q(\mem[309][7] ) );
  DFF_X1 \mem_reg[309][6]  ( .D(n23628), .CK(clk), .Q(\mem[309][6] ) );
  DFF_X1 \mem_reg[309][5]  ( .D(n23629), .CK(clk), .Q(\mem[309][5] ) );
  DFF_X1 \mem_reg[309][4]  ( .D(n23630), .CK(clk), .Q(\mem[309][4] ) );
  DFF_X1 \mem_reg[309][3]  ( .D(n23631), .CK(clk), .Q(\mem[309][3] ) );
  DFF_X1 \mem_reg[309][2]  ( .D(n23632), .CK(clk), .Q(\mem[309][2] ) );
  DFF_X1 \mem_reg[309][1]  ( .D(n23633), .CK(clk), .Q(\mem[309][1] ) );
  DFF_X1 \mem_reg[309][0]  ( .D(n23634), .CK(clk), .Q(\mem[309][0] ) );
  DFF_X1 \mem_reg[308][7]  ( .D(n23635), .CK(clk), .Q(\mem[308][7] ) );
  DFF_X1 \mem_reg[308][6]  ( .D(n23636), .CK(clk), .Q(\mem[308][6] ) );
  DFF_X1 \mem_reg[308][5]  ( .D(n23637), .CK(clk), .Q(\mem[308][5] ) );
  DFF_X1 \mem_reg[308][4]  ( .D(n23638), .CK(clk), .Q(\mem[308][4] ) );
  DFF_X1 \mem_reg[308][3]  ( .D(n23639), .CK(clk), .Q(\mem[308][3] ) );
  DFF_X1 \mem_reg[308][2]  ( .D(n23640), .CK(clk), .Q(\mem[308][2] ) );
  DFF_X1 \mem_reg[308][1]  ( .D(n23641), .CK(clk), .Q(\mem[308][1] ) );
  DFF_X1 \mem_reg[308][0]  ( .D(n23642), .CK(clk), .Q(\mem[308][0] ) );
  DFF_X1 \mem_reg[307][7]  ( .D(n23643), .CK(clk), .Q(\mem[307][7] ) );
  DFF_X1 \mem_reg[307][6]  ( .D(n23644), .CK(clk), .Q(\mem[307][6] ) );
  DFF_X1 \mem_reg[307][5]  ( .D(n23645), .CK(clk), .Q(\mem[307][5] ) );
  DFF_X1 \mem_reg[307][4]  ( .D(n23646), .CK(clk), .Q(\mem[307][4] ) );
  DFF_X1 \mem_reg[307][3]  ( .D(n23647), .CK(clk), .Q(\mem[307][3] ) );
  DFF_X1 \mem_reg[307][2]  ( .D(n23648), .CK(clk), .Q(\mem[307][2] ) );
  DFF_X1 \mem_reg[307][1]  ( .D(n23649), .CK(clk), .Q(\mem[307][1] ) );
  DFF_X1 \mem_reg[307][0]  ( .D(n23650), .CK(clk), .Q(\mem[307][0] ) );
  DFF_X1 \mem_reg[306][7]  ( .D(n23651), .CK(clk), .Q(\mem[306][7] ) );
  DFF_X1 \mem_reg[306][6]  ( .D(n23652), .CK(clk), .Q(\mem[306][6] ) );
  DFF_X1 \mem_reg[306][5]  ( .D(n23653), .CK(clk), .Q(\mem[306][5] ) );
  DFF_X1 \mem_reg[306][4]  ( .D(n23654), .CK(clk), .Q(\mem[306][4] ) );
  DFF_X1 \mem_reg[306][3]  ( .D(n23655), .CK(clk), .Q(\mem[306][3] ) );
  DFF_X1 \mem_reg[306][2]  ( .D(n23656), .CK(clk), .Q(\mem[306][2] ) );
  DFF_X1 \mem_reg[306][1]  ( .D(n23657), .CK(clk), .Q(\mem[306][1] ) );
  DFF_X1 \mem_reg[306][0]  ( .D(n23658), .CK(clk), .Q(\mem[306][0] ) );
  DFF_X1 \mem_reg[305][7]  ( .D(n23659), .CK(clk), .Q(\mem[305][7] ) );
  DFF_X1 \mem_reg[305][6]  ( .D(n23660), .CK(clk), .Q(\mem[305][6] ) );
  DFF_X1 \mem_reg[305][5]  ( .D(n23661), .CK(clk), .Q(\mem[305][5] ) );
  DFF_X1 \mem_reg[305][4]  ( .D(n23662), .CK(clk), .Q(\mem[305][4] ) );
  DFF_X1 \mem_reg[305][3]  ( .D(n23663), .CK(clk), .Q(\mem[305][3] ) );
  DFF_X1 \mem_reg[305][2]  ( .D(n23664), .CK(clk), .Q(\mem[305][2] ) );
  DFF_X1 \mem_reg[305][1]  ( .D(n23665), .CK(clk), .Q(\mem[305][1] ) );
  DFF_X1 \mem_reg[305][0]  ( .D(n23666), .CK(clk), .Q(\mem[305][0] ) );
  DFF_X1 \mem_reg[304][7]  ( .D(n23667), .CK(clk), .Q(\mem[304][7] ) );
  DFF_X1 \mem_reg[304][6]  ( .D(n23668), .CK(clk), .Q(\mem[304][6] ) );
  DFF_X1 \mem_reg[304][5]  ( .D(n23669), .CK(clk), .Q(\mem[304][5] ) );
  DFF_X1 \mem_reg[304][4]  ( .D(n23670), .CK(clk), .Q(\mem[304][4] ) );
  DFF_X1 \mem_reg[304][3]  ( .D(n23671), .CK(clk), .Q(\mem[304][3] ) );
  DFF_X1 \mem_reg[304][2]  ( .D(n23672), .CK(clk), .Q(\mem[304][2] ) );
  DFF_X1 \mem_reg[304][1]  ( .D(n23673), .CK(clk), .Q(\mem[304][1] ) );
  DFF_X1 \mem_reg[304][0]  ( .D(n23674), .CK(clk), .Q(\mem[304][0] ) );
  DFF_X1 \mem_reg[303][7]  ( .D(n23675), .CK(clk), .Q(\mem[303][7] ) );
  DFF_X1 \mem_reg[303][6]  ( .D(n23676), .CK(clk), .Q(\mem[303][6] ) );
  DFF_X1 \mem_reg[303][5]  ( .D(n23677), .CK(clk), .Q(\mem[303][5] ) );
  DFF_X1 \mem_reg[303][4]  ( .D(n23678), .CK(clk), .Q(\mem[303][4] ) );
  DFF_X1 \mem_reg[303][3]  ( .D(n23679), .CK(clk), .Q(\mem[303][3] ) );
  DFF_X1 \mem_reg[303][2]  ( .D(n23680), .CK(clk), .Q(\mem[303][2] ) );
  DFF_X1 \mem_reg[303][1]  ( .D(n23681), .CK(clk), .Q(\mem[303][1] ) );
  DFF_X1 \mem_reg[303][0]  ( .D(n23682), .CK(clk), .Q(\mem[303][0] ) );
  DFF_X1 \mem_reg[302][7]  ( .D(n23683), .CK(clk), .Q(\mem[302][7] ) );
  DFF_X1 \mem_reg[302][6]  ( .D(n23684), .CK(clk), .Q(\mem[302][6] ) );
  DFF_X1 \mem_reg[302][5]  ( .D(n23685), .CK(clk), .Q(\mem[302][5] ) );
  DFF_X1 \mem_reg[302][4]  ( .D(n23686), .CK(clk), .Q(\mem[302][4] ) );
  DFF_X1 \mem_reg[302][3]  ( .D(n23687), .CK(clk), .Q(\mem[302][3] ) );
  DFF_X1 \mem_reg[302][2]  ( .D(n23688), .CK(clk), .Q(\mem[302][2] ) );
  DFF_X1 \mem_reg[302][1]  ( .D(n23689), .CK(clk), .Q(\mem[302][1] ) );
  DFF_X1 \mem_reg[302][0]  ( .D(n23690), .CK(clk), .Q(\mem[302][0] ) );
  DFF_X1 \mem_reg[301][7]  ( .D(n23691), .CK(clk), .Q(\mem[301][7] ) );
  DFF_X1 \mem_reg[301][6]  ( .D(n23692), .CK(clk), .Q(\mem[301][6] ) );
  DFF_X1 \mem_reg[301][5]  ( .D(n23693), .CK(clk), .Q(\mem[301][5] ) );
  DFF_X1 \mem_reg[301][4]  ( .D(n23694), .CK(clk), .Q(\mem[301][4] ) );
  DFF_X1 \mem_reg[301][3]  ( .D(n23695), .CK(clk), .Q(\mem[301][3] ) );
  DFF_X1 \mem_reg[301][2]  ( .D(n23696), .CK(clk), .Q(\mem[301][2] ) );
  DFF_X1 \mem_reg[301][1]  ( .D(n23697), .CK(clk), .Q(\mem[301][1] ) );
  DFF_X1 \mem_reg[301][0]  ( .D(n23698), .CK(clk), .Q(\mem[301][0] ) );
  DFF_X1 \mem_reg[300][7]  ( .D(n23699), .CK(clk), .Q(\mem[300][7] ) );
  DFF_X1 \mem_reg[300][6]  ( .D(n23700), .CK(clk), .Q(\mem[300][6] ) );
  DFF_X1 \mem_reg[300][5]  ( .D(n23701), .CK(clk), .Q(\mem[300][5] ) );
  DFF_X1 \mem_reg[300][4]  ( .D(n23702), .CK(clk), .Q(\mem[300][4] ) );
  DFF_X1 \mem_reg[300][3]  ( .D(n23703), .CK(clk), .Q(\mem[300][3] ) );
  DFF_X1 \mem_reg[300][2]  ( .D(n23704), .CK(clk), .Q(\mem[300][2] ) );
  DFF_X1 \mem_reg[300][1]  ( .D(n23705), .CK(clk), .Q(\mem[300][1] ) );
  DFF_X1 \mem_reg[300][0]  ( .D(n23706), .CK(clk), .Q(\mem[300][0] ) );
  DFF_X1 \mem_reg[299][7]  ( .D(n23707), .CK(clk), .Q(\mem[299][7] ) );
  DFF_X1 \mem_reg[299][6]  ( .D(n23708), .CK(clk), .Q(\mem[299][6] ) );
  DFF_X1 \mem_reg[299][5]  ( .D(n23709), .CK(clk), .Q(\mem[299][5] ) );
  DFF_X1 \mem_reg[299][4]  ( .D(n23710), .CK(clk), .Q(\mem[299][4] ) );
  DFF_X1 \mem_reg[299][3]  ( .D(n23711), .CK(clk), .Q(\mem[299][3] ) );
  DFF_X1 \mem_reg[299][2]  ( .D(n23712), .CK(clk), .Q(\mem[299][2] ) );
  DFF_X1 \mem_reg[299][1]  ( .D(n23713), .CK(clk), .Q(\mem[299][1] ) );
  DFF_X1 \mem_reg[299][0]  ( .D(n23714), .CK(clk), .Q(\mem[299][0] ) );
  DFF_X1 \mem_reg[298][7]  ( .D(n23715), .CK(clk), .Q(\mem[298][7] ) );
  DFF_X1 \mem_reg[298][6]  ( .D(n23716), .CK(clk), .Q(\mem[298][6] ) );
  DFF_X1 \mem_reg[298][5]  ( .D(n23717), .CK(clk), .Q(\mem[298][5] ) );
  DFF_X1 \mem_reg[298][4]  ( .D(n23718), .CK(clk), .Q(\mem[298][4] ) );
  DFF_X1 \mem_reg[298][3]  ( .D(n23719), .CK(clk), .Q(\mem[298][3] ) );
  DFF_X1 \mem_reg[298][2]  ( .D(n23720), .CK(clk), .Q(\mem[298][2] ) );
  DFF_X1 \mem_reg[298][1]  ( .D(n23721), .CK(clk), .Q(\mem[298][1] ) );
  DFF_X1 \mem_reg[298][0]  ( .D(n23722), .CK(clk), .Q(\mem[298][0] ) );
  DFF_X1 \mem_reg[297][7]  ( .D(n23723), .CK(clk), .Q(\mem[297][7] ) );
  DFF_X1 \mem_reg[297][6]  ( .D(n23724), .CK(clk), .Q(\mem[297][6] ) );
  DFF_X1 \mem_reg[297][5]  ( .D(n23725), .CK(clk), .Q(\mem[297][5] ) );
  DFF_X1 \mem_reg[297][4]  ( .D(n23726), .CK(clk), .Q(\mem[297][4] ) );
  DFF_X1 \mem_reg[297][3]  ( .D(n23727), .CK(clk), .Q(\mem[297][3] ) );
  DFF_X1 \mem_reg[297][2]  ( .D(n23728), .CK(clk), .Q(\mem[297][2] ) );
  DFF_X1 \mem_reg[297][1]  ( .D(n23729), .CK(clk), .Q(\mem[297][1] ) );
  DFF_X1 \mem_reg[297][0]  ( .D(n23730), .CK(clk), .Q(\mem[297][0] ) );
  DFF_X1 \mem_reg[296][7]  ( .D(n23731), .CK(clk), .Q(\mem[296][7] ) );
  DFF_X1 \mem_reg[296][6]  ( .D(n23732), .CK(clk), .Q(\mem[296][6] ) );
  DFF_X1 \mem_reg[296][5]  ( .D(n23733), .CK(clk), .Q(\mem[296][5] ) );
  DFF_X1 \mem_reg[296][4]  ( .D(n23734), .CK(clk), .Q(\mem[296][4] ) );
  DFF_X1 \mem_reg[296][3]  ( .D(n23735), .CK(clk), .Q(\mem[296][3] ) );
  DFF_X1 \mem_reg[296][2]  ( .D(n23736), .CK(clk), .Q(\mem[296][2] ) );
  DFF_X1 \mem_reg[296][1]  ( .D(n23737), .CK(clk), .Q(\mem[296][1] ) );
  DFF_X1 \mem_reg[296][0]  ( .D(n23738), .CK(clk), .Q(\mem[296][0] ) );
  DFF_X1 \mem_reg[295][7]  ( .D(n23739), .CK(clk), .Q(\mem[295][7] ) );
  DFF_X1 \mem_reg[295][6]  ( .D(n23740), .CK(clk), .Q(\mem[295][6] ) );
  DFF_X1 \mem_reg[295][5]  ( .D(n23741), .CK(clk), .Q(\mem[295][5] ) );
  DFF_X1 \mem_reg[295][4]  ( .D(n23742), .CK(clk), .Q(\mem[295][4] ) );
  DFF_X1 \mem_reg[295][3]  ( .D(n23743), .CK(clk), .Q(\mem[295][3] ) );
  DFF_X1 \mem_reg[295][2]  ( .D(n23744), .CK(clk), .Q(\mem[295][2] ) );
  DFF_X1 \mem_reg[295][1]  ( .D(n23745), .CK(clk), .Q(\mem[295][1] ) );
  DFF_X1 \mem_reg[295][0]  ( .D(n23746), .CK(clk), .Q(\mem[295][0] ) );
  DFF_X1 \mem_reg[294][7]  ( .D(n23747), .CK(clk), .Q(\mem[294][7] ) );
  DFF_X1 \mem_reg[294][6]  ( .D(n23748), .CK(clk), .Q(\mem[294][6] ) );
  DFF_X1 \mem_reg[294][5]  ( .D(n23749), .CK(clk), .Q(\mem[294][5] ) );
  DFF_X1 \mem_reg[294][4]  ( .D(n23750), .CK(clk), .Q(\mem[294][4] ) );
  DFF_X1 \mem_reg[294][3]  ( .D(n23751), .CK(clk), .Q(\mem[294][3] ) );
  DFF_X1 \mem_reg[294][2]  ( .D(n23752), .CK(clk), .Q(\mem[294][2] ) );
  DFF_X1 \mem_reg[294][1]  ( .D(n23753), .CK(clk), .Q(\mem[294][1] ) );
  DFF_X1 \mem_reg[294][0]  ( .D(n23754), .CK(clk), .Q(\mem[294][0] ) );
  DFF_X1 \mem_reg[293][7]  ( .D(n23755), .CK(clk), .Q(\mem[293][7] ) );
  DFF_X1 \mem_reg[293][6]  ( .D(n23756), .CK(clk), .Q(\mem[293][6] ) );
  DFF_X1 \mem_reg[293][5]  ( .D(n23757), .CK(clk), .Q(\mem[293][5] ) );
  DFF_X1 \mem_reg[293][4]  ( .D(n23758), .CK(clk), .Q(\mem[293][4] ) );
  DFF_X1 \mem_reg[293][3]  ( .D(n23759), .CK(clk), .Q(\mem[293][3] ) );
  DFF_X1 \mem_reg[293][2]  ( .D(n23760), .CK(clk), .Q(\mem[293][2] ) );
  DFF_X1 \mem_reg[293][1]  ( .D(n23761), .CK(clk), .Q(\mem[293][1] ) );
  DFF_X1 \mem_reg[293][0]  ( .D(n23762), .CK(clk), .Q(\mem[293][0] ) );
  DFF_X1 \mem_reg[292][7]  ( .D(n23763), .CK(clk), .Q(\mem[292][7] ) );
  DFF_X1 \mem_reg[292][6]  ( .D(n23764), .CK(clk), .Q(\mem[292][6] ) );
  DFF_X1 \mem_reg[292][5]  ( .D(n23765), .CK(clk), .Q(\mem[292][5] ) );
  DFF_X1 \mem_reg[292][4]  ( .D(n23766), .CK(clk), .Q(\mem[292][4] ) );
  DFF_X1 \mem_reg[292][3]  ( .D(n23767), .CK(clk), .Q(\mem[292][3] ) );
  DFF_X1 \mem_reg[292][2]  ( .D(n23768), .CK(clk), .Q(\mem[292][2] ) );
  DFF_X1 \mem_reg[292][1]  ( .D(n23769), .CK(clk), .Q(\mem[292][1] ) );
  DFF_X1 \mem_reg[292][0]  ( .D(n23770), .CK(clk), .Q(\mem[292][0] ) );
  DFF_X1 \mem_reg[291][7]  ( .D(n23771), .CK(clk), .Q(\mem[291][7] ) );
  DFF_X1 \mem_reg[291][6]  ( .D(n23772), .CK(clk), .Q(\mem[291][6] ) );
  DFF_X1 \mem_reg[291][5]  ( .D(n23773), .CK(clk), .Q(\mem[291][5] ) );
  DFF_X1 \mem_reg[291][4]  ( .D(n23774), .CK(clk), .Q(\mem[291][4] ) );
  DFF_X1 \mem_reg[291][3]  ( .D(n23775), .CK(clk), .Q(\mem[291][3] ) );
  DFF_X1 \mem_reg[291][2]  ( .D(n23776), .CK(clk), .Q(\mem[291][2] ) );
  DFF_X1 \mem_reg[291][1]  ( .D(n23777), .CK(clk), .Q(\mem[291][1] ) );
  DFF_X1 \mem_reg[291][0]  ( .D(n23778), .CK(clk), .Q(\mem[291][0] ) );
  DFF_X1 \mem_reg[290][7]  ( .D(n23779), .CK(clk), .Q(\mem[290][7] ) );
  DFF_X1 \mem_reg[290][6]  ( .D(n23780), .CK(clk), .Q(\mem[290][6] ) );
  DFF_X1 \mem_reg[290][5]  ( .D(n23781), .CK(clk), .Q(\mem[290][5] ) );
  DFF_X1 \mem_reg[290][4]  ( .D(n23782), .CK(clk), .Q(\mem[290][4] ) );
  DFF_X1 \mem_reg[290][3]  ( .D(n23783), .CK(clk), .Q(\mem[290][3] ) );
  DFF_X1 \mem_reg[290][2]  ( .D(n23784), .CK(clk), .Q(\mem[290][2] ) );
  DFF_X1 \mem_reg[290][1]  ( .D(n23785), .CK(clk), .Q(\mem[290][1] ) );
  DFF_X1 \mem_reg[290][0]  ( .D(n23786), .CK(clk), .Q(\mem[290][0] ) );
  DFF_X1 \mem_reg[289][7]  ( .D(n23787), .CK(clk), .Q(\mem[289][7] ) );
  DFF_X1 \mem_reg[289][6]  ( .D(n23788), .CK(clk), .Q(\mem[289][6] ) );
  DFF_X1 \mem_reg[289][5]  ( .D(n23789), .CK(clk), .Q(\mem[289][5] ) );
  DFF_X1 \mem_reg[289][4]  ( .D(n23790), .CK(clk), .Q(\mem[289][4] ) );
  DFF_X1 \mem_reg[289][3]  ( .D(n23791), .CK(clk), .Q(\mem[289][3] ) );
  DFF_X1 \mem_reg[289][2]  ( .D(n23792), .CK(clk), .Q(\mem[289][2] ) );
  DFF_X1 \mem_reg[289][1]  ( .D(n23793), .CK(clk), .Q(\mem[289][1] ) );
  DFF_X1 \mem_reg[289][0]  ( .D(n23794), .CK(clk), .Q(\mem[289][0] ) );
  DFF_X1 \mem_reg[288][7]  ( .D(n23795), .CK(clk), .Q(\mem[288][7] ) );
  DFF_X1 \mem_reg[288][6]  ( .D(n23796), .CK(clk), .Q(\mem[288][6] ) );
  DFF_X1 \mem_reg[288][5]  ( .D(n23797), .CK(clk), .Q(\mem[288][5] ) );
  DFF_X1 \mem_reg[288][4]  ( .D(n23798), .CK(clk), .Q(\mem[288][4] ) );
  DFF_X1 \mem_reg[288][3]  ( .D(n23799), .CK(clk), .Q(\mem[288][3] ) );
  DFF_X1 \mem_reg[288][2]  ( .D(n23800), .CK(clk), .Q(\mem[288][2] ) );
  DFF_X1 \mem_reg[288][1]  ( .D(n23801), .CK(clk), .Q(\mem[288][1] ) );
  DFF_X1 \mem_reg[288][0]  ( .D(n23802), .CK(clk), .Q(\mem[288][0] ) );
  DFF_X1 \mem_reg[287][7]  ( .D(n23803), .CK(clk), .Q(\mem[287][7] ) );
  DFF_X1 \mem_reg[287][6]  ( .D(n23804), .CK(clk), .Q(\mem[287][6] ) );
  DFF_X1 \mem_reg[287][5]  ( .D(n23805), .CK(clk), .Q(\mem[287][5] ) );
  DFF_X1 \mem_reg[287][4]  ( .D(n23806), .CK(clk), .Q(\mem[287][4] ) );
  DFF_X1 \mem_reg[287][3]  ( .D(n23807), .CK(clk), .Q(\mem[287][3] ) );
  DFF_X1 \mem_reg[287][2]  ( .D(n23808), .CK(clk), .Q(\mem[287][2] ) );
  DFF_X1 \mem_reg[287][1]  ( .D(n23809), .CK(clk), .Q(\mem[287][1] ) );
  DFF_X1 \mem_reg[287][0]  ( .D(n23810), .CK(clk), .Q(\mem[287][0] ) );
  DFF_X1 \mem_reg[286][7]  ( .D(n23811), .CK(clk), .Q(\mem[286][7] ) );
  DFF_X1 \mem_reg[286][6]  ( .D(n23812), .CK(clk), .Q(\mem[286][6] ) );
  DFF_X1 \mem_reg[286][5]  ( .D(n23813), .CK(clk), .Q(\mem[286][5] ) );
  DFF_X1 \mem_reg[286][4]  ( .D(n23814), .CK(clk), .Q(\mem[286][4] ) );
  DFF_X1 \mem_reg[286][3]  ( .D(n23815), .CK(clk), .Q(\mem[286][3] ) );
  DFF_X1 \mem_reg[286][2]  ( .D(n23816), .CK(clk), .Q(\mem[286][2] ) );
  DFF_X1 \mem_reg[286][1]  ( .D(n23817), .CK(clk), .Q(\mem[286][1] ) );
  DFF_X1 \mem_reg[286][0]  ( .D(n23818), .CK(clk), .Q(\mem[286][0] ) );
  DFF_X1 \mem_reg[285][7]  ( .D(n23819), .CK(clk), .Q(\mem[285][7] ) );
  DFF_X1 \mem_reg[285][6]  ( .D(n23820), .CK(clk), .Q(\mem[285][6] ) );
  DFF_X1 \mem_reg[285][5]  ( .D(n23821), .CK(clk), .Q(\mem[285][5] ) );
  DFF_X1 \mem_reg[285][4]  ( .D(n23822), .CK(clk), .Q(\mem[285][4] ) );
  DFF_X1 \mem_reg[285][3]  ( .D(n23823), .CK(clk), .Q(\mem[285][3] ) );
  DFF_X1 \mem_reg[285][2]  ( .D(n23824), .CK(clk), .Q(\mem[285][2] ) );
  DFF_X1 \mem_reg[285][1]  ( .D(n23825), .CK(clk), .Q(\mem[285][1] ) );
  DFF_X1 \mem_reg[285][0]  ( .D(n23826), .CK(clk), .Q(\mem[285][0] ) );
  DFF_X1 \mem_reg[284][7]  ( .D(n23827), .CK(clk), .Q(\mem[284][7] ) );
  DFF_X1 \mem_reg[284][6]  ( .D(n23828), .CK(clk), .Q(\mem[284][6] ) );
  DFF_X1 \mem_reg[284][5]  ( .D(n23829), .CK(clk), .Q(\mem[284][5] ) );
  DFF_X1 \mem_reg[284][4]  ( .D(n23830), .CK(clk), .Q(\mem[284][4] ) );
  DFF_X1 \mem_reg[284][3]  ( .D(n23831), .CK(clk), .Q(\mem[284][3] ) );
  DFF_X1 \mem_reg[284][2]  ( .D(n23832), .CK(clk), .Q(\mem[284][2] ) );
  DFF_X1 \mem_reg[284][1]  ( .D(n23833), .CK(clk), .Q(\mem[284][1] ) );
  DFF_X1 \mem_reg[284][0]  ( .D(n23834), .CK(clk), .Q(\mem[284][0] ) );
  DFF_X1 \mem_reg[283][7]  ( .D(n23835), .CK(clk), .Q(\mem[283][7] ) );
  DFF_X1 \mem_reg[283][6]  ( .D(n23836), .CK(clk), .Q(\mem[283][6] ) );
  DFF_X1 \mem_reg[283][5]  ( .D(n23837), .CK(clk), .Q(\mem[283][5] ) );
  DFF_X1 \mem_reg[283][4]  ( .D(n23838), .CK(clk), .Q(\mem[283][4] ) );
  DFF_X1 \mem_reg[283][3]  ( .D(n23839), .CK(clk), .Q(\mem[283][3] ) );
  DFF_X1 \mem_reg[283][2]  ( .D(n23840), .CK(clk), .Q(\mem[283][2] ) );
  DFF_X1 \mem_reg[283][1]  ( .D(n23841), .CK(clk), .Q(\mem[283][1] ) );
  DFF_X1 \mem_reg[283][0]  ( .D(n23842), .CK(clk), .Q(\mem[283][0] ) );
  DFF_X1 \mem_reg[282][7]  ( .D(n23843), .CK(clk), .Q(\mem[282][7] ) );
  DFF_X1 \mem_reg[282][6]  ( .D(n23844), .CK(clk), .Q(\mem[282][6] ) );
  DFF_X1 \mem_reg[282][5]  ( .D(n23845), .CK(clk), .Q(\mem[282][5] ) );
  DFF_X1 \mem_reg[282][4]  ( .D(n23846), .CK(clk), .Q(\mem[282][4] ) );
  DFF_X1 \mem_reg[282][3]  ( .D(n23847), .CK(clk), .Q(\mem[282][3] ) );
  DFF_X1 \mem_reg[282][2]  ( .D(n23848), .CK(clk), .Q(\mem[282][2] ) );
  DFF_X1 \mem_reg[282][1]  ( .D(n23849), .CK(clk), .Q(\mem[282][1] ) );
  DFF_X1 \mem_reg[282][0]  ( .D(n23850), .CK(clk), .Q(\mem[282][0] ) );
  DFF_X1 \mem_reg[281][7]  ( .D(n23851), .CK(clk), .Q(\mem[281][7] ) );
  DFF_X1 \mem_reg[281][6]  ( .D(n23852), .CK(clk), .Q(\mem[281][6] ) );
  DFF_X1 \mem_reg[281][5]  ( .D(n23853), .CK(clk), .Q(\mem[281][5] ) );
  DFF_X1 \mem_reg[281][4]  ( .D(n23854), .CK(clk), .Q(\mem[281][4] ) );
  DFF_X1 \mem_reg[281][3]  ( .D(n23855), .CK(clk), .Q(\mem[281][3] ) );
  DFF_X1 \mem_reg[281][2]  ( .D(n23856), .CK(clk), .Q(\mem[281][2] ) );
  DFF_X1 \mem_reg[281][1]  ( .D(n23857), .CK(clk), .Q(\mem[281][1] ) );
  DFF_X1 \mem_reg[281][0]  ( .D(n23858), .CK(clk), .Q(\mem[281][0] ) );
  DFF_X1 \mem_reg[280][7]  ( .D(n23859), .CK(clk), .Q(\mem[280][7] ) );
  DFF_X1 \mem_reg[280][6]  ( .D(n23860), .CK(clk), .Q(\mem[280][6] ) );
  DFF_X1 \mem_reg[280][5]  ( .D(n23861), .CK(clk), .Q(\mem[280][5] ) );
  DFF_X1 \mem_reg[280][4]  ( .D(n23862), .CK(clk), .Q(\mem[280][4] ) );
  DFF_X1 \mem_reg[280][3]  ( .D(n23863), .CK(clk), .Q(\mem[280][3] ) );
  DFF_X1 \mem_reg[280][2]  ( .D(n23864), .CK(clk), .Q(\mem[280][2] ) );
  DFF_X1 \mem_reg[280][1]  ( .D(n23865), .CK(clk), .Q(\mem[280][1] ) );
  DFF_X1 \mem_reg[280][0]  ( .D(n23866), .CK(clk), .Q(\mem[280][0] ) );
  DFF_X1 \mem_reg[279][7]  ( .D(n23867), .CK(clk), .Q(\mem[279][7] ) );
  DFF_X1 \mem_reg[279][6]  ( .D(n23868), .CK(clk), .Q(\mem[279][6] ) );
  DFF_X1 \mem_reg[279][5]  ( .D(n23869), .CK(clk), .Q(\mem[279][5] ) );
  DFF_X1 \mem_reg[279][4]  ( .D(n23870), .CK(clk), .Q(\mem[279][4] ) );
  DFF_X1 \mem_reg[279][3]  ( .D(n23871), .CK(clk), .Q(\mem[279][3] ) );
  DFF_X1 \mem_reg[279][2]  ( .D(n23872), .CK(clk), .Q(\mem[279][2] ) );
  DFF_X1 \mem_reg[279][1]  ( .D(n23873), .CK(clk), .Q(\mem[279][1] ) );
  DFF_X1 \mem_reg[279][0]  ( .D(n23874), .CK(clk), .Q(\mem[279][0] ) );
  DFF_X1 \mem_reg[278][7]  ( .D(n23875), .CK(clk), .Q(\mem[278][7] ) );
  DFF_X1 \mem_reg[278][6]  ( .D(n23876), .CK(clk), .Q(\mem[278][6] ) );
  DFF_X1 \mem_reg[278][5]  ( .D(n23877), .CK(clk), .Q(\mem[278][5] ) );
  DFF_X1 \mem_reg[278][4]  ( .D(n23878), .CK(clk), .Q(\mem[278][4] ) );
  DFF_X1 \mem_reg[278][3]  ( .D(n23879), .CK(clk), .Q(\mem[278][3] ) );
  DFF_X1 \mem_reg[278][2]  ( .D(n23880), .CK(clk), .Q(\mem[278][2] ) );
  DFF_X1 \mem_reg[278][1]  ( .D(n23881), .CK(clk), .Q(\mem[278][1] ) );
  DFF_X1 \mem_reg[278][0]  ( .D(n23882), .CK(clk), .Q(\mem[278][0] ) );
  DFF_X1 \mem_reg[277][7]  ( .D(n23883), .CK(clk), .Q(\mem[277][7] ) );
  DFF_X1 \mem_reg[277][6]  ( .D(n23884), .CK(clk), .Q(\mem[277][6] ) );
  DFF_X1 \mem_reg[277][5]  ( .D(n23885), .CK(clk), .Q(\mem[277][5] ) );
  DFF_X1 \mem_reg[277][4]  ( .D(n23886), .CK(clk), .Q(\mem[277][4] ) );
  DFF_X1 \mem_reg[277][3]  ( .D(n23887), .CK(clk), .Q(\mem[277][3] ) );
  DFF_X1 \mem_reg[277][2]  ( .D(n23888), .CK(clk), .Q(\mem[277][2] ) );
  DFF_X1 \mem_reg[277][1]  ( .D(n23889), .CK(clk), .Q(\mem[277][1] ) );
  DFF_X1 \mem_reg[277][0]  ( .D(n23890), .CK(clk), .Q(\mem[277][0] ) );
  DFF_X1 \mem_reg[276][7]  ( .D(n23891), .CK(clk), .Q(\mem[276][7] ) );
  DFF_X1 \mem_reg[276][6]  ( .D(n23892), .CK(clk), .Q(\mem[276][6] ) );
  DFF_X1 \mem_reg[276][5]  ( .D(n23893), .CK(clk), .Q(\mem[276][5] ) );
  DFF_X1 \mem_reg[276][4]  ( .D(n23894), .CK(clk), .Q(\mem[276][4] ) );
  DFF_X1 \mem_reg[276][3]  ( .D(n23895), .CK(clk), .Q(\mem[276][3] ) );
  DFF_X1 \mem_reg[276][2]  ( .D(n23896), .CK(clk), .Q(\mem[276][2] ) );
  DFF_X1 \mem_reg[276][1]  ( .D(n23897), .CK(clk), .Q(\mem[276][1] ) );
  DFF_X1 \mem_reg[276][0]  ( .D(n23898), .CK(clk), .Q(\mem[276][0] ) );
  DFF_X1 \mem_reg[275][7]  ( .D(n23899), .CK(clk), .Q(\mem[275][7] ) );
  DFF_X1 \mem_reg[275][6]  ( .D(n23900), .CK(clk), .Q(\mem[275][6] ) );
  DFF_X1 \mem_reg[275][5]  ( .D(n23901), .CK(clk), .Q(\mem[275][5] ) );
  DFF_X1 \mem_reg[275][4]  ( .D(n23902), .CK(clk), .Q(\mem[275][4] ) );
  DFF_X1 \mem_reg[275][3]  ( .D(n23903), .CK(clk), .Q(\mem[275][3] ) );
  DFF_X1 \mem_reg[275][2]  ( .D(n23904), .CK(clk), .Q(\mem[275][2] ) );
  DFF_X1 \mem_reg[275][1]  ( .D(n23905), .CK(clk), .Q(\mem[275][1] ) );
  DFF_X1 \mem_reg[275][0]  ( .D(n23906), .CK(clk), .Q(\mem[275][0] ) );
  DFF_X1 \mem_reg[274][7]  ( .D(n23907), .CK(clk), .Q(\mem[274][7] ) );
  DFF_X1 \mem_reg[274][6]  ( .D(n23908), .CK(clk), .Q(\mem[274][6] ) );
  DFF_X1 \mem_reg[274][5]  ( .D(n23909), .CK(clk), .Q(\mem[274][5] ) );
  DFF_X1 \mem_reg[274][4]  ( .D(n23910), .CK(clk), .Q(\mem[274][4] ) );
  DFF_X1 \mem_reg[274][3]  ( .D(n23911), .CK(clk), .Q(\mem[274][3] ) );
  DFF_X1 \mem_reg[274][2]  ( .D(n23912), .CK(clk), .Q(\mem[274][2] ) );
  DFF_X1 \mem_reg[274][1]  ( .D(n23913), .CK(clk), .Q(\mem[274][1] ) );
  DFF_X1 \mem_reg[274][0]  ( .D(n23914), .CK(clk), .Q(\mem[274][0] ) );
  DFF_X1 \mem_reg[273][7]  ( .D(n23915), .CK(clk), .Q(\mem[273][7] ) );
  DFF_X1 \mem_reg[273][6]  ( .D(n23916), .CK(clk), .Q(\mem[273][6] ) );
  DFF_X1 \mem_reg[273][5]  ( .D(n23917), .CK(clk), .Q(\mem[273][5] ) );
  DFF_X1 \mem_reg[273][4]  ( .D(n23918), .CK(clk), .Q(\mem[273][4] ) );
  DFF_X1 \mem_reg[273][3]  ( .D(n23919), .CK(clk), .Q(\mem[273][3] ) );
  DFF_X1 \mem_reg[273][2]  ( .D(n23920), .CK(clk), .Q(\mem[273][2] ) );
  DFF_X1 \mem_reg[273][1]  ( .D(n23921), .CK(clk), .Q(\mem[273][1] ) );
  DFF_X1 \mem_reg[273][0]  ( .D(n23922), .CK(clk), .Q(\mem[273][0] ) );
  DFF_X1 \mem_reg[272][7]  ( .D(n23923), .CK(clk), .Q(\mem[272][7] ) );
  DFF_X1 \mem_reg[272][6]  ( .D(n23924), .CK(clk), .Q(\mem[272][6] ) );
  DFF_X1 \mem_reg[272][5]  ( .D(n23925), .CK(clk), .Q(\mem[272][5] ) );
  DFF_X1 \mem_reg[272][4]  ( .D(n23926), .CK(clk), .Q(\mem[272][4] ) );
  DFF_X1 \mem_reg[272][3]  ( .D(n23927), .CK(clk), .Q(\mem[272][3] ) );
  DFF_X1 \mem_reg[272][2]  ( .D(n23928), .CK(clk), .Q(\mem[272][2] ) );
  DFF_X1 \mem_reg[272][1]  ( .D(n23929), .CK(clk), .Q(\mem[272][1] ) );
  DFF_X1 \mem_reg[272][0]  ( .D(n23930), .CK(clk), .Q(\mem[272][0] ) );
  DFF_X1 \mem_reg[271][7]  ( .D(n23931), .CK(clk), .Q(\mem[271][7] ) );
  DFF_X1 \mem_reg[271][6]  ( .D(n23932), .CK(clk), .Q(\mem[271][6] ) );
  DFF_X1 \mem_reg[271][5]  ( .D(n23933), .CK(clk), .Q(\mem[271][5] ) );
  DFF_X1 \mem_reg[271][4]  ( .D(n23934), .CK(clk), .Q(\mem[271][4] ) );
  DFF_X1 \mem_reg[271][3]  ( .D(n23935), .CK(clk), .Q(\mem[271][3] ) );
  DFF_X1 \mem_reg[271][2]  ( .D(n23936), .CK(clk), .Q(\mem[271][2] ) );
  DFF_X1 \mem_reg[271][1]  ( .D(n23937), .CK(clk), .Q(\mem[271][1] ) );
  DFF_X1 \mem_reg[271][0]  ( .D(n23938), .CK(clk), .Q(\mem[271][0] ) );
  DFF_X1 \mem_reg[270][7]  ( .D(n23939), .CK(clk), .Q(\mem[270][7] ) );
  DFF_X1 \mem_reg[270][6]  ( .D(n23940), .CK(clk), .Q(\mem[270][6] ) );
  DFF_X1 \mem_reg[270][5]  ( .D(n23941), .CK(clk), .Q(\mem[270][5] ) );
  DFF_X1 \mem_reg[270][4]  ( .D(n23942), .CK(clk), .Q(\mem[270][4] ) );
  DFF_X1 \mem_reg[270][3]  ( .D(n23943), .CK(clk), .Q(\mem[270][3] ) );
  DFF_X1 \mem_reg[270][2]  ( .D(n23944), .CK(clk), .Q(\mem[270][2] ) );
  DFF_X1 \mem_reg[270][1]  ( .D(n23945), .CK(clk), .Q(\mem[270][1] ) );
  DFF_X1 \mem_reg[270][0]  ( .D(n23946), .CK(clk), .Q(\mem[270][0] ) );
  DFF_X1 \mem_reg[269][7]  ( .D(n23947), .CK(clk), .Q(\mem[269][7] ) );
  DFF_X1 \mem_reg[269][6]  ( .D(n23948), .CK(clk), .Q(\mem[269][6] ) );
  DFF_X1 \mem_reg[269][5]  ( .D(n23949), .CK(clk), .Q(\mem[269][5] ) );
  DFF_X1 \mem_reg[269][4]  ( .D(n23950), .CK(clk), .Q(\mem[269][4] ) );
  DFF_X1 \mem_reg[269][3]  ( .D(n23951), .CK(clk), .Q(\mem[269][3] ) );
  DFF_X1 \mem_reg[269][2]  ( .D(n23952), .CK(clk), .Q(\mem[269][2] ) );
  DFF_X1 \mem_reg[269][1]  ( .D(n23953), .CK(clk), .Q(\mem[269][1] ) );
  DFF_X1 \mem_reg[269][0]  ( .D(n23954), .CK(clk), .Q(\mem[269][0] ) );
  DFF_X1 \mem_reg[268][7]  ( .D(n23955), .CK(clk), .Q(\mem[268][7] ) );
  DFF_X1 \mem_reg[268][6]  ( .D(n23956), .CK(clk), .Q(\mem[268][6] ) );
  DFF_X1 \mem_reg[268][5]  ( .D(n23957), .CK(clk), .Q(\mem[268][5] ) );
  DFF_X1 \mem_reg[268][4]  ( .D(n23958), .CK(clk), .Q(\mem[268][4] ) );
  DFF_X1 \mem_reg[268][3]  ( .D(n23959), .CK(clk), .Q(\mem[268][3] ) );
  DFF_X1 \mem_reg[268][2]  ( .D(n23960), .CK(clk), .Q(\mem[268][2] ) );
  DFF_X1 \mem_reg[268][1]  ( .D(n23961), .CK(clk), .Q(\mem[268][1] ) );
  DFF_X1 \mem_reg[268][0]  ( .D(n23962), .CK(clk), .Q(\mem[268][0] ) );
  DFF_X1 \mem_reg[267][7]  ( .D(n23963), .CK(clk), .Q(\mem[267][7] ) );
  DFF_X1 \mem_reg[267][6]  ( .D(n23964), .CK(clk), .Q(\mem[267][6] ) );
  DFF_X1 \mem_reg[267][5]  ( .D(n23965), .CK(clk), .Q(\mem[267][5] ) );
  DFF_X1 \mem_reg[267][4]  ( .D(n23966), .CK(clk), .Q(\mem[267][4] ) );
  DFF_X1 \mem_reg[267][3]  ( .D(n23967), .CK(clk), .Q(\mem[267][3] ) );
  DFF_X1 \mem_reg[267][2]  ( .D(n23968), .CK(clk), .Q(\mem[267][2] ) );
  DFF_X1 \mem_reg[267][1]  ( .D(n23969), .CK(clk), .Q(\mem[267][1] ) );
  DFF_X1 \mem_reg[267][0]  ( .D(n23970), .CK(clk), .Q(\mem[267][0] ) );
  DFF_X1 \mem_reg[266][7]  ( .D(n23971), .CK(clk), .Q(\mem[266][7] ) );
  DFF_X1 \mem_reg[266][6]  ( .D(n23972), .CK(clk), .Q(\mem[266][6] ) );
  DFF_X1 \mem_reg[266][5]  ( .D(n23973), .CK(clk), .Q(\mem[266][5] ) );
  DFF_X1 \mem_reg[266][4]  ( .D(n23974), .CK(clk), .Q(\mem[266][4] ) );
  DFF_X1 \mem_reg[266][3]  ( .D(n23975), .CK(clk), .Q(\mem[266][3] ) );
  DFF_X1 \mem_reg[266][2]  ( .D(n23976), .CK(clk), .Q(\mem[266][2] ) );
  DFF_X1 \mem_reg[266][1]  ( .D(n23977), .CK(clk), .Q(\mem[266][1] ) );
  DFF_X1 \mem_reg[266][0]  ( .D(n23978), .CK(clk), .Q(\mem[266][0] ) );
  DFF_X1 \mem_reg[265][7]  ( .D(n23979), .CK(clk), .Q(\mem[265][7] ) );
  DFF_X1 \mem_reg[265][6]  ( .D(n23980), .CK(clk), .Q(\mem[265][6] ) );
  DFF_X1 \mem_reg[265][5]  ( .D(n23981), .CK(clk), .Q(\mem[265][5] ) );
  DFF_X1 \mem_reg[265][4]  ( .D(n23982), .CK(clk), .Q(\mem[265][4] ) );
  DFF_X1 \mem_reg[265][3]  ( .D(n23983), .CK(clk), .Q(\mem[265][3] ) );
  DFF_X1 \mem_reg[265][2]  ( .D(n23984), .CK(clk), .Q(\mem[265][2] ) );
  DFF_X1 \mem_reg[265][1]  ( .D(n23985), .CK(clk), .Q(\mem[265][1] ) );
  DFF_X1 \mem_reg[265][0]  ( .D(n23986), .CK(clk), .Q(\mem[265][0] ) );
  DFF_X1 \mem_reg[264][7]  ( .D(n23987), .CK(clk), .Q(\mem[264][7] ) );
  DFF_X1 \mem_reg[264][6]  ( .D(n23988), .CK(clk), .Q(\mem[264][6] ) );
  DFF_X1 \mem_reg[264][5]  ( .D(n23989), .CK(clk), .Q(\mem[264][5] ) );
  DFF_X1 \mem_reg[264][4]  ( .D(n23990), .CK(clk), .Q(\mem[264][4] ) );
  DFF_X1 \mem_reg[264][3]  ( .D(n23991), .CK(clk), .Q(\mem[264][3] ) );
  DFF_X1 \mem_reg[264][2]  ( .D(n23992), .CK(clk), .Q(\mem[264][2] ) );
  DFF_X1 \mem_reg[264][1]  ( .D(n23993), .CK(clk), .Q(\mem[264][1] ) );
  DFF_X1 \mem_reg[264][0]  ( .D(n23994), .CK(clk), .Q(\mem[264][0] ) );
  DFF_X1 \mem_reg[263][7]  ( .D(n23995), .CK(clk), .Q(\mem[263][7] ) );
  DFF_X1 \mem_reg[263][6]  ( .D(n23996), .CK(clk), .Q(\mem[263][6] ) );
  DFF_X1 \mem_reg[263][5]  ( .D(n23997), .CK(clk), .Q(\mem[263][5] ) );
  DFF_X1 \mem_reg[263][4]  ( .D(n23998), .CK(clk), .Q(\mem[263][4] ) );
  DFF_X1 \mem_reg[263][3]  ( .D(n23999), .CK(clk), .Q(\mem[263][3] ) );
  DFF_X1 \mem_reg[263][2]  ( .D(n24000), .CK(clk), .Q(\mem[263][2] ) );
  DFF_X1 \mem_reg[263][1]  ( .D(n24001), .CK(clk), .Q(\mem[263][1] ) );
  DFF_X1 \mem_reg[263][0]  ( .D(n24002), .CK(clk), .Q(\mem[263][0] ) );
  DFF_X1 \mem_reg[262][7]  ( .D(n24003), .CK(clk), .Q(\mem[262][7] ) );
  DFF_X1 \mem_reg[262][6]  ( .D(n24004), .CK(clk), .Q(\mem[262][6] ) );
  DFF_X1 \mem_reg[262][5]  ( .D(n24005), .CK(clk), .Q(\mem[262][5] ) );
  DFF_X1 \mem_reg[262][4]  ( .D(n24006), .CK(clk), .Q(\mem[262][4] ) );
  DFF_X1 \mem_reg[262][3]  ( .D(n24007), .CK(clk), .Q(\mem[262][3] ) );
  DFF_X1 \mem_reg[262][2]  ( .D(n24008), .CK(clk), .Q(\mem[262][2] ) );
  DFF_X1 \mem_reg[262][1]  ( .D(n24009), .CK(clk), .Q(\mem[262][1] ) );
  DFF_X1 \mem_reg[262][0]  ( .D(n24010), .CK(clk), .Q(\mem[262][0] ) );
  DFF_X1 \mem_reg[261][7]  ( .D(n24011), .CK(clk), .Q(\mem[261][7] ) );
  DFF_X1 \mem_reg[261][6]  ( .D(n24012), .CK(clk), .Q(\mem[261][6] ) );
  DFF_X1 \mem_reg[261][5]  ( .D(n24013), .CK(clk), .Q(\mem[261][5] ) );
  DFF_X1 \mem_reg[261][4]  ( .D(n24014), .CK(clk), .Q(\mem[261][4] ) );
  DFF_X1 \mem_reg[261][3]  ( .D(n24015), .CK(clk), .Q(\mem[261][3] ) );
  DFF_X1 \mem_reg[261][2]  ( .D(n24016), .CK(clk), .Q(\mem[261][2] ) );
  DFF_X1 \mem_reg[261][1]  ( .D(n24017), .CK(clk), .Q(\mem[261][1] ) );
  DFF_X1 \mem_reg[261][0]  ( .D(n24018), .CK(clk), .Q(\mem[261][0] ) );
  DFF_X1 \mem_reg[260][7]  ( .D(n24019), .CK(clk), .Q(\mem[260][7] ) );
  DFF_X1 \mem_reg[260][6]  ( .D(n24020), .CK(clk), .Q(\mem[260][6] ) );
  DFF_X1 \mem_reg[260][5]  ( .D(n24021), .CK(clk), .Q(\mem[260][5] ) );
  DFF_X1 \mem_reg[260][4]  ( .D(n24022), .CK(clk), .Q(\mem[260][4] ) );
  DFF_X1 \mem_reg[260][3]  ( .D(n24023), .CK(clk), .Q(\mem[260][3] ) );
  DFF_X1 \mem_reg[260][2]  ( .D(n24024), .CK(clk), .Q(\mem[260][2] ) );
  DFF_X1 \mem_reg[260][1]  ( .D(n24025), .CK(clk), .Q(\mem[260][1] ) );
  DFF_X1 \mem_reg[260][0]  ( .D(n24026), .CK(clk), .Q(\mem[260][0] ) );
  DFF_X1 \mem_reg[259][7]  ( .D(n24027), .CK(clk), .Q(\mem[259][7] ) );
  DFF_X1 \mem_reg[259][6]  ( .D(n24028), .CK(clk), .Q(\mem[259][6] ) );
  DFF_X1 \mem_reg[259][5]  ( .D(n24029), .CK(clk), .Q(\mem[259][5] ) );
  DFF_X1 \mem_reg[259][4]  ( .D(n24030), .CK(clk), .Q(\mem[259][4] ) );
  DFF_X1 \mem_reg[259][3]  ( .D(n24031), .CK(clk), .Q(\mem[259][3] ) );
  DFF_X1 \mem_reg[259][2]  ( .D(n24032), .CK(clk), .Q(\mem[259][2] ) );
  DFF_X1 \mem_reg[259][1]  ( .D(n24033), .CK(clk), .Q(\mem[259][1] ) );
  DFF_X1 \mem_reg[259][0]  ( .D(n24034), .CK(clk), .Q(\mem[259][0] ) );
  DFF_X1 \mem_reg[258][7]  ( .D(n24035), .CK(clk), .Q(\mem[258][7] ) );
  DFF_X1 \mem_reg[258][6]  ( .D(n24036), .CK(clk), .Q(\mem[258][6] ) );
  DFF_X1 \mem_reg[258][5]  ( .D(n24037), .CK(clk), .Q(\mem[258][5] ) );
  DFF_X1 \mem_reg[258][4]  ( .D(n24038), .CK(clk), .Q(\mem[258][4] ) );
  DFF_X1 \mem_reg[258][3]  ( .D(n24039), .CK(clk), .Q(\mem[258][3] ) );
  DFF_X1 \mem_reg[258][2]  ( .D(n24040), .CK(clk), .Q(\mem[258][2] ) );
  DFF_X1 \mem_reg[258][1]  ( .D(n24041), .CK(clk), .Q(\mem[258][1] ) );
  DFF_X1 \mem_reg[258][0]  ( .D(n24042), .CK(clk), .Q(\mem[258][0] ) );
  DFF_X1 \mem_reg[257][7]  ( .D(n24043), .CK(clk), .Q(\mem[257][7] ) );
  DFF_X1 \mem_reg[257][6]  ( .D(n24044), .CK(clk), .Q(\mem[257][6] ) );
  DFF_X1 \mem_reg[257][5]  ( .D(n24045), .CK(clk), .Q(\mem[257][5] ) );
  DFF_X1 \mem_reg[257][4]  ( .D(n24046), .CK(clk), .Q(\mem[257][4] ) );
  DFF_X1 \mem_reg[257][3]  ( .D(n24047), .CK(clk), .Q(\mem[257][3] ) );
  DFF_X1 \mem_reg[257][2]  ( .D(n24048), .CK(clk), .Q(\mem[257][2] ) );
  DFF_X1 \mem_reg[257][1]  ( .D(n24049), .CK(clk), .Q(\mem[257][1] ) );
  DFF_X1 \mem_reg[257][0]  ( .D(n24050), .CK(clk), .Q(\mem[257][0] ) );
  DFF_X1 \mem_reg[256][7]  ( .D(n24051), .CK(clk), .Q(\mem[256][7] ) );
  DFF_X1 \mem_reg[256][6]  ( .D(n24052), .CK(clk), .Q(\mem[256][6] ) );
  DFF_X1 \mem_reg[256][5]  ( .D(n24053), .CK(clk), .Q(\mem[256][5] ) );
  DFF_X1 \mem_reg[256][4]  ( .D(n24054), .CK(clk), .Q(\mem[256][4] ) );
  DFF_X1 \mem_reg[256][3]  ( .D(n24055), .CK(clk), .Q(\mem[256][3] ) );
  DFF_X1 \mem_reg[256][2]  ( .D(n24056), .CK(clk), .Q(\mem[256][2] ) );
  DFF_X1 \mem_reg[256][1]  ( .D(n24057), .CK(clk), .Q(\mem[256][1] ) );
  DFF_X1 \mem_reg[256][0]  ( .D(n24058), .CK(clk), .Q(\mem[256][0] ) );
  DFF_X1 \mem_reg[255][7]  ( .D(n24059), .CK(clk), .Q(\mem[255][7] ) );
  DFF_X1 \mem_reg[255][6]  ( .D(n24060), .CK(clk), .Q(\mem[255][6] ) );
  DFF_X1 \mem_reg[255][5]  ( .D(n24061), .CK(clk), .Q(\mem[255][5] ) );
  DFF_X1 \mem_reg[255][4]  ( .D(n24062), .CK(clk), .Q(\mem[255][4] ) );
  DFF_X1 \mem_reg[255][3]  ( .D(n24063), .CK(clk), .Q(\mem[255][3] ) );
  DFF_X1 \mem_reg[255][2]  ( .D(n24064), .CK(clk), .Q(\mem[255][2] ) );
  DFF_X1 \mem_reg[255][1]  ( .D(n24065), .CK(clk), .Q(\mem[255][1] ) );
  DFF_X1 \mem_reg[255][0]  ( .D(n24066), .CK(clk), .Q(\mem[255][0] ) );
  DFF_X1 \mem_reg[254][7]  ( .D(n24067), .CK(clk), .Q(\mem[254][7] ) );
  DFF_X1 \mem_reg[254][6]  ( .D(n24068), .CK(clk), .Q(\mem[254][6] ) );
  DFF_X1 \mem_reg[254][5]  ( .D(n24069), .CK(clk), .Q(\mem[254][5] ) );
  DFF_X1 \mem_reg[254][4]  ( .D(n24070), .CK(clk), .Q(\mem[254][4] ) );
  DFF_X1 \mem_reg[254][3]  ( .D(n24071), .CK(clk), .Q(\mem[254][3] ) );
  DFF_X1 \mem_reg[254][2]  ( .D(n24072), .CK(clk), .Q(\mem[254][2] ) );
  DFF_X1 \mem_reg[254][1]  ( .D(n24073), .CK(clk), .Q(\mem[254][1] ) );
  DFF_X1 \mem_reg[254][0]  ( .D(n24074), .CK(clk), .Q(\mem[254][0] ) );
  DFF_X1 \mem_reg[253][7]  ( .D(n24075), .CK(clk), .Q(\mem[253][7] ) );
  DFF_X1 \mem_reg[253][6]  ( .D(n24076), .CK(clk), .Q(\mem[253][6] ) );
  DFF_X1 \mem_reg[253][5]  ( .D(n24077), .CK(clk), .Q(\mem[253][5] ) );
  DFF_X1 \mem_reg[253][4]  ( .D(n24078), .CK(clk), .Q(\mem[253][4] ) );
  DFF_X1 \mem_reg[253][3]  ( .D(n24079), .CK(clk), .Q(\mem[253][3] ) );
  DFF_X1 \mem_reg[253][2]  ( .D(n24080), .CK(clk), .Q(\mem[253][2] ) );
  DFF_X1 \mem_reg[253][1]  ( .D(n24081), .CK(clk), .Q(\mem[253][1] ) );
  DFF_X1 \mem_reg[253][0]  ( .D(n24082), .CK(clk), .Q(\mem[253][0] ) );
  DFF_X1 \mem_reg[252][7]  ( .D(n24083), .CK(clk), .Q(\mem[252][7] ) );
  DFF_X1 \mem_reg[252][6]  ( .D(n24084), .CK(clk), .Q(\mem[252][6] ) );
  DFF_X1 \mem_reg[252][5]  ( .D(n24085), .CK(clk), .Q(\mem[252][5] ) );
  DFF_X1 \mem_reg[252][4]  ( .D(n24086), .CK(clk), .Q(\mem[252][4] ) );
  DFF_X1 \mem_reg[252][3]  ( .D(n24087), .CK(clk), .Q(\mem[252][3] ) );
  DFF_X1 \mem_reg[252][2]  ( .D(n24088), .CK(clk), .Q(\mem[252][2] ) );
  DFF_X1 \mem_reg[252][1]  ( .D(n24089), .CK(clk), .Q(\mem[252][1] ) );
  DFF_X1 \mem_reg[252][0]  ( .D(n24090), .CK(clk), .Q(\mem[252][0] ) );
  DFF_X1 \mem_reg[251][7]  ( .D(n24091), .CK(clk), .Q(\mem[251][7] ) );
  DFF_X1 \mem_reg[251][6]  ( .D(n24092), .CK(clk), .Q(\mem[251][6] ) );
  DFF_X1 \mem_reg[251][5]  ( .D(n24093), .CK(clk), .Q(\mem[251][5] ) );
  DFF_X1 \mem_reg[251][4]  ( .D(n24094), .CK(clk), .Q(\mem[251][4] ) );
  DFF_X1 \mem_reg[251][3]  ( .D(n24095), .CK(clk), .Q(\mem[251][3] ) );
  DFF_X1 \mem_reg[251][2]  ( .D(n24096), .CK(clk), .Q(\mem[251][2] ) );
  DFF_X1 \mem_reg[251][1]  ( .D(n24097), .CK(clk), .Q(\mem[251][1] ) );
  DFF_X1 \mem_reg[251][0]  ( .D(n24098), .CK(clk), .Q(\mem[251][0] ) );
  DFF_X1 \mem_reg[250][7]  ( .D(n24099), .CK(clk), .Q(\mem[250][7] ) );
  DFF_X1 \mem_reg[250][6]  ( .D(n24100), .CK(clk), .Q(\mem[250][6] ) );
  DFF_X1 \mem_reg[250][5]  ( .D(n24101), .CK(clk), .Q(\mem[250][5] ) );
  DFF_X1 \mem_reg[250][4]  ( .D(n24102), .CK(clk), .Q(\mem[250][4] ) );
  DFF_X1 \mem_reg[250][3]  ( .D(n24103), .CK(clk), .Q(\mem[250][3] ) );
  DFF_X1 \mem_reg[250][2]  ( .D(n24104), .CK(clk), .Q(\mem[250][2] ) );
  DFF_X1 \mem_reg[250][1]  ( .D(n24105), .CK(clk), .Q(\mem[250][1] ) );
  DFF_X1 \mem_reg[250][0]  ( .D(n24106), .CK(clk), .Q(\mem[250][0] ) );
  DFF_X1 \mem_reg[249][7]  ( .D(n24107), .CK(clk), .Q(\mem[249][7] ) );
  DFF_X1 \mem_reg[249][6]  ( .D(n24108), .CK(clk), .Q(\mem[249][6] ) );
  DFF_X1 \mem_reg[249][5]  ( .D(n24109), .CK(clk), .Q(\mem[249][5] ) );
  DFF_X1 \mem_reg[249][4]  ( .D(n24110), .CK(clk), .Q(\mem[249][4] ) );
  DFF_X1 \mem_reg[249][3]  ( .D(n24111), .CK(clk), .Q(\mem[249][3] ) );
  DFF_X1 \mem_reg[249][2]  ( .D(n24112), .CK(clk), .Q(\mem[249][2] ) );
  DFF_X1 \mem_reg[249][1]  ( .D(n24113), .CK(clk), .Q(\mem[249][1] ) );
  DFF_X1 \mem_reg[249][0]  ( .D(n24114), .CK(clk), .Q(\mem[249][0] ) );
  DFF_X1 \mem_reg[248][7]  ( .D(n24115), .CK(clk), .Q(\mem[248][7] ) );
  DFF_X1 \mem_reg[248][6]  ( .D(n24116), .CK(clk), .Q(\mem[248][6] ) );
  DFF_X1 \mem_reg[248][5]  ( .D(n24117), .CK(clk), .Q(\mem[248][5] ) );
  DFF_X1 \mem_reg[248][4]  ( .D(n24118), .CK(clk), .Q(\mem[248][4] ) );
  DFF_X1 \mem_reg[248][3]  ( .D(n24119), .CK(clk), .Q(\mem[248][3] ) );
  DFF_X1 \mem_reg[248][2]  ( .D(n24120), .CK(clk), .Q(\mem[248][2] ) );
  DFF_X1 \mem_reg[248][1]  ( .D(n24121), .CK(clk), .Q(\mem[248][1] ) );
  DFF_X1 \mem_reg[248][0]  ( .D(n24122), .CK(clk), .Q(\mem[248][0] ) );
  DFF_X1 \mem_reg[247][7]  ( .D(n24123), .CK(clk), .Q(\mem[247][7] ) );
  DFF_X1 \mem_reg[247][6]  ( .D(n24124), .CK(clk), .Q(\mem[247][6] ) );
  DFF_X1 \mem_reg[247][5]  ( .D(n24125), .CK(clk), .Q(\mem[247][5] ) );
  DFF_X1 \mem_reg[247][4]  ( .D(n24126), .CK(clk), .Q(\mem[247][4] ) );
  DFF_X1 \mem_reg[247][3]  ( .D(n24127), .CK(clk), .Q(\mem[247][3] ) );
  DFF_X1 \mem_reg[247][2]  ( .D(n24128), .CK(clk), .Q(\mem[247][2] ) );
  DFF_X1 \mem_reg[247][1]  ( .D(n24129), .CK(clk), .Q(\mem[247][1] ) );
  DFF_X1 \mem_reg[247][0]  ( .D(n24130), .CK(clk), .Q(\mem[247][0] ) );
  DFF_X1 \mem_reg[246][7]  ( .D(n24131), .CK(clk), .Q(\mem[246][7] ) );
  DFF_X1 \mem_reg[246][6]  ( .D(n24132), .CK(clk), .Q(\mem[246][6] ) );
  DFF_X1 \mem_reg[246][5]  ( .D(n24133), .CK(clk), .Q(\mem[246][5] ) );
  DFF_X1 \mem_reg[246][4]  ( .D(n24134), .CK(clk), .Q(\mem[246][4] ) );
  DFF_X1 \mem_reg[246][3]  ( .D(n24135), .CK(clk), .Q(\mem[246][3] ) );
  DFF_X1 \mem_reg[246][2]  ( .D(n24136), .CK(clk), .Q(\mem[246][2] ) );
  DFF_X1 \mem_reg[246][1]  ( .D(n24137), .CK(clk), .Q(\mem[246][1] ) );
  DFF_X1 \mem_reg[246][0]  ( .D(n24138), .CK(clk), .Q(\mem[246][0] ) );
  DFF_X1 \mem_reg[245][7]  ( .D(n24139), .CK(clk), .Q(\mem[245][7] ) );
  DFF_X1 \mem_reg[245][6]  ( .D(n24140), .CK(clk), .Q(\mem[245][6] ) );
  DFF_X1 \mem_reg[245][5]  ( .D(n24141), .CK(clk), .Q(\mem[245][5] ) );
  DFF_X1 \mem_reg[245][4]  ( .D(n24142), .CK(clk), .Q(\mem[245][4] ) );
  DFF_X1 \mem_reg[245][3]  ( .D(n24143), .CK(clk), .Q(\mem[245][3] ) );
  DFF_X1 \mem_reg[245][2]  ( .D(n24144), .CK(clk), .Q(\mem[245][2] ) );
  DFF_X1 \mem_reg[245][1]  ( .D(n24145), .CK(clk), .Q(\mem[245][1] ) );
  DFF_X1 \mem_reg[245][0]  ( .D(n24146), .CK(clk), .Q(\mem[245][0] ) );
  DFF_X1 \mem_reg[244][7]  ( .D(n24147), .CK(clk), .Q(\mem[244][7] ) );
  DFF_X1 \mem_reg[244][6]  ( .D(n24148), .CK(clk), .Q(\mem[244][6] ) );
  DFF_X1 \mem_reg[244][5]  ( .D(n24149), .CK(clk), .Q(\mem[244][5] ) );
  DFF_X1 \mem_reg[244][4]  ( .D(n24150), .CK(clk), .Q(\mem[244][4] ) );
  DFF_X1 \mem_reg[244][3]  ( .D(n24151), .CK(clk), .Q(\mem[244][3] ) );
  DFF_X1 \mem_reg[244][2]  ( .D(n24152), .CK(clk), .Q(\mem[244][2] ) );
  DFF_X1 \mem_reg[244][1]  ( .D(n24153), .CK(clk), .Q(\mem[244][1] ) );
  DFF_X1 \mem_reg[244][0]  ( .D(n24154), .CK(clk), .Q(\mem[244][0] ) );
  DFF_X1 \mem_reg[243][7]  ( .D(n24155), .CK(clk), .Q(\mem[243][7] ) );
  DFF_X1 \mem_reg[243][6]  ( .D(n24156), .CK(clk), .Q(\mem[243][6] ) );
  DFF_X1 \mem_reg[243][5]  ( .D(n24157), .CK(clk), .Q(\mem[243][5] ) );
  DFF_X1 \mem_reg[243][4]  ( .D(n24158), .CK(clk), .Q(\mem[243][4] ) );
  DFF_X1 \mem_reg[243][3]  ( .D(n24159), .CK(clk), .Q(\mem[243][3] ) );
  DFF_X1 \mem_reg[243][2]  ( .D(n24160), .CK(clk), .Q(\mem[243][2] ) );
  DFF_X1 \mem_reg[243][1]  ( .D(n24161), .CK(clk), .Q(\mem[243][1] ) );
  DFF_X1 \mem_reg[243][0]  ( .D(n24162), .CK(clk), .Q(\mem[243][0] ) );
  DFF_X1 \mem_reg[242][7]  ( .D(n24163), .CK(clk), .Q(\mem[242][7] ) );
  DFF_X1 \mem_reg[242][6]  ( .D(n24164), .CK(clk), .Q(\mem[242][6] ) );
  DFF_X1 \mem_reg[242][5]  ( .D(n24165), .CK(clk), .Q(\mem[242][5] ) );
  DFF_X1 \mem_reg[242][4]  ( .D(n24166), .CK(clk), .Q(\mem[242][4] ) );
  DFF_X1 \mem_reg[242][3]  ( .D(n24167), .CK(clk), .Q(\mem[242][3] ) );
  DFF_X1 \mem_reg[242][2]  ( .D(n24168), .CK(clk), .Q(\mem[242][2] ) );
  DFF_X1 \mem_reg[242][1]  ( .D(n24169), .CK(clk), .Q(\mem[242][1] ) );
  DFF_X1 \mem_reg[242][0]  ( .D(n24170), .CK(clk), .Q(\mem[242][0] ) );
  DFF_X1 \mem_reg[241][7]  ( .D(n24171), .CK(clk), .Q(\mem[241][7] ) );
  DFF_X1 \mem_reg[241][6]  ( .D(n24172), .CK(clk), .Q(\mem[241][6] ) );
  DFF_X1 \mem_reg[241][5]  ( .D(n24173), .CK(clk), .Q(\mem[241][5] ) );
  DFF_X1 \mem_reg[241][4]  ( .D(n24174), .CK(clk), .Q(\mem[241][4] ) );
  DFF_X1 \mem_reg[241][3]  ( .D(n24175), .CK(clk), .Q(\mem[241][3] ) );
  DFF_X1 \mem_reg[241][2]  ( .D(n24176), .CK(clk), .Q(\mem[241][2] ) );
  DFF_X1 \mem_reg[241][1]  ( .D(n24177), .CK(clk), .Q(\mem[241][1] ) );
  DFF_X1 \mem_reg[241][0]  ( .D(n24178), .CK(clk), .Q(\mem[241][0] ) );
  DFF_X1 \mem_reg[240][7]  ( .D(n24179), .CK(clk), .Q(\mem[240][7] ) );
  DFF_X1 \mem_reg[240][6]  ( .D(n24180), .CK(clk), .Q(\mem[240][6] ) );
  DFF_X1 \mem_reg[240][5]  ( .D(n24181), .CK(clk), .Q(\mem[240][5] ) );
  DFF_X1 \mem_reg[240][4]  ( .D(n24182), .CK(clk), .Q(\mem[240][4] ) );
  DFF_X1 \mem_reg[240][3]  ( .D(n24183), .CK(clk), .Q(\mem[240][3] ) );
  DFF_X1 \mem_reg[240][2]  ( .D(n24184), .CK(clk), .Q(\mem[240][2] ) );
  DFF_X1 \mem_reg[240][1]  ( .D(n24185), .CK(clk), .Q(\mem[240][1] ) );
  DFF_X1 \mem_reg[240][0]  ( .D(n24186), .CK(clk), .Q(\mem[240][0] ) );
  DFF_X1 \mem_reg[239][7]  ( .D(n24187), .CK(clk), .Q(\mem[239][7] ) );
  DFF_X1 \mem_reg[239][6]  ( .D(n24188), .CK(clk), .Q(\mem[239][6] ) );
  DFF_X1 \mem_reg[239][5]  ( .D(n24189), .CK(clk), .Q(\mem[239][5] ) );
  DFF_X1 \mem_reg[239][4]  ( .D(n24190), .CK(clk), .Q(\mem[239][4] ) );
  DFF_X1 \mem_reg[239][3]  ( .D(n24191), .CK(clk), .Q(\mem[239][3] ) );
  DFF_X1 \mem_reg[239][2]  ( .D(n24192), .CK(clk), .Q(\mem[239][2] ) );
  DFF_X1 \mem_reg[239][1]  ( .D(n24193), .CK(clk), .Q(\mem[239][1] ) );
  DFF_X1 \mem_reg[239][0]  ( .D(n24194), .CK(clk), .Q(\mem[239][0] ) );
  DFF_X1 \mem_reg[238][7]  ( .D(n24195), .CK(clk), .Q(\mem[238][7] ) );
  DFF_X1 \mem_reg[238][6]  ( .D(n24196), .CK(clk), .Q(\mem[238][6] ) );
  DFF_X1 \mem_reg[238][5]  ( .D(n24197), .CK(clk), .Q(\mem[238][5] ) );
  DFF_X1 \mem_reg[238][4]  ( .D(n24198), .CK(clk), .Q(\mem[238][4] ) );
  DFF_X1 \mem_reg[238][3]  ( .D(n24199), .CK(clk), .Q(\mem[238][3] ) );
  DFF_X1 \mem_reg[238][2]  ( .D(n24200), .CK(clk), .Q(\mem[238][2] ) );
  DFF_X1 \mem_reg[238][1]  ( .D(n24201), .CK(clk), .Q(\mem[238][1] ) );
  DFF_X1 \mem_reg[238][0]  ( .D(n24202), .CK(clk), .Q(\mem[238][0] ) );
  DFF_X1 \mem_reg[237][7]  ( .D(n24203), .CK(clk), .Q(\mem[237][7] ) );
  DFF_X1 \mem_reg[237][6]  ( .D(n24204), .CK(clk), .Q(\mem[237][6] ) );
  DFF_X1 \mem_reg[237][5]  ( .D(n24205), .CK(clk), .Q(\mem[237][5] ) );
  DFF_X1 \mem_reg[237][4]  ( .D(n24206), .CK(clk), .Q(\mem[237][4] ) );
  DFF_X1 \mem_reg[237][3]  ( .D(n24207), .CK(clk), .Q(\mem[237][3] ) );
  DFF_X1 \mem_reg[237][2]  ( .D(n24208), .CK(clk), .Q(\mem[237][2] ) );
  DFF_X1 \mem_reg[237][1]  ( .D(n24209), .CK(clk), .Q(\mem[237][1] ) );
  DFF_X1 \mem_reg[237][0]  ( .D(n24210), .CK(clk), .Q(\mem[237][0] ) );
  DFF_X1 \mem_reg[236][7]  ( .D(n24211), .CK(clk), .Q(\mem[236][7] ) );
  DFF_X1 \mem_reg[236][6]  ( .D(n24212), .CK(clk), .Q(\mem[236][6] ) );
  DFF_X1 \mem_reg[236][5]  ( .D(n24213), .CK(clk), .Q(\mem[236][5] ) );
  DFF_X1 \mem_reg[236][4]  ( .D(n24214), .CK(clk), .Q(\mem[236][4] ) );
  DFF_X1 \mem_reg[236][3]  ( .D(n24215), .CK(clk), .Q(\mem[236][3] ) );
  DFF_X1 \mem_reg[236][2]  ( .D(n24216), .CK(clk), .Q(\mem[236][2] ) );
  DFF_X1 \mem_reg[236][1]  ( .D(n24217), .CK(clk), .Q(\mem[236][1] ) );
  DFF_X1 \mem_reg[236][0]  ( .D(n24218), .CK(clk), .Q(\mem[236][0] ) );
  DFF_X1 \mem_reg[235][7]  ( .D(n24219), .CK(clk), .Q(\mem[235][7] ) );
  DFF_X1 \mem_reg[235][6]  ( .D(n24220), .CK(clk), .Q(\mem[235][6] ) );
  DFF_X1 \mem_reg[235][5]  ( .D(n24221), .CK(clk), .Q(\mem[235][5] ) );
  DFF_X1 \mem_reg[235][4]  ( .D(n24222), .CK(clk), .Q(\mem[235][4] ) );
  DFF_X1 \mem_reg[235][3]  ( .D(n24223), .CK(clk), .Q(\mem[235][3] ) );
  DFF_X1 \mem_reg[235][2]  ( .D(n24224), .CK(clk), .Q(\mem[235][2] ) );
  DFF_X1 \mem_reg[235][1]  ( .D(n24225), .CK(clk), .Q(\mem[235][1] ) );
  DFF_X1 \mem_reg[235][0]  ( .D(n24226), .CK(clk), .Q(\mem[235][0] ) );
  DFF_X1 \mem_reg[234][7]  ( .D(n24227), .CK(clk), .Q(\mem[234][7] ) );
  DFF_X1 \mem_reg[234][6]  ( .D(n24228), .CK(clk), .Q(\mem[234][6] ) );
  DFF_X1 \mem_reg[234][5]  ( .D(n24229), .CK(clk), .Q(\mem[234][5] ) );
  DFF_X1 \mem_reg[234][4]  ( .D(n24230), .CK(clk), .Q(\mem[234][4] ) );
  DFF_X1 \mem_reg[234][3]  ( .D(n24231), .CK(clk), .Q(\mem[234][3] ) );
  DFF_X1 \mem_reg[234][2]  ( .D(n24232), .CK(clk), .Q(\mem[234][2] ) );
  DFF_X1 \mem_reg[234][1]  ( .D(n24233), .CK(clk), .Q(\mem[234][1] ) );
  DFF_X1 \mem_reg[234][0]  ( .D(n24234), .CK(clk), .Q(\mem[234][0] ) );
  DFF_X1 \mem_reg[233][7]  ( .D(n24235), .CK(clk), .Q(\mem[233][7] ) );
  DFF_X1 \mem_reg[233][6]  ( .D(n24236), .CK(clk), .Q(\mem[233][6] ) );
  DFF_X1 \mem_reg[233][5]  ( .D(n24237), .CK(clk), .Q(\mem[233][5] ) );
  DFF_X1 \mem_reg[233][4]  ( .D(n24238), .CK(clk), .Q(\mem[233][4] ) );
  DFF_X1 \mem_reg[233][3]  ( .D(n24239), .CK(clk), .Q(\mem[233][3] ) );
  DFF_X1 \mem_reg[233][2]  ( .D(n24240), .CK(clk), .Q(\mem[233][2] ) );
  DFF_X1 \mem_reg[233][1]  ( .D(n24241), .CK(clk), .Q(\mem[233][1] ) );
  DFF_X1 \mem_reg[233][0]  ( .D(n24242), .CK(clk), .Q(\mem[233][0] ) );
  DFF_X1 \mem_reg[232][7]  ( .D(n24243), .CK(clk), .Q(\mem[232][7] ) );
  DFF_X1 \mem_reg[232][6]  ( .D(n24244), .CK(clk), .Q(\mem[232][6] ) );
  DFF_X1 \mem_reg[232][5]  ( .D(n24245), .CK(clk), .Q(\mem[232][5] ) );
  DFF_X1 \mem_reg[232][4]  ( .D(n24246), .CK(clk), .Q(\mem[232][4] ) );
  DFF_X1 \mem_reg[232][3]  ( .D(n24247), .CK(clk), .Q(\mem[232][3] ) );
  DFF_X1 \mem_reg[232][2]  ( .D(n24248), .CK(clk), .Q(\mem[232][2] ) );
  DFF_X1 \mem_reg[232][1]  ( .D(n24249), .CK(clk), .Q(\mem[232][1] ) );
  DFF_X1 \mem_reg[232][0]  ( .D(n24250), .CK(clk), .Q(\mem[232][0] ) );
  DFF_X1 \mem_reg[231][7]  ( .D(n24251), .CK(clk), .Q(\mem[231][7] ) );
  DFF_X1 \mem_reg[231][6]  ( .D(n24252), .CK(clk), .Q(\mem[231][6] ) );
  DFF_X1 \mem_reg[231][5]  ( .D(n24253), .CK(clk), .Q(\mem[231][5] ) );
  DFF_X1 \mem_reg[231][4]  ( .D(n24254), .CK(clk), .Q(\mem[231][4] ) );
  DFF_X1 \mem_reg[231][3]  ( .D(n24255), .CK(clk), .Q(\mem[231][3] ) );
  DFF_X1 \mem_reg[231][2]  ( .D(n24256), .CK(clk), .Q(\mem[231][2] ) );
  DFF_X1 \mem_reg[231][1]  ( .D(n24257), .CK(clk), .Q(\mem[231][1] ) );
  DFF_X1 \mem_reg[231][0]  ( .D(n24258), .CK(clk), .Q(\mem[231][0] ) );
  DFF_X1 \mem_reg[230][7]  ( .D(n24259), .CK(clk), .Q(\mem[230][7] ) );
  DFF_X1 \mem_reg[230][6]  ( .D(n24260), .CK(clk), .Q(\mem[230][6] ) );
  DFF_X1 \mem_reg[230][5]  ( .D(n24261), .CK(clk), .Q(\mem[230][5] ) );
  DFF_X1 \mem_reg[230][4]  ( .D(n24262), .CK(clk), .Q(\mem[230][4] ) );
  DFF_X1 \mem_reg[230][3]  ( .D(n24263), .CK(clk), .Q(\mem[230][3] ) );
  DFF_X1 \mem_reg[230][2]  ( .D(n24264), .CK(clk), .Q(\mem[230][2] ) );
  DFF_X1 \mem_reg[230][1]  ( .D(n24265), .CK(clk), .Q(\mem[230][1] ) );
  DFF_X1 \mem_reg[230][0]  ( .D(n24266), .CK(clk), .Q(\mem[230][0] ) );
  DFF_X1 \mem_reg[229][7]  ( .D(n24267), .CK(clk), .Q(\mem[229][7] ) );
  DFF_X1 \mem_reg[229][6]  ( .D(n24268), .CK(clk), .Q(\mem[229][6] ) );
  DFF_X1 \mem_reg[229][5]  ( .D(n24269), .CK(clk), .Q(\mem[229][5] ) );
  DFF_X1 \mem_reg[229][4]  ( .D(n24270), .CK(clk), .Q(\mem[229][4] ) );
  DFF_X1 \mem_reg[229][3]  ( .D(n24271), .CK(clk), .Q(\mem[229][3] ) );
  DFF_X1 \mem_reg[229][2]  ( .D(n24272), .CK(clk), .Q(\mem[229][2] ) );
  DFF_X1 \mem_reg[229][1]  ( .D(n24273), .CK(clk), .Q(\mem[229][1] ) );
  DFF_X1 \mem_reg[229][0]  ( .D(n24274), .CK(clk), .Q(\mem[229][0] ) );
  DFF_X1 \mem_reg[228][7]  ( .D(n24275), .CK(clk), .Q(\mem[228][7] ) );
  DFF_X1 \mem_reg[228][6]  ( .D(n24276), .CK(clk), .Q(\mem[228][6] ) );
  DFF_X1 \mem_reg[228][5]  ( .D(n24277), .CK(clk), .Q(\mem[228][5] ) );
  DFF_X1 \mem_reg[228][4]  ( .D(n24278), .CK(clk), .Q(\mem[228][4] ) );
  DFF_X1 \mem_reg[228][3]  ( .D(n24279), .CK(clk), .Q(\mem[228][3] ) );
  DFF_X1 \mem_reg[228][2]  ( .D(n24280), .CK(clk), .Q(\mem[228][2] ) );
  DFF_X1 \mem_reg[228][1]  ( .D(n24281), .CK(clk), .Q(\mem[228][1] ) );
  DFF_X1 \mem_reg[228][0]  ( .D(n24282), .CK(clk), .Q(\mem[228][0] ) );
  DFF_X1 \mem_reg[227][7]  ( .D(n24283), .CK(clk), .Q(\mem[227][7] ) );
  DFF_X1 \mem_reg[227][6]  ( .D(n24284), .CK(clk), .Q(\mem[227][6] ) );
  DFF_X1 \mem_reg[227][5]  ( .D(n24285), .CK(clk), .Q(\mem[227][5] ) );
  DFF_X1 \mem_reg[227][4]  ( .D(n24286), .CK(clk), .Q(\mem[227][4] ) );
  DFF_X1 \mem_reg[227][3]  ( .D(n24287), .CK(clk), .Q(\mem[227][3] ) );
  DFF_X1 \mem_reg[227][2]  ( .D(n24288), .CK(clk), .Q(\mem[227][2] ) );
  DFF_X1 \mem_reg[227][1]  ( .D(n24289), .CK(clk), .Q(\mem[227][1] ) );
  DFF_X1 \mem_reg[227][0]  ( .D(n24290), .CK(clk), .Q(\mem[227][0] ) );
  DFF_X1 \mem_reg[226][7]  ( .D(n24291), .CK(clk), .Q(\mem[226][7] ) );
  DFF_X1 \mem_reg[226][6]  ( .D(n24292), .CK(clk), .Q(\mem[226][6] ) );
  DFF_X1 \mem_reg[226][5]  ( .D(n24293), .CK(clk), .Q(\mem[226][5] ) );
  DFF_X1 \mem_reg[226][4]  ( .D(n24294), .CK(clk), .Q(\mem[226][4] ) );
  DFF_X1 \mem_reg[226][3]  ( .D(n24295), .CK(clk), .Q(\mem[226][3] ) );
  DFF_X1 \mem_reg[226][2]  ( .D(n24296), .CK(clk), .Q(\mem[226][2] ) );
  DFF_X1 \mem_reg[226][1]  ( .D(n24297), .CK(clk), .Q(\mem[226][1] ) );
  DFF_X1 \mem_reg[226][0]  ( .D(n24298), .CK(clk), .Q(\mem[226][0] ) );
  DFF_X1 \mem_reg[225][7]  ( .D(n24299), .CK(clk), .Q(\mem[225][7] ) );
  DFF_X1 \mem_reg[225][6]  ( .D(n24300), .CK(clk), .Q(\mem[225][6] ) );
  DFF_X1 \mem_reg[225][5]  ( .D(n24301), .CK(clk), .Q(\mem[225][5] ) );
  DFF_X1 \mem_reg[225][4]  ( .D(n24302), .CK(clk), .Q(\mem[225][4] ) );
  DFF_X1 \mem_reg[225][3]  ( .D(n24303), .CK(clk), .Q(\mem[225][3] ) );
  DFF_X1 \mem_reg[225][2]  ( .D(n24304), .CK(clk), .Q(\mem[225][2] ) );
  DFF_X1 \mem_reg[225][1]  ( .D(n24305), .CK(clk), .Q(\mem[225][1] ) );
  DFF_X1 \mem_reg[225][0]  ( .D(n24306), .CK(clk), .Q(\mem[225][0] ) );
  DFF_X1 \mem_reg[224][7]  ( .D(n24307), .CK(clk), .Q(\mem[224][7] ) );
  DFF_X1 \mem_reg[224][6]  ( .D(n24308), .CK(clk), .Q(\mem[224][6] ) );
  DFF_X1 \mem_reg[224][5]  ( .D(n24309), .CK(clk), .Q(\mem[224][5] ) );
  DFF_X1 \mem_reg[224][4]  ( .D(n24310), .CK(clk), .Q(\mem[224][4] ) );
  DFF_X1 \mem_reg[224][3]  ( .D(n24311), .CK(clk), .Q(\mem[224][3] ) );
  DFF_X1 \mem_reg[224][2]  ( .D(n24312), .CK(clk), .Q(\mem[224][2] ) );
  DFF_X1 \mem_reg[224][1]  ( .D(n24313), .CK(clk), .Q(\mem[224][1] ) );
  DFF_X1 \mem_reg[224][0]  ( .D(n24314), .CK(clk), .Q(\mem[224][0] ) );
  DFF_X1 \mem_reg[223][7]  ( .D(n24315), .CK(clk), .Q(\mem[223][7] ) );
  DFF_X1 \mem_reg[223][6]  ( .D(n24316), .CK(clk), .Q(\mem[223][6] ) );
  DFF_X1 \mem_reg[223][5]  ( .D(n24317), .CK(clk), .Q(\mem[223][5] ) );
  DFF_X1 \mem_reg[223][4]  ( .D(n24318), .CK(clk), .Q(\mem[223][4] ) );
  DFF_X1 \mem_reg[223][3]  ( .D(n24319), .CK(clk), .Q(\mem[223][3] ) );
  DFF_X1 \mem_reg[223][2]  ( .D(n24320), .CK(clk), .Q(\mem[223][2] ) );
  DFF_X1 \mem_reg[223][1]  ( .D(n24321), .CK(clk), .Q(\mem[223][1] ) );
  DFF_X1 \mem_reg[223][0]  ( .D(n24322), .CK(clk), .Q(\mem[223][0] ) );
  DFF_X1 \mem_reg[222][7]  ( .D(n24323), .CK(clk), .Q(\mem[222][7] ) );
  DFF_X1 \mem_reg[222][6]  ( .D(n24324), .CK(clk), .Q(\mem[222][6] ) );
  DFF_X1 \mem_reg[222][5]  ( .D(n24325), .CK(clk), .Q(\mem[222][5] ) );
  DFF_X1 \mem_reg[222][4]  ( .D(n24326), .CK(clk), .Q(\mem[222][4] ) );
  DFF_X1 \mem_reg[222][3]  ( .D(n24327), .CK(clk), .Q(\mem[222][3] ) );
  DFF_X1 \mem_reg[222][2]  ( .D(n24328), .CK(clk), .Q(\mem[222][2] ) );
  DFF_X1 \mem_reg[222][1]  ( .D(n24329), .CK(clk), .Q(\mem[222][1] ) );
  DFF_X1 \mem_reg[222][0]  ( .D(n24330), .CK(clk), .Q(\mem[222][0] ) );
  DFF_X1 \mem_reg[221][7]  ( .D(n24331), .CK(clk), .Q(\mem[221][7] ) );
  DFF_X1 \mem_reg[221][6]  ( .D(n24332), .CK(clk), .Q(\mem[221][6] ) );
  DFF_X1 \mem_reg[221][5]  ( .D(n24333), .CK(clk), .Q(\mem[221][5] ) );
  DFF_X1 \mem_reg[221][4]  ( .D(n24334), .CK(clk), .Q(\mem[221][4] ) );
  DFF_X1 \mem_reg[221][3]  ( .D(n24335), .CK(clk), .Q(\mem[221][3] ) );
  DFF_X1 \mem_reg[221][2]  ( .D(n24336), .CK(clk), .Q(\mem[221][2] ) );
  DFF_X1 \mem_reg[221][1]  ( .D(n24337), .CK(clk), .Q(\mem[221][1] ) );
  DFF_X1 \mem_reg[221][0]  ( .D(n24338), .CK(clk), .Q(\mem[221][0] ) );
  DFF_X1 \mem_reg[220][7]  ( .D(n24339), .CK(clk), .Q(\mem[220][7] ) );
  DFF_X1 \mem_reg[220][6]  ( .D(n24340), .CK(clk), .Q(\mem[220][6] ) );
  DFF_X1 \mem_reg[220][5]  ( .D(n24341), .CK(clk), .Q(\mem[220][5] ) );
  DFF_X1 \mem_reg[220][4]  ( .D(n24342), .CK(clk), .Q(\mem[220][4] ) );
  DFF_X1 \mem_reg[220][3]  ( .D(n24343), .CK(clk), .Q(\mem[220][3] ) );
  DFF_X1 \mem_reg[220][2]  ( .D(n24344), .CK(clk), .Q(\mem[220][2] ) );
  DFF_X1 \mem_reg[220][1]  ( .D(n24345), .CK(clk), .Q(\mem[220][1] ) );
  DFF_X1 \mem_reg[220][0]  ( .D(n24346), .CK(clk), .Q(\mem[220][0] ) );
  DFF_X1 \mem_reg[219][7]  ( .D(n24347), .CK(clk), .Q(\mem[219][7] ) );
  DFF_X1 \mem_reg[219][6]  ( .D(n24348), .CK(clk), .Q(\mem[219][6] ) );
  DFF_X1 \mem_reg[219][5]  ( .D(n24349), .CK(clk), .Q(\mem[219][5] ) );
  DFF_X1 \mem_reg[219][4]  ( .D(n24350), .CK(clk), .Q(\mem[219][4] ) );
  DFF_X1 \mem_reg[219][3]  ( .D(n24351), .CK(clk), .Q(\mem[219][3] ) );
  DFF_X1 \mem_reg[219][2]  ( .D(n24352), .CK(clk), .Q(\mem[219][2] ) );
  DFF_X1 \mem_reg[219][1]  ( .D(n24353), .CK(clk), .Q(\mem[219][1] ) );
  DFF_X1 \mem_reg[219][0]  ( .D(n24354), .CK(clk), .Q(\mem[219][0] ) );
  DFF_X1 \mem_reg[218][7]  ( .D(n24355), .CK(clk), .Q(\mem[218][7] ) );
  DFF_X1 \mem_reg[218][6]  ( .D(n24356), .CK(clk), .Q(\mem[218][6] ) );
  DFF_X1 \mem_reg[218][5]  ( .D(n24357), .CK(clk), .Q(\mem[218][5] ) );
  DFF_X1 \mem_reg[218][4]  ( .D(n24358), .CK(clk), .Q(\mem[218][4] ) );
  DFF_X1 \mem_reg[218][3]  ( .D(n24359), .CK(clk), .Q(\mem[218][3] ) );
  DFF_X1 \mem_reg[218][2]  ( .D(n24360), .CK(clk), .Q(\mem[218][2] ) );
  DFF_X1 \mem_reg[218][1]  ( .D(n24361), .CK(clk), .Q(\mem[218][1] ) );
  DFF_X1 \mem_reg[218][0]  ( .D(n24362), .CK(clk), .Q(\mem[218][0] ) );
  DFF_X1 \mem_reg[217][7]  ( .D(n24363), .CK(clk), .Q(\mem[217][7] ) );
  DFF_X1 \mem_reg[217][6]  ( .D(n24364), .CK(clk), .Q(\mem[217][6] ) );
  DFF_X1 \mem_reg[217][5]  ( .D(n24365), .CK(clk), .Q(\mem[217][5] ) );
  DFF_X1 \mem_reg[217][4]  ( .D(n24366), .CK(clk), .Q(\mem[217][4] ) );
  DFF_X1 \mem_reg[217][3]  ( .D(n24367), .CK(clk), .Q(\mem[217][3] ) );
  DFF_X1 \mem_reg[217][2]  ( .D(n24368), .CK(clk), .Q(\mem[217][2] ) );
  DFF_X1 \mem_reg[217][1]  ( .D(n24369), .CK(clk), .Q(\mem[217][1] ) );
  DFF_X1 \mem_reg[217][0]  ( .D(n24370), .CK(clk), .Q(\mem[217][0] ) );
  DFF_X1 \mem_reg[216][7]  ( .D(n24371), .CK(clk), .Q(\mem[216][7] ) );
  DFF_X1 \mem_reg[216][6]  ( .D(n24372), .CK(clk), .Q(\mem[216][6] ) );
  DFF_X1 \mem_reg[216][5]  ( .D(n24373), .CK(clk), .Q(\mem[216][5] ) );
  DFF_X1 \mem_reg[216][4]  ( .D(n24374), .CK(clk), .Q(\mem[216][4] ) );
  DFF_X1 \mem_reg[216][3]  ( .D(n24375), .CK(clk), .Q(\mem[216][3] ) );
  DFF_X1 \mem_reg[216][2]  ( .D(n24376), .CK(clk), .Q(\mem[216][2] ) );
  DFF_X1 \mem_reg[216][1]  ( .D(n24377), .CK(clk), .Q(\mem[216][1] ) );
  DFF_X1 \mem_reg[216][0]  ( .D(n24378), .CK(clk), .Q(\mem[216][0] ) );
  DFF_X1 \mem_reg[215][7]  ( .D(n24379), .CK(clk), .Q(\mem[215][7] ) );
  DFF_X1 \mem_reg[215][6]  ( .D(n24380), .CK(clk), .Q(\mem[215][6] ) );
  DFF_X1 \mem_reg[215][5]  ( .D(n24381), .CK(clk), .Q(\mem[215][5] ) );
  DFF_X1 \mem_reg[215][4]  ( .D(n24382), .CK(clk), .Q(\mem[215][4] ) );
  DFF_X1 \mem_reg[215][3]  ( .D(n24383), .CK(clk), .Q(\mem[215][3] ) );
  DFF_X1 \mem_reg[215][2]  ( .D(n24384), .CK(clk), .Q(\mem[215][2] ) );
  DFF_X1 \mem_reg[215][1]  ( .D(n24385), .CK(clk), .Q(\mem[215][1] ) );
  DFF_X1 \mem_reg[215][0]  ( .D(n24386), .CK(clk), .Q(\mem[215][0] ) );
  DFF_X1 \mem_reg[214][7]  ( .D(n24387), .CK(clk), .Q(\mem[214][7] ) );
  DFF_X1 \mem_reg[214][6]  ( .D(n24388), .CK(clk), .Q(\mem[214][6] ) );
  DFF_X1 \mem_reg[214][5]  ( .D(n24389), .CK(clk), .Q(\mem[214][5] ) );
  DFF_X1 \mem_reg[214][4]  ( .D(n24390), .CK(clk), .Q(\mem[214][4] ) );
  DFF_X1 \mem_reg[214][3]  ( .D(n24391), .CK(clk), .Q(\mem[214][3] ) );
  DFF_X1 \mem_reg[214][2]  ( .D(n24392), .CK(clk), .Q(\mem[214][2] ) );
  DFF_X1 \mem_reg[214][1]  ( .D(n24393), .CK(clk), .Q(\mem[214][1] ) );
  DFF_X1 \mem_reg[214][0]  ( .D(n24394), .CK(clk), .Q(\mem[214][0] ) );
  DFF_X1 \mem_reg[213][7]  ( .D(n24395), .CK(clk), .Q(\mem[213][7] ) );
  DFF_X1 \mem_reg[213][6]  ( .D(n24396), .CK(clk), .Q(\mem[213][6] ) );
  DFF_X1 \mem_reg[213][5]  ( .D(n24397), .CK(clk), .Q(\mem[213][5] ) );
  DFF_X1 \mem_reg[213][4]  ( .D(n24398), .CK(clk), .Q(\mem[213][4] ) );
  DFF_X1 \mem_reg[213][3]  ( .D(n24399), .CK(clk), .Q(\mem[213][3] ) );
  DFF_X1 \mem_reg[213][2]  ( .D(n24400), .CK(clk), .Q(\mem[213][2] ) );
  DFF_X1 \mem_reg[213][1]  ( .D(n24401), .CK(clk), .Q(\mem[213][1] ) );
  DFF_X1 \mem_reg[213][0]  ( .D(n24402), .CK(clk), .Q(\mem[213][0] ) );
  DFF_X1 \mem_reg[212][7]  ( .D(n24403), .CK(clk), .Q(\mem[212][7] ) );
  DFF_X1 \mem_reg[212][6]  ( .D(n24404), .CK(clk), .Q(\mem[212][6] ) );
  DFF_X1 \mem_reg[212][5]  ( .D(n24405), .CK(clk), .Q(\mem[212][5] ) );
  DFF_X1 \mem_reg[212][4]  ( .D(n24406), .CK(clk), .Q(\mem[212][4] ) );
  DFF_X1 \mem_reg[212][3]  ( .D(n24407), .CK(clk), .Q(\mem[212][3] ) );
  DFF_X1 \mem_reg[212][2]  ( .D(n24408), .CK(clk), .Q(\mem[212][2] ) );
  DFF_X1 \mem_reg[212][1]  ( .D(n24409), .CK(clk), .Q(\mem[212][1] ) );
  DFF_X1 \mem_reg[212][0]  ( .D(n24410), .CK(clk), .Q(\mem[212][0] ) );
  DFF_X1 \mem_reg[211][7]  ( .D(n24411), .CK(clk), .Q(\mem[211][7] ) );
  DFF_X1 \mem_reg[211][6]  ( .D(n24412), .CK(clk), .Q(\mem[211][6] ) );
  DFF_X1 \mem_reg[211][5]  ( .D(n24413), .CK(clk), .Q(\mem[211][5] ) );
  DFF_X1 \mem_reg[211][4]  ( .D(n24414), .CK(clk), .Q(\mem[211][4] ) );
  DFF_X1 \mem_reg[211][3]  ( .D(n24415), .CK(clk), .Q(\mem[211][3] ) );
  DFF_X1 \mem_reg[211][2]  ( .D(n24416), .CK(clk), .Q(\mem[211][2] ) );
  DFF_X1 \mem_reg[211][1]  ( .D(n24417), .CK(clk), .Q(\mem[211][1] ) );
  DFF_X1 \mem_reg[211][0]  ( .D(n24418), .CK(clk), .Q(\mem[211][0] ) );
  DFF_X1 \mem_reg[210][7]  ( .D(n24419), .CK(clk), .Q(\mem[210][7] ) );
  DFF_X1 \mem_reg[210][6]  ( .D(n24420), .CK(clk), .Q(\mem[210][6] ) );
  DFF_X1 \mem_reg[210][5]  ( .D(n24421), .CK(clk), .Q(\mem[210][5] ) );
  DFF_X1 \mem_reg[210][4]  ( .D(n24422), .CK(clk), .Q(\mem[210][4] ) );
  DFF_X1 \mem_reg[210][3]  ( .D(n24423), .CK(clk), .Q(\mem[210][3] ) );
  DFF_X1 \mem_reg[210][2]  ( .D(n24424), .CK(clk), .Q(\mem[210][2] ) );
  DFF_X1 \mem_reg[210][1]  ( .D(n24425), .CK(clk), .Q(\mem[210][1] ) );
  DFF_X1 \mem_reg[210][0]  ( .D(n24426), .CK(clk), .Q(\mem[210][0] ) );
  DFF_X1 \mem_reg[209][7]  ( .D(n24427), .CK(clk), .Q(\mem[209][7] ) );
  DFF_X1 \mem_reg[209][6]  ( .D(n24428), .CK(clk), .Q(\mem[209][6] ) );
  DFF_X1 \mem_reg[209][5]  ( .D(n24429), .CK(clk), .Q(\mem[209][5] ) );
  DFF_X1 \mem_reg[209][4]  ( .D(n24430), .CK(clk), .Q(\mem[209][4] ) );
  DFF_X1 \mem_reg[209][3]  ( .D(n24431), .CK(clk), .Q(\mem[209][3] ) );
  DFF_X1 \mem_reg[209][2]  ( .D(n24432), .CK(clk), .Q(\mem[209][2] ) );
  DFF_X1 \mem_reg[209][1]  ( .D(n24433), .CK(clk), .Q(\mem[209][1] ) );
  DFF_X1 \mem_reg[209][0]  ( .D(n24434), .CK(clk), .Q(\mem[209][0] ) );
  DFF_X1 \mem_reg[208][7]  ( .D(n24435), .CK(clk), .Q(\mem[208][7] ) );
  DFF_X1 \mem_reg[208][6]  ( .D(n24436), .CK(clk), .Q(\mem[208][6] ) );
  DFF_X1 \mem_reg[208][5]  ( .D(n24437), .CK(clk), .Q(\mem[208][5] ) );
  DFF_X1 \mem_reg[208][4]  ( .D(n24438), .CK(clk), .Q(\mem[208][4] ) );
  DFF_X1 \mem_reg[208][3]  ( .D(n24439), .CK(clk), .Q(\mem[208][3] ) );
  DFF_X1 \mem_reg[208][2]  ( .D(n24440), .CK(clk), .Q(\mem[208][2] ) );
  DFF_X1 \mem_reg[208][1]  ( .D(n24441), .CK(clk), .Q(\mem[208][1] ) );
  DFF_X1 \mem_reg[208][0]  ( .D(n24442), .CK(clk), .Q(\mem[208][0] ) );
  DFF_X1 \mem_reg[207][7]  ( .D(n24443), .CK(clk), .Q(\mem[207][7] ) );
  DFF_X1 \mem_reg[207][6]  ( .D(n24444), .CK(clk), .Q(\mem[207][6] ) );
  DFF_X1 \mem_reg[207][5]  ( .D(n24445), .CK(clk), .Q(\mem[207][5] ) );
  DFF_X1 \mem_reg[207][4]  ( .D(n24446), .CK(clk), .Q(\mem[207][4] ) );
  DFF_X1 \mem_reg[207][3]  ( .D(n24447), .CK(clk), .Q(\mem[207][3] ) );
  DFF_X1 \mem_reg[207][2]  ( .D(n24448), .CK(clk), .Q(\mem[207][2] ) );
  DFF_X1 \mem_reg[207][1]  ( .D(n24449), .CK(clk), .Q(\mem[207][1] ) );
  DFF_X1 \mem_reg[207][0]  ( .D(n24450), .CK(clk), .Q(\mem[207][0] ) );
  DFF_X1 \mem_reg[206][7]  ( .D(n24451), .CK(clk), .Q(\mem[206][7] ) );
  DFF_X1 \mem_reg[206][6]  ( .D(n24452), .CK(clk), .Q(\mem[206][6] ) );
  DFF_X1 \mem_reg[206][5]  ( .D(n24453), .CK(clk), .Q(\mem[206][5] ) );
  DFF_X1 \mem_reg[206][4]  ( .D(n24454), .CK(clk), .Q(\mem[206][4] ) );
  DFF_X1 \mem_reg[206][3]  ( .D(n24455), .CK(clk), .Q(\mem[206][3] ) );
  DFF_X1 \mem_reg[206][2]  ( .D(n24456), .CK(clk), .Q(\mem[206][2] ) );
  DFF_X1 \mem_reg[206][1]  ( .D(n24457), .CK(clk), .Q(\mem[206][1] ) );
  DFF_X1 \mem_reg[206][0]  ( .D(n24458), .CK(clk), .Q(\mem[206][0] ) );
  DFF_X1 \mem_reg[205][7]  ( .D(n24459), .CK(clk), .Q(\mem[205][7] ) );
  DFF_X1 \mem_reg[205][6]  ( .D(n24460), .CK(clk), .Q(\mem[205][6] ) );
  DFF_X1 \mem_reg[205][5]  ( .D(n24461), .CK(clk), .Q(\mem[205][5] ) );
  DFF_X1 \mem_reg[205][4]  ( .D(n24462), .CK(clk), .Q(\mem[205][4] ) );
  DFF_X1 \mem_reg[205][3]  ( .D(n24463), .CK(clk), .Q(\mem[205][3] ) );
  DFF_X1 \mem_reg[205][2]  ( .D(n24464), .CK(clk), .Q(\mem[205][2] ) );
  DFF_X1 \mem_reg[205][1]  ( .D(n24465), .CK(clk), .Q(\mem[205][1] ) );
  DFF_X1 \mem_reg[205][0]  ( .D(n24466), .CK(clk), .Q(\mem[205][0] ) );
  DFF_X1 \mem_reg[204][7]  ( .D(n24467), .CK(clk), .Q(\mem[204][7] ) );
  DFF_X1 \mem_reg[204][6]  ( .D(n24468), .CK(clk), .Q(\mem[204][6] ) );
  DFF_X1 \mem_reg[204][5]  ( .D(n24469), .CK(clk), .Q(\mem[204][5] ) );
  DFF_X1 \mem_reg[204][4]  ( .D(n24470), .CK(clk), .Q(\mem[204][4] ) );
  DFF_X1 \mem_reg[204][3]  ( .D(n24471), .CK(clk), .Q(\mem[204][3] ) );
  DFF_X1 \mem_reg[204][2]  ( .D(n24472), .CK(clk), .Q(\mem[204][2] ) );
  DFF_X1 \mem_reg[204][1]  ( .D(n24473), .CK(clk), .Q(\mem[204][1] ) );
  DFF_X1 \mem_reg[204][0]  ( .D(n24474), .CK(clk), .Q(\mem[204][0] ) );
  DFF_X1 \mem_reg[203][7]  ( .D(n24475), .CK(clk), .Q(\mem[203][7] ) );
  DFF_X1 \mem_reg[203][6]  ( .D(n24476), .CK(clk), .Q(\mem[203][6] ) );
  DFF_X1 \mem_reg[203][5]  ( .D(n24477), .CK(clk), .Q(\mem[203][5] ) );
  DFF_X1 \mem_reg[203][4]  ( .D(n24478), .CK(clk), .Q(\mem[203][4] ) );
  DFF_X1 \mem_reg[203][3]  ( .D(n24479), .CK(clk), .Q(\mem[203][3] ) );
  DFF_X1 \mem_reg[203][2]  ( .D(n24480), .CK(clk), .Q(\mem[203][2] ) );
  DFF_X1 \mem_reg[203][1]  ( .D(n24481), .CK(clk), .Q(\mem[203][1] ) );
  DFF_X1 \mem_reg[203][0]  ( .D(n24482), .CK(clk), .Q(\mem[203][0] ) );
  DFF_X1 \mem_reg[202][7]  ( .D(n24483), .CK(clk), .Q(\mem[202][7] ) );
  DFF_X1 \mem_reg[202][6]  ( .D(n24484), .CK(clk), .Q(\mem[202][6] ) );
  DFF_X1 \mem_reg[202][5]  ( .D(n24485), .CK(clk), .Q(\mem[202][5] ) );
  DFF_X1 \mem_reg[202][4]  ( .D(n24486), .CK(clk), .Q(\mem[202][4] ) );
  DFF_X1 \mem_reg[202][3]  ( .D(n24487), .CK(clk), .Q(\mem[202][3] ) );
  DFF_X1 \mem_reg[202][2]  ( .D(n24488), .CK(clk), .Q(\mem[202][2] ) );
  DFF_X1 \mem_reg[202][1]  ( .D(n24489), .CK(clk), .Q(\mem[202][1] ) );
  DFF_X1 \mem_reg[202][0]  ( .D(n24490), .CK(clk), .Q(\mem[202][0] ) );
  DFF_X1 \mem_reg[201][7]  ( .D(n24491), .CK(clk), .Q(\mem[201][7] ) );
  DFF_X1 \mem_reg[201][6]  ( .D(n24492), .CK(clk), .Q(\mem[201][6] ) );
  DFF_X1 \mem_reg[201][5]  ( .D(n24493), .CK(clk), .Q(\mem[201][5] ) );
  DFF_X1 \mem_reg[201][4]  ( .D(n24494), .CK(clk), .Q(\mem[201][4] ) );
  DFF_X1 \mem_reg[201][3]  ( .D(n24495), .CK(clk), .Q(\mem[201][3] ) );
  DFF_X1 \mem_reg[201][2]  ( .D(n24496), .CK(clk), .Q(\mem[201][2] ) );
  DFF_X1 \mem_reg[201][1]  ( .D(n24497), .CK(clk), .Q(\mem[201][1] ) );
  DFF_X1 \mem_reg[201][0]  ( .D(n24498), .CK(clk), .Q(\mem[201][0] ) );
  DFF_X1 \mem_reg[200][7]  ( .D(n24499), .CK(clk), .Q(\mem[200][7] ) );
  DFF_X1 \mem_reg[200][6]  ( .D(n24500), .CK(clk), .Q(\mem[200][6] ) );
  DFF_X1 \mem_reg[200][5]  ( .D(n24501), .CK(clk), .Q(\mem[200][5] ) );
  DFF_X1 \mem_reg[200][4]  ( .D(n24502), .CK(clk), .Q(\mem[200][4] ) );
  DFF_X1 \mem_reg[200][3]  ( .D(n24503), .CK(clk), .Q(\mem[200][3] ) );
  DFF_X1 \mem_reg[200][2]  ( .D(n24504), .CK(clk), .Q(\mem[200][2] ) );
  DFF_X1 \mem_reg[200][1]  ( .D(n24505), .CK(clk), .Q(\mem[200][1] ) );
  DFF_X1 \mem_reg[200][0]  ( .D(n24506), .CK(clk), .Q(\mem[200][0] ) );
  DFF_X1 \mem_reg[199][7]  ( .D(n24507), .CK(clk), .Q(\mem[199][7] ) );
  DFF_X1 \mem_reg[199][6]  ( .D(n24508), .CK(clk), .Q(\mem[199][6] ) );
  DFF_X1 \mem_reg[199][5]  ( .D(n24509), .CK(clk), .Q(\mem[199][5] ) );
  DFF_X1 \mem_reg[199][4]  ( .D(n24510), .CK(clk), .Q(\mem[199][4] ) );
  DFF_X1 \mem_reg[199][3]  ( .D(n24511), .CK(clk), .Q(\mem[199][3] ) );
  DFF_X1 \mem_reg[199][2]  ( .D(n24512), .CK(clk), .Q(\mem[199][2] ) );
  DFF_X1 \mem_reg[199][1]  ( .D(n24513), .CK(clk), .Q(\mem[199][1] ) );
  DFF_X1 \mem_reg[199][0]  ( .D(n24514), .CK(clk), .Q(\mem[199][0] ) );
  DFF_X1 \mem_reg[198][7]  ( .D(n24515), .CK(clk), .Q(\mem[198][7] ) );
  DFF_X1 \mem_reg[198][6]  ( .D(n24516), .CK(clk), .Q(\mem[198][6] ) );
  DFF_X1 \mem_reg[198][5]  ( .D(n24517), .CK(clk), .Q(\mem[198][5] ) );
  DFF_X1 \mem_reg[198][4]  ( .D(n24518), .CK(clk), .Q(\mem[198][4] ) );
  DFF_X1 \mem_reg[198][3]  ( .D(n24519), .CK(clk), .Q(\mem[198][3] ) );
  DFF_X1 \mem_reg[198][2]  ( .D(n24520), .CK(clk), .Q(\mem[198][2] ) );
  DFF_X1 \mem_reg[198][1]  ( .D(n24521), .CK(clk), .Q(\mem[198][1] ) );
  DFF_X1 \mem_reg[198][0]  ( .D(n24522), .CK(clk), .Q(\mem[198][0] ) );
  DFF_X1 \mem_reg[197][7]  ( .D(n24523), .CK(clk), .Q(\mem[197][7] ) );
  DFF_X1 \mem_reg[197][6]  ( .D(n24524), .CK(clk), .Q(\mem[197][6] ) );
  DFF_X1 \mem_reg[197][5]  ( .D(n24525), .CK(clk), .Q(\mem[197][5] ) );
  DFF_X1 \mem_reg[197][4]  ( .D(n24526), .CK(clk), .Q(\mem[197][4] ) );
  DFF_X1 \mem_reg[197][3]  ( .D(n24527), .CK(clk), .Q(\mem[197][3] ) );
  DFF_X1 \mem_reg[197][2]  ( .D(n24528), .CK(clk), .Q(\mem[197][2] ) );
  DFF_X1 \mem_reg[197][1]  ( .D(n24529), .CK(clk), .Q(\mem[197][1] ) );
  DFF_X1 \mem_reg[197][0]  ( .D(n24530), .CK(clk), .Q(\mem[197][0] ) );
  DFF_X1 \mem_reg[196][7]  ( .D(n24531), .CK(clk), .Q(\mem[196][7] ) );
  DFF_X1 \mem_reg[196][6]  ( .D(n24532), .CK(clk), .Q(\mem[196][6] ) );
  DFF_X1 \mem_reg[196][5]  ( .D(n24533), .CK(clk), .Q(\mem[196][5] ) );
  DFF_X1 \mem_reg[196][4]  ( .D(n24534), .CK(clk), .Q(\mem[196][4] ) );
  DFF_X1 \mem_reg[196][3]  ( .D(n24535), .CK(clk), .Q(\mem[196][3] ) );
  DFF_X1 \mem_reg[196][2]  ( .D(n24536), .CK(clk), .Q(\mem[196][2] ) );
  DFF_X1 \mem_reg[196][1]  ( .D(n24537), .CK(clk), .Q(\mem[196][1] ) );
  DFF_X1 \mem_reg[196][0]  ( .D(n24538), .CK(clk), .Q(\mem[196][0] ) );
  DFF_X1 \mem_reg[195][7]  ( .D(n24539), .CK(clk), .Q(\mem[195][7] ) );
  DFF_X1 \mem_reg[195][6]  ( .D(n24540), .CK(clk), .Q(\mem[195][6] ) );
  DFF_X1 \mem_reg[195][5]  ( .D(n24541), .CK(clk), .Q(\mem[195][5] ) );
  DFF_X1 \mem_reg[195][4]  ( .D(n24542), .CK(clk), .Q(\mem[195][4] ) );
  DFF_X1 \mem_reg[195][3]  ( .D(n24543), .CK(clk), .Q(\mem[195][3] ) );
  DFF_X1 \mem_reg[195][2]  ( .D(n24544), .CK(clk), .Q(\mem[195][2] ) );
  DFF_X1 \mem_reg[195][1]  ( .D(n24545), .CK(clk), .Q(\mem[195][1] ) );
  DFF_X1 \mem_reg[195][0]  ( .D(n24546), .CK(clk), .Q(\mem[195][0] ) );
  DFF_X1 \mem_reg[194][7]  ( .D(n24547), .CK(clk), .Q(\mem[194][7] ) );
  DFF_X1 \mem_reg[194][6]  ( .D(n24548), .CK(clk), .Q(\mem[194][6] ) );
  DFF_X1 \mem_reg[194][5]  ( .D(n24549), .CK(clk), .Q(\mem[194][5] ) );
  DFF_X1 \mem_reg[194][4]  ( .D(n24550), .CK(clk), .Q(\mem[194][4] ) );
  DFF_X1 \mem_reg[194][3]  ( .D(n24551), .CK(clk), .Q(\mem[194][3] ) );
  DFF_X1 \mem_reg[194][2]  ( .D(n24552), .CK(clk), .Q(\mem[194][2] ) );
  DFF_X1 \mem_reg[194][1]  ( .D(n24553), .CK(clk), .Q(\mem[194][1] ) );
  DFF_X1 \mem_reg[194][0]  ( .D(n24554), .CK(clk), .Q(\mem[194][0] ) );
  DFF_X1 \mem_reg[193][7]  ( .D(n24555), .CK(clk), .Q(\mem[193][7] ) );
  DFF_X1 \mem_reg[193][6]  ( .D(n24556), .CK(clk), .Q(\mem[193][6] ) );
  DFF_X1 \mem_reg[193][5]  ( .D(n24557), .CK(clk), .Q(\mem[193][5] ) );
  DFF_X1 \mem_reg[193][4]  ( .D(n24558), .CK(clk), .Q(\mem[193][4] ) );
  DFF_X1 \mem_reg[193][3]  ( .D(n24559), .CK(clk), .Q(\mem[193][3] ) );
  DFF_X1 \mem_reg[193][2]  ( .D(n24560), .CK(clk), .Q(\mem[193][2] ) );
  DFF_X1 \mem_reg[193][1]  ( .D(n24561), .CK(clk), .Q(\mem[193][1] ) );
  DFF_X1 \mem_reg[193][0]  ( .D(n24562), .CK(clk), .Q(\mem[193][0] ) );
  DFF_X1 \mem_reg[192][7]  ( .D(n24563), .CK(clk), .Q(\mem[192][7] ) );
  DFF_X1 \mem_reg[192][6]  ( .D(n24564), .CK(clk), .Q(\mem[192][6] ) );
  DFF_X1 \mem_reg[192][5]  ( .D(n24565), .CK(clk), .Q(\mem[192][5] ) );
  DFF_X1 \mem_reg[192][4]  ( .D(n24566), .CK(clk), .Q(\mem[192][4] ) );
  DFF_X1 \mem_reg[192][3]  ( .D(n24567), .CK(clk), .Q(\mem[192][3] ) );
  DFF_X1 \mem_reg[192][2]  ( .D(n24568), .CK(clk), .Q(\mem[192][2] ) );
  DFF_X1 \mem_reg[192][1]  ( .D(n24569), .CK(clk), .Q(\mem[192][1] ) );
  DFF_X1 \mem_reg[192][0]  ( .D(n24570), .CK(clk), .Q(\mem[192][0] ) );
  DFF_X1 \mem_reg[191][7]  ( .D(n24571), .CK(clk), .Q(\mem[191][7] ) );
  DFF_X1 \mem_reg[191][6]  ( .D(n24572), .CK(clk), .Q(\mem[191][6] ) );
  DFF_X1 \mem_reg[191][5]  ( .D(n24573), .CK(clk), .Q(\mem[191][5] ) );
  DFF_X1 \mem_reg[191][4]  ( .D(n24574), .CK(clk), .Q(\mem[191][4] ) );
  DFF_X1 \mem_reg[191][3]  ( .D(n24575), .CK(clk), .Q(\mem[191][3] ) );
  DFF_X1 \mem_reg[191][2]  ( .D(n24576), .CK(clk), .Q(\mem[191][2] ) );
  DFF_X1 \mem_reg[191][1]  ( .D(n24577), .CK(clk), .Q(\mem[191][1] ) );
  DFF_X1 \mem_reg[191][0]  ( .D(n24578), .CK(clk), .Q(\mem[191][0] ) );
  DFF_X1 \mem_reg[190][7]  ( .D(n24579), .CK(clk), .Q(\mem[190][7] ) );
  DFF_X1 \mem_reg[190][6]  ( .D(n24580), .CK(clk), .Q(\mem[190][6] ) );
  DFF_X1 \mem_reg[190][5]  ( .D(n24581), .CK(clk), .Q(\mem[190][5] ) );
  DFF_X1 \mem_reg[190][4]  ( .D(n24582), .CK(clk), .Q(\mem[190][4] ) );
  DFF_X1 \mem_reg[190][3]  ( .D(n24583), .CK(clk), .Q(\mem[190][3] ) );
  DFF_X1 \mem_reg[190][2]  ( .D(n24584), .CK(clk), .Q(\mem[190][2] ) );
  DFF_X1 \mem_reg[190][1]  ( .D(n24585), .CK(clk), .Q(\mem[190][1] ) );
  DFF_X1 \mem_reg[190][0]  ( .D(n24586), .CK(clk), .Q(\mem[190][0] ) );
  DFF_X1 \mem_reg[189][7]  ( .D(n24587), .CK(clk), .Q(\mem[189][7] ) );
  DFF_X1 \mem_reg[189][6]  ( .D(n24588), .CK(clk), .Q(\mem[189][6] ) );
  DFF_X1 \mem_reg[189][5]  ( .D(n24589), .CK(clk), .Q(\mem[189][5] ) );
  DFF_X1 \mem_reg[189][4]  ( .D(n24590), .CK(clk), .Q(\mem[189][4] ) );
  DFF_X1 \mem_reg[189][3]  ( .D(n24591), .CK(clk), .Q(\mem[189][3] ) );
  DFF_X1 \mem_reg[189][2]  ( .D(n24592), .CK(clk), .Q(\mem[189][2] ) );
  DFF_X1 \mem_reg[189][1]  ( .D(n24593), .CK(clk), .Q(\mem[189][1] ) );
  DFF_X1 \mem_reg[189][0]  ( .D(n24594), .CK(clk), .Q(\mem[189][0] ) );
  DFF_X1 \mem_reg[188][7]  ( .D(n24595), .CK(clk), .Q(\mem[188][7] ) );
  DFF_X1 \mem_reg[188][6]  ( .D(n24596), .CK(clk), .Q(\mem[188][6] ) );
  DFF_X1 \mem_reg[188][5]  ( .D(n24597), .CK(clk), .Q(\mem[188][5] ) );
  DFF_X1 \mem_reg[188][4]  ( .D(n24598), .CK(clk), .Q(\mem[188][4] ) );
  DFF_X1 \mem_reg[188][3]  ( .D(n24599), .CK(clk), .Q(\mem[188][3] ) );
  DFF_X1 \mem_reg[188][2]  ( .D(n24600), .CK(clk), .Q(\mem[188][2] ) );
  DFF_X1 \mem_reg[188][1]  ( .D(n24601), .CK(clk), .Q(\mem[188][1] ) );
  DFF_X1 \mem_reg[188][0]  ( .D(n24602), .CK(clk), .Q(\mem[188][0] ) );
  DFF_X1 \mem_reg[187][7]  ( .D(n24603), .CK(clk), .Q(\mem[187][7] ) );
  DFF_X1 \mem_reg[187][6]  ( .D(n24604), .CK(clk), .Q(\mem[187][6] ) );
  DFF_X1 \mem_reg[187][5]  ( .D(n24605), .CK(clk), .Q(\mem[187][5] ) );
  DFF_X1 \mem_reg[187][4]  ( .D(n24606), .CK(clk), .Q(\mem[187][4] ) );
  DFF_X1 \mem_reg[187][3]  ( .D(n24607), .CK(clk), .Q(\mem[187][3] ) );
  DFF_X1 \mem_reg[187][2]  ( .D(n24608), .CK(clk), .Q(\mem[187][2] ) );
  DFF_X1 \mem_reg[187][1]  ( .D(n24609), .CK(clk), .Q(\mem[187][1] ) );
  DFF_X1 \mem_reg[187][0]  ( .D(n24610), .CK(clk), .Q(\mem[187][0] ) );
  DFF_X1 \mem_reg[186][7]  ( .D(n24611), .CK(clk), .Q(\mem[186][7] ) );
  DFF_X1 \mem_reg[186][6]  ( .D(n24612), .CK(clk), .Q(\mem[186][6] ) );
  DFF_X1 \mem_reg[186][5]  ( .D(n24613), .CK(clk), .Q(\mem[186][5] ) );
  DFF_X1 \mem_reg[186][4]  ( .D(n24614), .CK(clk), .Q(\mem[186][4] ) );
  DFF_X1 \mem_reg[186][3]  ( .D(n24615), .CK(clk), .Q(\mem[186][3] ) );
  DFF_X1 \mem_reg[186][2]  ( .D(n24616), .CK(clk), .Q(\mem[186][2] ) );
  DFF_X1 \mem_reg[186][1]  ( .D(n24617), .CK(clk), .Q(\mem[186][1] ) );
  DFF_X1 \mem_reg[186][0]  ( .D(n24618), .CK(clk), .Q(\mem[186][0] ) );
  DFF_X1 \mem_reg[185][7]  ( .D(n24619), .CK(clk), .Q(\mem[185][7] ) );
  DFF_X1 \mem_reg[185][6]  ( .D(n24620), .CK(clk), .Q(\mem[185][6] ) );
  DFF_X1 \mem_reg[185][5]  ( .D(n24621), .CK(clk), .Q(\mem[185][5] ) );
  DFF_X1 \mem_reg[185][4]  ( .D(n24622), .CK(clk), .Q(\mem[185][4] ) );
  DFF_X1 \mem_reg[185][3]  ( .D(n24623), .CK(clk), .Q(\mem[185][3] ) );
  DFF_X1 \mem_reg[185][2]  ( .D(n24624), .CK(clk), .Q(\mem[185][2] ) );
  DFF_X1 \mem_reg[185][1]  ( .D(n24625), .CK(clk), .Q(\mem[185][1] ) );
  DFF_X1 \mem_reg[185][0]  ( .D(n24626), .CK(clk), .Q(\mem[185][0] ) );
  DFF_X1 \mem_reg[184][7]  ( .D(n24627), .CK(clk), .Q(\mem[184][7] ) );
  DFF_X1 \mem_reg[184][6]  ( .D(n24628), .CK(clk), .Q(\mem[184][6] ) );
  DFF_X1 \mem_reg[184][5]  ( .D(n24629), .CK(clk), .Q(\mem[184][5] ) );
  DFF_X1 \mem_reg[184][4]  ( .D(n24630), .CK(clk), .Q(\mem[184][4] ) );
  DFF_X1 \mem_reg[184][3]  ( .D(n24631), .CK(clk), .Q(\mem[184][3] ) );
  DFF_X1 \mem_reg[184][2]  ( .D(n24632), .CK(clk), .Q(\mem[184][2] ) );
  DFF_X1 \mem_reg[184][1]  ( .D(n24633), .CK(clk), .Q(\mem[184][1] ) );
  DFF_X1 \mem_reg[184][0]  ( .D(n24634), .CK(clk), .Q(\mem[184][0] ) );
  DFF_X1 \mem_reg[183][7]  ( .D(n24635), .CK(clk), .Q(\mem[183][7] ) );
  DFF_X1 \mem_reg[183][6]  ( .D(n24636), .CK(clk), .Q(\mem[183][6] ) );
  DFF_X1 \mem_reg[183][5]  ( .D(n24637), .CK(clk), .Q(\mem[183][5] ) );
  DFF_X1 \mem_reg[183][4]  ( .D(n24638), .CK(clk), .Q(\mem[183][4] ) );
  DFF_X1 \mem_reg[183][3]  ( .D(n24639), .CK(clk), .Q(\mem[183][3] ) );
  DFF_X1 \mem_reg[183][2]  ( .D(n24640), .CK(clk), .Q(\mem[183][2] ) );
  DFF_X1 \mem_reg[183][1]  ( .D(n24641), .CK(clk), .Q(\mem[183][1] ) );
  DFF_X1 \mem_reg[183][0]  ( .D(n24642), .CK(clk), .Q(\mem[183][0] ) );
  DFF_X1 \mem_reg[182][7]  ( .D(n24643), .CK(clk), .Q(\mem[182][7] ) );
  DFF_X1 \mem_reg[182][6]  ( .D(n24644), .CK(clk), .Q(\mem[182][6] ) );
  DFF_X1 \mem_reg[182][5]  ( .D(n24645), .CK(clk), .Q(\mem[182][5] ) );
  DFF_X1 \mem_reg[182][4]  ( .D(n24646), .CK(clk), .Q(\mem[182][4] ) );
  DFF_X1 \mem_reg[182][3]  ( .D(n24647), .CK(clk), .Q(\mem[182][3] ) );
  DFF_X1 \mem_reg[182][2]  ( .D(n24648), .CK(clk), .Q(\mem[182][2] ) );
  DFF_X1 \mem_reg[182][1]  ( .D(n24649), .CK(clk), .Q(\mem[182][1] ) );
  DFF_X1 \mem_reg[182][0]  ( .D(n24650), .CK(clk), .Q(\mem[182][0] ) );
  DFF_X1 \mem_reg[181][7]  ( .D(n24651), .CK(clk), .Q(\mem[181][7] ) );
  DFF_X1 \mem_reg[181][6]  ( .D(n24652), .CK(clk), .Q(\mem[181][6] ) );
  DFF_X1 \mem_reg[181][5]  ( .D(n24653), .CK(clk), .Q(\mem[181][5] ) );
  DFF_X1 \mem_reg[181][4]  ( .D(n24654), .CK(clk), .Q(\mem[181][4] ) );
  DFF_X1 \mem_reg[181][3]  ( .D(n24655), .CK(clk), .Q(\mem[181][3] ) );
  DFF_X1 \mem_reg[181][2]  ( .D(n24656), .CK(clk), .Q(\mem[181][2] ) );
  DFF_X1 \mem_reg[181][1]  ( .D(n24657), .CK(clk), .Q(\mem[181][1] ) );
  DFF_X1 \mem_reg[181][0]  ( .D(n24658), .CK(clk), .Q(\mem[181][0] ) );
  DFF_X1 \mem_reg[180][7]  ( .D(n24659), .CK(clk), .Q(\mem[180][7] ) );
  DFF_X1 \mem_reg[180][6]  ( .D(n24660), .CK(clk), .Q(\mem[180][6] ) );
  DFF_X1 \mem_reg[180][5]  ( .D(n24661), .CK(clk), .Q(\mem[180][5] ) );
  DFF_X1 \mem_reg[180][4]  ( .D(n24662), .CK(clk), .Q(\mem[180][4] ) );
  DFF_X1 \mem_reg[180][3]  ( .D(n24663), .CK(clk), .Q(\mem[180][3] ) );
  DFF_X1 \mem_reg[180][2]  ( .D(n24664), .CK(clk), .Q(\mem[180][2] ) );
  DFF_X1 \mem_reg[180][1]  ( .D(n24665), .CK(clk), .Q(\mem[180][1] ) );
  DFF_X1 \mem_reg[180][0]  ( .D(n24666), .CK(clk), .Q(\mem[180][0] ) );
  DFF_X1 \mem_reg[179][7]  ( .D(n24667), .CK(clk), .Q(\mem[179][7] ) );
  DFF_X1 \mem_reg[179][6]  ( .D(n24668), .CK(clk), .Q(\mem[179][6] ) );
  DFF_X1 \mem_reg[179][5]  ( .D(n24669), .CK(clk), .Q(\mem[179][5] ) );
  DFF_X1 \mem_reg[179][4]  ( .D(n24670), .CK(clk), .Q(\mem[179][4] ) );
  DFF_X1 \mem_reg[179][3]  ( .D(n24671), .CK(clk), .Q(\mem[179][3] ) );
  DFF_X1 \mem_reg[179][2]  ( .D(n24672), .CK(clk), .Q(\mem[179][2] ) );
  DFF_X1 \mem_reg[179][1]  ( .D(n24673), .CK(clk), .Q(\mem[179][1] ) );
  DFF_X1 \mem_reg[179][0]  ( .D(n24674), .CK(clk), .Q(\mem[179][0] ) );
  DFF_X1 \mem_reg[178][7]  ( .D(n24675), .CK(clk), .Q(\mem[178][7] ) );
  DFF_X1 \mem_reg[178][6]  ( .D(n24676), .CK(clk), .Q(\mem[178][6] ) );
  DFF_X1 \mem_reg[178][5]  ( .D(n24677), .CK(clk), .Q(\mem[178][5] ) );
  DFF_X1 \mem_reg[178][4]  ( .D(n24678), .CK(clk), .Q(\mem[178][4] ) );
  DFF_X1 \mem_reg[178][3]  ( .D(n24679), .CK(clk), .Q(\mem[178][3] ) );
  DFF_X1 \mem_reg[178][2]  ( .D(n24680), .CK(clk), .Q(\mem[178][2] ) );
  DFF_X1 \mem_reg[178][1]  ( .D(n24681), .CK(clk), .Q(\mem[178][1] ) );
  DFF_X1 \mem_reg[178][0]  ( .D(n24682), .CK(clk), .Q(\mem[178][0] ) );
  DFF_X1 \mem_reg[177][7]  ( .D(n24683), .CK(clk), .Q(\mem[177][7] ) );
  DFF_X1 \mem_reg[177][6]  ( .D(n24684), .CK(clk), .Q(\mem[177][6] ) );
  DFF_X1 \mem_reg[177][5]  ( .D(n24685), .CK(clk), .Q(\mem[177][5] ) );
  DFF_X1 \mem_reg[177][4]  ( .D(n24686), .CK(clk), .Q(\mem[177][4] ) );
  DFF_X1 \mem_reg[177][3]  ( .D(n24687), .CK(clk), .Q(\mem[177][3] ) );
  DFF_X1 \mem_reg[177][2]  ( .D(n24688), .CK(clk), .Q(\mem[177][2] ) );
  DFF_X1 \mem_reg[177][1]  ( .D(n24689), .CK(clk), .Q(\mem[177][1] ) );
  DFF_X1 \mem_reg[177][0]  ( .D(n24690), .CK(clk), .Q(\mem[177][0] ) );
  DFF_X1 \mem_reg[176][7]  ( .D(n24691), .CK(clk), .Q(\mem[176][7] ) );
  DFF_X1 \mem_reg[176][6]  ( .D(n24692), .CK(clk), .Q(\mem[176][6] ) );
  DFF_X1 \mem_reg[176][5]  ( .D(n24693), .CK(clk), .Q(\mem[176][5] ) );
  DFF_X1 \mem_reg[176][4]  ( .D(n24694), .CK(clk), .Q(\mem[176][4] ) );
  DFF_X1 \mem_reg[176][3]  ( .D(n24695), .CK(clk), .Q(\mem[176][3] ) );
  DFF_X1 \mem_reg[176][2]  ( .D(n24696), .CK(clk), .Q(\mem[176][2] ) );
  DFF_X1 \mem_reg[176][1]  ( .D(n24697), .CK(clk), .Q(\mem[176][1] ) );
  DFF_X1 \mem_reg[176][0]  ( .D(n24698), .CK(clk), .Q(\mem[176][0] ) );
  DFF_X1 \mem_reg[175][7]  ( .D(n24699), .CK(clk), .Q(\mem[175][7] ) );
  DFF_X1 \mem_reg[175][6]  ( .D(n24700), .CK(clk), .Q(\mem[175][6] ) );
  DFF_X1 \mem_reg[175][5]  ( .D(n24701), .CK(clk), .Q(\mem[175][5] ) );
  DFF_X1 \mem_reg[175][4]  ( .D(n24702), .CK(clk), .Q(\mem[175][4] ) );
  DFF_X1 \mem_reg[175][3]  ( .D(n24703), .CK(clk), .Q(\mem[175][3] ) );
  DFF_X1 \mem_reg[175][2]  ( .D(n24704), .CK(clk), .Q(\mem[175][2] ) );
  DFF_X1 \mem_reg[175][1]  ( .D(n24705), .CK(clk), .Q(\mem[175][1] ) );
  DFF_X1 \mem_reg[175][0]  ( .D(n24706), .CK(clk), .Q(\mem[175][0] ) );
  DFF_X1 \mem_reg[174][7]  ( .D(n24707), .CK(clk), .Q(\mem[174][7] ) );
  DFF_X1 \mem_reg[174][6]  ( .D(n24708), .CK(clk), .Q(\mem[174][6] ) );
  DFF_X1 \mem_reg[174][5]  ( .D(n24709), .CK(clk), .Q(\mem[174][5] ) );
  DFF_X1 \mem_reg[174][4]  ( .D(n24710), .CK(clk), .Q(\mem[174][4] ) );
  DFF_X1 \mem_reg[174][3]  ( .D(n24711), .CK(clk), .Q(\mem[174][3] ) );
  DFF_X1 \mem_reg[174][2]  ( .D(n24712), .CK(clk), .Q(\mem[174][2] ) );
  DFF_X1 \mem_reg[174][1]  ( .D(n24713), .CK(clk), .Q(\mem[174][1] ) );
  DFF_X1 \mem_reg[174][0]  ( .D(n24714), .CK(clk), .Q(\mem[174][0] ) );
  DFF_X1 \mem_reg[173][7]  ( .D(n24715), .CK(clk), .Q(\mem[173][7] ) );
  DFF_X1 \mem_reg[173][6]  ( .D(n24716), .CK(clk), .Q(\mem[173][6] ) );
  DFF_X1 \mem_reg[173][5]  ( .D(n24717), .CK(clk), .Q(\mem[173][5] ) );
  DFF_X1 \mem_reg[173][4]  ( .D(n24718), .CK(clk), .Q(\mem[173][4] ) );
  DFF_X1 \mem_reg[173][3]  ( .D(n24719), .CK(clk), .Q(\mem[173][3] ) );
  DFF_X1 \mem_reg[173][2]  ( .D(n24720), .CK(clk), .Q(\mem[173][2] ) );
  DFF_X1 \mem_reg[173][1]  ( .D(n24721), .CK(clk), .Q(\mem[173][1] ) );
  DFF_X1 \mem_reg[173][0]  ( .D(n24722), .CK(clk), .Q(\mem[173][0] ) );
  DFF_X1 \mem_reg[172][7]  ( .D(n24723), .CK(clk), .Q(\mem[172][7] ) );
  DFF_X1 \mem_reg[172][6]  ( .D(n24724), .CK(clk), .Q(\mem[172][6] ) );
  DFF_X1 \mem_reg[172][5]  ( .D(n24725), .CK(clk), .Q(\mem[172][5] ) );
  DFF_X1 \mem_reg[172][4]  ( .D(n24726), .CK(clk), .Q(\mem[172][4] ) );
  DFF_X1 \mem_reg[172][3]  ( .D(n24727), .CK(clk), .Q(\mem[172][3] ) );
  DFF_X1 \mem_reg[172][2]  ( .D(n24728), .CK(clk), .Q(\mem[172][2] ) );
  DFF_X1 \mem_reg[172][1]  ( .D(n24729), .CK(clk), .Q(\mem[172][1] ) );
  DFF_X1 \mem_reg[172][0]  ( .D(n24730), .CK(clk), .Q(\mem[172][0] ) );
  DFF_X1 \mem_reg[171][7]  ( .D(n24731), .CK(clk), .Q(\mem[171][7] ) );
  DFF_X1 \mem_reg[171][6]  ( .D(n24732), .CK(clk), .Q(\mem[171][6] ) );
  DFF_X1 \mem_reg[171][5]  ( .D(n24733), .CK(clk), .Q(\mem[171][5] ) );
  DFF_X1 \mem_reg[171][4]  ( .D(n24734), .CK(clk), .Q(\mem[171][4] ) );
  DFF_X1 \mem_reg[171][3]  ( .D(n24735), .CK(clk), .Q(\mem[171][3] ) );
  DFF_X1 \mem_reg[171][2]  ( .D(n24736), .CK(clk), .Q(\mem[171][2] ) );
  DFF_X1 \mem_reg[171][1]  ( .D(n24737), .CK(clk), .Q(\mem[171][1] ) );
  DFF_X1 \mem_reg[171][0]  ( .D(n24738), .CK(clk), .Q(\mem[171][0] ) );
  DFF_X1 \mem_reg[170][7]  ( .D(n24739), .CK(clk), .Q(\mem[170][7] ) );
  DFF_X1 \mem_reg[170][6]  ( .D(n24740), .CK(clk), .Q(\mem[170][6] ) );
  DFF_X1 \mem_reg[170][5]  ( .D(n24741), .CK(clk), .Q(\mem[170][5] ) );
  DFF_X1 \mem_reg[170][4]  ( .D(n24742), .CK(clk), .Q(\mem[170][4] ) );
  DFF_X1 \mem_reg[170][3]  ( .D(n24743), .CK(clk), .Q(\mem[170][3] ) );
  DFF_X1 \mem_reg[170][2]  ( .D(n24744), .CK(clk), .Q(\mem[170][2] ) );
  DFF_X1 \mem_reg[170][1]  ( .D(n24745), .CK(clk), .Q(\mem[170][1] ) );
  DFF_X1 \mem_reg[170][0]  ( .D(n24746), .CK(clk), .Q(\mem[170][0] ) );
  DFF_X1 \mem_reg[169][7]  ( .D(n24747), .CK(clk), .Q(\mem[169][7] ) );
  DFF_X1 \mem_reg[169][6]  ( .D(n24748), .CK(clk), .Q(\mem[169][6] ) );
  DFF_X1 \mem_reg[169][5]  ( .D(n24749), .CK(clk), .Q(\mem[169][5] ) );
  DFF_X1 \mem_reg[169][4]  ( .D(n24750), .CK(clk), .Q(\mem[169][4] ) );
  DFF_X1 \mem_reg[169][3]  ( .D(n24751), .CK(clk), .Q(\mem[169][3] ) );
  DFF_X1 \mem_reg[169][2]  ( .D(n24752), .CK(clk), .Q(\mem[169][2] ) );
  DFF_X1 \mem_reg[169][1]  ( .D(n24753), .CK(clk), .Q(\mem[169][1] ) );
  DFF_X1 \mem_reg[169][0]  ( .D(n24754), .CK(clk), .Q(\mem[169][0] ) );
  DFF_X1 \mem_reg[168][7]  ( .D(n24755), .CK(clk), .Q(\mem[168][7] ) );
  DFF_X1 \mem_reg[168][6]  ( .D(n24756), .CK(clk), .Q(\mem[168][6] ) );
  DFF_X1 \mem_reg[168][5]  ( .D(n24757), .CK(clk), .Q(\mem[168][5] ) );
  DFF_X1 \mem_reg[168][4]  ( .D(n24758), .CK(clk), .Q(\mem[168][4] ) );
  DFF_X1 \mem_reg[168][3]  ( .D(n24759), .CK(clk), .Q(\mem[168][3] ) );
  DFF_X1 \mem_reg[168][2]  ( .D(n24760), .CK(clk), .Q(\mem[168][2] ) );
  DFF_X1 \mem_reg[168][1]  ( .D(n24761), .CK(clk), .Q(\mem[168][1] ) );
  DFF_X1 \mem_reg[168][0]  ( .D(n24762), .CK(clk), .Q(\mem[168][0] ) );
  DFF_X1 \mem_reg[167][7]  ( .D(n24763), .CK(clk), .Q(\mem[167][7] ) );
  DFF_X1 \mem_reg[167][6]  ( .D(n24764), .CK(clk), .Q(\mem[167][6] ) );
  DFF_X1 \mem_reg[167][5]  ( .D(n24765), .CK(clk), .Q(\mem[167][5] ) );
  DFF_X1 \mem_reg[167][4]  ( .D(n24766), .CK(clk), .Q(\mem[167][4] ) );
  DFF_X1 \mem_reg[167][3]  ( .D(n24767), .CK(clk), .Q(\mem[167][3] ) );
  DFF_X1 \mem_reg[167][2]  ( .D(n24768), .CK(clk), .Q(\mem[167][2] ) );
  DFF_X1 \mem_reg[167][1]  ( .D(n24769), .CK(clk), .Q(\mem[167][1] ) );
  DFF_X1 \mem_reg[167][0]  ( .D(n24770), .CK(clk), .Q(\mem[167][0] ) );
  DFF_X1 \mem_reg[166][7]  ( .D(n24771), .CK(clk), .Q(\mem[166][7] ) );
  DFF_X1 \mem_reg[166][6]  ( .D(n24772), .CK(clk), .Q(\mem[166][6] ) );
  DFF_X1 \mem_reg[166][5]  ( .D(n24773), .CK(clk), .Q(\mem[166][5] ) );
  DFF_X1 \mem_reg[166][4]  ( .D(n24774), .CK(clk), .Q(\mem[166][4] ) );
  DFF_X1 \mem_reg[166][3]  ( .D(n24775), .CK(clk), .Q(\mem[166][3] ) );
  DFF_X1 \mem_reg[166][2]  ( .D(n24776), .CK(clk), .Q(\mem[166][2] ) );
  DFF_X1 \mem_reg[166][1]  ( .D(n24777), .CK(clk), .Q(\mem[166][1] ) );
  DFF_X1 \mem_reg[166][0]  ( .D(n24778), .CK(clk), .Q(\mem[166][0] ) );
  DFF_X1 \mem_reg[165][7]  ( .D(n24779), .CK(clk), .Q(\mem[165][7] ) );
  DFF_X1 \mem_reg[165][6]  ( .D(n24780), .CK(clk), .Q(\mem[165][6] ) );
  DFF_X1 \mem_reg[165][5]  ( .D(n24781), .CK(clk), .Q(\mem[165][5] ) );
  DFF_X1 \mem_reg[165][4]  ( .D(n24782), .CK(clk), .Q(\mem[165][4] ) );
  DFF_X1 \mem_reg[165][3]  ( .D(n24783), .CK(clk), .Q(\mem[165][3] ) );
  DFF_X1 \mem_reg[165][2]  ( .D(n24784), .CK(clk), .Q(\mem[165][2] ) );
  DFF_X1 \mem_reg[165][1]  ( .D(n24785), .CK(clk), .Q(\mem[165][1] ) );
  DFF_X1 \mem_reg[165][0]  ( .D(n24786), .CK(clk), .Q(\mem[165][0] ) );
  DFF_X1 \mem_reg[164][7]  ( .D(n24787), .CK(clk), .Q(\mem[164][7] ) );
  DFF_X1 \mem_reg[164][6]  ( .D(n24788), .CK(clk), .Q(\mem[164][6] ) );
  DFF_X1 \mem_reg[164][5]  ( .D(n24789), .CK(clk), .Q(\mem[164][5] ) );
  DFF_X1 \mem_reg[164][4]  ( .D(n24790), .CK(clk), .Q(\mem[164][4] ) );
  DFF_X1 \mem_reg[164][3]  ( .D(n24791), .CK(clk), .Q(\mem[164][3] ) );
  DFF_X1 \mem_reg[164][2]  ( .D(n24792), .CK(clk), .Q(\mem[164][2] ) );
  DFF_X1 \mem_reg[164][1]  ( .D(n24793), .CK(clk), .Q(\mem[164][1] ) );
  DFF_X1 \mem_reg[164][0]  ( .D(n24794), .CK(clk), .Q(\mem[164][0] ) );
  DFF_X1 \mem_reg[163][7]  ( .D(n24795), .CK(clk), .Q(\mem[163][7] ) );
  DFF_X1 \mem_reg[163][6]  ( .D(n24796), .CK(clk), .Q(\mem[163][6] ) );
  DFF_X1 \mem_reg[163][5]  ( .D(n24797), .CK(clk), .Q(\mem[163][5] ) );
  DFF_X1 \mem_reg[163][4]  ( .D(n24798), .CK(clk), .Q(\mem[163][4] ) );
  DFF_X1 \mem_reg[163][3]  ( .D(n24799), .CK(clk), .Q(\mem[163][3] ) );
  DFF_X1 \mem_reg[163][2]  ( .D(n24800), .CK(clk), .Q(\mem[163][2] ) );
  DFF_X1 \mem_reg[163][1]  ( .D(n24801), .CK(clk), .Q(\mem[163][1] ) );
  DFF_X1 \mem_reg[163][0]  ( .D(n24802), .CK(clk), .Q(\mem[163][0] ) );
  DFF_X1 \mem_reg[162][7]  ( .D(n24803), .CK(clk), .Q(\mem[162][7] ) );
  DFF_X1 \mem_reg[162][6]  ( .D(n24804), .CK(clk), .Q(\mem[162][6] ) );
  DFF_X1 \mem_reg[162][5]  ( .D(n24805), .CK(clk), .Q(\mem[162][5] ) );
  DFF_X1 \mem_reg[162][4]  ( .D(n24806), .CK(clk), .Q(\mem[162][4] ) );
  DFF_X1 \mem_reg[162][3]  ( .D(n24807), .CK(clk), .Q(\mem[162][3] ) );
  DFF_X1 \mem_reg[162][2]  ( .D(n24808), .CK(clk), .Q(\mem[162][2] ) );
  DFF_X1 \mem_reg[162][1]  ( .D(n24809), .CK(clk), .Q(\mem[162][1] ) );
  DFF_X1 \mem_reg[162][0]  ( .D(n24810), .CK(clk), .Q(\mem[162][0] ) );
  DFF_X1 \mem_reg[161][7]  ( .D(n24811), .CK(clk), .Q(\mem[161][7] ) );
  DFF_X1 \mem_reg[161][6]  ( .D(n24812), .CK(clk), .Q(\mem[161][6] ) );
  DFF_X1 \mem_reg[161][5]  ( .D(n24813), .CK(clk), .Q(\mem[161][5] ) );
  DFF_X1 \mem_reg[161][4]  ( .D(n24814), .CK(clk), .Q(\mem[161][4] ) );
  DFF_X1 \mem_reg[161][3]  ( .D(n24815), .CK(clk), .Q(\mem[161][3] ) );
  DFF_X1 \mem_reg[161][2]  ( .D(n24816), .CK(clk), .Q(\mem[161][2] ) );
  DFF_X1 \mem_reg[161][1]  ( .D(n24817), .CK(clk), .Q(\mem[161][1] ) );
  DFF_X1 \mem_reg[161][0]  ( .D(n24818), .CK(clk), .Q(\mem[161][0] ) );
  DFF_X1 \mem_reg[160][7]  ( .D(n24819), .CK(clk), .Q(\mem[160][7] ) );
  DFF_X1 \mem_reg[160][6]  ( .D(n24820), .CK(clk), .Q(\mem[160][6] ) );
  DFF_X1 \mem_reg[160][5]  ( .D(n24821), .CK(clk), .Q(\mem[160][5] ) );
  DFF_X1 \mem_reg[160][4]  ( .D(n24822), .CK(clk), .Q(\mem[160][4] ) );
  DFF_X1 \mem_reg[160][3]  ( .D(n24823), .CK(clk), .Q(\mem[160][3] ) );
  DFF_X1 \mem_reg[160][2]  ( .D(n24824), .CK(clk), .Q(\mem[160][2] ) );
  DFF_X1 \mem_reg[160][1]  ( .D(n24825), .CK(clk), .Q(\mem[160][1] ) );
  DFF_X1 \mem_reg[160][0]  ( .D(n24826), .CK(clk), .Q(\mem[160][0] ) );
  DFF_X1 \mem_reg[159][7]  ( .D(n24827), .CK(clk), .Q(\mem[159][7] ) );
  DFF_X1 \mem_reg[159][6]  ( .D(n24828), .CK(clk), .Q(\mem[159][6] ) );
  DFF_X1 \mem_reg[159][5]  ( .D(n24829), .CK(clk), .Q(\mem[159][5] ) );
  DFF_X1 \mem_reg[159][4]  ( .D(n24830), .CK(clk), .Q(\mem[159][4] ) );
  DFF_X1 \mem_reg[159][3]  ( .D(n24831), .CK(clk), .Q(\mem[159][3] ) );
  DFF_X1 \mem_reg[159][2]  ( .D(n24832), .CK(clk), .Q(\mem[159][2] ) );
  DFF_X1 \mem_reg[159][1]  ( .D(n24833), .CK(clk), .Q(\mem[159][1] ) );
  DFF_X1 \mem_reg[159][0]  ( .D(n24834), .CK(clk), .Q(\mem[159][0] ) );
  DFF_X1 \mem_reg[158][7]  ( .D(n24835), .CK(clk), .Q(\mem[158][7] ) );
  DFF_X1 \mem_reg[158][6]  ( .D(n24836), .CK(clk), .Q(\mem[158][6] ) );
  DFF_X1 \mem_reg[158][5]  ( .D(n24837), .CK(clk), .Q(\mem[158][5] ) );
  DFF_X1 \mem_reg[158][4]  ( .D(n24838), .CK(clk), .Q(\mem[158][4] ) );
  DFF_X1 \mem_reg[158][3]  ( .D(n24839), .CK(clk), .Q(\mem[158][3] ) );
  DFF_X1 \mem_reg[158][2]  ( .D(n24840), .CK(clk), .Q(\mem[158][2] ) );
  DFF_X1 \mem_reg[158][1]  ( .D(n24841), .CK(clk), .Q(\mem[158][1] ) );
  DFF_X1 \mem_reg[158][0]  ( .D(n24842), .CK(clk), .Q(\mem[158][0] ) );
  DFF_X1 \mem_reg[157][7]  ( .D(n24843), .CK(clk), .Q(\mem[157][7] ) );
  DFF_X1 \mem_reg[157][6]  ( .D(n24844), .CK(clk), .Q(\mem[157][6] ) );
  DFF_X1 \mem_reg[157][5]  ( .D(n24845), .CK(clk), .Q(\mem[157][5] ) );
  DFF_X1 \mem_reg[157][4]  ( .D(n24846), .CK(clk), .Q(\mem[157][4] ) );
  DFF_X1 \mem_reg[157][3]  ( .D(n24847), .CK(clk), .Q(\mem[157][3] ) );
  DFF_X1 \mem_reg[157][2]  ( .D(n24848), .CK(clk), .Q(\mem[157][2] ) );
  DFF_X1 \mem_reg[157][1]  ( .D(n24849), .CK(clk), .Q(\mem[157][1] ) );
  DFF_X1 \mem_reg[157][0]  ( .D(n24850), .CK(clk), .Q(\mem[157][0] ) );
  DFF_X1 \mem_reg[156][7]  ( .D(n24851), .CK(clk), .Q(\mem[156][7] ) );
  DFF_X1 \mem_reg[156][6]  ( .D(n24852), .CK(clk), .Q(\mem[156][6] ) );
  DFF_X1 \mem_reg[156][5]  ( .D(n24853), .CK(clk), .Q(\mem[156][5] ) );
  DFF_X1 \mem_reg[156][4]  ( .D(n24854), .CK(clk), .Q(\mem[156][4] ) );
  DFF_X1 \mem_reg[156][3]  ( .D(n24855), .CK(clk), .Q(\mem[156][3] ) );
  DFF_X1 \mem_reg[156][2]  ( .D(n24856), .CK(clk), .Q(\mem[156][2] ) );
  DFF_X1 \mem_reg[156][1]  ( .D(n24857), .CK(clk), .Q(\mem[156][1] ) );
  DFF_X1 \mem_reg[156][0]  ( .D(n24858), .CK(clk), .Q(\mem[156][0] ) );
  DFF_X1 \mem_reg[155][7]  ( .D(n24859), .CK(clk), .Q(\mem[155][7] ) );
  DFF_X1 \mem_reg[155][6]  ( .D(n24860), .CK(clk), .Q(\mem[155][6] ) );
  DFF_X1 \mem_reg[155][5]  ( .D(n24861), .CK(clk), .Q(\mem[155][5] ) );
  DFF_X1 \mem_reg[155][4]  ( .D(n24862), .CK(clk), .Q(\mem[155][4] ) );
  DFF_X1 \mem_reg[155][3]  ( .D(n24863), .CK(clk), .Q(\mem[155][3] ) );
  DFF_X1 \mem_reg[155][2]  ( .D(n24864), .CK(clk), .Q(\mem[155][2] ) );
  DFF_X1 \mem_reg[155][1]  ( .D(n24865), .CK(clk), .Q(\mem[155][1] ) );
  DFF_X1 \mem_reg[155][0]  ( .D(n24866), .CK(clk), .Q(\mem[155][0] ) );
  DFF_X1 \mem_reg[154][7]  ( .D(n24867), .CK(clk), .Q(\mem[154][7] ) );
  DFF_X1 \mem_reg[154][6]  ( .D(n24868), .CK(clk), .Q(\mem[154][6] ) );
  DFF_X1 \mem_reg[154][5]  ( .D(n24869), .CK(clk), .Q(\mem[154][5] ) );
  DFF_X1 \mem_reg[154][4]  ( .D(n24870), .CK(clk), .Q(\mem[154][4] ) );
  DFF_X1 \mem_reg[154][3]  ( .D(n24871), .CK(clk), .Q(\mem[154][3] ) );
  DFF_X1 \mem_reg[154][2]  ( .D(n24872), .CK(clk), .Q(\mem[154][2] ) );
  DFF_X1 \mem_reg[154][1]  ( .D(n24873), .CK(clk), .Q(\mem[154][1] ) );
  DFF_X1 \mem_reg[154][0]  ( .D(n24874), .CK(clk), .Q(\mem[154][0] ) );
  DFF_X1 \mem_reg[153][7]  ( .D(n24875), .CK(clk), .Q(\mem[153][7] ) );
  DFF_X1 \mem_reg[153][6]  ( .D(n24876), .CK(clk), .Q(\mem[153][6] ) );
  DFF_X1 \mem_reg[153][5]  ( .D(n24877), .CK(clk), .Q(\mem[153][5] ) );
  DFF_X1 \mem_reg[153][4]  ( .D(n24878), .CK(clk), .Q(\mem[153][4] ) );
  DFF_X1 \mem_reg[153][3]  ( .D(n24879), .CK(clk), .Q(\mem[153][3] ) );
  DFF_X1 \mem_reg[153][2]  ( .D(n24880), .CK(clk), .Q(\mem[153][2] ) );
  DFF_X1 \mem_reg[153][1]  ( .D(n24881), .CK(clk), .Q(\mem[153][1] ) );
  DFF_X1 \mem_reg[153][0]  ( .D(n24882), .CK(clk), .Q(\mem[153][0] ) );
  DFF_X1 \mem_reg[152][7]  ( .D(n24883), .CK(clk), .Q(\mem[152][7] ) );
  DFF_X1 \mem_reg[152][6]  ( .D(n24884), .CK(clk), .Q(\mem[152][6] ) );
  DFF_X1 \mem_reg[152][5]  ( .D(n24885), .CK(clk), .Q(\mem[152][5] ) );
  DFF_X1 \mem_reg[152][4]  ( .D(n24886), .CK(clk), .Q(\mem[152][4] ) );
  DFF_X1 \mem_reg[152][3]  ( .D(n24887), .CK(clk), .Q(\mem[152][3] ) );
  DFF_X1 \mem_reg[152][2]  ( .D(n24888), .CK(clk), .Q(\mem[152][2] ) );
  DFF_X1 \mem_reg[152][1]  ( .D(n24889), .CK(clk), .Q(\mem[152][1] ) );
  DFF_X1 \mem_reg[152][0]  ( .D(n24890), .CK(clk), .Q(\mem[152][0] ) );
  DFF_X1 \mem_reg[151][7]  ( .D(n24891), .CK(clk), .Q(\mem[151][7] ) );
  DFF_X1 \mem_reg[151][6]  ( .D(n24892), .CK(clk), .Q(\mem[151][6] ) );
  DFF_X1 \mem_reg[151][5]  ( .D(n24893), .CK(clk), .Q(\mem[151][5] ) );
  DFF_X1 \mem_reg[151][4]  ( .D(n24894), .CK(clk), .Q(\mem[151][4] ) );
  DFF_X1 \mem_reg[151][3]  ( .D(n24895), .CK(clk), .Q(\mem[151][3] ) );
  DFF_X1 \mem_reg[151][2]  ( .D(n24896), .CK(clk), .Q(\mem[151][2] ) );
  DFF_X1 \mem_reg[151][1]  ( .D(n24897), .CK(clk), .Q(\mem[151][1] ) );
  DFF_X1 \mem_reg[151][0]  ( .D(n24898), .CK(clk), .Q(\mem[151][0] ) );
  DFF_X1 \mem_reg[150][7]  ( .D(n24899), .CK(clk), .Q(\mem[150][7] ) );
  DFF_X1 \mem_reg[150][6]  ( .D(n24900), .CK(clk), .Q(\mem[150][6] ) );
  DFF_X1 \mem_reg[150][5]  ( .D(n24901), .CK(clk), .Q(\mem[150][5] ) );
  DFF_X1 \mem_reg[150][4]  ( .D(n24902), .CK(clk), .Q(\mem[150][4] ) );
  DFF_X1 \mem_reg[150][3]  ( .D(n24903), .CK(clk), .Q(\mem[150][3] ) );
  DFF_X1 \mem_reg[150][2]  ( .D(n24904), .CK(clk), .Q(\mem[150][2] ) );
  DFF_X1 \mem_reg[150][1]  ( .D(n24905), .CK(clk), .Q(\mem[150][1] ) );
  DFF_X1 \mem_reg[150][0]  ( .D(n24906), .CK(clk), .Q(\mem[150][0] ) );
  DFF_X1 \mem_reg[149][7]  ( .D(n24907), .CK(clk), .Q(\mem[149][7] ) );
  DFF_X1 \mem_reg[149][6]  ( .D(n24908), .CK(clk), .Q(\mem[149][6] ) );
  DFF_X1 \mem_reg[149][5]  ( .D(n24909), .CK(clk), .Q(\mem[149][5] ) );
  DFF_X1 \mem_reg[149][4]  ( .D(n24910), .CK(clk), .Q(\mem[149][4] ) );
  DFF_X1 \mem_reg[149][3]  ( .D(n24911), .CK(clk), .Q(\mem[149][3] ) );
  DFF_X1 \mem_reg[149][2]  ( .D(n24912), .CK(clk), .Q(\mem[149][2] ) );
  DFF_X1 \mem_reg[149][1]  ( .D(n24913), .CK(clk), .Q(\mem[149][1] ) );
  DFF_X1 \mem_reg[149][0]  ( .D(n24914), .CK(clk), .Q(\mem[149][0] ) );
  DFF_X1 \mem_reg[148][7]  ( .D(n24915), .CK(clk), .Q(\mem[148][7] ) );
  DFF_X1 \mem_reg[148][6]  ( .D(n24916), .CK(clk), .Q(\mem[148][6] ) );
  DFF_X1 \mem_reg[148][5]  ( .D(n24917), .CK(clk), .Q(\mem[148][5] ) );
  DFF_X1 \mem_reg[148][4]  ( .D(n24918), .CK(clk), .Q(\mem[148][4] ) );
  DFF_X1 \mem_reg[148][3]  ( .D(n24919), .CK(clk), .Q(\mem[148][3] ) );
  DFF_X1 \mem_reg[148][2]  ( .D(n24920), .CK(clk), .Q(\mem[148][2] ) );
  DFF_X1 \mem_reg[148][1]  ( .D(n24921), .CK(clk), .Q(\mem[148][1] ) );
  DFF_X1 \mem_reg[148][0]  ( .D(n24922), .CK(clk), .Q(\mem[148][0] ) );
  DFF_X1 \mem_reg[147][7]  ( .D(n24923), .CK(clk), .Q(\mem[147][7] ) );
  DFF_X1 \mem_reg[147][6]  ( .D(n24924), .CK(clk), .Q(\mem[147][6] ) );
  DFF_X1 \mem_reg[147][5]  ( .D(n24925), .CK(clk), .Q(\mem[147][5] ) );
  DFF_X1 \mem_reg[147][4]  ( .D(n24926), .CK(clk), .Q(\mem[147][4] ) );
  DFF_X1 \mem_reg[147][3]  ( .D(n24927), .CK(clk), .Q(\mem[147][3] ) );
  DFF_X1 \mem_reg[147][2]  ( .D(n24928), .CK(clk), .Q(\mem[147][2] ) );
  DFF_X1 \mem_reg[147][1]  ( .D(n24929), .CK(clk), .Q(\mem[147][1] ) );
  DFF_X1 \mem_reg[147][0]  ( .D(n24930), .CK(clk), .Q(\mem[147][0] ) );
  DFF_X1 \mem_reg[146][7]  ( .D(n24931), .CK(clk), .Q(\mem[146][7] ) );
  DFF_X1 \mem_reg[146][6]  ( .D(n24932), .CK(clk), .Q(\mem[146][6] ) );
  DFF_X1 \mem_reg[146][5]  ( .D(n24933), .CK(clk), .Q(\mem[146][5] ) );
  DFF_X1 \mem_reg[146][4]  ( .D(n24934), .CK(clk), .Q(\mem[146][4] ) );
  DFF_X1 \mem_reg[146][3]  ( .D(n24935), .CK(clk), .Q(\mem[146][3] ) );
  DFF_X1 \mem_reg[146][2]  ( .D(n24936), .CK(clk), .Q(\mem[146][2] ) );
  DFF_X1 \mem_reg[146][1]  ( .D(n24937), .CK(clk), .Q(\mem[146][1] ) );
  DFF_X1 \mem_reg[146][0]  ( .D(n24938), .CK(clk), .Q(\mem[146][0] ) );
  DFF_X1 \mem_reg[145][7]  ( .D(n24939), .CK(clk), .Q(\mem[145][7] ) );
  DFF_X1 \mem_reg[145][6]  ( .D(n24940), .CK(clk), .Q(\mem[145][6] ) );
  DFF_X1 \mem_reg[145][5]  ( .D(n24941), .CK(clk), .Q(\mem[145][5] ) );
  DFF_X1 \mem_reg[145][4]  ( .D(n24942), .CK(clk), .Q(\mem[145][4] ) );
  DFF_X1 \mem_reg[145][3]  ( .D(n24943), .CK(clk), .Q(\mem[145][3] ) );
  DFF_X1 \mem_reg[145][2]  ( .D(n24944), .CK(clk), .Q(\mem[145][2] ) );
  DFF_X1 \mem_reg[145][1]  ( .D(n24945), .CK(clk), .Q(\mem[145][1] ) );
  DFF_X1 \mem_reg[145][0]  ( .D(n24946), .CK(clk), .Q(\mem[145][0] ) );
  DFF_X1 \mem_reg[144][7]  ( .D(n24947), .CK(clk), .Q(\mem[144][7] ) );
  DFF_X1 \mem_reg[144][6]  ( .D(n24948), .CK(clk), .Q(\mem[144][6] ) );
  DFF_X1 \mem_reg[144][5]  ( .D(n24949), .CK(clk), .Q(\mem[144][5] ) );
  DFF_X1 \mem_reg[144][4]  ( .D(n24950), .CK(clk), .Q(\mem[144][4] ) );
  DFF_X1 \mem_reg[144][3]  ( .D(n24951), .CK(clk), .Q(\mem[144][3] ) );
  DFF_X1 \mem_reg[144][2]  ( .D(n24952), .CK(clk), .Q(\mem[144][2] ) );
  DFF_X1 \mem_reg[144][1]  ( .D(n24953), .CK(clk), .Q(\mem[144][1] ) );
  DFF_X1 \mem_reg[144][0]  ( .D(n24954), .CK(clk), .Q(\mem[144][0] ) );
  DFF_X1 \mem_reg[143][7]  ( .D(n24955), .CK(clk), .Q(\mem[143][7] ) );
  DFF_X1 \mem_reg[143][6]  ( .D(n24956), .CK(clk), .Q(\mem[143][6] ) );
  DFF_X1 \mem_reg[143][5]  ( .D(n24957), .CK(clk), .Q(\mem[143][5] ) );
  DFF_X1 \mem_reg[143][4]  ( .D(n24958), .CK(clk), .Q(\mem[143][4] ) );
  DFF_X1 \mem_reg[143][3]  ( .D(n24959), .CK(clk), .Q(\mem[143][3] ) );
  DFF_X1 \mem_reg[143][2]  ( .D(n24960), .CK(clk), .Q(\mem[143][2] ) );
  DFF_X1 \mem_reg[143][1]  ( .D(n24961), .CK(clk), .Q(\mem[143][1] ) );
  DFF_X1 \mem_reg[143][0]  ( .D(n24962), .CK(clk), .Q(\mem[143][0] ) );
  DFF_X1 \mem_reg[142][7]  ( .D(n24963), .CK(clk), .Q(\mem[142][7] ) );
  DFF_X1 \mem_reg[142][6]  ( .D(n24964), .CK(clk), .Q(\mem[142][6] ) );
  DFF_X1 \mem_reg[142][5]  ( .D(n24965), .CK(clk), .Q(\mem[142][5] ) );
  DFF_X1 \mem_reg[142][4]  ( .D(n24966), .CK(clk), .Q(\mem[142][4] ) );
  DFF_X1 \mem_reg[142][3]  ( .D(n24967), .CK(clk), .Q(\mem[142][3] ) );
  DFF_X1 \mem_reg[142][2]  ( .D(n24968), .CK(clk), .Q(\mem[142][2] ) );
  DFF_X1 \mem_reg[142][1]  ( .D(n24969), .CK(clk), .Q(\mem[142][1] ) );
  DFF_X1 \mem_reg[142][0]  ( .D(n24970), .CK(clk), .Q(\mem[142][0] ) );
  DFF_X1 \mem_reg[141][7]  ( .D(n24971), .CK(clk), .Q(\mem[141][7] ) );
  DFF_X1 \mem_reg[141][6]  ( .D(n24972), .CK(clk), .Q(\mem[141][6] ) );
  DFF_X1 \mem_reg[141][5]  ( .D(n24973), .CK(clk), .Q(\mem[141][5] ) );
  DFF_X1 \mem_reg[141][4]  ( .D(n24974), .CK(clk), .Q(\mem[141][4] ) );
  DFF_X1 \mem_reg[141][3]  ( .D(n24975), .CK(clk), .Q(\mem[141][3] ) );
  DFF_X1 \mem_reg[141][2]  ( .D(n24976), .CK(clk), .Q(\mem[141][2] ) );
  DFF_X1 \mem_reg[141][1]  ( .D(n24977), .CK(clk), .Q(\mem[141][1] ) );
  DFF_X1 \mem_reg[141][0]  ( .D(n24978), .CK(clk), .Q(\mem[141][0] ) );
  DFF_X1 \mem_reg[140][7]  ( .D(n24979), .CK(clk), .Q(\mem[140][7] ) );
  DFF_X1 \mem_reg[140][6]  ( .D(n24980), .CK(clk), .Q(\mem[140][6] ) );
  DFF_X1 \mem_reg[140][5]  ( .D(n24981), .CK(clk), .Q(\mem[140][5] ) );
  DFF_X1 \mem_reg[140][4]  ( .D(n24982), .CK(clk), .Q(\mem[140][4] ) );
  DFF_X1 \mem_reg[140][3]  ( .D(n24983), .CK(clk), .Q(\mem[140][3] ) );
  DFF_X1 \mem_reg[140][2]  ( .D(n24984), .CK(clk), .Q(\mem[140][2] ) );
  DFF_X1 \mem_reg[140][1]  ( .D(n24985), .CK(clk), .Q(\mem[140][1] ) );
  DFF_X1 \mem_reg[140][0]  ( .D(n24986), .CK(clk), .Q(\mem[140][0] ) );
  DFF_X1 \mem_reg[139][7]  ( .D(n24987), .CK(clk), .Q(\mem[139][7] ) );
  DFF_X1 \mem_reg[139][6]  ( .D(n24988), .CK(clk), .Q(\mem[139][6] ) );
  DFF_X1 \mem_reg[139][5]  ( .D(n24989), .CK(clk), .Q(\mem[139][5] ) );
  DFF_X1 \mem_reg[139][4]  ( .D(n24990), .CK(clk), .Q(\mem[139][4] ) );
  DFF_X1 \mem_reg[139][3]  ( .D(n24991), .CK(clk), .Q(\mem[139][3] ) );
  DFF_X1 \mem_reg[139][2]  ( .D(n24992), .CK(clk), .Q(\mem[139][2] ) );
  DFF_X1 \mem_reg[139][1]  ( .D(n24993), .CK(clk), .Q(\mem[139][1] ) );
  DFF_X1 \mem_reg[139][0]  ( .D(n24994), .CK(clk), .Q(\mem[139][0] ) );
  DFF_X1 \mem_reg[138][7]  ( .D(n24995), .CK(clk), .Q(\mem[138][7] ) );
  DFF_X1 \mem_reg[138][6]  ( .D(n24996), .CK(clk), .Q(\mem[138][6] ) );
  DFF_X1 \mem_reg[138][5]  ( .D(n24997), .CK(clk), .Q(\mem[138][5] ) );
  DFF_X1 \mem_reg[138][4]  ( .D(n24998), .CK(clk), .Q(\mem[138][4] ) );
  DFF_X1 \mem_reg[138][3]  ( .D(n24999), .CK(clk), .Q(\mem[138][3] ) );
  DFF_X1 \mem_reg[138][2]  ( .D(n25000), .CK(clk), .Q(\mem[138][2] ) );
  DFF_X1 \mem_reg[138][1]  ( .D(n25001), .CK(clk), .Q(\mem[138][1] ) );
  DFF_X1 \mem_reg[138][0]  ( .D(n25002), .CK(clk), .Q(\mem[138][0] ) );
  DFF_X1 \mem_reg[137][7]  ( .D(n25003), .CK(clk), .Q(\mem[137][7] ) );
  DFF_X1 \mem_reg[137][6]  ( .D(n25004), .CK(clk), .Q(\mem[137][6] ) );
  DFF_X1 \mem_reg[137][5]  ( .D(n25005), .CK(clk), .Q(\mem[137][5] ) );
  DFF_X1 \mem_reg[137][4]  ( .D(n25006), .CK(clk), .Q(\mem[137][4] ) );
  DFF_X1 \mem_reg[137][3]  ( .D(n25007), .CK(clk), .Q(\mem[137][3] ) );
  DFF_X1 \mem_reg[137][2]  ( .D(n25008), .CK(clk), .Q(\mem[137][2] ) );
  DFF_X1 \mem_reg[137][1]  ( .D(n25009), .CK(clk), .Q(\mem[137][1] ) );
  DFF_X1 \mem_reg[137][0]  ( .D(n25010), .CK(clk), .Q(\mem[137][0] ) );
  DFF_X1 \mem_reg[136][7]  ( .D(n25011), .CK(clk), .Q(\mem[136][7] ) );
  DFF_X1 \mem_reg[136][6]  ( .D(n25012), .CK(clk), .Q(\mem[136][6] ) );
  DFF_X1 \mem_reg[136][5]  ( .D(n25013), .CK(clk), .Q(\mem[136][5] ) );
  DFF_X1 \mem_reg[136][4]  ( .D(n25014), .CK(clk), .Q(\mem[136][4] ) );
  DFF_X1 \mem_reg[136][3]  ( .D(n25015), .CK(clk), .Q(\mem[136][3] ) );
  DFF_X1 \mem_reg[136][2]  ( .D(n25016), .CK(clk), .Q(\mem[136][2] ) );
  DFF_X1 \mem_reg[136][1]  ( .D(n25017), .CK(clk), .Q(\mem[136][1] ) );
  DFF_X1 \mem_reg[136][0]  ( .D(n25018), .CK(clk), .Q(\mem[136][0] ) );
  DFF_X1 \mem_reg[135][7]  ( .D(n25019), .CK(clk), .Q(\mem[135][7] ) );
  DFF_X1 \mem_reg[135][6]  ( .D(n25020), .CK(clk), .Q(\mem[135][6] ) );
  DFF_X1 \mem_reg[135][5]  ( .D(n25021), .CK(clk), .Q(\mem[135][5] ) );
  DFF_X1 \mem_reg[135][4]  ( .D(n25022), .CK(clk), .Q(\mem[135][4] ) );
  DFF_X1 \mem_reg[135][3]  ( .D(n25023), .CK(clk), .Q(\mem[135][3] ) );
  DFF_X1 \mem_reg[135][2]  ( .D(n25024), .CK(clk), .Q(\mem[135][2] ) );
  DFF_X1 \mem_reg[135][1]  ( .D(n25025), .CK(clk), .Q(\mem[135][1] ) );
  DFF_X1 \mem_reg[135][0]  ( .D(n25026), .CK(clk), .Q(\mem[135][0] ) );
  DFF_X1 \mem_reg[134][7]  ( .D(n25027), .CK(clk), .Q(\mem[134][7] ) );
  DFF_X1 \mem_reg[134][6]  ( .D(n25028), .CK(clk), .Q(\mem[134][6] ) );
  DFF_X1 \mem_reg[134][5]  ( .D(n25029), .CK(clk), .Q(\mem[134][5] ) );
  DFF_X1 \mem_reg[134][4]  ( .D(n25030), .CK(clk), .Q(\mem[134][4] ) );
  DFF_X1 \mem_reg[134][3]  ( .D(n25031), .CK(clk), .Q(\mem[134][3] ) );
  DFF_X1 \mem_reg[134][2]  ( .D(n25032), .CK(clk), .Q(\mem[134][2] ) );
  DFF_X1 \mem_reg[134][1]  ( .D(n25033), .CK(clk), .Q(\mem[134][1] ) );
  DFF_X1 \mem_reg[134][0]  ( .D(n25034), .CK(clk), .Q(\mem[134][0] ) );
  DFF_X1 \mem_reg[133][7]  ( .D(n25035), .CK(clk), .Q(\mem[133][7] ) );
  DFF_X1 \mem_reg[133][6]  ( .D(n25036), .CK(clk), .Q(\mem[133][6] ) );
  DFF_X1 \mem_reg[133][5]  ( .D(n25037), .CK(clk), .Q(\mem[133][5] ) );
  DFF_X1 \mem_reg[133][4]  ( .D(n25038), .CK(clk), .Q(\mem[133][4] ) );
  DFF_X1 \mem_reg[133][3]  ( .D(n25039), .CK(clk), .Q(\mem[133][3] ) );
  DFF_X1 \mem_reg[133][2]  ( .D(n25040), .CK(clk), .Q(\mem[133][2] ) );
  DFF_X1 \mem_reg[133][1]  ( .D(n25041), .CK(clk), .Q(\mem[133][1] ) );
  DFF_X1 \mem_reg[133][0]  ( .D(n25042), .CK(clk), .Q(\mem[133][0] ) );
  DFF_X1 \mem_reg[132][7]  ( .D(n25043), .CK(clk), .Q(\mem[132][7] ) );
  DFF_X1 \mem_reg[132][6]  ( .D(n25044), .CK(clk), .Q(\mem[132][6] ) );
  DFF_X1 \mem_reg[132][5]  ( .D(n25045), .CK(clk), .Q(\mem[132][5] ) );
  DFF_X1 \mem_reg[132][4]  ( .D(n25046), .CK(clk), .Q(\mem[132][4] ) );
  DFF_X1 \mem_reg[132][3]  ( .D(n25047), .CK(clk), .Q(\mem[132][3] ) );
  DFF_X1 \mem_reg[132][2]  ( .D(n25048), .CK(clk), .Q(\mem[132][2] ) );
  DFF_X1 \mem_reg[132][1]  ( .D(n25049), .CK(clk), .Q(\mem[132][1] ) );
  DFF_X1 \mem_reg[132][0]  ( .D(n25050), .CK(clk), .Q(\mem[132][0] ) );
  DFF_X1 \mem_reg[131][7]  ( .D(n25051), .CK(clk), .Q(\mem[131][7] ) );
  DFF_X1 \mem_reg[131][6]  ( .D(n25052), .CK(clk), .Q(\mem[131][6] ) );
  DFF_X1 \mem_reg[131][5]  ( .D(n25053), .CK(clk), .Q(\mem[131][5] ) );
  DFF_X1 \mem_reg[131][4]  ( .D(n25054), .CK(clk), .Q(\mem[131][4] ) );
  DFF_X1 \mem_reg[131][3]  ( .D(n25055), .CK(clk), .Q(\mem[131][3] ) );
  DFF_X1 \mem_reg[131][2]  ( .D(n25056), .CK(clk), .Q(\mem[131][2] ) );
  DFF_X1 \mem_reg[131][1]  ( .D(n25057), .CK(clk), .Q(\mem[131][1] ) );
  DFF_X1 \mem_reg[131][0]  ( .D(n25058), .CK(clk), .Q(\mem[131][0] ) );
  DFF_X1 \mem_reg[130][7]  ( .D(n25059), .CK(clk), .Q(\mem[130][7] ) );
  DFF_X1 \mem_reg[130][6]  ( .D(n25060), .CK(clk), .Q(\mem[130][6] ) );
  DFF_X1 \mem_reg[130][5]  ( .D(n25061), .CK(clk), .Q(\mem[130][5] ) );
  DFF_X1 \mem_reg[130][4]  ( .D(n25062), .CK(clk), .Q(\mem[130][4] ) );
  DFF_X1 \mem_reg[130][3]  ( .D(n25063), .CK(clk), .Q(\mem[130][3] ) );
  DFF_X1 \mem_reg[130][2]  ( .D(n25064), .CK(clk), .Q(\mem[130][2] ) );
  DFF_X1 \mem_reg[130][1]  ( .D(n25065), .CK(clk), .Q(\mem[130][1] ) );
  DFF_X1 \mem_reg[130][0]  ( .D(n25066), .CK(clk), .Q(\mem[130][0] ) );
  DFF_X1 \mem_reg[129][7]  ( .D(n25067), .CK(clk), .Q(\mem[129][7] ) );
  DFF_X1 \mem_reg[129][6]  ( .D(n25068), .CK(clk), .Q(\mem[129][6] ) );
  DFF_X1 \mem_reg[129][5]  ( .D(n25069), .CK(clk), .Q(\mem[129][5] ) );
  DFF_X1 \mem_reg[129][4]  ( .D(n25070), .CK(clk), .Q(\mem[129][4] ) );
  DFF_X1 \mem_reg[129][3]  ( .D(n25071), .CK(clk), .Q(\mem[129][3] ) );
  DFF_X1 \mem_reg[129][2]  ( .D(n25072), .CK(clk), .Q(\mem[129][2] ) );
  DFF_X1 \mem_reg[129][1]  ( .D(n25073), .CK(clk), .Q(\mem[129][1] ) );
  DFF_X1 \mem_reg[129][0]  ( .D(n25074), .CK(clk), .Q(\mem[129][0] ) );
  DFF_X1 \mem_reg[128][7]  ( .D(n25075), .CK(clk), .Q(\mem[128][7] ) );
  DFF_X1 \mem_reg[128][6]  ( .D(n25076), .CK(clk), .Q(\mem[128][6] ) );
  DFF_X1 \mem_reg[128][5]  ( .D(n25077), .CK(clk), .Q(\mem[128][5] ) );
  DFF_X1 \mem_reg[128][4]  ( .D(n25078), .CK(clk), .Q(\mem[128][4] ) );
  DFF_X1 \mem_reg[128][3]  ( .D(n25079), .CK(clk), .Q(\mem[128][3] ) );
  DFF_X1 \mem_reg[128][2]  ( .D(n25080), .CK(clk), .Q(\mem[128][2] ) );
  DFF_X1 \mem_reg[128][1]  ( .D(n25081), .CK(clk), .Q(\mem[128][1] ) );
  DFF_X1 \mem_reg[128][0]  ( .D(n25082), .CK(clk), .Q(\mem[128][0] ) );
  DFF_X1 \mem_reg[127][7]  ( .D(n25083), .CK(clk), .Q(\mem[127][7] ) );
  DFF_X1 \mem_reg[127][6]  ( .D(n25084), .CK(clk), .Q(\mem[127][6] ) );
  DFF_X1 \mem_reg[127][5]  ( .D(n25085), .CK(clk), .Q(\mem[127][5] ) );
  DFF_X1 \mem_reg[127][4]  ( .D(n25086), .CK(clk), .Q(\mem[127][4] ) );
  DFF_X1 \mem_reg[127][3]  ( .D(n25087), .CK(clk), .Q(\mem[127][3] ) );
  DFF_X1 \mem_reg[127][2]  ( .D(n25088), .CK(clk), .Q(\mem[127][2] ) );
  DFF_X1 \mem_reg[127][1]  ( .D(n25089), .CK(clk), .Q(\mem[127][1] ) );
  DFF_X1 \mem_reg[127][0]  ( .D(n25090), .CK(clk), .Q(\mem[127][0] ) );
  DFF_X1 \mem_reg[126][7]  ( .D(n25091), .CK(clk), .Q(\mem[126][7] ) );
  DFF_X1 \mem_reg[126][6]  ( .D(n25092), .CK(clk), .Q(\mem[126][6] ) );
  DFF_X1 \mem_reg[126][5]  ( .D(n25093), .CK(clk), .Q(\mem[126][5] ) );
  DFF_X1 \mem_reg[126][4]  ( .D(n25094), .CK(clk), .Q(\mem[126][4] ) );
  DFF_X1 \mem_reg[126][3]  ( .D(n25095), .CK(clk), .Q(\mem[126][3] ) );
  DFF_X1 \mem_reg[126][2]  ( .D(n25096), .CK(clk), .Q(\mem[126][2] ) );
  DFF_X1 \mem_reg[126][1]  ( .D(n25097), .CK(clk), .Q(\mem[126][1] ) );
  DFF_X1 \mem_reg[126][0]  ( .D(n25098), .CK(clk), .Q(\mem[126][0] ) );
  DFF_X1 \mem_reg[125][7]  ( .D(n25099), .CK(clk), .Q(\mem[125][7] ) );
  DFF_X1 \mem_reg[125][6]  ( .D(n25100), .CK(clk), .Q(\mem[125][6] ) );
  DFF_X1 \mem_reg[125][5]  ( .D(n25101), .CK(clk), .Q(\mem[125][5] ) );
  DFF_X1 \mem_reg[125][4]  ( .D(n25102), .CK(clk), .Q(\mem[125][4] ) );
  DFF_X1 \mem_reg[125][3]  ( .D(n25103), .CK(clk), .Q(\mem[125][3] ) );
  DFF_X1 \mem_reg[125][2]  ( .D(n25104), .CK(clk), .Q(\mem[125][2] ) );
  DFF_X1 \mem_reg[125][1]  ( .D(n25105), .CK(clk), .Q(\mem[125][1] ) );
  DFF_X1 \mem_reg[125][0]  ( .D(n25106), .CK(clk), .Q(\mem[125][0] ) );
  DFF_X1 \mem_reg[124][7]  ( .D(n25107), .CK(clk), .Q(\mem[124][7] ) );
  DFF_X1 \mem_reg[124][6]  ( .D(n25108), .CK(clk), .Q(\mem[124][6] ) );
  DFF_X1 \mem_reg[124][5]  ( .D(n25109), .CK(clk), .Q(\mem[124][5] ) );
  DFF_X1 \mem_reg[124][4]  ( .D(n25110), .CK(clk), .Q(\mem[124][4] ) );
  DFF_X1 \mem_reg[124][3]  ( .D(n25111), .CK(clk), .Q(\mem[124][3] ) );
  DFF_X1 \mem_reg[124][2]  ( .D(n25112), .CK(clk), .Q(\mem[124][2] ) );
  DFF_X1 \mem_reg[124][1]  ( .D(n25113), .CK(clk), .Q(\mem[124][1] ) );
  DFF_X1 \mem_reg[124][0]  ( .D(n25114), .CK(clk), .Q(\mem[124][0] ) );
  DFF_X1 \mem_reg[123][7]  ( .D(n25115), .CK(clk), .Q(\mem[123][7] ) );
  DFF_X1 \mem_reg[123][6]  ( .D(n25116), .CK(clk), .Q(\mem[123][6] ) );
  DFF_X1 \mem_reg[123][5]  ( .D(n25117), .CK(clk), .Q(\mem[123][5] ) );
  DFF_X1 \mem_reg[123][4]  ( .D(n25118), .CK(clk), .Q(\mem[123][4] ) );
  DFF_X1 \mem_reg[123][3]  ( .D(n25119), .CK(clk), .Q(\mem[123][3] ) );
  DFF_X1 \mem_reg[123][2]  ( .D(n25120), .CK(clk), .Q(\mem[123][2] ) );
  DFF_X1 \mem_reg[123][1]  ( .D(n25121), .CK(clk), .Q(\mem[123][1] ) );
  DFF_X1 \mem_reg[123][0]  ( .D(n25122), .CK(clk), .Q(\mem[123][0] ) );
  DFF_X1 \mem_reg[122][7]  ( .D(n25123), .CK(clk), .Q(\mem[122][7] ) );
  DFF_X1 \mem_reg[122][6]  ( .D(n25124), .CK(clk), .Q(\mem[122][6] ) );
  DFF_X1 \mem_reg[122][5]  ( .D(n25125), .CK(clk), .Q(\mem[122][5] ) );
  DFF_X1 \mem_reg[122][4]  ( .D(n25126), .CK(clk), .Q(\mem[122][4] ) );
  DFF_X1 \mem_reg[122][3]  ( .D(n25127), .CK(clk), .Q(\mem[122][3] ) );
  DFF_X1 \mem_reg[122][2]  ( .D(n25128), .CK(clk), .Q(\mem[122][2] ) );
  DFF_X1 \mem_reg[122][1]  ( .D(n25129), .CK(clk), .Q(\mem[122][1] ) );
  DFF_X1 \mem_reg[122][0]  ( .D(n25130), .CK(clk), .Q(\mem[122][0] ) );
  DFF_X1 \mem_reg[121][7]  ( .D(n25131), .CK(clk), .Q(\mem[121][7] ) );
  DFF_X1 \mem_reg[121][6]  ( .D(n25132), .CK(clk), .Q(\mem[121][6] ) );
  DFF_X1 \mem_reg[121][5]  ( .D(n25133), .CK(clk), .Q(\mem[121][5] ) );
  DFF_X1 \mem_reg[121][4]  ( .D(n25134), .CK(clk), .Q(\mem[121][4] ) );
  DFF_X1 \mem_reg[121][3]  ( .D(n25135), .CK(clk), .Q(\mem[121][3] ) );
  DFF_X1 \mem_reg[121][2]  ( .D(n25136), .CK(clk), .Q(\mem[121][2] ) );
  DFF_X1 \mem_reg[121][1]  ( .D(n25137), .CK(clk), .Q(\mem[121][1] ) );
  DFF_X1 \mem_reg[121][0]  ( .D(n25138), .CK(clk), .Q(\mem[121][0] ) );
  DFF_X1 \mem_reg[120][7]  ( .D(n25139), .CK(clk), .Q(\mem[120][7] ) );
  DFF_X1 \mem_reg[120][6]  ( .D(n25140), .CK(clk), .Q(\mem[120][6] ) );
  DFF_X1 \mem_reg[120][5]  ( .D(n25141), .CK(clk), .Q(\mem[120][5] ) );
  DFF_X1 \mem_reg[120][4]  ( .D(n25142), .CK(clk), .Q(\mem[120][4] ) );
  DFF_X1 \mem_reg[120][3]  ( .D(n25143), .CK(clk), .Q(\mem[120][3] ) );
  DFF_X1 \mem_reg[120][2]  ( .D(n25144), .CK(clk), .Q(\mem[120][2] ) );
  DFF_X1 \mem_reg[120][1]  ( .D(n25145), .CK(clk), .Q(\mem[120][1] ) );
  DFF_X1 \mem_reg[120][0]  ( .D(n25146), .CK(clk), .Q(\mem[120][0] ) );
  DFF_X1 \mem_reg[119][7]  ( .D(n25147), .CK(clk), .Q(\mem[119][7] ) );
  DFF_X1 \mem_reg[119][6]  ( .D(n25148), .CK(clk), .Q(\mem[119][6] ) );
  DFF_X1 \mem_reg[119][5]  ( .D(n25149), .CK(clk), .Q(\mem[119][5] ) );
  DFF_X1 \mem_reg[119][4]  ( .D(n25150), .CK(clk), .Q(\mem[119][4] ) );
  DFF_X1 \mem_reg[119][3]  ( .D(n25151), .CK(clk), .Q(\mem[119][3] ) );
  DFF_X1 \mem_reg[119][2]  ( .D(n25152), .CK(clk), .Q(\mem[119][2] ) );
  DFF_X1 \mem_reg[119][1]  ( .D(n25153), .CK(clk), .Q(\mem[119][1] ) );
  DFF_X1 \mem_reg[119][0]  ( .D(n25154), .CK(clk), .Q(\mem[119][0] ) );
  DFF_X1 \mem_reg[118][7]  ( .D(n25155), .CK(clk), .Q(\mem[118][7] ) );
  DFF_X1 \mem_reg[118][6]  ( .D(n25156), .CK(clk), .Q(\mem[118][6] ) );
  DFF_X1 \mem_reg[118][5]  ( .D(n25157), .CK(clk), .Q(\mem[118][5] ) );
  DFF_X1 \mem_reg[118][4]  ( .D(n25158), .CK(clk), .Q(\mem[118][4] ) );
  DFF_X1 \mem_reg[118][3]  ( .D(n25159), .CK(clk), .Q(\mem[118][3] ) );
  DFF_X1 \mem_reg[118][2]  ( .D(n25160), .CK(clk), .Q(\mem[118][2] ) );
  DFF_X1 \mem_reg[118][1]  ( .D(n25161), .CK(clk), .Q(\mem[118][1] ) );
  DFF_X1 \mem_reg[118][0]  ( .D(n25162), .CK(clk), .Q(\mem[118][0] ) );
  DFF_X1 \mem_reg[117][7]  ( .D(n25163), .CK(clk), .Q(\mem[117][7] ) );
  DFF_X1 \mem_reg[117][6]  ( .D(n25164), .CK(clk), .Q(\mem[117][6] ) );
  DFF_X1 \mem_reg[117][5]  ( .D(n25165), .CK(clk), .Q(\mem[117][5] ) );
  DFF_X1 \mem_reg[117][4]  ( .D(n25166), .CK(clk), .Q(\mem[117][4] ) );
  DFF_X1 \mem_reg[117][3]  ( .D(n25167), .CK(clk), .Q(\mem[117][3] ) );
  DFF_X1 \mem_reg[117][2]  ( .D(n25168), .CK(clk), .Q(\mem[117][2] ) );
  DFF_X1 \mem_reg[117][1]  ( .D(n25169), .CK(clk), .Q(\mem[117][1] ) );
  DFF_X1 \mem_reg[117][0]  ( .D(n25170), .CK(clk), .Q(\mem[117][0] ) );
  DFF_X1 \mem_reg[116][7]  ( .D(n25171), .CK(clk), .Q(\mem[116][7] ) );
  DFF_X1 \mem_reg[116][6]  ( .D(n25172), .CK(clk), .Q(\mem[116][6] ) );
  DFF_X1 \mem_reg[116][5]  ( .D(n25173), .CK(clk), .Q(\mem[116][5] ) );
  DFF_X1 \mem_reg[116][4]  ( .D(n25174), .CK(clk), .Q(\mem[116][4] ) );
  DFF_X1 \mem_reg[116][3]  ( .D(n25175), .CK(clk), .Q(\mem[116][3] ) );
  DFF_X1 \mem_reg[116][2]  ( .D(n25176), .CK(clk), .Q(\mem[116][2] ) );
  DFF_X1 \mem_reg[116][1]  ( .D(n25177), .CK(clk), .Q(\mem[116][1] ) );
  DFF_X1 \mem_reg[116][0]  ( .D(n25178), .CK(clk), .Q(\mem[116][0] ) );
  DFF_X1 \mem_reg[115][7]  ( .D(n25179), .CK(clk), .Q(\mem[115][7] ) );
  DFF_X1 \mem_reg[115][6]  ( .D(n25180), .CK(clk), .Q(\mem[115][6] ) );
  DFF_X1 \mem_reg[115][5]  ( .D(n25181), .CK(clk), .Q(\mem[115][5] ) );
  DFF_X1 \mem_reg[115][4]  ( .D(n25182), .CK(clk), .Q(\mem[115][4] ) );
  DFF_X1 \mem_reg[115][3]  ( .D(n25183), .CK(clk), .Q(\mem[115][3] ) );
  DFF_X1 \mem_reg[115][2]  ( .D(n25184), .CK(clk), .Q(\mem[115][2] ) );
  DFF_X1 \mem_reg[115][1]  ( .D(n25185), .CK(clk), .Q(\mem[115][1] ) );
  DFF_X1 \mem_reg[115][0]  ( .D(n25186), .CK(clk), .Q(\mem[115][0] ) );
  DFF_X1 \mem_reg[114][7]  ( .D(n25187), .CK(clk), .Q(\mem[114][7] ) );
  DFF_X1 \mem_reg[114][6]  ( .D(n25188), .CK(clk), .Q(\mem[114][6] ) );
  DFF_X1 \mem_reg[114][5]  ( .D(n25189), .CK(clk), .Q(\mem[114][5] ) );
  DFF_X1 \mem_reg[114][4]  ( .D(n25190), .CK(clk), .Q(\mem[114][4] ) );
  DFF_X1 \mem_reg[114][3]  ( .D(n25191), .CK(clk), .Q(\mem[114][3] ) );
  DFF_X1 \mem_reg[114][2]  ( .D(n25192), .CK(clk), .Q(\mem[114][2] ) );
  DFF_X1 \mem_reg[114][1]  ( .D(n25193), .CK(clk), .Q(\mem[114][1] ) );
  DFF_X1 \mem_reg[114][0]  ( .D(n25194), .CK(clk), .Q(\mem[114][0] ) );
  DFF_X1 \mem_reg[113][7]  ( .D(n25195), .CK(clk), .Q(\mem[113][7] ) );
  DFF_X1 \mem_reg[113][6]  ( .D(n25196), .CK(clk), .Q(\mem[113][6] ) );
  DFF_X1 \mem_reg[113][5]  ( .D(n25197), .CK(clk), .Q(\mem[113][5] ) );
  DFF_X1 \mem_reg[113][4]  ( .D(n25198), .CK(clk), .Q(\mem[113][4] ) );
  DFF_X1 \mem_reg[113][3]  ( .D(n25199), .CK(clk), .Q(\mem[113][3] ) );
  DFF_X1 \mem_reg[113][2]  ( .D(n25200), .CK(clk), .Q(\mem[113][2] ) );
  DFF_X1 \mem_reg[113][1]  ( .D(n25201), .CK(clk), .Q(\mem[113][1] ) );
  DFF_X1 \mem_reg[113][0]  ( .D(n25202), .CK(clk), .Q(\mem[113][0] ) );
  DFF_X1 \mem_reg[112][7]  ( .D(n25203), .CK(clk), .Q(\mem[112][7] ) );
  DFF_X1 \mem_reg[112][6]  ( .D(n25204), .CK(clk), .Q(\mem[112][6] ) );
  DFF_X1 \mem_reg[112][5]  ( .D(n25205), .CK(clk), .Q(\mem[112][5] ) );
  DFF_X1 \mem_reg[112][4]  ( .D(n25206), .CK(clk), .Q(\mem[112][4] ) );
  DFF_X1 \mem_reg[112][3]  ( .D(n25207), .CK(clk), .Q(\mem[112][3] ) );
  DFF_X1 \mem_reg[112][2]  ( .D(n25208), .CK(clk), .Q(\mem[112][2] ) );
  DFF_X1 \mem_reg[112][1]  ( .D(n25209), .CK(clk), .Q(\mem[112][1] ) );
  DFF_X1 \mem_reg[112][0]  ( .D(n25210), .CK(clk), .Q(\mem[112][0] ) );
  DFF_X1 \mem_reg[111][7]  ( .D(n25211), .CK(clk), .Q(\mem[111][7] ) );
  DFF_X1 \mem_reg[111][6]  ( .D(n25212), .CK(clk), .Q(\mem[111][6] ) );
  DFF_X1 \mem_reg[111][5]  ( .D(n25213), .CK(clk), .Q(\mem[111][5] ) );
  DFF_X1 \mem_reg[111][4]  ( .D(n25214), .CK(clk), .Q(\mem[111][4] ) );
  DFF_X1 \mem_reg[111][3]  ( .D(n25215), .CK(clk), .Q(\mem[111][3] ) );
  DFF_X1 \mem_reg[111][2]  ( .D(n25216), .CK(clk), .Q(\mem[111][2] ) );
  DFF_X1 \mem_reg[111][1]  ( .D(n25217), .CK(clk), .Q(\mem[111][1] ) );
  DFF_X1 \mem_reg[111][0]  ( .D(n25218), .CK(clk), .Q(\mem[111][0] ) );
  DFF_X1 \mem_reg[110][7]  ( .D(n25219), .CK(clk), .Q(\mem[110][7] ) );
  DFF_X1 \mem_reg[110][6]  ( .D(n25220), .CK(clk), .Q(\mem[110][6] ) );
  DFF_X1 \mem_reg[110][5]  ( .D(n25221), .CK(clk), .Q(\mem[110][5] ) );
  DFF_X1 \mem_reg[110][4]  ( .D(n25222), .CK(clk), .Q(\mem[110][4] ) );
  DFF_X1 \mem_reg[110][3]  ( .D(n25223), .CK(clk), .Q(\mem[110][3] ) );
  DFF_X1 \mem_reg[110][2]  ( .D(n25224), .CK(clk), .Q(\mem[110][2] ) );
  DFF_X1 \mem_reg[110][1]  ( .D(n25225), .CK(clk), .Q(\mem[110][1] ) );
  DFF_X1 \mem_reg[110][0]  ( .D(n25226), .CK(clk), .Q(\mem[110][0] ) );
  DFF_X1 \mem_reg[109][7]  ( .D(n25227), .CK(clk), .Q(\mem[109][7] ) );
  DFF_X1 \mem_reg[109][6]  ( .D(n25228), .CK(clk), .Q(\mem[109][6] ) );
  DFF_X1 \mem_reg[109][5]  ( .D(n25229), .CK(clk), .Q(\mem[109][5] ) );
  DFF_X1 \mem_reg[109][4]  ( .D(n25230), .CK(clk), .Q(\mem[109][4] ) );
  DFF_X1 \mem_reg[109][3]  ( .D(n25231), .CK(clk), .Q(\mem[109][3] ) );
  DFF_X1 \mem_reg[109][2]  ( .D(n25232), .CK(clk), .Q(\mem[109][2] ) );
  DFF_X1 \mem_reg[109][1]  ( .D(n25233), .CK(clk), .Q(\mem[109][1] ) );
  DFF_X1 \mem_reg[109][0]  ( .D(n25234), .CK(clk), .Q(\mem[109][0] ) );
  DFF_X1 \mem_reg[108][7]  ( .D(n25235), .CK(clk), .Q(\mem[108][7] ) );
  DFF_X1 \mem_reg[108][6]  ( .D(n25236), .CK(clk), .Q(\mem[108][6] ) );
  DFF_X1 \mem_reg[108][5]  ( .D(n25237), .CK(clk), .Q(\mem[108][5] ) );
  DFF_X1 \mem_reg[108][4]  ( .D(n25238), .CK(clk), .Q(\mem[108][4] ) );
  DFF_X1 \mem_reg[108][3]  ( .D(n25239), .CK(clk), .Q(\mem[108][3] ) );
  DFF_X1 \mem_reg[108][2]  ( .D(n25240), .CK(clk), .Q(\mem[108][2] ) );
  DFF_X1 \mem_reg[108][1]  ( .D(n25241), .CK(clk), .Q(\mem[108][1] ) );
  DFF_X1 \mem_reg[108][0]  ( .D(n25242), .CK(clk), .Q(\mem[108][0] ) );
  DFF_X1 \mem_reg[107][7]  ( .D(n25243), .CK(clk), .Q(\mem[107][7] ) );
  DFF_X1 \mem_reg[107][6]  ( .D(n25244), .CK(clk), .Q(\mem[107][6] ) );
  DFF_X1 \mem_reg[107][5]  ( .D(n25245), .CK(clk), .Q(\mem[107][5] ) );
  DFF_X1 \mem_reg[107][4]  ( .D(n25246), .CK(clk), .Q(\mem[107][4] ) );
  DFF_X1 \mem_reg[107][3]  ( .D(n25247), .CK(clk), .Q(\mem[107][3] ) );
  DFF_X1 \mem_reg[107][2]  ( .D(n25248), .CK(clk), .Q(\mem[107][2] ) );
  DFF_X1 \mem_reg[107][1]  ( .D(n25249), .CK(clk), .Q(\mem[107][1] ) );
  DFF_X1 \mem_reg[107][0]  ( .D(n25250), .CK(clk), .Q(\mem[107][0] ) );
  DFF_X1 \mem_reg[106][7]  ( .D(n25251), .CK(clk), .Q(\mem[106][7] ) );
  DFF_X1 \mem_reg[106][6]  ( .D(n25252), .CK(clk), .Q(\mem[106][6] ) );
  DFF_X1 \mem_reg[106][5]  ( .D(n25253), .CK(clk), .Q(\mem[106][5] ) );
  DFF_X1 \mem_reg[106][4]  ( .D(n25254), .CK(clk), .Q(\mem[106][4] ) );
  DFF_X1 \mem_reg[106][3]  ( .D(n25255), .CK(clk), .Q(\mem[106][3] ) );
  DFF_X1 \mem_reg[106][2]  ( .D(n25256), .CK(clk), .Q(\mem[106][2] ) );
  DFF_X1 \mem_reg[106][1]  ( .D(n25257), .CK(clk), .Q(\mem[106][1] ) );
  DFF_X1 \mem_reg[106][0]  ( .D(n25258), .CK(clk), .Q(\mem[106][0] ) );
  DFF_X1 \mem_reg[105][7]  ( .D(n25259), .CK(clk), .Q(\mem[105][7] ) );
  DFF_X1 \mem_reg[105][6]  ( .D(n25260), .CK(clk), .Q(\mem[105][6] ) );
  DFF_X1 \mem_reg[105][5]  ( .D(n25261), .CK(clk), .Q(\mem[105][5] ) );
  DFF_X1 \mem_reg[105][4]  ( .D(n25262), .CK(clk), .Q(\mem[105][4] ) );
  DFF_X1 \mem_reg[105][3]  ( .D(n25263), .CK(clk), .Q(\mem[105][3] ) );
  DFF_X1 \mem_reg[105][2]  ( .D(n25264), .CK(clk), .Q(\mem[105][2] ) );
  DFF_X1 \mem_reg[105][1]  ( .D(n25265), .CK(clk), .Q(\mem[105][1] ) );
  DFF_X1 \mem_reg[105][0]  ( .D(n25266), .CK(clk), .Q(\mem[105][0] ) );
  DFF_X1 \mem_reg[104][7]  ( .D(n25267), .CK(clk), .Q(\mem[104][7] ) );
  DFF_X1 \mem_reg[104][6]  ( .D(n25268), .CK(clk), .Q(\mem[104][6] ) );
  DFF_X1 \mem_reg[104][5]  ( .D(n25269), .CK(clk), .Q(\mem[104][5] ) );
  DFF_X1 \mem_reg[104][4]  ( .D(n25270), .CK(clk), .Q(\mem[104][4] ) );
  DFF_X1 \mem_reg[104][3]  ( .D(n25271), .CK(clk), .Q(\mem[104][3] ) );
  DFF_X1 \mem_reg[104][2]  ( .D(n25272), .CK(clk), .Q(\mem[104][2] ) );
  DFF_X1 \mem_reg[104][1]  ( .D(n25273), .CK(clk), .Q(\mem[104][1] ) );
  DFF_X1 \mem_reg[104][0]  ( .D(n25274), .CK(clk), .Q(\mem[104][0] ) );
  DFF_X1 \mem_reg[103][7]  ( .D(n25275), .CK(clk), .Q(\mem[103][7] ) );
  DFF_X1 \mem_reg[103][6]  ( .D(n25276), .CK(clk), .Q(\mem[103][6] ) );
  DFF_X1 \mem_reg[103][5]  ( .D(n25277), .CK(clk), .Q(\mem[103][5] ) );
  DFF_X1 \mem_reg[103][4]  ( .D(n25278), .CK(clk), .Q(\mem[103][4] ) );
  DFF_X1 \mem_reg[103][3]  ( .D(n25279), .CK(clk), .Q(\mem[103][3] ) );
  DFF_X1 \mem_reg[103][2]  ( .D(n25280), .CK(clk), .Q(\mem[103][2] ) );
  DFF_X1 \mem_reg[103][1]  ( .D(n25281), .CK(clk), .Q(\mem[103][1] ) );
  DFF_X1 \mem_reg[103][0]  ( .D(n25282), .CK(clk), .Q(\mem[103][0] ) );
  DFF_X1 \mem_reg[102][7]  ( .D(n25283), .CK(clk), .Q(\mem[102][7] ) );
  DFF_X1 \mem_reg[102][6]  ( .D(n25284), .CK(clk), .Q(\mem[102][6] ) );
  DFF_X1 \mem_reg[102][5]  ( .D(n25285), .CK(clk), .Q(\mem[102][5] ) );
  DFF_X1 \mem_reg[102][4]  ( .D(n25286), .CK(clk), .Q(\mem[102][4] ) );
  DFF_X1 \mem_reg[102][3]  ( .D(n25287), .CK(clk), .Q(\mem[102][3] ) );
  DFF_X1 \mem_reg[102][2]  ( .D(n25288), .CK(clk), .Q(\mem[102][2] ) );
  DFF_X1 \mem_reg[102][1]  ( .D(n25289), .CK(clk), .Q(\mem[102][1] ) );
  DFF_X1 \mem_reg[102][0]  ( .D(n25290), .CK(clk), .Q(\mem[102][0] ) );
  DFF_X1 \mem_reg[101][7]  ( .D(n25291), .CK(clk), .Q(\mem[101][7] ) );
  DFF_X1 \mem_reg[101][6]  ( .D(n25292), .CK(clk), .Q(\mem[101][6] ) );
  DFF_X1 \mem_reg[101][5]  ( .D(n25293), .CK(clk), .Q(\mem[101][5] ) );
  DFF_X1 \mem_reg[101][4]  ( .D(n25294), .CK(clk), .Q(\mem[101][4] ) );
  DFF_X1 \mem_reg[101][3]  ( .D(n25295), .CK(clk), .Q(\mem[101][3] ) );
  DFF_X1 \mem_reg[101][2]  ( .D(n25296), .CK(clk), .Q(\mem[101][2] ) );
  DFF_X1 \mem_reg[101][1]  ( .D(n25297), .CK(clk), .Q(\mem[101][1] ) );
  DFF_X1 \mem_reg[101][0]  ( .D(n25298), .CK(clk), .Q(\mem[101][0] ) );
  DFF_X1 \mem_reg[100][7]  ( .D(n25299), .CK(clk), .Q(\mem[100][7] ) );
  DFF_X1 \mem_reg[100][6]  ( .D(n25300), .CK(clk), .Q(\mem[100][6] ) );
  DFF_X1 \mem_reg[100][5]  ( .D(n25301), .CK(clk), .Q(\mem[100][5] ) );
  DFF_X1 \mem_reg[100][4]  ( .D(n25302), .CK(clk), .Q(\mem[100][4] ) );
  DFF_X1 \mem_reg[100][3]  ( .D(n25303), .CK(clk), .Q(\mem[100][3] ) );
  DFF_X1 \mem_reg[100][2]  ( .D(n25304), .CK(clk), .Q(\mem[100][2] ) );
  DFF_X1 \mem_reg[100][1]  ( .D(n25305), .CK(clk), .Q(\mem[100][1] ) );
  DFF_X1 \mem_reg[100][0]  ( .D(n25306), .CK(clk), .Q(\mem[100][0] ) );
  DFF_X1 \mem_reg[99][7]  ( .D(n25307), .CK(clk), .Q(\mem[99][7] ) );
  DFF_X1 \mem_reg[99][6]  ( .D(n25308), .CK(clk), .Q(\mem[99][6] ) );
  DFF_X1 \mem_reg[99][5]  ( .D(n25309), .CK(clk), .Q(\mem[99][5] ) );
  DFF_X1 \mem_reg[99][4]  ( .D(n25310), .CK(clk), .Q(\mem[99][4] ) );
  DFF_X1 \mem_reg[99][3]  ( .D(n25311), .CK(clk), .Q(\mem[99][3] ) );
  DFF_X1 \mem_reg[99][2]  ( .D(n25312), .CK(clk), .Q(\mem[99][2] ) );
  DFF_X1 \mem_reg[99][1]  ( .D(n25313), .CK(clk), .Q(\mem[99][1] ) );
  DFF_X1 \mem_reg[99][0]  ( .D(n25314), .CK(clk), .Q(\mem[99][0] ) );
  DFF_X1 \mem_reg[98][7]  ( .D(n25315), .CK(clk), .Q(\mem[98][7] ) );
  DFF_X1 \mem_reg[98][6]  ( .D(n25316), .CK(clk), .Q(\mem[98][6] ) );
  DFF_X1 \mem_reg[98][5]  ( .D(n25317), .CK(clk), .Q(\mem[98][5] ) );
  DFF_X1 \mem_reg[98][4]  ( .D(n25318), .CK(clk), .Q(\mem[98][4] ) );
  DFF_X1 \mem_reg[98][3]  ( .D(n25319), .CK(clk), .Q(\mem[98][3] ) );
  DFF_X1 \mem_reg[98][2]  ( .D(n25320), .CK(clk), .Q(\mem[98][2] ) );
  DFF_X1 \mem_reg[98][1]  ( .D(n25321), .CK(clk), .Q(\mem[98][1] ) );
  DFF_X1 \mem_reg[98][0]  ( .D(n25322), .CK(clk), .Q(\mem[98][0] ) );
  DFF_X1 \mem_reg[97][7]  ( .D(n25323), .CK(clk), .Q(\mem[97][7] ) );
  DFF_X1 \mem_reg[97][6]  ( .D(n25324), .CK(clk), .Q(\mem[97][6] ) );
  DFF_X1 \mem_reg[97][5]  ( .D(n25325), .CK(clk), .Q(\mem[97][5] ) );
  DFF_X1 \mem_reg[97][4]  ( .D(n25326), .CK(clk), .Q(\mem[97][4] ) );
  DFF_X1 \mem_reg[97][3]  ( .D(n25327), .CK(clk), .Q(\mem[97][3] ) );
  DFF_X1 \mem_reg[97][2]  ( .D(n25328), .CK(clk), .Q(\mem[97][2] ) );
  DFF_X1 \mem_reg[97][1]  ( .D(n25329), .CK(clk), .Q(\mem[97][1] ) );
  DFF_X1 \mem_reg[97][0]  ( .D(n25330), .CK(clk), .Q(\mem[97][0] ) );
  DFF_X1 \mem_reg[96][7]  ( .D(n25331), .CK(clk), .Q(\mem[96][7] ) );
  DFF_X1 \mem_reg[96][6]  ( .D(n25332), .CK(clk), .Q(\mem[96][6] ) );
  DFF_X1 \mem_reg[96][5]  ( .D(n25333), .CK(clk), .Q(\mem[96][5] ) );
  DFF_X1 \mem_reg[96][4]  ( .D(n25334), .CK(clk), .Q(\mem[96][4] ) );
  DFF_X1 \mem_reg[96][3]  ( .D(n25335), .CK(clk), .Q(\mem[96][3] ) );
  DFF_X1 \mem_reg[96][2]  ( .D(n25336), .CK(clk), .Q(\mem[96][2] ) );
  DFF_X1 \mem_reg[96][1]  ( .D(n25337), .CK(clk), .Q(\mem[96][1] ) );
  DFF_X1 \mem_reg[96][0]  ( .D(n25338), .CK(clk), .Q(\mem[96][0] ) );
  DFF_X1 \mem_reg[95][7]  ( .D(n25339), .CK(clk), .Q(\mem[95][7] ) );
  DFF_X1 \mem_reg[95][6]  ( .D(n25340), .CK(clk), .Q(\mem[95][6] ) );
  DFF_X1 \mem_reg[95][5]  ( .D(n25341), .CK(clk), .Q(\mem[95][5] ) );
  DFF_X1 \mem_reg[95][4]  ( .D(n25342), .CK(clk), .Q(\mem[95][4] ) );
  DFF_X1 \mem_reg[95][3]  ( .D(n25343), .CK(clk), .Q(\mem[95][3] ) );
  DFF_X1 \mem_reg[95][2]  ( .D(n25344), .CK(clk), .Q(\mem[95][2] ) );
  DFF_X1 \mem_reg[95][1]  ( .D(n25345), .CK(clk), .Q(\mem[95][1] ) );
  DFF_X1 \mem_reg[95][0]  ( .D(n25346), .CK(clk), .Q(\mem[95][0] ) );
  DFF_X1 \mem_reg[94][7]  ( .D(n25347), .CK(clk), .Q(\mem[94][7] ) );
  DFF_X1 \mem_reg[94][6]  ( .D(n25348), .CK(clk), .Q(\mem[94][6] ) );
  DFF_X1 \mem_reg[94][5]  ( .D(n25349), .CK(clk), .Q(\mem[94][5] ) );
  DFF_X1 \mem_reg[94][4]  ( .D(n25350), .CK(clk), .Q(\mem[94][4] ) );
  DFF_X1 \mem_reg[94][3]  ( .D(n25351), .CK(clk), .Q(\mem[94][3] ) );
  DFF_X1 \mem_reg[94][2]  ( .D(n25352), .CK(clk), .Q(\mem[94][2] ) );
  DFF_X1 \mem_reg[94][1]  ( .D(n25353), .CK(clk), .Q(\mem[94][1] ) );
  DFF_X1 \mem_reg[94][0]  ( .D(n25354), .CK(clk), .Q(\mem[94][0] ) );
  DFF_X1 \mem_reg[93][7]  ( .D(n25355), .CK(clk), .Q(\mem[93][7] ) );
  DFF_X1 \mem_reg[93][6]  ( .D(n25356), .CK(clk), .Q(\mem[93][6] ) );
  DFF_X1 \mem_reg[93][5]  ( .D(n25357), .CK(clk), .Q(\mem[93][5] ) );
  DFF_X1 \mem_reg[93][4]  ( .D(n25358), .CK(clk), .Q(\mem[93][4] ) );
  DFF_X1 \mem_reg[93][3]  ( .D(n25359), .CK(clk), .Q(\mem[93][3] ) );
  DFF_X1 \mem_reg[93][2]  ( .D(n25360), .CK(clk), .Q(\mem[93][2] ) );
  DFF_X1 \mem_reg[93][1]  ( .D(n25361), .CK(clk), .Q(\mem[93][1] ) );
  DFF_X1 \mem_reg[93][0]  ( .D(n25362), .CK(clk), .Q(\mem[93][0] ) );
  DFF_X1 \mem_reg[92][7]  ( .D(n25363), .CK(clk), .Q(\mem[92][7] ) );
  DFF_X1 \mem_reg[92][6]  ( .D(n25364), .CK(clk), .Q(\mem[92][6] ) );
  DFF_X1 \mem_reg[92][5]  ( .D(n25365), .CK(clk), .Q(\mem[92][5] ) );
  DFF_X1 \mem_reg[92][4]  ( .D(n25366), .CK(clk), .Q(\mem[92][4] ) );
  DFF_X1 \mem_reg[92][3]  ( .D(n25367), .CK(clk), .Q(\mem[92][3] ) );
  DFF_X1 \mem_reg[92][2]  ( .D(n25368), .CK(clk), .Q(\mem[92][2] ) );
  DFF_X1 \mem_reg[92][1]  ( .D(n25369), .CK(clk), .Q(\mem[92][1] ) );
  DFF_X1 \mem_reg[92][0]  ( .D(n25370), .CK(clk), .Q(\mem[92][0] ) );
  DFF_X1 \mem_reg[91][7]  ( .D(n25371), .CK(clk), .Q(\mem[91][7] ) );
  DFF_X1 \mem_reg[91][6]  ( .D(n25372), .CK(clk), .Q(\mem[91][6] ) );
  DFF_X1 \mem_reg[91][5]  ( .D(n25373), .CK(clk), .Q(\mem[91][5] ) );
  DFF_X1 \mem_reg[91][4]  ( .D(n25374), .CK(clk), .Q(\mem[91][4] ) );
  DFF_X1 \mem_reg[91][3]  ( .D(n25375), .CK(clk), .Q(\mem[91][3] ) );
  DFF_X1 \mem_reg[91][2]  ( .D(n25376), .CK(clk), .Q(\mem[91][2] ) );
  DFF_X1 \mem_reg[91][1]  ( .D(n25377), .CK(clk), .Q(\mem[91][1] ) );
  DFF_X1 \mem_reg[91][0]  ( .D(n25378), .CK(clk), .Q(\mem[91][0] ) );
  DFF_X1 \mem_reg[90][7]  ( .D(n25379), .CK(clk), .Q(\mem[90][7] ) );
  DFF_X1 \mem_reg[90][6]  ( .D(n25380), .CK(clk), .Q(\mem[90][6] ) );
  DFF_X1 \mem_reg[90][5]  ( .D(n25381), .CK(clk), .Q(\mem[90][5] ) );
  DFF_X1 \mem_reg[90][4]  ( .D(n25382), .CK(clk), .Q(\mem[90][4] ) );
  DFF_X1 \mem_reg[90][3]  ( .D(n25383), .CK(clk), .Q(\mem[90][3] ) );
  DFF_X1 \mem_reg[90][2]  ( .D(n25384), .CK(clk), .Q(\mem[90][2] ) );
  DFF_X1 \mem_reg[90][1]  ( .D(n25385), .CK(clk), .Q(\mem[90][1] ) );
  DFF_X1 \mem_reg[90][0]  ( .D(n25386), .CK(clk), .Q(\mem[90][0] ) );
  DFF_X1 \mem_reg[89][7]  ( .D(n25387), .CK(clk), .Q(\mem[89][7] ) );
  DFF_X1 \mem_reg[89][6]  ( .D(n25388), .CK(clk), .Q(\mem[89][6] ) );
  DFF_X1 \mem_reg[89][5]  ( .D(n25389), .CK(clk), .Q(\mem[89][5] ) );
  DFF_X1 \mem_reg[89][4]  ( .D(n25390), .CK(clk), .Q(\mem[89][4] ) );
  DFF_X1 \mem_reg[89][3]  ( .D(n25391), .CK(clk), .Q(\mem[89][3] ) );
  DFF_X1 \mem_reg[89][2]  ( .D(n25392), .CK(clk), .Q(\mem[89][2] ) );
  DFF_X1 \mem_reg[89][1]  ( .D(n25393), .CK(clk), .Q(\mem[89][1] ) );
  DFF_X1 \mem_reg[89][0]  ( .D(n25394), .CK(clk), .Q(\mem[89][0] ) );
  DFF_X1 \mem_reg[88][7]  ( .D(n25395), .CK(clk), .Q(\mem[88][7] ) );
  DFF_X1 \mem_reg[88][6]  ( .D(n25396), .CK(clk), .Q(\mem[88][6] ) );
  DFF_X1 \mem_reg[88][5]  ( .D(n25397), .CK(clk), .Q(\mem[88][5] ) );
  DFF_X1 \mem_reg[88][4]  ( .D(n25398), .CK(clk), .Q(\mem[88][4] ) );
  DFF_X1 \mem_reg[88][3]  ( .D(n25399), .CK(clk), .Q(\mem[88][3] ) );
  DFF_X1 \mem_reg[88][2]  ( .D(n25400), .CK(clk), .Q(\mem[88][2] ) );
  DFF_X1 \mem_reg[88][1]  ( .D(n25401), .CK(clk), .Q(\mem[88][1] ) );
  DFF_X1 \mem_reg[88][0]  ( .D(n25402), .CK(clk), .Q(\mem[88][0] ) );
  DFF_X1 \mem_reg[87][7]  ( .D(n25403), .CK(clk), .Q(\mem[87][7] ) );
  DFF_X1 \mem_reg[87][6]  ( .D(n25404), .CK(clk), .Q(\mem[87][6] ) );
  DFF_X1 \mem_reg[87][5]  ( .D(n25405), .CK(clk), .Q(\mem[87][5] ) );
  DFF_X1 \mem_reg[87][4]  ( .D(n25406), .CK(clk), .Q(\mem[87][4] ) );
  DFF_X1 \mem_reg[87][3]  ( .D(n25407), .CK(clk), .Q(\mem[87][3] ) );
  DFF_X1 \mem_reg[87][2]  ( .D(n25408), .CK(clk), .Q(\mem[87][2] ) );
  DFF_X1 \mem_reg[87][1]  ( .D(n25409), .CK(clk), .Q(\mem[87][1] ) );
  DFF_X1 \mem_reg[87][0]  ( .D(n25410), .CK(clk), .Q(\mem[87][0] ) );
  DFF_X1 \mem_reg[86][7]  ( .D(n25411), .CK(clk), .Q(\mem[86][7] ) );
  DFF_X1 \mem_reg[86][6]  ( .D(n25412), .CK(clk), .Q(\mem[86][6] ) );
  DFF_X1 \mem_reg[86][5]  ( .D(n25413), .CK(clk), .Q(\mem[86][5] ) );
  DFF_X1 \mem_reg[86][4]  ( .D(n25414), .CK(clk), .Q(\mem[86][4] ) );
  DFF_X1 \mem_reg[86][3]  ( .D(n25415), .CK(clk), .Q(\mem[86][3] ) );
  DFF_X1 \mem_reg[86][2]  ( .D(n25416), .CK(clk), .Q(\mem[86][2] ) );
  DFF_X1 \mem_reg[86][1]  ( .D(n25417), .CK(clk), .Q(\mem[86][1] ) );
  DFF_X1 \mem_reg[86][0]  ( .D(n25418), .CK(clk), .Q(\mem[86][0] ) );
  DFF_X1 \mem_reg[85][7]  ( .D(n25419), .CK(clk), .Q(\mem[85][7] ) );
  DFF_X1 \mem_reg[85][6]  ( .D(n25420), .CK(clk), .Q(\mem[85][6] ) );
  DFF_X1 \mem_reg[85][5]  ( .D(n25421), .CK(clk), .Q(\mem[85][5] ) );
  DFF_X1 \mem_reg[85][4]  ( .D(n25422), .CK(clk), .Q(\mem[85][4] ) );
  DFF_X1 \mem_reg[85][3]  ( .D(n25423), .CK(clk), .Q(\mem[85][3] ) );
  DFF_X1 \mem_reg[85][2]  ( .D(n25424), .CK(clk), .Q(\mem[85][2] ) );
  DFF_X1 \mem_reg[85][1]  ( .D(n25425), .CK(clk), .Q(\mem[85][1] ) );
  DFF_X1 \mem_reg[85][0]  ( .D(n25426), .CK(clk), .Q(\mem[85][0] ) );
  DFF_X1 \mem_reg[84][7]  ( .D(n25427), .CK(clk), .Q(\mem[84][7] ) );
  DFF_X1 \mem_reg[84][6]  ( .D(n25428), .CK(clk), .Q(\mem[84][6] ) );
  DFF_X1 \mem_reg[84][5]  ( .D(n25429), .CK(clk), .Q(\mem[84][5] ) );
  DFF_X1 \mem_reg[84][4]  ( .D(n25430), .CK(clk), .Q(\mem[84][4] ) );
  DFF_X1 \mem_reg[84][3]  ( .D(n25431), .CK(clk), .Q(\mem[84][3] ) );
  DFF_X1 \mem_reg[84][2]  ( .D(n25432), .CK(clk), .Q(\mem[84][2] ) );
  DFF_X1 \mem_reg[84][1]  ( .D(n25433), .CK(clk), .Q(\mem[84][1] ) );
  DFF_X1 \mem_reg[84][0]  ( .D(n25434), .CK(clk), .Q(\mem[84][0] ) );
  DFF_X1 \mem_reg[83][7]  ( .D(n25435), .CK(clk), .Q(\mem[83][7] ) );
  DFF_X1 \mem_reg[83][6]  ( .D(n25436), .CK(clk), .Q(\mem[83][6] ) );
  DFF_X1 \mem_reg[83][5]  ( .D(n25437), .CK(clk), .Q(\mem[83][5] ) );
  DFF_X1 \mem_reg[83][4]  ( .D(n25438), .CK(clk), .Q(\mem[83][4] ) );
  DFF_X1 \mem_reg[83][3]  ( .D(n25439), .CK(clk), .Q(\mem[83][3] ) );
  DFF_X1 \mem_reg[83][2]  ( .D(n25440), .CK(clk), .Q(\mem[83][2] ) );
  DFF_X1 \mem_reg[83][1]  ( .D(n25441), .CK(clk), .Q(\mem[83][1] ) );
  DFF_X1 \mem_reg[83][0]  ( .D(n25442), .CK(clk), .Q(\mem[83][0] ) );
  DFF_X1 \mem_reg[82][7]  ( .D(n25443), .CK(clk), .Q(\mem[82][7] ) );
  DFF_X1 \mem_reg[82][6]  ( .D(n25444), .CK(clk), .Q(\mem[82][6] ) );
  DFF_X1 \mem_reg[82][5]  ( .D(n25445), .CK(clk), .Q(\mem[82][5] ) );
  DFF_X1 \mem_reg[82][4]  ( .D(n25446), .CK(clk), .Q(\mem[82][4] ) );
  DFF_X1 \mem_reg[82][3]  ( .D(n25447), .CK(clk), .Q(\mem[82][3] ) );
  DFF_X1 \mem_reg[82][2]  ( .D(n25448), .CK(clk), .Q(\mem[82][2] ) );
  DFF_X1 \mem_reg[82][1]  ( .D(n25449), .CK(clk), .Q(\mem[82][1] ) );
  DFF_X1 \mem_reg[82][0]  ( .D(n25450), .CK(clk), .Q(\mem[82][0] ) );
  DFF_X1 \mem_reg[81][7]  ( .D(n25451), .CK(clk), .Q(\mem[81][7] ) );
  DFF_X1 \mem_reg[81][6]  ( .D(n25452), .CK(clk), .Q(\mem[81][6] ) );
  DFF_X1 \mem_reg[81][5]  ( .D(n25453), .CK(clk), .Q(\mem[81][5] ) );
  DFF_X1 \mem_reg[81][4]  ( .D(n25454), .CK(clk), .Q(\mem[81][4] ) );
  DFF_X1 \mem_reg[81][3]  ( .D(n25455), .CK(clk), .Q(\mem[81][3] ) );
  DFF_X1 \mem_reg[81][2]  ( .D(n25456), .CK(clk), .Q(\mem[81][2] ) );
  DFF_X1 \mem_reg[81][1]  ( .D(n25457), .CK(clk), .Q(\mem[81][1] ) );
  DFF_X1 \mem_reg[81][0]  ( .D(n25458), .CK(clk), .Q(\mem[81][0] ) );
  DFF_X1 \mem_reg[80][7]  ( .D(n25459), .CK(clk), .Q(\mem[80][7] ) );
  DFF_X1 \mem_reg[80][6]  ( .D(n25460), .CK(clk), .Q(\mem[80][6] ) );
  DFF_X1 \mem_reg[80][5]  ( .D(n25461), .CK(clk), .Q(\mem[80][5] ) );
  DFF_X1 \mem_reg[80][4]  ( .D(n25462), .CK(clk), .Q(\mem[80][4] ) );
  DFF_X1 \mem_reg[80][3]  ( .D(n25463), .CK(clk), .Q(\mem[80][3] ) );
  DFF_X1 \mem_reg[80][2]  ( .D(n25464), .CK(clk), .Q(\mem[80][2] ) );
  DFF_X1 \mem_reg[80][1]  ( .D(n25465), .CK(clk), .Q(\mem[80][1] ) );
  DFF_X1 \mem_reg[80][0]  ( .D(n25466), .CK(clk), .Q(\mem[80][0] ) );
  DFF_X1 \mem_reg[79][7]  ( .D(n25467), .CK(clk), .Q(\mem[79][7] ) );
  DFF_X1 \mem_reg[79][6]  ( .D(n25468), .CK(clk), .Q(\mem[79][6] ) );
  DFF_X1 \mem_reg[79][5]  ( .D(n25469), .CK(clk), .Q(\mem[79][5] ) );
  DFF_X1 \mem_reg[79][4]  ( .D(n25470), .CK(clk), .Q(\mem[79][4] ) );
  DFF_X1 \mem_reg[79][3]  ( .D(n25471), .CK(clk), .Q(\mem[79][3] ) );
  DFF_X1 \mem_reg[79][2]  ( .D(n25472), .CK(clk), .Q(\mem[79][2] ) );
  DFF_X1 \mem_reg[79][1]  ( .D(n25473), .CK(clk), .Q(\mem[79][1] ) );
  DFF_X1 \mem_reg[79][0]  ( .D(n25474), .CK(clk), .Q(\mem[79][0] ) );
  DFF_X1 \mem_reg[78][7]  ( .D(n25475), .CK(clk), .Q(\mem[78][7] ) );
  DFF_X1 \mem_reg[78][6]  ( .D(n25476), .CK(clk), .Q(\mem[78][6] ) );
  DFF_X1 \mem_reg[78][5]  ( .D(n25477), .CK(clk), .Q(\mem[78][5] ) );
  DFF_X1 \mem_reg[78][4]  ( .D(n25478), .CK(clk), .Q(\mem[78][4] ) );
  DFF_X1 \mem_reg[78][3]  ( .D(n25479), .CK(clk), .Q(\mem[78][3] ) );
  DFF_X1 \mem_reg[78][2]  ( .D(n25480), .CK(clk), .Q(\mem[78][2] ) );
  DFF_X1 \mem_reg[78][1]  ( .D(n25481), .CK(clk), .Q(\mem[78][1] ) );
  DFF_X1 \mem_reg[78][0]  ( .D(n25482), .CK(clk), .Q(\mem[78][0] ) );
  DFF_X1 \mem_reg[77][7]  ( .D(n25483), .CK(clk), .Q(\mem[77][7] ) );
  DFF_X1 \mem_reg[77][6]  ( .D(n25484), .CK(clk), .Q(\mem[77][6] ) );
  DFF_X1 \mem_reg[77][5]  ( .D(n25485), .CK(clk), .Q(\mem[77][5] ) );
  DFF_X1 \mem_reg[77][4]  ( .D(n25486), .CK(clk), .Q(\mem[77][4] ) );
  DFF_X1 \mem_reg[77][3]  ( .D(n25487), .CK(clk), .Q(\mem[77][3] ) );
  DFF_X1 \mem_reg[77][2]  ( .D(n25488), .CK(clk), .Q(\mem[77][2] ) );
  DFF_X1 \mem_reg[77][1]  ( .D(n25489), .CK(clk), .Q(\mem[77][1] ) );
  DFF_X1 \mem_reg[77][0]  ( .D(n25490), .CK(clk), .Q(\mem[77][0] ) );
  DFF_X1 \mem_reg[76][7]  ( .D(n25491), .CK(clk), .Q(\mem[76][7] ) );
  DFF_X1 \mem_reg[76][6]  ( .D(n25492), .CK(clk), .Q(\mem[76][6] ) );
  DFF_X1 \mem_reg[76][5]  ( .D(n25493), .CK(clk), .Q(\mem[76][5] ) );
  DFF_X1 \mem_reg[76][4]  ( .D(n25494), .CK(clk), .Q(\mem[76][4] ) );
  DFF_X1 \mem_reg[76][3]  ( .D(n25495), .CK(clk), .Q(\mem[76][3] ) );
  DFF_X1 \mem_reg[76][2]  ( .D(n25496), .CK(clk), .Q(\mem[76][2] ) );
  DFF_X1 \mem_reg[76][1]  ( .D(n25497), .CK(clk), .Q(\mem[76][1] ) );
  DFF_X1 \mem_reg[76][0]  ( .D(n25498), .CK(clk), .Q(\mem[76][0] ) );
  DFF_X1 \mem_reg[75][7]  ( .D(n25499), .CK(clk), .Q(\mem[75][7] ) );
  DFF_X1 \mem_reg[75][6]  ( .D(n25500), .CK(clk), .Q(\mem[75][6] ) );
  DFF_X1 \mem_reg[75][5]  ( .D(n25501), .CK(clk), .Q(\mem[75][5] ) );
  DFF_X1 \mem_reg[75][4]  ( .D(n25502), .CK(clk), .Q(\mem[75][4] ) );
  DFF_X1 \mem_reg[75][3]  ( .D(n25503), .CK(clk), .Q(\mem[75][3] ) );
  DFF_X1 \mem_reg[75][2]  ( .D(n25504), .CK(clk), .Q(\mem[75][2] ) );
  DFF_X1 \mem_reg[75][1]  ( .D(n25505), .CK(clk), .Q(\mem[75][1] ) );
  DFF_X1 \mem_reg[75][0]  ( .D(n25506), .CK(clk), .Q(\mem[75][0] ) );
  DFF_X1 \mem_reg[74][7]  ( .D(n25507), .CK(clk), .Q(\mem[74][7] ) );
  DFF_X1 \mem_reg[74][6]  ( .D(n25508), .CK(clk), .Q(\mem[74][6] ) );
  DFF_X1 \mem_reg[74][5]  ( .D(n25509), .CK(clk), .Q(\mem[74][5] ) );
  DFF_X1 \mem_reg[74][4]  ( .D(n25510), .CK(clk), .Q(\mem[74][4] ) );
  DFF_X1 \mem_reg[74][3]  ( .D(n25511), .CK(clk), .Q(\mem[74][3] ) );
  DFF_X1 \mem_reg[74][2]  ( .D(n25512), .CK(clk), .Q(\mem[74][2] ) );
  DFF_X1 \mem_reg[74][1]  ( .D(n25513), .CK(clk), .Q(\mem[74][1] ) );
  DFF_X1 \mem_reg[74][0]  ( .D(n25514), .CK(clk), .Q(\mem[74][0] ) );
  DFF_X1 \mem_reg[73][7]  ( .D(n25515), .CK(clk), .Q(\mem[73][7] ) );
  DFF_X1 \mem_reg[73][6]  ( .D(n25516), .CK(clk), .Q(\mem[73][6] ) );
  DFF_X1 \mem_reg[73][5]  ( .D(n25517), .CK(clk), .Q(\mem[73][5] ) );
  DFF_X1 \mem_reg[73][4]  ( .D(n25518), .CK(clk), .Q(\mem[73][4] ) );
  DFF_X1 \mem_reg[73][3]  ( .D(n25519), .CK(clk), .Q(\mem[73][3] ) );
  DFF_X1 \mem_reg[73][2]  ( .D(n25520), .CK(clk), .Q(\mem[73][2] ) );
  DFF_X1 \mem_reg[73][1]  ( .D(n25521), .CK(clk), .Q(\mem[73][1] ) );
  DFF_X1 \mem_reg[73][0]  ( .D(n25522), .CK(clk), .Q(\mem[73][0] ) );
  DFF_X1 \mem_reg[72][7]  ( .D(n25523), .CK(clk), .Q(\mem[72][7] ) );
  DFF_X1 \mem_reg[72][6]  ( .D(n25524), .CK(clk), .Q(\mem[72][6] ) );
  DFF_X1 \mem_reg[72][5]  ( .D(n25525), .CK(clk), .Q(\mem[72][5] ) );
  DFF_X1 \mem_reg[72][4]  ( .D(n25526), .CK(clk), .Q(\mem[72][4] ) );
  DFF_X1 \mem_reg[72][3]  ( .D(n25527), .CK(clk), .Q(\mem[72][3] ) );
  DFF_X1 \mem_reg[72][2]  ( .D(n25528), .CK(clk), .Q(\mem[72][2] ) );
  DFF_X1 \mem_reg[72][1]  ( .D(n25529), .CK(clk), .Q(\mem[72][1] ) );
  DFF_X1 \mem_reg[72][0]  ( .D(n25530), .CK(clk), .Q(\mem[72][0] ) );
  DFF_X1 \mem_reg[71][7]  ( .D(n25531), .CK(clk), .Q(\mem[71][7] ) );
  DFF_X1 \mem_reg[71][6]  ( .D(n25532), .CK(clk), .Q(\mem[71][6] ) );
  DFF_X1 \mem_reg[71][5]  ( .D(n25533), .CK(clk), .Q(\mem[71][5] ) );
  DFF_X1 \mem_reg[71][4]  ( .D(n25534), .CK(clk), .Q(\mem[71][4] ) );
  DFF_X1 \mem_reg[71][3]  ( .D(n25535), .CK(clk), .Q(\mem[71][3] ) );
  DFF_X1 \mem_reg[71][2]  ( .D(n25536), .CK(clk), .Q(\mem[71][2] ) );
  DFF_X1 \mem_reg[71][1]  ( .D(n25537), .CK(clk), .Q(\mem[71][1] ) );
  DFF_X1 \mem_reg[71][0]  ( .D(n25538), .CK(clk), .Q(\mem[71][0] ) );
  DFF_X1 \mem_reg[70][7]  ( .D(n25539), .CK(clk), .Q(\mem[70][7] ) );
  DFF_X1 \mem_reg[70][6]  ( .D(n25540), .CK(clk), .Q(\mem[70][6] ) );
  DFF_X1 \mem_reg[70][5]  ( .D(n25541), .CK(clk), .Q(\mem[70][5] ) );
  DFF_X1 \mem_reg[70][4]  ( .D(n25542), .CK(clk), .Q(\mem[70][4] ) );
  DFF_X1 \mem_reg[70][3]  ( .D(n25543), .CK(clk), .Q(\mem[70][3] ) );
  DFF_X1 \mem_reg[70][2]  ( .D(n25544), .CK(clk), .Q(\mem[70][2] ) );
  DFF_X1 \mem_reg[70][1]  ( .D(n25545), .CK(clk), .Q(\mem[70][1] ) );
  DFF_X1 \mem_reg[70][0]  ( .D(n25546), .CK(clk), .Q(\mem[70][0] ) );
  DFF_X1 \mem_reg[69][7]  ( .D(n25547), .CK(clk), .Q(\mem[69][7] ) );
  DFF_X1 \mem_reg[69][6]  ( .D(n25548), .CK(clk), .Q(\mem[69][6] ) );
  DFF_X1 \mem_reg[69][5]  ( .D(n25549), .CK(clk), .Q(\mem[69][5] ) );
  DFF_X1 \mem_reg[69][4]  ( .D(n25550), .CK(clk), .Q(\mem[69][4] ) );
  DFF_X1 \mem_reg[69][3]  ( .D(n25551), .CK(clk), .Q(\mem[69][3] ) );
  DFF_X1 \mem_reg[69][2]  ( .D(n25552), .CK(clk), .Q(\mem[69][2] ) );
  DFF_X1 \mem_reg[69][1]  ( .D(n25553), .CK(clk), .Q(\mem[69][1] ) );
  DFF_X1 \mem_reg[69][0]  ( .D(n25554), .CK(clk), .Q(\mem[69][0] ) );
  DFF_X1 \mem_reg[68][7]  ( .D(n25555), .CK(clk), .Q(\mem[68][7] ) );
  DFF_X1 \mem_reg[68][6]  ( .D(n25556), .CK(clk), .Q(\mem[68][6] ) );
  DFF_X1 \mem_reg[68][5]  ( .D(n25557), .CK(clk), .Q(\mem[68][5] ) );
  DFF_X1 \mem_reg[68][4]  ( .D(n25558), .CK(clk), .Q(\mem[68][4] ) );
  DFF_X1 \mem_reg[68][3]  ( .D(n25559), .CK(clk), .Q(\mem[68][3] ) );
  DFF_X1 \mem_reg[68][2]  ( .D(n25560), .CK(clk), .Q(\mem[68][2] ) );
  DFF_X1 \mem_reg[68][1]  ( .D(n25561), .CK(clk), .Q(\mem[68][1] ) );
  DFF_X1 \mem_reg[68][0]  ( .D(n25562), .CK(clk), .Q(\mem[68][0] ) );
  DFF_X1 \mem_reg[67][7]  ( .D(n25563), .CK(clk), .Q(\mem[67][7] ) );
  DFF_X1 \mem_reg[67][6]  ( .D(n25564), .CK(clk), .Q(\mem[67][6] ) );
  DFF_X1 \mem_reg[67][5]  ( .D(n25565), .CK(clk), .Q(\mem[67][5] ) );
  DFF_X1 \mem_reg[67][4]  ( .D(n25566), .CK(clk), .Q(\mem[67][4] ) );
  DFF_X1 \mem_reg[67][3]  ( .D(n25567), .CK(clk), .Q(\mem[67][3] ) );
  DFF_X1 \mem_reg[67][2]  ( .D(n25568), .CK(clk), .Q(\mem[67][2] ) );
  DFF_X1 \mem_reg[67][1]  ( .D(n25569), .CK(clk), .Q(\mem[67][1] ) );
  DFF_X1 \mem_reg[67][0]  ( .D(n25570), .CK(clk), .Q(\mem[67][0] ) );
  DFF_X1 \mem_reg[66][7]  ( .D(n25571), .CK(clk), .Q(\mem[66][7] ) );
  DFF_X1 \mem_reg[66][6]  ( .D(n25572), .CK(clk), .Q(\mem[66][6] ) );
  DFF_X1 \mem_reg[66][5]  ( .D(n25573), .CK(clk), .Q(\mem[66][5] ) );
  DFF_X1 \mem_reg[66][4]  ( .D(n25574), .CK(clk), .Q(\mem[66][4] ) );
  DFF_X1 \mem_reg[66][3]  ( .D(n25575), .CK(clk), .Q(\mem[66][3] ) );
  DFF_X1 \mem_reg[66][2]  ( .D(n25576), .CK(clk), .Q(\mem[66][2] ) );
  DFF_X1 \mem_reg[66][1]  ( .D(n25577), .CK(clk), .Q(\mem[66][1] ) );
  DFF_X1 \mem_reg[66][0]  ( .D(n25578), .CK(clk), .Q(\mem[66][0] ) );
  DFF_X1 \mem_reg[65][7]  ( .D(n25579), .CK(clk), .Q(\mem[65][7] ) );
  DFF_X1 \mem_reg[65][6]  ( .D(n25580), .CK(clk), .Q(\mem[65][6] ) );
  DFF_X1 \mem_reg[65][5]  ( .D(n25581), .CK(clk), .Q(\mem[65][5] ) );
  DFF_X1 \mem_reg[65][4]  ( .D(n25582), .CK(clk), .Q(\mem[65][4] ) );
  DFF_X1 \mem_reg[65][3]  ( .D(n25583), .CK(clk), .Q(\mem[65][3] ) );
  DFF_X1 \mem_reg[65][2]  ( .D(n25584), .CK(clk), .Q(\mem[65][2] ) );
  DFF_X1 \mem_reg[65][1]  ( .D(n25585), .CK(clk), .Q(\mem[65][1] ) );
  DFF_X1 \mem_reg[65][0]  ( .D(n25586), .CK(clk), .Q(\mem[65][0] ) );
  DFF_X1 \mem_reg[64][7]  ( .D(n25587), .CK(clk), .Q(\mem[64][7] ) );
  DFF_X1 \mem_reg[64][6]  ( .D(n25588), .CK(clk), .Q(\mem[64][6] ) );
  DFF_X1 \mem_reg[64][5]  ( .D(n25589), .CK(clk), .Q(\mem[64][5] ) );
  DFF_X1 \mem_reg[64][4]  ( .D(n25590), .CK(clk), .Q(\mem[64][4] ) );
  DFF_X1 \mem_reg[64][3]  ( .D(n25591), .CK(clk), .Q(\mem[64][3] ) );
  DFF_X1 \mem_reg[64][2]  ( .D(n25592), .CK(clk), .Q(\mem[64][2] ) );
  DFF_X1 \mem_reg[64][1]  ( .D(n25593), .CK(clk), .Q(\mem[64][1] ) );
  DFF_X1 \mem_reg[64][0]  ( .D(n25594), .CK(clk), .Q(\mem[64][0] ) );
  DFF_X1 \mem_reg[63][7]  ( .D(n25595), .CK(clk), .Q(\mem[63][7] ) );
  DFF_X1 \mem_reg[63][6]  ( .D(n25596), .CK(clk), .Q(\mem[63][6] ) );
  DFF_X1 \mem_reg[63][5]  ( .D(n25597), .CK(clk), .Q(\mem[63][5] ) );
  DFF_X1 \mem_reg[63][4]  ( .D(n25598), .CK(clk), .Q(\mem[63][4] ) );
  DFF_X1 \mem_reg[63][3]  ( .D(n25599), .CK(clk), .Q(\mem[63][3] ) );
  DFF_X1 \mem_reg[63][2]  ( .D(n25600), .CK(clk), .Q(\mem[63][2] ) );
  DFF_X1 \mem_reg[63][1]  ( .D(n25601), .CK(clk), .Q(\mem[63][1] ) );
  DFF_X1 \mem_reg[63][0]  ( .D(n25602), .CK(clk), .Q(\mem[63][0] ) );
  DFF_X1 \mem_reg[62][7]  ( .D(n25603), .CK(clk), .Q(\mem[62][7] ) );
  DFF_X1 \mem_reg[62][6]  ( .D(n25604), .CK(clk), .Q(\mem[62][6] ) );
  DFF_X1 \mem_reg[62][5]  ( .D(n25605), .CK(clk), .Q(\mem[62][5] ) );
  DFF_X1 \mem_reg[62][4]  ( .D(n25606), .CK(clk), .Q(\mem[62][4] ) );
  DFF_X1 \mem_reg[62][3]  ( .D(n25607), .CK(clk), .Q(\mem[62][3] ) );
  DFF_X1 \mem_reg[62][2]  ( .D(n25608), .CK(clk), .Q(\mem[62][2] ) );
  DFF_X1 \mem_reg[62][1]  ( .D(n25609), .CK(clk), .Q(\mem[62][1] ) );
  DFF_X1 \mem_reg[62][0]  ( .D(n25610), .CK(clk), .Q(\mem[62][0] ) );
  DFF_X1 \mem_reg[61][7]  ( .D(n25611), .CK(clk), .Q(\mem[61][7] ) );
  DFF_X1 \mem_reg[61][6]  ( .D(n25612), .CK(clk), .Q(\mem[61][6] ) );
  DFF_X1 \mem_reg[61][5]  ( .D(n25613), .CK(clk), .Q(\mem[61][5] ) );
  DFF_X1 \mem_reg[61][4]  ( .D(n25614), .CK(clk), .Q(\mem[61][4] ) );
  DFF_X1 \mem_reg[61][3]  ( .D(n25615), .CK(clk), .Q(\mem[61][3] ) );
  DFF_X1 \mem_reg[61][2]  ( .D(n25616), .CK(clk), .Q(\mem[61][2] ) );
  DFF_X1 \mem_reg[61][1]  ( .D(n25617), .CK(clk), .Q(\mem[61][1] ) );
  DFF_X1 \mem_reg[61][0]  ( .D(n25618), .CK(clk), .Q(\mem[61][0] ) );
  DFF_X1 \mem_reg[60][7]  ( .D(n25619), .CK(clk), .Q(\mem[60][7] ) );
  DFF_X1 \mem_reg[60][6]  ( .D(n25620), .CK(clk), .Q(\mem[60][6] ) );
  DFF_X1 \mem_reg[60][5]  ( .D(n25621), .CK(clk), .Q(\mem[60][5] ) );
  DFF_X1 \mem_reg[60][4]  ( .D(n25622), .CK(clk), .Q(\mem[60][4] ) );
  DFF_X1 \mem_reg[60][3]  ( .D(n25623), .CK(clk), .Q(\mem[60][3] ) );
  DFF_X1 \mem_reg[60][2]  ( .D(n25624), .CK(clk), .Q(\mem[60][2] ) );
  DFF_X1 \mem_reg[60][1]  ( .D(n25625), .CK(clk), .Q(\mem[60][1] ) );
  DFF_X1 \mem_reg[60][0]  ( .D(n25626), .CK(clk), .Q(\mem[60][0] ) );
  DFF_X1 \mem_reg[59][7]  ( .D(n25627), .CK(clk), .Q(\mem[59][7] ) );
  DFF_X1 \mem_reg[59][6]  ( .D(n25628), .CK(clk), .Q(\mem[59][6] ) );
  DFF_X1 \mem_reg[59][5]  ( .D(n25629), .CK(clk), .Q(\mem[59][5] ) );
  DFF_X1 \mem_reg[59][4]  ( .D(n25630), .CK(clk), .Q(\mem[59][4] ) );
  DFF_X1 \mem_reg[59][3]  ( .D(n25631), .CK(clk), .Q(\mem[59][3] ) );
  DFF_X1 \mem_reg[59][2]  ( .D(n25632), .CK(clk), .Q(\mem[59][2] ) );
  DFF_X1 \mem_reg[59][1]  ( .D(n25633), .CK(clk), .Q(\mem[59][1] ) );
  DFF_X1 \mem_reg[59][0]  ( .D(n25634), .CK(clk), .Q(\mem[59][0] ) );
  DFF_X1 \mem_reg[58][7]  ( .D(n25635), .CK(clk), .Q(\mem[58][7] ) );
  DFF_X1 \mem_reg[58][6]  ( .D(n25636), .CK(clk), .Q(\mem[58][6] ) );
  DFF_X1 \mem_reg[58][5]  ( .D(n25637), .CK(clk), .Q(\mem[58][5] ) );
  DFF_X1 \mem_reg[58][4]  ( .D(n25638), .CK(clk), .Q(\mem[58][4] ) );
  DFF_X1 \mem_reg[58][3]  ( .D(n25639), .CK(clk), .Q(\mem[58][3] ) );
  DFF_X1 \mem_reg[58][2]  ( .D(n25640), .CK(clk), .Q(\mem[58][2] ) );
  DFF_X1 \mem_reg[58][1]  ( .D(n25641), .CK(clk), .Q(\mem[58][1] ) );
  DFF_X1 \mem_reg[58][0]  ( .D(n25642), .CK(clk), .Q(\mem[58][0] ) );
  DFF_X1 \mem_reg[57][7]  ( .D(n25643), .CK(clk), .Q(\mem[57][7] ) );
  DFF_X1 \mem_reg[57][6]  ( .D(n25644), .CK(clk), .Q(\mem[57][6] ) );
  DFF_X1 \mem_reg[57][5]  ( .D(n25645), .CK(clk), .Q(\mem[57][5] ) );
  DFF_X1 \mem_reg[57][4]  ( .D(n25646), .CK(clk), .Q(\mem[57][4] ) );
  DFF_X1 \mem_reg[57][3]  ( .D(n25647), .CK(clk), .Q(\mem[57][3] ) );
  DFF_X1 \mem_reg[57][2]  ( .D(n25648), .CK(clk), .Q(\mem[57][2] ) );
  DFF_X1 \mem_reg[57][1]  ( .D(n25649), .CK(clk), .Q(\mem[57][1] ) );
  DFF_X1 \mem_reg[57][0]  ( .D(n25650), .CK(clk), .Q(\mem[57][0] ) );
  DFF_X1 \mem_reg[56][7]  ( .D(n25651), .CK(clk), .Q(\mem[56][7] ) );
  DFF_X1 \mem_reg[56][6]  ( .D(n25652), .CK(clk), .Q(\mem[56][6] ) );
  DFF_X1 \mem_reg[56][5]  ( .D(n25653), .CK(clk), .Q(\mem[56][5] ) );
  DFF_X1 \mem_reg[56][4]  ( .D(n25654), .CK(clk), .Q(\mem[56][4] ) );
  DFF_X1 \mem_reg[56][3]  ( .D(n25655), .CK(clk), .Q(\mem[56][3] ) );
  DFF_X1 \mem_reg[56][2]  ( .D(n25656), .CK(clk), .Q(\mem[56][2] ) );
  DFF_X1 \mem_reg[56][1]  ( .D(n25657), .CK(clk), .Q(\mem[56][1] ) );
  DFF_X1 \mem_reg[56][0]  ( .D(n25658), .CK(clk), .Q(\mem[56][0] ) );
  DFF_X1 \mem_reg[55][7]  ( .D(n25659), .CK(clk), .Q(\mem[55][7] ) );
  DFF_X1 \mem_reg[55][6]  ( .D(n25660), .CK(clk), .Q(\mem[55][6] ) );
  DFF_X1 \mem_reg[55][5]  ( .D(n25661), .CK(clk), .Q(\mem[55][5] ) );
  DFF_X1 \mem_reg[55][4]  ( .D(n25662), .CK(clk), .Q(\mem[55][4] ) );
  DFF_X1 \mem_reg[55][3]  ( .D(n25663), .CK(clk), .Q(\mem[55][3] ) );
  DFF_X1 \mem_reg[55][2]  ( .D(n25664), .CK(clk), .Q(\mem[55][2] ) );
  DFF_X1 \mem_reg[55][1]  ( .D(n25665), .CK(clk), .Q(\mem[55][1] ) );
  DFF_X1 \mem_reg[55][0]  ( .D(n25666), .CK(clk), .Q(\mem[55][0] ) );
  DFF_X1 \mem_reg[54][7]  ( .D(n25667), .CK(clk), .Q(\mem[54][7] ) );
  DFF_X1 \mem_reg[54][6]  ( .D(n25668), .CK(clk), .Q(\mem[54][6] ) );
  DFF_X1 \mem_reg[54][5]  ( .D(n25669), .CK(clk), .Q(\mem[54][5] ) );
  DFF_X1 \mem_reg[54][4]  ( .D(n25670), .CK(clk), .Q(\mem[54][4] ) );
  DFF_X1 \mem_reg[54][3]  ( .D(n25671), .CK(clk), .Q(\mem[54][3] ) );
  DFF_X1 \mem_reg[54][2]  ( .D(n25672), .CK(clk), .Q(\mem[54][2] ) );
  DFF_X1 \mem_reg[54][1]  ( .D(n25673), .CK(clk), .Q(\mem[54][1] ) );
  DFF_X1 \mem_reg[54][0]  ( .D(n25674), .CK(clk), .Q(\mem[54][0] ) );
  DFF_X1 \mem_reg[53][7]  ( .D(n25675), .CK(clk), .Q(\mem[53][7] ) );
  DFF_X1 \mem_reg[53][6]  ( .D(n25676), .CK(clk), .Q(\mem[53][6] ) );
  DFF_X1 \mem_reg[53][5]  ( .D(n25677), .CK(clk), .Q(\mem[53][5] ) );
  DFF_X1 \mem_reg[53][4]  ( .D(n25678), .CK(clk), .Q(\mem[53][4] ) );
  DFF_X1 \mem_reg[53][3]  ( .D(n25679), .CK(clk), .Q(\mem[53][3] ) );
  DFF_X1 \mem_reg[53][2]  ( .D(n25680), .CK(clk), .Q(\mem[53][2] ) );
  DFF_X1 \mem_reg[53][1]  ( .D(n25681), .CK(clk), .Q(\mem[53][1] ) );
  DFF_X1 \mem_reg[53][0]  ( .D(n25682), .CK(clk), .Q(\mem[53][0] ) );
  DFF_X1 \mem_reg[52][7]  ( .D(n25683), .CK(clk), .Q(\mem[52][7] ) );
  DFF_X1 \mem_reg[52][6]  ( .D(n25684), .CK(clk), .Q(\mem[52][6] ) );
  DFF_X1 \mem_reg[52][5]  ( .D(n25685), .CK(clk), .Q(\mem[52][5] ) );
  DFF_X1 \mem_reg[52][4]  ( .D(n25686), .CK(clk), .Q(\mem[52][4] ) );
  DFF_X1 \mem_reg[52][3]  ( .D(n25687), .CK(clk), .Q(\mem[52][3] ) );
  DFF_X1 \mem_reg[52][2]  ( .D(n25688), .CK(clk), .Q(\mem[52][2] ) );
  DFF_X1 \mem_reg[52][1]  ( .D(n25689), .CK(clk), .Q(\mem[52][1] ) );
  DFF_X1 \mem_reg[52][0]  ( .D(n25690), .CK(clk), .Q(\mem[52][0] ) );
  DFF_X1 \mem_reg[51][7]  ( .D(n25691), .CK(clk), .Q(\mem[51][7] ) );
  DFF_X1 \mem_reg[51][6]  ( .D(n25692), .CK(clk), .Q(\mem[51][6] ) );
  DFF_X1 \mem_reg[51][5]  ( .D(n25693), .CK(clk), .Q(\mem[51][5] ) );
  DFF_X1 \mem_reg[51][4]  ( .D(n25694), .CK(clk), .Q(\mem[51][4] ) );
  DFF_X1 \mem_reg[51][3]  ( .D(n25695), .CK(clk), .Q(\mem[51][3] ) );
  DFF_X1 \mem_reg[51][2]  ( .D(n25696), .CK(clk), .Q(\mem[51][2] ) );
  DFF_X1 \mem_reg[51][1]  ( .D(n25697), .CK(clk), .Q(\mem[51][1] ) );
  DFF_X1 \mem_reg[51][0]  ( .D(n25698), .CK(clk), .Q(\mem[51][0] ) );
  DFF_X1 \mem_reg[50][7]  ( .D(n25699), .CK(clk), .Q(\mem[50][7] ) );
  DFF_X1 \mem_reg[50][6]  ( .D(n25700), .CK(clk), .Q(\mem[50][6] ) );
  DFF_X1 \mem_reg[50][5]  ( .D(n25701), .CK(clk), .Q(\mem[50][5] ) );
  DFF_X1 \mem_reg[50][4]  ( .D(n25702), .CK(clk), .Q(\mem[50][4] ) );
  DFF_X1 \mem_reg[50][3]  ( .D(n25703), .CK(clk), .Q(\mem[50][3] ) );
  DFF_X1 \mem_reg[50][2]  ( .D(n25704), .CK(clk), .Q(\mem[50][2] ) );
  DFF_X1 \mem_reg[50][1]  ( .D(n25705), .CK(clk), .Q(\mem[50][1] ) );
  DFF_X1 \mem_reg[50][0]  ( .D(n25706), .CK(clk), .Q(\mem[50][0] ) );
  DFF_X1 \mem_reg[49][7]  ( .D(n25707), .CK(clk), .Q(\mem[49][7] ) );
  DFF_X1 \mem_reg[49][6]  ( .D(n25708), .CK(clk), .Q(\mem[49][6] ) );
  DFF_X1 \mem_reg[49][5]  ( .D(n25709), .CK(clk), .Q(\mem[49][5] ) );
  DFF_X1 \mem_reg[49][4]  ( .D(n25710), .CK(clk), .Q(\mem[49][4] ) );
  DFF_X1 \mem_reg[49][3]  ( .D(n25711), .CK(clk), .Q(\mem[49][3] ) );
  DFF_X1 \mem_reg[49][2]  ( .D(n25712), .CK(clk), .Q(\mem[49][2] ) );
  DFF_X1 \mem_reg[49][1]  ( .D(n25713), .CK(clk), .Q(\mem[49][1] ) );
  DFF_X1 \mem_reg[49][0]  ( .D(n25714), .CK(clk), .Q(\mem[49][0] ) );
  DFF_X1 \mem_reg[48][7]  ( .D(n25715), .CK(clk), .Q(\mem[48][7] ) );
  DFF_X1 \mem_reg[48][6]  ( .D(n25716), .CK(clk), .Q(\mem[48][6] ) );
  DFF_X1 \mem_reg[48][5]  ( .D(n25717), .CK(clk), .Q(\mem[48][5] ) );
  DFF_X1 \mem_reg[48][4]  ( .D(n25718), .CK(clk), .Q(\mem[48][4] ) );
  DFF_X1 \mem_reg[48][3]  ( .D(n25719), .CK(clk), .Q(\mem[48][3] ) );
  DFF_X1 \mem_reg[48][2]  ( .D(n25720), .CK(clk), .Q(\mem[48][2] ) );
  DFF_X1 \mem_reg[48][1]  ( .D(n25721), .CK(clk), .Q(\mem[48][1] ) );
  DFF_X1 \mem_reg[48][0]  ( .D(n25722), .CK(clk), .Q(\mem[48][0] ) );
  DFF_X1 \mem_reg[47][7]  ( .D(n25723), .CK(clk), .Q(\mem[47][7] ) );
  DFF_X1 \mem_reg[47][6]  ( .D(n25724), .CK(clk), .Q(\mem[47][6] ) );
  DFF_X1 \mem_reg[47][5]  ( .D(n25725), .CK(clk), .Q(\mem[47][5] ) );
  DFF_X1 \mem_reg[47][4]  ( .D(n25726), .CK(clk), .Q(\mem[47][4] ) );
  DFF_X1 \mem_reg[47][3]  ( .D(n25727), .CK(clk), .Q(\mem[47][3] ) );
  DFF_X1 \mem_reg[47][2]  ( .D(n25728), .CK(clk), .Q(\mem[47][2] ) );
  DFF_X1 \mem_reg[47][1]  ( .D(n25729), .CK(clk), .Q(\mem[47][1] ) );
  DFF_X1 \mem_reg[47][0]  ( .D(n25730), .CK(clk), .Q(\mem[47][0] ) );
  DFF_X1 \mem_reg[46][7]  ( .D(n25731), .CK(clk), .Q(\mem[46][7] ) );
  DFF_X1 \mem_reg[46][6]  ( .D(n25732), .CK(clk), .Q(\mem[46][6] ) );
  DFF_X1 \mem_reg[46][5]  ( .D(n25733), .CK(clk), .Q(\mem[46][5] ) );
  DFF_X1 \mem_reg[46][4]  ( .D(n25734), .CK(clk), .Q(\mem[46][4] ) );
  DFF_X1 \mem_reg[46][3]  ( .D(n25735), .CK(clk), .Q(\mem[46][3] ) );
  DFF_X1 \mem_reg[46][2]  ( .D(n25736), .CK(clk), .Q(\mem[46][2] ) );
  DFF_X1 \mem_reg[46][1]  ( .D(n25737), .CK(clk), .Q(\mem[46][1] ) );
  DFF_X1 \mem_reg[46][0]  ( .D(n25738), .CK(clk), .Q(\mem[46][0] ) );
  DFF_X1 \mem_reg[45][7]  ( .D(n25739), .CK(clk), .Q(\mem[45][7] ) );
  DFF_X1 \mem_reg[45][6]  ( .D(n25740), .CK(clk), .Q(\mem[45][6] ) );
  DFF_X1 \mem_reg[45][5]  ( .D(n25741), .CK(clk), .Q(\mem[45][5] ) );
  DFF_X1 \mem_reg[45][4]  ( .D(n25742), .CK(clk), .Q(\mem[45][4] ) );
  DFF_X1 \mem_reg[45][3]  ( .D(n25743), .CK(clk), .Q(\mem[45][3] ) );
  DFF_X1 \mem_reg[45][2]  ( .D(n25744), .CK(clk), .Q(\mem[45][2] ) );
  DFF_X1 \mem_reg[45][1]  ( .D(n25745), .CK(clk), .Q(\mem[45][1] ) );
  DFF_X1 \mem_reg[45][0]  ( .D(n25746), .CK(clk), .Q(\mem[45][0] ) );
  DFF_X1 \mem_reg[44][7]  ( .D(n25747), .CK(clk), .Q(\mem[44][7] ) );
  DFF_X1 \mem_reg[44][6]  ( .D(n25748), .CK(clk), .Q(\mem[44][6] ) );
  DFF_X1 \mem_reg[44][5]  ( .D(n25749), .CK(clk), .Q(\mem[44][5] ) );
  DFF_X1 \mem_reg[44][4]  ( .D(n25750), .CK(clk), .Q(\mem[44][4] ) );
  DFF_X1 \mem_reg[44][3]  ( .D(n25751), .CK(clk), .Q(\mem[44][3] ) );
  DFF_X1 \mem_reg[44][2]  ( .D(n25752), .CK(clk), .Q(\mem[44][2] ) );
  DFF_X1 \mem_reg[44][1]  ( .D(n25753), .CK(clk), .Q(\mem[44][1] ) );
  DFF_X1 \mem_reg[44][0]  ( .D(n25754), .CK(clk), .Q(\mem[44][0] ) );
  DFF_X1 \mem_reg[43][7]  ( .D(n25755), .CK(clk), .Q(\mem[43][7] ) );
  DFF_X1 \mem_reg[43][6]  ( .D(n25756), .CK(clk), .Q(\mem[43][6] ) );
  DFF_X1 \mem_reg[43][5]  ( .D(n25757), .CK(clk), .Q(\mem[43][5] ) );
  DFF_X1 \mem_reg[43][4]  ( .D(n25758), .CK(clk), .Q(\mem[43][4] ) );
  DFF_X1 \mem_reg[43][3]  ( .D(n25759), .CK(clk), .Q(\mem[43][3] ) );
  DFF_X1 \mem_reg[43][2]  ( .D(n25760), .CK(clk), .Q(\mem[43][2] ) );
  DFF_X1 \mem_reg[43][1]  ( .D(n25761), .CK(clk), .Q(\mem[43][1] ) );
  DFF_X1 \mem_reg[43][0]  ( .D(n25762), .CK(clk), .Q(\mem[43][0] ) );
  DFF_X1 \mem_reg[42][7]  ( .D(n25763), .CK(clk), .Q(\mem[42][7] ) );
  DFF_X1 \mem_reg[42][6]  ( .D(n25764), .CK(clk), .Q(\mem[42][6] ) );
  DFF_X1 \mem_reg[42][5]  ( .D(n25765), .CK(clk), .Q(\mem[42][5] ) );
  DFF_X1 \mem_reg[42][4]  ( .D(n25766), .CK(clk), .Q(\mem[42][4] ) );
  DFF_X1 \mem_reg[42][3]  ( .D(n25767), .CK(clk), .Q(\mem[42][3] ) );
  DFF_X1 \mem_reg[42][2]  ( .D(n25768), .CK(clk), .Q(\mem[42][2] ) );
  DFF_X1 \mem_reg[42][1]  ( .D(n25769), .CK(clk), .Q(\mem[42][1] ) );
  DFF_X1 \mem_reg[42][0]  ( .D(n25770), .CK(clk), .Q(\mem[42][0] ) );
  DFF_X1 \mem_reg[41][7]  ( .D(n25771), .CK(clk), .Q(\mem[41][7] ) );
  DFF_X1 \mem_reg[41][6]  ( .D(n25772), .CK(clk), .Q(\mem[41][6] ) );
  DFF_X1 \mem_reg[41][5]  ( .D(n25773), .CK(clk), .Q(\mem[41][5] ) );
  DFF_X1 \mem_reg[41][4]  ( .D(n25774), .CK(clk), .Q(\mem[41][4] ) );
  DFF_X1 \mem_reg[41][3]  ( .D(n25775), .CK(clk), .Q(\mem[41][3] ) );
  DFF_X1 \mem_reg[41][2]  ( .D(n25776), .CK(clk), .Q(\mem[41][2] ) );
  DFF_X1 \mem_reg[41][1]  ( .D(n25777), .CK(clk), .Q(\mem[41][1] ) );
  DFF_X1 \mem_reg[41][0]  ( .D(n25778), .CK(clk), .Q(\mem[41][0] ) );
  DFF_X1 \mem_reg[40][7]  ( .D(n25779), .CK(clk), .Q(\mem[40][7] ) );
  DFF_X1 \mem_reg[40][6]  ( .D(n25780), .CK(clk), .Q(\mem[40][6] ) );
  DFF_X1 \mem_reg[40][5]  ( .D(n25781), .CK(clk), .Q(\mem[40][5] ) );
  DFF_X1 \mem_reg[40][4]  ( .D(n25782), .CK(clk), .Q(\mem[40][4] ) );
  DFF_X1 \mem_reg[40][3]  ( .D(n25783), .CK(clk), .Q(\mem[40][3] ) );
  DFF_X1 \mem_reg[40][2]  ( .D(n25784), .CK(clk), .Q(\mem[40][2] ) );
  DFF_X1 \mem_reg[40][1]  ( .D(n25785), .CK(clk), .Q(\mem[40][1] ) );
  DFF_X1 \mem_reg[40][0]  ( .D(n25786), .CK(clk), .Q(\mem[40][0] ) );
  DFF_X1 \mem_reg[39][7]  ( .D(n25787), .CK(clk), .Q(\mem[39][7] ) );
  DFF_X1 \mem_reg[39][6]  ( .D(n25788), .CK(clk), .Q(\mem[39][6] ) );
  DFF_X1 \mem_reg[39][5]  ( .D(n25789), .CK(clk), .Q(\mem[39][5] ) );
  DFF_X1 \mem_reg[39][4]  ( .D(n25790), .CK(clk), .Q(\mem[39][4] ) );
  DFF_X1 \mem_reg[39][3]  ( .D(n25791), .CK(clk), .Q(\mem[39][3] ) );
  DFF_X1 \mem_reg[39][2]  ( .D(n25792), .CK(clk), .Q(\mem[39][2] ) );
  DFF_X1 \mem_reg[39][1]  ( .D(n25793), .CK(clk), .Q(\mem[39][1] ) );
  DFF_X1 \mem_reg[39][0]  ( .D(n25794), .CK(clk), .Q(\mem[39][0] ) );
  DFF_X1 \mem_reg[38][7]  ( .D(n25795), .CK(clk), .Q(\mem[38][7] ) );
  DFF_X1 \mem_reg[38][6]  ( .D(n25796), .CK(clk), .Q(\mem[38][6] ) );
  DFF_X1 \mem_reg[38][5]  ( .D(n25797), .CK(clk), .Q(\mem[38][5] ) );
  DFF_X1 \mem_reg[38][4]  ( .D(n25798), .CK(clk), .Q(\mem[38][4] ) );
  DFF_X1 \mem_reg[38][3]  ( .D(n25799), .CK(clk), .Q(\mem[38][3] ) );
  DFF_X1 \mem_reg[38][2]  ( .D(n25800), .CK(clk), .Q(\mem[38][2] ) );
  DFF_X1 \mem_reg[38][1]  ( .D(n25801), .CK(clk), .Q(\mem[38][1] ) );
  DFF_X1 \mem_reg[38][0]  ( .D(n25802), .CK(clk), .Q(\mem[38][0] ) );
  DFF_X1 \mem_reg[37][7]  ( .D(n25803), .CK(clk), .Q(\mem[37][7] ) );
  DFF_X1 \mem_reg[37][6]  ( .D(n25804), .CK(clk), .Q(\mem[37][6] ) );
  DFF_X1 \mem_reg[37][5]  ( .D(n25805), .CK(clk), .Q(\mem[37][5] ) );
  DFF_X1 \mem_reg[37][4]  ( .D(n25806), .CK(clk), .Q(\mem[37][4] ) );
  DFF_X1 \mem_reg[37][3]  ( .D(n25807), .CK(clk), .Q(\mem[37][3] ) );
  DFF_X1 \mem_reg[37][2]  ( .D(n25808), .CK(clk), .Q(\mem[37][2] ) );
  DFF_X1 \mem_reg[37][1]  ( .D(n25809), .CK(clk), .Q(\mem[37][1] ) );
  DFF_X1 \mem_reg[37][0]  ( .D(n25810), .CK(clk), .Q(\mem[37][0] ) );
  DFF_X1 \mem_reg[36][7]  ( .D(n25811), .CK(clk), .Q(\mem[36][7] ) );
  DFF_X1 \mem_reg[36][6]  ( .D(n25812), .CK(clk), .Q(\mem[36][6] ) );
  DFF_X1 \mem_reg[36][5]  ( .D(n25813), .CK(clk), .Q(\mem[36][5] ) );
  DFF_X1 \mem_reg[36][4]  ( .D(n25814), .CK(clk), .Q(\mem[36][4] ) );
  DFF_X1 \mem_reg[36][3]  ( .D(n25815), .CK(clk), .Q(\mem[36][3] ) );
  DFF_X1 \mem_reg[36][2]  ( .D(n25816), .CK(clk), .Q(\mem[36][2] ) );
  DFF_X1 \mem_reg[36][1]  ( .D(n25817), .CK(clk), .Q(\mem[36][1] ) );
  DFF_X1 \mem_reg[36][0]  ( .D(n25818), .CK(clk), .Q(\mem[36][0] ) );
  DFF_X1 \mem_reg[35][7]  ( .D(n25819), .CK(clk), .Q(\mem[35][7] ) );
  DFF_X1 \mem_reg[35][6]  ( .D(n25820), .CK(clk), .Q(\mem[35][6] ) );
  DFF_X1 \mem_reg[35][5]  ( .D(n25821), .CK(clk), .Q(\mem[35][5] ) );
  DFF_X1 \mem_reg[35][4]  ( .D(n25822), .CK(clk), .Q(\mem[35][4] ) );
  DFF_X1 \mem_reg[35][3]  ( .D(n25823), .CK(clk), .Q(\mem[35][3] ) );
  DFF_X1 \mem_reg[35][2]  ( .D(n25824), .CK(clk), .Q(\mem[35][2] ) );
  DFF_X1 \mem_reg[35][1]  ( .D(n25825), .CK(clk), .Q(\mem[35][1] ) );
  DFF_X1 \mem_reg[35][0]  ( .D(n25826), .CK(clk), .Q(\mem[35][0] ) );
  DFF_X1 \mem_reg[34][7]  ( .D(n25827), .CK(clk), .Q(\mem[34][7] ) );
  DFF_X1 \mem_reg[34][6]  ( .D(n25828), .CK(clk), .Q(\mem[34][6] ) );
  DFF_X1 \mem_reg[34][5]  ( .D(n25829), .CK(clk), .Q(\mem[34][5] ) );
  DFF_X1 \mem_reg[34][4]  ( .D(n25830), .CK(clk), .Q(\mem[34][4] ) );
  DFF_X1 \mem_reg[34][3]  ( .D(n25831), .CK(clk), .Q(\mem[34][3] ) );
  DFF_X1 \mem_reg[34][2]  ( .D(n25832), .CK(clk), .Q(\mem[34][2] ) );
  DFF_X1 \mem_reg[34][1]  ( .D(n25833), .CK(clk), .Q(\mem[34][1] ) );
  DFF_X1 \mem_reg[34][0]  ( .D(n25834), .CK(clk), .Q(\mem[34][0] ) );
  DFF_X1 \mem_reg[33][7]  ( .D(n25835), .CK(clk), .Q(\mem[33][7] ) );
  DFF_X1 \mem_reg[33][6]  ( .D(n25836), .CK(clk), .Q(\mem[33][6] ) );
  DFF_X1 \mem_reg[33][5]  ( .D(n25837), .CK(clk), .Q(\mem[33][5] ) );
  DFF_X1 \mem_reg[33][4]  ( .D(n25838), .CK(clk), .Q(\mem[33][4] ) );
  DFF_X1 \mem_reg[33][3]  ( .D(n25839), .CK(clk), .Q(\mem[33][3] ) );
  DFF_X1 \mem_reg[33][2]  ( .D(n25840), .CK(clk), .Q(\mem[33][2] ) );
  DFF_X1 \mem_reg[33][1]  ( .D(n25841), .CK(clk), .Q(\mem[33][1] ) );
  DFF_X1 \mem_reg[33][0]  ( .D(n25842), .CK(clk), .Q(\mem[33][0] ) );
  DFF_X1 \mem_reg[32][7]  ( .D(n25843), .CK(clk), .Q(\mem[32][7] ) );
  DFF_X1 \mem_reg[32][6]  ( .D(n25844), .CK(clk), .Q(\mem[32][6] ) );
  DFF_X1 \mem_reg[32][5]  ( .D(n25845), .CK(clk), .Q(\mem[32][5] ) );
  DFF_X1 \mem_reg[32][4]  ( .D(n25846), .CK(clk), .Q(\mem[32][4] ) );
  DFF_X1 \mem_reg[32][3]  ( .D(n25847), .CK(clk), .Q(\mem[32][3] ) );
  DFF_X1 \mem_reg[32][2]  ( .D(n25848), .CK(clk), .Q(\mem[32][2] ) );
  DFF_X1 \mem_reg[32][1]  ( .D(n25849), .CK(clk), .Q(\mem[32][1] ) );
  DFF_X1 \mem_reg[32][0]  ( .D(n25850), .CK(clk), .Q(\mem[32][0] ) );
  DFF_X1 \mem_reg[31][7]  ( .D(n25851), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n25852), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n25853), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n25854), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n25855), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n25856), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n25857), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n25858), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n25859), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n25860), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n25861), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n25862), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n25863), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n25864), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n25865), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n25866), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n25867), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n25868), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n25869), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n25870), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n25871), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n25872), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n25873), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n25874), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n25875), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n25876), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n25877), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n25878), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n25879), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n25880), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n25881), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n25882), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n25883), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n25884), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n25885), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n25886), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n25887), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n25888), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n25889), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n25890), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n25891), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n25892), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n25893), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n25894), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n25895), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n25896), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n25897), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n25898), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n25899), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n25900), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n25901), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n25902), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n25903), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n25904), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n25905), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n25906), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n25907), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n25908), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n25909), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n25910), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n25911), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n25912), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n25913), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n25914), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n25915), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n25916), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n25917), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n25918), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n25919), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n25920), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n25921), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n25922), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n25923), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n25924), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n25925), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n25926), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n25927), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n25928), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n25929), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n25930), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n25931), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n25932), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n25933), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n25934), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n25935), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n25936), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n25937), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n25938), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n25939), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n25940), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n25941), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n25942), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n25943), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n25944), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n25945), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n25946), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n25947), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n25948), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n25949), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n25950), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n25951), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n25952), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n25953), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n25954), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n25955), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n25956), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n25957), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n25958), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n25959), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n25960), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n25961), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n25962), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n25963), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n25964), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n25965), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n25966), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n25967), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n25968), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n25969), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n25970), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n25971), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n25972), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n25973), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n25974), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n25975), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n25976), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n25977), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n25978), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n25979), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n25980), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n25981), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n25982), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n25983), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n25984), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n25985), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n25986), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n25987), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n25988), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n25989), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n25990), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n25991), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n25992), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n25993), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n25994), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n25995), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n25996), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n25997), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n25998), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n25999), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n26000), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n26001), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n26002), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n26003), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n26004), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n26005), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n26006), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n26007), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n26008), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n26009), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n26010), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n26011), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n26012), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n26013), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n26014), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n26015), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n26016), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n26017), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n26018), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n26019), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n26020), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n26021), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n26022), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n26023), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n26024), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n26025), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n26026), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n26027), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n26028), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n26029), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n26030), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n26031), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n26032), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n26033), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n26034), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n26035), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n26036), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n26037), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n26038), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n26039), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n26040), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n26041), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n26042), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n26043), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n26044), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n26045), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n26046), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n26047), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n26048), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n26049), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n26050), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n26051), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n26052), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n26053), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n26054), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n26055), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n26056), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n26057), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n26058), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n26059), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n26060), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n26061), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n26062), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n26063), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n26064), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n26065), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n26066), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n26067), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n26068), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n26069), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n26070), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n26071), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n26072), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n26073), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n26074), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n26075), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n26076), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n26077), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n26078), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n26079), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n26080), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n26081), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n26082), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n26083), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n26084), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n26085), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n26086), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n26087), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n26088), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n26089), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n26090), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n26091), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n26092), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n26093), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n26094), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n26095), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n26096), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n26097), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n26098), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n26099), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n26100), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n26101), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n26102), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n26103), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n26104), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n26105), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n26106), .CK(clk), .Q(\mem[0][0] ) );
  BUF_X1 U3 ( .A(n8508), .Z(n8409) );
  BUF_X1 U4 ( .A(n8516), .Z(n8410) );
  BUF_X1 U5 ( .A(n8385), .Z(n8414) );
  BUF_X1 U6 ( .A(n8385), .Z(n8415) );
  BUF_X1 U7 ( .A(n8385), .Z(n8416) );
  BUF_X1 U8 ( .A(n8384), .Z(n8420) );
  BUF_X1 U9 ( .A(n8384), .Z(n8421) );
  BUF_X1 U10 ( .A(n8384), .Z(n8422) );
  BUF_X1 U11 ( .A(n8383), .Z(n8426) );
  BUF_X1 U12 ( .A(n8383), .Z(n8427) );
  BUF_X1 U13 ( .A(n8383), .Z(n8428) );
  BUF_X1 U14 ( .A(n8382), .Z(n8432) );
  BUF_X1 U15 ( .A(n8382), .Z(n8433) );
  BUF_X1 U16 ( .A(n8382), .Z(n8434) );
  BUF_X1 U17 ( .A(n8381), .Z(n8438) );
  BUF_X1 U18 ( .A(n8381), .Z(n8439) );
  BUF_X1 U19 ( .A(n8381), .Z(n8440) );
  BUF_X1 U20 ( .A(n8380), .Z(n8444) );
  BUF_X1 U21 ( .A(n8380), .Z(n8445) );
  BUF_X1 U22 ( .A(n8380), .Z(n8446) );
  BUF_X1 U23 ( .A(n8379), .Z(n8450) );
  BUF_X1 U24 ( .A(n8379), .Z(n8451) );
  BUF_X1 U25 ( .A(n8379), .Z(n8452) );
  BUF_X1 U26 ( .A(n8378), .Z(n8456) );
  BUF_X1 U27 ( .A(n8378), .Z(n8457) );
  BUF_X1 U28 ( .A(n8378), .Z(n8458) );
  BUF_X1 U29 ( .A(n8377), .Z(n8462) );
  BUF_X1 U30 ( .A(n8377), .Z(n8463) );
  BUF_X1 U31 ( .A(n8377), .Z(n8464) );
  BUF_X1 U32 ( .A(n8376), .Z(n8468) );
  BUF_X1 U33 ( .A(n8376), .Z(n8469) );
  BUF_X1 U34 ( .A(n8376), .Z(n8470) );
  BUF_X1 U35 ( .A(n8375), .Z(n8474) );
  BUF_X1 U36 ( .A(n8375), .Z(n8475) );
  BUF_X1 U37 ( .A(n8375), .Z(n8476) );
  BUF_X1 U38 ( .A(n8374), .Z(n8480) );
  BUF_X1 U39 ( .A(n8374), .Z(n8481) );
  BUF_X1 U40 ( .A(n8374), .Z(n8482) );
  BUF_X1 U41 ( .A(n8373), .Z(n8486) );
  BUF_X1 U42 ( .A(n8373), .Z(n8487) );
  BUF_X1 U43 ( .A(n8373), .Z(n8488) );
  BUF_X1 U44 ( .A(n8372), .Z(n8492) );
  BUF_X1 U45 ( .A(n8372), .Z(n8493) );
  BUF_X1 U46 ( .A(n8372), .Z(n8494) );
  BUF_X1 U47 ( .A(n8371), .Z(n8498) );
  BUF_X1 U48 ( .A(n8371), .Z(n8499) );
  BUF_X1 U49 ( .A(n8371), .Z(n8500) );
  BUF_X1 U50 ( .A(n8370), .Z(n8504) );
  BUF_X1 U51 ( .A(n8370), .Z(n8505) );
  BUF_X1 U52 ( .A(n8370), .Z(n8506) );
  BUF_X1 U53 ( .A(n8369), .Z(n8510) );
  BUF_X1 U54 ( .A(n8369), .Z(n8511) );
  BUF_X1 U55 ( .A(n8369), .Z(n8512) );
  BUF_X1 U56 ( .A(n8368), .Z(n8516) );
  BUF_X1 U57 ( .A(n8368), .Z(n8517) );
  BUF_X1 U58 ( .A(n8368), .Z(n8518) );
  BUF_X1 U59 ( .A(n8367), .Z(n8522) );
  BUF_X1 U60 ( .A(n8367), .Z(n8523) );
  BUF_X1 U61 ( .A(n8367), .Z(n8524) );
  BUF_X1 U62 ( .A(n8366), .Z(n8528) );
  BUF_X1 U63 ( .A(n8366), .Z(n8529) );
  BUF_X1 U64 ( .A(n8366), .Z(n8530) );
  BUF_X1 U65 ( .A(n8365), .Z(n8534) );
  BUF_X1 U66 ( .A(n8365), .Z(n8535) );
  BUF_X1 U67 ( .A(n8365), .Z(n8536) );
  BUF_X1 U68 ( .A(n8321), .Z(n8283) );
  BUF_X1 U69 ( .A(n8281), .Z(n8290) );
  BUF_X1 U70 ( .A(n8281), .Z(n8291) );
  BUF_X1 U71 ( .A(n8281), .Z(n8292) );
  BUF_X1 U72 ( .A(n8280), .Z(n8296) );
  BUF_X1 U73 ( .A(n8280), .Z(n8297) );
  BUF_X1 U74 ( .A(n8280), .Z(n8298) );
  BUF_X1 U75 ( .A(n8279), .Z(n8302) );
  BUF_X1 U76 ( .A(n8279), .Z(n8303) );
  BUF_X1 U77 ( .A(n8279), .Z(n8304) );
  BUF_X1 U78 ( .A(n8278), .Z(n8308) );
  BUF_X1 U79 ( .A(n8278), .Z(n8309) );
  BUF_X1 U80 ( .A(n8278), .Z(n8310) );
  BUF_X1 U81 ( .A(n8277), .Z(n8314) );
  BUF_X1 U82 ( .A(n8277), .Z(n8315) );
  BUF_X1 U83 ( .A(n8277), .Z(n8316) );
  BUF_X1 U84 ( .A(n8276), .Z(n8320) );
  BUF_X1 U85 ( .A(n8276), .Z(n8321) );
  BUF_X1 U86 ( .A(n8276), .Z(n8322) );
  BUF_X1 U87 ( .A(n8275), .Z(n8326) );
  BUF_X1 U88 ( .A(n8275), .Z(n8327) );
  BUF_X1 U89 ( .A(n8275), .Z(n8328) );
  BUF_X1 U90 ( .A(n8274), .Z(n8332) );
  BUF_X1 U91 ( .A(n8274), .Z(n8333) );
  BUF_X1 U92 ( .A(n8274), .Z(n8334) );
  BUF_X1 U93 ( .A(n8273), .Z(n8338) );
  BUF_X1 U94 ( .A(n8273), .Z(n8339) );
  BUF_X1 U95 ( .A(n8273), .Z(n8340) );
  BUF_X1 U96 ( .A(n8272), .Z(n8344) );
  BUF_X1 U97 ( .A(n8272), .Z(n8345) );
  BUF_X1 U98 ( .A(n8272), .Z(n8346) );
  BUF_X1 U99 ( .A(n8271), .Z(n8350) );
  BUF_X1 U100 ( .A(n8271), .Z(n8351) );
  BUF_X1 U101 ( .A(n8271), .Z(n8352) );
  BUF_X1 U102 ( .A(n8517), .Z(n8407) );
  BUF_X1 U103 ( .A(n8518), .Z(n8408) );
  BUF_X1 U104 ( .A(n8385), .Z(n8411) );
  BUF_X1 U105 ( .A(n8385), .Z(n8412) );
  BUF_X1 U106 ( .A(n8385), .Z(n8413) );
  BUF_X1 U107 ( .A(n8384), .Z(n8417) );
  BUF_X1 U108 ( .A(n8384), .Z(n8418) );
  BUF_X1 U109 ( .A(n8384), .Z(n8419) );
  BUF_X1 U110 ( .A(n8383), .Z(n8423) );
  BUF_X1 U111 ( .A(n8383), .Z(n8424) );
  BUF_X1 U112 ( .A(n8383), .Z(n8425) );
  BUF_X1 U113 ( .A(n8382), .Z(n8429) );
  BUF_X1 U114 ( .A(n8382), .Z(n8430) );
  BUF_X1 U115 ( .A(n8382), .Z(n8431) );
  BUF_X1 U116 ( .A(n8381), .Z(n8435) );
  BUF_X1 U117 ( .A(n8381), .Z(n8436) );
  BUF_X1 U118 ( .A(n8381), .Z(n8437) );
  BUF_X1 U119 ( .A(n8380), .Z(n8441) );
  BUF_X1 U120 ( .A(n8380), .Z(n8442) );
  BUF_X1 U121 ( .A(n8380), .Z(n8443) );
  BUF_X1 U122 ( .A(n8379), .Z(n8447) );
  BUF_X1 U123 ( .A(n8379), .Z(n8448) );
  BUF_X1 U124 ( .A(n8379), .Z(n8449) );
  BUF_X1 U125 ( .A(n8378), .Z(n8453) );
  BUF_X1 U126 ( .A(n8378), .Z(n8454) );
  BUF_X1 U127 ( .A(n8378), .Z(n8455) );
  BUF_X1 U128 ( .A(n8377), .Z(n8459) );
  BUF_X1 U129 ( .A(n8377), .Z(n8460) );
  BUF_X1 U130 ( .A(n8377), .Z(n8461) );
  BUF_X1 U131 ( .A(n8376), .Z(n8465) );
  BUF_X1 U132 ( .A(n8376), .Z(n8466) );
  BUF_X1 U133 ( .A(n8376), .Z(n8467) );
  BUF_X1 U134 ( .A(n8375), .Z(n8471) );
  BUF_X1 U135 ( .A(n8375), .Z(n8472) );
  BUF_X1 U136 ( .A(n8375), .Z(n8473) );
  BUF_X1 U137 ( .A(n8374), .Z(n8477) );
  BUF_X1 U138 ( .A(n8374), .Z(n8478) );
  BUF_X1 U139 ( .A(n8374), .Z(n8479) );
  BUF_X1 U140 ( .A(n8373), .Z(n8483) );
  BUF_X1 U141 ( .A(n8373), .Z(n8484) );
  BUF_X1 U142 ( .A(n8373), .Z(n8485) );
  BUF_X1 U143 ( .A(n8372), .Z(n8489) );
  BUF_X1 U144 ( .A(n8372), .Z(n8490) );
  BUF_X1 U145 ( .A(n8372), .Z(n8491) );
  BUF_X1 U146 ( .A(n8371), .Z(n8495) );
  BUF_X1 U147 ( .A(n8371), .Z(n8496) );
  BUF_X1 U148 ( .A(n8371), .Z(n8497) );
  BUF_X1 U149 ( .A(n8370), .Z(n8501) );
  BUF_X1 U150 ( .A(n8370), .Z(n8502) );
  BUF_X1 U151 ( .A(n8370), .Z(n8503) );
  BUF_X1 U152 ( .A(n8369), .Z(n8507) );
  BUF_X1 U153 ( .A(n8369), .Z(n8508) );
  BUF_X1 U154 ( .A(n8369), .Z(n8509) );
  BUF_X1 U155 ( .A(n8368), .Z(n8513) );
  BUF_X1 U156 ( .A(n8368), .Z(n8514) );
  BUF_X1 U157 ( .A(n8368), .Z(n8515) );
  BUF_X1 U158 ( .A(n8367), .Z(n8519) );
  BUF_X1 U159 ( .A(n8367), .Z(n8520) );
  BUF_X1 U160 ( .A(n8367), .Z(n8521) );
  BUF_X1 U161 ( .A(n8366), .Z(n8525) );
  BUF_X1 U162 ( .A(n8366), .Z(n8526) );
  BUF_X1 U163 ( .A(n8366), .Z(n8527) );
  BUF_X1 U164 ( .A(n8365), .Z(n8531) );
  BUF_X1 U165 ( .A(n8365), .Z(n8532) );
  BUF_X1 U166 ( .A(n8365), .Z(n8533) );
  BUF_X1 U167 ( .A(n8282), .Z(n8284) );
  BUF_X1 U168 ( .A(n8282), .Z(n8285) );
  BUF_X1 U169 ( .A(n8282), .Z(n8286) );
  BUF_X1 U170 ( .A(n8281), .Z(n8287) );
  BUF_X1 U171 ( .A(n8281), .Z(n8288) );
  BUF_X1 U172 ( .A(n8281), .Z(n8289) );
  BUF_X1 U173 ( .A(n8280), .Z(n8293) );
  BUF_X1 U174 ( .A(n8280), .Z(n8294) );
  BUF_X1 U175 ( .A(n8280), .Z(n8295) );
  BUF_X1 U176 ( .A(n8279), .Z(n8299) );
  BUF_X1 U177 ( .A(n8279), .Z(n8300) );
  BUF_X1 U178 ( .A(n8279), .Z(n8301) );
  BUF_X1 U179 ( .A(n8278), .Z(n8305) );
  BUF_X1 U180 ( .A(n8278), .Z(n8306) );
  BUF_X1 U181 ( .A(n8278), .Z(n8307) );
  BUF_X1 U182 ( .A(n8277), .Z(n8311) );
  BUF_X1 U183 ( .A(n8277), .Z(n8312) );
  BUF_X1 U184 ( .A(n8277), .Z(n8313) );
  BUF_X1 U185 ( .A(n8276), .Z(n8317) );
  BUF_X1 U186 ( .A(n8276), .Z(n8318) );
  BUF_X1 U187 ( .A(n8276), .Z(n8319) );
  BUF_X1 U188 ( .A(n8275), .Z(n8323) );
  BUF_X1 U189 ( .A(n8275), .Z(n8324) );
  BUF_X1 U190 ( .A(n8275), .Z(n8325) );
  BUF_X1 U191 ( .A(n8274), .Z(n8329) );
  BUF_X1 U192 ( .A(n8274), .Z(n8330) );
  BUF_X1 U193 ( .A(n8274), .Z(n8331) );
  BUF_X1 U194 ( .A(n8273), .Z(n8335) );
  BUF_X1 U195 ( .A(n8273), .Z(n8336) );
  BUF_X1 U196 ( .A(n8273), .Z(n8337) );
  BUF_X1 U197 ( .A(n8272), .Z(n8341) );
  BUF_X1 U198 ( .A(n8272), .Z(n8342) );
  BUF_X1 U199 ( .A(n8272), .Z(n8343) );
  BUF_X1 U200 ( .A(n8271), .Z(n8347) );
  BUF_X1 U201 ( .A(n8271), .Z(n8348) );
  BUF_X1 U202 ( .A(n8271), .Z(n8349) );
  BUF_X1 U203 ( .A(n8270), .Z(n8353) );
  BUF_X1 U204 ( .A(n8270), .Z(n8354) );
  BUF_X1 U205 ( .A(n8270), .Z(n8355) );
  INV_X1 U206 ( .A(n9224), .ZN(n27130) );
  INV_X1 U207 ( .A(n9235), .ZN(n27129) );
  INV_X1 U208 ( .A(n9245), .ZN(n27128) );
  INV_X1 U209 ( .A(n9255), .ZN(n27127) );
  INV_X1 U210 ( .A(n9265), .ZN(n27126) );
  INV_X1 U211 ( .A(n9275), .ZN(n27125) );
  INV_X1 U212 ( .A(n9285), .ZN(n27124) );
  INV_X1 U213 ( .A(n9295), .ZN(n27123) );
  INV_X1 U214 ( .A(n9305), .ZN(n27122) );
  INV_X1 U215 ( .A(n9315), .ZN(n27121) );
  INV_X1 U216 ( .A(n9325), .ZN(n27120) );
  INV_X1 U217 ( .A(n9335), .ZN(n27119) );
  INV_X1 U218 ( .A(n9345), .ZN(n27118) );
  INV_X1 U219 ( .A(n9355), .ZN(n27117) );
  INV_X1 U220 ( .A(n9365), .ZN(n27116) );
  INV_X1 U221 ( .A(n9375), .ZN(n27115) );
  INV_X1 U222 ( .A(n9385), .ZN(n27114) );
  INV_X1 U223 ( .A(n9395), .ZN(n27113) );
  INV_X1 U224 ( .A(n9405), .ZN(n27112) );
  INV_X1 U225 ( .A(n9415), .ZN(n27111) );
  INV_X1 U226 ( .A(n9425), .ZN(n27110) );
  INV_X1 U227 ( .A(n9435), .ZN(n27109) );
  INV_X1 U228 ( .A(n9445), .ZN(n27108) );
  INV_X1 U229 ( .A(n9455), .ZN(n27107) );
  INV_X1 U230 ( .A(n9465), .ZN(n27106) );
  INV_X1 U231 ( .A(n9475), .ZN(n27105) );
  INV_X1 U232 ( .A(n9485), .ZN(n27104) );
  INV_X1 U233 ( .A(n9495), .ZN(n27103) );
  INV_X1 U234 ( .A(n9505), .ZN(n27102) );
  INV_X1 U235 ( .A(n9515), .ZN(n27101) );
  INV_X1 U236 ( .A(n9525), .ZN(n27100) );
  INV_X1 U237 ( .A(n9535), .ZN(n27099) );
  INV_X1 U238 ( .A(n9621), .ZN(n27090) );
  INV_X1 U239 ( .A(n9630), .ZN(n27089) );
  INV_X1 U240 ( .A(n9639), .ZN(n27088) );
  INV_X1 U241 ( .A(n9648), .ZN(n27087) );
  INV_X1 U242 ( .A(n9657), .ZN(n27086) );
  INV_X1 U243 ( .A(n9666), .ZN(n27085) );
  INV_X1 U244 ( .A(n9675), .ZN(n27084) );
  INV_X1 U245 ( .A(n9684), .ZN(n27083) );
  INV_X1 U246 ( .A(n9693), .ZN(n27082) );
  INV_X1 U247 ( .A(n9702), .ZN(n27081) );
  INV_X1 U248 ( .A(n9711), .ZN(n27080) );
  INV_X1 U249 ( .A(n9720), .ZN(n27079) );
  INV_X1 U250 ( .A(n9729), .ZN(n27078) );
  INV_X1 U251 ( .A(n9738), .ZN(n27077) );
  INV_X1 U252 ( .A(n9747), .ZN(n27076) );
  INV_X1 U253 ( .A(n9756), .ZN(n27075) );
  INV_X1 U254 ( .A(n9765), .ZN(n27074) );
  INV_X1 U255 ( .A(n9774), .ZN(n27073) );
  INV_X1 U256 ( .A(n9783), .ZN(n27072) );
  INV_X1 U257 ( .A(n9792), .ZN(n27071) );
  INV_X1 U258 ( .A(n9801), .ZN(n27070) );
  INV_X1 U259 ( .A(n9810), .ZN(n27069) );
  INV_X1 U260 ( .A(n9819), .ZN(n27068) );
  INV_X1 U261 ( .A(n9828), .ZN(n27067) );
  INV_X1 U262 ( .A(n9911), .ZN(n27058) );
  INV_X1 U263 ( .A(n9920), .ZN(n27057) );
  INV_X1 U264 ( .A(n9929), .ZN(n27056) );
  INV_X1 U265 ( .A(n9938), .ZN(n27055) );
  INV_X1 U266 ( .A(n9947), .ZN(n27054) );
  INV_X1 U267 ( .A(n9956), .ZN(n27053) );
  INV_X1 U268 ( .A(n9965), .ZN(n27052) );
  INV_X1 U269 ( .A(n9974), .ZN(n27051) );
  INV_X1 U270 ( .A(n9983), .ZN(n27050) );
  INV_X1 U271 ( .A(n9992), .ZN(n27049) );
  INV_X1 U272 ( .A(n10001), .ZN(n27048) );
  INV_X1 U273 ( .A(n10010), .ZN(n27047) );
  INV_X1 U274 ( .A(n10019), .ZN(n27046) );
  INV_X1 U275 ( .A(n10028), .ZN(n27045) );
  INV_X1 U276 ( .A(n10037), .ZN(n27044) );
  INV_X1 U277 ( .A(n10046), .ZN(n27043) );
  INV_X1 U278 ( .A(n10055), .ZN(n27042) );
  INV_X1 U279 ( .A(n10064), .ZN(n27041) );
  INV_X1 U280 ( .A(n10073), .ZN(n27040) );
  INV_X1 U281 ( .A(n10082), .ZN(n27039) );
  INV_X1 U282 ( .A(n10091), .ZN(n27038) );
  INV_X1 U283 ( .A(n10100), .ZN(n27037) );
  INV_X1 U284 ( .A(n10109), .ZN(n27036) );
  INV_X1 U285 ( .A(n10118), .ZN(n27035) );
  INV_X1 U286 ( .A(n10201), .ZN(n27026) );
  INV_X1 U287 ( .A(n10210), .ZN(n27025) );
  INV_X1 U288 ( .A(n10219), .ZN(n27024) );
  INV_X1 U289 ( .A(n10228), .ZN(n27023) );
  INV_X1 U290 ( .A(n10237), .ZN(n27022) );
  INV_X1 U291 ( .A(n10246), .ZN(n27021) );
  INV_X1 U292 ( .A(n10255), .ZN(n27020) );
  INV_X1 U293 ( .A(n10264), .ZN(n27019) );
  INV_X1 U294 ( .A(n10273), .ZN(n27018) );
  INV_X1 U295 ( .A(n10282), .ZN(n27017) );
  INV_X1 U296 ( .A(n10291), .ZN(n27016) );
  INV_X1 U297 ( .A(n10300), .ZN(n27015) );
  INV_X1 U298 ( .A(n10309), .ZN(n27014) );
  INV_X1 U299 ( .A(n10318), .ZN(n27013) );
  INV_X1 U300 ( .A(n10327), .ZN(n27012) );
  INV_X1 U301 ( .A(n10336), .ZN(n27011) );
  INV_X1 U302 ( .A(n10345), .ZN(n27010) );
  INV_X1 U303 ( .A(n10354), .ZN(n27009) );
  INV_X1 U304 ( .A(n10363), .ZN(n27008) );
  INV_X1 U305 ( .A(n10372), .ZN(n27007) );
  INV_X1 U306 ( .A(n10381), .ZN(n27006) );
  INV_X1 U307 ( .A(n10390), .ZN(n27005) );
  INV_X1 U308 ( .A(n10399), .ZN(n27004) );
  INV_X1 U309 ( .A(n10408), .ZN(n27003) );
  INV_X1 U310 ( .A(n10491), .ZN(n26994) );
  INV_X1 U311 ( .A(n10500), .ZN(n26993) );
  INV_X1 U312 ( .A(n10509), .ZN(n26992) );
  INV_X1 U313 ( .A(n10518), .ZN(n26991) );
  INV_X1 U314 ( .A(n10527), .ZN(n26990) );
  INV_X1 U315 ( .A(n10536), .ZN(n26989) );
  INV_X1 U316 ( .A(n10545), .ZN(n26988) );
  INV_X1 U317 ( .A(n10554), .ZN(n26987) );
  INV_X1 U318 ( .A(n10563), .ZN(n26986) );
  INV_X1 U319 ( .A(n10572), .ZN(n26985) );
  INV_X1 U320 ( .A(n10581), .ZN(n26984) );
  INV_X1 U321 ( .A(n10590), .ZN(n26983) );
  INV_X1 U322 ( .A(n10599), .ZN(n26982) );
  INV_X1 U323 ( .A(n10608), .ZN(n26981) );
  INV_X1 U324 ( .A(n10617), .ZN(n26980) );
  INV_X1 U325 ( .A(n10626), .ZN(n26979) );
  INV_X1 U326 ( .A(n10635), .ZN(n26978) );
  INV_X1 U327 ( .A(n10644), .ZN(n26977) );
  INV_X1 U328 ( .A(n10653), .ZN(n26976) );
  INV_X1 U329 ( .A(n10662), .ZN(n26975) );
  INV_X1 U330 ( .A(n10671), .ZN(n26974) );
  INV_X1 U331 ( .A(n10680), .ZN(n26973) );
  INV_X1 U332 ( .A(n10689), .ZN(n26972) );
  INV_X1 U333 ( .A(n10698), .ZN(n26971) );
  INV_X1 U334 ( .A(n10781), .ZN(n26962) );
  INV_X1 U335 ( .A(n10790), .ZN(n26961) );
  INV_X1 U336 ( .A(n10799), .ZN(n26960) );
  INV_X1 U337 ( .A(n10808), .ZN(n26959) );
  INV_X1 U338 ( .A(n10817), .ZN(n26958) );
  INV_X1 U339 ( .A(n10826), .ZN(n26957) );
  INV_X1 U340 ( .A(n10835), .ZN(n26956) );
  INV_X1 U341 ( .A(n10844), .ZN(n26955) );
  INV_X1 U342 ( .A(n10853), .ZN(n26954) );
  INV_X1 U343 ( .A(n10862), .ZN(n26953) );
  INV_X1 U344 ( .A(n10871), .ZN(n26952) );
  INV_X1 U345 ( .A(n10880), .ZN(n26951) );
  INV_X1 U346 ( .A(n10889), .ZN(n26950) );
  INV_X1 U347 ( .A(n10898), .ZN(n26949) );
  INV_X1 U348 ( .A(n10907), .ZN(n26948) );
  INV_X1 U349 ( .A(n10916), .ZN(n26947) );
  INV_X1 U350 ( .A(n10925), .ZN(n26946) );
  INV_X1 U351 ( .A(n10934), .ZN(n26945) );
  INV_X1 U352 ( .A(n10943), .ZN(n26944) );
  INV_X1 U353 ( .A(n10952), .ZN(n26943) );
  INV_X1 U354 ( .A(n10961), .ZN(n26942) );
  INV_X1 U355 ( .A(n10970), .ZN(n26941) );
  INV_X1 U356 ( .A(n10979), .ZN(n26940) );
  INV_X1 U357 ( .A(n10988), .ZN(n26939) );
  INV_X1 U358 ( .A(n11071), .ZN(n26930) );
  INV_X1 U359 ( .A(n11080), .ZN(n26929) );
  INV_X1 U360 ( .A(n11089), .ZN(n26928) );
  INV_X1 U361 ( .A(n11098), .ZN(n26927) );
  INV_X1 U362 ( .A(n11107), .ZN(n26926) );
  INV_X1 U363 ( .A(n11116), .ZN(n26925) );
  INV_X1 U364 ( .A(n11125), .ZN(n26924) );
  INV_X1 U365 ( .A(n11134), .ZN(n26923) );
  INV_X1 U366 ( .A(n11143), .ZN(n26922) );
  INV_X1 U367 ( .A(n11152), .ZN(n26921) );
  INV_X1 U368 ( .A(n11161), .ZN(n26920) );
  INV_X1 U369 ( .A(n11170), .ZN(n26919) );
  INV_X1 U370 ( .A(n11179), .ZN(n26918) );
  INV_X1 U371 ( .A(n11188), .ZN(n26917) );
  INV_X1 U372 ( .A(n11197), .ZN(n26916) );
  INV_X1 U373 ( .A(n11206), .ZN(n26915) );
  INV_X1 U374 ( .A(n11215), .ZN(n26914) );
  INV_X1 U375 ( .A(n11224), .ZN(n26913) );
  INV_X1 U376 ( .A(n11233), .ZN(n26912) );
  INV_X1 U377 ( .A(n11242), .ZN(n26911) );
  INV_X1 U378 ( .A(n11251), .ZN(n26910) );
  INV_X1 U379 ( .A(n11260), .ZN(n26909) );
  INV_X1 U380 ( .A(n11269), .ZN(n26908) );
  INV_X1 U381 ( .A(n11278), .ZN(n26907) );
  INV_X1 U382 ( .A(n11361), .ZN(n26898) );
  INV_X1 U383 ( .A(n11370), .ZN(n26897) );
  INV_X1 U384 ( .A(n11379), .ZN(n26896) );
  INV_X1 U385 ( .A(n11388), .ZN(n26895) );
  INV_X1 U386 ( .A(n11397), .ZN(n26894) );
  INV_X1 U387 ( .A(n11406), .ZN(n26893) );
  INV_X1 U388 ( .A(n11415), .ZN(n26892) );
  INV_X1 U389 ( .A(n11424), .ZN(n26891) );
  INV_X1 U390 ( .A(n11433), .ZN(n26890) );
  INV_X1 U391 ( .A(n11442), .ZN(n26889) );
  INV_X1 U392 ( .A(n11451), .ZN(n26888) );
  INV_X1 U393 ( .A(n11460), .ZN(n26887) );
  INV_X1 U394 ( .A(n11469), .ZN(n26886) );
  INV_X1 U395 ( .A(n11478), .ZN(n26885) );
  INV_X1 U396 ( .A(n11487), .ZN(n26884) );
  INV_X1 U397 ( .A(n11496), .ZN(n26883) );
  INV_X1 U398 ( .A(n11505), .ZN(n26882) );
  INV_X1 U399 ( .A(n11514), .ZN(n26881) );
  INV_X1 U400 ( .A(n11523), .ZN(n26880) );
  INV_X1 U401 ( .A(n11532), .ZN(n26879) );
  INV_X1 U402 ( .A(n11541), .ZN(n26878) );
  INV_X1 U403 ( .A(n11550), .ZN(n26877) );
  INV_X1 U404 ( .A(n11559), .ZN(n26876) );
  INV_X1 U405 ( .A(n11568), .ZN(n26875) );
  INV_X1 U406 ( .A(n11651), .ZN(n26866) );
  INV_X1 U407 ( .A(n11660), .ZN(n26865) );
  INV_X1 U408 ( .A(n11669), .ZN(n26864) );
  INV_X1 U409 ( .A(n11678), .ZN(n26863) );
  INV_X1 U410 ( .A(n11687), .ZN(n26862) );
  INV_X1 U411 ( .A(n11696), .ZN(n26861) );
  INV_X1 U412 ( .A(n11705), .ZN(n26860) );
  INV_X1 U413 ( .A(n11714), .ZN(n26859) );
  INV_X1 U414 ( .A(n11723), .ZN(n26858) );
  INV_X1 U415 ( .A(n11732), .ZN(n26857) );
  INV_X1 U416 ( .A(n11741), .ZN(n26856) );
  INV_X1 U417 ( .A(n11750), .ZN(n26855) );
  INV_X1 U418 ( .A(n11759), .ZN(n26854) );
  INV_X1 U419 ( .A(n11768), .ZN(n26853) );
  INV_X1 U420 ( .A(n11777), .ZN(n26852) );
  INV_X1 U421 ( .A(n11786), .ZN(n26851) );
  INV_X1 U422 ( .A(n11795), .ZN(n26850) );
  INV_X1 U423 ( .A(n11804), .ZN(n26849) );
  INV_X1 U424 ( .A(n11813), .ZN(n26848) );
  INV_X1 U425 ( .A(n11822), .ZN(n26847) );
  INV_X1 U426 ( .A(n11831), .ZN(n26846) );
  INV_X1 U427 ( .A(n11840), .ZN(n26845) );
  INV_X1 U428 ( .A(n11849), .ZN(n26844) );
  INV_X1 U429 ( .A(n11858), .ZN(n26843) );
  INV_X1 U430 ( .A(n11941), .ZN(n26834) );
  INV_X1 U431 ( .A(n11950), .ZN(n26833) );
  INV_X1 U432 ( .A(n11959), .ZN(n26832) );
  INV_X1 U433 ( .A(n11968), .ZN(n26831) );
  INV_X1 U434 ( .A(n11977), .ZN(n26830) );
  INV_X1 U435 ( .A(n11986), .ZN(n26829) );
  INV_X1 U436 ( .A(n11995), .ZN(n26828) );
  INV_X1 U437 ( .A(n12004), .ZN(n26827) );
  INV_X1 U438 ( .A(n12013), .ZN(n26826) );
  INV_X1 U439 ( .A(n12022), .ZN(n26825) );
  INV_X1 U440 ( .A(n12031), .ZN(n26824) );
  INV_X1 U441 ( .A(n12040), .ZN(n26823) );
  INV_X1 U442 ( .A(n12049), .ZN(n26822) );
  INV_X1 U443 ( .A(n12058), .ZN(n26821) );
  INV_X1 U444 ( .A(n12067), .ZN(n26820) );
  INV_X1 U445 ( .A(n12076), .ZN(n26819) );
  INV_X1 U446 ( .A(n12085), .ZN(n26818) );
  INV_X1 U447 ( .A(n12094), .ZN(n26817) );
  INV_X1 U448 ( .A(n12103), .ZN(n26816) );
  INV_X1 U449 ( .A(n12112), .ZN(n26815) );
  INV_X1 U450 ( .A(n12121), .ZN(n26814) );
  INV_X1 U451 ( .A(n12130), .ZN(n26813) );
  INV_X1 U452 ( .A(n12139), .ZN(n26812) );
  INV_X1 U453 ( .A(n12148), .ZN(n26811) );
  INV_X1 U454 ( .A(n12230), .ZN(n26802) );
  INV_X1 U455 ( .A(n12239), .ZN(n26801) );
  INV_X1 U456 ( .A(n12248), .ZN(n26800) );
  INV_X1 U457 ( .A(n12257), .ZN(n26799) );
  INV_X1 U458 ( .A(n12266), .ZN(n26798) );
  INV_X1 U459 ( .A(n12275), .ZN(n26797) );
  INV_X1 U460 ( .A(n12284), .ZN(n26796) );
  INV_X1 U461 ( .A(n12293), .ZN(n26795) );
  INV_X1 U462 ( .A(n12302), .ZN(n26794) );
  INV_X1 U463 ( .A(n12311), .ZN(n26793) );
  INV_X1 U464 ( .A(n12320), .ZN(n26792) );
  INV_X1 U465 ( .A(n12329), .ZN(n26791) );
  INV_X1 U466 ( .A(n12338), .ZN(n26790) );
  INV_X1 U467 ( .A(n12347), .ZN(n26789) );
  INV_X1 U468 ( .A(n12356), .ZN(n26788) );
  INV_X1 U469 ( .A(n12365), .ZN(n26787) );
  INV_X1 U470 ( .A(n12374), .ZN(n26786) );
  INV_X1 U471 ( .A(n12383), .ZN(n26785) );
  INV_X1 U472 ( .A(n12392), .ZN(n26784) );
  INV_X1 U473 ( .A(n12401), .ZN(n26783) );
  INV_X1 U474 ( .A(n12410), .ZN(n26782) );
  INV_X1 U475 ( .A(n12419), .ZN(n26781) );
  INV_X1 U476 ( .A(n12428), .ZN(n26780) );
  INV_X1 U477 ( .A(n12437), .ZN(n26779) );
  INV_X1 U478 ( .A(n12519), .ZN(n26770) );
  INV_X1 U479 ( .A(n12528), .ZN(n26769) );
  INV_X1 U480 ( .A(n12537), .ZN(n26768) );
  INV_X1 U481 ( .A(n12546), .ZN(n26767) );
  INV_X1 U482 ( .A(n12555), .ZN(n26766) );
  INV_X1 U483 ( .A(n12564), .ZN(n26765) );
  INV_X1 U484 ( .A(n12573), .ZN(n26764) );
  INV_X1 U485 ( .A(n12582), .ZN(n26763) );
  INV_X1 U486 ( .A(n12591), .ZN(n26762) );
  INV_X1 U487 ( .A(n12600), .ZN(n26761) );
  INV_X1 U488 ( .A(n12609), .ZN(n26760) );
  INV_X1 U489 ( .A(n12618), .ZN(n26759) );
  INV_X1 U490 ( .A(n12627), .ZN(n26758) );
  INV_X1 U491 ( .A(n12636), .ZN(n26757) );
  INV_X1 U492 ( .A(n12645), .ZN(n26756) );
  INV_X1 U493 ( .A(n12654), .ZN(n26755) );
  INV_X1 U494 ( .A(n12663), .ZN(n26754) );
  INV_X1 U495 ( .A(n12672), .ZN(n26753) );
  INV_X1 U496 ( .A(n12681), .ZN(n26752) );
  INV_X1 U497 ( .A(n12690), .ZN(n26751) );
  INV_X1 U498 ( .A(n12699), .ZN(n26750) );
  INV_X1 U499 ( .A(n12708), .ZN(n26749) );
  INV_X1 U500 ( .A(n12717), .ZN(n26748) );
  INV_X1 U501 ( .A(n12726), .ZN(n26747) );
  INV_X1 U502 ( .A(n12808), .ZN(n26738) );
  INV_X1 U503 ( .A(n12817), .ZN(n26737) );
  INV_X1 U504 ( .A(n12826), .ZN(n26736) );
  INV_X1 U505 ( .A(n12835), .ZN(n26735) );
  INV_X1 U506 ( .A(n12844), .ZN(n26734) );
  INV_X1 U507 ( .A(n12853), .ZN(n26733) );
  INV_X1 U508 ( .A(n12862), .ZN(n26732) );
  INV_X1 U509 ( .A(n12871), .ZN(n26731) );
  INV_X1 U510 ( .A(n12880), .ZN(n26730) );
  INV_X1 U511 ( .A(n12889), .ZN(n26729) );
  INV_X1 U512 ( .A(n12898), .ZN(n26728) );
  INV_X1 U513 ( .A(n12907), .ZN(n26727) );
  INV_X1 U514 ( .A(n12916), .ZN(n26726) );
  INV_X1 U515 ( .A(n12925), .ZN(n26725) );
  INV_X1 U516 ( .A(n12934), .ZN(n26724) );
  INV_X1 U517 ( .A(n12943), .ZN(n26723) );
  INV_X1 U518 ( .A(n12952), .ZN(n26722) );
  INV_X1 U519 ( .A(n12961), .ZN(n26721) );
  INV_X1 U520 ( .A(n12970), .ZN(n26720) );
  INV_X1 U521 ( .A(n12979), .ZN(n26719) );
  INV_X1 U522 ( .A(n12988), .ZN(n26718) );
  INV_X1 U523 ( .A(n12997), .ZN(n26717) );
  INV_X1 U524 ( .A(n13006), .ZN(n26716) );
  INV_X1 U525 ( .A(n13015), .ZN(n26715) );
  INV_X1 U526 ( .A(n13097), .ZN(n26706) );
  INV_X1 U527 ( .A(n13106), .ZN(n26705) );
  INV_X1 U528 ( .A(n13115), .ZN(n26704) );
  INV_X1 U529 ( .A(n13124), .ZN(n26703) );
  INV_X1 U530 ( .A(n13133), .ZN(n26702) );
  INV_X1 U531 ( .A(n13142), .ZN(n26701) );
  INV_X1 U532 ( .A(n13151), .ZN(n26700) );
  INV_X1 U533 ( .A(n13160), .ZN(n26699) );
  INV_X1 U534 ( .A(n13169), .ZN(n26698) );
  INV_X1 U535 ( .A(n13178), .ZN(n26697) );
  INV_X1 U536 ( .A(n13187), .ZN(n26696) );
  INV_X1 U537 ( .A(n13196), .ZN(n26695) );
  INV_X1 U538 ( .A(n13205), .ZN(n26694) );
  INV_X1 U539 ( .A(n13214), .ZN(n26693) );
  INV_X1 U540 ( .A(n13223), .ZN(n26692) );
  INV_X1 U541 ( .A(n13232), .ZN(n26691) );
  INV_X1 U542 ( .A(n13241), .ZN(n26690) );
  INV_X1 U543 ( .A(n13250), .ZN(n26689) );
  INV_X1 U544 ( .A(n13259), .ZN(n26688) );
  INV_X1 U545 ( .A(n13268), .ZN(n26687) );
  INV_X1 U546 ( .A(n13277), .ZN(n26686) );
  INV_X1 U547 ( .A(n13286), .ZN(n26685) );
  INV_X1 U548 ( .A(n13295), .ZN(n26684) );
  INV_X1 U549 ( .A(n13304), .ZN(n26683) );
  INV_X1 U550 ( .A(n13386), .ZN(n26674) );
  INV_X1 U551 ( .A(n13395), .ZN(n26673) );
  INV_X1 U552 ( .A(n13404), .ZN(n26672) );
  INV_X1 U553 ( .A(n13413), .ZN(n26671) );
  INV_X1 U554 ( .A(n13422), .ZN(n26670) );
  INV_X1 U555 ( .A(n13431), .ZN(n26669) );
  INV_X1 U556 ( .A(n13440), .ZN(n26668) );
  INV_X1 U557 ( .A(n13449), .ZN(n26667) );
  INV_X1 U558 ( .A(n13458), .ZN(n26666) );
  INV_X1 U559 ( .A(n13467), .ZN(n26665) );
  INV_X1 U560 ( .A(n13476), .ZN(n26664) );
  INV_X1 U561 ( .A(n13485), .ZN(n26663) );
  INV_X1 U562 ( .A(n13494), .ZN(n26662) );
  INV_X1 U563 ( .A(n13503), .ZN(n26661) );
  INV_X1 U564 ( .A(n13512), .ZN(n26660) );
  INV_X1 U565 ( .A(n13521), .ZN(n26659) );
  INV_X1 U566 ( .A(n13530), .ZN(n26658) );
  INV_X1 U567 ( .A(n13539), .ZN(n26657) );
  INV_X1 U568 ( .A(n13548), .ZN(n26656) );
  INV_X1 U569 ( .A(n13557), .ZN(n26655) );
  INV_X1 U570 ( .A(n13566), .ZN(n26654) );
  INV_X1 U571 ( .A(n13575), .ZN(n26653) );
  INV_X1 U572 ( .A(n13584), .ZN(n26652) );
  INV_X1 U573 ( .A(n13593), .ZN(n26651) );
  INV_X1 U574 ( .A(n13675), .ZN(n26642) );
  INV_X1 U575 ( .A(n13684), .ZN(n26641) );
  INV_X1 U576 ( .A(n13693), .ZN(n26640) );
  INV_X1 U577 ( .A(n13702), .ZN(n26639) );
  INV_X1 U578 ( .A(n13711), .ZN(n26638) );
  INV_X1 U579 ( .A(n13720), .ZN(n26637) );
  INV_X1 U580 ( .A(n13729), .ZN(n26636) );
  INV_X1 U581 ( .A(n13738), .ZN(n26635) );
  INV_X1 U582 ( .A(n13747), .ZN(n26634) );
  INV_X1 U583 ( .A(n13756), .ZN(n26633) );
  INV_X1 U584 ( .A(n13765), .ZN(n26632) );
  INV_X1 U585 ( .A(n13774), .ZN(n26631) );
  INV_X1 U586 ( .A(n13783), .ZN(n26630) );
  INV_X1 U587 ( .A(n13792), .ZN(n26629) );
  INV_X1 U588 ( .A(n13801), .ZN(n26628) );
  INV_X1 U589 ( .A(n13810), .ZN(n26627) );
  INV_X1 U590 ( .A(n13819), .ZN(n26626) );
  INV_X1 U591 ( .A(n13828), .ZN(n26625) );
  INV_X1 U592 ( .A(n13837), .ZN(n26624) );
  INV_X1 U593 ( .A(n13846), .ZN(n26623) );
  INV_X1 U594 ( .A(n13855), .ZN(n26622) );
  INV_X1 U595 ( .A(n13864), .ZN(n26621) );
  INV_X1 U596 ( .A(n13873), .ZN(n26620) );
  INV_X1 U597 ( .A(n13882), .ZN(n26619) );
  INV_X1 U598 ( .A(n13964), .ZN(n26610) );
  INV_X1 U599 ( .A(n13973), .ZN(n26609) );
  INV_X1 U600 ( .A(n13982), .ZN(n26608) );
  INV_X1 U601 ( .A(n13991), .ZN(n26607) );
  INV_X1 U602 ( .A(n14000), .ZN(n26606) );
  INV_X1 U603 ( .A(n14009), .ZN(n26605) );
  INV_X1 U604 ( .A(n14018), .ZN(n26604) );
  INV_X1 U605 ( .A(n14027), .ZN(n26603) );
  INV_X1 U606 ( .A(n14036), .ZN(n26602) );
  INV_X1 U607 ( .A(n14045), .ZN(n26601) );
  INV_X1 U608 ( .A(n14054), .ZN(n26600) );
  INV_X1 U609 ( .A(n14063), .ZN(n26599) );
  INV_X1 U610 ( .A(n14072), .ZN(n26598) );
  INV_X1 U611 ( .A(n14081), .ZN(n26597) );
  INV_X1 U612 ( .A(n14090), .ZN(n26596) );
  INV_X1 U613 ( .A(n14099), .ZN(n26595) );
  INV_X1 U614 ( .A(n14108), .ZN(n26594) );
  INV_X1 U615 ( .A(n14117), .ZN(n26593) );
  INV_X1 U616 ( .A(n14126), .ZN(n26592) );
  INV_X1 U617 ( .A(n14135), .ZN(n26591) );
  INV_X1 U618 ( .A(n14144), .ZN(n26590) );
  INV_X1 U619 ( .A(n14153), .ZN(n26589) );
  INV_X1 U620 ( .A(n14162), .ZN(n26588) );
  INV_X1 U621 ( .A(n14171), .ZN(n26587) );
  INV_X1 U622 ( .A(n14254), .ZN(n26578) );
  INV_X1 U623 ( .A(n14263), .ZN(n26577) );
  INV_X1 U624 ( .A(n14272), .ZN(n26576) );
  INV_X1 U625 ( .A(n14281), .ZN(n26575) );
  INV_X1 U626 ( .A(n14290), .ZN(n26574) );
  INV_X1 U627 ( .A(n14299), .ZN(n26573) );
  INV_X1 U628 ( .A(n14308), .ZN(n26572) );
  INV_X1 U629 ( .A(n14317), .ZN(n26571) );
  INV_X1 U630 ( .A(n14326), .ZN(n26570) );
  INV_X1 U631 ( .A(n14335), .ZN(n26569) );
  INV_X1 U632 ( .A(n14344), .ZN(n26568) );
  INV_X1 U633 ( .A(n14353), .ZN(n26567) );
  INV_X1 U634 ( .A(n14362), .ZN(n26566) );
  INV_X1 U635 ( .A(n14371), .ZN(n26565) );
  INV_X1 U636 ( .A(n14380), .ZN(n26564) );
  INV_X1 U637 ( .A(n14389), .ZN(n26563) );
  INV_X1 U638 ( .A(n14398), .ZN(n26562) );
  INV_X1 U639 ( .A(n14407), .ZN(n26561) );
  INV_X1 U640 ( .A(n14416), .ZN(n26560) );
  INV_X1 U641 ( .A(n14425), .ZN(n26559) );
  INV_X1 U642 ( .A(n14434), .ZN(n26558) );
  INV_X1 U643 ( .A(n14443), .ZN(n26557) );
  INV_X1 U644 ( .A(n14452), .ZN(n26556) );
  INV_X1 U645 ( .A(n14461), .ZN(n26555) );
  INV_X1 U646 ( .A(n14543), .ZN(n26546) );
  INV_X1 U647 ( .A(n14552), .ZN(n26545) );
  INV_X1 U648 ( .A(n14561), .ZN(n26544) );
  INV_X1 U649 ( .A(n14570), .ZN(n26543) );
  INV_X1 U650 ( .A(n14579), .ZN(n26542) );
  INV_X1 U651 ( .A(n14588), .ZN(n26541) );
  INV_X1 U652 ( .A(n14597), .ZN(n26540) );
  INV_X1 U653 ( .A(n14606), .ZN(n26539) );
  INV_X1 U654 ( .A(n14615), .ZN(n26538) );
  INV_X1 U655 ( .A(n14624), .ZN(n26537) );
  INV_X1 U656 ( .A(n14633), .ZN(n26536) );
  INV_X1 U657 ( .A(n14642), .ZN(n26535) );
  INV_X1 U658 ( .A(n14651), .ZN(n26534) );
  INV_X1 U659 ( .A(n14660), .ZN(n26533) );
  INV_X1 U660 ( .A(n14669), .ZN(n26532) );
  INV_X1 U661 ( .A(n14678), .ZN(n26531) );
  INV_X1 U662 ( .A(n14687), .ZN(n26530) );
  INV_X1 U663 ( .A(n14696), .ZN(n26529) );
  INV_X1 U664 ( .A(n14705), .ZN(n26528) );
  INV_X1 U665 ( .A(n14714), .ZN(n26527) );
  INV_X1 U666 ( .A(n14723), .ZN(n26526) );
  INV_X1 U667 ( .A(n14732), .ZN(n26525) );
  INV_X1 U668 ( .A(n14741), .ZN(n26524) );
  INV_X1 U669 ( .A(n14750), .ZN(n26523) );
  INV_X1 U670 ( .A(n14832), .ZN(n26514) );
  INV_X1 U671 ( .A(n14841), .ZN(n26513) );
  INV_X1 U672 ( .A(n14850), .ZN(n26512) );
  INV_X1 U673 ( .A(n14859), .ZN(n26511) );
  INV_X1 U674 ( .A(n14868), .ZN(n26510) );
  INV_X1 U675 ( .A(n14877), .ZN(n26509) );
  INV_X1 U676 ( .A(n14886), .ZN(n26508) );
  INV_X1 U677 ( .A(n14895), .ZN(n26507) );
  INV_X1 U678 ( .A(n14904), .ZN(n26506) );
  INV_X1 U679 ( .A(n14913), .ZN(n26505) );
  INV_X1 U680 ( .A(n14922), .ZN(n26504) );
  INV_X1 U681 ( .A(n14931), .ZN(n26503) );
  INV_X1 U682 ( .A(n14940), .ZN(n26502) );
  INV_X1 U683 ( .A(n14949), .ZN(n26501) );
  INV_X1 U684 ( .A(n14958), .ZN(n26500) );
  INV_X1 U685 ( .A(n14967), .ZN(n26499) );
  INV_X1 U686 ( .A(n14976), .ZN(n26498) );
  INV_X1 U687 ( .A(n14985), .ZN(n26497) );
  INV_X1 U688 ( .A(n14994), .ZN(n26496) );
  INV_X1 U689 ( .A(n15003), .ZN(n26495) );
  INV_X1 U690 ( .A(n15012), .ZN(n26494) );
  INV_X1 U691 ( .A(n15021), .ZN(n26493) );
  INV_X1 U692 ( .A(n15030), .ZN(n26492) );
  INV_X1 U693 ( .A(n15039), .ZN(n26491) );
  INV_X1 U694 ( .A(n15121), .ZN(n26482) );
  INV_X1 U695 ( .A(n15130), .ZN(n26481) );
  INV_X1 U696 ( .A(n15139), .ZN(n26480) );
  INV_X1 U697 ( .A(n15148), .ZN(n26479) );
  INV_X1 U698 ( .A(n15157), .ZN(n26478) );
  INV_X1 U699 ( .A(n15166), .ZN(n26477) );
  INV_X1 U700 ( .A(n15175), .ZN(n26476) );
  INV_X1 U701 ( .A(n15184), .ZN(n26475) );
  INV_X1 U702 ( .A(n15193), .ZN(n26474) );
  INV_X1 U703 ( .A(n15202), .ZN(n26473) );
  INV_X1 U704 ( .A(n15211), .ZN(n26472) );
  INV_X1 U705 ( .A(n15220), .ZN(n26471) );
  INV_X1 U706 ( .A(n15229), .ZN(n26470) );
  INV_X1 U707 ( .A(n15238), .ZN(n26469) );
  INV_X1 U708 ( .A(n15247), .ZN(n26468) );
  INV_X1 U709 ( .A(n15256), .ZN(n26467) );
  INV_X1 U710 ( .A(n15265), .ZN(n26466) );
  INV_X1 U711 ( .A(n15274), .ZN(n26465) );
  INV_X1 U712 ( .A(n15283), .ZN(n26464) );
  INV_X1 U713 ( .A(n15292), .ZN(n26463) );
  INV_X1 U714 ( .A(n15301), .ZN(n26462) );
  INV_X1 U715 ( .A(n15310), .ZN(n26461) );
  INV_X1 U716 ( .A(n15319), .ZN(n26460) );
  INV_X1 U717 ( .A(n15328), .ZN(n26459) );
  INV_X1 U718 ( .A(n15410), .ZN(n26450) );
  INV_X1 U719 ( .A(n15419), .ZN(n26449) );
  INV_X1 U720 ( .A(n15428), .ZN(n26448) );
  INV_X1 U721 ( .A(n15437), .ZN(n26447) );
  INV_X1 U722 ( .A(n15446), .ZN(n26446) );
  INV_X1 U723 ( .A(n15455), .ZN(n26445) );
  INV_X1 U724 ( .A(n15464), .ZN(n26444) );
  INV_X1 U725 ( .A(n15473), .ZN(n26443) );
  INV_X1 U726 ( .A(n15482), .ZN(n26442) );
  INV_X1 U727 ( .A(n15491), .ZN(n26441) );
  INV_X1 U728 ( .A(n15500), .ZN(n26440) );
  INV_X1 U729 ( .A(n15509), .ZN(n26439) );
  INV_X1 U730 ( .A(n15518), .ZN(n26438) );
  INV_X1 U731 ( .A(n15527), .ZN(n26437) );
  INV_X1 U732 ( .A(n15536), .ZN(n26436) );
  INV_X1 U733 ( .A(n15545), .ZN(n26435) );
  INV_X1 U734 ( .A(n15554), .ZN(n26434) );
  INV_X1 U735 ( .A(n15563), .ZN(n26433) );
  INV_X1 U736 ( .A(n15572), .ZN(n26432) );
  INV_X1 U737 ( .A(n15581), .ZN(n26431) );
  INV_X1 U738 ( .A(n15590), .ZN(n26430) );
  INV_X1 U739 ( .A(n15599), .ZN(n26429) );
  INV_X1 U740 ( .A(n15608), .ZN(n26428) );
  INV_X1 U741 ( .A(n15617), .ZN(n26427) );
  INV_X1 U742 ( .A(n15699), .ZN(n26418) );
  INV_X1 U743 ( .A(n15708), .ZN(n26417) );
  INV_X1 U744 ( .A(n15717), .ZN(n26416) );
  INV_X1 U745 ( .A(n15726), .ZN(n26415) );
  INV_X1 U746 ( .A(n15735), .ZN(n26414) );
  INV_X1 U747 ( .A(n15744), .ZN(n26413) );
  INV_X1 U748 ( .A(n15753), .ZN(n26412) );
  INV_X1 U749 ( .A(n15762), .ZN(n26411) );
  INV_X1 U750 ( .A(n15771), .ZN(n26410) );
  INV_X1 U751 ( .A(n15780), .ZN(n26409) );
  INV_X1 U752 ( .A(n15789), .ZN(n26408) );
  INV_X1 U753 ( .A(n15798), .ZN(n26407) );
  INV_X1 U754 ( .A(n15807), .ZN(n26406) );
  INV_X1 U755 ( .A(n15816), .ZN(n26405) );
  INV_X1 U756 ( .A(n15825), .ZN(n26404) );
  INV_X1 U757 ( .A(n15834), .ZN(n26403) );
  INV_X1 U758 ( .A(n15843), .ZN(n26402) );
  INV_X1 U759 ( .A(n15852), .ZN(n26401) );
  INV_X1 U760 ( .A(n15861), .ZN(n26400) );
  INV_X1 U761 ( .A(n15870), .ZN(n26399) );
  INV_X1 U762 ( .A(n15879), .ZN(n26398) );
  INV_X1 U763 ( .A(n15888), .ZN(n26397) );
  INV_X1 U764 ( .A(n15897), .ZN(n26396) );
  INV_X1 U765 ( .A(n15906), .ZN(n26395) );
  INV_X1 U766 ( .A(n15988), .ZN(n26386) );
  INV_X1 U767 ( .A(n15997), .ZN(n26385) );
  INV_X1 U768 ( .A(n16006), .ZN(n26384) );
  INV_X1 U769 ( .A(n16015), .ZN(n26383) );
  INV_X1 U770 ( .A(n16024), .ZN(n26382) );
  INV_X1 U771 ( .A(n16033), .ZN(n26381) );
  INV_X1 U772 ( .A(n16042), .ZN(n26380) );
  INV_X1 U773 ( .A(n16051), .ZN(n26379) );
  INV_X1 U774 ( .A(n16060), .ZN(n26378) );
  INV_X1 U775 ( .A(n16069), .ZN(n26377) );
  INV_X1 U776 ( .A(n16078), .ZN(n26376) );
  INV_X1 U777 ( .A(n16087), .ZN(n26375) );
  INV_X1 U778 ( .A(n16096), .ZN(n26374) );
  INV_X1 U779 ( .A(n16105), .ZN(n26373) );
  INV_X1 U780 ( .A(n16114), .ZN(n26372) );
  INV_X1 U781 ( .A(n16123), .ZN(n26371) );
  INV_X1 U782 ( .A(n16132), .ZN(n26370) );
  INV_X1 U783 ( .A(n16141), .ZN(n26369) );
  INV_X1 U784 ( .A(n16150), .ZN(n26368) );
  INV_X1 U785 ( .A(n16159), .ZN(n26367) );
  INV_X1 U786 ( .A(n16168), .ZN(n26366) );
  INV_X1 U787 ( .A(n16177), .ZN(n26365) );
  INV_X1 U788 ( .A(n16186), .ZN(n26364) );
  INV_X1 U789 ( .A(n16195), .ZN(n26363) );
  INV_X1 U790 ( .A(n16277), .ZN(n26354) );
  INV_X1 U791 ( .A(n16286), .ZN(n26353) );
  INV_X1 U792 ( .A(n16295), .ZN(n26352) );
  INV_X1 U793 ( .A(n16304), .ZN(n26351) );
  INV_X1 U794 ( .A(n16313), .ZN(n26350) );
  INV_X1 U795 ( .A(n16322), .ZN(n26349) );
  INV_X1 U796 ( .A(n16331), .ZN(n26348) );
  INV_X1 U797 ( .A(n16340), .ZN(n26347) );
  INV_X1 U798 ( .A(n16349), .ZN(n26346) );
  INV_X1 U799 ( .A(n16358), .ZN(n26345) );
  INV_X1 U800 ( .A(n16367), .ZN(n26344) );
  INV_X1 U801 ( .A(n16376), .ZN(n26343) );
  INV_X1 U802 ( .A(n16385), .ZN(n26342) );
  INV_X1 U803 ( .A(n16394), .ZN(n26341) );
  INV_X1 U804 ( .A(n16403), .ZN(n26340) );
  INV_X1 U805 ( .A(n16412), .ZN(n26339) );
  INV_X1 U806 ( .A(n16421), .ZN(n26338) );
  INV_X1 U807 ( .A(n16430), .ZN(n26337) );
  INV_X1 U808 ( .A(n16439), .ZN(n26336) );
  INV_X1 U809 ( .A(n16448), .ZN(n26335) );
  INV_X1 U810 ( .A(n16457), .ZN(n26334) );
  INV_X1 U811 ( .A(n16466), .ZN(n26333) );
  INV_X1 U812 ( .A(n16475), .ZN(n26332) );
  INV_X1 U813 ( .A(n16484), .ZN(n26331) );
  INV_X1 U814 ( .A(n16567), .ZN(n26322) );
  INV_X1 U815 ( .A(n16576), .ZN(n26321) );
  INV_X1 U816 ( .A(n16585), .ZN(n26320) );
  INV_X1 U817 ( .A(n16594), .ZN(n26319) );
  INV_X1 U818 ( .A(n16603), .ZN(n26318) );
  INV_X1 U819 ( .A(n16612), .ZN(n26317) );
  INV_X1 U820 ( .A(n16621), .ZN(n26316) );
  INV_X1 U821 ( .A(n16630), .ZN(n26315) );
  INV_X1 U822 ( .A(n16639), .ZN(n26314) );
  INV_X1 U823 ( .A(n16648), .ZN(n26313) );
  INV_X1 U824 ( .A(n16657), .ZN(n26312) );
  INV_X1 U825 ( .A(n16666), .ZN(n26311) );
  INV_X1 U826 ( .A(n16675), .ZN(n26310) );
  INV_X1 U827 ( .A(n16684), .ZN(n26309) );
  INV_X1 U828 ( .A(n16693), .ZN(n26308) );
  INV_X1 U829 ( .A(n16702), .ZN(n26307) );
  INV_X1 U830 ( .A(n16711), .ZN(n26306) );
  INV_X1 U831 ( .A(n16720), .ZN(n26305) );
  INV_X1 U832 ( .A(n16729), .ZN(n26304) );
  INV_X1 U833 ( .A(n16738), .ZN(n26303) );
  INV_X1 U834 ( .A(n16747), .ZN(n26302) );
  INV_X1 U835 ( .A(n16756), .ZN(n26301) );
  INV_X1 U836 ( .A(n16765), .ZN(n26300) );
  INV_X1 U837 ( .A(n16774), .ZN(n26299) );
  INV_X1 U838 ( .A(n16856), .ZN(n26290) );
  INV_X1 U839 ( .A(n16865), .ZN(n26289) );
  INV_X1 U840 ( .A(n16874), .ZN(n26288) );
  INV_X1 U841 ( .A(n16883), .ZN(n26287) );
  INV_X1 U842 ( .A(n16892), .ZN(n26286) );
  INV_X1 U843 ( .A(n16901), .ZN(n26285) );
  INV_X1 U844 ( .A(n16910), .ZN(n26284) );
  INV_X1 U845 ( .A(n16919), .ZN(n26283) );
  INV_X1 U846 ( .A(n16928), .ZN(n26282) );
  INV_X1 U847 ( .A(n16937), .ZN(n26281) );
  INV_X1 U848 ( .A(n16946), .ZN(n26280) );
  INV_X1 U849 ( .A(n16955), .ZN(n26279) );
  INV_X1 U850 ( .A(n16964), .ZN(n26278) );
  INV_X1 U851 ( .A(n16973), .ZN(n26277) );
  INV_X1 U852 ( .A(n16982), .ZN(n26276) );
  INV_X1 U853 ( .A(n16991), .ZN(n26275) );
  INV_X1 U854 ( .A(n17000), .ZN(n26274) );
  INV_X1 U855 ( .A(n17009), .ZN(n26273) );
  INV_X1 U856 ( .A(n17018), .ZN(n26272) );
  INV_X1 U857 ( .A(n17027), .ZN(n26271) );
  INV_X1 U858 ( .A(n17036), .ZN(n26270) );
  INV_X1 U859 ( .A(n17045), .ZN(n26269) );
  INV_X1 U860 ( .A(n17054), .ZN(n26268) );
  INV_X1 U861 ( .A(n17063), .ZN(n26267) );
  INV_X1 U862 ( .A(n17145), .ZN(n26258) );
  INV_X1 U863 ( .A(n17154), .ZN(n26257) );
  INV_X1 U864 ( .A(n17163), .ZN(n26256) );
  INV_X1 U865 ( .A(n17172), .ZN(n26255) );
  INV_X1 U866 ( .A(n17181), .ZN(n26254) );
  INV_X1 U867 ( .A(n17190), .ZN(n26253) );
  INV_X1 U868 ( .A(n17199), .ZN(n26252) );
  INV_X1 U869 ( .A(n17208), .ZN(n26251) );
  INV_X1 U870 ( .A(n17217), .ZN(n26250) );
  INV_X1 U871 ( .A(n17226), .ZN(n26249) );
  INV_X1 U872 ( .A(n17235), .ZN(n26248) );
  INV_X1 U873 ( .A(n17244), .ZN(n26247) );
  INV_X1 U874 ( .A(n17253), .ZN(n26246) );
  INV_X1 U875 ( .A(n17262), .ZN(n26245) );
  INV_X1 U876 ( .A(n17271), .ZN(n26244) );
  INV_X1 U877 ( .A(n17280), .ZN(n26243) );
  INV_X1 U878 ( .A(n17289), .ZN(n26242) );
  INV_X1 U879 ( .A(n17298), .ZN(n26241) );
  INV_X1 U880 ( .A(n17307), .ZN(n26240) );
  INV_X1 U881 ( .A(n17316), .ZN(n26239) );
  INV_X1 U882 ( .A(n17325), .ZN(n26238) );
  INV_X1 U883 ( .A(n17334), .ZN(n26237) );
  INV_X1 U884 ( .A(n17343), .ZN(n26236) );
  INV_X1 U885 ( .A(n17352), .ZN(n26235) );
  INV_X1 U886 ( .A(n17434), .ZN(n26226) );
  INV_X1 U887 ( .A(n17443), .ZN(n26225) );
  INV_X1 U888 ( .A(n17452), .ZN(n26224) );
  INV_X1 U889 ( .A(n17461), .ZN(n26223) );
  INV_X1 U890 ( .A(n17470), .ZN(n26222) );
  INV_X1 U891 ( .A(n17479), .ZN(n26221) );
  INV_X1 U892 ( .A(n17488), .ZN(n26220) );
  INV_X1 U893 ( .A(n17497), .ZN(n26219) );
  INV_X1 U894 ( .A(n17506), .ZN(n26218) );
  INV_X1 U895 ( .A(n17515), .ZN(n26217) );
  INV_X1 U896 ( .A(n17524), .ZN(n26216) );
  INV_X1 U897 ( .A(n17533), .ZN(n26215) );
  INV_X1 U898 ( .A(n17542), .ZN(n26214) );
  INV_X1 U899 ( .A(n17551), .ZN(n26213) );
  INV_X1 U900 ( .A(n17560), .ZN(n26212) );
  INV_X1 U901 ( .A(n17569), .ZN(n26211) );
  INV_X1 U902 ( .A(n17578), .ZN(n26210) );
  INV_X1 U903 ( .A(n17587), .ZN(n26209) );
  INV_X1 U904 ( .A(n17596), .ZN(n26208) );
  INV_X1 U905 ( .A(n17605), .ZN(n26207) );
  INV_X1 U906 ( .A(n17614), .ZN(n26206) );
  INV_X1 U907 ( .A(n17623), .ZN(n26205) );
  INV_X1 U908 ( .A(n17632), .ZN(n26204) );
  INV_X1 U909 ( .A(n17641), .ZN(n26203) );
  INV_X1 U910 ( .A(n17723), .ZN(n26194) );
  INV_X1 U911 ( .A(n17732), .ZN(n26193) );
  INV_X1 U912 ( .A(n17741), .ZN(n26192) );
  INV_X1 U913 ( .A(n17750), .ZN(n26191) );
  INV_X1 U914 ( .A(n17759), .ZN(n26190) );
  INV_X1 U915 ( .A(n17768), .ZN(n26189) );
  INV_X1 U916 ( .A(n17777), .ZN(n26188) );
  INV_X1 U917 ( .A(n17786), .ZN(n26187) );
  INV_X1 U918 ( .A(n17795), .ZN(n26186) );
  INV_X1 U919 ( .A(n17804), .ZN(n26185) );
  INV_X1 U920 ( .A(n17813), .ZN(n26184) );
  INV_X1 U921 ( .A(n17822), .ZN(n26183) );
  INV_X1 U922 ( .A(n17831), .ZN(n26182) );
  INV_X1 U923 ( .A(n17840), .ZN(n26181) );
  INV_X1 U924 ( .A(n17849), .ZN(n26180) );
  INV_X1 U925 ( .A(n17858), .ZN(n26179) );
  INV_X1 U926 ( .A(n17867), .ZN(n26178) );
  INV_X1 U927 ( .A(n17876), .ZN(n26177) );
  INV_X1 U928 ( .A(n17885), .ZN(n26176) );
  INV_X1 U929 ( .A(n17894), .ZN(n26175) );
  INV_X1 U930 ( .A(n17903), .ZN(n26174) );
  INV_X1 U931 ( .A(n17912), .ZN(n26173) );
  INV_X1 U932 ( .A(n17921), .ZN(n26172) );
  INV_X1 U933 ( .A(n17930), .ZN(n26171) );
  INV_X1 U934 ( .A(n18012), .ZN(n26162) );
  INV_X1 U935 ( .A(n18021), .ZN(n26161) );
  INV_X1 U936 ( .A(n18030), .ZN(n26160) );
  INV_X1 U937 ( .A(n18039), .ZN(n26159) );
  INV_X1 U938 ( .A(n18048), .ZN(n26158) );
  INV_X1 U939 ( .A(n18057), .ZN(n26157) );
  INV_X1 U940 ( .A(n18066), .ZN(n26156) );
  INV_X1 U941 ( .A(n18075), .ZN(n26155) );
  INV_X1 U942 ( .A(n18084), .ZN(n26154) );
  INV_X1 U943 ( .A(n18093), .ZN(n26153) );
  INV_X1 U944 ( .A(n18102), .ZN(n26152) );
  INV_X1 U945 ( .A(n18111), .ZN(n26151) );
  INV_X1 U946 ( .A(n18120), .ZN(n26150) );
  INV_X1 U947 ( .A(n18129), .ZN(n26149) );
  INV_X1 U948 ( .A(n18138), .ZN(n26148) );
  INV_X1 U949 ( .A(n18147), .ZN(n26147) );
  INV_X1 U950 ( .A(n18156), .ZN(n26146) );
  INV_X1 U951 ( .A(n18165), .ZN(n26145) );
  INV_X1 U952 ( .A(n18174), .ZN(n26144) );
  INV_X1 U953 ( .A(n18183), .ZN(n26143) );
  INV_X1 U954 ( .A(n18192), .ZN(n26142) );
  INV_X1 U955 ( .A(n18201), .ZN(n26141) );
  INV_X1 U956 ( .A(n18210), .ZN(n26140) );
  INV_X1 U957 ( .A(n18219), .ZN(n26139) );
  INV_X1 U958 ( .A(n18310), .ZN(n26130) );
  INV_X1 U959 ( .A(n18320), .ZN(n26129) );
  INV_X1 U960 ( .A(n18329), .ZN(n26128) );
  INV_X1 U961 ( .A(n18338), .ZN(n26127) );
  INV_X1 U962 ( .A(n18347), .ZN(n26126) );
  INV_X1 U963 ( .A(n18356), .ZN(n26125) );
  INV_X1 U964 ( .A(n18365), .ZN(n26124) );
  INV_X1 U965 ( .A(n18374), .ZN(n26123) );
  INV_X1 U966 ( .A(n18383), .ZN(n26122) );
  INV_X1 U967 ( .A(n18393), .ZN(n26121) );
  INV_X1 U968 ( .A(n18402), .ZN(n26120) );
  INV_X1 U969 ( .A(n18411), .ZN(n26119) );
  INV_X1 U970 ( .A(n18420), .ZN(n26118) );
  INV_X1 U971 ( .A(n18429), .ZN(n26117) );
  INV_X1 U972 ( .A(n18438), .ZN(n26116) );
  INV_X1 U973 ( .A(n18447), .ZN(n26115) );
  INV_X1 U974 ( .A(n18456), .ZN(n26114) );
  INV_X1 U975 ( .A(n18466), .ZN(n26113) );
  INV_X1 U976 ( .A(n18475), .ZN(n26112) );
  INV_X1 U977 ( .A(n18484), .ZN(n26111) );
  INV_X1 U978 ( .A(n18493), .ZN(n26110) );
  INV_X1 U979 ( .A(n18502), .ZN(n26109) );
  INV_X1 U980 ( .A(n18511), .ZN(n26108) );
  INV_X1 U981 ( .A(n18520), .ZN(n26107) );
  INV_X1 U982 ( .A(n9548), .ZN(n27098) );
  INV_X1 U983 ( .A(n9558), .ZN(n27097) );
  INV_X1 U984 ( .A(n9567), .ZN(n27096) );
  INV_X1 U985 ( .A(n9576), .ZN(n27095) );
  INV_X1 U986 ( .A(n9585), .ZN(n27094) );
  INV_X1 U987 ( .A(n9594), .ZN(n27093) );
  INV_X1 U988 ( .A(n9603), .ZN(n27092) );
  INV_X1 U989 ( .A(n9612), .ZN(n27091) );
  INV_X1 U990 ( .A(n9838), .ZN(n27066) );
  INV_X1 U991 ( .A(n9848), .ZN(n27065) );
  INV_X1 U992 ( .A(n9857), .ZN(n27064) );
  INV_X1 U993 ( .A(n9866), .ZN(n27063) );
  INV_X1 U994 ( .A(n9875), .ZN(n27062) );
  INV_X1 U995 ( .A(n9884), .ZN(n27061) );
  INV_X1 U996 ( .A(n9893), .ZN(n27060) );
  INV_X1 U997 ( .A(n9902), .ZN(n27059) );
  INV_X1 U998 ( .A(n10128), .ZN(n27034) );
  INV_X1 U999 ( .A(n10138), .ZN(n27033) );
  INV_X1 U1000 ( .A(n10147), .ZN(n27032) );
  INV_X1 U1001 ( .A(n10156), .ZN(n27031) );
  INV_X1 U1002 ( .A(n10165), .ZN(n27030) );
  INV_X1 U1003 ( .A(n10174), .ZN(n27029) );
  INV_X1 U1004 ( .A(n10183), .ZN(n27028) );
  INV_X1 U1005 ( .A(n10192), .ZN(n27027) );
  INV_X1 U1006 ( .A(n10418), .ZN(n27002) );
  INV_X1 U1007 ( .A(n10428), .ZN(n27001) );
  INV_X1 U1008 ( .A(n10437), .ZN(n27000) );
  INV_X1 U1009 ( .A(n10446), .ZN(n26999) );
  INV_X1 U1010 ( .A(n10455), .ZN(n26998) );
  INV_X1 U1011 ( .A(n10464), .ZN(n26997) );
  INV_X1 U1012 ( .A(n10473), .ZN(n26996) );
  INV_X1 U1013 ( .A(n10482), .ZN(n26995) );
  INV_X1 U1014 ( .A(n10708), .ZN(n26970) );
  INV_X1 U1015 ( .A(n10718), .ZN(n26969) );
  INV_X1 U1016 ( .A(n10727), .ZN(n26968) );
  INV_X1 U1017 ( .A(n10736), .ZN(n26967) );
  INV_X1 U1018 ( .A(n10745), .ZN(n26966) );
  INV_X1 U1019 ( .A(n10754), .ZN(n26965) );
  INV_X1 U1020 ( .A(n10763), .ZN(n26964) );
  INV_X1 U1021 ( .A(n10772), .ZN(n26963) );
  INV_X1 U1022 ( .A(n10998), .ZN(n26938) );
  INV_X1 U1023 ( .A(n11008), .ZN(n26937) );
  INV_X1 U1024 ( .A(n11017), .ZN(n26936) );
  INV_X1 U1025 ( .A(n11026), .ZN(n26935) );
  INV_X1 U1026 ( .A(n11035), .ZN(n26934) );
  INV_X1 U1027 ( .A(n11044), .ZN(n26933) );
  INV_X1 U1028 ( .A(n11053), .ZN(n26932) );
  INV_X1 U1029 ( .A(n11062), .ZN(n26931) );
  INV_X1 U1030 ( .A(n11288), .ZN(n26906) );
  INV_X1 U1031 ( .A(n11298), .ZN(n26905) );
  INV_X1 U1032 ( .A(n11307), .ZN(n26904) );
  INV_X1 U1033 ( .A(n11316), .ZN(n26903) );
  INV_X1 U1034 ( .A(n11325), .ZN(n26902) );
  INV_X1 U1035 ( .A(n11334), .ZN(n26901) );
  INV_X1 U1036 ( .A(n11343), .ZN(n26900) );
  INV_X1 U1037 ( .A(n11352), .ZN(n26899) );
  INV_X1 U1038 ( .A(n11578), .ZN(n26874) );
  INV_X1 U1039 ( .A(n11588), .ZN(n26873) );
  INV_X1 U1040 ( .A(n11597), .ZN(n26872) );
  INV_X1 U1041 ( .A(n11606), .ZN(n26871) );
  INV_X1 U1042 ( .A(n11615), .ZN(n26870) );
  INV_X1 U1043 ( .A(n11624), .ZN(n26869) );
  INV_X1 U1044 ( .A(n11633), .ZN(n26868) );
  INV_X1 U1045 ( .A(n11642), .ZN(n26867) );
  INV_X1 U1046 ( .A(n11868), .ZN(n26842) );
  INV_X1 U1047 ( .A(n11878), .ZN(n26841) );
  INV_X1 U1048 ( .A(n11887), .ZN(n26840) );
  INV_X1 U1049 ( .A(n11896), .ZN(n26839) );
  INV_X1 U1050 ( .A(n11905), .ZN(n26838) );
  INV_X1 U1051 ( .A(n11914), .ZN(n26837) );
  INV_X1 U1052 ( .A(n11923), .ZN(n26836) );
  INV_X1 U1053 ( .A(n11932), .ZN(n26835) );
  INV_X1 U1054 ( .A(n12157), .ZN(n26810) );
  INV_X1 U1055 ( .A(n12167), .ZN(n26809) );
  INV_X1 U1056 ( .A(n12176), .ZN(n26808) );
  INV_X1 U1057 ( .A(n12185), .ZN(n26807) );
  INV_X1 U1058 ( .A(n12194), .ZN(n26806) );
  INV_X1 U1059 ( .A(n12203), .ZN(n26805) );
  INV_X1 U1060 ( .A(n12212), .ZN(n26804) );
  INV_X1 U1061 ( .A(n12221), .ZN(n26803) );
  INV_X1 U1062 ( .A(n12446), .ZN(n26778) );
  INV_X1 U1063 ( .A(n12456), .ZN(n26777) );
  INV_X1 U1064 ( .A(n12465), .ZN(n26776) );
  INV_X1 U1065 ( .A(n12474), .ZN(n26775) );
  INV_X1 U1066 ( .A(n12483), .ZN(n26774) );
  INV_X1 U1067 ( .A(n12492), .ZN(n26773) );
  INV_X1 U1068 ( .A(n12501), .ZN(n26772) );
  INV_X1 U1069 ( .A(n12510), .ZN(n26771) );
  INV_X1 U1070 ( .A(n12735), .ZN(n26746) );
  INV_X1 U1071 ( .A(n12745), .ZN(n26745) );
  INV_X1 U1072 ( .A(n12754), .ZN(n26744) );
  INV_X1 U1073 ( .A(n12763), .ZN(n26743) );
  INV_X1 U1074 ( .A(n12772), .ZN(n26742) );
  INV_X1 U1075 ( .A(n12781), .ZN(n26741) );
  INV_X1 U1076 ( .A(n12790), .ZN(n26740) );
  INV_X1 U1077 ( .A(n12799), .ZN(n26739) );
  INV_X1 U1078 ( .A(n13024), .ZN(n26714) );
  INV_X1 U1079 ( .A(n13034), .ZN(n26713) );
  INV_X1 U1080 ( .A(n13043), .ZN(n26712) );
  INV_X1 U1081 ( .A(n13052), .ZN(n26711) );
  INV_X1 U1082 ( .A(n13061), .ZN(n26710) );
  INV_X1 U1083 ( .A(n13070), .ZN(n26709) );
  INV_X1 U1084 ( .A(n13079), .ZN(n26708) );
  INV_X1 U1085 ( .A(n13088), .ZN(n26707) );
  INV_X1 U1086 ( .A(n13313), .ZN(n26682) );
  INV_X1 U1087 ( .A(n13323), .ZN(n26681) );
  INV_X1 U1088 ( .A(n13332), .ZN(n26680) );
  INV_X1 U1089 ( .A(n13341), .ZN(n26679) );
  INV_X1 U1090 ( .A(n13350), .ZN(n26678) );
  INV_X1 U1091 ( .A(n13359), .ZN(n26677) );
  INV_X1 U1092 ( .A(n13368), .ZN(n26676) );
  INV_X1 U1093 ( .A(n13377), .ZN(n26675) );
  INV_X1 U1094 ( .A(n13602), .ZN(n26650) );
  INV_X1 U1095 ( .A(n13612), .ZN(n26649) );
  INV_X1 U1096 ( .A(n13621), .ZN(n26648) );
  INV_X1 U1097 ( .A(n13630), .ZN(n26647) );
  INV_X1 U1098 ( .A(n13639), .ZN(n26646) );
  INV_X1 U1099 ( .A(n13648), .ZN(n26645) );
  INV_X1 U1100 ( .A(n13657), .ZN(n26644) );
  INV_X1 U1101 ( .A(n13666), .ZN(n26643) );
  INV_X1 U1102 ( .A(n13891), .ZN(n26618) );
  INV_X1 U1103 ( .A(n13901), .ZN(n26617) );
  INV_X1 U1104 ( .A(n13910), .ZN(n26616) );
  INV_X1 U1105 ( .A(n13919), .ZN(n26615) );
  INV_X1 U1106 ( .A(n13928), .ZN(n26614) );
  INV_X1 U1107 ( .A(n13937), .ZN(n26613) );
  INV_X1 U1108 ( .A(n13946), .ZN(n26612) );
  INV_X1 U1109 ( .A(n13955), .ZN(n26611) );
  INV_X1 U1110 ( .A(n14181), .ZN(n26586) );
  INV_X1 U1111 ( .A(n14191), .ZN(n26585) );
  INV_X1 U1112 ( .A(n14200), .ZN(n26584) );
  INV_X1 U1113 ( .A(n14209), .ZN(n26583) );
  INV_X1 U1114 ( .A(n14218), .ZN(n26582) );
  INV_X1 U1115 ( .A(n14227), .ZN(n26581) );
  INV_X1 U1116 ( .A(n14236), .ZN(n26580) );
  INV_X1 U1117 ( .A(n14245), .ZN(n26579) );
  INV_X1 U1118 ( .A(n14470), .ZN(n26554) );
  INV_X1 U1119 ( .A(n14480), .ZN(n26553) );
  INV_X1 U1120 ( .A(n14489), .ZN(n26552) );
  INV_X1 U1121 ( .A(n14498), .ZN(n26551) );
  INV_X1 U1122 ( .A(n14507), .ZN(n26550) );
  INV_X1 U1123 ( .A(n14516), .ZN(n26549) );
  INV_X1 U1124 ( .A(n14525), .ZN(n26548) );
  INV_X1 U1125 ( .A(n14534), .ZN(n26547) );
  INV_X1 U1126 ( .A(n14759), .ZN(n26522) );
  INV_X1 U1127 ( .A(n14769), .ZN(n26521) );
  INV_X1 U1128 ( .A(n14778), .ZN(n26520) );
  INV_X1 U1129 ( .A(n14787), .ZN(n26519) );
  INV_X1 U1130 ( .A(n14796), .ZN(n26518) );
  INV_X1 U1131 ( .A(n14805), .ZN(n26517) );
  INV_X1 U1132 ( .A(n14814), .ZN(n26516) );
  INV_X1 U1133 ( .A(n14823), .ZN(n26515) );
  INV_X1 U1134 ( .A(n15048), .ZN(n26490) );
  INV_X1 U1135 ( .A(n15058), .ZN(n26489) );
  INV_X1 U1136 ( .A(n15067), .ZN(n26488) );
  INV_X1 U1137 ( .A(n15076), .ZN(n26487) );
  INV_X1 U1138 ( .A(n15085), .ZN(n26486) );
  INV_X1 U1139 ( .A(n15094), .ZN(n26485) );
  INV_X1 U1140 ( .A(n15103), .ZN(n26484) );
  INV_X1 U1141 ( .A(n15112), .ZN(n26483) );
  INV_X1 U1142 ( .A(n15337), .ZN(n26458) );
  INV_X1 U1143 ( .A(n15347), .ZN(n26457) );
  INV_X1 U1144 ( .A(n15356), .ZN(n26456) );
  INV_X1 U1145 ( .A(n15365), .ZN(n26455) );
  INV_X1 U1146 ( .A(n15374), .ZN(n26454) );
  INV_X1 U1147 ( .A(n15383), .ZN(n26453) );
  INV_X1 U1148 ( .A(n15392), .ZN(n26452) );
  INV_X1 U1149 ( .A(n15401), .ZN(n26451) );
  INV_X1 U1150 ( .A(n15626), .ZN(n26426) );
  INV_X1 U1151 ( .A(n15636), .ZN(n26425) );
  INV_X1 U1152 ( .A(n15645), .ZN(n26424) );
  INV_X1 U1153 ( .A(n15654), .ZN(n26423) );
  INV_X1 U1154 ( .A(n15663), .ZN(n26422) );
  INV_X1 U1155 ( .A(n15672), .ZN(n26421) );
  INV_X1 U1156 ( .A(n15681), .ZN(n26420) );
  INV_X1 U1157 ( .A(n15690), .ZN(n26419) );
  INV_X1 U1158 ( .A(n15915), .ZN(n26394) );
  INV_X1 U1159 ( .A(n15925), .ZN(n26393) );
  INV_X1 U1160 ( .A(n15934), .ZN(n26392) );
  INV_X1 U1161 ( .A(n15943), .ZN(n26391) );
  INV_X1 U1162 ( .A(n15952), .ZN(n26390) );
  INV_X1 U1163 ( .A(n15961), .ZN(n26389) );
  INV_X1 U1164 ( .A(n15970), .ZN(n26388) );
  INV_X1 U1165 ( .A(n15979), .ZN(n26387) );
  INV_X1 U1166 ( .A(n16204), .ZN(n26362) );
  INV_X1 U1167 ( .A(n16214), .ZN(n26361) );
  INV_X1 U1168 ( .A(n16223), .ZN(n26360) );
  INV_X1 U1169 ( .A(n16232), .ZN(n26359) );
  INV_X1 U1170 ( .A(n16241), .ZN(n26358) );
  INV_X1 U1171 ( .A(n16250), .ZN(n26357) );
  INV_X1 U1172 ( .A(n16259), .ZN(n26356) );
  INV_X1 U1173 ( .A(n16268), .ZN(n26355) );
  INV_X1 U1174 ( .A(n16494), .ZN(n26330) );
  INV_X1 U1175 ( .A(n16504), .ZN(n26329) );
  INV_X1 U1176 ( .A(n16513), .ZN(n26328) );
  INV_X1 U1177 ( .A(n16522), .ZN(n26327) );
  INV_X1 U1178 ( .A(n16531), .ZN(n26326) );
  INV_X1 U1179 ( .A(n16540), .ZN(n26325) );
  INV_X1 U1180 ( .A(n16549), .ZN(n26324) );
  INV_X1 U1181 ( .A(n16558), .ZN(n26323) );
  INV_X1 U1182 ( .A(n16783), .ZN(n26298) );
  INV_X1 U1183 ( .A(n16793), .ZN(n26297) );
  INV_X1 U1184 ( .A(n16802), .ZN(n26296) );
  INV_X1 U1185 ( .A(n16811), .ZN(n26295) );
  INV_X1 U1186 ( .A(n16820), .ZN(n26294) );
  INV_X1 U1187 ( .A(n16829), .ZN(n26293) );
  INV_X1 U1188 ( .A(n16838), .ZN(n26292) );
  INV_X1 U1189 ( .A(n16847), .ZN(n26291) );
  INV_X1 U1190 ( .A(n17072), .ZN(n26266) );
  INV_X1 U1191 ( .A(n17082), .ZN(n26265) );
  INV_X1 U1192 ( .A(n17091), .ZN(n26264) );
  INV_X1 U1193 ( .A(n17100), .ZN(n26263) );
  INV_X1 U1194 ( .A(n17109), .ZN(n26262) );
  INV_X1 U1195 ( .A(n17118), .ZN(n26261) );
  INV_X1 U1196 ( .A(n17127), .ZN(n26260) );
  INV_X1 U1197 ( .A(n17136), .ZN(n26259) );
  INV_X1 U1198 ( .A(n17361), .ZN(n26234) );
  INV_X1 U1199 ( .A(n17371), .ZN(n26233) );
  INV_X1 U1200 ( .A(n17380), .ZN(n26232) );
  INV_X1 U1201 ( .A(n17389), .ZN(n26231) );
  INV_X1 U1202 ( .A(n17398), .ZN(n26230) );
  INV_X1 U1203 ( .A(n17407), .ZN(n26229) );
  INV_X1 U1204 ( .A(n17416), .ZN(n26228) );
  INV_X1 U1205 ( .A(n17425), .ZN(n26227) );
  INV_X1 U1206 ( .A(n17650), .ZN(n26202) );
  INV_X1 U1207 ( .A(n17660), .ZN(n26201) );
  INV_X1 U1208 ( .A(n17669), .ZN(n26200) );
  INV_X1 U1209 ( .A(n17678), .ZN(n26199) );
  INV_X1 U1210 ( .A(n17687), .ZN(n26198) );
  INV_X1 U1211 ( .A(n17696), .ZN(n26197) );
  INV_X1 U1212 ( .A(n17705), .ZN(n26196) );
  INV_X1 U1213 ( .A(n17714), .ZN(n26195) );
  INV_X1 U1214 ( .A(n17939), .ZN(n26170) );
  INV_X1 U1215 ( .A(n17949), .ZN(n26169) );
  INV_X1 U1216 ( .A(n17958), .ZN(n26168) );
  INV_X1 U1217 ( .A(n17967), .ZN(n26167) );
  INV_X1 U1218 ( .A(n17976), .ZN(n26166) );
  INV_X1 U1219 ( .A(n17985), .ZN(n26165) );
  INV_X1 U1220 ( .A(n17994), .ZN(n26164) );
  INV_X1 U1221 ( .A(n18003), .ZN(n26163) );
  INV_X1 U1222 ( .A(n18228), .ZN(n26138) );
  INV_X1 U1223 ( .A(n18240), .ZN(n26137) );
  INV_X1 U1224 ( .A(n18250), .ZN(n26136) );
  INV_X1 U1225 ( .A(n18260), .ZN(n26135) );
  INV_X1 U1226 ( .A(n18270), .ZN(n26134) );
  INV_X1 U1227 ( .A(n18280), .ZN(n26133) );
  INV_X1 U1228 ( .A(n18290), .ZN(n26132) );
  INV_X1 U1229 ( .A(n18300), .ZN(n26131) );
  BUF_X1 U1230 ( .A(n8387), .Z(n8398) );
  BUF_X1 U1231 ( .A(n8387), .Z(n8399) );
  BUF_X1 U1232 ( .A(n8387), .Z(n8400) );
  BUF_X1 U1233 ( .A(n8386), .Z(n8404) );
  BUF_X1 U1234 ( .A(n8386), .Z(n8405) );
  BUF_X1 U1235 ( .A(n8386), .Z(n8406) );
  BUF_X1 U1236 ( .A(n8224), .Z(n8235) );
  BUF_X1 U1237 ( .A(n8224), .Z(n8236) );
  BUF_X1 U1238 ( .A(n8224), .Z(n8237) );
  BUF_X1 U1239 ( .A(n8223), .Z(n8241) );
  BUF_X1 U1240 ( .A(n8223), .Z(n8242) );
  BUF_X1 U1241 ( .A(n8223), .Z(n8243) );
  BUF_X1 U1242 ( .A(n8222), .Z(n8247) );
  BUF_X1 U1243 ( .A(n8222), .Z(n8248) );
  BUF_X1 U1244 ( .A(n8222), .Z(n8249) );
  BUF_X1 U1245 ( .A(n8221), .Z(n8253) );
  BUF_X1 U1246 ( .A(n8221), .Z(n8254) );
  BUF_X1 U1247 ( .A(n8221), .Z(n8255) );
  BUF_X1 U1248 ( .A(n8220), .Z(n8259) );
  BUF_X1 U1249 ( .A(n8220), .Z(n8260) );
  BUF_X1 U1250 ( .A(n8220), .Z(n8261) );
  BUF_X1 U1251 ( .A(n8215), .Z(n8201) );
  BUF_X1 U1252 ( .A(n8200), .Z(n8202) );
  BUF_X1 U1253 ( .A(n8200), .Z(n8203) );
  BUF_X1 U1254 ( .A(n8200), .Z(n8204) );
  BUF_X1 U1255 ( .A(n8200), .Z(n8205) );
  BUF_X1 U1256 ( .A(n8199), .Z(n8207) );
  BUF_X1 U1257 ( .A(n8199), .Z(n8208) );
  BUF_X1 U1258 ( .A(n8199), .Z(n8209) );
  BUF_X1 U1259 ( .A(n8199), .Z(n8210) );
  BUF_X1 U1260 ( .A(n8198), .Z(n8212) );
  BUF_X1 U1261 ( .A(n8198), .Z(n8213) );
  BUF_X1 U1262 ( .A(n8198), .Z(n8214) );
  BUF_X1 U1263 ( .A(n8198), .Z(n8215) );
  BUF_X1 U1264 ( .A(n8388), .Z(n8393) );
  BUF_X1 U1265 ( .A(n8388), .Z(n8394) );
  BUF_X1 U1266 ( .A(n8225), .Z(n8230) );
  BUF_X1 U1267 ( .A(n8225), .Z(n8231) );
  BUF_X1 U1268 ( .A(n8387), .Z(n8395) );
  BUF_X1 U1269 ( .A(n8387), .Z(n8396) );
  BUF_X1 U1270 ( .A(n8387), .Z(n8397) );
  BUF_X1 U1271 ( .A(n8386), .Z(n8401) );
  BUF_X1 U1272 ( .A(n8386), .Z(n8402) );
  BUF_X1 U1273 ( .A(n8386), .Z(n8403) );
  BUF_X1 U1274 ( .A(n8224), .Z(n8232) );
  BUF_X1 U1275 ( .A(n8224), .Z(n8233) );
  BUF_X1 U1276 ( .A(n8224), .Z(n8234) );
  BUF_X1 U1277 ( .A(n8223), .Z(n8238) );
  BUF_X1 U1278 ( .A(n8223), .Z(n8239) );
  BUF_X1 U1279 ( .A(n8223), .Z(n8240) );
  BUF_X1 U1280 ( .A(n8222), .Z(n8244) );
  BUF_X1 U1281 ( .A(n8222), .Z(n8245) );
  BUF_X1 U1282 ( .A(n8222), .Z(n8246) );
  BUF_X1 U1283 ( .A(n8221), .Z(n8250) );
  BUF_X1 U1284 ( .A(n8221), .Z(n8251) );
  BUF_X1 U1285 ( .A(n8221), .Z(n8252) );
  BUF_X1 U1286 ( .A(n8220), .Z(n8256) );
  BUF_X1 U1287 ( .A(n8220), .Z(n8257) );
  BUF_X1 U1288 ( .A(n8220), .Z(n8258) );
  BUF_X1 U1289 ( .A(n8199), .Z(n8206) );
  BUF_X1 U1290 ( .A(n8198), .Z(n8211) );
  BUF_X1 U1291 ( .A(n8388), .Z(n8390) );
  BUF_X1 U1292 ( .A(n8388), .Z(n8391) );
  BUF_X1 U1293 ( .A(n8388), .Z(n8392) );
  BUF_X1 U1294 ( .A(n8225), .Z(n8227) );
  BUF_X1 U1295 ( .A(n8225), .Z(n8228) );
  BUF_X1 U1296 ( .A(n8225), .Z(n8229) );
  BUF_X1 U1297 ( .A(n8197), .Z(n8216) );
  BUF_X1 U1298 ( .A(n8197), .Z(n8217) );
  BUF_X1 U1299 ( .A(n8197), .Z(n8218) );
  BUF_X1 U1300 ( .A(n8237), .Z(n8262) );
  BUF_X1 U1301 ( .A(n8358), .Z(n8385) );
  BUF_X1 U1302 ( .A(n8358), .Z(n8384) );
  BUF_X1 U1303 ( .A(n8358), .Z(n8383) );
  BUF_X1 U1304 ( .A(n8359), .Z(n8382) );
  BUF_X1 U1305 ( .A(n8359), .Z(n8381) );
  BUF_X1 U1306 ( .A(n8359), .Z(n8380) );
  BUF_X1 U1307 ( .A(n8360), .Z(n8379) );
  BUF_X1 U1308 ( .A(n8360), .Z(n8378) );
  BUF_X1 U1309 ( .A(n8360), .Z(n8377) );
  BUF_X1 U1310 ( .A(n8361), .Z(n8376) );
  BUF_X1 U1311 ( .A(n8361), .Z(n8375) );
  BUF_X1 U1312 ( .A(n8361), .Z(n8374) );
  BUF_X1 U1313 ( .A(n8362), .Z(n8373) );
  BUF_X1 U1314 ( .A(n8362), .Z(n8372) );
  BUF_X1 U1315 ( .A(n8362), .Z(n8371) );
  BUF_X1 U1316 ( .A(n8363), .Z(n8370) );
  BUF_X1 U1317 ( .A(n8363), .Z(n8369) );
  BUF_X1 U1318 ( .A(n8363), .Z(n8368) );
  BUF_X1 U1319 ( .A(n8364), .Z(n8367) );
  BUF_X1 U1320 ( .A(n8364), .Z(n8366) );
  BUF_X1 U1321 ( .A(n8364), .Z(n8365) );
  BUF_X1 U1322 ( .A(n8270), .Z(n8282) );
  BUF_X1 U1323 ( .A(n8266), .Z(n8281) );
  BUF_X1 U1324 ( .A(n8266), .Z(n8280) );
  BUF_X1 U1325 ( .A(n8266), .Z(n8279) );
  BUF_X1 U1326 ( .A(n8267), .Z(n8278) );
  BUF_X1 U1327 ( .A(n8267), .Z(n8277) );
  BUF_X1 U1328 ( .A(n8267), .Z(n8276) );
  BUF_X1 U1329 ( .A(n8268), .Z(n8275) );
  BUF_X1 U1330 ( .A(n8268), .Z(n8274) );
  BUF_X1 U1331 ( .A(n8268), .Z(n8273) );
  BUF_X1 U1332 ( .A(n8269), .Z(n8272) );
  BUF_X1 U1333 ( .A(n8269), .Z(n8271) );
  BUF_X1 U1334 ( .A(n8269), .Z(n8270) );
  NAND2_X1 U1335 ( .A1(n9232), .A2(n9233), .ZN(n9224) );
  NAND2_X1 U1336 ( .A1(n9243), .A2(n9233), .ZN(n9235) );
  NAND2_X1 U1337 ( .A1(n9253), .A2(n9233), .ZN(n9245) );
  NAND2_X1 U1338 ( .A1(n9263), .A2(n9233), .ZN(n9255) );
  NAND2_X1 U1339 ( .A1(n9273), .A2(n9233), .ZN(n9265) );
  NAND2_X1 U1340 ( .A1(n9283), .A2(n9233), .ZN(n9275) );
  NAND2_X1 U1341 ( .A1(n9293), .A2(n9233), .ZN(n9285) );
  NAND2_X1 U1342 ( .A1(n8595), .A2(n9233), .ZN(n9295) );
  NAND2_X1 U1343 ( .A1(n9556), .A2(n9232), .ZN(n9548) );
  NAND2_X1 U1344 ( .A1(n9556), .A2(n9243), .ZN(n9558) );
  NAND2_X1 U1345 ( .A1(n9556), .A2(n9253), .ZN(n9567) );
  NAND2_X1 U1346 ( .A1(n9556), .A2(n9263), .ZN(n9576) );
  NAND2_X1 U1347 ( .A1(n9556), .A2(n8598), .ZN(n9585) );
  NAND2_X1 U1348 ( .A1(n9556), .A2(n9283), .ZN(n9594) );
  NAND2_X1 U1349 ( .A1(n9556), .A2(n9293), .ZN(n9603) );
  NAND2_X1 U1350 ( .A1(n9556), .A2(n8595), .ZN(n9612) );
  NAND2_X1 U1351 ( .A1(n9556), .A2(n9313), .ZN(n9621) );
  NAND2_X1 U1352 ( .A1(n9556), .A2(n9323), .ZN(n9630) );
  NAND2_X1 U1353 ( .A1(n9556), .A2(n9333), .ZN(n9639) );
  NAND2_X1 U1354 ( .A1(n9556), .A2(n9343), .ZN(n9648) );
  NAND2_X1 U1355 ( .A1(n9556), .A2(n9353), .ZN(n9657) );
  NAND2_X1 U1356 ( .A1(n9556), .A2(n9363), .ZN(n9666) );
  NAND2_X1 U1357 ( .A1(n9556), .A2(n8588), .ZN(n9675) );
  NAND2_X1 U1358 ( .A1(n9556), .A2(n9383), .ZN(n9684) );
  NAND2_X1 U1359 ( .A1(n9556), .A2(n9393), .ZN(n9693) );
  NAND2_X1 U1360 ( .A1(n9556), .A2(n8585), .ZN(n9702) );
  NAND2_X1 U1361 ( .A1(n9556), .A2(n9413), .ZN(n9711) );
  NAND2_X1 U1362 ( .A1(n9556), .A2(n9423), .ZN(n9720) );
  NAND2_X1 U1363 ( .A1(n8570), .A2(n9433), .ZN(n9729) );
  NAND2_X1 U1364 ( .A1(n8570), .A2(n9443), .ZN(n9738) );
  NAND2_X1 U1365 ( .A1(n8570), .A2(n9453), .ZN(n9747) );
  NAND2_X1 U1366 ( .A1(n8570), .A2(n9463), .ZN(n9756) );
  NAND2_X1 U1367 ( .A1(n8570), .A2(n8578), .ZN(n9765) );
  NAND2_X1 U1368 ( .A1(n8570), .A2(n9483), .ZN(n9774) );
  NAND2_X1 U1369 ( .A1(n8570), .A2(n9493), .ZN(n9783) );
  NAND2_X1 U1370 ( .A1(n8570), .A2(n8575), .ZN(n9792) );
  NAND2_X1 U1371 ( .A1(n8570), .A2(n9513), .ZN(n9801) );
  NAND2_X1 U1372 ( .A1(n8570), .A2(n9523), .ZN(n9810) );
  NAND2_X1 U1373 ( .A1(n8570), .A2(n9533), .ZN(n9819) );
  NAND2_X1 U1374 ( .A1(n8570), .A2(n9543), .ZN(n9828) );
  NAND2_X1 U1375 ( .A1(n9846), .A2(n9232), .ZN(n9838) );
  NAND2_X1 U1376 ( .A1(n9846), .A2(n9243), .ZN(n9848) );
  NAND2_X1 U1377 ( .A1(n9846), .A2(n9253), .ZN(n9857) );
  NAND2_X1 U1378 ( .A1(n9846), .A2(n9263), .ZN(n9866) );
  NAND2_X1 U1379 ( .A1(n9846), .A2(n9273), .ZN(n9875) );
  NAND2_X1 U1380 ( .A1(n9846), .A2(n9283), .ZN(n9884) );
  NAND2_X1 U1381 ( .A1(n9846), .A2(n9293), .ZN(n9893) );
  NAND2_X1 U1382 ( .A1(n9846), .A2(n8595), .ZN(n9902) );
  NAND2_X1 U1383 ( .A1(n8569), .A2(n9313), .ZN(n9911) );
  NAND2_X1 U1384 ( .A1(n8569), .A2(n9323), .ZN(n9920) );
  NAND2_X1 U1385 ( .A1(n8569), .A2(n9333), .ZN(n9929) );
  NAND2_X1 U1386 ( .A1(n8569), .A2(n9343), .ZN(n9938) );
  NAND2_X1 U1387 ( .A1(n8569), .A2(n9353), .ZN(n9947) );
  NAND2_X1 U1388 ( .A1(n8569), .A2(n9363), .ZN(n9956) );
  NAND2_X1 U1389 ( .A1(n8569), .A2(n9373), .ZN(n9965) );
  NAND2_X1 U1390 ( .A1(n8569), .A2(n9383), .ZN(n9974) );
  NAND2_X1 U1391 ( .A1(n8569), .A2(n9393), .ZN(n9983) );
  NAND2_X1 U1392 ( .A1(n8569), .A2(n8585), .ZN(n9992) );
  NAND2_X1 U1393 ( .A1(n8569), .A2(n9413), .ZN(n10001) );
  NAND2_X1 U1394 ( .A1(n8569), .A2(n9423), .ZN(n10010) );
  NAND2_X1 U1395 ( .A1(n9846), .A2(n9433), .ZN(n10019) );
  NAND2_X1 U1396 ( .A1(n9846), .A2(n9443), .ZN(n10028) );
  NAND2_X1 U1397 ( .A1(n9846), .A2(n9453), .ZN(n10037) );
  NAND2_X1 U1398 ( .A1(n9846), .A2(n9463), .ZN(n10046) );
  NAND2_X1 U1399 ( .A1(n9846), .A2(n9473), .ZN(n10055) );
  NAND2_X1 U1400 ( .A1(n9846), .A2(n9483), .ZN(n10064) );
  NAND2_X1 U1401 ( .A1(n9846), .A2(n9493), .ZN(n10073) );
  NAND2_X1 U1402 ( .A1(n9846), .A2(n8575), .ZN(n10082) );
  NAND2_X1 U1403 ( .A1(n9846), .A2(n9513), .ZN(n10091) );
  NAND2_X1 U1404 ( .A1(n9846), .A2(n9523), .ZN(n10100) );
  NAND2_X1 U1405 ( .A1(n9846), .A2(n9533), .ZN(n10109) );
  NAND2_X1 U1406 ( .A1(n9846), .A2(n9543), .ZN(n10118) );
  NAND2_X1 U1407 ( .A1(n10136), .A2(n9232), .ZN(n10128) );
  NAND2_X1 U1408 ( .A1(n10136), .A2(n9243), .ZN(n10138) );
  NAND2_X1 U1409 ( .A1(n10136), .A2(n9253), .ZN(n10147) );
  NAND2_X1 U1410 ( .A1(n10136), .A2(n9263), .ZN(n10156) );
  NAND2_X1 U1411 ( .A1(n10136), .A2(n8598), .ZN(n10165) );
  NAND2_X1 U1412 ( .A1(n10136), .A2(n9283), .ZN(n10174) );
  NAND2_X1 U1413 ( .A1(n10136), .A2(n9293), .ZN(n10183) );
  NAND2_X1 U1414 ( .A1(n10136), .A2(n8595), .ZN(n10192) );
  NAND2_X1 U1415 ( .A1(n8568), .A2(n9313), .ZN(n10201) );
  NAND2_X1 U1416 ( .A1(n8568), .A2(n9323), .ZN(n10210) );
  NAND2_X1 U1417 ( .A1(n8568), .A2(n9333), .ZN(n10219) );
  NAND2_X1 U1418 ( .A1(n8568), .A2(n9343), .ZN(n10228) );
  NAND2_X1 U1419 ( .A1(n8568), .A2(n9353), .ZN(n10237) );
  NAND2_X1 U1420 ( .A1(n8568), .A2(n9363), .ZN(n10246) );
  NAND2_X1 U1421 ( .A1(n8568), .A2(n8588), .ZN(n10255) );
  NAND2_X1 U1422 ( .A1(n8568), .A2(n9383), .ZN(n10264) );
  NAND2_X1 U1423 ( .A1(n8568), .A2(n9393), .ZN(n10273) );
  NAND2_X1 U1424 ( .A1(n8568), .A2(n8585), .ZN(n10282) );
  NAND2_X1 U1425 ( .A1(n8568), .A2(n9413), .ZN(n10291) );
  NAND2_X1 U1426 ( .A1(n8568), .A2(n9423), .ZN(n10300) );
  NAND2_X1 U1427 ( .A1(n10136), .A2(n9433), .ZN(n10309) );
  NAND2_X1 U1428 ( .A1(n10136), .A2(n9443), .ZN(n10318) );
  NAND2_X1 U1429 ( .A1(n10136), .A2(n9453), .ZN(n10327) );
  NAND2_X1 U1430 ( .A1(n10136), .A2(n9463), .ZN(n10336) );
  NAND2_X1 U1431 ( .A1(n10136), .A2(n8578), .ZN(n10345) );
  NAND2_X1 U1432 ( .A1(n10136), .A2(n9483), .ZN(n10354) );
  NAND2_X1 U1433 ( .A1(n10136), .A2(n9493), .ZN(n10363) );
  NAND2_X1 U1434 ( .A1(n10136), .A2(n8575), .ZN(n10372) );
  NAND2_X1 U1435 ( .A1(n10136), .A2(n9513), .ZN(n10381) );
  NAND2_X1 U1436 ( .A1(n10136), .A2(n9523), .ZN(n10390) );
  NAND2_X1 U1437 ( .A1(n10136), .A2(n9533), .ZN(n10399) );
  NAND2_X1 U1438 ( .A1(n10136), .A2(n9543), .ZN(n10408) );
  NAND2_X1 U1439 ( .A1(n8567), .A2(n9232), .ZN(n10418) );
  NAND2_X1 U1440 ( .A1(n8567), .A2(n9243), .ZN(n10428) );
  NAND2_X1 U1441 ( .A1(n8567), .A2(n9253), .ZN(n10437) );
  NAND2_X1 U1442 ( .A1(n8567), .A2(n9263), .ZN(n10446) );
  NAND2_X1 U1443 ( .A1(n8567), .A2(n9273), .ZN(n10455) );
  NAND2_X1 U1444 ( .A1(n8567), .A2(n9283), .ZN(n10464) );
  NAND2_X1 U1445 ( .A1(n8567), .A2(n9293), .ZN(n10473) );
  NAND2_X1 U1446 ( .A1(n8567), .A2(n8595), .ZN(n10482) );
  NAND2_X1 U1447 ( .A1(n10426), .A2(n9313), .ZN(n10491) );
  NAND2_X1 U1448 ( .A1(n10426), .A2(n9323), .ZN(n10500) );
  NAND2_X1 U1449 ( .A1(n10426), .A2(n9333), .ZN(n10509) );
  NAND2_X1 U1450 ( .A1(n10426), .A2(n9343), .ZN(n10518) );
  NAND2_X1 U1451 ( .A1(n10426), .A2(n9353), .ZN(n10527) );
  NAND2_X1 U1452 ( .A1(n10426), .A2(n9363), .ZN(n10536) );
  NAND2_X1 U1453 ( .A1(n10426), .A2(n9373), .ZN(n10545) );
  NAND2_X1 U1454 ( .A1(n10426), .A2(n9383), .ZN(n10554) );
  NAND2_X1 U1455 ( .A1(n10426), .A2(n9393), .ZN(n10563) );
  NAND2_X1 U1456 ( .A1(n10426), .A2(n8585), .ZN(n10572) );
  NAND2_X1 U1457 ( .A1(n10426), .A2(n9413), .ZN(n10581) );
  NAND2_X1 U1458 ( .A1(n10426), .A2(n9423), .ZN(n10590) );
  NAND2_X1 U1459 ( .A1(n8567), .A2(n9433), .ZN(n10599) );
  NAND2_X1 U1460 ( .A1(n8567), .A2(n9443), .ZN(n10608) );
  NAND2_X1 U1461 ( .A1(n8567), .A2(n9453), .ZN(n10617) );
  NAND2_X1 U1462 ( .A1(n8567), .A2(n9463), .ZN(n10626) );
  NAND2_X1 U1463 ( .A1(n10426), .A2(n9473), .ZN(n10635) );
  NAND2_X1 U1464 ( .A1(n10426), .A2(n9483), .ZN(n10644) );
  NAND2_X1 U1465 ( .A1(n10426), .A2(n9493), .ZN(n10653) );
  NAND2_X1 U1466 ( .A1(n10426), .A2(n8575), .ZN(n10662) );
  NAND2_X1 U1467 ( .A1(n10426), .A2(n9513), .ZN(n10671) );
  NAND2_X1 U1468 ( .A1(n10426), .A2(n9523), .ZN(n10680) );
  NAND2_X1 U1469 ( .A1(n10426), .A2(n9533), .ZN(n10689) );
  NAND2_X1 U1470 ( .A1(n10426), .A2(n9543), .ZN(n10698) );
  NAND2_X1 U1471 ( .A1(n10716), .A2(n9232), .ZN(n10708) );
  NAND2_X1 U1472 ( .A1(n10716), .A2(n9243), .ZN(n10718) );
  NAND2_X1 U1473 ( .A1(n10716), .A2(n9253), .ZN(n10727) );
  NAND2_X1 U1474 ( .A1(n10716), .A2(n9263), .ZN(n10736) );
  NAND2_X1 U1475 ( .A1(n10716), .A2(n8598), .ZN(n10745) );
  NAND2_X1 U1476 ( .A1(n10716), .A2(n9283), .ZN(n10754) );
  NAND2_X1 U1477 ( .A1(n10716), .A2(n9293), .ZN(n10763) );
  NAND2_X1 U1478 ( .A1(n10716), .A2(n8595), .ZN(n10772) );
  NAND2_X1 U1479 ( .A1(n8566), .A2(n9313), .ZN(n10781) );
  NAND2_X1 U1480 ( .A1(n8566), .A2(n9323), .ZN(n10790) );
  NAND2_X1 U1481 ( .A1(n8566), .A2(n9333), .ZN(n10799) );
  NAND2_X1 U1482 ( .A1(n8566), .A2(n9343), .ZN(n10808) );
  NAND2_X1 U1483 ( .A1(n8566), .A2(n9353), .ZN(n10817) );
  NAND2_X1 U1484 ( .A1(n8566), .A2(n9363), .ZN(n10826) );
  NAND2_X1 U1485 ( .A1(n8566), .A2(n8588), .ZN(n10835) );
  NAND2_X1 U1486 ( .A1(n8566), .A2(n9383), .ZN(n10844) );
  NAND2_X1 U1487 ( .A1(n8566), .A2(n9393), .ZN(n10853) );
  NAND2_X1 U1488 ( .A1(n8566), .A2(n8585), .ZN(n10862) );
  NAND2_X1 U1489 ( .A1(n8566), .A2(n9413), .ZN(n10871) );
  NAND2_X1 U1490 ( .A1(n8566), .A2(n9423), .ZN(n10880) );
  NAND2_X1 U1491 ( .A1(n10716), .A2(n9433), .ZN(n10889) );
  NAND2_X1 U1492 ( .A1(n10716), .A2(n9443), .ZN(n10898) );
  NAND2_X1 U1493 ( .A1(n10716), .A2(n9453), .ZN(n10907) );
  NAND2_X1 U1494 ( .A1(n10716), .A2(n9463), .ZN(n10916) );
  NAND2_X1 U1495 ( .A1(n10716), .A2(n8578), .ZN(n10925) );
  NAND2_X1 U1496 ( .A1(n10716), .A2(n9483), .ZN(n10934) );
  NAND2_X1 U1497 ( .A1(n10716), .A2(n9493), .ZN(n10943) );
  NAND2_X1 U1498 ( .A1(n10716), .A2(n8575), .ZN(n10952) );
  NAND2_X1 U1499 ( .A1(n10716), .A2(n9513), .ZN(n10961) );
  NAND2_X1 U1500 ( .A1(n10716), .A2(n9523), .ZN(n10970) );
  NAND2_X1 U1501 ( .A1(n10716), .A2(n9533), .ZN(n10979) );
  NAND2_X1 U1502 ( .A1(n10716), .A2(n9543), .ZN(n10988) );
  NAND2_X1 U1503 ( .A1(n11006), .A2(n9232), .ZN(n10998) );
  NAND2_X1 U1504 ( .A1(n11006), .A2(n9243), .ZN(n11008) );
  NAND2_X1 U1505 ( .A1(n11006), .A2(n9253), .ZN(n11017) );
  NAND2_X1 U1506 ( .A1(n11006), .A2(n9263), .ZN(n11026) );
  NAND2_X1 U1507 ( .A1(n11006), .A2(n9273), .ZN(n11035) );
  NAND2_X1 U1508 ( .A1(n11006), .A2(n9283), .ZN(n11044) );
  NAND2_X1 U1509 ( .A1(n11006), .A2(n9293), .ZN(n11053) );
  NAND2_X1 U1510 ( .A1(n11006), .A2(n8595), .ZN(n11062) );
  NAND2_X1 U1511 ( .A1(n8565), .A2(n9313), .ZN(n11071) );
  NAND2_X1 U1512 ( .A1(n8565), .A2(n9323), .ZN(n11080) );
  NAND2_X1 U1513 ( .A1(n8565), .A2(n9333), .ZN(n11089) );
  NAND2_X1 U1514 ( .A1(n8565), .A2(n9343), .ZN(n11098) );
  NAND2_X1 U1515 ( .A1(n8565), .A2(n9353), .ZN(n11107) );
  NAND2_X1 U1516 ( .A1(n8565), .A2(n9363), .ZN(n11116) );
  NAND2_X1 U1517 ( .A1(n8565), .A2(n9373), .ZN(n11125) );
  NAND2_X1 U1518 ( .A1(n8565), .A2(n9383), .ZN(n11134) );
  NAND2_X1 U1519 ( .A1(n8565), .A2(n9393), .ZN(n11143) );
  NAND2_X1 U1520 ( .A1(n8565), .A2(n8585), .ZN(n11152) );
  NAND2_X1 U1521 ( .A1(n8565), .A2(n9413), .ZN(n11161) );
  NAND2_X1 U1522 ( .A1(n8565), .A2(n9423), .ZN(n11170) );
  NAND2_X1 U1523 ( .A1(n11006), .A2(n9433), .ZN(n11179) );
  NAND2_X1 U1524 ( .A1(n11006), .A2(n9443), .ZN(n11188) );
  NAND2_X1 U1525 ( .A1(n11006), .A2(n9453), .ZN(n11197) );
  NAND2_X1 U1526 ( .A1(n11006), .A2(n9463), .ZN(n11206) );
  NAND2_X1 U1527 ( .A1(n11006), .A2(n9473), .ZN(n11215) );
  NAND2_X1 U1528 ( .A1(n11006), .A2(n9483), .ZN(n11224) );
  NAND2_X1 U1529 ( .A1(n11006), .A2(n9493), .ZN(n11233) );
  NAND2_X1 U1530 ( .A1(n11006), .A2(n8575), .ZN(n11242) );
  NAND2_X1 U1531 ( .A1(n11006), .A2(n9513), .ZN(n11251) );
  NAND2_X1 U1532 ( .A1(n11006), .A2(n9523), .ZN(n11260) );
  NAND2_X1 U1533 ( .A1(n11006), .A2(n9533), .ZN(n11269) );
  NAND2_X1 U1534 ( .A1(n11006), .A2(n9543), .ZN(n11278) );
  NAND2_X1 U1535 ( .A1(n11296), .A2(n9232), .ZN(n11288) );
  NAND2_X1 U1536 ( .A1(n11296), .A2(n9243), .ZN(n11298) );
  NAND2_X1 U1537 ( .A1(n11296), .A2(n9253), .ZN(n11307) );
  NAND2_X1 U1538 ( .A1(n11296), .A2(n9263), .ZN(n11316) );
  NAND2_X1 U1539 ( .A1(n11296), .A2(n8598), .ZN(n11325) );
  NAND2_X1 U1540 ( .A1(n11296), .A2(n9283), .ZN(n11334) );
  NAND2_X1 U1541 ( .A1(n11296), .A2(n9293), .ZN(n11343) );
  NAND2_X1 U1542 ( .A1(n11296), .A2(n8595), .ZN(n11352) );
  NAND2_X1 U1543 ( .A1(n8564), .A2(n9313), .ZN(n11361) );
  NAND2_X1 U1544 ( .A1(n8564), .A2(n9323), .ZN(n11370) );
  NAND2_X1 U1545 ( .A1(n8564), .A2(n9333), .ZN(n11379) );
  NAND2_X1 U1546 ( .A1(n8564), .A2(n9343), .ZN(n11388) );
  NAND2_X1 U1547 ( .A1(n8564), .A2(n9353), .ZN(n11397) );
  NAND2_X1 U1548 ( .A1(n8564), .A2(n9363), .ZN(n11406) );
  NAND2_X1 U1549 ( .A1(n8564), .A2(n8588), .ZN(n11415) );
  NAND2_X1 U1550 ( .A1(n8564), .A2(n9383), .ZN(n11424) );
  NAND2_X1 U1551 ( .A1(n8564), .A2(n9393), .ZN(n11433) );
  NAND2_X1 U1552 ( .A1(n8564), .A2(n8585), .ZN(n11442) );
  NAND2_X1 U1553 ( .A1(n8564), .A2(n9413), .ZN(n11451) );
  NAND2_X1 U1554 ( .A1(n8564), .A2(n9423), .ZN(n11460) );
  NAND2_X1 U1555 ( .A1(n11296), .A2(n9433), .ZN(n11469) );
  NAND2_X1 U1556 ( .A1(n11296), .A2(n9443), .ZN(n11478) );
  NAND2_X1 U1557 ( .A1(n11296), .A2(n9453), .ZN(n11487) );
  NAND2_X1 U1558 ( .A1(n11296), .A2(n9463), .ZN(n11496) );
  NAND2_X1 U1559 ( .A1(n11296), .A2(n8578), .ZN(n11505) );
  NAND2_X1 U1560 ( .A1(n11296), .A2(n9483), .ZN(n11514) );
  NAND2_X1 U1561 ( .A1(n11296), .A2(n9493), .ZN(n11523) );
  NAND2_X1 U1562 ( .A1(n11296), .A2(n8575), .ZN(n11532) );
  NAND2_X1 U1563 ( .A1(n11296), .A2(n9513), .ZN(n11541) );
  NAND2_X1 U1564 ( .A1(n11296), .A2(n9523), .ZN(n11550) );
  NAND2_X1 U1565 ( .A1(n11296), .A2(n9533), .ZN(n11559) );
  NAND2_X1 U1566 ( .A1(n11296), .A2(n9543), .ZN(n11568) );
  NAND2_X1 U1567 ( .A1(n9313), .A2(n8602), .ZN(n9305) );
  NAND2_X1 U1568 ( .A1(n9323), .A2(n8602), .ZN(n9315) );
  NAND2_X1 U1569 ( .A1(n9333), .A2(n8602), .ZN(n9325) );
  NAND2_X1 U1570 ( .A1(n9343), .A2(n8602), .ZN(n9335) );
  NAND2_X1 U1571 ( .A1(n9353), .A2(n8602), .ZN(n9345) );
  NAND2_X1 U1572 ( .A1(n9363), .A2(n8602), .ZN(n9355) );
  NAND2_X1 U1573 ( .A1(n9373), .A2(n8602), .ZN(n9365) );
  NAND2_X1 U1574 ( .A1(n9383), .A2(n8602), .ZN(n9375) );
  NAND2_X1 U1575 ( .A1(n9393), .A2(n8602), .ZN(n9385) );
  NAND2_X1 U1576 ( .A1(n8585), .A2(n8602), .ZN(n9395) );
  NAND2_X1 U1577 ( .A1(n9413), .A2(n8602), .ZN(n9405) );
  NAND2_X1 U1578 ( .A1(n9423), .A2(n8602), .ZN(n9415) );
  NAND2_X1 U1579 ( .A1(n9433), .A2(n9233), .ZN(n9425) );
  NAND2_X1 U1580 ( .A1(n9443), .A2(n9233), .ZN(n9435) );
  NAND2_X1 U1581 ( .A1(n9453), .A2(n9233), .ZN(n9445) );
  NAND2_X1 U1582 ( .A1(n9463), .A2(n9233), .ZN(n9455) );
  NAND2_X1 U1583 ( .A1(n9473), .A2(n9233), .ZN(n9465) );
  NAND2_X1 U1584 ( .A1(n9483), .A2(n9233), .ZN(n9475) );
  NAND2_X1 U1585 ( .A1(n9493), .A2(n9233), .ZN(n9485) );
  NAND2_X1 U1586 ( .A1(n8575), .A2(n9233), .ZN(n9495) );
  NAND2_X1 U1587 ( .A1(n9513), .A2(n9233), .ZN(n9505) );
  NAND2_X1 U1588 ( .A1(n9523), .A2(n9233), .ZN(n9515) );
  NAND2_X1 U1589 ( .A1(n9533), .A2(n9233), .ZN(n9525) );
  NAND2_X1 U1590 ( .A1(n9543), .A2(n9233), .ZN(n9535) );
  NAND2_X1 U1591 ( .A1(n11586), .A2(n8603), .ZN(n11578) );
  NAND2_X1 U1592 ( .A1(n11586), .A2(n8601), .ZN(n11588) );
  NAND2_X1 U1593 ( .A1(n11586), .A2(n8600), .ZN(n11597) );
  NAND2_X1 U1594 ( .A1(n11586), .A2(n8599), .ZN(n11606) );
  NAND2_X1 U1595 ( .A1(n11586), .A2(n9273), .ZN(n11615) );
  NAND2_X1 U1596 ( .A1(n11586), .A2(n8597), .ZN(n11624) );
  NAND2_X1 U1597 ( .A1(n11586), .A2(n8596), .ZN(n11633) );
  NAND2_X1 U1598 ( .A1(n11586), .A2(n9303), .ZN(n11642) );
  NAND2_X1 U1599 ( .A1(n8563), .A2(n8594), .ZN(n11651) );
  NAND2_X1 U1600 ( .A1(n8563), .A2(n8593), .ZN(n11660) );
  NAND2_X1 U1601 ( .A1(n8563), .A2(n8592), .ZN(n11669) );
  NAND2_X1 U1602 ( .A1(n8563), .A2(n8591), .ZN(n11678) );
  NAND2_X1 U1603 ( .A1(n8563), .A2(n8590), .ZN(n11687) );
  NAND2_X1 U1604 ( .A1(n8563), .A2(n8589), .ZN(n11696) );
  NAND2_X1 U1605 ( .A1(n8563), .A2(n9373), .ZN(n11705) );
  NAND2_X1 U1606 ( .A1(n8563), .A2(n8587), .ZN(n11714) );
  NAND2_X1 U1607 ( .A1(n8563), .A2(n8586), .ZN(n11723) );
  NAND2_X1 U1608 ( .A1(n8563), .A2(n9403), .ZN(n11732) );
  NAND2_X1 U1609 ( .A1(n8563), .A2(n8584), .ZN(n11741) );
  NAND2_X1 U1610 ( .A1(n8563), .A2(n8583), .ZN(n11750) );
  NAND2_X1 U1611 ( .A1(n11586), .A2(n8582), .ZN(n11759) );
  NAND2_X1 U1612 ( .A1(n11586), .A2(n8581), .ZN(n11768) );
  NAND2_X1 U1613 ( .A1(n11586), .A2(n8580), .ZN(n11777) );
  NAND2_X1 U1614 ( .A1(n11586), .A2(n8579), .ZN(n11786) );
  NAND2_X1 U1615 ( .A1(n11586), .A2(n9473), .ZN(n11795) );
  NAND2_X1 U1616 ( .A1(n11586), .A2(n8577), .ZN(n11804) );
  NAND2_X1 U1617 ( .A1(n11586), .A2(n8576), .ZN(n11813) );
  NAND2_X1 U1618 ( .A1(n11586), .A2(n9503), .ZN(n11822) );
  NAND2_X1 U1619 ( .A1(n11586), .A2(n8574), .ZN(n11831) );
  NAND2_X1 U1620 ( .A1(n11586), .A2(n8573), .ZN(n11840) );
  NAND2_X1 U1621 ( .A1(n11586), .A2(n8572), .ZN(n11849) );
  NAND2_X1 U1622 ( .A1(n11586), .A2(n8571), .ZN(n11858) );
  NAND2_X1 U1623 ( .A1(n11876), .A2(n8603), .ZN(n11868) );
  NAND2_X1 U1624 ( .A1(n11876), .A2(n8601), .ZN(n11878) );
  NAND2_X1 U1625 ( .A1(n11876), .A2(n8600), .ZN(n11887) );
  NAND2_X1 U1626 ( .A1(n11876), .A2(n8599), .ZN(n11896) );
  NAND2_X1 U1627 ( .A1(n11876), .A2(n9273), .ZN(n11905) );
  NAND2_X1 U1628 ( .A1(n11876), .A2(n8597), .ZN(n11914) );
  NAND2_X1 U1629 ( .A1(n11876), .A2(n8596), .ZN(n11923) );
  NAND2_X1 U1630 ( .A1(n11876), .A2(n9303), .ZN(n11932) );
  NAND2_X1 U1631 ( .A1(n8562), .A2(n8594), .ZN(n11941) );
  NAND2_X1 U1632 ( .A1(n8562), .A2(n8593), .ZN(n11950) );
  NAND2_X1 U1633 ( .A1(n8562), .A2(n8592), .ZN(n11959) );
  NAND2_X1 U1634 ( .A1(n8562), .A2(n8591), .ZN(n11968) );
  NAND2_X1 U1635 ( .A1(n8562), .A2(n8590), .ZN(n11977) );
  NAND2_X1 U1636 ( .A1(n8562), .A2(n8589), .ZN(n11986) );
  NAND2_X1 U1637 ( .A1(n8562), .A2(n9373), .ZN(n11995) );
  NAND2_X1 U1638 ( .A1(n8562), .A2(n8587), .ZN(n12004) );
  NAND2_X1 U1639 ( .A1(n8562), .A2(n8586), .ZN(n12013) );
  NAND2_X1 U1640 ( .A1(n8562), .A2(n9403), .ZN(n12022) );
  NAND2_X1 U1641 ( .A1(n8562), .A2(n8584), .ZN(n12031) );
  NAND2_X1 U1642 ( .A1(n8562), .A2(n8583), .ZN(n12040) );
  NAND2_X1 U1643 ( .A1(n11876), .A2(n8582), .ZN(n12049) );
  NAND2_X1 U1644 ( .A1(n11876), .A2(n8581), .ZN(n12058) );
  NAND2_X1 U1645 ( .A1(n11876), .A2(n8580), .ZN(n12067) );
  NAND2_X1 U1646 ( .A1(n11876), .A2(n8579), .ZN(n12076) );
  NAND2_X1 U1647 ( .A1(n11876), .A2(n9473), .ZN(n12085) );
  NAND2_X1 U1648 ( .A1(n11876), .A2(n8577), .ZN(n12094) );
  NAND2_X1 U1649 ( .A1(n11876), .A2(n8576), .ZN(n12103) );
  NAND2_X1 U1650 ( .A1(n11876), .A2(n9503), .ZN(n12112) );
  NAND2_X1 U1651 ( .A1(n11876), .A2(n8574), .ZN(n12121) );
  NAND2_X1 U1652 ( .A1(n11876), .A2(n8573), .ZN(n12130) );
  NAND2_X1 U1653 ( .A1(n11876), .A2(n8572), .ZN(n12139) );
  NAND2_X1 U1654 ( .A1(n11876), .A2(n8571), .ZN(n12148) );
  NAND2_X1 U1655 ( .A1(n12165), .A2(n8603), .ZN(n12157) );
  NAND2_X1 U1656 ( .A1(n12165), .A2(n8601), .ZN(n12167) );
  NAND2_X1 U1657 ( .A1(n12165), .A2(n8600), .ZN(n12176) );
  NAND2_X1 U1658 ( .A1(n12165), .A2(n8599), .ZN(n12185) );
  NAND2_X1 U1659 ( .A1(n12165), .A2(n9273), .ZN(n12194) );
  NAND2_X1 U1660 ( .A1(n12165), .A2(n8597), .ZN(n12203) );
  NAND2_X1 U1661 ( .A1(n12165), .A2(n8596), .ZN(n12212) );
  NAND2_X1 U1662 ( .A1(n12165), .A2(n8595), .ZN(n12221) );
  NAND2_X1 U1663 ( .A1(n8561), .A2(n8594), .ZN(n12230) );
  NAND2_X1 U1664 ( .A1(n8561), .A2(n8593), .ZN(n12239) );
  NAND2_X1 U1665 ( .A1(n8561), .A2(n8592), .ZN(n12248) );
  NAND2_X1 U1666 ( .A1(n8561), .A2(n8591), .ZN(n12257) );
  NAND2_X1 U1667 ( .A1(n8561), .A2(n8590), .ZN(n12266) );
  NAND2_X1 U1668 ( .A1(n8561), .A2(n8589), .ZN(n12275) );
  NAND2_X1 U1669 ( .A1(n8561), .A2(n9373), .ZN(n12284) );
  NAND2_X1 U1670 ( .A1(n8561), .A2(n8587), .ZN(n12293) );
  NAND2_X1 U1671 ( .A1(n8561), .A2(n8586), .ZN(n12302) );
  NAND2_X1 U1672 ( .A1(n8561), .A2(n8585), .ZN(n12311) );
  NAND2_X1 U1673 ( .A1(n8561), .A2(n8584), .ZN(n12320) );
  NAND2_X1 U1674 ( .A1(n8561), .A2(n8583), .ZN(n12329) );
  NAND2_X1 U1675 ( .A1(n12165), .A2(n8582), .ZN(n12338) );
  NAND2_X1 U1676 ( .A1(n12165), .A2(n8581), .ZN(n12347) );
  NAND2_X1 U1677 ( .A1(n12165), .A2(n8580), .ZN(n12356) );
  NAND2_X1 U1678 ( .A1(n12165), .A2(n8579), .ZN(n12365) );
  NAND2_X1 U1679 ( .A1(n12165), .A2(n9473), .ZN(n12374) );
  NAND2_X1 U1680 ( .A1(n12165), .A2(n8577), .ZN(n12383) );
  NAND2_X1 U1681 ( .A1(n12165), .A2(n8576), .ZN(n12392) );
  NAND2_X1 U1682 ( .A1(n12165), .A2(n8575), .ZN(n12401) );
  NAND2_X1 U1683 ( .A1(n12165), .A2(n8574), .ZN(n12410) );
  NAND2_X1 U1684 ( .A1(n12165), .A2(n8573), .ZN(n12419) );
  NAND2_X1 U1685 ( .A1(n12165), .A2(n8572), .ZN(n12428) );
  NAND2_X1 U1686 ( .A1(n12165), .A2(n8571), .ZN(n12437) );
  NAND2_X1 U1687 ( .A1(n12454), .A2(n8603), .ZN(n12446) );
  NAND2_X1 U1688 ( .A1(n12454), .A2(n8601), .ZN(n12456) );
  NAND2_X1 U1689 ( .A1(n12454), .A2(n8600), .ZN(n12465) );
  NAND2_X1 U1690 ( .A1(n12454), .A2(n8599), .ZN(n12474) );
  NAND2_X1 U1691 ( .A1(n12454), .A2(n9273), .ZN(n12483) );
  NAND2_X1 U1692 ( .A1(n12454), .A2(n8597), .ZN(n12492) );
  NAND2_X1 U1693 ( .A1(n12454), .A2(n8596), .ZN(n12501) );
  NAND2_X1 U1694 ( .A1(n12454), .A2(n9303), .ZN(n12510) );
  NAND2_X1 U1695 ( .A1(n12454), .A2(n8594), .ZN(n12519) );
  NAND2_X1 U1696 ( .A1(n12454), .A2(n8593), .ZN(n12528) );
  NAND2_X1 U1697 ( .A1(n12454), .A2(n8592), .ZN(n12537) );
  NAND2_X1 U1698 ( .A1(n12454), .A2(n8591), .ZN(n12546) );
  NAND2_X1 U1699 ( .A1(n12454), .A2(n8590), .ZN(n12555) );
  NAND2_X1 U1700 ( .A1(n12454), .A2(n8589), .ZN(n12564) );
  NAND2_X1 U1701 ( .A1(n12454), .A2(n9373), .ZN(n12573) );
  NAND2_X1 U1702 ( .A1(n12454), .A2(n8587), .ZN(n12582) );
  NAND2_X1 U1703 ( .A1(n12454), .A2(n8586), .ZN(n12591) );
  NAND2_X1 U1704 ( .A1(n12454), .A2(n9403), .ZN(n12600) );
  NAND2_X1 U1705 ( .A1(n12454), .A2(n8584), .ZN(n12609) );
  NAND2_X1 U1706 ( .A1(n12454), .A2(n8583), .ZN(n12618) );
  NAND2_X1 U1707 ( .A1(n8560), .A2(n8582), .ZN(n12627) );
  NAND2_X1 U1708 ( .A1(n8560), .A2(n8581), .ZN(n12636) );
  NAND2_X1 U1709 ( .A1(n8560), .A2(n8580), .ZN(n12645) );
  NAND2_X1 U1710 ( .A1(n8560), .A2(n8579), .ZN(n12654) );
  NAND2_X1 U1711 ( .A1(n8560), .A2(n9473), .ZN(n12663) );
  NAND2_X1 U1712 ( .A1(n8560), .A2(n8577), .ZN(n12672) );
  NAND2_X1 U1713 ( .A1(n8560), .A2(n8576), .ZN(n12681) );
  NAND2_X1 U1714 ( .A1(n8560), .A2(n9503), .ZN(n12690) );
  NAND2_X1 U1715 ( .A1(n8560), .A2(n8574), .ZN(n12699) );
  NAND2_X1 U1716 ( .A1(n8560), .A2(n8573), .ZN(n12708) );
  NAND2_X1 U1717 ( .A1(n8560), .A2(n8572), .ZN(n12717) );
  NAND2_X1 U1718 ( .A1(n8560), .A2(n8571), .ZN(n12726) );
  NAND2_X1 U1719 ( .A1(n12743), .A2(n8603), .ZN(n12735) );
  NAND2_X1 U1720 ( .A1(n12743), .A2(n8601), .ZN(n12745) );
  NAND2_X1 U1721 ( .A1(n12743), .A2(n8600), .ZN(n12754) );
  NAND2_X1 U1722 ( .A1(n12743), .A2(n8599), .ZN(n12763) );
  NAND2_X1 U1723 ( .A1(n12743), .A2(n9273), .ZN(n12772) );
  NAND2_X1 U1724 ( .A1(n12743), .A2(n8597), .ZN(n12781) );
  NAND2_X1 U1725 ( .A1(n12743), .A2(n8596), .ZN(n12790) );
  NAND2_X1 U1726 ( .A1(n12743), .A2(n8595), .ZN(n12799) );
  NAND2_X1 U1727 ( .A1(n8559), .A2(n8594), .ZN(n12808) );
  NAND2_X1 U1728 ( .A1(n8559), .A2(n8593), .ZN(n12817) );
  NAND2_X1 U1729 ( .A1(n8559), .A2(n8592), .ZN(n12826) );
  NAND2_X1 U1730 ( .A1(n8559), .A2(n8591), .ZN(n12835) );
  NAND2_X1 U1731 ( .A1(n8559), .A2(n8590), .ZN(n12844) );
  NAND2_X1 U1732 ( .A1(n8559), .A2(n8589), .ZN(n12853) );
  NAND2_X1 U1733 ( .A1(n8559), .A2(n9373), .ZN(n12862) );
  NAND2_X1 U1734 ( .A1(n8559), .A2(n8587), .ZN(n12871) );
  NAND2_X1 U1735 ( .A1(n8559), .A2(n8586), .ZN(n12880) );
  NAND2_X1 U1736 ( .A1(n8559), .A2(n8585), .ZN(n12889) );
  NAND2_X1 U1737 ( .A1(n8559), .A2(n8584), .ZN(n12898) );
  NAND2_X1 U1738 ( .A1(n8559), .A2(n8583), .ZN(n12907) );
  NAND2_X1 U1739 ( .A1(n12743), .A2(n8582), .ZN(n12916) );
  NAND2_X1 U1740 ( .A1(n12743), .A2(n8581), .ZN(n12925) );
  NAND2_X1 U1741 ( .A1(n12743), .A2(n8580), .ZN(n12934) );
  NAND2_X1 U1742 ( .A1(n12743), .A2(n8579), .ZN(n12943) );
  NAND2_X1 U1743 ( .A1(n12743), .A2(n9473), .ZN(n12952) );
  NAND2_X1 U1744 ( .A1(n12743), .A2(n8577), .ZN(n12961) );
  NAND2_X1 U1745 ( .A1(n12743), .A2(n8576), .ZN(n12970) );
  NAND2_X1 U1746 ( .A1(n12743), .A2(n8575), .ZN(n12979) );
  NAND2_X1 U1747 ( .A1(n12743), .A2(n8574), .ZN(n12988) );
  NAND2_X1 U1748 ( .A1(n12743), .A2(n8573), .ZN(n12997) );
  NAND2_X1 U1749 ( .A1(n12743), .A2(n8572), .ZN(n13006) );
  NAND2_X1 U1750 ( .A1(n12743), .A2(n8571), .ZN(n13015) );
  NAND2_X1 U1751 ( .A1(n13032), .A2(n8603), .ZN(n13024) );
  NAND2_X1 U1752 ( .A1(n13032), .A2(n8601), .ZN(n13034) );
  NAND2_X1 U1753 ( .A1(n13032), .A2(n8600), .ZN(n13043) );
  NAND2_X1 U1754 ( .A1(n13032), .A2(n8599), .ZN(n13052) );
  NAND2_X1 U1755 ( .A1(n13032), .A2(n9273), .ZN(n13061) );
  NAND2_X1 U1756 ( .A1(n13032), .A2(n8597), .ZN(n13070) );
  NAND2_X1 U1757 ( .A1(n13032), .A2(n8596), .ZN(n13079) );
  NAND2_X1 U1758 ( .A1(n13032), .A2(n9303), .ZN(n13088) );
  NAND2_X1 U1759 ( .A1(n8558), .A2(n8594), .ZN(n13097) );
  NAND2_X1 U1760 ( .A1(n8558), .A2(n8593), .ZN(n13106) );
  NAND2_X1 U1761 ( .A1(n8558), .A2(n8592), .ZN(n13115) );
  NAND2_X1 U1762 ( .A1(n8558), .A2(n8591), .ZN(n13124) );
  NAND2_X1 U1763 ( .A1(n8558), .A2(n8590), .ZN(n13133) );
  NAND2_X1 U1764 ( .A1(n8558), .A2(n8589), .ZN(n13142) );
  NAND2_X1 U1765 ( .A1(n8558), .A2(n9373), .ZN(n13151) );
  NAND2_X1 U1766 ( .A1(n8558), .A2(n8587), .ZN(n13160) );
  NAND2_X1 U1767 ( .A1(n8558), .A2(n8586), .ZN(n13169) );
  NAND2_X1 U1768 ( .A1(n8558), .A2(n9403), .ZN(n13178) );
  NAND2_X1 U1769 ( .A1(n8558), .A2(n8584), .ZN(n13187) );
  NAND2_X1 U1770 ( .A1(n8558), .A2(n8583), .ZN(n13196) );
  NAND2_X1 U1771 ( .A1(n13032), .A2(n8582), .ZN(n13205) );
  NAND2_X1 U1772 ( .A1(n13032), .A2(n8581), .ZN(n13214) );
  NAND2_X1 U1773 ( .A1(n13032), .A2(n8580), .ZN(n13223) );
  NAND2_X1 U1774 ( .A1(n13032), .A2(n8579), .ZN(n13232) );
  NAND2_X1 U1775 ( .A1(n13032), .A2(n9473), .ZN(n13241) );
  NAND2_X1 U1776 ( .A1(n13032), .A2(n8577), .ZN(n13250) );
  NAND2_X1 U1777 ( .A1(n13032), .A2(n8576), .ZN(n13259) );
  NAND2_X1 U1778 ( .A1(n13032), .A2(n9503), .ZN(n13268) );
  NAND2_X1 U1779 ( .A1(n13032), .A2(n8574), .ZN(n13277) );
  NAND2_X1 U1780 ( .A1(n13032), .A2(n8573), .ZN(n13286) );
  NAND2_X1 U1781 ( .A1(n13032), .A2(n8572), .ZN(n13295) );
  NAND2_X1 U1782 ( .A1(n13032), .A2(n8571), .ZN(n13304) );
  NAND2_X1 U1783 ( .A1(n8557), .A2(n8603), .ZN(n13313) );
  NAND2_X1 U1784 ( .A1(n8557), .A2(n8601), .ZN(n13323) );
  NAND2_X1 U1785 ( .A1(n8557), .A2(n8600), .ZN(n13332) );
  NAND2_X1 U1786 ( .A1(n8557), .A2(n8599), .ZN(n13341) );
  NAND2_X1 U1787 ( .A1(n8557), .A2(n9273), .ZN(n13350) );
  NAND2_X1 U1788 ( .A1(n8557), .A2(n8597), .ZN(n13359) );
  NAND2_X1 U1789 ( .A1(n8557), .A2(n8596), .ZN(n13368) );
  NAND2_X1 U1790 ( .A1(n8557), .A2(n8595), .ZN(n13377) );
  NAND2_X1 U1791 ( .A1(n13321), .A2(n8594), .ZN(n13386) );
  NAND2_X1 U1792 ( .A1(n13321), .A2(n8593), .ZN(n13395) );
  NAND2_X1 U1793 ( .A1(n13321), .A2(n8592), .ZN(n13404) );
  NAND2_X1 U1794 ( .A1(n13321), .A2(n8591), .ZN(n13413) );
  NAND2_X1 U1795 ( .A1(n13321), .A2(n8590), .ZN(n13422) );
  NAND2_X1 U1796 ( .A1(n13321), .A2(n8589), .ZN(n13431) );
  NAND2_X1 U1797 ( .A1(n13321), .A2(n9373), .ZN(n13440) );
  NAND2_X1 U1798 ( .A1(n13321), .A2(n8587), .ZN(n13449) );
  NAND2_X1 U1799 ( .A1(n13321), .A2(n8586), .ZN(n13458) );
  NAND2_X1 U1800 ( .A1(n13321), .A2(n8585), .ZN(n13467) );
  NAND2_X1 U1801 ( .A1(n13321), .A2(n8584), .ZN(n13476) );
  NAND2_X1 U1802 ( .A1(n13321), .A2(n8583), .ZN(n13485) );
  NAND2_X1 U1803 ( .A1(n8557), .A2(n8582), .ZN(n13494) );
  NAND2_X1 U1804 ( .A1(n8557), .A2(n8581), .ZN(n13503) );
  NAND2_X1 U1805 ( .A1(n8557), .A2(n8580), .ZN(n13512) );
  NAND2_X1 U1806 ( .A1(n8557), .A2(n8579), .ZN(n13521) );
  NAND2_X1 U1807 ( .A1(n13321), .A2(n9473), .ZN(n13530) );
  NAND2_X1 U1808 ( .A1(n13321), .A2(n8577), .ZN(n13539) );
  NAND2_X1 U1809 ( .A1(n13321), .A2(n8576), .ZN(n13548) );
  NAND2_X1 U1810 ( .A1(n13321), .A2(n8575), .ZN(n13557) );
  NAND2_X1 U1811 ( .A1(n13321), .A2(n8574), .ZN(n13566) );
  NAND2_X1 U1812 ( .A1(n13321), .A2(n8573), .ZN(n13575) );
  NAND2_X1 U1813 ( .A1(n13321), .A2(n8572), .ZN(n13584) );
  NAND2_X1 U1814 ( .A1(n13321), .A2(n8571), .ZN(n13593) );
  NAND2_X1 U1815 ( .A1(n13610), .A2(n8603), .ZN(n13602) );
  NAND2_X1 U1816 ( .A1(n13610), .A2(n8601), .ZN(n13612) );
  NAND2_X1 U1817 ( .A1(n13610), .A2(n8600), .ZN(n13621) );
  NAND2_X1 U1818 ( .A1(n13610), .A2(n8599), .ZN(n13630) );
  NAND2_X1 U1819 ( .A1(n13610), .A2(n9273), .ZN(n13639) );
  NAND2_X1 U1820 ( .A1(n13610), .A2(n8597), .ZN(n13648) );
  NAND2_X1 U1821 ( .A1(n13610), .A2(n8596), .ZN(n13657) );
  NAND2_X1 U1822 ( .A1(n13610), .A2(n9303), .ZN(n13666) );
  NAND2_X1 U1823 ( .A1(n8556), .A2(n8594), .ZN(n13675) );
  NAND2_X1 U1824 ( .A1(n8556), .A2(n8593), .ZN(n13684) );
  NAND2_X1 U1825 ( .A1(n8556), .A2(n8592), .ZN(n13693) );
  NAND2_X1 U1826 ( .A1(n8556), .A2(n8591), .ZN(n13702) );
  NAND2_X1 U1827 ( .A1(n8556), .A2(n8590), .ZN(n13711) );
  NAND2_X1 U1828 ( .A1(n8556), .A2(n8589), .ZN(n13720) );
  NAND2_X1 U1829 ( .A1(n8556), .A2(n9373), .ZN(n13729) );
  NAND2_X1 U1830 ( .A1(n8556), .A2(n8587), .ZN(n13738) );
  NAND2_X1 U1831 ( .A1(n8556), .A2(n8586), .ZN(n13747) );
  NAND2_X1 U1832 ( .A1(n8556), .A2(n9403), .ZN(n13756) );
  NAND2_X1 U1833 ( .A1(n8556), .A2(n8584), .ZN(n13765) );
  NAND2_X1 U1834 ( .A1(n8556), .A2(n8583), .ZN(n13774) );
  NAND2_X1 U1835 ( .A1(n13610), .A2(n8582), .ZN(n13783) );
  NAND2_X1 U1836 ( .A1(n13610), .A2(n8581), .ZN(n13792) );
  NAND2_X1 U1837 ( .A1(n13610), .A2(n8580), .ZN(n13801) );
  NAND2_X1 U1838 ( .A1(n13610), .A2(n8579), .ZN(n13810) );
  NAND2_X1 U1839 ( .A1(n13610), .A2(n9473), .ZN(n13819) );
  NAND2_X1 U1840 ( .A1(n13610), .A2(n8577), .ZN(n13828) );
  NAND2_X1 U1841 ( .A1(n13610), .A2(n8576), .ZN(n13837) );
  NAND2_X1 U1842 ( .A1(n13610), .A2(n9503), .ZN(n13846) );
  NAND2_X1 U1843 ( .A1(n13610), .A2(n8574), .ZN(n13855) );
  NAND2_X1 U1844 ( .A1(n13610), .A2(n8573), .ZN(n13864) );
  NAND2_X1 U1845 ( .A1(n13610), .A2(n8572), .ZN(n13873) );
  NAND2_X1 U1846 ( .A1(n13610), .A2(n8571), .ZN(n13882) );
  NAND2_X1 U1847 ( .A1(n8555), .A2(n8603), .ZN(n13891) );
  NAND2_X1 U1848 ( .A1(n8555), .A2(n8601), .ZN(n13901) );
  NAND2_X1 U1849 ( .A1(n8555), .A2(n8600), .ZN(n13910) );
  NAND2_X1 U1850 ( .A1(n8555), .A2(n8599), .ZN(n13919) );
  NAND2_X1 U1851 ( .A1(n8555), .A2(n9273), .ZN(n13928) );
  NAND2_X1 U1852 ( .A1(n8555), .A2(n8597), .ZN(n13937) );
  NAND2_X1 U1853 ( .A1(n8555), .A2(n8596), .ZN(n13946) );
  NAND2_X1 U1854 ( .A1(n8555), .A2(n8595), .ZN(n13955) );
  NAND2_X1 U1855 ( .A1(n13899), .A2(n8594), .ZN(n13964) );
  NAND2_X1 U1856 ( .A1(n13899), .A2(n8593), .ZN(n13973) );
  NAND2_X1 U1857 ( .A1(n13899), .A2(n8592), .ZN(n13982) );
  NAND2_X1 U1858 ( .A1(n13899), .A2(n8591), .ZN(n13991) );
  NAND2_X1 U1859 ( .A1(n13899), .A2(n8590), .ZN(n14000) );
  NAND2_X1 U1860 ( .A1(n13899), .A2(n8589), .ZN(n14009) );
  NAND2_X1 U1861 ( .A1(n13899), .A2(n9373), .ZN(n14018) );
  NAND2_X1 U1862 ( .A1(n13899), .A2(n8587), .ZN(n14027) );
  NAND2_X1 U1863 ( .A1(n13899), .A2(n8586), .ZN(n14036) );
  NAND2_X1 U1864 ( .A1(n13899), .A2(n8585), .ZN(n14045) );
  NAND2_X1 U1865 ( .A1(n13899), .A2(n8584), .ZN(n14054) );
  NAND2_X1 U1866 ( .A1(n13899), .A2(n8583), .ZN(n14063) );
  NAND2_X1 U1867 ( .A1(n8555), .A2(n8582), .ZN(n14072) );
  NAND2_X1 U1868 ( .A1(n8555), .A2(n8581), .ZN(n14081) );
  NAND2_X1 U1869 ( .A1(n8555), .A2(n8580), .ZN(n14090) );
  NAND2_X1 U1870 ( .A1(n8555), .A2(n8579), .ZN(n14099) );
  NAND2_X1 U1871 ( .A1(n13899), .A2(n9473), .ZN(n14108) );
  NAND2_X1 U1872 ( .A1(n13899), .A2(n8577), .ZN(n14117) );
  NAND2_X1 U1873 ( .A1(n13899), .A2(n8576), .ZN(n14126) );
  NAND2_X1 U1874 ( .A1(n13899), .A2(n8575), .ZN(n14135) );
  NAND2_X1 U1875 ( .A1(n13899), .A2(n8574), .ZN(n14144) );
  NAND2_X1 U1876 ( .A1(n13899), .A2(n8573), .ZN(n14153) );
  NAND2_X1 U1877 ( .A1(n13899), .A2(n8572), .ZN(n14162) );
  NAND2_X1 U1878 ( .A1(n13899), .A2(n8571), .ZN(n14171) );
  NAND2_X1 U1879 ( .A1(n14189), .A2(n8603), .ZN(n14181) );
  NAND2_X1 U1880 ( .A1(n14189), .A2(n8601), .ZN(n14191) );
  NAND2_X1 U1881 ( .A1(n14189), .A2(n8600), .ZN(n14200) );
  NAND2_X1 U1882 ( .A1(n14189), .A2(n8599), .ZN(n14209) );
  NAND2_X1 U1883 ( .A1(n14189), .A2(n9273), .ZN(n14218) );
  NAND2_X1 U1884 ( .A1(n14189), .A2(n8597), .ZN(n14227) );
  NAND2_X1 U1885 ( .A1(n14189), .A2(n8596), .ZN(n14236) );
  NAND2_X1 U1886 ( .A1(n14189), .A2(n9303), .ZN(n14245) );
  NAND2_X1 U1887 ( .A1(n8554), .A2(n8594), .ZN(n14254) );
  NAND2_X1 U1888 ( .A1(n8554), .A2(n8593), .ZN(n14263) );
  NAND2_X1 U1889 ( .A1(n8554), .A2(n8592), .ZN(n14272) );
  NAND2_X1 U1890 ( .A1(n8554), .A2(n8591), .ZN(n14281) );
  NAND2_X1 U1891 ( .A1(n8554), .A2(n8590), .ZN(n14290) );
  NAND2_X1 U1892 ( .A1(n8554), .A2(n8589), .ZN(n14299) );
  NAND2_X1 U1893 ( .A1(n8554), .A2(n9373), .ZN(n14308) );
  NAND2_X1 U1894 ( .A1(n8554), .A2(n8587), .ZN(n14317) );
  NAND2_X1 U1895 ( .A1(n8554), .A2(n8586), .ZN(n14326) );
  NAND2_X1 U1896 ( .A1(n8554), .A2(n9403), .ZN(n14335) );
  NAND2_X1 U1897 ( .A1(n8554), .A2(n8584), .ZN(n14344) );
  NAND2_X1 U1898 ( .A1(n8554), .A2(n8583), .ZN(n14353) );
  NAND2_X1 U1899 ( .A1(n14189), .A2(n8582), .ZN(n14362) );
  NAND2_X1 U1900 ( .A1(n14189), .A2(n8581), .ZN(n14371) );
  NAND2_X1 U1901 ( .A1(n14189), .A2(n8580), .ZN(n14380) );
  NAND2_X1 U1902 ( .A1(n14189), .A2(n8579), .ZN(n14389) );
  NAND2_X1 U1903 ( .A1(n14189), .A2(n9473), .ZN(n14398) );
  NAND2_X1 U1904 ( .A1(n14189), .A2(n8577), .ZN(n14407) );
  NAND2_X1 U1905 ( .A1(n14189), .A2(n8576), .ZN(n14416) );
  NAND2_X1 U1906 ( .A1(n14189), .A2(n9503), .ZN(n14425) );
  NAND2_X1 U1907 ( .A1(n14189), .A2(n8574), .ZN(n14434) );
  NAND2_X1 U1908 ( .A1(n14189), .A2(n8573), .ZN(n14443) );
  NAND2_X1 U1909 ( .A1(n14189), .A2(n8572), .ZN(n14452) );
  NAND2_X1 U1910 ( .A1(n14189), .A2(n8571), .ZN(n14461) );
  NAND2_X1 U1911 ( .A1(n14478), .A2(n8603), .ZN(n14470) );
  NAND2_X1 U1912 ( .A1(n14478), .A2(n8601), .ZN(n14480) );
  NAND2_X1 U1913 ( .A1(n14478), .A2(n8600), .ZN(n14489) );
  NAND2_X1 U1914 ( .A1(n14478), .A2(n8599), .ZN(n14498) );
  NAND2_X1 U1915 ( .A1(n14478), .A2(n9273), .ZN(n14507) );
  NAND2_X1 U1916 ( .A1(n14478), .A2(n8597), .ZN(n14516) );
  NAND2_X1 U1917 ( .A1(n14478), .A2(n8596), .ZN(n14525) );
  NAND2_X1 U1918 ( .A1(n14478), .A2(n8595), .ZN(n14534) );
  NAND2_X1 U1919 ( .A1(n8553), .A2(n8594), .ZN(n14543) );
  NAND2_X1 U1920 ( .A1(n8553), .A2(n8593), .ZN(n14552) );
  NAND2_X1 U1921 ( .A1(n8553), .A2(n8592), .ZN(n14561) );
  NAND2_X1 U1922 ( .A1(n8553), .A2(n8591), .ZN(n14570) );
  NAND2_X1 U1923 ( .A1(n8553), .A2(n8590), .ZN(n14579) );
  NAND2_X1 U1924 ( .A1(n8553), .A2(n8589), .ZN(n14588) );
  NAND2_X1 U1925 ( .A1(n8553), .A2(n9373), .ZN(n14597) );
  NAND2_X1 U1926 ( .A1(n8553), .A2(n8587), .ZN(n14606) );
  NAND2_X1 U1927 ( .A1(n8553), .A2(n8586), .ZN(n14615) );
  NAND2_X1 U1928 ( .A1(n8553), .A2(n8585), .ZN(n14624) );
  NAND2_X1 U1929 ( .A1(n8553), .A2(n8584), .ZN(n14633) );
  NAND2_X1 U1930 ( .A1(n8553), .A2(n8583), .ZN(n14642) );
  NAND2_X1 U1931 ( .A1(n14478), .A2(n8582), .ZN(n14651) );
  NAND2_X1 U1932 ( .A1(n14478), .A2(n8581), .ZN(n14660) );
  NAND2_X1 U1933 ( .A1(n14478), .A2(n8580), .ZN(n14669) );
  NAND2_X1 U1934 ( .A1(n14478), .A2(n8579), .ZN(n14678) );
  NAND2_X1 U1935 ( .A1(n14478), .A2(n9473), .ZN(n14687) );
  NAND2_X1 U1936 ( .A1(n14478), .A2(n8577), .ZN(n14696) );
  NAND2_X1 U1937 ( .A1(n14478), .A2(n8576), .ZN(n14705) );
  NAND2_X1 U1938 ( .A1(n14478), .A2(n8575), .ZN(n14714) );
  NAND2_X1 U1939 ( .A1(n14478), .A2(n8574), .ZN(n14723) );
  NAND2_X1 U1940 ( .A1(n14478), .A2(n8573), .ZN(n14732) );
  NAND2_X1 U1941 ( .A1(n14478), .A2(n8572), .ZN(n14741) );
  NAND2_X1 U1942 ( .A1(n14478), .A2(n8571), .ZN(n14750) );
  NAND2_X1 U1943 ( .A1(n14767), .A2(n8603), .ZN(n14759) );
  NAND2_X1 U1944 ( .A1(n14767), .A2(n8601), .ZN(n14769) );
  NAND2_X1 U1945 ( .A1(n14767), .A2(n8600), .ZN(n14778) );
  NAND2_X1 U1946 ( .A1(n14767), .A2(n8599), .ZN(n14787) );
  NAND2_X1 U1947 ( .A1(n14767), .A2(n9273), .ZN(n14796) );
  NAND2_X1 U1948 ( .A1(n14767), .A2(n8597), .ZN(n14805) );
  NAND2_X1 U1949 ( .A1(n14767), .A2(n8596), .ZN(n14814) );
  NAND2_X1 U1950 ( .A1(n14767), .A2(n9303), .ZN(n14823) );
  NAND2_X1 U1951 ( .A1(n8552), .A2(n8594), .ZN(n14832) );
  NAND2_X1 U1952 ( .A1(n8552), .A2(n8593), .ZN(n14841) );
  NAND2_X1 U1953 ( .A1(n8552), .A2(n8592), .ZN(n14850) );
  NAND2_X1 U1954 ( .A1(n8552), .A2(n8591), .ZN(n14859) );
  NAND2_X1 U1955 ( .A1(n8552), .A2(n8590), .ZN(n14868) );
  NAND2_X1 U1956 ( .A1(n8552), .A2(n8589), .ZN(n14877) );
  NAND2_X1 U1957 ( .A1(n8552), .A2(n9373), .ZN(n14886) );
  NAND2_X1 U1958 ( .A1(n8552), .A2(n8587), .ZN(n14895) );
  NAND2_X1 U1959 ( .A1(n8552), .A2(n8586), .ZN(n14904) );
  NAND2_X1 U1960 ( .A1(n8552), .A2(n9403), .ZN(n14913) );
  NAND2_X1 U1961 ( .A1(n8552), .A2(n8584), .ZN(n14922) );
  NAND2_X1 U1962 ( .A1(n8552), .A2(n8583), .ZN(n14931) );
  NAND2_X1 U1963 ( .A1(n14767), .A2(n8582), .ZN(n14940) );
  NAND2_X1 U1964 ( .A1(n14767), .A2(n8581), .ZN(n14949) );
  NAND2_X1 U1965 ( .A1(n14767), .A2(n8580), .ZN(n14958) );
  NAND2_X1 U1966 ( .A1(n14767), .A2(n8579), .ZN(n14967) );
  NAND2_X1 U1967 ( .A1(n14767), .A2(n9473), .ZN(n14976) );
  NAND2_X1 U1968 ( .A1(n14767), .A2(n8577), .ZN(n14985) );
  NAND2_X1 U1969 ( .A1(n14767), .A2(n8576), .ZN(n14994) );
  NAND2_X1 U1970 ( .A1(n14767), .A2(n9503), .ZN(n15003) );
  NAND2_X1 U1971 ( .A1(n14767), .A2(n8574), .ZN(n15012) );
  NAND2_X1 U1972 ( .A1(n14767), .A2(n8573), .ZN(n15021) );
  NAND2_X1 U1973 ( .A1(n14767), .A2(n8572), .ZN(n15030) );
  NAND2_X1 U1974 ( .A1(n14767), .A2(n8571), .ZN(n15039) );
  NAND2_X1 U1975 ( .A1(n15056), .A2(n9232), .ZN(n15048) );
  NAND2_X1 U1976 ( .A1(n15056), .A2(n9243), .ZN(n15058) );
  NAND2_X1 U1977 ( .A1(n15056), .A2(n9253), .ZN(n15067) );
  NAND2_X1 U1978 ( .A1(n15056), .A2(n9263), .ZN(n15076) );
  NAND2_X1 U1979 ( .A1(n15056), .A2(n8598), .ZN(n15085) );
  NAND2_X1 U1980 ( .A1(n15056), .A2(n9283), .ZN(n15094) );
  NAND2_X1 U1981 ( .A1(n15056), .A2(n9293), .ZN(n15103) );
  NAND2_X1 U1982 ( .A1(n15056), .A2(n9303), .ZN(n15112) );
  NAND2_X1 U1983 ( .A1(n8551), .A2(n9313), .ZN(n15121) );
  NAND2_X1 U1984 ( .A1(n8551), .A2(n9323), .ZN(n15130) );
  NAND2_X1 U1985 ( .A1(n8551), .A2(n9333), .ZN(n15139) );
  NAND2_X1 U1986 ( .A1(n8551), .A2(n9343), .ZN(n15148) );
  NAND2_X1 U1987 ( .A1(n8551), .A2(n9353), .ZN(n15157) );
  NAND2_X1 U1988 ( .A1(n8551), .A2(n9363), .ZN(n15166) );
  NAND2_X1 U1989 ( .A1(n8551), .A2(n8588), .ZN(n15175) );
  NAND2_X1 U1990 ( .A1(n8551), .A2(n9383), .ZN(n15184) );
  NAND2_X1 U1991 ( .A1(n8551), .A2(n9393), .ZN(n15193) );
  NAND2_X1 U1992 ( .A1(n8551), .A2(n9403), .ZN(n15202) );
  NAND2_X1 U1993 ( .A1(n8551), .A2(n9413), .ZN(n15211) );
  NAND2_X1 U1994 ( .A1(n8551), .A2(n9423), .ZN(n15220) );
  NAND2_X1 U1995 ( .A1(n15056), .A2(n9433), .ZN(n15229) );
  NAND2_X1 U1996 ( .A1(n15056), .A2(n9443), .ZN(n15238) );
  NAND2_X1 U1997 ( .A1(n15056), .A2(n9453), .ZN(n15247) );
  NAND2_X1 U1998 ( .A1(n15056), .A2(n9463), .ZN(n15256) );
  NAND2_X1 U1999 ( .A1(n15056), .A2(n8578), .ZN(n15265) );
  NAND2_X1 U2000 ( .A1(n15056), .A2(n9483), .ZN(n15274) );
  NAND2_X1 U2001 ( .A1(n15056), .A2(n9493), .ZN(n15283) );
  NAND2_X1 U2002 ( .A1(n15056), .A2(n9503), .ZN(n15292) );
  NAND2_X1 U2003 ( .A1(n15056), .A2(n9513), .ZN(n15301) );
  NAND2_X1 U2004 ( .A1(n15056), .A2(n9523), .ZN(n15310) );
  NAND2_X1 U2005 ( .A1(n15056), .A2(n9533), .ZN(n15319) );
  NAND2_X1 U2006 ( .A1(n15056), .A2(n9543), .ZN(n15328) );
  NAND2_X1 U2007 ( .A1(n15345), .A2(n9232), .ZN(n15337) );
  NAND2_X1 U2008 ( .A1(n15345), .A2(n9243), .ZN(n15347) );
  NAND2_X1 U2009 ( .A1(n15345), .A2(n9253), .ZN(n15356) );
  NAND2_X1 U2010 ( .A1(n15345), .A2(n9263), .ZN(n15365) );
  NAND2_X1 U2011 ( .A1(n15345), .A2(n8598), .ZN(n15374) );
  NAND2_X1 U2012 ( .A1(n15345), .A2(n9283), .ZN(n15383) );
  NAND2_X1 U2013 ( .A1(n15345), .A2(n9293), .ZN(n15392) );
  NAND2_X1 U2014 ( .A1(n15345), .A2(n9303), .ZN(n15401) );
  NAND2_X1 U2015 ( .A1(n8550), .A2(n9313), .ZN(n15410) );
  NAND2_X1 U2016 ( .A1(n8550), .A2(n9323), .ZN(n15419) );
  NAND2_X1 U2017 ( .A1(n8550), .A2(n9333), .ZN(n15428) );
  NAND2_X1 U2018 ( .A1(n8550), .A2(n9343), .ZN(n15437) );
  NAND2_X1 U2019 ( .A1(n8550), .A2(n9353), .ZN(n15446) );
  NAND2_X1 U2020 ( .A1(n8550), .A2(n9363), .ZN(n15455) );
  NAND2_X1 U2021 ( .A1(n8550), .A2(n8588), .ZN(n15464) );
  NAND2_X1 U2022 ( .A1(n8550), .A2(n9383), .ZN(n15473) );
  NAND2_X1 U2023 ( .A1(n8550), .A2(n9393), .ZN(n15482) );
  NAND2_X1 U2024 ( .A1(n8550), .A2(n9403), .ZN(n15491) );
  NAND2_X1 U2025 ( .A1(n8550), .A2(n9413), .ZN(n15500) );
  NAND2_X1 U2026 ( .A1(n8550), .A2(n9423), .ZN(n15509) );
  NAND2_X1 U2027 ( .A1(n15345), .A2(n9433), .ZN(n15518) );
  NAND2_X1 U2028 ( .A1(n15345), .A2(n9443), .ZN(n15527) );
  NAND2_X1 U2029 ( .A1(n15345), .A2(n9453), .ZN(n15536) );
  NAND2_X1 U2030 ( .A1(n15345), .A2(n9463), .ZN(n15545) );
  NAND2_X1 U2031 ( .A1(n15345), .A2(n8578), .ZN(n15554) );
  NAND2_X1 U2032 ( .A1(n15345), .A2(n9483), .ZN(n15563) );
  NAND2_X1 U2033 ( .A1(n15345), .A2(n9493), .ZN(n15572) );
  NAND2_X1 U2034 ( .A1(n15345), .A2(n9503), .ZN(n15581) );
  NAND2_X1 U2035 ( .A1(n15345), .A2(n9513), .ZN(n15590) );
  NAND2_X1 U2036 ( .A1(n15345), .A2(n9523), .ZN(n15599) );
  NAND2_X1 U2037 ( .A1(n15345), .A2(n9533), .ZN(n15608) );
  NAND2_X1 U2038 ( .A1(n15345), .A2(n9543), .ZN(n15617) );
  NAND2_X1 U2039 ( .A1(n15634), .A2(n9232), .ZN(n15626) );
  NAND2_X1 U2040 ( .A1(n15634), .A2(n9243), .ZN(n15636) );
  NAND2_X1 U2041 ( .A1(n15634), .A2(n9253), .ZN(n15645) );
  NAND2_X1 U2042 ( .A1(n15634), .A2(n9263), .ZN(n15654) );
  NAND2_X1 U2043 ( .A1(n15634), .A2(n8598), .ZN(n15663) );
  NAND2_X1 U2044 ( .A1(n15634), .A2(n9283), .ZN(n15672) );
  NAND2_X1 U2045 ( .A1(n15634), .A2(n9293), .ZN(n15681) );
  NAND2_X1 U2046 ( .A1(n15634), .A2(n9303), .ZN(n15690) );
  NAND2_X1 U2047 ( .A1(n8549), .A2(n9313), .ZN(n15699) );
  NAND2_X1 U2048 ( .A1(n8549), .A2(n9323), .ZN(n15708) );
  NAND2_X1 U2049 ( .A1(n8549), .A2(n9333), .ZN(n15717) );
  NAND2_X1 U2050 ( .A1(n8549), .A2(n9343), .ZN(n15726) );
  NAND2_X1 U2051 ( .A1(n8549), .A2(n9353), .ZN(n15735) );
  NAND2_X1 U2052 ( .A1(n8549), .A2(n9363), .ZN(n15744) );
  NAND2_X1 U2053 ( .A1(n8549), .A2(n8588), .ZN(n15753) );
  NAND2_X1 U2054 ( .A1(n8549), .A2(n9383), .ZN(n15762) );
  NAND2_X1 U2055 ( .A1(n8549), .A2(n9393), .ZN(n15771) );
  NAND2_X1 U2056 ( .A1(n8549), .A2(n9403), .ZN(n15780) );
  NAND2_X1 U2057 ( .A1(n8549), .A2(n9413), .ZN(n15789) );
  NAND2_X1 U2058 ( .A1(n8549), .A2(n9423), .ZN(n15798) );
  NAND2_X1 U2059 ( .A1(n15634), .A2(n9433), .ZN(n15807) );
  NAND2_X1 U2060 ( .A1(n15634), .A2(n9443), .ZN(n15816) );
  NAND2_X1 U2061 ( .A1(n15634), .A2(n9453), .ZN(n15825) );
  NAND2_X1 U2062 ( .A1(n15634), .A2(n9463), .ZN(n15834) );
  NAND2_X1 U2063 ( .A1(n15634), .A2(n8578), .ZN(n15843) );
  NAND2_X1 U2064 ( .A1(n15634), .A2(n9483), .ZN(n15852) );
  NAND2_X1 U2065 ( .A1(n15634), .A2(n9493), .ZN(n15861) );
  NAND2_X1 U2066 ( .A1(n15634), .A2(n9503), .ZN(n15870) );
  NAND2_X1 U2067 ( .A1(n15634), .A2(n9513), .ZN(n15879) );
  NAND2_X1 U2068 ( .A1(n15634), .A2(n9523), .ZN(n15888) );
  NAND2_X1 U2069 ( .A1(n15634), .A2(n9533), .ZN(n15897) );
  NAND2_X1 U2070 ( .A1(n15634), .A2(n9543), .ZN(n15906) );
  NAND2_X1 U2071 ( .A1(n15923), .A2(n9232), .ZN(n15915) );
  NAND2_X1 U2072 ( .A1(n15923), .A2(n9243), .ZN(n15925) );
  NAND2_X1 U2073 ( .A1(n15923), .A2(n9253), .ZN(n15934) );
  NAND2_X1 U2074 ( .A1(n15923), .A2(n9263), .ZN(n15943) );
  NAND2_X1 U2075 ( .A1(n15923), .A2(n8598), .ZN(n15952) );
  NAND2_X1 U2076 ( .A1(n15923), .A2(n9283), .ZN(n15961) );
  NAND2_X1 U2077 ( .A1(n15923), .A2(n9293), .ZN(n15970) );
  NAND2_X1 U2078 ( .A1(n15923), .A2(n9303), .ZN(n15979) );
  NAND2_X1 U2079 ( .A1(n15923), .A2(n9313), .ZN(n15988) );
  NAND2_X1 U2080 ( .A1(n15923), .A2(n9323), .ZN(n15997) );
  NAND2_X1 U2081 ( .A1(n15923), .A2(n9333), .ZN(n16006) );
  NAND2_X1 U2082 ( .A1(n15923), .A2(n9343), .ZN(n16015) );
  NAND2_X1 U2083 ( .A1(n15923), .A2(n9353), .ZN(n16024) );
  NAND2_X1 U2084 ( .A1(n15923), .A2(n9363), .ZN(n16033) );
  NAND2_X1 U2085 ( .A1(n15923), .A2(n8588), .ZN(n16042) );
  NAND2_X1 U2086 ( .A1(n15923), .A2(n9383), .ZN(n16051) );
  NAND2_X1 U2087 ( .A1(n15923), .A2(n9393), .ZN(n16060) );
  NAND2_X1 U2088 ( .A1(n15923), .A2(n9403), .ZN(n16069) );
  NAND2_X1 U2089 ( .A1(n15923), .A2(n9413), .ZN(n16078) );
  NAND2_X1 U2090 ( .A1(n15923), .A2(n9423), .ZN(n16087) );
  NAND2_X1 U2091 ( .A1(n8548), .A2(n9433), .ZN(n16096) );
  NAND2_X1 U2092 ( .A1(n8548), .A2(n9443), .ZN(n16105) );
  NAND2_X1 U2093 ( .A1(n8548), .A2(n9453), .ZN(n16114) );
  NAND2_X1 U2094 ( .A1(n8548), .A2(n9463), .ZN(n16123) );
  NAND2_X1 U2095 ( .A1(n8548), .A2(n8578), .ZN(n16132) );
  NAND2_X1 U2096 ( .A1(n8548), .A2(n9483), .ZN(n16141) );
  NAND2_X1 U2097 ( .A1(n8548), .A2(n9493), .ZN(n16150) );
  NAND2_X1 U2098 ( .A1(n8548), .A2(n9503), .ZN(n16159) );
  NAND2_X1 U2099 ( .A1(n8548), .A2(n9513), .ZN(n16168) );
  NAND2_X1 U2100 ( .A1(n8548), .A2(n9523), .ZN(n16177) );
  NAND2_X1 U2101 ( .A1(n8548), .A2(n9533), .ZN(n16186) );
  NAND2_X1 U2102 ( .A1(n8548), .A2(n9543), .ZN(n16195) );
  NAND2_X1 U2103 ( .A1(n16212), .A2(n8603), .ZN(n16204) );
  NAND2_X1 U2104 ( .A1(n16212), .A2(n8601), .ZN(n16214) );
  NAND2_X1 U2105 ( .A1(n16212), .A2(n8600), .ZN(n16223) );
  NAND2_X1 U2106 ( .A1(n16212), .A2(n8599), .ZN(n16232) );
  NAND2_X1 U2107 ( .A1(n16212), .A2(n8598), .ZN(n16241) );
  NAND2_X1 U2108 ( .A1(n16212), .A2(n8597), .ZN(n16250) );
  NAND2_X1 U2109 ( .A1(n16212), .A2(n8596), .ZN(n16259) );
  NAND2_X1 U2110 ( .A1(n16212), .A2(n9303), .ZN(n16268) );
  NAND2_X1 U2111 ( .A1(n8547), .A2(n8594), .ZN(n16277) );
  NAND2_X1 U2112 ( .A1(n8547), .A2(n8593), .ZN(n16286) );
  NAND2_X1 U2113 ( .A1(n8547), .A2(n8592), .ZN(n16295) );
  NAND2_X1 U2114 ( .A1(n8547), .A2(n8591), .ZN(n16304) );
  NAND2_X1 U2115 ( .A1(n8547), .A2(n8590), .ZN(n16313) );
  NAND2_X1 U2116 ( .A1(n8547), .A2(n8589), .ZN(n16322) );
  NAND2_X1 U2117 ( .A1(n8547), .A2(n8588), .ZN(n16331) );
  NAND2_X1 U2118 ( .A1(n8547), .A2(n8587), .ZN(n16340) );
  NAND2_X1 U2119 ( .A1(n8547), .A2(n8586), .ZN(n16349) );
  NAND2_X1 U2120 ( .A1(n8547), .A2(n9403), .ZN(n16358) );
  NAND2_X1 U2121 ( .A1(n8547), .A2(n8584), .ZN(n16367) );
  NAND2_X1 U2122 ( .A1(n8547), .A2(n8583), .ZN(n16376) );
  NAND2_X1 U2123 ( .A1(n16212), .A2(n8582), .ZN(n16385) );
  NAND2_X1 U2124 ( .A1(n16212), .A2(n8581), .ZN(n16394) );
  NAND2_X1 U2125 ( .A1(n16212), .A2(n8580), .ZN(n16403) );
  NAND2_X1 U2126 ( .A1(n16212), .A2(n8579), .ZN(n16412) );
  NAND2_X1 U2127 ( .A1(n16212), .A2(n8578), .ZN(n16421) );
  NAND2_X1 U2128 ( .A1(n16212), .A2(n8577), .ZN(n16430) );
  NAND2_X1 U2129 ( .A1(n16212), .A2(n8576), .ZN(n16439) );
  NAND2_X1 U2130 ( .A1(n16212), .A2(n9503), .ZN(n16448) );
  NAND2_X1 U2131 ( .A1(n16212), .A2(n8574), .ZN(n16457) );
  NAND2_X1 U2132 ( .A1(n16212), .A2(n8573), .ZN(n16466) );
  NAND2_X1 U2133 ( .A1(n16212), .A2(n8572), .ZN(n16475) );
  NAND2_X1 U2134 ( .A1(n16212), .A2(n8571), .ZN(n16484) );
  NAND2_X1 U2135 ( .A1(n16502), .A2(n9232), .ZN(n16494) );
  NAND2_X1 U2136 ( .A1(n16502), .A2(n9243), .ZN(n16504) );
  NAND2_X1 U2137 ( .A1(n16502), .A2(n9253), .ZN(n16513) );
  NAND2_X1 U2138 ( .A1(n16502), .A2(n9263), .ZN(n16522) );
  NAND2_X1 U2139 ( .A1(n16502), .A2(n8598), .ZN(n16531) );
  NAND2_X1 U2140 ( .A1(n16502), .A2(n9283), .ZN(n16540) );
  NAND2_X1 U2141 ( .A1(n16502), .A2(n9293), .ZN(n16549) );
  NAND2_X1 U2142 ( .A1(n16502), .A2(n9303), .ZN(n16558) );
  NAND2_X1 U2143 ( .A1(n8546), .A2(n9313), .ZN(n16567) );
  NAND2_X1 U2144 ( .A1(n8546), .A2(n9323), .ZN(n16576) );
  NAND2_X1 U2145 ( .A1(n8546), .A2(n9333), .ZN(n16585) );
  NAND2_X1 U2146 ( .A1(n8546), .A2(n9343), .ZN(n16594) );
  NAND2_X1 U2147 ( .A1(n8546), .A2(n9353), .ZN(n16603) );
  NAND2_X1 U2148 ( .A1(n8546), .A2(n9363), .ZN(n16612) );
  NAND2_X1 U2149 ( .A1(n8546), .A2(n8588), .ZN(n16621) );
  NAND2_X1 U2150 ( .A1(n8546), .A2(n9383), .ZN(n16630) );
  NAND2_X1 U2151 ( .A1(n8546), .A2(n9393), .ZN(n16639) );
  NAND2_X1 U2152 ( .A1(n8546), .A2(n9403), .ZN(n16648) );
  NAND2_X1 U2153 ( .A1(n8546), .A2(n9413), .ZN(n16657) );
  NAND2_X1 U2154 ( .A1(n8546), .A2(n9423), .ZN(n16666) );
  NAND2_X1 U2155 ( .A1(n16502), .A2(n9433), .ZN(n16675) );
  NAND2_X1 U2156 ( .A1(n16502), .A2(n9443), .ZN(n16684) );
  NAND2_X1 U2157 ( .A1(n16502), .A2(n9453), .ZN(n16693) );
  NAND2_X1 U2158 ( .A1(n16502), .A2(n9463), .ZN(n16702) );
  NAND2_X1 U2159 ( .A1(n16502), .A2(n8578), .ZN(n16711) );
  NAND2_X1 U2160 ( .A1(n16502), .A2(n9483), .ZN(n16720) );
  NAND2_X1 U2161 ( .A1(n16502), .A2(n9493), .ZN(n16729) );
  NAND2_X1 U2162 ( .A1(n16502), .A2(n9503), .ZN(n16738) );
  NAND2_X1 U2163 ( .A1(n16502), .A2(n9513), .ZN(n16747) );
  NAND2_X1 U2164 ( .A1(n16502), .A2(n9523), .ZN(n16756) );
  NAND2_X1 U2165 ( .A1(n16502), .A2(n9533), .ZN(n16765) );
  NAND2_X1 U2166 ( .A1(n16502), .A2(n9543), .ZN(n16774) );
  NAND2_X1 U2167 ( .A1(n16791), .A2(n8603), .ZN(n16783) );
  NAND2_X1 U2168 ( .A1(n16791), .A2(n8601), .ZN(n16793) );
  NAND2_X1 U2169 ( .A1(n16791), .A2(n8600), .ZN(n16802) );
  NAND2_X1 U2170 ( .A1(n16791), .A2(n8599), .ZN(n16811) );
  NAND2_X1 U2171 ( .A1(n16791), .A2(n8598), .ZN(n16820) );
  NAND2_X1 U2172 ( .A1(n16791), .A2(n8597), .ZN(n16829) );
  NAND2_X1 U2173 ( .A1(n16791), .A2(n8596), .ZN(n16838) );
  NAND2_X1 U2174 ( .A1(n16791), .A2(n9303), .ZN(n16847) );
  NAND2_X1 U2175 ( .A1(n8545), .A2(n8594), .ZN(n16856) );
  NAND2_X1 U2176 ( .A1(n8545), .A2(n8593), .ZN(n16865) );
  NAND2_X1 U2177 ( .A1(n8545), .A2(n8592), .ZN(n16874) );
  NAND2_X1 U2178 ( .A1(n8545), .A2(n8591), .ZN(n16883) );
  NAND2_X1 U2179 ( .A1(n8545), .A2(n8590), .ZN(n16892) );
  NAND2_X1 U2180 ( .A1(n8545), .A2(n8589), .ZN(n16901) );
  NAND2_X1 U2181 ( .A1(n8545), .A2(n8588), .ZN(n16910) );
  NAND2_X1 U2182 ( .A1(n8545), .A2(n8587), .ZN(n16919) );
  NAND2_X1 U2183 ( .A1(n8545), .A2(n8586), .ZN(n16928) );
  NAND2_X1 U2184 ( .A1(n8545), .A2(n9403), .ZN(n16937) );
  NAND2_X1 U2185 ( .A1(n8545), .A2(n8584), .ZN(n16946) );
  NAND2_X1 U2186 ( .A1(n8545), .A2(n8583), .ZN(n16955) );
  NAND2_X1 U2187 ( .A1(n16791), .A2(n8582), .ZN(n16964) );
  NAND2_X1 U2188 ( .A1(n16791), .A2(n8581), .ZN(n16973) );
  NAND2_X1 U2189 ( .A1(n16791), .A2(n8580), .ZN(n16982) );
  NAND2_X1 U2190 ( .A1(n16791), .A2(n8579), .ZN(n16991) );
  NAND2_X1 U2191 ( .A1(n16791), .A2(n8578), .ZN(n17000) );
  NAND2_X1 U2192 ( .A1(n16791), .A2(n8577), .ZN(n17009) );
  NAND2_X1 U2193 ( .A1(n16791), .A2(n8576), .ZN(n17018) );
  NAND2_X1 U2194 ( .A1(n16791), .A2(n9503), .ZN(n17027) );
  NAND2_X1 U2195 ( .A1(n16791), .A2(n8574), .ZN(n17036) );
  NAND2_X1 U2196 ( .A1(n16791), .A2(n8573), .ZN(n17045) );
  NAND2_X1 U2197 ( .A1(n16791), .A2(n8572), .ZN(n17054) );
  NAND2_X1 U2198 ( .A1(n16791), .A2(n8571), .ZN(n17063) );
  NAND2_X1 U2199 ( .A1(n17080), .A2(n9232), .ZN(n17072) );
  NAND2_X1 U2200 ( .A1(n17080), .A2(n9243), .ZN(n17082) );
  NAND2_X1 U2201 ( .A1(n17080), .A2(n9253), .ZN(n17091) );
  NAND2_X1 U2202 ( .A1(n17080), .A2(n9263), .ZN(n17100) );
  NAND2_X1 U2203 ( .A1(n17080), .A2(n8598), .ZN(n17109) );
  NAND2_X1 U2204 ( .A1(n17080), .A2(n9283), .ZN(n17118) );
  NAND2_X1 U2205 ( .A1(n17080), .A2(n9293), .ZN(n17127) );
  NAND2_X1 U2206 ( .A1(n17080), .A2(n8595), .ZN(n17136) );
  NAND2_X1 U2207 ( .A1(n8544), .A2(n9313), .ZN(n17145) );
  NAND2_X1 U2208 ( .A1(n8544), .A2(n9323), .ZN(n17154) );
  NAND2_X1 U2209 ( .A1(n8544), .A2(n9333), .ZN(n17163) );
  NAND2_X1 U2210 ( .A1(n8544), .A2(n9343), .ZN(n17172) );
  NAND2_X1 U2211 ( .A1(n8544), .A2(n9353), .ZN(n17181) );
  NAND2_X1 U2212 ( .A1(n8544), .A2(n9363), .ZN(n17190) );
  NAND2_X1 U2213 ( .A1(n8544), .A2(n8588), .ZN(n17199) );
  NAND2_X1 U2214 ( .A1(n8544), .A2(n9383), .ZN(n17208) );
  NAND2_X1 U2215 ( .A1(n8544), .A2(n9393), .ZN(n17217) );
  NAND2_X1 U2216 ( .A1(n8544), .A2(n8585), .ZN(n17226) );
  NAND2_X1 U2217 ( .A1(n8544), .A2(n9413), .ZN(n17235) );
  NAND2_X1 U2218 ( .A1(n8544), .A2(n9423), .ZN(n17244) );
  NAND2_X1 U2219 ( .A1(n17080), .A2(n9433), .ZN(n17253) );
  NAND2_X1 U2220 ( .A1(n17080), .A2(n9443), .ZN(n17262) );
  NAND2_X1 U2221 ( .A1(n17080), .A2(n9453), .ZN(n17271) );
  NAND2_X1 U2222 ( .A1(n17080), .A2(n9463), .ZN(n17280) );
  NAND2_X1 U2223 ( .A1(n17080), .A2(n8578), .ZN(n17289) );
  NAND2_X1 U2224 ( .A1(n17080), .A2(n9483), .ZN(n17298) );
  NAND2_X1 U2225 ( .A1(n17080), .A2(n9493), .ZN(n17307) );
  NAND2_X1 U2226 ( .A1(n17080), .A2(n8575), .ZN(n17316) );
  NAND2_X1 U2227 ( .A1(n17080), .A2(n9513), .ZN(n17325) );
  NAND2_X1 U2228 ( .A1(n17080), .A2(n9523), .ZN(n17334) );
  NAND2_X1 U2229 ( .A1(n17080), .A2(n9533), .ZN(n17343) );
  NAND2_X1 U2230 ( .A1(n17080), .A2(n9543), .ZN(n17352) );
  NAND2_X1 U2231 ( .A1(n17369), .A2(n8603), .ZN(n17361) );
  NAND2_X1 U2232 ( .A1(n17369), .A2(n8601), .ZN(n17371) );
  NAND2_X1 U2233 ( .A1(n17369), .A2(n8600), .ZN(n17380) );
  NAND2_X1 U2234 ( .A1(n17369), .A2(n8599), .ZN(n17389) );
  NAND2_X1 U2235 ( .A1(n17369), .A2(n8598), .ZN(n17398) );
  NAND2_X1 U2236 ( .A1(n17369), .A2(n8597), .ZN(n17407) );
  NAND2_X1 U2237 ( .A1(n17369), .A2(n8596), .ZN(n17416) );
  NAND2_X1 U2238 ( .A1(n17369), .A2(n9303), .ZN(n17425) );
  NAND2_X1 U2239 ( .A1(n8543), .A2(n8594), .ZN(n17434) );
  NAND2_X1 U2240 ( .A1(n8543), .A2(n8593), .ZN(n17443) );
  NAND2_X1 U2241 ( .A1(n8543), .A2(n8592), .ZN(n17452) );
  NAND2_X1 U2242 ( .A1(n8543), .A2(n8591), .ZN(n17461) );
  NAND2_X1 U2243 ( .A1(n8543), .A2(n8590), .ZN(n17470) );
  NAND2_X1 U2244 ( .A1(n8543), .A2(n8589), .ZN(n17479) );
  NAND2_X1 U2245 ( .A1(n8543), .A2(n8588), .ZN(n17488) );
  NAND2_X1 U2246 ( .A1(n8543), .A2(n8587), .ZN(n17497) );
  NAND2_X1 U2247 ( .A1(n8543), .A2(n8586), .ZN(n17506) );
  NAND2_X1 U2248 ( .A1(n8543), .A2(n9403), .ZN(n17515) );
  NAND2_X1 U2249 ( .A1(n8543), .A2(n8584), .ZN(n17524) );
  NAND2_X1 U2250 ( .A1(n8543), .A2(n8583), .ZN(n17533) );
  NAND2_X1 U2251 ( .A1(n17369), .A2(n8582), .ZN(n17542) );
  NAND2_X1 U2252 ( .A1(n17369), .A2(n8581), .ZN(n17551) );
  NAND2_X1 U2253 ( .A1(n17369), .A2(n8580), .ZN(n17560) );
  NAND2_X1 U2254 ( .A1(n17369), .A2(n8579), .ZN(n17569) );
  NAND2_X1 U2255 ( .A1(n17369), .A2(n8578), .ZN(n17578) );
  NAND2_X1 U2256 ( .A1(n17369), .A2(n8577), .ZN(n17587) );
  NAND2_X1 U2257 ( .A1(n17369), .A2(n8576), .ZN(n17596) );
  NAND2_X1 U2258 ( .A1(n17369), .A2(n9503), .ZN(n17605) );
  NAND2_X1 U2259 ( .A1(n17369), .A2(n8574), .ZN(n17614) );
  NAND2_X1 U2260 ( .A1(n17369), .A2(n8573), .ZN(n17623) );
  NAND2_X1 U2261 ( .A1(n17369), .A2(n8572), .ZN(n17632) );
  NAND2_X1 U2262 ( .A1(n17369), .A2(n8571), .ZN(n17641) );
  NAND2_X1 U2263 ( .A1(n17658), .A2(n9232), .ZN(n17650) );
  NAND2_X1 U2264 ( .A1(n17658), .A2(n9243), .ZN(n17660) );
  NAND2_X1 U2265 ( .A1(n17658), .A2(n9253), .ZN(n17669) );
  NAND2_X1 U2266 ( .A1(n17658), .A2(n9263), .ZN(n17678) );
  NAND2_X1 U2267 ( .A1(n17658), .A2(n8598), .ZN(n17687) );
  NAND2_X1 U2268 ( .A1(n17658), .A2(n9283), .ZN(n17696) );
  NAND2_X1 U2269 ( .A1(n17658), .A2(n9293), .ZN(n17705) );
  NAND2_X1 U2270 ( .A1(n17658), .A2(n8595), .ZN(n17714) );
  NAND2_X1 U2271 ( .A1(n17658), .A2(n9313), .ZN(n17723) );
  NAND2_X1 U2272 ( .A1(n17658), .A2(n9323), .ZN(n17732) );
  NAND2_X1 U2273 ( .A1(n17658), .A2(n9333), .ZN(n17741) );
  NAND2_X1 U2274 ( .A1(n17658), .A2(n9343), .ZN(n17750) );
  NAND2_X1 U2275 ( .A1(n17658), .A2(n9353), .ZN(n17759) );
  NAND2_X1 U2276 ( .A1(n17658), .A2(n9363), .ZN(n17768) );
  NAND2_X1 U2277 ( .A1(n17658), .A2(n8588), .ZN(n17777) );
  NAND2_X1 U2278 ( .A1(n17658), .A2(n9383), .ZN(n17786) );
  NAND2_X1 U2279 ( .A1(n17658), .A2(n9393), .ZN(n17795) );
  NAND2_X1 U2280 ( .A1(n17658), .A2(n8585), .ZN(n17804) );
  NAND2_X1 U2281 ( .A1(n17658), .A2(n9413), .ZN(n17813) );
  NAND2_X1 U2282 ( .A1(n17658), .A2(n9423), .ZN(n17822) );
  NAND2_X1 U2283 ( .A1(n8542), .A2(n9433), .ZN(n17831) );
  NAND2_X1 U2284 ( .A1(n8542), .A2(n9443), .ZN(n17840) );
  NAND2_X1 U2285 ( .A1(n8542), .A2(n9453), .ZN(n17849) );
  NAND2_X1 U2286 ( .A1(n8542), .A2(n9463), .ZN(n17858) );
  NAND2_X1 U2287 ( .A1(n8542), .A2(n8578), .ZN(n17867) );
  NAND2_X1 U2288 ( .A1(n8542), .A2(n9483), .ZN(n17876) );
  NAND2_X1 U2289 ( .A1(n8542), .A2(n9493), .ZN(n17885) );
  NAND2_X1 U2290 ( .A1(n8542), .A2(n8575), .ZN(n17894) );
  NAND2_X1 U2291 ( .A1(n8542), .A2(n9513), .ZN(n17903) );
  NAND2_X1 U2292 ( .A1(n8542), .A2(n9523), .ZN(n17912) );
  NAND2_X1 U2293 ( .A1(n8542), .A2(n9533), .ZN(n17921) );
  NAND2_X1 U2294 ( .A1(n8542), .A2(n9543), .ZN(n17930) );
  NAND2_X1 U2295 ( .A1(n17947), .A2(n8603), .ZN(n17939) );
  NAND2_X1 U2296 ( .A1(n17947), .A2(n8601), .ZN(n17949) );
  NAND2_X1 U2297 ( .A1(n17947), .A2(n8600), .ZN(n17958) );
  NAND2_X1 U2298 ( .A1(n17947), .A2(n8599), .ZN(n17967) );
  NAND2_X1 U2299 ( .A1(n17947), .A2(n8598), .ZN(n17976) );
  NAND2_X1 U2300 ( .A1(n17947), .A2(n8597), .ZN(n17985) );
  NAND2_X1 U2301 ( .A1(n17947), .A2(n8596), .ZN(n17994) );
  NAND2_X1 U2302 ( .A1(n17947), .A2(n9303), .ZN(n18003) );
  NAND2_X1 U2303 ( .A1(n8541), .A2(n8594), .ZN(n18012) );
  NAND2_X1 U2304 ( .A1(n8541), .A2(n8593), .ZN(n18021) );
  NAND2_X1 U2305 ( .A1(n8541), .A2(n8592), .ZN(n18030) );
  NAND2_X1 U2306 ( .A1(n8541), .A2(n8591), .ZN(n18039) );
  NAND2_X1 U2307 ( .A1(n8541), .A2(n8590), .ZN(n18048) );
  NAND2_X1 U2308 ( .A1(n8541), .A2(n8589), .ZN(n18057) );
  NAND2_X1 U2309 ( .A1(n8541), .A2(n8588), .ZN(n18066) );
  NAND2_X1 U2310 ( .A1(n8541), .A2(n8587), .ZN(n18075) );
  NAND2_X1 U2311 ( .A1(n8541), .A2(n8586), .ZN(n18084) );
  NAND2_X1 U2312 ( .A1(n8541), .A2(n9403), .ZN(n18093) );
  NAND2_X1 U2313 ( .A1(n8541), .A2(n8584), .ZN(n18102) );
  NAND2_X1 U2314 ( .A1(n8541), .A2(n8583), .ZN(n18111) );
  NAND2_X1 U2315 ( .A1(n17947), .A2(n8582), .ZN(n18120) );
  NAND2_X1 U2316 ( .A1(n17947), .A2(n8581), .ZN(n18129) );
  NAND2_X1 U2317 ( .A1(n17947), .A2(n8580), .ZN(n18138) );
  NAND2_X1 U2318 ( .A1(n17947), .A2(n8579), .ZN(n18147) );
  NAND2_X1 U2319 ( .A1(n17947), .A2(n8578), .ZN(n18156) );
  NAND2_X1 U2320 ( .A1(n17947), .A2(n8577), .ZN(n18165) );
  NAND2_X1 U2321 ( .A1(n17947), .A2(n8576), .ZN(n18174) );
  NAND2_X1 U2322 ( .A1(n17947), .A2(n9503), .ZN(n18183) );
  NAND2_X1 U2323 ( .A1(n17947), .A2(n8574), .ZN(n18192) );
  NAND2_X1 U2324 ( .A1(n17947), .A2(n8573), .ZN(n18201) );
  NAND2_X1 U2325 ( .A1(n17947), .A2(n8572), .ZN(n18210) );
  NAND2_X1 U2326 ( .A1(n17947), .A2(n8571), .ZN(n18219) );
  NAND2_X1 U2327 ( .A1(n18236), .A2(n9232), .ZN(n18228) );
  NAND2_X1 U2328 ( .A1(n18236), .A2(n9243), .ZN(n18240) );
  NAND2_X1 U2329 ( .A1(n18236), .A2(n9253), .ZN(n18250) );
  NAND2_X1 U2330 ( .A1(n18236), .A2(n9263), .ZN(n18260) );
  NAND2_X1 U2331 ( .A1(n18236), .A2(n8598), .ZN(n18270) );
  NAND2_X1 U2332 ( .A1(n18236), .A2(n9283), .ZN(n18280) );
  NAND2_X1 U2333 ( .A1(n18236), .A2(n9293), .ZN(n18290) );
  NAND2_X1 U2334 ( .A1(n18236), .A2(n8595), .ZN(n18300) );
  NAND2_X1 U2335 ( .A1(n8540), .A2(n9313), .ZN(n18310) );
  NAND2_X1 U2336 ( .A1(n8540), .A2(n9323), .ZN(n18320) );
  NAND2_X1 U2337 ( .A1(n8540), .A2(n9333), .ZN(n18329) );
  NAND2_X1 U2338 ( .A1(n8540), .A2(n9343), .ZN(n18338) );
  NAND2_X1 U2339 ( .A1(n8540), .A2(n9353), .ZN(n18347) );
  NAND2_X1 U2340 ( .A1(n8540), .A2(n9363), .ZN(n18356) );
  NAND2_X1 U2341 ( .A1(n8540), .A2(n8588), .ZN(n18365) );
  NAND2_X1 U2342 ( .A1(n8540), .A2(n9383), .ZN(n18374) );
  NAND2_X1 U2343 ( .A1(n8540), .A2(n9393), .ZN(n18383) );
  NAND2_X1 U2344 ( .A1(n8540), .A2(n8585), .ZN(n18393) );
  NAND2_X1 U2345 ( .A1(n8540), .A2(n9413), .ZN(n18402) );
  NAND2_X1 U2346 ( .A1(n8540), .A2(n9423), .ZN(n18411) );
  NAND2_X1 U2347 ( .A1(n18236), .A2(n9433), .ZN(n18420) );
  NAND2_X1 U2348 ( .A1(n18236), .A2(n9443), .ZN(n18429) );
  NAND2_X1 U2349 ( .A1(n18236), .A2(n9453), .ZN(n18438) );
  NAND2_X1 U2350 ( .A1(n18236), .A2(n9463), .ZN(n18447) );
  NAND2_X1 U2351 ( .A1(n18236), .A2(n8578), .ZN(n18456) );
  NAND2_X1 U2352 ( .A1(n18236), .A2(n9483), .ZN(n18466) );
  NAND2_X1 U2353 ( .A1(n18236), .A2(n9493), .ZN(n18475) );
  NAND2_X1 U2354 ( .A1(n18236), .A2(n8575), .ZN(n18484) );
  NAND2_X1 U2355 ( .A1(n18236), .A2(n9513), .ZN(n18493) );
  NAND2_X1 U2356 ( .A1(n18236), .A2(n9523), .ZN(n18502) );
  NAND2_X1 U2357 ( .A1(n18236), .A2(n9533), .ZN(n18511) );
  NAND2_X1 U2358 ( .A1(n18236), .A2(n9543), .ZN(n18520) );
  BUF_X1 U2359 ( .A(n8185), .Z(n8181) );
  BUF_X1 U2360 ( .A(n8185), .Z(n8182) );
  BUF_X1 U2361 ( .A(n8185), .Z(n8183) );
  BUF_X1 U2362 ( .A(n8185), .Z(n8184) );
  BUF_X1 U2363 ( .A(N21), .Z(n8200) );
  BUF_X1 U2364 ( .A(n8219), .Z(n8199) );
  BUF_X1 U2365 ( .A(n8219), .Z(n8198) );
  BUF_X1 U2366 ( .A(n8357), .Z(n8387) );
  BUF_X1 U2367 ( .A(n8357), .Z(n8386) );
  BUF_X1 U2368 ( .A(n8265), .Z(n8224) );
  BUF_X1 U2369 ( .A(n8265), .Z(n8223) );
  BUF_X1 U2370 ( .A(n8264), .Z(n8222) );
  BUF_X1 U2371 ( .A(n8264), .Z(n8221) );
  BUF_X1 U2372 ( .A(n8264), .Z(n8220) );
  BUF_X1 U2373 ( .A(n8357), .Z(n8388) );
  BUF_X1 U2374 ( .A(n8265), .Z(n8225) );
  BUF_X1 U2375 ( .A(n8219), .Z(n8197) );
  BUF_X1 U2376 ( .A(n8460), .Z(n8358) );
  BUF_X1 U2377 ( .A(n8538), .Z(n8359) );
  BUF_X1 U2378 ( .A(n8538), .Z(n8360) );
  BUF_X1 U2379 ( .A(n8538), .Z(n8361) );
  BUF_X1 U2380 ( .A(n8539), .Z(n8362) );
  BUF_X1 U2381 ( .A(n8539), .Z(n8363) );
  BUF_X1 U2382 ( .A(n8539), .Z(n8364) );
  BUF_X1 U2383 ( .A(n8356), .Z(n8266) );
  BUF_X1 U2384 ( .A(n8356), .Z(n8267) );
  BUF_X1 U2385 ( .A(n8356), .Z(n8268) );
  BUF_X1 U2386 ( .A(n8356), .Z(n8269) );
  BUF_X1 U2387 ( .A(n9233), .Z(n8602) );
  BUF_X1 U2388 ( .A(n9556), .Z(n8570) );
  BUF_X1 U2389 ( .A(n9846), .Z(n8569) );
  BUF_X1 U2390 ( .A(n10136), .Z(n8568) );
  BUF_X1 U2391 ( .A(n10716), .Z(n8566) );
  BUF_X1 U2392 ( .A(n11006), .Z(n8565) );
  BUF_X1 U2393 ( .A(n11296), .Z(n8564) );
  BUF_X1 U2394 ( .A(n11586), .Z(n8563) );
  BUF_X1 U2395 ( .A(n11876), .Z(n8562) );
  BUF_X1 U2396 ( .A(n12165), .Z(n8561) );
  BUF_X1 U2397 ( .A(n12454), .Z(n8560) );
  BUF_X1 U2398 ( .A(n12743), .Z(n8559) );
  BUF_X1 U2399 ( .A(n13032), .Z(n8558) );
  BUF_X1 U2400 ( .A(n13610), .Z(n8556) );
  BUF_X1 U2401 ( .A(n14189), .Z(n8554) );
  BUF_X1 U2402 ( .A(n14478), .Z(n8553) );
  BUF_X1 U2403 ( .A(n14767), .Z(n8552) );
  BUF_X1 U2404 ( .A(n15056), .Z(n8551) );
  BUF_X1 U2405 ( .A(n15345), .Z(n8550) );
  BUF_X1 U2406 ( .A(n15634), .Z(n8549) );
  BUF_X1 U2407 ( .A(n15923), .Z(n8548) );
  BUF_X1 U2408 ( .A(n16212), .Z(n8547) );
  BUF_X1 U2409 ( .A(n16502), .Z(n8546) );
  BUF_X1 U2410 ( .A(n16791), .Z(n8545) );
  BUF_X1 U2411 ( .A(n17080), .Z(n8544) );
  BUF_X1 U2412 ( .A(n17369), .Z(n8543) );
  BUF_X1 U2413 ( .A(n17658), .Z(n8542) );
  BUF_X1 U2414 ( .A(n17947), .Z(n8541) );
  BUF_X1 U2415 ( .A(n18236), .Z(n8540) );
  BUF_X1 U2416 ( .A(n10426), .Z(n8567) );
  BUF_X1 U2417 ( .A(n13321), .Z(n8557) );
  BUF_X1 U2418 ( .A(n13899), .Z(n8555) );
  BUF_X1 U2419 ( .A(N24), .Z(n8179) );
  BUF_X1 U2420 ( .A(N24), .Z(n8180) );
  BUF_X1 U2421 ( .A(n8196), .Z(n8189) );
  BUF_X1 U2422 ( .A(n8196), .Z(n8192) );
  BUF_X1 U2423 ( .A(n8196), .Z(n8193) );
  BUF_X1 U2424 ( .A(n8196), .Z(n8194) );
  BUF_X1 U2425 ( .A(n9232), .Z(n8603) );
  BUF_X1 U2426 ( .A(n9243), .Z(n8601) );
  BUF_X1 U2427 ( .A(n9253), .Z(n8600) );
  BUF_X1 U2428 ( .A(n9263), .Z(n8599) );
  BUF_X1 U2429 ( .A(n9283), .Z(n8597) );
  BUF_X1 U2430 ( .A(n9293), .Z(n8596) );
  BUF_X1 U2431 ( .A(n9313), .Z(n8594) );
  BUF_X1 U2432 ( .A(n9323), .Z(n8593) );
  BUF_X1 U2433 ( .A(n9333), .Z(n8592) );
  BUF_X1 U2434 ( .A(n9343), .Z(n8591) );
  BUF_X1 U2435 ( .A(n9353), .Z(n8590) );
  BUF_X1 U2436 ( .A(n9363), .Z(n8589) );
  BUF_X1 U2437 ( .A(n9383), .Z(n8587) );
  BUF_X1 U2438 ( .A(n9393), .Z(n8586) );
  BUF_X1 U2439 ( .A(n9413), .Z(n8584) );
  BUF_X1 U2440 ( .A(n9423), .Z(n8583) );
  BUF_X1 U2441 ( .A(n9433), .Z(n8582) );
  BUF_X1 U2442 ( .A(n9443), .Z(n8581) );
  BUF_X1 U2443 ( .A(n9453), .Z(n8580) );
  BUF_X1 U2444 ( .A(n9463), .Z(n8579) );
  BUF_X1 U2445 ( .A(n9483), .Z(n8577) );
  BUF_X1 U2446 ( .A(n9493), .Z(n8576) );
  BUF_X1 U2447 ( .A(n9513), .Z(n8574) );
  BUF_X1 U2448 ( .A(n9523), .Z(n8573) );
  BUF_X1 U2449 ( .A(n9533), .Z(n8572) );
  BUF_X1 U2450 ( .A(n9543), .Z(n8571) );
  BUF_X1 U2451 ( .A(n9273), .Z(n8598) );
  BUF_X1 U2452 ( .A(n9373), .Z(n8588) );
  BUF_X1 U2453 ( .A(n9473), .Z(n8578) );
  BUF_X1 U2454 ( .A(n9303), .Z(n8595) );
  BUF_X1 U2455 ( .A(n9403), .Z(n8585) );
  BUF_X1 U2456 ( .A(n9503), .Z(n8575) );
  BUF_X1 U2457 ( .A(n8195), .Z(n8186) );
  BUF_X1 U2458 ( .A(n8192), .Z(n8187) );
  BUF_X1 U2459 ( .A(n8193), .Z(n8188) );
  BUF_X1 U2460 ( .A(n8196), .Z(n8190) );
  BUF_X1 U2461 ( .A(n8196), .Z(n8191) );
  BUF_X1 U2462 ( .A(N23), .Z(n8185) );
  BUF_X1 U2463 ( .A(N18), .Z(n8538) );
  BUF_X1 U2464 ( .A(N18), .Z(n8539) );
  BUF_X1 U2465 ( .A(N19), .Z(n8356) );
  BUF_X1 U2466 ( .A(N21), .Z(n8219) );
  BUF_X1 U2467 ( .A(n8537), .Z(n8357) );
  BUF_X1 U2468 ( .A(N18), .Z(n8537) );
  BUF_X1 U2469 ( .A(n8263), .Z(n8265) );
  BUF_X1 U2470 ( .A(n8263), .Z(n8264) );
  AND3_X1 U2471 ( .A1(n9544), .A2(n9545), .A3(n9546), .ZN(n9233) );
  AND3_X1 U2472 ( .A1(n9544), .A2(n9545), .A3(n9836), .ZN(n9556) );
  AND3_X1 U2473 ( .A1(n9544), .A2(n9545), .A3(n10126), .ZN(n9846) );
  AND3_X1 U2474 ( .A1(n9544), .A2(n9545), .A3(n10416), .ZN(n10136) );
  AND3_X1 U2475 ( .A1(n9544), .A2(n9545), .A3(n10706), .ZN(n10426) );
  AND3_X1 U2476 ( .A1(n9544), .A2(n9545), .A3(n10996), .ZN(n10716) );
  AND3_X1 U2477 ( .A1(n9544), .A2(n9545), .A3(n11286), .ZN(n11006) );
  AND3_X1 U2478 ( .A1(n9544), .A2(n9545), .A3(n11576), .ZN(n11296) );
  AND3_X1 U2479 ( .A1(n9546), .A2(n9545), .A3(n11866), .ZN(n11586) );
  AND3_X1 U2480 ( .A1(n9836), .A2(n9545), .A3(n11866), .ZN(n11876) );
  AND3_X1 U2481 ( .A1(n10126), .A2(n9545), .A3(n11866), .ZN(n12165) );
  AND3_X1 U2482 ( .A1(n10416), .A2(n9545), .A3(n11866), .ZN(n12454) );
  AND3_X1 U2483 ( .A1(n9546), .A2(n9545), .A3(n14179), .ZN(n13899) );
  AND3_X1 U2484 ( .A1(n9836), .A2(n9545), .A3(n14179), .ZN(n14189) );
  AND3_X1 U2485 ( .A1(n10126), .A2(n9545), .A3(n14179), .ZN(n14478) );
  AND3_X1 U2486 ( .A1(n10416), .A2(n9545), .A3(n14179), .ZN(n14767) );
  AND3_X1 U2487 ( .A1(n9546), .A2(n9545), .A3(n16492), .ZN(n16212) );
  AND3_X1 U2488 ( .A1(n9836), .A2(n9545), .A3(n16492), .ZN(n16502) );
  AND3_X1 U2489 ( .A1(n10126), .A2(n9545), .A3(n16492), .ZN(n16791) );
  AND3_X1 U2490 ( .A1(n10416), .A2(n9545), .A3(n16492), .ZN(n17080) );
  AND3_X1 U2491 ( .A1(n10706), .A2(n9545), .A3(n11866), .ZN(n12743) );
  AND3_X1 U2492 ( .A1(n10996), .A2(n9545), .A3(n11866), .ZN(n13032) );
  AND3_X1 U2493 ( .A1(n11286), .A2(n9545), .A3(n11866), .ZN(n13321) );
  AND3_X1 U2494 ( .A1(n11576), .A2(n9545), .A3(n11866), .ZN(n13610) );
  AND3_X1 U2495 ( .A1(n10706), .A2(n9545), .A3(n16492), .ZN(n17369) );
  AND3_X1 U2496 ( .A1(n10996), .A2(n9545), .A3(n16492), .ZN(n17658) );
  AND3_X1 U2497 ( .A1(n11286), .A2(n9545), .A3(n16492), .ZN(n17947) );
  AND3_X1 U2498 ( .A1(n11576), .A2(n9545), .A3(n16492), .ZN(n18236) );
  AND3_X1 U2499 ( .A1(n10706), .A2(n9545), .A3(n14179), .ZN(n15056) );
  AND3_X1 U2500 ( .A1(n10996), .A2(n9545), .A3(n14179), .ZN(n15345) );
  AND3_X1 U2501 ( .A1(n11286), .A2(n9545), .A3(n14179), .ZN(n15634) );
  AND3_X1 U2502 ( .A1(n11576), .A2(n9545), .A3(n14179), .ZN(n15923) );
  NOR3_X1 U2503 ( .A1(N19), .A2(N20), .A3(N18), .ZN(n18237) );
  NOR3_X1 U2504 ( .A1(N19), .A2(N20), .A3(n8604), .ZN(n18248) );
  NOR3_X1 U2505 ( .A1(N18), .A2(N20), .A3(n8605), .ZN(n18258) );
  NOR3_X1 U2506 ( .A1(n8604), .A2(N20), .A3(n8605), .ZN(n18268) );
  BUF_X1 U2507 ( .A(n8195), .Z(n8196) );
  AND3_X1 U2508 ( .A1(N18), .A2(n8605), .A3(N20), .ZN(n18288) );
  AND3_X1 U2509 ( .A1(N19), .A2(N18), .A3(N20), .ZN(n18308) );
  AND3_X1 U2510 ( .A1(N19), .A2(n8604), .A3(N20), .ZN(n18298) );
  AND3_X1 U2511 ( .A1(n8604), .A2(n8605), .A3(N20), .ZN(n18278) );
  AND2_X1 U2512 ( .A1(n18318), .A2(n18237), .ZN(n9313) );
  AND2_X1 U2513 ( .A1(n18318), .A2(n18248), .ZN(n9323) );
  AND2_X1 U2514 ( .A1(n18318), .A2(n18258), .ZN(n9333) );
  AND2_X1 U2515 ( .A1(n18318), .A2(n18268), .ZN(n9343) );
  AND2_X1 U2516 ( .A1(n18318), .A2(n18278), .ZN(n9353) );
  AND2_X1 U2517 ( .A1(n18318), .A2(n18288), .ZN(n9363) );
  AND2_X1 U2518 ( .A1(n18318), .A2(n18298), .ZN(n9373) );
  AND2_X1 U2519 ( .A1(n18318), .A2(n18308), .ZN(n9383) );
  AND2_X1 U2520 ( .A1(n18237), .A2(n18238), .ZN(n9232) );
  AND2_X1 U2521 ( .A1(n18248), .A2(n18238), .ZN(n9243) );
  AND2_X1 U2522 ( .A1(n18258), .A2(n18238), .ZN(n9253) );
  AND2_X1 U2523 ( .A1(n18268), .A2(n18238), .ZN(n9263) );
  AND2_X1 U2524 ( .A1(n18278), .A2(n18238), .ZN(n9273) );
  AND2_X1 U2525 ( .A1(n18288), .A2(n18238), .ZN(n9283) );
  AND2_X1 U2526 ( .A1(n18298), .A2(n18238), .ZN(n9293) );
  AND2_X1 U2527 ( .A1(n18308), .A2(n18238), .ZN(n9303) );
  AND2_X1 U2528 ( .A1(n18391), .A2(n18237), .ZN(n9393) );
  AND2_X1 U2529 ( .A1(n18391), .A2(n18248), .ZN(n9403) );
  AND2_X1 U2530 ( .A1(n18391), .A2(n18258), .ZN(n9413) );
  AND2_X1 U2531 ( .A1(n18391), .A2(n18268), .ZN(n9423) );
  AND2_X1 U2532 ( .A1(n18464), .A2(n18237), .ZN(n9473) );
  AND2_X1 U2533 ( .A1(n18464), .A2(n18248), .ZN(n9483) );
  AND2_X1 U2534 ( .A1(n18464), .A2(n18258), .ZN(n9493) );
  AND2_X1 U2535 ( .A1(n18464), .A2(n18268), .ZN(n9503) );
  AND2_X1 U2536 ( .A1(n18391), .A2(n18278), .ZN(n9433) );
  AND2_X1 U2537 ( .A1(n18391), .A2(n18288), .ZN(n9443) );
  AND2_X1 U2538 ( .A1(n18391), .A2(n18298), .ZN(n9453) );
  AND2_X1 U2539 ( .A1(n18391), .A2(n18308), .ZN(n9463) );
  AND2_X1 U2540 ( .A1(n18464), .A2(n18278), .ZN(n9513) );
  AND2_X1 U2541 ( .A1(n18464), .A2(n18288), .ZN(n9523) );
  AND2_X1 U2542 ( .A1(n18464), .A2(n18298), .ZN(n9533) );
  AND2_X1 U2543 ( .A1(n18464), .A2(n18308), .ZN(n9543) );
  BUF_X1 U2544 ( .A(N20), .Z(n8263) );
  AND2_X1 U2545 ( .A1(n18528), .A2(wr_en), .ZN(n9545) );
  NOR2_X1 U2546 ( .A1(addr[11]), .A2(addr[10]), .ZN(n18528) );
  INV_X1 U2547 ( .A(n9223), .ZN(n26106) );
  AOI22_X1 U2548 ( .A1(\mem[0][0] ), .A2(n9224), .B1(data_in[0]), .B2(n27130), 
        .ZN(n9223) );
  INV_X1 U2549 ( .A(n9225), .ZN(n26105) );
  AOI22_X1 U2550 ( .A1(\mem[0][1] ), .A2(n9224), .B1(data_in[1]), .B2(n27130), 
        .ZN(n9225) );
  INV_X1 U2551 ( .A(n9226), .ZN(n26104) );
  AOI22_X1 U2552 ( .A1(\mem[0][2] ), .A2(n9224), .B1(data_in[2]), .B2(n27130), 
        .ZN(n9226) );
  INV_X1 U2553 ( .A(n9227), .ZN(n26103) );
  AOI22_X1 U2554 ( .A1(\mem[0][3] ), .A2(n9224), .B1(data_in[3]), .B2(n27130), 
        .ZN(n9227) );
  INV_X1 U2555 ( .A(n9228), .ZN(n26102) );
  AOI22_X1 U2556 ( .A1(\mem[0][4] ), .A2(n9224), .B1(data_in[4]), .B2(n27130), 
        .ZN(n9228) );
  INV_X1 U2557 ( .A(n9229), .ZN(n26101) );
  AOI22_X1 U2558 ( .A1(\mem[0][5] ), .A2(n9224), .B1(data_in[5]), .B2(n27130), 
        .ZN(n9229) );
  INV_X1 U2559 ( .A(n9230), .ZN(n26100) );
  AOI22_X1 U2560 ( .A1(\mem[0][6] ), .A2(n9224), .B1(data_in[6]), .B2(n27130), 
        .ZN(n9230) );
  INV_X1 U2561 ( .A(n9231), .ZN(n26099) );
  AOI22_X1 U2562 ( .A1(\mem[0][7] ), .A2(n9224), .B1(data_in[7]), .B2(n27130), 
        .ZN(n9231) );
  INV_X1 U2563 ( .A(n9234), .ZN(n26098) );
  AOI22_X1 U2564 ( .A1(\mem[1][0] ), .A2(n9235), .B1(n27129), .B2(data_in[0]), 
        .ZN(n9234) );
  INV_X1 U2565 ( .A(n9236), .ZN(n26097) );
  AOI22_X1 U2566 ( .A1(\mem[1][1] ), .A2(n9235), .B1(n27129), .B2(data_in[1]), 
        .ZN(n9236) );
  INV_X1 U2567 ( .A(n9237), .ZN(n26096) );
  AOI22_X1 U2568 ( .A1(\mem[1][2] ), .A2(n9235), .B1(n27129), .B2(data_in[2]), 
        .ZN(n9237) );
  INV_X1 U2569 ( .A(n9238), .ZN(n26095) );
  AOI22_X1 U2570 ( .A1(\mem[1][3] ), .A2(n9235), .B1(n27129), .B2(data_in[3]), 
        .ZN(n9238) );
  INV_X1 U2571 ( .A(n9239), .ZN(n26094) );
  AOI22_X1 U2572 ( .A1(\mem[1][4] ), .A2(n9235), .B1(n27129), .B2(data_in[4]), 
        .ZN(n9239) );
  INV_X1 U2573 ( .A(n9240), .ZN(n26093) );
  AOI22_X1 U2574 ( .A1(\mem[1][5] ), .A2(n9235), .B1(n27129), .B2(data_in[5]), 
        .ZN(n9240) );
  INV_X1 U2575 ( .A(n9241), .ZN(n26092) );
  AOI22_X1 U2576 ( .A1(\mem[1][6] ), .A2(n9235), .B1(n27129), .B2(data_in[6]), 
        .ZN(n9241) );
  INV_X1 U2577 ( .A(n9242), .ZN(n26091) );
  AOI22_X1 U2578 ( .A1(\mem[1][7] ), .A2(n9235), .B1(n27129), .B2(data_in[7]), 
        .ZN(n9242) );
  INV_X1 U2579 ( .A(n9244), .ZN(n26090) );
  AOI22_X1 U2580 ( .A1(\mem[2][0] ), .A2(n9245), .B1(n27128), .B2(data_in[0]), 
        .ZN(n9244) );
  INV_X1 U2581 ( .A(n9246), .ZN(n26089) );
  AOI22_X1 U2582 ( .A1(\mem[2][1] ), .A2(n9245), .B1(n27128), .B2(data_in[1]), 
        .ZN(n9246) );
  INV_X1 U2583 ( .A(n9247), .ZN(n26088) );
  AOI22_X1 U2584 ( .A1(\mem[2][2] ), .A2(n9245), .B1(n27128), .B2(data_in[2]), 
        .ZN(n9247) );
  INV_X1 U2585 ( .A(n9248), .ZN(n26087) );
  AOI22_X1 U2586 ( .A1(\mem[2][3] ), .A2(n9245), .B1(n27128), .B2(data_in[3]), 
        .ZN(n9248) );
  INV_X1 U2587 ( .A(n9249), .ZN(n26086) );
  AOI22_X1 U2588 ( .A1(\mem[2][4] ), .A2(n9245), .B1(n27128), .B2(data_in[4]), 
        .ZN(n9249) );
  INV_X1 U2589 ( .A(n9250), .ZN(n26085) );
  AOI22_X1 U2590 ( .A1(\mem[2][5] ), .A2(n9245), .B1(n27128), .B2(data_in[5]), 
        .ZN(n9250) );
  INV_X1 U2591 ( .A(n9251), .ZN(n26084) );
  AOI22_X1 U2592 ( .A1(\mem[2][6] ), .A2(n9245), .B1(n27128), .B2(data_in[6]), 
        .ZN(n9251) );
  INV_X1 U2593 ( .A(n9252), .ZN(n26083) );
  AOI22_X1 U2594 ( .A1(\mem[2][7] ), .A2(n9245), .B1(n27128), .B2(data_in[7]), 
        .ZN(n9252) );
  INV_X1 U2595 ( .A(n9254), .ZN(n26082) );
  AOI22_X1 U2596 ( .A1(\mem[3][0] ), .A2(n9255), .B1(n27127), .B2(data_in[0]), 
        .ZN(n9254) );
  INV_X1 U2597 ( .A(n9256), .ZN(n26081) );
  AOI22_X1 U2598 ( .A1(\mem[3][1] ), .A2(n9255), .B1(n27127), .B2(data_in[1]), 
        .ZN(n9256) );
  INV_X1 U2599 ( .A(n9257), .ZN(n26080) );
  AOI22_X1 U2600 ( .A1(\mem[3][2] ), .A2(n9255), .B1(n27127), .B2(data_in[2]), 
        .ZN(n9257) );
  INV_X1 U2601 ( .A(n9258), .ZN(n26079) );
  AOI22_X1 U2602 ( .A1(\mem[3][3] ), .A2(n9255), .B1(n27127), .B2(data_in[3]), 
        .ZN(n9258) );
  INV_X1 U2603 ( .A(n9259), .ZN(n26078) );
  AOI22_X1 U2604 ( .A1(\mem[3][4] ), .A2(n9255), .B1(n27127), .B2(data_in[4]), 
        .ZN(n9259) );
  INV_X1 U2605 ( .A(n9260), .ZN(n26077) );
  AOI22_X1 U2606 ( .A1(\mem[3][5] ), .A2(n9255), .B1(n27127), .B2(data_in[5]), 
        .ZN(n9260) );
  INV_X1 U2607 ( .A(n9261), .ZN(n26076) );
  AOI22_X1 U2608 ( .A1(\mem[3][6] ), .A2(n9255), .B1(n27127), .B2(data_in[6]), 
        .ZN(n9261) );
  INV_X1 U2609 ( .A(n9262), .ZN(n26075) );
  AOI22_X1 U2610 ( .A1(\mem[3][7] ), .A2(n9255), .B1(n27127), .B2(data_in[7]), 
        .ZN(n9262) );
  INV_X1 U2611 ( .A(n9264), .ZN(n26074) );
  AOI22_X1 U2612 ( .A1(\mem[4][0] ), .A2(n9265), .B1(n27126), .B2(data_in[0]), 
        .ZN(n9264) );
  INV_X1 U2613 ( .A(n9266), .ZN(n26073) );
  AOI22_X1 U2614 ( .A1(\mem[4][1] ), .A2(n9265), .B1(n27126), .B2(data_in[1]), 
        .ZN(n9266) );
  INV_X1 U2615 ( .A(n9267), .ZN(n26072) );
  AOI22_X1 U2616 ( .A1(\mem[4][2] ), .A2(n9265), .B1(n27126), .B2(data_in[2]), 
        .ZN(n9267) );
  INV_X1 U2617 ( .A(n9268), .ZN(n26071) );
  AOI22_X1 U2618 ( .A1(\mem[4][3] ), .A2(n9265), .B1(n27126), .B2(data_in[3]), 
        .ZN(n9268) );
  INV_X1 U2619 ( .A(n9269), .ZN(n26070) );
  AOI22_X1 U2620 ( .A1(\mem[4][4] ), .A2(n9265), .B1(n27126), .B2(data_in[4]), 
        .ZN(n9269) );
  INV_X1 U2621 ( .A(n9270), .ZN(n26069) );
  AOI22_X1 U2622 ( .A1(\mem[4][5] ), .A2(n9265), .B1(n27126), .B2(data_in[5]), 
        .ZN(n9270) );
  INV_X1 U2623 ( .A(n9271), .ZN(n26068) );
  AOI22_X1 U2624 ( .A1(\mem[4][6] ), .A2(n9265), .B1(n27126), .B2(data_in[6]), 
        .ZN(n9271) );
  INV_X1 U2625 ( .A(n9272), .ZN(n26067) );
  AOI22_X1 U2626 ( .A1(\mem[4][7] ), .A2(n9265), .B1(n27126), .B2(data_in[7]), 
        .ZN(n9272) );
  INV_X1 U2627 ( .A(n9274), .ZN(n26066) );
  AOI22_X1 U2628 ( .A1(\mem[5][0] ), .A2(n9275), .B1(n27125), .B2(data_in[0]), 
        .ZN(n9274) );
  INV_X1 U2629 ( .A(n9276), .ZN(n26065) );
  AOI22_X1 U2630 ( .A1(\mem[5][1] ), .A2(n9275), .B1(n27125), .B2(data_in[1]), 
        .ZN(n9276) );
  INV_X1 U2631 ( .A(n9277), .ZN(n26064) );
  AOI22_X1 U2632 ( .A1(\mem[5][2] ), .A2(n9275), .B1(n27125), .B2(data_in[2]), 
        .ZN(n9277) );
  INV_X1 U2633 ( .A(n9278), .ZN(n26063) );
  AOI22_X1 U2634 ( .A1(\mem[5][3] ), .A2(n9275), .B1(n27125), .B2(data_in[3]), 
        .ZN(n9278) );
  INV_X1 U2635 ( .A(n9279), .ZN(n26062) );
  AOI22_X1 U2636 ( .A1(\mem[5][4] ), .A2(n9275), .B1(n27125), .B2(data_in[4]), 
        .ZN(n9279) );
  INV_X1 U2637 ( .A(n9280), .ZN(n26061) );
  AOI22_X1 U2638 ( .A1(\mem[5][5] ), .A2(n9275), .B1(n27125), .B2(data_in[5]), 
        .ZN(n9280) );
  INV_X1 U2639 ( .A(n9281), .ZN(n26060) );
  AOI22_X1 U2640 ( .A1(\mem[5][6] ), .A2(n9275), .B1(n27125), .B2(data_in[6]), 
        .ZN(n9281) );
  INV_X1 U2641 ( .A(n9282), .ZN(n26059) );
  AOI22_X1 U2642 ( .A1(\mem[5][7] ), .A2(n9275), .B1(n27125), .B2(data_in[7]), 
        .ZN(n9282) );
  INV_X1 U2643 ( .A(n9284), .ZN(n26058) );
  AOI22_X1 U2644 ( .A1(\mem[6][0] ), .A2(n9285), .B1(n27124), .B2(data_in[0]), 
        .ZN(n9284) );
  INV_X1 U2645 ( .A(n9286), .ZN(n26057) );
  AOI22_X1 U2646 ( .A1(\mem[6][1] ), .A2(n9285), .B1(n27124), .B2(data_in[1]), 
        .ZN(n9286) );
  INV_X1 U2647 ( .A(n9287), .ZN(n26056) );
  AOI22_X1 U2648 ( .A1(\mem[6][2] ), .A2(n9285), .B1(n27124), .B2(data_in[2]), 
        .ZN(n9287) );
  INV_X1 U2649 ( .A(n9288), .ZN(n26055) );
  AOI22_X1 U2650 ( .A1(\mem[6][3] ), .A2(n9285), .B1(n27124), .B2(data_in[3]), 
        .ZN(n9288) );
  INV_X1 U2651 ( .A(n9289), .ZN(n26054) );
  AOI22_X1 U2652 ( .A1(\mem[6][4] ), .A2(n9285), .B1(n27124), .B2(data_in[4]), 
        .ZN(n9289) );
  INV_X1 U2653 ( .A(n9290), .ZN(n26053) );
  AOI22_X1 U2654 ( .A1(\mem[6][5] ), .A2(n9285), .B1(n27124), .B2(data_in[5]), 
        .ZN(n9290) );
  INV_X1 U2655 ( .A(n9291), .ZN(n26052) );
  AOI22_X1 U2656 ( .A1(\mem[6][6] ), .A2(n9285), .B1(n27124), .B2(data_in[6]), 
        .ZN(n9291) );
  INV_X1 U2657 ( .A(n9292), .ZN(n26051) );
  AOI22_X1 U2658 ( .A1(\mem[6][7] ), .A2(n9285), .B1(n27124), .B2(data_in[7]), 
        .ZN(n9292) );
  INV_X1 U2659 ( .A(n9294), .ZN(n26050) );
  AOI22_X1 U2660 ( .A1(\mem[7][0] ), .A2(n9295), .B1(n27123), .B2(data_in[0]), 
        .ZN(n9294) );
  INV_X1 U2661 ( .A(n9296), .ZN(n26049) );
  AOI22_X1 U2662 ( .A1(\mem[7][1] ), .A2(n9295), .B1(n27123), .B2(data_in[1]), 
        .ZN(n9296) );
  INV_X1 U2663 ( .A(n9297), .ZN(n26048) );
  AOI22_X1 U2664 ( .A1(\mem[7][2] ), .A2(n9295), .B1(n27123), .B2(data_in[2]), 
        .ZN(n9297) );
  INV_X1 U2665 ( .A(n9298), .ZN(n26047) );
  AOI22_X1 U2666 ( .A1(\mem[7][3] ), .A2(n9295), .B1(n27123), .B2(data_in[3]), 
        .ZN(n9298) );
  INV_X1 U2667 ( .A(n9299), .ZN(n26046) );
  AOI22_X1 U2668 ( .A1(\mem[7][4] ), .A2(n9295), .B1(n27123), .B2(data_in[4]), 
        .ZN(n9299) );
  INV_X1 U2669 ( .A(n9300), .ZN(n26045) );
  AOI22_X1 U2670 ( .A1(\mem[7][5] ), .A2(n9295), .B1(n27123), .B2(data_in[5]), 
        .ZN(n9300) );
  INV_X1 U2671 ( .A(n9301), .ZN(n26044) );
  AOI22_X1 U2672 ( .A1(\mem[7][6] ), .A2(n9295), .B1(n27123), .B2(data_in[6]), 
        .ZN(n9301) );
  INV_X1 U2673 ( .A(n9302), .ZN(n26043) );
  AOI22_X1 U2674 ( .A1(\mem[7][7] ), .A2(n9295), .B1(n27123), .B2(data_in[7]), 
        .ZN(n9302) );
  INV_X1 U2675 ( .A(n9304), .ZN(n26042) );
  AOI22_X1 U2676 ( .A1(\mem[8][0] ), .A2(n9305), .B1(n27122), .B2(data_in[0]), 
        .ZN(n9304) );
  INV_X1 U2677 ( .A(n9306), .ZN(n26041) );
  AOI22_X1 U2678 ( .A1(\mem[8][1] ), .A2(n9305), .B1(n27122), .B2(data_in[1]), 
        .ZN(n9306) );
  INV_X1 U2679 ( .A(n9307), .ZN(n26040) );
  AOI22_X1 U2680 ( .A1(\mem[8][2] ), .A2(n9305), .B1(n27122), .B2(data_in[2]), 
        .ZN(n9307) );
  INV_X1 U2681 ( .A(n9308), .ZN(n26039) );
  AOI22_X1 U2682 ( .A1(\mem[8][3] ), .A2(n9305), .B1(n27122), .B2(data_in[3]), 
        .ZN(n9308) );
  INV_X1 U2683 ( .A(n9309), .ZN(n26038) );
  AOI22_X1 U2684 ( .A1(\mem[8][4] ), .A2(n9305), .B1(n27122), .B2(data_in[4]), 
        .ZN(n9309) );
  INV_X1 U2685 ( .A(n9310), .ZN(n26037) );
  AOI22_X1 U2686 ( .A1(\mem[8][5] ), .A2(n9305), .B1(n27122), .B2(data_in[5]), 
        .ZN(n9310) );
  INV_X1 U2687 ( .A(n9311), .ZN(n26036) );
  AOI22_X1 U2688 ( .A1(\mem[8][6] ), .A2(n9305), .B1(n27122), .B2(data_in[6]), 
        .ZN(n9311) );
  INV_X1 U2689 ( .A(n9312), .ZN(n26035) );
  AOI22_X1 U2690 ( .A1(\mem[8][7] ), .A2(n9305), .B1(n27122), .B2(data_in[7]), 
        .ZN(n9312) );
  INV_X1 U2691 ( .A(n9314), .ZN(n26034) );
  AOI22_X1 U2692 ( .A1(\mem[9][0] ), .A2(n9315), .B1(n27121), .B2(data_in[0]), 
        .ZN(n9314) );
  INV_X1 U2693 ( .A(n9316), .ZN(n26033) );
  AOI22_X1 U2694 ( .A1(\mem[9][1] ), .A2(n9315), .B1(n27121), .B2(data_in[1]), 
        .ZN(n9316) );
  INV_X1 U2695 ( .A(n9317), .ZN(n26032) );
  AOI22_X1 U2696 ( .A1(\mem[9][2] ), .A2(n9315), .B1(n27121), .B2(data_in[2]), 
        .ZN(n9317) );
  INV_X1 U2697 ( .A(n9318), .ZN(n26031) );
  AOI22_X1 U2698 ( .A1(\mem[9][3] ), .A2(n9315), .B1(n27121), .B2(data_in[3]), 
        .ZN(n9318) );
  INV_X1 U2699 ( .A(n9319), .ZN(n26030) );
  AOI22_X1 U2700 ( .A1(\mem[9][4] ), .A2(n9315), .B1(n27121), .B2(data_in[4]), 
        .ZN(n9319) );
  INV_X1 U2701 ( .A(n9320), .ZN(n26029) );
  AOI22_X1 U2702 ( .A1(\mem[9][5] ), .A2(n9315), .B1(n27121), .B2(data_in[5]), 
        .ZN(n9320) );
  INV_X1 U2703 ( .A(n9321), .ZN(n26028) );
  AOI22_X1 U2704 ( .A1(\mem[9][6] ), .A2(n9315), .B1(n27121), .B2(data_in[6]), 
        .ZN(n9321) );
  INV_X1 U2705 ( .A(n9322), .ZN(n26027) );
  AOI22_X1 U2706 ( .A1(\mem[9][7] ), .A2(n9315), .B1(n27121), .B2(data_in[7]), 
        .ZN(n9322) );
  INV_X1 U2707 ( .A(n9324), .ZN(n26026) );
  AOI22_X1 U2708 ( .A1(\mem[10][0] ), .A2(n9325), .B1(n27120), .B2(data_in[0]), 
        .ZN(n9324) );
  INV_X1 U2709 ( .A(n9326), .ZN(n26025) );
  AOI22_X1 U2710 ( .A1(\mem[10][1] ), .A2(n9325), .B1(n27120), .B2(data_in[1]), 
        .ZN(n9326) );
  INV_X1 U2711 ( .A(n9327), .ZN(n26024) );
  AOI22_X1 U2712 ( .A1(\mem[10][2] ), .A2(n9325), .B1(n27120), .B2(data_in[2]), 
        .ZN(n9327) );
  INV_X1 U2713 ( .A(n9328), .ZN(n26023) );
  AOI22_X1 U2714 ( .A1(\mem[10][3] ), .A2(n9325), .B1(n27120), .B2(data_in[3]), 
        .ZN(n9328) );
  INV_X1 U2715 ( .A(n9329), .ZN(n26022) );
  AOI22_X1 U2716 ( .A1(\mem[10][4] ), .A2(n9325), .B1(n27120), .B2(data_in[4]), 
        .ZN(n9329) );
  INV_X1 U2717 ( .A(n9330), .ZN(n26021) );
  AOI22_X1 U2718 ( .A1(\mem[10][5] ), .A2(n9325), .B1(n27120), .B2(data_in[5]), 
        .ZN(n9330) );
  INV_X1 U2719 ( .A(n9331), .ZN(n26020) );
  AOI22_X1 U2720 ( .A1(\mem[10][6] ), .A2(n9325), .B1(n27120), .B2(data_in[6]), 
        .ZN(n9331) );
  INV_X1 U2721 ( .A(n9332), .ZN(n26019) );
  AOI22_X1 U2722 ( .A1(\mem[10][7] ), .A2(n9325), .B1(n27120), .B2(data_in[7]), 
        .ZN(n9332) );
  INV_X1 U2723 ( .A(n9334), .ZN(n26018) );
  AOI22_X1 U2724 ( .A1(\mem[11][0] ), .A2(n9335), .B1(n27119), .B2(data_in[0]), 
        .ZN(n9334) );
  INV_X1 U2725 ( .A(n9336), .ZN(n26017) );
  AOI22_X1 U2726 ( .A1(\mem[11][1] ), .A2(n9335), .B1(n27119), .B2(data_in[1]), 
        .ZN(n9336) );
  INV_X1 U2727 ( .A(n9337), .ZN(n26016) );
  AOI22_X1 U2728 ( .A1(\mem[11][2] ), .A2(n9335), .B1(n27119), .B2(data_in[2]), 
        .ZN(n9337) );
  INV_X1 U2729 ( .A(n9338), .ZN(n26015) );
  AOI22_X1 U2730 ( .A1(\mem[11][3] ), .A2(n9335), .B1(n27119), .B2(data_in[3]), 
        .ZN(n9338) );
  INV_X1 U2731 ( .A(n9339), .ZN(n26014) );
  AOI22_X1 U2732 ( .A1(\mem[11][4] ), .A2(n9335), .B1(n27119), .B2(data_in[4]), 
        .ZN(n9339) );
  INV_X1 U2733 ( .A(n9340), .ZN(n26013) );
  AOI22_X1 U2734 ( .A1(\mem[11][5] ), .A2(n9335), .B1(n27119), .B2(data_in[5]), 
        .ZN(n9340) );
  INV_X1 U2735 ( .A(n9341), .ZN(n26012) );
  AOI22_X1 U2736 ( .A1(\mem[11][6] ), .A2(n9335), .B1(n27119), .B2(data_in[6]), 
        .ZN(n9341) );
  INV_X1 U2737 ( .A(n9342), .ZN(n26011) );
  AOI22_X1 U2738 ( .A1(\mem[11][7] ), .A2(n9335), .B1(n27119), .B2(data_in[7]), 
        .ZN(n9342) );
  INV_X1 U2739 ( .A(n9344), .ZN(n26010) );
  AOI22_X1 U2740 ( .A1(\mem[12][0] ), .A2(n9345), .B1(n27118), .B2(data_in[0]), 
        .ZN(n9344) );
  INV_X1 U2741 ( .A(n9346), .ZN(n26009) );
  AOI22_X1 U2742 ( .A1(\mem[12][1] ), .A2(n9345), .B1(n27118), .B2(data_in[1]), 
        .ZN(n9346) );
  INV_X1 U2743 ( .A(n9347), .ZN(n26008) );
  AOI22_X1 U2744 ( .A1(\mem[12][2] ), .A2(n9345), .B1(n27118), .B2(data_in[2]), 
        .ZN(n9347) );
  INV_X1 U2745 ( .A(n9348), .ZN(n26007) );
  AOI22_X1 U2746 ( .A1(\mem[12][3] ), .A2(n9345), .B1(n27118), .B2(data_in[3]), 
        .ZN(n9348) );
  INV_X1 U2747 ( .A(n9349), .ZN(n26006) );
  AOI22_X1 U2748 ( .A1(\mem[12][4] ), .A2(n9345), .B1(n27118), .B2(data_in[4]), 
        .ZN(n9349) );
  INV_X1 U2749 ( .A(n9350), .ZN(n26005) );
  AOI22_X1 U2750 ( .A1(\mem[12][5] ), .A2(n9345), .B1(n27118), .B2(data_in[5]), 
        .ZN(n9350) );
  INV_X1 U2751 ( .A(n9351), .ZN(n26004) );
  AOI22_X1 U2752 ( .A1(\mem[12][6] ), .A2(n9345), .B1(n27118), .B2(data_in[6]), 
        .ZN(n9351) );
  INV_X1 U2753 ( .A(n9352), .ZN(n26003) );
  AOI22_X1 U2754 ( .A1(\mem[12][7] ), .A2(n9345), .B1(n27118), .B2(data_in[7]), 
        .ZN(n9352) );
  INV_X1 U2755 ( .A(n9354), .ZN(n26002) );
  AOI22_X1 U2756 ( .A1(\mem[13][0] ), .A2(n9355), .B1(n27117), .B2(data_in[0]), 
        .ZN(n9354) );
  INV_X1 U2757 ( .A(n9356), .ZN(n26001) );
  AOI22_X1 U2758 ( .A1(\mem[13][1] ), .A2(n9355), .B1(n27117), .B2(data_in[1]), 
        .ZN(n9356) );
  INV_X1 U2759 ( .A(n9357), .ZN(n26000) );
  AOI22_X1 U2760 ( .A1(\mem[13][2] ), .A2(n9355), .B1(n27117), .B2(data_in[2]), 
        .ZN(n9357) );
  INV_X1 U2761 ( .A(n9358), .ZN(n25999) );
  AOI22_X1 U2762 ( .A1(\mem[13][3] ), .A2(n9355), .B1(n27117), .B2(data_in[3]), 
        .ZN(n9358) );
  INV_X1 U2763 ( .A(n9359), .ZN(n25998) );
  AOI22_X1 U2764 ( .A1(\mem[13][4] ), .A2(n9355), .B1(n27117), .B2(data_in[4]), 
        .ZN(n9359) );
  INV_X1 U2765 ( .A(n9360), .ZN(n25997) );
  AOI22_X1 U2766 ( .A1(\mem[13][5] ), .A2(n9355), .B1(n27117), .B2(data_in[5]), 
        .ZN(n9360) );
  INV_X1 U2767 ( .A(n9361), .ZN(n25996) );
  AOI22_X1 U2768 ( .A1(\mem[13][6] ), .A2(n9355), .B1(n27117), .B2(data_in[6]), 
        .ZN(n9361) );
  INV_X1 U2769 ( .A(n9362), .ZN(n25995) );
  AOI22_X1 U2770 ( .A1(\mem[13][7] ), .A2(n9355), .B1(n27117), .B2(data_in[7]), 
        .ZN(n9362) );
  INV_X1 U2771 ( .A(n9364), .ZN(n25994) );
  AOI22_X1 U2772 ( .A1(\mem[14][0] ), .A2(n9365), .B1(n27116), .B2(data_in[0]), 
        .ZN(n9364) );
  INV_X1 U2773 ( .A(n9366), .ZN(n25993) );
  AOI22_X1 U2774 ( .A1(\mem[14][1] ), .A2(n9365), .B1(n27116), .B2(data_in[1]), 
        .ZN(n9366) );
  INV_X1 U2775 ( .A(n9367), .ZN(n25992) );
  AOI22_X1 U2776 ( .A1(\mem[14][2] ), .A2(n9365), .B1(n27116), .B2(data_in[2]), 
        .ZN(n9367) );
  INV_X1 U2777 ( .A(n9368), .ZN(n25991) );
  AOI22_X1 U2778 ( .A1(\mem[14][3] ), .A2(n9365), .B1(n27116), .B2(data_in[3]), 
        .ZN(n9368) );
  INV_X1 U2779 ( .A(n9369), .ZN(n25990) );
  AOI22_X1 U2780 ( .A1(\mem[14][4] ), .A2(n9365), .B1(n27116), .B2(data_in[4]), 
        .ZN(n9369) );
  INV_X1 U2781 ( .A(n9370), .ZN(n25989) );
  AOI22_X1 U2782 ( .A1(\mem[14][5] ), .A2(n9365), .B1(n27116), .B2(data_in[5]), 
        .ZN(n9370) );
  INV_X1 U2783 ( .A(n9371), .ZN(n25988) );
  AOI22_X1 U2784 ( .A1(\mem[14][6] ), .A2(n9365), .B1(n27116), .B2(data_in[6]), 
        .ZN(n9371) );
  INV_X1 U2785 ( .A(n9372), .ZN(n25987) );
  AOI22_X1 U2786 ( .A1(\mem[14][7] ), .A2(n9365), .B1(n27116), .B2(data_in[7]), 
        .ZN(n9372) );
  INV_X1 U2787 ( .A(n9374), .ZN(n25986) );
  AOI22_X1 U2788 ( .A1(\mem[15][0] ), .A2(n9375), .B1(n27115), .B2(data_in[0]), 
        .ZN(n9374) );
  INV_X1 U2789 ( .A(n9376), .ZN(n25985) );
  AOI22_X1 U2790 ( .A1(\mem[15][1] ), .A2(n9375), .B1(n27115), .B2(data_in[1]), 
        .ZN(n9376) );
  INV_X1 U2791 ( .A(n9377), .ZN(n25984) );
  AOI22_X1 U2792 ( .A1(\mem[15][2] ), .A2(n9375), .B1(n27115), .B2(data_in[2]), 
        .ZN(n9377) );
  INV_X1 U2793 ( .A(n9378), .ZN(n25983) );
  AOI22_X1 U2794 ( .A1(\mem[15][3] ), .A2(n9375), .B1(n27115), .B2(data_in[3]), 
        .ZN(n9378) );
  INV_X1 U2795 ( .A(n9379), .ZN(n25982) );
  AOI22_X1 U2796 ( .A1(\mem[15][4] ), .A2(n9375), .B1(n27115), .B2(data_in[4]), 
        .ZN(n9379) );
  INV_X1 U2797 ( .A(n9380), .ZN(n25981) );
  AOI22_X1 U2798 ( .A1(\mem[15][5] ), .A2(n9375), .B1(n27115), .B2(data_in[5]), 
        .ZN(n9380) );
  INV_X1 U2799 ( .A(n9381), .ZN(n25980) );
  AOI22_X1 U2800 ( .A1(\mem[15][6] ), .A2(n9375), .B1(n27115), .B2(data_in[6]), 
        .ZN(n9381) );
  INV_X1 U2801 ( .A(n9382), .ZN(n25979) );
  AOI22_X1 U2802 ( .A1(\mem[15][7] ), .A2(n9375), .B1(n27115), .B2(data_in[7]), 
        .ZN(n9382) );
  INV_X1 U2803 ( .A(n9384), .ZN(n25978) );
  AOI22_X1 U2804 ( .A1(\mem[16][0] ), .A2(n9385), .B1(n27114), .B2(data_in[0]), 
        .ZN(n9384) );
  INV_X1 U2805 ( .A(n9386), .ZN(n25977) );
  AOI22_X1 U2806 ( .A1(\mem[16][1] ), .A2(n9385), .B1(n27114), .B2(data_in[1]), 
        .ZN(n9386) );
  INV_X1 U2807 ( .A(n9387), .ZN(n25976) );
  AOI22_X1 U2808 ( .A1(\mem[16][2] ), .A2(n9385), .B1(n27114), .B2(data_in[2]), 
        .ZN(n9387) );
  INV_X1 U2809 ( .A(n9388), .ZN(n25975) );
  AOI22_X1 U2810 ( .A1(\mem[16][3] ), .A2(n9385), .B1(n27114), .B2(data_in[3]), 
        .ZN(n9388) );
  INV_X1 U2811 ( .A(n9389), .ZN(n25974) );
  AOI22_X1 U2812 ( .A1(\mem[16][4] ), .A2(n9385), .B1(n27114), .B2(data_in[4]), 
        .ZN(n9389) );
  INV_X1 U2813 ( .A(n9390), .ZN(n25973) );
  AOI22_X1 U2814 ( .A1(\mem[16][5] ), .A2(n9385), .B1(n27114), .B2(data_in[5]), 
        .ZN(n9390) );
  INV_X1 U2815 ( .A(n9391), .ZN(n25972) );
  AOI22_X1 U2816 ( .A1(\mem[16][6] ), .A2(n9385), .B1(n27114), .B2(data_in[6]), 
        .ZN(n9391) );
  INV_X1 U2817 ( .A(n9392), .ZN(n25971) );
  AOI22_X1 U2818 ( .A1(\mem[16][7] ), .A2(n9385), .B1(n27114), .B2(data_in[7]), 
        .ZN(n9392) );
  INV_X1 U2819 ( .A(n9394), .ZN(n25970) );
  AOI22_X1 U2820 ( .A1(\mem[17][0] ), .A2(n9395), .B1(n27113), .B2(data_in[0]), 
        .ZN(n9394) );
  INV_X1 U2821 ( .A(n9396), .ZN(n25969) );
  AOI22_X1 U2822 ( .A1(\mem[17][1] ), .A2(n9395), .B1(n27113), .B2(data_in[1]), 
        .ZN(n9396) );
  INV_X1 U2823 ( .A(n9397), .ZN(n25968) );
  AOI22_X1 U2824 ( .A1(\mem[17][2] ), .A2(n9395), .B1(n27113), .B2(data_in[2]), 
        .ZN(n9397) );
  INV_X1 U2825 ( .A(n9398), .ZN(n25967) );
  AOI22_X1 U2826 ( .A1(\mem[17][3] ), .A2(n9395), .B1(n27113), .B2(data_in[3]), 
        .ZN(n9398) );
  INV_X1 U2827 ( .A(n9399), .ZN(n25966) );
  AOI22_X1 U2828 ( .A1(\mem[17][4] ), .A2(n9395), .B1(n27113), .B2(data_in[4]), 
        .ZN(n9399) );
  INV_X1 U2829 ( .A(n9400), .ZN(n25965) );
  AOI22_X1 U2830 ( .A1(\mem[17][5] ), .A2(n9395), .B1(n27113), .B2(data_in[5]), 
        .ZN(n9400) );
  INV_X1 U2831 ( .A(n9401), .ZN(n25964) );
  AOI22_X1 U2832 ( .A1(\mem[17][6] ), .A2(n9395), .B1(n27113), .B2(data_in[6]), 
        .ZN(n9401) );
  INV_X1 U2833 ( .A(n9402), .ZN(n25963) );
  AOI22_X1 U2834 ( .A1(\mem[17][7] ), .A2(n9395), .B1(n27113), .B2(data_in[7]), 
        .ZN(n9402) );
  INV_X1 U2835 ( .A(n9404), .ZN(n25962) );
  AOI22_X1 U2836 ( .A1(\mem[18][0] ), .A2(n9405), .B1(n27112), .B2(data_in[0]), 
        .ZN(n9404) );
  INV_X1 U2837 ( .A(n9406), .ZN(n25961) );
  AOI22_X1 U2838 ( .A1(\mem[18][1] ), .A2(n9405), .B1(n27112), .B2(data_in[1]), 
        .ZN(n9406) );
  INV_X1 U2839 ( .A(n9407), .ZN(n25960) );
  AOI22_X1 U2840 ( .A1(\mem[18][2] ), .A2(n9405), .B1(n27112), .B2(data_in[2]), 
        .ZN(n9407) );
  INV_X1 U2841 ( .A(n9408), .ZN(n25959) );
  AOI22_X1 U2842 ( .A1(\mem[18][3] ), .A2(n9405), .B1(n27112), .B2(data_in[3]), 
        .ZN(n9408) );
  INV_X1 U2843 ( .A(n9409), .ZN(n25958) );
  AOI22_X1 U2844 ( .A1(\mem[18][4] ), .A2(n9405), .B1(n27112), .B2(data_in[4]), 
        .ZN(n9409) );
  INV_X1 U2845 ( .A(n9410), .ZN(n25957) );
  AOI22_X1 U2846 ( .A1(\mem[18][5] ), .A2(n9405), .B1(n27112), .B2(data_in[5]), 
        .ZN(n9410) );
  INV_X1 U2847 ( .A(n9411), .ZN(n25956) );
  AOI22_X1 U2848 ( .A1(\mem[18][6] ), .A2(n9405), .B1(n27112), .B2(data_in[6]), 
        .ZN(n9411) );
  INV_X1 U2849 ( .A(n9412), .ZN(n25955) );
  AOI22_X1 U2850 ( .A1(\mem[18][7] ), .A2(n9405), .B1(n27112), .B2(data_in[7]), 
        .ZN(n9412) );
  INV_X1 U2851 ( .A(n9414), .ZN(n25954) );
  AOI22_X1 U2852 ( .A1(\mem[19][0] ), .A2(n9415), .B1(n27111), .B2(data_in[0]), 
        .ZN(n9414) );
  INV_X1 U2853 ( .A(n9416), .ZN(n25953) );
  AOI22_X1 U2854 ( .A1(\mem[19][1] ), .A2(n9415), .B1(n27111), .B2(data_in[1]), 
        .ZN(n9416) );
  INV_X1 U2855 ( .A(n9417), .ZN(n25952) );
  AOI22_X1 U2856 ( .A1(\mem[19][2] ), .A2(n9415), .B1(n27111), .B2(data_in[2]), 
        .ZN(n9417) );
  INV_X1 U2857 ( .A(n9418), .ZN(n25951) );
  AOI22_X1 U2858 ( .A1(\mem[19][3] ), .A2(n9415), .B1(n27111), .B2(data_in[3]), 
        .ZN(n9418) );
  INV_X1 U2859 ( .A(n9419), .ZN(n25950) );
  AOI22_X1 U2860 ( .A1(\mem[19][4] ), .A2(n9415), .B1(n27111), .B2(data_in[4]), 
        .ZN(n9419) );
  INV_X1 U2861 ( .A(n9420), .ZN(n25949) );
  AOI22_X1 U2862 ( .A1(\mem[19][5] ), .A2(n9415), .B1(n27111), .B2(data_in[5]), 
        .ZN(n9420) );
  INV_X1 U2863 ( .A(n9421), .ZN(n25948) );
  AOI22_X1 U2864 ( .A1(\mem[19][6] ), .A2(n9415), .B1(n27111), .B2(data_in[6]), 
        .ZN(n9421) );
  INV_X1 U2865 ( .A(n9422), .ZN(n25947) );
  AOI22_X1 U2866 ( .A1(\mem[19][7] ), .A2(n9415), .B1(n27111), .B2(data_in[7]), 
        .ZN(n9422) );
  INV_X1 U2867 ( .A(n9424), .ZN(n25946) );
  AOI22_X1 U2868 ( .A1(\mem[20][0] ), .A2(n9425), .B1(n27110), .B2(data_in[0]), 
        .ZN(n9424) );
  INV_X1 U2869 ( .A(n9426), .ZN(n25945) );
  AOI22_X1 U2870 ( .A1(\mem[20][1] ), .A2(n9425), .B1(n27110), .B2(data_in[1]), 
        .ZN(n9426) );
  INV_X1 U2871 ( .A(n9427), .ZN(n25944) );
  AOI22_X1 U2872 ( .A1(\mem[20][2] ), .A2(n9425), .B1(n27110), .B2(data_in[2]), 
        .ZN(n9427) );
  INV_X1 U2873 ( .A(n9428), .ZN(n25943) );
  AOI22_X1 U2874 ( .A1(\mem[20][3] ), .A2(n9425), .B1(n27110), .B2(data_in[3]), 
        .ZN(n9428) );
  INV_X1 U2875 ( .A(n9429), .ZN(n25942) );
  AOI22_X1 U2876 ( .A1(\mem[20][4] ), .A2(n9425), .B1(n27110), .B2(data_in[4]), 
        .ZN(n9429) );
  INV_X1 U2877 ( .A(n9430), .ZN(n25941) );
  AOI22_X1 U2878 ( .A1(\mem[20][5] ), .A2(n9425), .B1(n27110), .B2(data_in[5]), 
        .ZN(n9430) );
  INV_X1 U2879 ( .A(n9431), .ZN(n25940) );
  AOI22_X1 U2880 ( .A1(\mem[20][6] ), .A2(n9425), .B1(n27110), .B2(data_in[6]), 
        .ZN(n9431) );
  INV_X1 U2881 ( .A(n9432), .ZN(n25939) );
  AOI22_X1 U2882 ( .A1(\mem[20][7] ), .A2(n9425), .B1(n27110), .B2(data_in[7]), 
        .ZN(n9432) );
  INV_X1 U2883 ( .A(n9434), .ZN(n25938) );
  AOI22_X1 U2884 ( .A1(\mem[21][0] ), .A2(n9435), .B1(n27109), .B2(data_in[0]), 
        .ZN(n9434) );
  INV_X1 U2885 ( .A(n9436), .ZN(n25937) );
  AOI22_X1 U2886 ( .A1(\mem[21][1] ), .A2(n9435), .B1(n27109), .B2(data_in[1]), 
        .ZN(n9436) );
  INV_X1 U2887 ( .A(n9437), .ZN(n25936) );
  AOI22_X1 U2888 ( .A1(\mem[21][2] ), .A2(n9435), .B1(n27109), .B2(data_in[2]), 
        .ZN(n9437) );
  INV_X1 U2889 ( .A(n9438), .ZN(n25935) );
  AOI22_X1 U2890 ( .A1(\mem[21][3] ), .A2(n9435), .B1(n27109), .B2(data_in[3]), 
        .ZN(n9438) );
  INV_X1 U2891 ( .A(n9439), .ZN(n25934) );
  AOI22_X1 U2892 ( .A1(\mem[21][4] ), .A2(n9435), .B1(n27109), .B2(data_in[4]), 
        .ZN(n9439) );
  INV_X1 U2893 ( .A(n9440), .ZN(n25933) );
  AOI22_X1 U2894 ( .A1(\mem[21][5] ), .A2(n9435), .B1(n27109), .B2(data_in[5]), 
        .ZN(n9440) );
  INV_X1 U2895 ( .A(n9441), .ZN(n25932) );
  AOI22_X1 U2896 ( .A1(\mem[21][6] ), .A2(n9435), .B1(n27109), .B2(data_in[6]), 
        .ZN(n9441) );
  INV_X1 U2897 ( .A(n9442), .ZN(n25931) );
  AOI22_X1 U2898 ( .A1(\mem[21][7] ), .A2(n9435), .B1(n27109), .B2(data_in[7]), 
        .ZN(n9442) );
  INV_X1 U2899 ( .A(n9444), .ZN(n25930) );
  AOI22_X1 U2900 ( .A1(\mem[22][0] ), .A2(n9445), .B1(n27108), .B2(data_in[0]), 
        .ZN(n9444) );
  INV_X1 U2901 ( .A(n9446), .ZN(n25929) );
  AOI22_X1 U2902 ( .A1(\mem[22][1] ), .A2(n9445), .B1(n27108), .B2(data_in[1]), 
        .ZN(n9446) );
  INV_X1 U2903 ( .A(n9447), .ZN(n25928) );
  AOI22_X1 U2904 ( .A1(\mem[22][2] ), .A2(n9445), .B1(n27108), .B2(data_in[2]), 
        .ZN(n9447) );
  INV_X1 U2905 ( .A(n9448), .ZN(n25927) );
  AOI22_X1 U2906 ( .A1(\mem[22][3] ), .A2(n9445), .B1(n27108), .B2(data_in[3]), 
        .ZN(n9448) );
  INV_X1 U2907 ( .A(n9449), .ZN(n25926) );
  AOI22_X1 U2908 ( .A1(\mem[22][4] ), .A2(n9445), .B1(n27108), .B2(data_in[4]), 
        .ZN(n9449) );
  INV_X1 U2909 ( .A(n9450), .ZN(n25925) );
  AOI22_X1 U2910 ( .A1(\mem[22][5] ), .A2(n9445), .B1(n27108), .B2(data_in[5]), 
        .ZN(n9450) );
  INV_X1 U2911 ( .A(n9451), .ZN(n25924) );
  AOI22_X1 U2912 ( .A1(\mem[22][6] ), .A2(n9445), .B1(n27108), .B2(data_in[6]), 
        .ZN(n9451) );
  INV_X1 U2913 ( .A(n9452), .ZN(n25923) );
  AOI22_X1 U2914 ( .A1(\mem[22][7] ), .A2(n9445), .B1(n27108), .B2(data_in[7]), 
        .ZN(n9452) );
  INV_X1 U2915 ( .A(n9454), .ZN(n25922) );
  AOI22_X1 U2916 ( .A1(\mem[23][0] ), .A2(n9455), .B1(n27107), .B2(data_in[0]), 
        .ZN(n9454) );
  INV_X1 U2917 ( .A(n9456), .ZN(n25921) );
  AOI22_X1 U2918 ( .A1(\mem[23][1] ), .A2(n9455), .B1(n27107), .B2(data_in[1]), 
        .ZN(n9456) );
  INV_X1 U2919 ( .A(n9457), .ZN(n25920) );
  AOI22_X1 U2920 ( .A1(\mem[23][2] ), .A2(n9455), .B1(n27107), .B2(data_in[2]), 
        .ZN(n9457) );
  INV_X1 U2921 ( .A(n9458), .ZN(n25919) );
  AOI22_X1 U2922 ( .A1(\mem[23][3] ), .A2(n9455), .B1(n27107), .B2(data_in[3]), 
        .ZN(n9458) );
  INV_X1 U2923 ( .A(n9459), .ZN(n25918) );
  AOI22_X1 U2924 ( .A1(\mem[23][4] ), .A2(n9455), .B1(n27107), .B2(data_in[4]), 
        .ZN(n9459) );
  INV_X1 U2925 ( .A(n9460), .ZN(n25917) );
  AOI22_X1 U2926 ( .A1(\mem[23][5] ), .A2(n9455), .B1(n27107), .B2(data_in[5]), 
        .ZN(n9460) );
  INV_X1 U2927 ( .A(n9461), .ZN(n25916) );
  AOI22_X1 U2928 ( .A1(\mem[23][6] ), .A2(n9455), .B1(n27107), .B2(data_in[6]), 
        .ZN(n9461) );
  INV_X1 U2929 ( .A(n9462), .ZN(n25915) );
  AOI22_X1 U2930 ( .A1(\mem[23][7] ), .A2(n9455), .B1(n27107), .B2(data_in[7]), 
        .ZN(n9462) );
  INV_X1 U2931 ( .A(n9464), .ZN(n25914) );
  AOI22_X1 U2932 ( .A1(\mem[24][0] ), .A2(n9465), .B1(n27106), .B2(data_in[0]), 
        .ZN(n9464) );
  INV_X1 U2933 ( .A(n9466), .ZN(n25913) );
  AOI22_X1 U2934 ( .A1(\mem[24][1] ), .A2(n9465), .B1(n27106), .B2(data_in[1]), 
        .ZN(n9466) );
  INV_X1 U2935 ( .A(n9467), .ZN(n25912) );
  AOI22_X1 U2936 ( .A1(\mem[24][2] ), .A2(n9465), .B1(n27106), .B2(data_in[2]), 
        .ZN(n9467) );
  INV_X1 U2937 ( .A(n9468), .ZN(n25911) );
  AOI22_X1 U2938 ( .A1(\mem[24][3] ), .A2(n9465), .B1(n27106), .B2(data_in[3]), 
        .ZN(n9468) );
  INV_X1 U2939 ( .A(n9469), .ZN(n25910) );
  AOI22_X1 U2940 ( .A1(\mem[24][4] ), .A2(n9465), .B1(n27106), .B2(data_in[4]), 
        .ZN(n9469) );
  INV_X1 U2941 ( .A(n9470), .ZN(n25909) );
  AOI22_X1 U2942 ( .A1(\mem[24][5] ), .A2(n9465), .B1(n27106), .B2(data_in[5]), 
        .ZN(n9470) );
  INV_X1 U2943 ( .A(n9471), .ZN(n25908) );
  AOI22_X1 U2944 ( .A1(\mem[24][6] ), .A2(n9465), .B1(n27106), .B2(data_in[6]), 
        .ZN(n9471) );
  INV_X1 U2945 ( .A(n9472), .ZN(n25907) );
  AOI22_X1 U2946 ( .A1(\mem[24][7] ), .A2(n9465), .B1(n27106), .B2(data_in[7]), 
        .ZN(n9472) );
  INV_X1 U2947 ( .A(n9474), .ZN(n25906) );
  AOI22_X1 U2948 ( .A1(\mem[25][0] ), .A2(n9475), .B1(n27105), .B2(data_in[0]), 
        .ZN(n9474) );
  INV_X1 U2949 ( .A(n9476), .ZN(n25905) );
  AOI22_X1 U2950 ( .A1(\mem[25][1] ), .A2(n9475), .B1(n27105), .B2(data_in[1]), 
        .ZN(n9476) );
  INV_X1 U2951 ( .A(n9477), .ZN(n25904) );
  AOI22_X1 U2952 ( .A1(\mem[25][2] ), .A2(n9475), .B1(n27105), .B2(data_in[2]), 
        .ZN(n9477) );
  INV_X1 U2953 ( .A(n9478), .ZN(n25903) );
  AOI22_X1 U2954 ( .A1(\mem[25][3] ), .A2(n9475), .B1(n27105), .B2(data_in[3]), 
        .ZN(n9478) );
  INV_X1 U2955 ( .A(n9479), .ZN(n25902) );
  AOI22_X1 U2956 ( .A1(\mem[25][4] ), .A2(n9475), .B1(n27105), .B2(data_in[4]), 
        .ZN(n9479) );
  INV_X1 U2957 ( .A(n9480), .ZN(n25901) );
  AOI22_X1 U2958 ( .A1(\mem[25][5] ), .A2(n9475), .B1(n27105), .B2(data_in[5]), 
        .ZN(n9480) );
  INV_X1 U2959 ( .A(n9481), .ZN(n25900) );
  AOI22_X1 U2960 ( .A1(\mem[25][6] ), .A2(n9475), .B1(n27105), .B2(data_in[6]), 
        .ZN(n9481) );
  INV_X1 U2961 ( .A(n9482), .ZN(n25899) );
  AOI22_X1 U2962 ( .A1(\mem[25][7] ), .A2(n9475), .B1(n27105), .B2(data_in[7]), 
        .ZN(n9482) );
  INV_X1 U2963 ( .A(n9484), .ZN(n25898) );
  AOI22_X1 U2964 ( .A1(\mem[26][0] ), .A2(n9485), .B1(n27104), .B2(data_in[0]), 
        .ZN(n9484) );
  INV_X1 U2965 ( .A(n9486), .ZN(n25897) );
  AOI22_X1 U2966 ( .A1(\mem[26][1] ), .A2(n9485), .B1(n27104), .B2(data_in[1]), 
        .ZN(n9486) );
  INV_X1 U2967 ( .A(n9487), .ZN(n25896) );
  AOI22_X1 U2968 ( .A1(\mem[26][2] ), .A2(n9485), .B1(n27104), .B2(data_in[2]), 
        .ZN(n9487) );
  INV_X1 U2969 ( .A(n9488), .ZN(n25895) );
  AOI22_X1 U2970 ( .A1(\mem[26][3] ), .A2(n9485), .B1(n27104), .B2(data_in[3]), 
        .ZN(n9488) );
  INV_X1 U2971 ( .A(n9489), .ZN(n25894) );
  AOI22_X1 U2972 ( .A1(\mem[26][4] ), .A2(n9485), .B1(n27104), .B2(data_in[4]), 
        .ZN(n9489) );
  INV_X1 U2973 ( .A(n9490), .ZN(n25893) );
  AOI22_X1 U2974 ( .A1(\mem[26][5] ), .A2(n9485), .B1(n27104), .B2(data_in[5]), 
        .ZN(n9490) );
  INV_X1 U2975 ( .A(n9491), .ZN(n25892) );
  AOI22_X1 U2976 ( .A1(\mem[26][6] ), .A2(n9485), .B1(n27104), .B2(data_in[6]), 
        .ZN(n9491) );
  INV_X1 U2977 ( .A(n9492), .ZN(n25891) );
  AOI22_X1 U2978 ( .A1(\mem[26][7] ), .A2(n9485), .B1(n27104), .B2(data_in[7]), 
        .ZN(n9492) );
  INV_X1 U2979 ( .A(n9494), .ZN(n25890) );
  AOI22_X1 U2980 ( .A1(\mem[27][0] ), .A2(n9495), .B1(n27103), .B2(data_in[0]), 
        .ZN(n9494) );
  INV_X1 U2981 ( .A(n9496), .ZN(n25889) );
  AOI22_X1 U2982 ( .A1(\mem[27][1] ), .A2(n9495), .B1(n27103), .B2(data_in[1]), 
        .ZN(n9496) );
  INV_X1 U2983 ( .A(n9497), .ZN(n25888) );
  AOI22_X1 U2984 ( .A1(\mem[27][2] ), .A2(n9495), .B1(n27103), .B2(data_in[2]), 
        .ZN(n9497) );
  INV_X1 U2985 ( .A(n9498), .ZN(n25887) );
  AOI22_X1 U2986 ( .A1(\mem[27][3] ), .A2(n9495), .B1(n27103), .B2(data_in[3]), 
        .ZN(n9498) );
  INV_X1 U2987 ( .A(n9499), .ZN(n25886) );
  AOI22_X1 U2988 ( .A1(\mem[27][4] ), .A2(n9495), .B1(n27103), .B2(data_in[4]), 
        .ZN(n9499) );
  INV_X1 U2989 ( .A(n9500), .ZN(n25885) );
  AOI22_X1 U2990 ( .A1(\mem[27][5] ), .A2(n9495), .B1(n27103), .B2(data_in[5]), 
        .ZN(n9500) );
  INV_X1 U2991 ( .A(n9501), .ZN(n25884) );
  AOI22_X1 U2992 ( .A1(\mem[27][6] ), .A2(n9495), .B1(n27103), .B2(data_in[6]), 
        .ZN(n9501) );
  INV_X1 U2993 ( .A(n9502), .ZN(n25883) );
  AOI22_X1 U2994 ( .A1(\mem[27][7] ), .A2(n9495), .B1(n27103), .B2(data_in[7]), 
        .ZN(n9502) );
  INV_X1 U2995 ( .A(n9504), .ZN(n25882) );
  AOI22_X1 U2996 ( .A1(\mem[28][0] ), .A2(n9505), .B1(n27102), .B2(data_in[0]), 
        .ZN(n9504) );
  INV_X1 U2997 ( .A(n9506), .ZN(n25881) );
  AOI22_X1 U2998 ( .A1(\mem[28][1] ), .A2(n9505), .B1(n27102), .B2(data_in[1]), 
        .ZN(n9506) );
  INV_X1 U2999 ( .A(n9507), .ZN(n25880) );
  AOI22_X1 U3000 ( .A1(\mem[28][2] ), .A2(n9505), .B1(n27102), .B2(data_in[2]), 
        .ZN(n9507) );
  INV_X1 U3001 ( .A(n9508), .ZN(n25879) );
  AOI22_X1 U3002 ( .A1(\mem[28][3] ), .A2(n9505), .B1(n27102), .B2(data_in[3]), 
        .ZN(n9508) );
  INV_X1 U3003 ( .A(n9509), .ZN(n25878) );
  AOI22_X1 U3004 ( .A1(\mem[28][4] ), .A2(n9505), .B1(n27102), .B2(data_in[4]), 
        .ZN(n9509) );
  INV_X1 U3005 ( .A(n9510), .ZN(n25877) );
  AOI22_X1 U3006 ( .A1(\mem[28][5] ), .A2(n9505), .B1(n27102), .B2(data_in[5]), 
        .ZN(n9510) );
  INV_X1 U3007 ( .A(n9511), .ZN(n25876) );
  AOI22_X1 U3008 ( .A1(\mem[28][6] ), .A2(n9505), .B1(n27102), .B2(data_in[6]), 
        .ZN(n9511) );
  INV_X1 U3009 ( .A(n9512), .ZN(n25875) );
  AOI22_X1 U3010 ( .A1(\mem[28][7] ), .A2(n9505), .B1(n27102), .B2(data_in[7]), 
        .ZN(n9512) );
  INV_X1 U3011 ( .A(n9514), .ZN(n25874) );
  AOI22_X1 U3012 ( .A1(\mem[29][0] ), .A2(n9515), .B1(n27101), .B2(data_in[0]), 
        .ZN(n9514) );
  INV_X1 U3013 ( .A(n9516), .ZN(n25873) );
  AOI22_X1 U3014 ( .A1(\mem[29][1] ), .A2(n9515), .B1(n27101), .B2(data_in[1]), 
        .ZN(n9516) );
  INV_X1 U3015 ( .A(n9517), .ZN(n25872) );
  AOI22_X1 U3016 ( .A1(\mem[29][2] ), .A2(n9515), .B1(n27101), .B2(data_in[2]), 
        .ZN(n9517) );
  INV_X1 U3017 ( .A(n9518), .ZN(n25871) );
  AOI22_X1 U3018 ( .A1(\mem[29][3] ), .A2(n9515), .B1(n27101), .B2(data_in[3]), 
        .ZN(n9518) );
  INV_X1 U3019 ( .A(n9519), .ZN(n25870) );
  AOI22_X1 U3020 ( .A1(\mem[29][4] ), .A2(n9515), .B1(n27101), .B2(data_in[4]), 
        .ZN(n9519) );
  INV_X1 U3021 ( .A(n9520), .ZN(n25869) );
  AOI22_X1 U3022 ( .A1(\mem[29][5] ), .A2(n9515), .B1(n27101), .B2(data_in[5]), 
        .ZN(n9520) );
  INV_X1 U3023 ( .A(n9521), .ZN(n25868) );
  AOI22_X1 U3024 ( .A1(\mem[29][6] ), .A2(n9515), .B1(n27101), .B2(data_in[6]), 
        .ZN(n9521) );
  INV_X1 U3025 ( .A(n9522), .ZN(n25867) );
  AOI22_X1 U3026 ( .A1(\mem[29][7] ), .A2(n9515), .B1(n27101), .B2(data_in[7]), 
        .ZN(n9522) );
  INV_X1 U3027 ( .A(n9524), .ZN(n25866) );
  AOI22_X1 U3028 ( .A1(\mem[30][0] ), .A2(n9525), .B1(n27100), .B2(data_in[0]), 
        .ZN(n9524) );
  INV_X1 U3029 ( .A(n9526), .ZN(n25865) );
  AOI22_X1 U3030 ( .A1(\mem[30][1] ), .A2(n9525), .B1(n27100), .B2(data_in[1]), 
        .ZN(n9526) );
  INV_X1 U3031 ( .A(n9527), .ZN(n25864) );
  AOI22_X1 U3032 ( .A1(\mem[30][2] ), .A2(n9525), .B1(n27100), .B2(data_in[2]), 
        .ZN(n9527) );
  INV_X1 U3033 ( .A(n9528), .ZN(n25863) );
  AOI22_X1 U3034 ( .A1(\mem[30][3] ), .A2(n9525), .B1(n27100), .B2(data_in[3]), 
        .ZN(n9528) );
  INV_X1 U3035 ( .A(n9529), .ZN(n25862) );
  AOI22_X1 U3036 ( .A1(\mem[30][4] ), .A2(n9525), .B1(n27100), .B2(data_in[4]), 
        .ZN(n9529) );
  INV_X1 U3037 ( .A(n9530), .ZN(n25861) );
  AOI22_X1 U3038 ( .A1(\mem[30][5] ), .A2(n9525), .B1(n27100), .B2(data_in[5]), 
        .ZN(n9530) );
  INV_X1 U3039 ( .A(n9531), .ZN(n25860) );
  AOI22_X1 U3040 ( .A1(\mem[30][6] ), .A2(n9525), .B1(n27100), .B2(data_in[6]), 
        .ZN(n9531) );
  INV_X1 U3041 ( .A(n9532), .ZN(n25859) );
  AOI22_X1 U3042 ( .A1(\mem[30][7] ), .A2(n9525), .B1(n27100), .B2(data_in[7]), 
        .ZN(n9532) );
  INV_X1 U3043 ( .A(n9534), .ZN(n25858) );
  AOI22_X1 U3044 ( .A1(\mem[31][0] ), .A2(n9535), .B1(n27099), .B2(data_in[0]), 
        .ZN(n9534) );
  INV_X1 U3045 ( .A(n9536), .ZN(n25857) );
  AOI22_X1 U3046 ( .A1(\mem[31][1] ), .A2(n9535), .B1(n27099), .B2(data_in[1]), 
        .ZN(n9536) );
  INV_X1 U3047 ( .A(n9537), .ZN(n25856) );
  AOI22_X1 U3048 ( .A1(\mem[31][2] ), .A2(n9535), .B1(n27099), .B2(data_in[2]), 
        .ZN(n9537) );
  INV_X1 U3049 ( .A(n9538), .ZN(n25855) );
  AOI22_X1 U3050 ( .A1(\mem[31][3] ), .A2(n9535), .B1(n27099), .B2(data_in[3]), 
        .ZN(n9538) );
  INV_X1 U3051 ( .A(n9539), .ZN(n25854) );
  AOI22_X1 U3052 ( .A1(\mem[31][4] ), .A2(n9535), .B1(n27099), .B2(data_in[4]), 
        .ZN(n9539) );
  INV_X1 U3053 ( .A(n9540), .ZN(n25853) );
  AOI22_X1 U3054 ( .A1(\mem[31][5] ), .A2(n9535), .B1(n27099), .B2(data_in[5]), 
        .ZN(n9540) );
  INV_X1 U3055 ( .A(n9541), .ZN(n25852) );
  AOI22_X1 U3056 ( .A1(\mem[31][6] ), .A2(n9535), .B1(n27099), .B2(data_in[6]), 
        .ZN(n9541) );
  INV_X1 U3057 ( .A(n9542), .ZN(n25851) );
  AOI22_X1 U3058 ( .A1(\mem[31][7] ), .A2(n9535), .B1(n27099), .B2(data_in[7]), 
        .ZN(n9542) );
  INV_X1 U3059 ( .A(n9620), .ZN(n25786) );
  AOI22_X1 U3060 ( .A1(\mem[40][0] ), .A2(n9621), .B1(n27090), .B2(data_in[0]), 
        .ZN(n9620) );
  INV_X1 U3061 ( .A(n9622), .ZN(n25785) );
  AOI22_X1 U3062 ( .A1(\mem[40][1] ), .A2(n9621), .B1(n27090), .B2(data_in[1]), 
        .ZN(n9622) );
  INV_X1 U3063 ( .A(n9623), .ZN(n25784) );
  AOI22_X1 U3064 ( .A1(\mem[40][2] ), .A2(n9621), .B1(n27090), .B2(data_in[2]), 
        .ZN(n9623) );
  INV_X1 U3065 ( .A(n9624), .ZN(n25783) );
  AOI22_X1 U3066 ( .A1(\mem[40][3] ), .A2(n9621), .B1(n27090), .B2(data_in[3]), 
        .ZN(n9624) );
  INV_X1 U3067 ( .A(n9625), .ZN(n25782) );
  AOI22_X1 U3068 ( .A1(\mem[40][4] ), .A2(n9621), .B1(n27090), .B2(data_in[4]), 
        .ZN(n9625) );
  INV_X1 U3069 ( .A(n9626), .ZN(n25781) );
  AOI22_X1 U3070 ( .A1(\mem[40][5] ), .A2(n9621), .B1(n27090), .B2(data_in[5]), 
        .ZN(n9626) );
  INV_X1 U3071 ( .A(n9627), .ZN(n25780) );
  AOI22_X1 U3072 ( .A1(\mem[40][6] ), .A2(n9621), .B1(n27090), .B2(data_in[6]), 
        .ZN(n9627) );
  INV_X1 U3073 ( .A(n9628), .ZN(n25779) );
  AOI22_X1 U3074 ( .A1(\mem[40][7] ), .A2(n9621), .B1(n27090), .B2(data_in[7]), 
        .ZN(n9628) );
  INV_X1 U3075 ( .A(n9629), .ZN(n25778) );
  AOI22_X1 U3076 ( .A1(\mem[41][0] ), .A2(n9630), .B1(n27089), .B2(data_in[0]), 
        .ZN(n9629) );
  INV_X1 U3077 ( .A(n9631), .ZN(n25777) );
  AOI22_X1 U3078 ( .A1(\mem[41][1] ), .A2(n9630), .B1(n27089), .B2(data_in[1]), 
        .ZN(n9631) );
  INV_X1 U3079 ( .A(n9632), .ZN(n25776) );
  AOI22_X1 U3080 ( .A1(\mem[41][2] ), .A2(n9630), .B1(n27089), .B2(data_in[2]), 
        .ZN(n9632) );
  INV_X1 U3081 ( .A(n9633), .ZN(n25775) );
  AOI22_X1 U3082 ( .A1(\mem[41][3] ), .A2(n9630), .B1(n27089), .B2(data_in[3]), 
        .ZN(n9633) );
  INV_X1 U3083 ( .A(n9634), .ZN(n25774) );
  AOI22_X1 U3084 ( .A1(\mem[41][4] ), .A2(n9630), .B1(n27089), .B2(data_in[4]), 
        .ZN(n9634) );
  INV_X1 U3085 ( .A(n9635), .ZN(n25773) );
  AOI22_X1 U3086 ( .A1(\mem[41][5] ), .A2(n9630), .B1(n27089), .B2(data_in[5]), 
        .ZN(n9635) );
  INV_X1 U3087 ( .A(n9636), .ZN(n25772) );
  AOI22_X1 U3088 ( .A1(\mem[41][6] ), .A2(n9630), .B1(n27089), .B2(data_in[6]), 
        .ZN(n9636) );
  INV_X1 U3089 ( .A(n9637), .ZN(n25771) );
  AOI22_X1 U3090 ( .A1(\mem[41][7] ), .A2(n9630), .B1(n27089), .B2(data_in[7]), 
        .ZN(n9637) );
  INV_X1 U3091 ( .A(n9638), .ZN(n25770) );
  AOI22_X1 U3092 ( .A1(\mem[42][0] ), .A2(n9639), .B1(n27088), .B2(data_in[0]), 
        .ZN(n9638) );
  INV_X1 U3093 ( .A(n9640), .ZN(n25769) );
  AOI22_X1 U3094 ( .A1(\mem[42][1] ), .A2(n9639), .B1(n27088), .B2(data_in[1]), 
        .ZN(n9640) );
  INV_X1 U3095 ( .A(n9641), .ZN(n25768) );
  AOI22_X1 U3096 ( .A1(\mem[42][2] ), .A2(n9639), .B1(n27088), .B2(data_in[2]), 
        .ZN(n9641) );
  INV_X1 U3097 ( .A(n9642), .ZN(n25767) );
  AOI22_X1 U3098 ( .A1(\mem[42][3] ), .A2(n9639), .B1(n27088), .B2(data_in[3]), 
        .ZN(n9642) );
  INV_X1 U3099 ( .A(n9643), .ZN(n25766) );
  AOI22_X1 U3100 ( .A1(\mem[42][4] ), .A2(n9639), .B1(n27088), .B2(data_in[4]), 
        .ZN(n9643) );
  INV_X1 U3101 ( .A(n9644), .ZN(n25765) );
  AOI22_X1 U3102 ( .A1(\mem[42][5] ), .A2(n9639), .B1(n27088), .B2(data_in[5]), 
        .ZN(n9644) );
  INV_X1 U3103 ( .A(n9645), .ZN(n25764) );
  AOI22_X1 U3104 ( .A1(\mem[42][6] ), .A2(n9639), .B1(n27088), .B2(data_in[6]), 
        .ZN(n9645) );
  INV_X1 U3105 ( .A(n9646), .ZN(n25763) );
  AOI22_X1 U3106 ( .A1(\mem[42][7] ), .A2(n9639), .B1(n27088), .B2(data_in[7]), 
        .ZN(n9646) );
  INV_X1 U3107 ( .A(n9647), .ZN(n25762) );
  AOI22_X1 U3108 ( .A1(\mem[43][0] ), .A2(n9648), .B1(n27087), .B2(data_in[0]), 
        .ZN(n9647) );
  INV_X1 U3109 ( .A(n9649), .ZN(n25761) );
  AOI22_X1 U3110 ( .A1(\mem[43][1] ), .A2(n9648), .B1(n27087), .B2(data_in[1]), 
        .ZN(n9649) );
  INV_X1 U3111 ( .A(n9650), .ZN(n25760) );
  AOI22_X1 U3112 ( .A1(\mem[43][2] ), .A2(n9648), .B1(n27087), .B2(data_in[2]), 
        .ZN(n9650) );
  INV_X1 U3113 ( .A(n9651), .ZN(n25759) );
  AOI22_X1 U3114 ( .A1(\mem[43][3] ), .A2(n9648), .B1(n27087), .B2(data_in[3]), 
        .ZN(n9651) );
  INV_X1 U3115 ( .A(n9652), .ZN(n25758) );
  AOI22_X1 U3116 ( .A1(\mem[43][4] ), .A2(n9648), .B1(n27087), .B2(data_in[4]), 
        .ZN(n9652) );
  INV_X1 U3117 ( .A(n9653), .ZN(n25757) );
  AOI22_X1 U3118 ( .A1(\mem[43][5] ), .A2(n9648), .B1(n27087), .B2(data_in[5]), 
        .ZN(n9653) );
  INV_X1 U3119 ( .A(n9654), .ZN(n25756) );
  AOI22_X1 U3120 ( .A1(\mem[43][6] ), .A2(n9648), .B1(n27087), .B2(data_in[6]), 
        .ZN(n9654) );
  INV_X1 U3121 ( .A(n9655), .ZN(n25755) );
  AOI22_X1 U3122 ( .A1(\mem[43][7] ), .A2(n9648), .B1(n27087), .B2(data_in[7]), 
        .ZN(n9655) );
  INV_X1 U3123 ( .A(n9656), .ZN(n25754) );
  AOI22_X1 U3124 ( .A1(\mem[44][0] ), .A2(n9657), .B1(n27086), .B2(data_in[0]), 
        .ZN(n9656) );
  INV_X1 U3125 ( .A(n9658), .ZN(n25753) );
  AOI22_X1 U3126 ( .A1(\mem[44][1] ), .A2(n9657), .B1(n27086), .B2(data_in[1]), 
        .ZN(n9658) );
  INV_X1 U3127 ( .A(n9659), .ZN(n25752) );
  AOI22_X1 U3128 ( .A1(\mem[44][2] ), .A2(n9657), .B1(n27086), .B2(data_in[2]), 
        .ZN(n9659) );
  INV_X1 U3129 ( .A(n9660), .ZN(n25751) );
  AOI22_X1 U3130 ( .A1(\mem[44][3] ), .A2(n9657), .B1(n27086), .B2(data_in[3]), 
        .ZN(n9660) );
  INV_X1 U3131 ( .A(n9661), .ZN(n25750) );
  AOI22_X1 U3132 ( .A1(\mem[44][4] ), .A2(n9657), .B1(n27086), .B2(data_in[4]), 
        .ZN(n9661) );
  INV_X1 U3133 ( .A(n9662), .ZN(n25749) );
  AOI22_X1 U3134 ( .A1(\mem[44][5] ), .A2(n9657), .B1(n27086), .B2(data_in[5]), 
        .ZN(n9662) );
  INV_X1 U3135 ( .A(n9663), .ZN(n25748) );
  AOI22_X1 U3136 ( .A1(\mem[44][6] ), .A2(n9657), .B1(n27086), .B2(data_in[6]), 
        .ZN(n9663) );
  INV_X1 U3137 ( .A(n9664), .ZN(n25747) );
  AOI22_X1 U3138 ( .A1(\mem[44][7] ), .A2(n9657), .B1(n27086), .B2(data_in[7]), 
        .ZN(n9664) );
  INV_X1 U3139 ( .A(n9665), .ZN(n25746) );
  AOI22_X1 U3140 ( .A1(\mem[45][0] ), .A2(n9666), .B1(n27085), .B2(data_in[0]), 
        .ZN(n9665) );
  INV_X1 U3141 ( .A(n9667), .ZN(n25745) );
  AOI22_X1 U3142 ( .A1(\mem[45][1] ), .A2(n9666), .B1(n27085), .B2(data_in[1]), 
        .ZN(n9667) );
  INV_X1 U3143 ( .A(n9668), .ZN(n25744) );
  AOI22_X1 U3144 ( .A1(\mem[45][2] ), .A2(n9666), .B1(n27085), .B2(data_in[2]), 
        .ZN(n9668) );
  INV_X1 U3145 ( .A(n9669), .ZN(n25743) );
  AOI22_X1 U3146 ( .A1(\mem[45][3] ), .A2(n9666), .B1(n27085), .B2(data_in[3]), 
        .ZN(n9669) );
  INV_X1 U3147 ( .A(n9670), .ZN(n25742) );
  AOI22_X1 U3148 ( .A1(\mem[45][4] ), .A2(n9666), .B1(n27085), .B2(data_in[4]), 
        .ZN(n9670) );
  INV_X1 U3149 ( .A(n9671), .ZN(n25741) );
  AOI22_X1 U3150 ( .A1(\mem[45][5] ), .A2(n9666), .B1(n27085), .B2(data_in[5]), 
        .ZN(n9671) );
  INV_X1 U3151 ( .A(n9672), .ZN(n25740) );
  AOI22_X1 U3152 ( .A1(\mem[45][6] ), .A2(n9666), .B1(n27085), .B2(data_in[6]), 
        .ZN(n9672) );
  INV_X1 U3153 ( .A(n9673), .ZN(n25739) );
  AOI22_X1 U3154 ( .A1(\mem[45][7] ), .A2(n9666), .B1(n27085), .B2(data_in[7]), 
        .ZN(n9673) );
  INV_X1 U3155 ( .A(n9674), .ZN(n25738) );
  AOI22_X1 U3156 ( .A1(\mem[46][0] ), .A2(n9675), .B1(n27084), .B2(data_in[0]), 
        .ZN(n9674) );
  INV_X1 U3157 ( .A(n9676), .ZN(n25737) );
  AOI22_X1 U3158 ( .A1(\mem[46][1] ), .A2(n9675), .B1(n27084), .B2(data_in[1]), 
        .ZN(n9676) );
  INV_X1 U3159 ( .A(n9677), .ZN(n25736) );
  AOI22_X1 U3160 ( .A1(\mem[46][2] ), .A2(n9675), .B1(n27084), .B2(data_in[2]), 
        .ZN(n9677) );
  INV_X1 U3161 ( .A(n9678), .ZN(n25735) );
  AOI22_X1 U3162 ( .A1(\mem[46][3] ), .A2(n9675), .B1(n27084), .B2(data_in[3]), 
        .ZN(n9678) );
  INV_X1 U3163 ( .A(n9679), .ZN(n25734) );
  AOI22_X1 U3164 ( .A1(\mem[46][4] ), .A2(n9675), .B1(n27084), .B2(data_in[4]), 
        .ZN(n9679) );
  INV_X1 U3165 ( .A(n9680), .ZN(n25733) );
  AOI22_X1 U3166 ( .A1(\mem[46][5] ), .A2(n9675), .B1(n27084), .B2(data_in[5]), 
        .ZN(n9680) );
  INV_X1 U3167 ( .A(n9681), .ZN(n25732) );
  AOI22_X1 U3168 ( .A1(\mem[46][6] ), .A2(n9675), .B1(n27084), .B2(data_in[6]), 
        .ZN(n9681) );
  INV_X1 U3169 ( .A(n9682), .ZN(n25731) );
  AOI22_X1 U3170 ( .A1(\mem[46][7] ), .A2(n9675), .B1(n27084), .B2(data_in[7]), 
        .ZN(n9682) );
  INV_X1 U3171 ( .A(n9683), .ZN(n25730) );
  AOI22_X1 U3172 ( .A1(\mem[47][0] ), .A2(n9684), .B1(n27083), .B2(data_in[0]), 
        .ZN(n9683) );
  INV_X1 U3173 ( .A(n9685), .ZN(n25729) );
  AOI22_X1 U3174 ( .A1(\mem[47][1] ), .A2(n9684), .B1(n27083), .B2(data_in[1]), 
        .ZN(n9685) );
  INV_X1 U3175 ( .A(n9686), .ZN(n25728) );
  AOI22_X1 U3176 ( .A1(\mem[47][2] ), .A2(n9684), .B1(n27083), .B2(data_in[2]), 
        .ZN(n9686) );
  INV_X1 U3177 ( .A(n9687), .ZN(n25727) );
  AOI22_X1 U3178 ( .A1(\mem[47][3] ), .A2(n9684), .B1(n27083), .B2(data_in[3]), 
        .ZN(n9687) );
  INV_X1 U3179 ( .A(n9688), .ZN(n25726) );
  AOI22_X1 U3180 ( .A1(\mem[47][4] ), .A2(n9684), .B1(n27083), .B2(data_in[4]), 
        .ZN(n9688) );
  INV_X1 U3181 ( .A(n9689), .ZN(n25725) );
  AOI22_X1 U3182 ( .A1(\mem[47][5] ), .A2(n9684), .B1(n27083), .B2(data_in[5]), 
        .ZN(n9689) );
  INV_X1 U3183 ( .A(n9690), .ZN(n25724) );
  AOI22_X1 U3184 ( .A1(\mem[47][6] ), .A2(n9684), .B1(n27083), .B2(data_in[6]), 
        .ZN(n9690) );
  INV_X1 U3185 ( .A(n9691), .ZN(n25723) );
  AOI22_X1 U3186 ( .A1(\mem[47][7] ), .A2(n9684), .B1(n27083), .B2(data_in[7]), 
        .ZN(n9691) );
  INV_X1 U3187 ( .A(n9692), .ZN(n25722) );
  AOI22_X1 U3188 ( .A1(\mem[48][0] ), .A2(n9693), .B1(n27082), .B2(data_in[0]), 
        .ZN(n9692) );
  INV_X1 U3189 ( .A(n9694), .ZN(n25721) );
  AOI22_X1 U3190 ( .A1(\mem[48][1] ), .A2(n9693), .B1(n27082), .B2(data_in[1]), 
        .ZN(n9694) );
  INV_X1 U3191 ( .A(n9695), .ZN(n25720) );
  AOI22_X1 U3192 ( .A1(\mem[48][2] ), .A2(n9693), .B1(n27082), .B2(data_in[2]), 
        .ZN(n9695) );
  INV_X1 U3193 ( .A(n9696), .ZN(n25719) );
  AOI22_X1 U3194 ( .A1(\mem[48][3] ), .A2(n9693), .B1(n27082), .B2(data_in[3]), 
        .ZN(n9696) );
  INV_X1 U3195 ( .A(n9697), .ZN(n25718) );
  AOI22_X1 U3196 ( .A1(\mem[48][4] ), .A2(n9693), .B1(n27082), .B2(data_in[4]), 
        .ZN(n9697) );
  INV_X1 U3197 ( .A(n9698), .ZN(n25717) );
  AOI22_X1 U3198 ( .A1(\mem[48][5] ), .A2(n9693), .B1(n27082), .B2(data_in[5]), 
        .ZN(n9698) );
  INV_X1 U3199 ( .A(n9699), .ZN(n25716) );
  AOI22_X1 U3200 ( .A1(\mem[48][6] ), .A2(n9693), .B1(n27082), .B2(data_in[6]), 
        .ZN(n9699) );
  INV_X1 U3201 ( .A(n9700), .ZN(n25715) );
  AOI22_X1 U3202 ( .A1(\mem[48][7] ), .A2(n9693), .B1(n27082), .B2(data_in[7]), 
        .ZN(n9700) );
  INV_X1 U3203 ( .A(n9701), .ZN(n25714) );
  AOI22_X1 U3204 ( .A1(\mem[49][0] ), .A2(n9702), .B1(n27081), .B2(data_in[0]), 
        .ZN(n9701) );
  INV_X1 U3205 ( .A(n9703), .ZN(n25713) );
  AOI22_X1 U3206 ( .A1(\mem[49][1] ), .A2(n9702), .B1(n27081), .B2(data_in[1]), 
        .ZN(n9703) );
  INV_X1 U3207 ( .A(n9704), .ZN(n25712) );
  AOI22_X1 U3208 ( .A1(\mem[49][2] ), .A2(n9702), .B1(n27081), .B2(data_in[2]), 
        .ZN(n9704) );
  INV_X1 U3209 ( .A(n9705), .ZN(n25711) );
  AOI22_X1 U3210 ( .A1(\mem[49][3] ), .A2(n9702), .B1(n27081), .B2(data_in[3]), 
        .ZN(n9705) );
  INV_X1 U3211 ( .A(n9706), .ZN(n25710) );
  AOI22_X1 U3212 ( .A1(\mem[49][4] ), .A2(n9702), .B1(n27081), .B2(data_in[4]), 
        .ZN(n9706) );
  INV_X1 U3213 ( .A(n9707), .ZN(n25709) );
  AOI22_X1 U3214 ( .A1(\mem[49][5] ), .A2(n9702), .B1(n27081), .B2(data_in[5]), 
        .ZN(n9707) );
  INV_X1 U3215 ( .A(n9708), .ZN(n25708) );
  AOI22_X1 U3216 ( .A1(\mem[49][6] ), .A2(n9702), .B1(n27081), .B2(data_in[6]), 
        .ZN(n9708) );
  INV_X1 U3217 ( .A(n9709), .ZN(n25707) );
  AOI22_X1 U3218 ( .A1(\mem[49][7] ), .A2(n9702), .B1(n27081), .B2(data_in[7]), 
        .ZN(n9709) );
  INV_X1 U3219 ( .A(n9710), .ZN(n25706) );
  AOI22_X1 U3220 ( .A1(\mem[50][0] ), .A2(n9711), .B1(n27080), .B2(data_in[0]), 
        .ZN(n9710) );
  INV_X1 U3221 ( .A(n9712), .ZN(n25705) );
  AOI22_X1 U3222 ( .A1(\mem[50][1] ), .A2(n9711), .B1(n27080), .B2(data_in[1]), 
        .ZN(n9712) );
  INV_X1 U3223 ( .A(n9713), .ZN(n25704) );
  AOI22_X1 U3224 ( .A1(\mem[50][2] ), .A2(n9711), .B1(n27080), .B2(data_in[2]), 
        .ZN(n9713) );
  INV_X1 U3225 ( .A(n9714), .ZN(n25703) );
  AOI22_X1 U3226 ( .A1(\mem[50][3] ), .A2(n9711), .B1(n27080), .B2(data_in[3]), 
        .ZN(n9714) );
  INV_X1 U3227 ( .A(n9715), .ZN(n25702) );
  AOI22_X1 U3228 ( .A1(\mem[50][4] ), .A2(n9711), .B1(n27080), .B2(data_in[4]), 
        .ZN(n9715) );
  INV_X1 U3229 ( .A(n9716), .ZN(n25701) );
  AOI22_X1 U3230 ( .A1(\mem[50][5] ), .A2(n9711), .B1(n27080), .B2(data_in[5]), 
        .ZN(n9716) );
  INV_X1 U3231 ( .A(n9717), .ZN(n25700) );
  AOI22_X1 U3232 ( .A1(\mem[50][6] ), .A2(n9711), .B1(n27080), .B2(data_in[6]), 
        .ZN(n9717) );
  INV_X1 U3233 ( .A(n9718), .ZN(n25699) );
  AOI22_X1 U3234 ( .A1(\mem[50][7] ), .A2(n9711), .B1(n27080), .B2(data_in[7]), 
        .ZN(n9718) );
  INV_X1 U3235 ( .A(n9719), .ZN(n25698) );
  AOI22_X1 U3236 ( .A1(\mem[51][0] ), .A2(n9720), .B1(n27079), .B2(data_in[0]), 
        .ZN(n9719) );
  INV_X1 U3237 ( .A(n9721), .ZN(n25697) );
  AOI22_X1 U3238 ( .A1(\mem[51][1] ), .A2(n9720), .B1(n27079), .B2(data_in[1]), 
        .ZN(n9721) );
  INV_X1 U3239 ( .A(n9722), .ZN(n25696) );
  AOI22_X1 U3240 ( .A1(\mem[51][2] ), .A2(n9720), .B1(n27079), .B2(data_in[2]), 
        .ZN(n9722) );
  INV_X1 U3241 ( .A(n9723), .ZN(n25695) );
  AOI22_X1 U3242 ( .A1(\mem[51][3] ), .A2(n9720), .B1(n27079), .B2(data_in[3]), 
        .ZN(n9723) );
  INV_X1 U3243 ( .A(n9724), .ZN(n25694) );
  AOI22_X1 U3244 ( .A1(\mem[51][4] ), .A2(n9720), .B1(n27079), .B2(data_in[4]), 
        .ZN(n9724) );
  INV_X1 U3245 ( .A(n9725), .ZN(n25693) );
  AOI22_X1 U3246 ( .A1(\mem[51][5] ), .A2(n9720), .B1(n27079), .B2(data_in[5]), 
        .ZN(n9725) );
  INV_X1 U3247 ( .A(n9726), .ZN(n25692) );
  AOI22_X1 U3248 ( .A1(\mem[51][6] ), .A2(n9720), .B1(n27079), .B2(data_in[6]), 
        .ZN(n9726) );
  INV_X1 U3249 ( .A(n9727), .ZN(n25691) );
  AOI22_X1 U3250 ( .A1(\mem[51][7] ), .A2(n9720), .B1(n27079), .B2(data_in[7]), 
        .ZN(n9727) );
  INV_X1 U3251 ( .A(n9728), .ZN(n25690) );
  AOI22_X1 U3252 ( .A1(\mem[52][0] ), .A2(n9729), .B1(n27078), .B2(data_in[0]), 
        .ZN(n9728) );
  INV_X1 U3253 ( .A(n9730), .ZN(n25689) );
  AOI22_X1 U3254 ( .A1(\mem[52][1] ), .A2(n9729), .B1(n27078), .B2(data_in[1]), 
        .ZN(n9730) );
  INV_X1 U3255 ( .A(n9731), .ZN(n25688) );
  AOI22_X1 U3256 ( .A1(\mem[52][2] ), .A2(n9729), .B1(n27078), .B2(data_in[2]), 
        .ZN(n9731) );
  INV_X1 U3257 ( .A(n9732), .ZN(n25687) );
  AOI22_X1 U3258 ( .A1(\mem[52][3] ), .A2(n9729), .B1(n27078), .B2(data_in[3]), 
        .ZN(n9732) );
  INV_X1 U3259 ( .A(n9733), .ZN(n25686) );
  AOI22_X1 U3260 ( .A1(\mem[52][4] ), .A2(n9729), .B1(n27078), .B2(data_in[4]), 
        .ZN(n9733) );
  INV_X1 U3261 ( .A(n9734), .ZN(n25685) );
  AOI22_X1 U3262 ( .A1(\mem[52][5] ), .A2(n9729), .B1(n27078), .B2(data_in[5]), 
        .ZN(n9734) );
  INV_X1 U3263 ( .A(n9735), .ZN(n25684) );
  AOI22_X1 U3264 ( .A1(\mem[52][6] ), .A2(n9729), .B1(n27078), .B2(data_in[6]), 
        .ZN(n9735) );
  INV_X1 U3265 ( .A(n9736), .ZN(n25683) );
  AOI22_X1 U3266 ( .A1(\mem[52][7] ), .A2(n9729), .B1(n27078), .B2(data_in[7]), 
        .ZN(n9736) );
  INV_X1 U3267 ( .A(n9737), .ZN(n25682) );
  AOI22_X1 U3268 ( .A1(\mem[53][0] ), .A2(n9738), .B1(n27077), .B2(data_in[0]), 
        .ZN(n9737) );
  INV_X1 U3269 ( .A(n9739), .ZN(n25681) );
  AOI22_X1 U3270 ( .A1(\mem[53][1] ), .A2(n9738), .B1(n27077), .B2(data_in[1]), 
        .ZN(n9739) );
  INV_X1 U3271 ( .A(n9740), .ZN(n25680) );
  AOI22_X1 U3272 ( .A1(\mem[53][2] ), .A2(n9738), .B1(n27077), .B2(data_in[2]), 
        .ZN(n9740) );
  INV_X1 U3273 ( .A(n9741), .ZN(n25679) );
  AOI22_X1 U3274 ( .A1(\mem[53][3] ), .A2(n9738), .B1(n27077), .B2(data_in[3]), 
        .ZN(n9741) );
  INV_X1 U3275 ( .A(n9742), .ZN(n25678) );
  AOI22_X1 U3276 ( .A1(\mem[53][4] ), .A2(n9738), .B1(n27077), .B2(data_in[4]), 
        .ZN(n9742) );
  INV_X1 U3277 ( .A(n9743), .ZN(n25677) );
  AOI22_X1 U3278 ( .A1(\mem[53][5] ), .A2(n9738), .B1(n27077), .B2(data_in[5]), 
        .ZN(n9743) );
  INV_X1 U3279 ( .A(n9744), .ZN(n25676) );
  AOI22_X1 U3280 ( .A1(\mem[53][6] ), .A2(n9738), .B1(n27077), .B2(data_in[6]), 
        .ZN(n9744) );
  INV_X1 U3281 ( .A(n9745), .ZN(n25675) );
  AOI22_X1 U3282 ( .A1(\mem[53][7] ), .A2(n9738), .B1(n27077), .B2(data_in[7]), 
        .ZN(n9745) );
  INV_X1 U3283 ( .A(n9746), .ZN(n25674) );
  AOI22_X1 U3284 ( .A1(\mem[54][0] ), .A2(n9747), .B1(n27076), .B2(data_in[0]), 
        .ZN(n9746) );
  INV_X1 U3285 ( .A(n9748), .ZN(n25673) );
  AOI22_X1 U3286 ( .A1(\mem[54][1] ), .A2(n9747), .B1(n27076), .B2(data_in[1]), 
        .ZN(n9748) );
  INV_X1 U3287 ( .A(n9749), .ZN(n25672) );
  AOI22_X1 U3288 ( .A1(\mem[54][2] ), .A2(n9747), .B1(n27076), .B2(data_in[2]), 
        .ZN(n9749) );
  INV_X1 U3289 ( .A(n9750), .ZN(n25671) );
  AOI22_X1 U3290 ( .A1(\mem[54][3] ), .A2(n9747), .B1(n27076), .B2(data_in[3]), 
        .ZN(n9750) );
  INV_X1 U3291 ( .A(n9751), .ZN(n25670) );
  AOI22_X1 U3292 ( .A1(\mem[54][4] ), .A2(n9747), .B1(n27076), .B2(data_in[4]), 
        .ZN(n9751) );
  INV_X1 U3293 ( .A(n9752), .ZN(n25669) );
  AOI22_X1 U3294 ( .A1(\mem[54][5] ), .A2(n9747), .B1(n27076), .B2(data_in[5]), 
        .ZN(n9752) );
  INV_X1 U3295 ( .A(n9753), .ZN(n25668) );
  AOI22_X1 U3296 ( .A1(\mem[54][6] ), .A2(n9747), .B1(n27076), .B2(data_in[6]), 
        .ZN(n9753) );
  INV_X1 U3297 ( .A(n9754), .ZN(n25667) );
  AOI22_X1 U3298 ( .A1(\mem[54][7] ), .A2(n9747), .B1(n27076), .B2(data_in[7]), 
        .ZN(n9754) );
  INV_X1 U3299 ( .A(n9755), .ZN(n25666) );
  AOI22_X1 U3300 ( .A1(\mem[55][0] ), .A2(n9756), .B1(n27075), .B2(data_in[0]), 
        .ZN(n9755) );
  INV_X1 U3301 ( .A(n9757), .ZN(n25665) );
  AOI22_X1 U3302 ( .A1(\mem[55][1] ), .A2(n9756), .B1(n27075), .B2(data_in[1]), 
        .ZN(n9757) );
  INV_X1 U3303 ( .A(n9758), .ZN(n25664) );
  AOI22_X1 U3304 ( .A1(\mem[55][2] ), .A2(n9756), .B1(n27075), .B2(data_in[2]), 
        .ZN(n9758) );
  INV_X1 U3305 ( .A(n9759), .ZN(n25663) );
  AOI22_X1 U3306 ( .A1(\mem[55][3] ), .A2(n9756), .B1(n27075), .B2(data_in[3]), 
        .ZN(n9759) );
  INV_X1 U3307 ( .A(n9760), .ZN(n25662) );
  AOI22_X1 U3308 ( .A1(\mem[55][4] ), .A2(n9756), .B1(n27075), .B2(data_in[4]), 
        .ZN(n9760) );
  INV_X1 U3309 ( .A(n9761), .ZN(n25661) );
  AOI22_X1 U3310 ( .A1(\mem[55][5] ), .A2(n9756), .B1(n27075), .B2(data_in[5]), 
        .ZN(n9761) );
  INV_X1 U3311 ( .A(n9762), .ZN(n25660) );
  AOI22_X1 U3312 ( .A1(\mem[55][6] ), .A2(n9756), .B1(n27075), .B2(data_in[6]), 
        .ZN(n9762) );
  INV_X1 U3313 ( .A(n9763), .ZN(n25659) );
  AOI22_X1 U3314 ( .A1(\mem[55][7] ), .A2(n9756), .B1(n27075), .B2(data_in[7]), 
        .ZN(n9763) );
  INV_X1 U3315 ( .A(n9764), .ZN(n25658) );
  AOI22_X1 U3316 ( .A1(\mem[56][0] ), .A2(n9765), .B1(n27074), .B2(data_in[0]), 
        .ZN(n9764) );
  INV_X1 U3317 ( .A(n9766), .ZN(n25657) );
  AOI22_X1 U3318 ( .A1(\mem[56][1] ), .A2(n9765), .B1(n27074), .B2(data_in[1]), 
        .ZN(n9766) );
  INV_X1 U3319 ( .A(n9767), .ZN(n25656) );
  AOI22_X1 U3320 ( .A1(\mem[56][2] ), .A2(n9765), .B1(n27074), .B2(data_in[2]), 
        .ZN(n9767) );
  INV_X1 U3321 ( .A(n9768), .ZN(n25655) );
  AOI22_X1 U3322 ( .A1(\mem[56][3] ), .A2(n9765), .B1(n27074), .B2(data_in[3]), 
        .ZN(n9768) );
  INV_X1 U3323 ( .A(n9769), .ZN(n25654) );
  AOI22_X1 U3324 ( .A1(\mem[56][4] ), .A2(n9765), .B1(n27074), .B2(data_in[4]), 
        .ZN(n9769) );
  INV_X1 U3325 ( .A(n9770), .ZN(n25653) );
  AOI22_X1 U3326 ( .A1(\mem[56][5] ), .A2(n9765), .B1(n27074), .B2(data_in[5]), 
        .ZN(n9770) );
  INV_X1 U3327 ( .A(n9771), .ZN(n25652) );
  AOI22_X1 U3328 ( .A1(\mem[56][6] ), .A2(n9765), .B1(n27074), .B2(data_in[6]), 
        .ZN(n9771) );
  INV_X1 U3329 ( .A(n9772), .ZN(n25651) );
  AOI22_X1 U3330 ( .A1(\mem[56][7] ), .A2(n9765), .B1(n27074), .B2(data_in[7]), 
        .ZN(n9772) );
  INV_X1 U3331 ( .A(n9773), .ZN(n25650) );
  AOI22_X1 U3332 ( .A1(\mem[57][0] ), .A2(n9774), .B1(n27073), .B2(data_in[0]), 
        .ZN(n9773) );
  INV_X1 U3333 ( .A(n9775), .ZN(n25649) );
  AOI22_X1 U3334 ( .A1(\mem[57][1] ), .A2(n9774), .B1(n27073), .B2(data_in[1]), 
        .ZN(n9775) );
  INV_X1 U3335 ( .A(n9776), .ZN(n25648) );
  AOI22_X1 U3336 ( .A1(\mem[57][2] ), .A2(n9774), .B1(n27073), .B2(data_in[2]), 
        .ZN(n9776) );
  INV_X1 U3337 ( .A(n9777), .ZN(n25647) );
  AOI22_X1 U3338 ( .A1(\mem[57][3] ), .A2(n9774), .B1(n27073), .B2(data_in[3]), 
        .ZN(n9777) );
  INV_X1 U3339 ( .A(n9778), .ZN(n25646) );
  AOI22_X1 U3340 ( .A1(\mem[57][4] ), .A2(n9774), .B1(n27073), .B2(data_in[4]), 
        .ZN(n9778) );
  INV_X1 U3341 ( .A(n9779), .ZN(n25645) );
  AOI22_X1 U3342 ( .A1(\mem[57][5] ), .A2(n9774), .B1(n27073), .B2(data_in[5]), 
        .ZN(n9779) );
  INV_X1 U3343 ( .A(n9780), .ZN(n25644) );
  AOI22_X1 U3344 ( .A1(\mem[57][6] ), .A2(n9774), .B1(n27073), .B2(data_in[6]), 
        .ZN(n9780) );
  INV_X1 U3345 ( .A(n9781), .ZN(n25643) );
  AOI22_X1 U3346 ( .A1(\mem[57][7] ), .A2(n9774), .B1(n27073), .B2(data_in[7]), 
        .ZN(n9781) );
  INV_X1 U3347 ( .A(n9782), .ZN(n25642) );
  AOI22_X1 U3348 ( .A1(\mem[58][0] ), .A2(n9783), .B1(n27072), .B2(data_in[0]), 
        .ZN(n9782) );
  INV_X1 U3349 ( .A(n9784), .ZN(n25641) );
  AOI22_X1 U3350 ( .A1(\mem[58][1] ), .A2(n9783), .B1(n27072), .B2(data_in[1]), 
        .ZN(n9784) );
  INV_X1 U3351 ( .A(n9785), .ZN(n25640) );
  AOI22_X1 U3352 ( .A1(\mem[58][2] ), .A2(n9783), .B1(n27072), .B2(data_in[2]), 
        .ZN(n9785) );
  INV_X1 U3353 ( .A(n9786), .ZN(n25639) );
  AOI22_X1 U3354 ( .A1(\mem[58][3] ), .A2(n9783), .B1(n27072), .B2(data_in[3]), 
        .ZN(n9786) );
  INV_X1 U3355 ( .A(n9787), .ZN(n25638) );
  AOI22_X1 U3356 ( .A1(\mem[58][4] ), .A2(n9783), .B1(n27072), .B2(data_in[4]), 
        .ZN(n9787) );
  INV_X1 U3357 ( .A(n9788), .ZN(n25637) );
  AOI22_X1 U3358 ( .A1(\mem[58][5] ), .A2(n9783), .B1(n27072), .B2(data_in[5]), 
        .ZN(n9788) );
  INV_X1 U3359 ( .A(n9789), .ZN(n25636) );
  AOI22_X1 U3360 ( .A1(\mem[58][6] ), .A2(n9783), .B1(n27072), .B2(data_in[6]), 
        .ZN(n9789) );
  INV_X1 U3361 ( .A(n9790), .ZN(n25635) );
  AOI22_X1 U3362 ( .A1(\mem[58][7] ), .A2(n9783), .B1(n27072), .B2(data_in[7]), 
        .ZN(n9790) );
  INV_X1 U3363 ( .A(n9791), .ZN(n25634) );
  AOI22_X1 U3364 ( .A1(\mem[59][0] ), .A2(n9792), .B1(n27071), .B2(data_in[0]), 
        .ZN(n9791) );
  INV_X1 U3365 ( .A(n9793), .ZN(n25633) );
  AOI22_X1 U3366 ( .A1(\mem[59][1] ), .A2(n9792), .B1(n27071), .B2(data_in[1]), 
        .ZN(n9793) );
  INV_X1 U3367 ( .A(n9794), .ZN(n25632) );
  AOI22_X1 U3368 ( .A1(\mem[59][2] ), .A2(n9792), .B1(n27071), .B2(data_in[2]), 
        .ZN(n9794) );
  INV_X1 U3369 ( .A(n9795), .ZN(n25631) );
  AOI22_X1 U3370 ( .A1(\mem[59][3] ), .A2(n9792), .B1(n27071), .B2(data_in[3]), 
        .ZN(n9795) );
  INV_X1 U3371 ( .A(n9796), .ZN(n25630) );
  AOI22_X1 U3372 ( .A1(\mem[59][4] ), .A2(n9792), .B1(n27071), .B2(data_in[4]), 
        .ZN(n9796) );
  INV_X1 U3373 ( .A(n9797), .ZN(n25629) );
  AOI22_X1 U3374 ( .A1(\mem[59][5] ), .A2(n9792), .B1(n27071), .B2(data_in[5]), 
        .ZN(n9797) );
  INV_X1 U3375 ( .A(n9798), .ZN(n25628) );
  AOI22_X1 U3376 ( .A1(\mem[59][6] ), .A2(n9792), .B1(n27071), .B2(data_in[6]), 
        .ZN(n9798) );
  INV_X1 U3377 ( .A(n9799), .ZN(n25627) );
  AOI22_X1 U3378 ( .A1(\mem[59][7] ), .A2(n9792), .B1(n27071), .B2(data_in[7]), 
        .ZN(n9799) );
  INV_X1 U3379 ( .A(n9800), .ZN(n25626) );
  AOI22_X1 U3380 ( .A1(\mem[60][0] ), .A2(n9801), .B1(n27070), .B2(data_in[0]), 
        .ZN(n9800) );
  INV_X1 U3381 ( .A(n9802), .ZN(n25625) );
  AOI22_X1 U3382 ( .A1(\mem[60][1] ), .A2(n9801), .B1(n27070), .B2(data_in[1]), 
        .ZN(n9802) );
  INV_X1 U3383 ( .A(n9803), .ZN(n25624) );
  AOI22_X1 U3384 ( .A1(\mem[60][2] ), .A2(n9801), .B1(n27070), .B2(data_in[2]), 
        .ZN(n9803) );
  INV_X1 U3385 ( .A(n9804), .ZN(n25623) );
  AOI22_X1 U3386 ( .A1(\mem[60][3] ), .A2(n9801), .B1(n27070), .B2(data_in[3]), 
        .ZN(n9804) );
  INV_X1 U3387 ( .A(n9805), .ZN(n25622) );
  AOI22_X1 U3388 ( .A1(\mem[60][4] ), .A2(n9801), .B1(n27070), .B2(data_in[4]), 
        .ZN(n9805) );
  INV_X1 U3389 ( .A(n9806), .ZN(n25621) );
  AOI22_X1 U3390 ( .A1(\mem[60][5] ), .A2(n9801), .B1(n27070), .B2(data_in[5]), 
        .ZN(n9806) );
  INV_X1 U3391 ( .A(n9807), .ZN(n25620) );
  AOI22_X1 U3392 ( .A1(\mem[60][6] ), .A2(n9801), .B1(n27070), .B2(data_in[6]), 
        .ZN(n9807) );
  INV_X1 U3393 ( .A(n9808), .ZN(n25619) );
  AOI22_X1 U3394 ( .A1(\mem[60][7] ), .A2(n9801), .B1(n27070), .B2(data_in[7]), 
        .ZN(n9808) );
  INV_X1 U3395 ( .A(n9809), .ZN(n25618) );
  AOI22_X1 U3396 ( .A1(\mem[61][0] ), .A2(n9810), .B1(n27069), .B2(data_in[0]), 
        .ZN(n9809) );
  INV_X1 U3397 ( .A(n9811), .ZN(n25617) );
  AOI22_X1 U3398 ( .A1(\mem[61][1] ), .A2(n9810), .B1(n27069), .B2(data_in[1]), 
        .ZN(n9811) );
  INV_X1 U3399 ( .A(n9812), .ZN(n25616) );
  AOI22_X1 U3400 ( .A1(\mem[61][2] ), .A2(n9810), .B1(n27069), .B2(data_in[2]), 
        .ZN(n9812) );
  INV_X1 U3401 ( .A(n9813), .ZN(n25615) );
  AOI22_X1 U3402 ( .A1(\mem[61][3] ), .A2(n9810), .B1(n27069), .B2(data_in[3]), 
        .ZN(n9813) );
  INV_X1 U3403 ( .A(n9814), .ZN(n25614) );
  AOI22_X1 U3404 ( .A1(\mem[61][4] ), .A2(n9810), .B1(n27069), .B2(data_in[4]), 
        .ZN(n9814) );
  INV_X1 U3405 ( .A(n9815), .ZN(n25613) );
  AOI22_X1 U3406 ( .A1(\mem[61][5] ), .A2(n9810), .B1(n27069), .B2(data_in[5]), 
        .ZN(n9815) );
  INV_X1 U3407 ( .A(n9816), .ZN(n25612) );
  AOI22_X1 U3408 ( .A1(\mem[61][6] ), .A2(n9810), .B1(n27069), .B2(data_in[6]), 
        .ZN(n9816) );
  INV_X1 U3409 ( .A(n9817), .ZN(n25611) );
  AOI22_X1 U3410 ( .A1(\mem[61][7] ), .A2(n9810), .B1(n27069), .B2(data_in[7]), 
        .ZN(n9817) );
  INV_X1 U3411 ( .A(n9818), .ZN(n25610) );
  AOI22_X1 U3412 ( .A1(\mem[62][0] ), .A2(n9819), .B1(n27068), .B2(data_in[0]), 
        .ZN(n9818) );
  INV_X1 U3413 ( .A(n9820), .ZN(n25609) );
  AOI22_X1 U3414 ( .A1(\mem[62][1] ), .A2(n9819), .B1(n27068), .B2(data_in[1]), 
        .ZN(n9820) );
  INV_X1 U3415 ( .A(n9821), .ZN(n25608) );
  AOI22_X1 U3416 ( .A1(\mem[62][2] ), .A2(n9819), .B1(n27068), .B2(data_in[2]), 
        .ZN(n9821) );
  INV_X1 U3417 ( .A(n9822), .ZN(n25607) );
  AOI22_X1 U3418 ( .A1(\mem[62][3] ), .A2(n9819), .B1(n27068), .B2(data_in[3]), 
        .ZN(n9822) );
  INV_X1 U3419 ( .A(n9823), .ZN(n25606) );
  AOI22_X1 U3420 ( .A1(\mem[62][4] ), .A2(n9819), .B1(n27068), .B2(data_in[4]), 
        .ZN(n9823) );
  INV_X1 U3421 ( .A(n9824), .ZN(n25605) );
  AOI22_X1 U3422 ( .A1(\mem[62][5] ), .A2(n9819), .B1(n27068), .B2(data_in[5]), 
        .ZN(n9824) );
  INV_X1 U3423 ( .A(n9825), .ZN(n25604) );
  AOI22_X1 U3424 ( .A1(\mem[62][6] ), .A2(n9819), .B1(n27068), .B2(data_in[6]), 
        .ZN(n9825) );
  INV_X1 U3425 ( .A(n9826), .ZN(n25603) );
  AOI22_X1 U3426 ( .A1(\mem[62][7] ), .A2(n9819), .B1(n27068), .B2(data_in[7]), 
        .ZN(n9826) );
  INV_X1 U3427 ( .A(n9827), .ZN(n25602) );
  AOI22_X1 U3428 ( .A1(\mem[63][0] ), .A2(n9828), .B1(n27067), .B2(data_in[0]), 
        .ZN(n9827) );
  INV_X1 U3429 ( .A(n9829), .ZN(n25601) );
  AOI22_X1 U3430 ( .A1(\mem[63][1] ), .A2(n9828), .B1(n27067), .B2(data_in[1]), 
        .ZN(n9829) );
  INV_X1 U3431 ( .A(n9830), .ZN(n25600) );
  AOI22_X1 U3432 ( .A1(\mem[63][2] ), .A2(n9828), .B1(n27067), .B2(data_in[2]), 
        .ZN(n9830) );
  INV_X1 U3433 ( .A(n9831), .ZN(n25599) );
  AOI22_X1 U3434 ( .A1(\mem[63][3] ), .A2(n9828), .B1(n27067), .B2(data_in[3]), 
        .ZN(n9831) );
  INV_X1 U3435 ( .A(n9832), .ZN(n25598) );
  AOI22_X1 U3436 ( .A1(\mem[63][4] ), .A2(n9828), .B1(n27067), .B2(data_in[4]), 
        .ZN(n9832) );
  INV_X1 U3437 ( .A(n9833), .ZN(n25597) );
  AOI22_X1 U3438 ( .A1(\mem[63][5] ), .A2(n9828), .B1(n27067), .B2(data_in[5]), 
        .ZN(n9833) );
  INV_X1 U3439 ( .A(n9834), .ZN(n25596) );
  AOI22_X1 U3440 ( .A1(\mem[63][6] ), .A2(n9828), .B1(n27067), .B2(data_in[6]), 
        .ZN(n9834) );
  INV_X1 U3441 ( .A(n9835), .ZN(n25595) );
  AOI22_X1 U3442 ( .A1(\mem[63][7] ), .A2(n9828), .B1(n27067), .B2(data_in[7]), 
        .ZN(n9835) );
  INV_X1 U3443 ( .A(n9910), .ZN(n25530) );
  AOI22_X1 U3444 ( .A1(\mem[72][0] ), .A2(n9911), .B1(n27058), .B2(data_in[0]), 
        .ZN(n9910) );
  INV_X1 U3445 ( .A(n9912), .ZN(n25529) );
  AOI22_X1 U3446 ( .A1(\mem[72][1] ), .A2(n9911), .B1(n27058), .B2(data_in[1]), 
        .ZN(n9912) );
  INV_X1 U3447 ( .A(n9913), .ZN(n25528) );
  AOI22_X1 U3448 ( .A1(\mem[72][2] ), .A2(n9911), .B1(n27058), .B2(data_in[2]), 
        .ZN(n9913) );
  INV_X1 U3449 ( .A(n9914), .ZN(n25527) );
  AOI22_X1 U3450 ( .A1(\mem[72][3] ), .A2(n9911), .B1(n27058), .B2(data_in[3]), 
        .ZN(n9914) );
  INV_X1 U3451 ( .A(n9915), .ZN(n25526) );
  AOI22_X1 U3452 ( .A1(\mem[72][4] ), .A2(n9911), .B1(n27058), .B2(data_in[4]), 
        .ZN(n9915) );
  INV_X1 U3453 ( .A(n9916), .ZN(n25525) );
  AOI22_X1 U3454 ( .A1(\mem[72][5] ), .A2(n9911), .B1(n27058), .B2(data_in[5]), 
        .ZN(n9916) );
  INV_X1 U3455 ( .A(n9917), .ZN(n25524) );
  AOI22_X1 U3456 ( .A1(\mem[72][6] ), .A2(n9911), .B1(n27058), .B2(data_in[6]), 
        .ZN(n9917) );
  INV_X1 U3457 ( .A(n9918), .ZN(n25523) );
  AOI22_X1 U3458 ( .A1(\mem[72][7] ), .A2(n9911), .B1(n27058), .B2(data_in[7]), 
        .ZN(n9918) );
  INV_X1 U3459 ( .A(n9919), .ZN(n25522) );
  AOI22_X1 U3460 ( .A1(\mem[73][0] ), .A2(n9920), .B1(n27057), .B2(data_in[0]), 
        .ZN(n9919) );
  INV_X1 U3461 ( .A(n9921), .ZN(n25521) );
  AOI22_X1 U3462 ( .A1(\mem[73][1] ), .A2(n9920), .B1(n27057), .B2(data_in[1]), 
        .ZN(n9921) );
  INV_X1 U3463 ( .A(n9922), .ZN(n25520) );
  AOI22_X1 U3464 ( .A1(\mem[73][2] ), .A2(n9920), .B1(n27057), .B2(data_in[2]), 
        .ZN(n9922) );
  INV_X1 U3465 ( .A(n9923), .ZN(n25519) );
  AOI22_X1 U3466 ( .A1(\mem[73][3] ), .A2(n9920), .B1(n27057), .B2(data_in[3]), 
        .ZN(n9923) );
  INV_X1 U3467 ( .A(n9924), .ZN(n25518) );
  AOI22_X1 U3468 ( .A1(\mem[73][4] ), .A2(n9920), .B1(n27057), .B2(data_in[4]), 
        .ZN(n9924) );
  INV_X1 U3469 ( .A(n9925), .ZN(n25517) );
  AOI22_X1 U3470 ( .A1(\mem[73][5] ), .A2(n9920), .B1(n27057), .B2(data_in[5]), 
        .ZN(n9925) );
  INV_X1 U3471 ( .A(n9926), .ZN(n25516) );
  AOI22_X1 U3472 ( .A1(\mem[73][6] ), .A2(n9920), .B1(n27057), .B2(data_in[6]), 
        .ZN(n9926) );
  INV_X1 U3473 ( .A(n9927), .ZN(n25515) );
  AOI22_X1 U3474 ( .A1(\mem[73][7] ), .A2(n9920), .B1(n27057), .B2(data_in[7]), 
        .ZN(n9927) );
  INV_X1 U3475 ( .A(n9928), .ZN(n25514) );
  AOI22_X1 U3476 ( .A1(\mem[74][0] ), .A2(n9929), .B1(n27056), .B2(data_in[0]), 
        .ZN(n9928) );
  INV_X1 U3477 ( .A(n9930), .ZN(n25513) );
  AOI22_X1 U3478 ( .A1(\mem[74][1] ), .A2(n9929), .B1(n27056), .B2(data_in[1]), 
        .ZN(n9930) );
  INV_X1 U3479 ( .A(n9931), .ZN(n25512) );
  AOI22_X1 U3480 ( .A1(\mem[74][2] ), .A2(n9929), .B1(n27056), .B2(data_in[2]), 
        .ZN(n9931) );
  INV_X1 U3481 ( .A(n9932), .ZN(n25511) );
  AOI22_X1 U3482 ( .A1(\mem[74][3] ), .A2(n9929), .B1(n27056), .B2(data_in[3]), 
        .ZN(n9932) );
  INV_X1 U3483 ( .A(n9933), .ZN(n25510) );
  AOI22_X1 U3484 ( .A1(\mem[74][4] ), .A2(n9929), .B1(n27056), .B2(data_in[4]), 
        .ZN(n9933) );
  INV_X1 U3485 ( .A(n9934), .ZN(n25509) );
  AOI22_X1 U3486 ( .A1(\mem[74][5] ), .A2(n9929), .B1(n27056), .B2(data_in[5]), 
        .ZN(n9934) );
  INV_X1 U3487 ( .A(n9935), .ZN(n25508) );
  AOI22_X1 U3488 ( .A1(\mem[74][6] ), .A2(n9929), .B1(n27056), .B2(data_in[6]), 
        .ZN(n9935) );
  INV_X1 U3489 ( .A(n9936), .ZN(n25507) );
  AOI22_X1 U3490 ( .A1(\mem[74][7] ), .A2(n9929), .B1(n27056), .B2(data_in[7]), 
        .ZN(n9936) );
  INV_X1 U3491 ( .A(n9937), .ZN(n25506) );
  AOI22_X1 U3492 ( .A1(\mem[75][0] ), .A2(n9938), .B1(n27055), .B2(data_in[0]), 
        .ZN(n9937) );
  INV_X1 U3493 ( .A(n9939), .ZN(n25505) );
  AOI22_X1 U3494 ( .A1(\mem[75][1] ), .A2(n9938), .B1(n27055), .B2(data_in[1]), 
        .ZN(n9939) );
  INV_X1 U3495 ( .A(n9940), .ZN(n25504) );
  AOI22_X1 U3496 ( .A1(\mem[75][2] ), .A2(n9938), .B1(n27055), .B2(data_in[2]), 
        .ZN(n9940) );
  INV_X1 U3497 ( .A(n9941), .ZN(n25503) );
  AOI22_X1 U3498 ( .A1(\mem[75][3] ), .A2(n9938), .B1(n27055), .B2(data_in[3]), 
        .ZN(n9941) );
  INV_X1 U3499 ( .A(n9942), .ZN(n25502) );
  AOI22_X1 U3500 ( .A1(\mem[75][4] ), .A2(n9938), .B1(n27055), .B2(data_in[4]), 
        .ZN(n9942) );
  INV_X1 U3501 ( .A(n9943), .ZN(n25501) );
  AOI22_X1 U3502 ( .A1(\mem[75][5] ), .A2(n9938), .B1(n27055), .B2(data_in[5]), 
        .ZN(n9943) );
  INV_X1 U3503 ( .A(n9944), .ZN(n25500) );
  AOI22_X1 U3504 ( .A1(\mem[75][6] ), .A2(n9938), .B1(n27055), .B2(data_in[6]), 
        .ZN(n9944) );
  INV_X1 U3505 ( .A(n9945), .ZN(n25499) );
  AOI22_X1 U3506 ( .A1(\mem[75][7] ), .A2(n9938), .B1(n27055), .B2(data_in[7]), 
        .ZN(n9945) );
  INV_X1 U3507 ( .A(n9946), .ZN(n25498) );
  AOI22_X1 U3508 ( .A1(\mem[76][0] ), .A2(n9947), .B1(n27054), .B2(data_in[0]), 
        .ZN(n9946) );
  INV_X1 U3509 ( .A(n9948), .ZN(n25497) );
  AOI22_X1 U3510 ( .A1(\mem[76][1] ), .A2(n9947), .B1(n27054), .B2(data_in[1]), 
        .ZN(n9948) );
  INV_X1 U3511 ( .A(n9949), .ZN(n25496) );
  AOI22_X1 U3512 ( .A1(\mem[76][2] ), .A2(n9947), .B1(n27054), .B2(data_in[2]), 
        .ZN(n9949) );
  INV_X1 U3513 ( .A(n9950), .ZN(n25495) );
  AOI22_X1 U3514 ( .A1(\mem[76][3] ), .A2(n9947), .B1(n27054), .B2(data_in[3]), 
        .ZN(n9950) );
  INV_X1 U3515 ( .A(n9951), .ZN(n25494) );
  AOI22_X1 U3516 ( .A1(\mem[76][4] ), .A2(n9947), .B1(n27054), .B2(data_in[4]), 
        .ZN(n9951) );
  INV_X1 U3517 ( .A(n9952), .ZN(n25493) );
  AOI22_X1 U3518 ( .A1(\mem[76][5] ), .A2(n9947), .B1(n27054), .B2(data_in[5]), 
        .ZN(n9952) );
  INV_X1 U3519 ( .A(n9953), .ZN(n25492) );
  AOI22_X1 U3520 ( .A1(\mem[76][6] ), .A2(n9947), .B1(n27054), .B2(data_in[6]), 
        .ZN(n9953) );
  INV_X1 U3521 ( .A(n9954), .ZN(n25491) );
  AOI22_X1 U3522 ( .A1(\mem[76][7] ), .A2(n9947), .B1(n27054), .B2(data_in[7]), 
        .ZN(n9954) );
  INV_X1 U3523 ( .A(n9955), .ZN(n25490) );
  AOI22_X1 U3524 ( .A1(\mem[77][0] ), .A2(n9956), .B1(n27053), .B2(data_in[0]), 
        .ZN(n9955) );
  INV_X1 U3525 ( .A(n9957), .ZN(n25489) );
  AOI22_X1 U3526 ( .A1(\mem[77][1] ), .A2(n9956), .B1(n27053), .B2(data_in[1]), 
        .ZN(n9957) );
  INV_X1 U3527 ( .A(n9958), .ZN(n25488) );
  AOI22_X1 U3528 ( .A1(\mem[77][2] ), .A2(n9956), .B1(n27053), .B2(data_in[2]), 
        .ZN(n9958) );
  INV_X1 U3529 ( .A(n9959), .ZN(n25487) );
  AOI22_X1 U3530 ( .A1(\mem[77][3] ), .A2(n9956), .B1(n27053), .B2(data_in[3]), 
        .ZN(n9959) );
  INV_X1 U3531 ( .A(n9960), .ZN(n25486) );
  AOI22_X1 U3532 ( .A1(\mem[77][4] ), .A2(n9956), .B1(n27053), .B2(data_in[4]), 
        .ZN(n9960) );
  INV_X1 U3533 ( .A(n9961), .ZN(n25485) );
  AOI22_X1 U3534 ( .A1(\mem[77][5] ), .A2(n9956), .B1(n27053), .B2(data_in[5]), 
        .ZN(n9961) );
  INV_X1 U3535 ( .A(n9962), .ZN(n25484) );
  AOI22_X1 U3536 ( .A1(\mem[77][6] ), .A2(n9956), .B1(n27053), .B2(data_in[6]), 
        .ZN(n9962) );
  INV_X1 U3537 ( .A(n9963), .ZN(n25483) );
  AOI22_X1 U3538 ( .A1(\mem[77][7] ), .A2(n9956), .B1(n27053), .B2(data_in[7]), 
        .ZN(n9963) );
  INV_X1 U3539 ( .A(n9964), .ZN(n25482) );
  AOI22_X1 U3540 ( .A1(\mem[78][0] ), .A2(n9965), .B1(n27052), .B2(data_in[0]), 
        .ZN(n9964) );
  INV_X1 U3541 ( .A(n9966), .ZN(n25481) );
  AOI22_X1 U3542 ( .A1(\mem[78][1] ), .A2(n9965), .B1(n27052), .B2(data_in[1]), 
        .ZN(n9966) );
  INV_X1 U3543 ( .A(n9967), .ZN(n25480) );
  AOI22_X1 U3544 ( .A1(\mem[78][2] ), .A2(n9965), .B1(n27052), .B2(data_in[2]), 
        .ZN(n9967) );
  INV_X1 U3545 ( .A(n9968), .ZN(n25479) );
  AOI22_X1 U3546 ( .A1(\mem[78][3] ), .A2(n9965), .B1(n27052), .B2(data_in[3]), 
        .ZN(n9968) );
  INV_X1 U3547 ( .A(n9969), .ZN(n25478) );
  AOI22_X1 U3548 ( .A1(\mem[78][4] ), .A2(n9965), .B1(n27052), .B2(data_in[4]), 
        .ZN(n9969) );
  INV_X1 U3549 ( .A(n9970), .ZN(n25477) );
  AOI22_X1 U3550 ( .A1(\mem[78][5] ), .A2(n9965), .B1(n27052), .B2(data_in[5]), 
        .ZN(n9970) );
  INV_X1 U3551 ( .A(n9971), .ZN(n25476) );
  AOI22_X1 U3552 ( .A1(\mem[78][6] ), .A2(n9965), .B1(n27052), .B2(data_in[6]), 
        .ZN(n9971) );
  INV_X1 U3553 ( .A(n9972), .ZN(n25475) );
  AOI22_X1 U3554 ( .A1(\mem[78][7] ), .A2(n9965), .B1(n27052), .B2(data_in[7]), 
        .ZN(n9972) );
  INV_X1 U3555 ( .A(n9973), .ZN(n25474) );
  AOI22_X1 U3556 ( .A1(\mem[79][0] ), .A2(n9974), .B1(n27051), .B2(data_in[0]), 
        .ZN(n9973) );
  INV_X1 U3557 ( .A(n9975), .ZN(n25473) );
  AOI22_X1 U3558 ( .A1(\mem[79][1] ), .A2(n9974), .B1(n27051), .B2(data_in[1]), 
        .ZN(n9975) );
  INV_X1 U3559 ( .A(n9976), .ZN(n25472) );
  AOI22_X1 U3560 ( .A1(\mem[79][2] ), .A2(n9974), .B1(n27051), .B2(data_in[2]), 
        .ZN(n9976) );
  INV_X1 U3561 ( .A(n9977), .ZN(n25471) );
  AOI22_X1 U3562 ( .A1(\mem[79][3] ), .A2(n9974), .B1(n27051), .B2(data_in[3]), 
        .ZN(n9977) );
  INV_X1 U3563 ( .A(n9978), .ZN(n25470) );
  AOI22_X1 U3564 ( .A1(\mem[79][4] ), .A2(n9974), .B1(n27051), .B2(data_in[4]), 
        .ZN(n9978) );
  INV_X1 U3565 ( .A(n9979), .ZN(n25469) );
  AOI22_X1 U3566 ( .A1(\mem[79][5] ), .A2(n9974), .B1(n27051), .B2(data_in[5]), 
        .ZN(n9979) );
  INV_X1 U3567 ( .A(n9980), .ZN(n25468) );
  AOI22_X1 U3568 ( .A1(\mem[79][6] ), .A2(n9974), .B1(n27051), .B2(data_in[6]), 
        .ZN(n9980) );
  INV_X1 U3569 ( .A(n9981), .ZN(n25467) );
  AOI22_X1 U3570 ( .A1(\mem[79][7] ), .A2(n9974), .B1(n27051), .B2(data_in[7]), 
        .ZN(n9981) );
  INV_X1 U3571 ( .A(n9982), .ZN(n25466) );
  AOI22_X1 U3572 ( .A1(\mem[80][0] ), .A2(n9983), .B1(n27050), .B2(data_in[0]), 
        .ZN(n9982) );
  INV_X1 U3573 ( .A(n9984), .ZN(n25465) );
  AOI22_X1 U3574 ( .A1(\mem[80][1] ), .A2(n9983), .B1(n27050), .B2(data_in[1]), 
        .ZN(n9984) );
  INV_X1 U3575 ( .A(n9985), .ZN(n25464) );
  AOI22_X1 U3576 ( .A1(\mem[80][2] ), .A2(n9983), .B1(n27050), .B2(data_in[2]), 
        .ZN(n9985) );
  INV_X1 U3577 ( .A(n9986), .ZN(n25463) );
  AOI22_X1 U3578 ( .A1(\mem[80][3] ), .A2(n9983), .B1(n27050), .B2(data_in[3]), 
        .ZN(n9986) );
  INV_X1 U3579 ( .A(n9987), .ZN(n25462) );
  AOI22_X1 U3580 ( .A1(\mem[80][4] ), .A2(n9983), .B1(n27050), .B2(data_in[4]), 
        .ZN(n9987) );
  INV_X1 U3581 ( .A(n9988), .ZN(n25461) );
  AOI22_X1 U3582 ( .A1(\mem[80][5] ), .A2(n9983), .B1(n27050), .B2(data_in[5]), 
        .ZN(n9988) );
  INV_X1 U3583 ( .A(n9989), .ZN(n25460) );
  AOI22_X1 U3584 ( .A1(\mem[80][6] ), .A2(n9983), .B1(n27050), .B2(data_in[6]), 
        .ZN(n9989) );
  INV_X1 U3585 ( .A(n9990), .ZN(n25459) );
  AOI22_X1 U3586 ( .A1(\mem[80][7] ), .A2(n9983), .B1(n27050), .B2(data_in[7]), 
        .ZN(n9990) );
  INV_X1 U3587 ( .A(n9991), .ZN(n25458) );
  AOI22_X1 U3588 ( .A1(\mem[81][0] ), .A2(n9992), .B1(n27049), .B2(data_in[0]), 
        .ZN(n9991) );
  INV_X1 U3589 ( .A(n9993), .ZN(n25457) );
  AOI22_X1 U3590 ( .A1(\mem[81][1] ), .A2(n9992), .B1(n27049), .B2(data_in[1]), 
        .ZN(n9993) );
  INV_X1 U3591 ( .A(n9994), .ZN(n25456) );
  AOI22_X1 U3592 ( .A1(\mem[81][2] ), .A2(n9992), .B1(n27049), .B2(data_in[2]), 
        .ZN(n9994) );
  INV_X1 U3593 ( .A(n9995), .ZN(n25455) );
  AOI22_X1 U3594 ( .A1(\mem[81][3] ), .A2(n9992), .B1(n27049), .B2(data_in[3]), 
        .ZN(n9995) );
  INV_X1 U3595 ( .A(n9996), .ZN(n25454) );
  AOI22_X1 U3596 ( .A1(\mem[81][4] ), .A2(n9992), .B1(n27049), .B2(data_in[4]), 
        .ZN(n9996) );
  INV_X1 U3597 ( .A(n9997), .ZN(n25453) );
  AOI22_X1 U3598 ( .A1(\mem[81][5] ), .A2(n9992), .B1(n27049), .B2(data_in[5]), 
        .ZN(n9997) );
  INV_X1 U3599 ( .A(n9998), .ZN(n25452) );
  AOI22_X1 U3600 ( .A1(\mem[81][6] ), .A2(n9992), .B1(n27049), .B2(data_in[6]), 
        .ZN(n9998) );
  INV_X1 U3601 ( .A(n9999), .ZN(n25451) );
  AOI22_X1 U3602 ( .A1(\mem[81][7] ), .A2(n9992), .B1(n27049), .B2(data_in[7]), 
        .ZN(n9999) );
  INV_X1 U3603 ( .A(n10000), .ZN(n25450) );
  AOI22_X1 U3604 ( .A1(\mem[82][0] ), .A2(n10001), .B1(n27048), .B2(data_in[0]), .ZN(n10000) );
  INV_X1 U3605 ( .A(n10002), .ZN(n25449) );
  AOI22_X1 U3606 ( .A1(\mem[82][1] ), .A2(n10001), .B1(n27048), .B2(data_in[1]), .ZN(n10002) );
  INV_X1 U3607 ( .A(n10003), .ZN(n25448) );
  AOI22_X1 U3608 ( .A1(\mem[82][2] ), .A2(n10001), .B1(n27048), .B2(data_in[2]), .ZN(n10003) );
  INV_X1 U3609 ( .A(n10004), .ZN(n25447) );
  AOI22_X1 U3610 ( .A1(\mem[82][3] ), .A2(n10001), .B1(n27048), .B2(data_in[3]), .ZN(n10004) );
  INV_X1 U3611 ( .A(n10005), .ZN(n25446) );
  AOI22_X1 U3612 ( .A1(\mem[82][4] ), .A2(n10001), .B1(n27048), .B2(data_in[4]), .ZN(n10005) );
  INV_X1 U3613 ( .A(n10006), .ZN(n25445) );
  AOI22_X1 U3614 ( .A1(\mem[82][5] ), .A2(n10001), .B1(n27048), .B2(data_in[5]), .ZN(n10006) );
  INV_X1 U3615 ( .A(n10007), .ZN(n25444) );
  AOI22_X1 U3616 ( .A1(\mem[82][6] ), .A2(n10001), .B1(n27048), .B2(data_in[6]), .ZN(n10007) );
  INV_X1 U3617 ( .A(n10008), .ZN(n25443) );
  AOI22_X1 U3618 ( .A1(\mem[82][7] ), .A2(n10001), .B1(n27048), .B2(data_in[7]), .ZN(n10008) );
  INV_X1 U3619 ( .A(n10009), .ZN(n25442) );
  AOI22_X1 U3620 ( .A1(\mem[83][0] ), .A2(n10010), .B1(n27047), .B2(data_in[0]), .ZN(n10009) );
  INV_X1 U3621 ( .A(n10011), .ZN(n25441) );
  AOI22_X1 U3622 ( .A1(\mem[83][1] ), .A2(n10010), .B1(n27047), .B2(data_in[1]), .ZN(n10011) );
  INV_X1 U3623 ( .A(n10012), .ZN(n25440) );
  AOI22_X1 U3624 ( .A1(\mem[83][2] ), .A2(n10010), .B1(n27047), .B2(data_in[2]), .ZN(n10012) );
  INV_X1 U3625 ( .A(n10013), .ZN(n25439) );
  AOI22_X1 U3626 ( .A1(\mem[83][3] ), .A2(n10010), .B1(n27047), .B2(data_in[3]), .ZN(n10013) );
  INV_X1 U3627 ( .A(n10014), .ZN(n25438) );
  AOI22_X1 U3628 ( .A1(\mem[83][4] ), .A2(n10010), .B1(n27047), .B2(data_in[4]), .ZN(n10014) );
  INV_X1 U3629 ( .A(n10015), .ZN(n25437) );
  AOI22_X1 U3630 ( .A1(\mem[83][5] ), .A2(n10010), .B1(n27047), .B2(data_in[5]), .ZN(n10015) );
  INV_X1 U3631 ( .A(n10016), .ZN(n25436) );
  AOI22_X1 U3632 ( .A1(\mem[83][6] ), .A2(n10010), .B1(n27047), .B2(data_in[6]), .ZN(n10016) );
  INV_X1 U3633 ( .A(n10017), .ZN(n25435) );
  AOI22_X1 U3634 ( .A1(\mem[83][7] ), .A2(n10010), .B1(n27047), .B2(data_in[7]), .ZN(n10017) );
  INV_X1 U3635 ( .A(n10018), .ZN(n25434) );
  AOI22_X1 U3636 ( .A1(\mem[84][0] ), .A2(n10019), .B1(n27046), .B2(data_in[0]), .ZN(n10018) );
  INV_X1 U3637 ( .A(n10020), .ZN(n25433) );
  AOI22_X1 U3638 ( .A1(\mem[84][1] ), .A2(n10019), .B1(n27046), .B2(data_in[1]), .ZN(n10020) );
  INV_X1 U3639 ( .A(n10021), .ZN(n25432) );
  AOI22_X1 U3640 ( .A1(\mem[84][2] ), .A2(n10019), .B1(n27046), .B2(data_in[2]), .ZN(n10021) );
  INV_X1 U3641 ( .A(n10022), .ZN(n25431) );
  AOI22_X1 U3642 ( .A1(\mem[84][3] ), .A2(n10019), .B1(n27046), .B2(data_in[3]), .ZN(n10022) );
  INV_X1 U3643 ( .A(n10023), .ZN(n25430) );
  AOI22_X1 U3644 ( .A1(\mem[84][4] ), .A2(n10019), .B1(n27046), .B2(data_in[4]), .ZN(n10023) );
  INV_X1 U3645 ( .A(n10024), .ZN(n25429) );
  AOI22_X1 U3646 ( .A1(\mem[84][5] ), .A2(n10019), .B1(n27046), .B2(data_in[5]), .ZN(n10024) );
  INV_X1 U3647 ( .A(n10025), .ZN(n25428) );
  AOI22_X1 U3648 ( .A1(\mem[84][6] ), .A2(n10019), .B1(n27046), .B2(data_in[6]), .ZN(n10025) );
  INV_X1 U3649 ( .A(n10026), .ZN(n25427) );
  AOI22_X1 U3650 ( .A1(\mem[84][7] ), .A2(n10019), .B1(n27046), .B2(data_in[7]), .ZN(n10026) );
  INV_X1 U3651 ( .A(n10027), .ZN(n25426) );
  AOI22_X1 U3652 ( .A1(\mem[85][0] ), .A2(n10028), .B1(n27045), .B2(data_in[0]), .ZN(n10027) );
  INV_X1 U3653 ( .A(n10029), .ZN(n25425) );
  AOI22_X1 U3654 ( .A1(\mem[85][1] ), .A2(n10028), .B1(n27045), .B2(data_in[1]), .ZN(n10029) );
  INV_X1 U3655 ( .A(n10030), .ZN(n25424) );
  AOI22_X1 U3656 ( .A1(\mem[85][2] ), .A2(n10028), .B1(n27045), .B2(data_in[2]), .ZN(n10030) );
  INV_X1 U3657 ( .A(n10031), .ZN(n25423) );
  AOI22_X1 U3658 ( .A1(\mem[85][3] ), .A2(n10028), .B1(n27045), .B2(data_in[3]), .ZN(n10031) );
  INV_X1 U3659 ( .A(n10032), .ZN(n25422) );
  AOI22_X1 U3660 ( .A1(\mem[85][4] ), .A2(n10028), .B1(n27045), .B2(data_in[4]), .ZN(n10032) );
  INV_X1 U3661 ( .A(n10033), .ZN(n25421) );
  AOI22_X1 U3662 ( .A1(\mem[85][5] ), .A2(n10028), .B1(n27045), .B2(data_in[5]), .ZN(n10033) );
  INV_X1 U3663 ( .A(n10034), .ZN(n25420) );
  AOI22_X1 U3664 ( .A1(\mem[85][6] ), .A2(n10028), .B1(n27045), .B2(data_in[6]), .ZN(n10034) );
  INV_X1 U3665 ( .A(n10035), .ZN(n25419) );
  AOI22_X1 U3666 ( .A1(\mem[85][7] ), .A2(n10028), .B1(n27045), .B2(data_in[7]), .ZN(n10035) );
  INV_X1 U3667 ( .A(n10036), .ZN(n25418) );
  AOI22_X1 U3668 ( .A1(\mem[86][0] ), .A2(n10037), .B1(n27044), .B2(data_in[0]), .ZN(n10036) );
  INV_X1 U3669 ( .A(n10038), .ZN(n25417) );
  AOI22_X1 U3670 ( .A1(\mem[86][1] ), .A2(n10037), .B1(n27044), .B2(data_in[1]), .ZN(n10038) );
  INV_X1 U3671 ( .A(n10039), .ZN(n25416) );
  AOI22_X1 U3672 ( .A1(\mem[86][2] ), .A2(n10037), .B1(n27044), .B2(data_in[2]), .ZN(n10039) );
  INV_X1 U3673 ( .A(n10040), .ZN(n25415) );
  AOI22_X1 U3674 ( .A1(\mem[86][3] ), .A2(n10037), .B1(n27044), .B2(data_in[3]), .ZN(n10040) );
  INV_X1 U3675 ( .A(n10041), .ZN(n25414) );
  AOI22_X1 U3676 ( .A1(\mem[86][4] ), .A2(n10037), .B1(n27044), .B2(data_in[4]), .ZN(n10041) );
  INV_X1 U3677 ( .A(n10042), .ZN(n25413) );
  AOI22_X1 U3678 ( .A1(\mem[86][5] ), .A2(n10037), .B1(n27044), .B2(data_in[5]), .ZN(n10042) );
  INV_X1 U3679 ( .A(n10043), .ZN(n25412) );
  AOI22_X1 U3680 ( .A1(\mem[86][6] ), .A2(n10037), .B1(n27044), .B2(data_in[6]), .ZN(n10043) );
  INV_X1 U3681 ( .A(n10044), .ZN(n25411) );
  AOI22_X1 U3682 ( .A1(\mem[86][7] ), .A2(n10037), .B1(n27044), .B2(data_in[7]), .ZN(n10044) );
  INV_X1 U3683 ( .A(n10045), .ZN(n25410) );
  AOI22_X1 U3684 ( .A1(\mem[87][0] ), .A2(n10046), .B1(n27043), .B2(data_in[0]), .ZN(n10045) );
  INV_X1 U3685 ( .A(n10047), .ZN(n25409) );
  AOI22_X1 U3686 ( .A1(\mem[87][1] ), .A2(n10046), .B1(n27043), .B2(data_in[1]), .ZN(n10047) );
  INV_X1 U3687 ( .A(n10048), .ZN(n25408) );
  AOI22_X1 U3688 ( .A1(\mem[87][2] ), .A2(n10046), .B1(n27043), .B2(data_in[2]), .ZN(n10048) );
  INV_X1 U3689 ( .A(n10049), .ZN(n25407) );
  AOI22_X1 U3690 ( .A1(\mem[87][3] ), .A2(n10046), .B1(n27043), .B2(data_in[3]), .ZN(n10049) );
  INV_X1 U3691 ( .A(n10050), .ZN(n25406) );
  AOI22_X1 U3692 ( .A1(\mem[87][4] ), .A2(n10046), .B1(n27043), .B2(data_in[4]), .ZN(n10050) );
  INV_X1 U3693 ( .A(n10051), .ZN(n25405) );
  AOI22_X1 U3694 ( .A1(\mem[87][5] ), .A2(n10046), .B1(n27043), .B2(data_in[5]), .ZN(n10051) );
  INV_X1 U3695 ( .A(n10052), .ZN(n25404) );
  AOI22_X1 U3696 ( .A1(\mem[87][6] ), .A2(n10046), .B1(n27043), .B2(data_in[6]), .ZN(n10052) );
  INV_X1 U3697 ( .A(n10053), .ZN(n25403) );
  AOI22_X1 U3698 ( .A1(\mem[87][7] ), .A2(n10046), .B1(n27043), .B2(data_in[7]), .ZN(n10053) );
  INV_X1 U3699 ( .A(n10054), .ZN(n25402) );
  AOI22_X1 U3700 ( .A1(\mem[88][0] ), .A2(n10055), .B1(n27042), .B2(data_in[0]), .ZN(n10054) );
  INV_X1 U3701 ( .A(n10056), .ZN(n25401) );
  AOI22_X1 U3702 ( .A1(\mem[88][1] ), .A2(n10055), .B1(n27042), .B2(data_in[1]), .ZN(n10056) );
  INV_X1 U3703 ( .A(n10057), .ZN(n25400) );
  AOI22_X1 U3704 ( .A1(\mem[88][2] ), .A2(n10055), .B1(n27042), .B2(data_in[2]), .ZN(n10057) );
  INV_X1 U3705 ( .A(n10058), .ZN(n25399) );
  AOI22_X1 U3706 ( .A1(\mem[88][3] ), .A2(n10055), .B1(n27042), .B2(data_in[3]), .ZN(n10058) );
  INV_X1 U3707 ( .A(n10059), .ZN(n25398) );
  AOI22_X1 U3708 ( .A1(\mem[88][4] ), .A2(n10055), .B1(n27042), .B2(data_in[4]), .ZN(n10059) );
  INV_X1 U3709 ( .A(n10060), .ZN(n25397) );
  AOI22_X1 U3710 ( .A1(\mem[88][5] ), .A2(n10055), .B1(n27042), .B2(data_in[5]), .ZN(n10060) );
  INV_X1 U3711 ( .A(n10061), .ZN(n25396) );
  AOI22_X1 U3712 ( .A1(\mem[88][6] ), .A2(n10055), .B1(n27042), .B2(data_in[6]), .ZN(n10061) );
  INV_X1 U3713 ( .A(n10062), .ZN(n25395) );
  AOI22_X1 U3714 ( .A1(\mem[88][7] ), .A2(n10055), .B1(n27042), .B2(data_in[7]), .ZN(n10062) );
  INV_X1 U3715 ( .A(n10063), .ZN(n25394) );
  AOI22_X1 U3716 ( .A1(\mem[89][0] ), .A2(n10064), .B1(n27041), .B2(data_in[0]), .ZN(n10063) );
  INV_X1 U3717 ( .A(n10065), .ZN(n25393) );
  AOI22_X1 U3718 ( .A1(\mem[89][1] ), .A2(n10064), .B1(n27041), .B2(data_in[1]), .ZN(n10065) );
  INV_X1 U3719 ( .A(n10066), .ZN(n25392) );
  AOI22_X1 U3720 ( .A1(\mem[89][2] ), .A2(n10064), .B1(n27041), .B2(data_in[2]), .ZN(n10066) );
  INV_X1 U3721 ( .A(n10067), .ZN(n25391) );
  AOI22_X1 U3722 ( .A1(\mem[89][3] ), .A2(n10064), .B1(n27041), .B2(data_in[3]), .ZN(n10067) );
  INV_X1 U3723 ( .A(n10068), .ZN(n25390) );
  AOI22_X1 U3724 ( .A1(\mem[89][4] ), .A2(n10064), .B1(n27041), .B2(data_in[4]), .ZN(n10068) );
  INV_X1 U3725 ( .A(n10069), .ZN(n25389) );
  AOI22_X1 U3726 ( .A1(\mem[89][5] ), .A2(n10064), .B1(n27041), .B2(data_in[5]), .ZN(n10069) );
  INV_X1 U3727 ( .A(n10070), .ZN(n25388) );
  AOI22_X1 U3728 ( .A1(\mem[89][6] ), .A2(n10064), .B1(n27041), .B2(data_in[6]), .ZN(n10070) );
  INV_X1 U3729 ( .A(n10071), .ZN(n25387) );
  AOI22_X1 U3730 ( .A1(\mem[89][7] ), .A2(n10064), .B1(n27041), .B2(data_in[7]), .ZN(n10071) );
  INV_X1 U3731 ( .A(n10072), .ZN(n25386) );
  AOI22_X1 U3732 ( .A1(\mem[90][0] ), .A2(n10073), .B1(n27040), .B2(data_in[0]), .ZN(n10072) );
  INV_X1 U3733 ( .A(n10074), .ZN(n25385) );
  AOI22_X1 U3734 ( .A1(\mem[90][1] ), .A2(n10073), .B1(n27040), .B2(data_in[1]), .ZN(n10074) );
  INV_X1 U3735 ( .A(n10075), .ZN(n25384) );
  AOI22_X1 U3736 ( .A1(\mem[90][2] ), .A2(n10073), .B1(n27040), .B2(data_in[2]), .ZN(n10075) );
  INV_X1 U3737 ( .A(n10076), .ZN(n25383) );
  AOI22_X1 U3738 ( .A1(\mem[90][3] ), .A2(n10073), .B1(n27040), .B2(data_in[3]), .ZN(n10076) );
  INV_X1 U3739 ( .A(n10077), .ZN(n25382) );
  AOI22_X1 U3740 ( .A1(\mem[90][4] ), .A2(n10073), .B1(n27040), .B2(data_in[4]), .ZN(n10077) );
  INV_X1 U3741 ( .A(n10078), .ZN(n25381) );
  AOI22_X1 U3742 ( .A1(\mem[90][5] ), .A2(n10073), .B1(n27040), .B2(data_in[5]), .ZN(n10078) );
  INV_X1 U3743 ( .A(n10079), .ZN(n25380) );
  AOI22_X1 U3744 ( .A1(\mem[90][6] ), .A2(n10073), .B1(n27040), .B2(data_in[6]), .ZN(n10079) );
  INV_X1 U3745 ( .A(n10080), .ZN(n25379) );
  AOI22_X1 U3746 ( .A1(\mem[90][7] ), .A2(n10073), .B1(n27040), .B2(data_in[7]), .ZN(n10080) );
  INV_X1 U3747 ( .A(n10081), .ZN(n25378) );
  AOI22_X1 U3748 ( .A1(\mem[91][0] ), .A2(n10082), .B1(n27039), .B2(data_in[0]), .ZN(n10081) );
  INV_X1 U3749 ( .A(n10083), .ZN(n25377) );
  AOI22_X1 U3750 ( .A1(\mem[91][1] ), .A2(n10082), .B1(n27039), .B2(data_in[1]), .ZN(n10083) );
  INV_X1 U3751 ( .A(n10084), .ZN(n25376) );
  AOI22_X1 U3752 ( .A1(\mem[91][2] ), .A2(n10082), .B1(n27039), .B2(data_in[2]), .ZN(n10084) );
  INV_X1 U3753 ( .A(n10085), .ZN(n25375) );
  AOI22_X1 U3754 ( .A1(\mem[91][3] ), .A2(n10082), .B1(n27039), .B2(data_in[3]), .ZN(n10085) );
  INV_X1 U3755 ( .A(n10086), .ZN(n25374) );
  AOI22_X1 U3756 ( .A1(\mem[91][4] ), .A2(n10082), .B1(n27039), .B2(data_in[4]), .ZN(n10086) );
  INV_X1 U3757 ( .A(n10087), .ZN(n25373) );
  AOI22_X1 U3758 ( .A1(\mem[91][5] ), .A2(n10082), .B1(n27039), .B2(data_in[5]), .ZN(n10087) );
  INV_X1 U3759 ( .A(n10088), .ZN(n25372) );
  AOI22_X1 U3760 ( .A1(\mem[91][6] ), .A2(n10082), .B1(n27039), .B2(data_in[6]), .ZN(n10088) );
  INV_X1 U3761 ( .A(n10089), .ZN(n25371) );
  AOI22_X1 U3762 ( .A1(\mem[91][7] ), .A2(n10082), .B1(n27039), .B2(data_in[7]), .ZN(n10089) );
  INV_X1 U3763 ( .A(n10090), .ZN(n25370) );
  AOI22_X1 U3764 ( .A1(\mem[92][0] ), .A2(n10091), .B1(n27038), .B2(data_in[0]), .ZN(n10090) );
  INV_X1 U3765 ( .A(n10092), .ZN(n25369) );
  AOI22_X1 U3766 ( .A1(\mem[92][1] ), .A2(n10091), .B1(n27038), .B2(data_in[1]), .ZN(n10092) );
  INV_X1 U3767 ( .A(n10093), .ZN(n25368) );
  AOI22_X1 U3768 ( .A1(\mem[92][2] ), .A2(n10091), .B1(n27038), .B2(data_in[2]), .ZN(n10093) );
  INV_X1 U3769 ( .A(n10094), .ZN(n25367) );
  AOI22_X1 U3770 ( .A1(\mem[92][3] ), .A2(n10091), .B1(n27038), .B2(data_in[3]), .ZN(n10094) );
  INV_X1 U3771 ( .A(n10095), .ZN(n25366) );
  AOI22_X1 U3772 ( .A1(\mem[92][4] ), .A2(n10091), .B1(n27038), .B2(data_in[4]), .ZN(n10095) );
  INV_X1 U3773 ( .A(n10096), .ZN(n25365) );
  AOI22_X1 U3774 ( .A1(\mem[92][5] ), .A2(n10091), .B1(n27038), .B2(data_in[5]), .ZN(n10096) );
  INV_X1 U3775 ( .A(n10097), .ZN(n25364) );
  AOI22_X1 U3776 ( .A1(\mem[92][6] ), .A2(n10091), .B1(n27038), .B2(data_in[6]), .ZN(n10097) );
  INV_X1 U3777 ( .A(n10098), .ZN(n25363) );
  AOI22_X1 U3778 ( .A1(\mem[92][7] ), .A2(n10091), .B1(n27038), .B2(data_in[7]), .ZN(n10098) );
  INV_X1 U3779 ( .A(n10099), .ZN(n25362) );
  AOI22_X1 U3780 ( .A1(\mem[93][0] ), .A2(n10100), .B1(n27037), .B2(data_in[0]), .ZN(n10099) );
  INV_X1 U3781 ( .A(n10101), .ZN(n25361) );
  AOI22_X1 U3782 ( .A1(\mem[93][1] ), .A2(n10100), .B1(n27037), .B2(data_in[1]), .ZN(n10101) );
  INV_X1 U3783 ( .A(n10102), .ZN(n25360) );
  AOI22_X1 U3784 ( .A1(\mem[93][2] ), .A2(n10100), .B1(n27037), .B2(data_in[2]), .ZN(n10102) );
  INV_X1 U3785 ( .A(n10103), .ZN(n25359) );
  AOI22_X1 U3786 ( .A1(\mem[93][3] ), .A2(n10100), .B1(n27037), .B2(data_in[3]), .ZN(n10103) );
  INV_X1 U3787 ( .A(n10104), .ZN(n25358) );
  AOI22_X1 U3788 ( .A1(\mem[93][4] ), .A2(n10100), .B1(n27037), .B2(data_in[4]), .ZN(n10104) );
  INV_X1 U3789 ( .A(n10105), .ZN(n25357) );
  AOI22_X1 U3790 ( .A1(\mem[93][5] ), .A2(n10100), .B1(n27037), .B2(data_in[5]), .ZN(n10105) );
  INV_X1 U3791 ( .A(n10106), .ZN(n25356) );
  AOI22_X1 U3792 ( .A1(\mem[93][6] ), .A2(n10100), .B1(n27037), .B2(data_in[6]), .ZN(n10106) );
  INV_X1 U3793 ( .A(n10107), .ZN(n25355) );
  AOI22_X1 U3794 ( .A1(\mem[93][7] ), .A2(n10100), .B1(n27037), .B2(data_in[7]), .ZN(n10107) );
  INV_X1 U3795 ( .A(n10108), .ZN(n25354) );
  AOI22_X1 U3796 ( .A1(\mem[94][0] ), .A2(n10109), .B1(n27036), .B2(data_in[0]), .ZN(n10108) );
  INV_X1 U3797 ( .A(n10110), .ZN(n25353) );
  AOI22_X1 U3798 ( .A1(\mem[94][1] ), .A2(n10109), .B1(n27036), .B2(data_in[1]), .ZN(n10110) );
  INV_X1 U3799 ( .A(n10111), .ZN(n25352) );
  AOI22_X1 U3800 ( .A1(\mem[94][2] ), .A2(n10109), .B1(n27036), .B2(data_in[2]), .ZN(n10111) );
  INV_X1 U3801 ( .A(n10112), .ZN(n25351) );
  AOI22_X1 U3802 ( .A1(\mem[94][3] ), .A2(n10109), .B1(n27036), .B2(data_in[3]), .ZN(n10112) );
  INV_X1 U3803 ( .A(n10113), .ZN(n25350) );
  AOI22_X1 U3804 ( .A1(\mem[94][4] ), .A2(n10109), .B1(n27036), .B2(data_in[4]), .ZN(n10113) );
  INV_X1 U3805 ( .A(n10114), .ZN(n25349) );
  AOI22_X1 U3806 ( .A1(\mem[94][5] ), .A2(n10109), .B1(n27036), .B2(data_in[5]), .ZN(n10114) );
  INV_X1 U3807 ( .A(n10115), .ZN(n25348) );
  AOI22_X1 U3808 ( .A1(\mem[94][6] ), .A2(n10109), .B1(n27036), .B2(data_in[6]), .ZN(n10115) );
  INV_X1 U3809 ( .A(n10116), .ZN(n25347) );
  AOI22_X1 U3810 ( .A1(\mem[94][7] ), .A2(n10109), .B1(n27036), .B2(data_in[7]), .ZN(n10116) );
  INV_X1 U3811 ( .A(n10117), .ZN(n25346) );
  AOI22_X1 U3812 ( .A1(\mem[95][0] ), .A2(n10118), .B1(n27035), .B2(data_in[0]), .ZN(n10117) );
  INV_X1 U3813 ( .A(n10119), .ZN(n25345) );
  AOI22_X1 U3814 ( .A1(\mem[95][1] ), .A2(n10118), .B1(n27035), .B2(data_in[1]), .ZN(n10119) );
  INV_X1 U3815 ( .A(n10120), .ZN(n25344) );
  AOI22_X1 U3816 ( .A1(\mem[95][2] ), .A2(n10118), .B1(n27035), .B2(data_in[2]), .ZN(n10120) );
  INV_X1 U3817 ( .A(n10121), .ZN(n25343) );
  AOI22_X1 U3818 ( .A1(\mem[95][3] ), .A2(n10118), .B1(n27035), .B2(data_in[3]), .ZN(n10121) );
  INV_X1 U3819 ( .A(n10122), .ZN(n25342) );
  AOI22_X1 U3820 ( .A1(\mem[95][4] ), .A2(n10118), .B1(n27035), .B2(data_in[4]), .ZN(n10122) );
  INV_X1 U3821 ( .A(n10123), .ZN(n25341) );
  AOI22_X1 U3822 ( .A1(\mem[95][5] ), .A2(n10118), .B1(n27035), .B2(data_in[5]), .ZN(n10123) );
  INV_X1 U3823 ( .A(n10124), .ZN(n25340) );
  AOI22_X1 U3824 ( .A1(\mem[95][6] ), .A2(n10118), .B1(n27035), .B2(data_in[6]), .ZN(n10124) );
  INV_X1 U3825 ( .A(n10125), .ZN(n25339) );
  AOI22_X1 U3826 ( .A1(\mem[95][7] ), .A2(n10118), .B1(n27035), .B2(data_in[7]), .ZN(n10125) );
  INV_X1 U3827 ( .A(n10200), .ZN(n25274) );
  AOI22_X1 U3828 ( .A1(\mem[104][0] ), .A2(n10201), .B1(n27026), .B2(
        data_in[0]), .ZN(n10200) );
  INV_X1 U3829 ( .A(n10202), .ZN(n25273) );
  AOI22_X1 U3830 ( .A1(\mem[104][1] ), .A2(n10201), .B1(n27026), .B2(
        data_in[1]), .ZN(n10202) );
  INV_X1 U3831 ( .A(n10203), .ZN(n25272) );
  AOI22_X1 U3832 ( .A1(\mem[104][2] ), .A2(n10201), .B1(n27026), .B2(
        data_in[2]), .ZN(n10203) );
  INV_X1 U3833 ( .A(n10204), .ZN(n25271) );
  AOI22_X1 U3834 ( .A1(\mem[104][3] ), .A2(n10201), .B1(n27026), .B2(
        data_in[3]), .ZN(n10204) );
  INV_X1 U3835 ( .A(n10205), .ZN(n25270) );
  AOI22_X1 U3836 ( .A1(\mem[104][4] ), .A2(n10201), .B1(n27026), .B2(
        data_in[4]), .ZN(n10205) );
  INV_X1 U3837 ( .A(n10206), .ZN(n25269) );
  AOI22_X1 U3838 ( .A1(\mem[104][5] ), .A2(n10201), .B1(n27026), .B2(
        data_in[5]), .ZN(n10206) );
  INV_X1 U3839 ( .A(n10207), .ZN(n25268) );
  AOI22_X1 U3840 ( .A1(\mem[104][6] ), .A2(n10201), .B1(n27026), .B2(
        data_in[6]), .ZN(n10207) );
  INV_X1 U3841 ( .A(n10208), .ZN(n25267) );
  AOI22_X1 U3842 ( .A1(\mem[104][7] ), .A2(n10201), .B1(n27026), .B2(
        data_in[7]), .ZN(n10208) );
  INV_X1 U3843 ( .A(n10209), .ZN(n25266) );
  AOI22_X1 U3844 ( .A1(\mem[105][0] ), .A2(n10210), .B1(n27025), .B2(
        data_in[0]), .ZN(n10209) );
  INV_X1 U3845 ( .A(n10211), .ZN(n25265) );
  AOI22_X1 U3846 ( .A1(\mem[105][1] ), .A2(n10210), .B1(n27025), .B2(
        data_in[1]), .ZN(n10211) );
  INV_X1 U3847 ( .A(n10212), .ZN(n25264) );
  AOI22_X1 U3848 ( .A1(\mem[105][2] ), .A2(n10210), .B1(n27025), .B2(
        data_in[2]), .ZN(n10212) );
  INV_X1 U3849 ( .A(n10213), .ZN(n25263) );
  AOI22_X1 U3850 ( .A1(\mem[105][3] ), .A2(n10210), .B1(n27025), .B2(
        data_in[3]), .ZN(n10213) );
  INV_X1 U3851 ( .A(n10214), .ZN(n25262) );
  AOI22_X1 U3852 ( .A1(\mem[105][4] ), .A2(n10210), .B1(n27025), .B2(
        data_in[4]), .ZN(n10214) );
  INV_X1 U3853 ( .A(n10215), .ZN(n25261) );
  AOI22_X1 U3854 ( .A1(\mem[105][5] ), .A2(n10210), .B1(n27025), .B2(
        data_in[5]), .ZN(n10215) );
  INV_X1 U3855 ( .A(n10216), .ZN(n25260) );
  AOI22_X1 U3856 ( .A1(\mem[105][6] ), .A2(n10210), .B1(n27025), .B2(
        data_in[6]), .ZN(n10216) );
  INV_X1 U3857 ( .A(n10217), .ZN(n25259) );
  AOI22_X1 U3858 ( .A1(\mem[105][7] ), .A2(n10210), .B1(n27025), .B2(
        data_in[7]), .ZN(n10217) );
  INV_X1 U3859 ( .A(n10218), .ZN(n25258) );
  AOI22_X1 U3860 ( .A1(\mem[106][0] ), .A2(n10219), .B1(n27024), .B2(
        data_in[0]), .ZN(n10218) );
  INV_X1 U3861 ( .A(n10220), .ZN(n25257) );
  AOI22_X1 U3862 ( .A1(\mem[106][1] ), .A2(n10219), .B1(n27024), .B2(
        data_in[1]), .ZN(n10220) );
  INV_X1 U3863 ( .A(n10221), .ZN(n25256) );
  AOI22_X1 U3864 ( .A1(\mem[106][2] ), .A2(n10219), .B1(n27024), .B2(
        data_in[2]), .ZN(n10221) );
  INV_X1 U3865 ( .A(n10222), .ZN(n25255) );
  AOI22_X1 U3866 ( .A1(\mem[106][3] ), .A2(n10219), .B1(n27024), .B2(
        data_in[3]), .ZN(n10222) );
  INV_X1 U3867 ( .A(n10223), .ZN(n25254) );
  AOI22_X1 U3868 ( .A1(\mem[106][4] ), .A2(n10219), .B1(n27024), .B2(
        data_in[4]), .ZN(n10223) );
  INV_X1 U3869 ( .A(n10224), .ZN(n25253) );
  AOI22_X1 U3870 ( .A1(\mem[106][5] ), .A2(n10219), .B1(n27024), .B2(
        data_in[5]), .ZN(n10224) );
  INV_X1 U3871 ( .A(n10225), .ZN(n25252) );
  AOI22_X1 U3872 ( .A1(\mem[106][6] ), .A2(n10219), .B1(n27024), .B2(
        data_in[6]), .ZN(n10225) );
  INV_X1 U3873 ( .A(n10226), .ZN(n25251) );
  AOI22_X1 U3874 ( .A1(\mem[106][7] ), .A2(n10219), .B1(n27024), .B2(
        data_in[7]), .ZN(n10226) );
  INV_X1 U3875 ( .A(n10227), .ZN(n25250) );
  AOI22_X1 U3876 ( .A1(\mem[107][0] ), .A2(n10228), .B1(n27023), .B2(
        data_in[0]), .ZN(n10227) );
  INV_X1 U3877 ( .A(n10229), .ZN(n25249) );
  AOI22_X1 U3878 ( .A1(\mem[107][1] ), .A2(n10228), .B1(n27023), .B2(
        data_in[1]), .ZN(n10229) );
  INV_X1 U3879 ( .A(n10230), .ZN(n25248) );
  AOI22_X1 U3880 ( .A1(\mem[107][2] ), .A2(n10228), .B1(n27023), .B2(
        data_in[2]), .ZN(n10230) );
  INV_X1 U3881 ( .A(n10231), .ZN(n25247) );
  AOI22_X1 U3882 ( .A1(\mem[107][3] ), .A2(n10228), .B1(n27023), .B2(
        data_in[3]), .ZN(n10231) );
  INV_X1 U3883 ( .A(n10232), .ZN(n25246) );
  AOI22_X1 U3884 ( .A1(\mem[107][4] ), .A2(n10228), .B1(n27023), .B2(
        data_in[4]), .ZN(n10232) );
  INV_X1 U3885 ( .A(n10233), .ZN(n25245) );
  AOI22_X1 U3886 ( .A1(\mem[107][5] ), .A2(n10228), .B1(n27023), .B2(
        data_in[5]), .ZN(n10233) );
  INV_X1 U3887 ( .A(n10234), .ZN(n25244) );
  AOI22_X1 U3888 ( .A1(\mem[107][6] ), .A2(n10228), .B1(n27023), .B2(
        data_in[6]), .ZN(n10234) );
  INV_X1 U3889 ( .A(n10235), .ZN(n25243) );
  AOI22_X1 U3890 ( .A1(\mem[107][7] ), .A2(n10228), .B1(n27023), .B2(
        data_in[7]), .ZN(n10235) );
  INV_X1 U3891 ( .A(n10236), .ZN(n25242) );
  AOI22_X1 U3892 ( .A1(\mem[108][0] ), .A2(n10237), .B1(n27022), .B2(
        data_in[0]), .ZN(n10236) );
  INV_X1 U3893 ( .A(n10238), .ZN(n25241) );
  AOI22_X1 U3894 ( .A1(\mem[108][1] ), .A2(n10237), .B1(n27022), .B2(
        data_in[1]), .ZN(n10238) );
  INV_X1 U3895 ( .A(n10239), .ZN(n25240) );
  AOI22_X1 U3896 ( .A1(\mem[108][2] ), .A2(n10237), .B1(n27022), .B2(
        data_in[2]), .ZN(n10239) );
  INV_X1 U3897 ( .A(n10240), .ZN(n25239) );
  AOI22_X1 U3898 ( .A1(\mem[108][3] ), .A2(n10237), .B1(n27022), .B2(
        data_in[3]), .ZN(n10240) );
  INV_X1 U3899 ( .A(n10241), .ZN(n25238) );
  AOI22_X1 U3900 ( .A1(\mem[108][4] ), .A2(n10237), .B1(n27022), .B2(
        data_in[4]), .ZN(n10241) );
  INV_X1 U3901 ( .A(n10242), .ZN(n25237) );
  AOI22_X1 U3902 ( .A1(\mem[108][5] ), .A2(n10237), .B1(n27022), .B2(
        data_in[5]), .ZN(n10242) );
  INV_X1 U3903 ( .A(n10243), .ZN(n25236) );
  AOI22_X1 U3904 ( .A1(\mem[108][6] ), .A2(n10237), .B1(n27022), .B2(
        data_in[6]), .ZN(n10243) );
  INV_X1 U3905 ( .A(n10244), .ZN(n25235) );
  AOI22_X1 U3906 ( .A1(\mem[108][7] ), .A2(n10237), .B1(n27022), .B2(
        data_in[7]), .ZN(n10244) );
  INV_X1 U3907 ( .A(n10245), .ZN(n25234) );
  AOI22_X1 U3908 ( .A1(\mem[109][0] ), .A2(n10246), .B1(n27021), .B2(
        data_in[0]), .ZN(n10245) );
  INV_X1 U3909 ( .A(n10247), .ZN(n25233) );
  AOI22_X1 U3910 ( .A1(\mem[109][1] ), .A2(n10246), .B1(n27021), .B2(
        data_in[1]), .ZN(n10247) );
  INV_X1 U3911 ( .A(n10248), .ZN(n25232) );
  AOI22_X1 U3912 ( .A1(\mem[109][2] ), .A2(n10246), .B1(n27021), .B2(
        data_in[2]), .ZN(n10248) );
  INV_X1 U3913 ( .A(n10249), .ZN(n25231) );
  AOI22_X1 U3914 ( .A1(\mem[109][3] ), .A2(n10246), .B1(n27021), .B2(
        data_in[3]), .ZN(n10249) );
  INV_X1 U3915 ( .A(n10250), .ZN(n25230) );
  AOI22_X1 U3916 ( .A1(\mem[109][4] ), .A2(n10246), .B1(n27021), .B2(
        data_in[4]), .ZN(n10250) );
  INV_X1 U3917 ( .A(n10251), .ZN(n25229) );
  AOI22_X1 U3918 ( .A1(\mem[109][5] ), .A2(n10246), .B1(n27021), .B2(
        data_in[5]), .ZN(n10251) );
  INV_X1 U3919 ( .A(n10252), .ZN(n25228) );
  AOI22_X1 U3920 ( .A1(\mem[109][6] ), .A2(n10246), .B1(n27021), .B2(
        data_in[6]), .ZN(n10252) );
  INV_X1 U3921 ( .A(n10253), .ZN(n25227) );
  AOI22_X1 U3922 ( .A1(\mem[109][7] ), .A2(n10246), .B1(n27021), .B2(
        data_in[7]), .ZN(n10253) );
  INV_X1 U3923 ( .A(n10254), .ZN(n25226) );
  AOI22_X1 U3924 ( .A1(\mem[110][0] ), .A2(n10255), .B1(n27020), .B2(
        data_in[0]), .ZN(n10254) );
  INV_X1 U3925 ( .A(n10256), .ZN(n25225) );
  AOI22_X1 U3926 ( .A1(\mem[110][1] ), .A2(n10255), .B1(n27020), .B2(
        data_in[1]), .ZN(n10256) );
  INV_X1 U3927 ( .A(n10257), .ZN(n25224) );
  AOI22_X1 U3928 ( .A1(\mem[110][2] ), .A2(n10255), .B1(n27020), .B2(
        data_in[2]), .ZN(n10257) );
  INV_X1 U3929 ( .A(n10258), .ZN(n25223) );
  AOI22_X1 U3930 ( .A1(\mem[110][3] ), .A2(n10255), .B1(n27020), .B2(
        data_in[3]), .ZN(n10258) );
  INV_X1 U3931 ( .A(n10259), .ZN(n25222) );
  AOI22_X1 U3932 ( .A1(\mem[110][4] ), .A2(n10255), .B1(n27020), .B2(
        data_in[4]), .ZN(n10259) );
  INV_X1 U3933 ( .A(n10260), .ZN(n25221) );
  AOI22_X1 U3934 ( .A1(\mem[110][5] ), .A2(n10255), .B1(n27020), .B2(
        data_in[5]), .ZN(n10260) );
  INV_X1 U3935 ( .A(n10261), .ZN(n25220) );
  AOI22_X1 U3936 ( .A1(\mem[110][6] ), .A2(n10255), .B1(n27020), .B2(
        data_in[6]), .ZN(n10261) );
  INV_X1 U3937 ( .A(n10262), .ZN(n25219) );
  AOI22_X1 U3938 ( .A1(\mem[110][7] ), .A2(n10255), .B1(n27020), .B2(
        data_in[7]), .ZN(n10262) );
  INV_X1 U3939 ( .A(n10263), .ZN(n25218) );
  AOI22_X1 U3940 ( .A1(\mem[111][0] ), .A2(n10264), .B1(n27019), .B2(
        data_in[0]), .ZN(n10263) );
  INV_X1 U3941 ( .A(n10265), .ZN(n25217) );
  AOI22_X1 U3942 ( .A1(\mem[111][1] ), .A2(n10264), .B1(n27019), .B2(
        data_in[1]), .ZN(n10265) );
  INV_X1 U3943 ( .A(n10266), .ZN(n25216) );
  AOI22_X1 U3944 ( .A1(\mem[111][2] ), .A2(n10264), .B1(n27019), .B2(
        data_in[2]), .ZN(n10266) );
  INV_X1 U3945 ( .A(n10267), .ZN(n25215) );
  AOI22_X1 U3946 ( .A1(\mem[111][3] ), .A2(n10264), .B1(n27019), .B2(
        data_in[3]), .ZN(n10267) );
  INV_X1 U3947 ( .A(n10268), .ZN(n25214) );
  AOI22_X1 U3948 ( .A1(\mem[111][4] ), .A2(n10264), .B1(n27019), .B2(
        data_in[4]), .ZN(n10268) );
  INV_X1 U3949 ( .A(n10269), .ZN(n25213) );
  AOI22_X1 U3950 ( .A1(\mem[111][5] ), .A2(n10264), .B1(n27019), .B2(
        data_in[5]), .ZN(n10269) );
  INV_X1 U3951 ( .A(n10270), .ZN(n25212) );
  AOI22_X1 U3952 ( .A1(\mem[111][6] ), .A2(n10264), .B1(n27019), .B2(
        data_in[6]), .ZN(n10270) );
  INV_X1 U3953 ( .A(n10271), .ZN(n25211) );
  AOI22_X1 U3954 ( .A1(\mem[111][7] ), .A2(n10264), .B1(n27019), .B2(
        data_in[7]), .ZN(n10271) );
  INV_X1 U3955 ( .A(n10272), .ZN(n25210) );
  AOI22_X1 U3956 ( .A1(\mem[112][0] ), .A2(n10273), .B1(n27018), .B2(
        data_in[0]), .ZN(n10272) );
  INV_X1 U3957 ( .A(n10274), .ZN(n25209) );
  AOI22_X1 U3958 ( .A1(\mem[112][1] ), .A2(n10273), .B1(n27018), .B2(
        data_in[1]), .ZN(n10274) );
  INV_X1 U3959 ( .A(n10275), .ZN(n25208) );
  AOI22_X1 U3960 ( .A1(\mem[112][2] ), .A2(n10273), .B1(n27018), .B2(
        data_in[2]), .ZN(n10275) );
  INV_X1 U3961 ( .A(n10276), .ZN(n25207) );
  AOI22_X1 U3962 ( .A1(\mem[112][3] ), .A2(n10273), .B1(n27018), .B2(
        data_in[3]), .ZN(n10276) );
  INV_X1 U3963 ( .A(n10277), .ZN(n25206) );
  AOI22_X1 U3964 ( .A1(\mem[112][4] ), .A2(n10273), .B1(n27018), .B2(
        data_in[4]), .ZN(n10277) );
  INV_X1 U3965 ( .A(n10278), .ZN(n25205) );
  AOI22_X1 U3966 ( .A1(\mem[112][5] ), .A2(n10273), .B1(n27018), .B2(
        data_in[5]), .ZN(n10278) );
  INV_X1 U3967 ( .A(n10279), .ZN(n25204) );
  AOI22_X1 U3968 ( .A1(\mem[112][6] ), .A2(n10273), .B1(n27018), .B2(
        data_in[6]), .ZN(n10279) );
  INV_X1 U3969 ( .A(n10280), .ZN(n25203) );
  AOI22_X1 U3970 ( .A1(\mem[112][7] ), .A2(n10273), .B1(n27018), .B2(
        data_in[7]), .ZN(n10280) );
  INV_X1 U3971 ( .A(n10281), .ZN(n25202) );
  AOI22_X1 U3972 ( .A1(\mem[113][0] ), .A2(n10282), .B1(n27017), .B2(
        data_in[0]), .ZN(n10281) );
  INV_X1 U3973 ( .A(n10283), .ZN(n25201) );
  AOI22_X1 U3974 ( .A1(\mem[113][1] ), .A2(n10282), .B1(n27017), .B2(
        data_in[1]), .ZN(n10283) );
  INV_X1 U3975 ( .A(n10284), .ZN(n25200) );
  AOI22_X1 U3976 ( .A1(\mem[113][2] ), .A2(n10282), .B1(n27017), .B2(
        data_in[2]), .ZN(n10284) );
  INV_X1 U3977 ( .A(n10285), .ZN(n25199) );
  AOI22_X1 U3978 ( .A1(\mem[113][3] ), .A2(n10282), .B1(n27017), .B2(
        data_in[3]), .ZN(n10285) );
  INV_X1 U3979 ( .A(n10286), .ZN(n25198) );
  AOI22_X1 U3980 ( .A1(\mem[113][4] ), .A2(n10282), .B1(n27017), .B2(
        data_in[4]), .ZN(n10286) );
  INV_X1 U3981 ( .A(n10287), .ZN(n25197) );
  AOI22_X1 U3982 ( .A1(\mem[113][5] ), .A2(n10282), .B1(n27017), .B2(
        data_in[5]), .ZN(n10287) );
  INV_X1 U3983 ( .A(n10288), .ZN(n25196) );
  AOI22_X1 U3984 ( .A1(\mem[113][6] ), .A2(n10282), .B1(n27017), .B2(
        data_in[6]), .ZN(n10288) );
  INV_X1 U3985 ( .A(n10289), .ZN(n25195) );
  AOI22_X1 U3986 ( .A1(\mem[113][7] ), .A2(n10282), .B1(n27017), .B2(
        data_in[7]), .ZN(n10289) );
  INV_X1 U3987 ( .A(n10290), .ZN(n25194) );
  AOI22_X1 U3988 ( .A1(\mem[114][0] ), .A2(n10291), .B1(n27016), .B2(
        data_in[0]), .ZN(n10290) );
  INV_X1 U3989 ( .A(n10292), .ZN(n25193) );
  AOI22_X1 U3990 ( .A1(\mem[114][1] ), .A2(n10291), .B1(n27016), .B2(
        data_in[1]), .ZN(n10292) );
  INV_X1 U3991 ( .A(n10293), .ZN(n25192) );
  AOI22_X1 U3992 ( .A1(\mem[114][2] ), .A2(n10291), .B1(n27016), .B2(
        data_in[2]), .ZN(n10293) );
  INV_X1 U3993 ( .A(n10294), .ZN(n25191) );
  AOI22_X1 U3994 ( .A1(\mem[114][3] ), .A2(n10291), .B1(n27016), .B2(
        data_in[3]), .ZN(n10294) );
  INV_X1 U3995 ( .A(n10295), .ZN(n25190) );
  AOI22_X1 U3996 ( .A1(\mem[114][4] ), .A2(n10291), .B1(n27016), .B2(
        data_in[4]), .ZN(n10295) );
  INV_X1 U3997 ( .A(n10296), .ZN(n25189) );
  AOI22_X1 U3998 ( .A1(\mem[114][5] ), .A2(n10291), .B1(n27016), .B2(
        data_in[5]), .ZN(n10296) );
  INV_X1 U3999 ( .A(n10297), .ZN(n25188) );
  AOI22_X1 U4000 ( .A1(\mem[114][6] ), .A2(n10291), .B1(n27016), .B2(
        data_in[6]), .ZN(n10297) );
  INV_X1 U4001 ( .A(n10298), .ZN(n25187) );
  AOI22_X1 U4002 ( .A1(\mem[114][7] ), .A2(n10291), .B1(n27016), .B2(
        data_in[7]), .ZN(n10298) );
  INV_X1 U4003 ( .A(n10299), .ZN(n25186) );
  AOI22_X1 U4004 ( .A1(\mem[115][0] ), .A2(n10300), .B1(n27015), .B2(
        data_in[0]), .ZN(n10299) );
  INV_X1 U4005 ( .A(n10301), .ZN(n25185) );
  AOI22_X1 U4006 ( .A1(\mem[115][1] ), .A2(n10300), .B1(n27015), .B2(
        data_in[1]), .ZN(n10301) );
  INV_X1 U4007 ( .A(n10302), .ZN(n25184) );
  AOI22_X1 U4008 ( .A1(\mem[115][2] ), .A2(n10300), .B1(n27015), .B2(
        data_in[2]), .ZN(n10302) );
  INV_X1 U4009 ( .A(n10303), .ZN(n25183) );
  AOI22_X1 U4010 ( .A1(\mem[115][3] ), .A2(n10300), .B1(n27015), .B2(
        data_in[3]), .ZN(n10303) );
  INV_X1 U4011 ( .A(n10304), .ZN(n25182) );
  AOI22_X1 U4012 ( .A1(\mem[115][4] ), .A2(n10300), .B1(n27015), .B2(
        data_in[4]), .ZN(n10304) );
  INV_X1 U4013 ( .A(n10305), .ZN(n25181) );
  AOI22_X1 U4014 ( .A1(\mem[115][5] ), .A2(n10300), .B1(n27015), .B2(
        data_in[5]), .ZN(n10305) );
  INV_X1 U4015 ( .A(n10306), .ZN(n25180) );
  AOI22_X1 U4016 ( .A1(\mem[115][6] ), .A2(n10300), .B1(n27015), .B2(
        data_in[6]), .ZN(n10306) );
  INV_X1 U4017 ( .A(n10307), .ZN(n25179) );
  AOI22_X1 U4018 ( .A1(\mem[115][7] ), .A2(n10300), .B1(n27015), .B2(
        data_in[7]), .ZN(n10307) );
  INV_X1 U4019 ( .A(n10308), .ZN(n25178) );
  AOI22_X1 U4020 ( .A1(\mem[116][0] ), .A2(n10309), .B1(n27014), .B2(
        data_in[0]), .ZN(n10308) );
  INV_X1 U4021 ( .A(n10310), .ZN(n25177) );
  AOI22_X1 U4022 ( .A1(\mem[116][1] ), .A2(n10309), .B1(n27014), .B2(
        data_in[1]), .ZN(n10310) );
  INV_X1 U4023 ( .A(n10311), .ZN(n25176) );
  AOI22_X1 U4024 ( .A1(\mem[116][2] ), .A2(n10309), .B1(n27014), .B2(
        data_in[2]), .ZN(n10311) );
  INV_X1 U4025 ( .A(n10312), .ZN(n25175) );
  AOI22_X1 U4026 ( .A1(\mem[116][3] ), .A2(n10309), .B1(n27014), .B2(
        data_in[3]), .ZN(n10312) );
  INV_X1 U4027 ( .A(n10313), .ZN(n25174) );
  AOI22_X1 U4028 ( .A1(\mem[116][4] ), .A2(n10309), .B1(n27014), .B2(
        data_in[4]), .ZN(n10313) );
  INV_X1 U4029 ( .A(n10314), .ZN(n25173) );
  AOI22_X1 U4030 ( .A1(\mem[116][5] ), .A2(n10309), .B1(n27014), .B2(
        data_in[5]), .ZN(n10314) );
  INV_X1 U4031 ( .A(n10315), .ZN(n25172) );
  AOI22_X1 U4032 ( .A1(\mem[116][6] ), .A2(n10309), .B1(n27014), .B2(
        data_in[6]), .ZN(n10315) );
  INV_X1 U4033 ( .A(n10316), .ZN(n25171) );
  AOI22_X1 U4034 ( .A1(\mem[116][7] ), .A2(n10309), .B1(n27014), .B2(
        data_in[7]), .ZN(n10316) );
  INV_X1 U4035 ( .A(n10317), .ZN(n25170) );
  AOI22_X1 U4036 ( .A1(\mem[117][0] ), .A2(n10318), .B1(n27013), .B2(
        data_in[0]), .ZN(n10317) );
  INV_X1 U4037 ( .A(n10319), .ZN(n25169) );
  AOI22_X1 U4038 ( .A1(\mem[117][1] ), .A2(n10318), .B1(n27013), .B2(
        data_in[1]), .ZN(n10319) );
  INV_X1 U4039 ( .A(n10320), .ZN(n25168) );
  AOI22_X1 U4040 ( .A1(\mem[117][2] ), .A2(n10318), .B1(n27013), .B2(
        data_in[2]), .ZN(n10320) );
  INV_X1 U4041 ( .A(n10321), .ZN(n25167) );
  AOI22_X1 U4042 ( .A1(\mem[117][3] ), .A2(n10318), .B1(n27013), .B2(
        data_in[3]), .ZN(n10321) );
  INV_X1 U4043 ( .A(n10322), .ZN(n25166) );
  AOI22_X1 U4044 ( .A1(\mem[117][4] ), .A2(n10318), .B1(n27013), .B2(
        data_in[4]), .ZN(n10322) );
  INV_X1 U4045 ( .A(n10323), .ZN(n25165) );
  AOI22_X1 U4046 ( .A1(\mem[117][5] ), .A2(n10318), .B1(n27013), .B2(
        data_in[5]), .ZN(n10323) );
  INV_X1 U4047 ( .A(n10324), .ZN(n25164) );
  AOI22_X1 U4048 ( .A1(\mem[117][6] ), .A2(n10318), .B1(n27013), .B2(
        data_in[6]), .ZN(n10324) );
  INV_X1 U4049 ( .A(n10325), .ZN(n25163) );
  AOI22_X1 U4050 ( .A1(\mem[117][7] ), .A2(n10318), .B1(n27013), .B2(
        data_in[7]), .ZN(n10325) );
  INV_X1 U4051 ( .A(n10326), .ZN(n25162) );
  AOI22_X1 U4052 ( .A1(\mem[118][0] ), .A2(n10327), .B1(n27012), .B2(
        data_in[0]), .ZN(n10326) );
  INV_X1 U4053 ( .A(n10328), .ZN(n25161) );
  AOI22_X1 U4054 ( .A1(\mem[118][1] ), .A2(n10327), .B1(n27012), .B2(
        data_in[1]), .ZN(n10328) );
  INV_X1 U4055 ( .A(n10329), .ZN(n25160) );
  AOI22_X1 U4056 ( .A1(\mem[118][2] ), .A2(n10327), .B1(n27012), .B2(
        data_in[2]), .ZN(n10329) );
  INV_X1 U4057 ( .A(n10330), .ZN(n25159) );
  AOI22_X1 U4058 ( .A1(\mem[118][3] ), .A2(n10327), .B1(n27012), .B2(
        data_in[3]), .ZN(n10330) );
  INV_X1 U4059 ( .A(n10331), .ZN(n25158) );
  AOI22_X1 U4060 ( .A1(\mem[118][4] ), .A2(n10327), .B1(n27012), .B2(
        data_in[4]), .ZN(n10331) );
  INV_X1 U4061 ( .A(n10332), .ZN(n25157) );
  AOI22_X1 U4062 ( .A1(\mem[118][5] ), .A2(n10327), .B1(n27012), .B2(
        data_in[5]), .ZN(n10332) );
  INV_X1 U4063 ( .A(n10333), .ZN(n25156) );
  AOI22_X1 U4064 ( .A1(\mem[118][6] ), .A2(n10327), .B1(n27012), .B2(
        data_in[6]), .ZN(n10333) );
  INV_X1 U4065 ( .A(n10334), .ZN(n25155) );
  AOI22_X1 U4066 ( .A1(\mem[118][7] ), .A2(n10327), .B1(n27012), .B2(
        data_in[7]), .ZN(n10334) );
  INV_X1 U4067 ( .A(n10335), .ZN(n25154) );
  AOI22_X1 U4068 ( .A1(\mem[119][0] ), .A2(n10336), .B1(n27011), .B2(
        data_in[0]), .ZN(n10335) );
  INV_X1 U4069 ( .A(n10337), .ZN(n25153) );
  AOI22_X1 U4070 ( .A1(\mem[119][1] ), .A2(n10336), .B1(n27011), .B2(
        data_in[1]), .ZN(n10337) );
  INV_X1 U4071 ( .A(n10338), .ZN(n25152) );
  AOI22_X1 U4072 ( .A1(\mem[119][2] ), .A2(n10336), .B1(n27011), .B2(
        data_in[2]), .ZN(n10338) );
  INV_X1 U4073 ( .A(n10339), .ZN(n25151) );
  AOI22_X1 U4074 ( .A1(\mem[119][3] ), .A2(n10336), .B1(n27011), .B2(
        data_in[3]), .ZN(n10339) );
  INV_X1 U4075 ( .A(n10340), .ZN(n25150) );
  AOI22_X1 U4076 ( .A1(\mem[119][4] ), .A2(n10336), .B1(n27011), .B2(
        data_in[4]), .ZN(n10340) );
  INV_X1 U4077 ( .A(n10341), .ZN(n25149) );
  AOI22_X1 U4078 ( .A1(\mem[119][5] ), .A2(n10336), .B1(n27011), .B2(
        data_in[5]), .ZN(n10341) );
  INV_X1 U4079 ( .A(n10342), .ZN(n25148) );
  AOI22_X1 U4080 ( .A1(\mem[119][6] ), .A2(n10336), .B1(n27011), .B2(
        data_in[6]), .ZN(n10342) );
  INV_X1 U4081 ( .A(n10343), .ZN(n25147) );
  AOI22_X1 U4082 ( .A1(\mem[119][7] ), .A2(n10336), .B1(n27011), .B2(
        data_in[7]), .ZN(n10343) );
  INV_X1 U4083 ( .A(n10344), .ZN(n25146) );
  AOI22_X1 U4084 ( .A1(\mem[120][0] ), .A2(n10345), .B1(n27010), .B2(
        data_in[0]), .ZN(n10344) );
  INV_X1 U4085 ( .A(n10346), .ZN(n25145) );
  AOI22_X1 U4086 ( .A1(\mem[120][1] ), .A2(n10345), .B1(n27010), .B2(
        data_in[1]), .ZN(n10346) );
  INV_X1 U4087 ( .A(n10347), .ZN(n25144) );
  AOI22_X1 U4088 ( .A1(\mem[120][2] ), .A2(n10345), .B1(n27010), .B2(
        data_in[2]), .ZN(n10347) );
  INV_X1 U4089 ( .A(n10348), .ZN(n25143) );
  AOI22_X1 U4090 ( .A1(\mem[120][3] ), .A2(n10345), .B1(n27010), .B2(
        data_in[3]), .ZN(n10348) );
  INV_X1 U4091 ( .A(n10349), .ZN(n25142) );
  AOI22_X1 U4092 ( .A1(\mem[120][4] ), .A2(n10345), .B1(n27010), .B2(
        data_in[4]), .ZN(n10349) );
  INV_X1 U4093 ( .A(n10350), .ZN(n25141) );
  AOI22_X1 U4094 ( .A1(\mem[120][5] ), .A2(n10345), .B1(n27010), .B2(
        data_in[5]), .ZN(n10350) );
  INV_X1 U4095 ( .A(n10351), .ZN(n25140) );
  AOI22_X1 U4096 ( .A1(\mem[120][6] ), .A2(n10345), .B1(n27010), .B2(
        data_in[6]), .ZN(n10351) );
  INV_X1 U4097 ( .A(n10352), .ZN(n25139) );
  AOI22_X1 U4098 ( .A1(\mem[120][7] ), .A2(n10345), .B1(n27010), .B2(
        data_in[7]), .ZN(n10352) );
  INV_X1 U4099 ( .A(n10353), .ZN(n25138) );
  AOI22_X1 U4100 ( .A1(\mem[121][0] ), .A2(n10354), .B1(n27009), .B2(
        data_in[0]), .ZN(n10353) );
  INV_X1 U4101 ( .A(n10355), .ZN(n25137) );
  AOI22_X1 U4102 ( .A1(\mem[121][1] ), .A2(n10354), .B1(n27009), .B2(
        data_in[1]), .ZN(n10355) );
  INV_X1 U4103 ( .A(n10356), .ZN(n25136) );
  AOI22_X1 U4104 ( .A1(\mem[121][2] ), .A2(n10354), .B1(n27009), .B2(
        data_in[2]), .ZN(n10356) );
  INV_X1 U4105 ( .A(n10357), .ZN(n25135) );
  AOI22_X1 U4106 ( .A1(\mem[121][3] ), .A2(n10354), .B1(n27009), .B2(
        data_in[3]), .ZN(n10357) );
  INV_X1 U4107 ( .A(n10358), .ZN(n25134) );
  AOI22_X1 U4108 ( .A1(\mem[121][4] ), .A2(n10354), .B1(n27009), .B2(
        data_in[4]), .ZN(n10358) );
  INV_X1 U4109 ( .A(n10359), .ZN(n25133) );
  AOI22_X1 U4110 ( .A1(\mem[121][5] ), .A2(n10354), .B1(n27009), .B2(
        data_in[5]), .ZN(n10359) );
  INV_X1 U4111 ( .A(n10360), .ZN(n25132) );
  AOI22_X1 U4112 ( .A1(\mem[121][6] ), .A2(n10354), .B1(n27009), .B2(
        data_in[6]), .ZN(n10360) );
  INV_X1 U4113 ( .A(n10361), .ZN(n25131) );
  AOI22_X1 U4114 ( .A1(\mem[121][7] ), .A2(n10354), .B1(n27009), .B2(
        data_in[7]), .ZN(n10361) );
  INV_X1 U4115 ( .A(n10362), .ZN(n25130) );
  AOI22_X1 U4116 ( .A1(\mem[122][0] ), .A2(n10363), .B1(n27008), .B2(
        data_in[0]), .ZN(n10362) );
  INV_X1 U4117 ( .A(n10364), .ZN(n25129) );
  AOI22_X1 U4118 ( .A1(\mem[122][1] ), .A2(n10363), .B1(n27008), .B2(
        data_in[1]), .ZN(n10364) );
  INV_X1 U4119 ( .A(n10365), .ZN(n25128) );
  AOI22_X1 U4120 ( .A1(\mem[122][2] ), .A2(n10363), .B1(n27008), .B2(
        data_in[2]), .ZN(n10365) );
  INV_X1 U4121 ( .A(n10366), .ZN(n25127) );
  AOI22_X1 U4122 ( .A1(\mem[122][3] ), .A2(n10363), .B1(n27008), .B2(
        data_in[3]), .ZN(n10366) );
  INV_X1 U4123 ( .A(n10367), .ZN(n25126) );
  AOI22_X1 U4124 ( .A1(\mem[122][4] ), .A2(n10363), .B1(n27008), .B2(
        data_in[4]), .ZN(n10367) );
  INV_X1 U4125 ( .A(n10368), .ZN(n25125) );
  AOI22_X1 U4126 ( .A1(\mem[122][5] ), .A2(n10363), .B1(n27008), .B2(
        data_in[5]), .ZN(n10368) );
  INV_X1 U4127 ( .A(n10369), .ZN(n25124) );
  AOI22_X1 U4128 ( .A1(\mem[122][6] ), .A2(n10363), .B1(n27008), .B2(
        data_in[6]), .ZN(n10369) );
  INV_X1 U4129 ( .A(n10370), .ZN(n25123) );
  AOI22_X1 U4130 ( .A1(\mem[122][7] ), .A2(n10363), .B1(n27008), .B2(
        data_in[7]), .ZN(n10370) );
  INV_X1 U4131 ( .A(n10371), .ZN(n25122) );
  AOI22_X1 U4132 ( .A1(\mem[123][0] ), .A2(n10372), .B1(n27007), .B2(
        data_in[0]), .ZN(n10371) );
  INV_X1 U4133 ( .A(n10373), .ZN(n25121) );
  AOI22_X1 U4134 ( .A1(\mem[123][1] ), .A2(n10372), .B1(n27007), .B2(
        data_in[1]), .ZN(n10373) );
  INV_X1 U4135 ( .A(n10374), .ZN(n25120) );
  AOI22_X1 U4136 ( .A1(\mem[123][2] ), .A2(n10372), .B1(n27007), .B2(
        data_in[2]), .ZN(n10374) );
  INV_X1 U4137 ( .A(n10375), .ZN(n25119) );
  AOI22_X1 U4138 ( .A1(\mem[123][3] ), .A2(n10372), .B1(n27007), .B2(
        data_in[3]), .ZN(n10375) );
  INV_X1 U4139 ( .A(n10376), .ZN(n25118) );
  AOI22_X1 U4140 ( .A1(\mem[123][4] ), .A2(n10372), .B1(n27007), .B2(
        data_in[4]), .ZN(n10376) );
  INV_X1 U4141 ( .A(n10377), .ZN(n25117) );
  AOI22_X1 U4142 ( .A1(\mem[123][5] ), .A2(n10372), .B1(n27007), .B2(
        data_in[5]), .ZN(n10377) );
  INV_X1 U4143 ( .A(n10378), .ZN(n25116) );
  AOI22_X1 U4144 ( .A1(\mem[123][6] ), .A2(n10372), .B1(n27007), .B2(
        data_in[6]), .ZN(n10378) );
  INV_X1 U4145 ( .A(n10379), .ZN(n25115) );
  AOI22_X1 U4146 ( .A1(\mem[123][7] ), .A2(n10372), .B1(n27007), .B2(
        data_in[7]), .ZN(n10379) );
  INV_X1 U4147 ( .A(n10380), .ZN(n25114) );
  AOI22_X1 U4148 ( .A1(\mem[124][0] ), .A2(n10381), .B1(n27006), .B2(
        data_in[0]), .ZN(n10380) );
  INV_X1 U4149 ( .A(n10382), .ZN(n25113) );
  AOI22_X1 U4150 ( .A1(\mem[124][1] ), .A2(n10381), .B1(n27006), .B2(
        data_in[1]), .ZN(n10382) );
  INV_X1 U4151 ( .A(n10383), .ZN(n25112) );
  AOI22_X1 U4152 ( .A1(\mem[124][2] ), .A2(n10381), .B1(n27006), .B2(
        data_in[2]), .ZN(n10383) );
  INV_X1 U4153 ( .A(n10384), .ZN(n25111) );
  AOI22_X1 U4154 ( .A1(\mem[124][3] ), .A2(n10381), .B1(n27006), .B2(
        data_in[3]), .ZN(n10384) );
  INV_X1 U4155 ( .A(n10385), .ZN(n25110) );
  AOI22_X1 U4156 ( .A1(\mem[124][4] ), .A2(n10381), .B1(n27006), .B2(
        data_in[4]), .ZN(n10385) );
  INV_X1 U4157 ( .A(n10386), .ZN(n25109) );
  AOI22_X1 U4158 ( .A1(\mem[124][5] ), .A2(n10381), .B1(n27006), .B2(
        data_in[5]), .ZN(n10386) );
  INV_X1 U4159 ( .A(n10387), .ZN(n25108) );
  AOI22_X1 U4160 ( .A1(\mem[124][6] ), .A2(n10381), .B1(n27006), .B2(
        data_in[6]), .ZN(n10387) );
  INV_X1 U4161 ( .A(n10388), .ZN(n25107) );
  AOI22_X1 U4162 ( .A1(\mem[124][7] ), .A2(n10381), .B1(n27006), .B2(
        data_in[7]), .ZN(n10388) );
  INV_X1 U4163 ( .A(n10389), .ZN(n25106) );
  AOI22_X1 U4164 ( .A1(\mem[125][0] ), .A2(n10390), .B1(n27005), .B2(
        data_in[0]), .ZN(n10389) );
  INV_X1 U4165 ( .A(n10391), .ZN(n25105) );
  AOI22_X1 U4166 ( .A1(\mem[125][1] ), .A2(n10390), .B1(n27005), .B2(
        data_in[1]), .ZN(n10391) );
  INV_X1 U4167 ( .A(n10392), .ZN(n25104) );
  AOI22_X1 U4168 ( .A1(\mem[125][2] ), .A2(n10390), .B1(n27005), .B2(
        data_in[2]), .ZN(n10392) );
  INV_X1 U4169 ( .A(n10393), .ZN(n25103) );
  AOI22_X1 U4170 ( .A1(\mem[125][3] ), .A2(n10390), .B1(n27005), .B2(
        data_in[3]), .ZN(n10393) );
  INV_X1 U4171 ( .A(n10394), .ZN(n25102) );
  AOI22_X1 U4172 ( .A1(\mem[125][4] ), .A2(n10390), .B1(n27005), .B2(
        data_in[4]), .ZN(n10394) );
  INV_X1 U4173 ( .A(n10395), .ZN(n25101) );
  AOI22_X1 U4174 ( .A1(\mem[125][5] ), .A2(n10390), .B1(n27005), .B2(
        data_in[5]), .ZN(n10395) );
  INV_X1 U4175 ( .A(n10396), .ZN(n25100) );
  AOI22_X1 U4176 ( .A1(\mem[125][6] ), .A2(n10390), .B1(n27005), .B2(
        data_in[6]), .ZN(n10396) );
  INV_X1 U4177 ( .A(n10397), .ZN(n25099) );
  AOI22_X1 U4178 ( .A1(\mem[125][7] ), .A2(n10390), .B1(n27005), .B2(
        data_in[7]), .ZN(n10397) );
  INV_X1 U4179 ( .A(n10398), .ZN(n25098) );
  AOI22_X1 U4180 ( .A1(\mem[126][0] ), .A2(n10399), .B1(n27004), .B2(
        data_in[0]), .ZN(n10398) );
  INV_X1 U4181 ( .A(n10400), .ZN(n25097) );
  AOI22_X1 U4182 ( .A1(\mem[126][1] ), .A2(n10399), .B1(n27004), .B2(
        data_in[1]), .ZN(n10400) );
  INV_X1 U4183 ( .A(n10401), .ZN(n25096) );
  AOI22_X1 U4184 ( .A1(\mem[126][2] ), .A2(n10399), .B1(n27004), .B2(
        data_in[2]), .ZN(n10401) );
  INV_X1 U4185 ( .A(n10402), .ZN(n25095) );
  AOI22_X1 U4186 ( .A1(\mem[126][3] ), .A2(n10399), .B1(n27004), .B2(
        data_in[3]), .ZN(n10402) );
  INV_X1 U4187 ( .A(n10403), .ZN(n25094) );
  AOI22_X1 U4188 ( .A1(\mem[126][4] ), .A2(n10399), .B1(n27004), .B2(
        data_in[4]), .ZN(n10403) );
  INV_X1 U4189 ( .A(n10404), .ZN(n25093) );
  AOI22_X1 U4190 ( .A1(\mem[126][5] ), .A2(n10399), .B1(n27004), .B2(
        data_in[5]), .ZN(n10404) );
  INV_X1 U4191 ( .A(n10405), .ZN(n25092) );
  AOI22_X1 U4192 ( .A1(\mem[126][6] ), .A2(n10399), .B1(n27004), .B2(
        data_in[6]), .ZN(n10405) );
  INV_X1 U4193 ( .A(n10406), .ZN(n25091) );
  AOI22_X1 U4194 ( .A1(\mem[126][7] ), .A2(n10399), .B1(n27004), .B2(
        data_in[7]), .ZN(n10406) );
  INV_X1 U4195 ( .A(n10407), .ZN(n25090) );
  AOI22_X1 U4196 ( .A1(\mem[127][0] ), .A2(n10408), .B1(n27003), .B2(
        data_in[0]), .ZN(n10407) );
  INV_X1 U4197 ( .A(n10409), .ZN(n25089) );
  AOI22_X1 U4198 ( .A1(\mem[127][1] ), .A2(n10408), .B1(n27003), .B2(
        data_in[1]), .ZN(n10409) );
  INV_X1 U4199 ( .A(n10410), .ZN(n25088) );
  AOI22_X1 U4200 ( .A1(\mem[127][2] ), .A2(n10408), .B1(n27003), .B2(
        data_in[2]), .ZN(n10410) );
  INV_X1 U4201 ( .A(n10411), .ZN(n25087) );
  AOI22_X1 U4202 ( .A1(\mem[127][3] ), .A2(n10408), .B1(n27003), .B2(
        data_in[3]), .ZN(n10411) );
  INV_X1 U4203 ( .A(n10412), .ZN(n25086) );
  AOI22_X1 U4204 ( .A1(\mem[127][4] ), .A2(n10408), .B1(n27003), .B2(
        data_in[4]), .ZN(n10412) );
  INV_X1 U4205 ( .A(n10413), .ZN(n25085) );
  AOI22_X1 U4206 ( .A1(\mem[127][5] ), .A2(n10408), .B1(n27003), .B2(
        data_in[5]), .ZN(n10413) );
  INV_X1 U4207 ( .A(n10414), .ZN(n25084) );
  AOI22_X1 U4208 ( .A1(\mem[127][6] ), .A2(n10408), .B1(n27003), .B2(
        data_in[6]), .ZN(n10414) );
  INV_X1 U4209 ( .A(n10415), .ZN(n25083) );
  AOI22_X1 U4210 ( .A1(\mem[127][7] ), .A2(n10408), .B1(n27003), .B2(
        data_in[7]), .ZN(n10415) );
  INV_X1 U4211 ( .A(n10490), .ZN(n25018) );
  AOI22_X1 U4212 ( .A1(\mem[136][0] ), .A2(n10491), .B1(n26994), .B2(
        data_in[0]), .ZN(n10490) );
  INV_X1 U4213 ( .A(n10492), .ZN(n25017) );
  AOI22_X1 U4214 ( .A1(\mem[136][1] ), .A2(n10491), .B1(n26994), .B2(
        data_in[1]), .ZN(n10492) );
  INV_X1 U4215 ( .A(n10493), .ZN(n25016) );
  AOI22_X1 U4216 ( .A1(\mem[136][2] ), .A2(n10491), .B1(n26994), .B2(
        data_in[2]), .ZN(n10493) );
  INV_X1 U4217 ( .A(n10494), .ZN(n25015) );
  AOI22_X1 U4218 ( .A1(\mem[136][3] ), .A2(n10491), .B1(n26994), .B2(
        data_in[3]), .ZN(n10494) );
  INV_X1 U4219 ( .A(n10495), .ZN(n25014) );
  AOI22_X1 U4220 ( .A1(\mem[136][4] ), .A2(n10491), .B1(n26994), .B2(
        data_in[4]), .ZN(n10495) );
  INV_X1 U4221 ( .A(n10496), .ZN(n25013) );
  AOI22_X1 U4222 ( .A1(\mem[136][5] ), .A2(n10491), .B1(n26994), .B2(
        data_in[5]), .ZN(n10496) );
  INV_X1 U4223 ( .A(n10497), .ZN(n25012) );
  AOI22_X1 U4224 ( .A1(\mem[136][6] ), .A2(n10491), .B1(n26994), .B2(
        data_in[6]), .ZN(n10497) );
  INV_X1 U4225 ( .A(n10498), .ZN(n25011) );
  AOI22_X1 U4226 ( .A1(\mem[136][7] ), .A2(n10491), .B1(n26994), .B2(
        data_in[7]), .ZN(n10498) );
  INV_X1 U4227 ( .A(n10499), .ZN(n25010) );
  AOI22_X1 U4228 ( .A1(\mem[137][0] ), .A2(n10500), .B1(n26993), .B2(
        data_in[0]), .ZN(n10499) );
  INV_X1 U4229 ( .A(n10501), .ZN(n25009) );
  AOI22_X1 U4230 ( .A1(\mem[137][1] ), .A2(n10500), .B1(n26993), .B2(
        data_in[1]), .ZN(n10501) );
  INV_X1 U4231 ( .A(n10502), .ZN(n25008) );
  AOI22_X1 U4232 ( .A1(\mem[137][2] ), .A2(n10500), .B1(n26993), .B2(
        data_in[2]), .ZN(n10502) );
  INV_X1 U4233 ( .A(n10503), .ZN(n25007) );
  AOI22_X1 U4234 ( .A1(\mem[137][3] ), .A2(n10500), .B1(n26993), .B2(
        data_in[3]), .ZN(n10503) );
  INV_X1 U4235 ( .A(n10504), .ZN(n25006) );
  AOI22_X1 U4236 ( .A1(\mem[137][4] ), .A2(n10500), .B1(n26993), .B2(
        data_in[4]), .ZN(n10504) );
  INV_X1 U4237 ( .A(n10505), .ZN(n25005) );
  AOI22_X1 U4238 ( .A1(\mem[137][5] ), .A2(n10500), .B1(n26993), .B2(
        data_in[5]), .ZN(n10505) );
  INV_X1 U4239 ( .A(n10506), .ZN(n25004) );
  AOI22_X1 U4240 ( .A1(\mem[137][6] ), .A2(n10500), .B1(n26993), .B2(
        data_in[6]), .ZN(n10506) );
  INV_X1 U4241 ( .A(n10507), .ZN(n25003) );
  AOI22_X1 U4242 ( .A1(\mem[137][7] ), .A2(n10500), .B1(n26993), .B2(
        data_in[7]), .ZN(n10507) );
  INV_X1 U4243 ( .A(n10508), .ZN(n25002) );
  AOI22_X1 U4244 ( .A1(\mem[138][0] ), .A2(n10509), .B1(n26992), .B2(
        data_in[0]), .ZN(n10508) );
  INV_X1 U4245 ( .A(n10510), .ZN(n25001) );
  AOI22_X1 U4246 ( .A1(\mem[138][1] ), .A2(n10509), .B1(n26992), .B2(
        data_in[1]), .ZN(n10510) );
  INV_X1 U4247 ( .A(n10511), .ZN(n25000) );
  AOI22_X1 U4248 ( .A1(\mem[138][2] ), .A2(n10509), .B1(n26992), .B2(
        data_in[2]), .ZN(n10511) );
  INV_X1 U4249 ( .A(n10512), .ZN(n24999) );
  AOI22_X1 U4250 ( .A1(\mem[138][3] ), .A2(n10509), .B1(n26992), .B2(
        data_in[3]), .ZN(n10512) );
  INV_X1 U4251 ( .A(n10513), .ZN(n24998) );
  AOI22_X1 U4252 ( .A1(\mem[138][4] ), .A2(n10509), .B1(n26992), .B2(
        data_in[4]), .ZN(n10513) );
  INV_X1 U4253 ( .A(n10514), .ZN(n24997) );
  AOI22_X1 U4254 ( .A1(\mem[138][5] ), .A2(n10509), .B1(n26992), .B2(
        data_in[5]), .ZN(n10514) );
  INV_X1 U4255 ( .A(n10515), .ZN(n24996) );
  AOI22_X1 U4256 ( .A1(\mem[138][6] ), .A2(n10509), .B1(n26992), .B2(
        data_in[6]), .ZN(n10515) );
  INV_X1 U4257 ( .A(n10516), .ZN(n24995) );
  AOI22_X1 U4258 ( .A1(\mem[138][7] ), .A2(n10509), .B1(n26992), .B2(
        data_in[7]), .ZN(n10516) );
  INV_X1 U4259 ( .A(n10517), .ZN(n24994) );
  AOI22_X1 U4260 ( .A1(\mem[139][0] ), .A2(n10518), .B1(n26991), .B2(
        data_in[0]), .ZN(n10517) );
  INV_X1 U4261 ( .A(n10519), .ZN(n24993) );
  AOI22_X1 U4262 ( .A1(\mem[139][1] ), .A2(n10518), .B1(n26991), .B2(
        data_in[1]), .ZN(n10519) );
  INV_X1 U4263 ( .A(n10520), .ZN(n24992) );
  AOI22_X1 U4264 ( .A1(\mem[139][2] ), .A2(n10518), .B1(n26991), .B2(
        data_in[2]), .ZN(n10520) );
  INV_X1 U4265 ( .A(n10521), .ZN(n24991) );
  AOI22_X1 U4266 ( .A1(\mem[139][3] ), .A2(n10518), .B1(n26991), .B2(
        data_in[3]), .ZN(n10521) );
  INV_X1 U4267 ( .A(n10522), .ZN(n24990) );
  AOI22_X1 U4268 ( .A1(\mem[139][4] ), .A2(n10518), .B1(n26991), .B2(
        data_in[4]), .ZN(n10522) );
  INV_X1 U4269 ( .A(n10523), .ZN(n24989) );
  AOI22_X1 U4270 ( .A1(\mem[139][5] ), .A2(n10518), .B1(n26991), .B2(
        data_in[5]), .ZN(n10523) );
  INV_X1 U4271 ( .A(n10524), .ZN(n24988) );
  AOI22_X1 U4272 ( .A1(\mem[139][6] ), .A2(n10518), .B1(n26991), .B2(
        data_in[6]), .ZN(n10524) );
  INV_X1 U4273 ( .A(n10525), .ZN(n24987) );
  AOI22_X1 U4274 ( .A1(\mem[139][7] ), .A2(n10518), .B1(n26991), .B2(
        data_in[7]), .ZN(n10525) );
  INV_X1 U4275 ( .A(n10526), .ZN(n24986) );
  AOI22_X1 U4276 ( .A1(\mem[140][0] ), .A2(n10527), .B1(n26990), .B2(
        data_in[0]), .ZN(n10526) );
  INV_X1 U4277 ( .A(n10528), .ZN(n24985) );
  AOI22_X1 U4278 ( .A1(\mem[140][1] ), .A2(n10527), .B1(n26990), .B2(
        data_in[1]), .ZN(n10528) );
  INV_X1 U4279 ( .A(n10529), .ZN(n24984) );
  AOI22_X1 U4280 ( .A1(\mem[140][2] ), .A2(n10527), .B1(n26990), .B2(
        data_in[2]), .ZN(n10529) );
  INV_X1 U4281 ( .A(n10530), .ZN(n24983) );
  AOI22_X1 U4282 ( .A1(\mem[140][3] ), .A2(n10527), .B1(n26990), .B2(
        data_in[3]), .ZN(n10530) );
  INV_X1 U4283 ( .A(n10531), .ZN(n24982) );
  AOI22_X1 U4284 ( .A1(\mem[140][4] ), .A2(n10527), .B1(n26990), .B2(
        data_in[4]), .ZN(n10531) );
  INV_X1 U4285 ( .A(n10532), .ZN(n24981) );
  AOI22_X1 U4286 ( .A1(\mem[140][5] ), .A2(n10527), .B1(n26990), .B2(
        data_in[5]), .ZN(n10532) );
  INV_X1 U4287 ( .A(n10533), .ZN(n24980) );
  AOI22_X1 U4288 ( .A1(\mem[140][6] ), .A2(n10527), .B1(n26990), .B2(
        data_in[6]), .ZN(n10533) );
  INV_X1 U4289 ( .A(n10534), .ZN(n24979) );
  AOI22_X1 U4290 ( .A1(\mem[140][7] ), .A2(n10527), .B1(n26990), .B2(
        data_in[7]), .ZN(n10534) );
  INV_X1 U4291 ( .A(n10535), .ZN(n24978) );
  AOI22_X1 U4292 ( .A1(\mem[141][0] ), .A2(n10536), .B1(n26989), .B2(
        data_in[0]), .ZN(n10535) );
  INV_X1 U4293 ( .A(n10537), .ZN(n24977) );
  AOI22_X1 U4294 ( .A1(\mem[141][1] ), .A2(n10536), .B1(n26989), .B2(
        data_in[1]), .ZN(n10537) );
  INV_X1 U4295 ( .A(n10538), .ZN(n24976) );
  AOI22_X1 U4296 ( .A1(\mem[141][2] ), .A2(n10536), .B1(n26989), .B2(
        data_in[2]), .ZN(n10538) );
  INV_X1 U4297 ( .A(n10539), .ZN(n24975) );
  AOI22_X1 U4298 ( .A1(\mem[141][3] ), .A2(n10536), .B1(n26989), .B2(
        data_in[3]), .ZN(n10539) );
  INV_X1 U4299 ( .A(n10540), .ZN(n24974) );
  AOI22_X1 U4300 ( .A1(\mem[141][4] ), .A2(n10536), .B1(n26989), .B2(
        data_in[4]), .ZN(n10540) );
  INV_X1 U4301 ( .A(n10541), .ZN(n24973) );
  AOI22_X1 U4302 ( .A1(\mem[141][5] ), .A2(n10536), .B1(n26989), .B2(
        data_in[5]), .ZN(n10541) );
  INV_X1 U4303 ( .A(n10542), .ZN(n24972) );
  AOI22_X1 U4304 ( .A1(\mem[141][6] ), .A2(n10536), .B1(n26989), .B2(
        data_in[6]), .ZN(n10542) );
  INV_X1 U4305 ( .A(n10543), .ZN(n24971) );
  AOI22_X1 U4306 ( .A1(\mem[141][7] ), .A2(n10536), .B1(n26989), .B2(
        data_in[7]), .ZN(n10543) );
  INV_X1 U4307 ( .A(n10544), .ZN(n24970) );
  AOI22_X1 U4308 ( .A1(\mem[142][0] ), .A2(n10545), .B1(n26988), .B2(
        data_in[0]), .ZN(n10544) );
  INV_X1 U4309 ( .A(n10546), .ZN(n24969) );
  AOI22_X1 U4310 ( .A1(\mem[142][1] ), .A2(n10545), .B1(n26988), .B2(
        data_in[1]), .ZN(n10546) );
  INV_X1 U4311 ( .A(n10547), .ZN(n24968) );
  AOI22_X1 U4312 ( .A1(\mem[142][2] ), .A2(n10545), .B1(n26988), .B2(
        data_in[2]), .ZN(n10547) );
  INV_X1 U4313 ( .A(n10548), .ZN(n24967) );
  AOI22_X1 U4314 ( .A1(\mem[142][3] ), .A2(n10545), .B1(n26988), .B2(
        data_in[3]), .ZN(n10548) );
  INV_X1 U4315 ( .A(n10549), .ZN(n24966) );
  AOI22_X1 U4316 ( .A1(\mem[142][4] ), .A2(n10545), .B1(n26988), .B2(
        data_in[4]), .ZN(n10549) );
  INV_X1 U4317 ( .A(n10550), .ZN(n24965) );
  AOI22_X1 U4318 ( .A1(\mem[142][5] ), .A2(n10545), .B1(n26988), .B2(
        data_in[5]), .ZN(n10550) );
  INV_X1 U4319 ( .A(n10551), .ZN(n24964) );
  AOI22_X1 U4320 ( .A1(\mem[142][6] ), .A2(n10545), .B1(n26988), .B2(
        data_in[6]), .ZN(n10551) );
  INV_X1 U4321 ( .A(n10552), .ZN(n24963) );
  AOI22_X1 U4322 ( .A1(\mem[142][7] ), .A2(n10545), .B1(n26988), .B2(
        data_in[7]), .ZN(n10552) );
  INV_X1 U4323 ( .A(n10553), .ZN(n24962) );
  AOI22_X1 U4324 ( .A1(\mem[143][0] ), .A2(n10554), .B1(n26987), .B2(
        data_in[0]), .ZN(n10553) );
  INV_X1 U4325 ( .A(n10555), .ZN(n24961) );
  AOI22_X1 U4326 ( .A1(\mem[143][1] ), .A2(n10554), .B1(n26987), .B2(
        data_in[1]), .ZN(n10555) );
  INV_X1 U4327 ( .A(n10556), .ZN(n24960) );
  AOI22_X1 U4328 ( .A1(\mem[143][2] ), .A2(n10554), .B1(n26987), .B2(
        data_in[2]), .ZN(n10556) );
  INV_X1 U4329 ( .A(n10557), .ZN(n24959) );
  AOI22_X1 U4330 ( .A1(\mem[143][3] ), .A2(n10554), .B1(n26987), .B2(
        data_in[3]), .ZN(n10557) );
  INV_X1 U4331 ( .A(n10558), .ZN(n24958) );
  AOI22_X1 U4332 ( .A1(\mem[143][4] ), .A2(n10554), .B1(n26987), .B2(
        data_in[4]), .ZN(n10558) );
  INV_X1 U4333 ( .A(n10559), .ZN(n24957) );
  AOI22_X1 U4334 ( .A1(\mem[143][5] ), .A2(n10554), .B1(n26987), .B2(
        data_in[5]), .ZN(n10559) );
  INV_X1 U4335 ( .A(n10560), .ZN(n24956) );
  AOI22_X1 U4336 ( .A1(\mem[143][6] ), .A2(n10554), .B1(n26987), .B2(
        data_in[6]), .ZN(n10560) );
  INV_X1 U4337 ( .A(n10561), .ZN(n24955) );
  AOI22_X1 U4338 ( .A1(\mem[143][7] ), .A2(n10554), .B1(n26987), .B2(
        data_in[7]), .ZN(n10561) );
  INV_X1 U4339 ( .A(n10562), .ZN(n24954) );
  AOI22_X1 U4340 ( .A1(\mem[144][0] ), .A2(n10563), .B1(n26986), .B2(
        data_in[0]), .ZN(n10562) );
  INV_X1 U4341 ( .A(n10564), .ZN(n24953) );
  AOI22_X1 U4342 ( .A1(\mem[144][1] ), .A2(n10563), .B1(n26986), .B2(
        data_in[1]), .ZN(n10564) );
  INV_X1 U4343 ( .A(n10565), .ZN(n24952) );
  AOI22_X1 U4344 ( .A1(\mem[144][2] ), .A2(n10563), .B1(n26986), .B2(
        data_in[2]), .ZN(n10565) );
  INV_X1 U4345 ( .A(n10566), .ZN(n24951) );
  AOI22_X1 U4346 ( .A1(\mem[144][3] ), .A2(n10563), .B1(n26986), .B2(
        data_in[3]), .ZN(n10566) );
  INV_X1 U4347 ( .A(n10567), .ZN(n24950) );
  AOI22_X1 U4348 ( .A1(\mem[144][4] ), .A2(n10563), .B1(n26986), .B2(
        data_in[4]), .ZN(n10567) );
  INV_X1 U4349 ( .A(n10568), .ZN(n24949) );
  AOI22_X1 U4350 ( .A1(\mem[144][5] ), .A2(n10563), .B1(n26986), .B2(
        data_in[5]), .ZN(n10568) );
  INV_X1 U4351 ( .A(n10569), .ZN(n24948) );
  AOI22_X1 U4352 ( .A1(\mem[144][6] ), .A2(n10563), .B1(n26986), .B2(
        data_in[6]), .ZN(n10569) );
  INV_X1 U4353 ( .A(n10570), .ZN(n24947) );
  AOI22_X1 U4354 ( .A1(\mem[144][7] ), .A2(n10563), .B1(n26986), .B2(
        data_in[7]), .ZN(n10570) );
  INV_X1 U4355 ( .A(n10571), .ZN(n24946) );
  AOI22_X1 U4356 ( .A1(\mem[145][0] ), .A2(n10572), .B1(n26985), .B2(
        data_in[0]), .ZN(n10571) );
  INV_X1 U4357 ( .A(n10573), .ZN(n24945) );
  AOI22_X1 U4358 ( .A1(\mem[145][1] ), .A2(n10572), .B1(n26985), .B2(
        data_in[1]), .ZN(n10573) );
  INV_X1 U4359 ( .A(n10574), .ZN(n24944) );
  AOI22_X1 U4360 ( .A1(\mem[145][2] ), .A2(n10572), .B1(n26985), .B2(
        data_in[2]), .ZN(n10574) );
  INV_X1 U4361 ( .A(n10575), .ZN(n24943) );
  AOI22_X1 U4362 ( .A1(\mem[145][3] ), .A2(n10572), .B1(n26985), .B2(
        data_in[3]), .ZN(n10575) );
  INV_X1 U4363 ( .A(n10576), .ZN(n24942) );
  AOI22_X1 U4364 ( .A1(\mem[145][4] ), .A2(n10572), .B1(n26985), .B2(
        data_in[4]), .ZN(n10576) );
  INV_X1 U4365 ( .A(n10577), .ZN(n24941) );
  AOI22_X1 U4366 ( .A1(\mem[145][5] ), .A2(n10572), .B1(n26985), .B2(
        data_in[5]), .ZN(n10577) );
  INV_X1 U4367 ( .A(n10578), .ZN(n24940) );
  AOI22_X1 U4368 ( .A1(\mem[145][6] ), .A2(n10572), .B1(n26985), .B2(
        data_in[6]), .ZN(n10578) );
  INV_X1 U4369 ( .A(n10579), .ZN(n24939) );
  AOI22_X1 U4370 ( .A1(\mem[145][7] ), .A2(n10572), .B1(n26985), .B2(
        data_in[7]), .ZN(n10579) );
  INV_X1 U4371 ( .A(n10580), .ZN(n24938) );
  AOI22_X1 U4372 ( .A1(\mem[146][0] ), .A2(n10581), .B1(n26984), .B2(
        data_in[0]), .ZN(n10580) );
  INV_X1 U4373 ( .A(n10582), .ZN(n24937) );
  AOI22_X1 U4374 ( .A1(\mem[146][1] ), .A2(n10581), .B1(n26984), .B2(
        data_in[1]), .ZN(n10582) );
  INV_X1 U4375 ( .A(n10583), .ZN(n24936) );
  AOI22_X1 U4376 ( .A1(\mem[146][2] ), .A2(n10581), .B1(n26984), .B2(
        data_in[2]), .ZN(n10583) );
  INV_X1 U4377 ( .A(n10584), .ZN(n24935) );
  AOI22_X1 U4378 ( .A1(\mem[146][3] ), .A2(n10581), .B1(n26984), .B2(
        data_in[3]), .ZN(n10584) );
  INV_X1 U4379 ( .A(n10585), .ZN(n24934) );
  AOI22_X1 U4380 ( .A1(\mem[146][4] ), .A2(n10581), .B1(n26984), .B2(
        data_in[4]), .ZN(n10585) );
  INV_X1 U4381 ( .A(n10586), .ZN(n24933) );
  AOI22_X1 U4382 ( .A1(\mem[146][5] ), .A2(n10581), .B1(n26984), .B2(
        data_in[5]), .ZN(n10586) );
  INV_X1 U4383 ( .A(n10587), .ZN(n24932) );
  AOI22_X1 U4384 ( .A1(\mem[146][6] ), .A2(n10581), .B1(n26984), .B2(
        data_in[6]), .ZN(n10587) );
  INV_X1 U4385 ( .A(n10588), .ZN(n24931) );
  AOI22_X1 U4386 ( .A1(\mem[146][7] ), .A2(n10581), .B1(n26984), .B2(
        data_in[7]), .ZN(n10588) );
  INV_X1 U4387 ( .A(n10589), .ZN(n24930) );
  AOI22_X1 U4388 ( .A1(\mem[147][0] ), .A2(n10590), .B1(n26983), .B2(
        data_in[0]), .ZN(n10589) );
  INV_X1 U4389 ( .A(n10591), .ZN(n24929) );
  AOI22_X1 U4390 ( .A1(\mem[147][1] ), .A2(n10590), .B1(n26983), .B2(
        data_in[1]), .ZN(n10591) );
  INV_X1 U4391 ( .A(n10592), .ZN(n24928) );
  AOI22_X1 U4392 ( .A1(\mem[147][2] ), .A2(n10590), .B1(n26983), .B2(
        data_in[2]), .ZN(n10592) );
  INV_X1 U4393 ( .A(n10593), .ZN(n24927) );
  AOI22_X1 U4394 ( .A1(\mem[147][3] ), .A2(n10590), .B1(n26983), .B2(
        data_in[3]), .ZN(n10593) );
  INV_X1 U4395 ( .A(n10594), .ZN(n24926) );
  AOI22_X1 U4396 ( .A1(\mem[147][4] ), .A2(n10590), .B1(n26983), .B2(
        data_in[4]), .ZN(n10594) );
  INV_X1 U4397 ( .A(n10595), .ZN(n24925) );
  AOI22_X1 U4398 ( .A1(\mem[147][5] ), .A2(n10590), .B1(n26983), .B2(
        data_in[5]), .ZN(n10595) );
  INV_X1 U4399 ( .A(n10596), .ZN(n24924) );
  AOI22_X1 U4400 ( .A1(\mem[147][6] ), .A2(n10590), .B1(n26983), .B2(
        data_in[6]), .ZN(n10596) );
  INV_X1 U4401 ( .A(n10597), .ZN(n24923) );
  AOI22_X1 U4402 ( .A1(\mem[147][7] ), .A2(n10590), .B1(n26983), .B2(
        data_in[7]), .ZN(n10597) );
  INV_X1 U4403 ( .A(n10598), .ZN(n24922) );
  AOI22_X1 U4404 ( .A1(\mem[148][0] ), .A2(n10599), .B1(n26982), .B2(
        data_in[0]), .ZN(n10598) );
  INV_X1 U4405 ( .A(n10600), .ZN(n24921) );
  AOI22_X1 U4406 ( .A1(\mem[148][1] ), .A2(n10599), .B1(n26982), .B2(
        data_in[1]), .ZN(n10600) );
  INV_X1 U4407 ( .A(n10601), .ZN(n24920) );
  AOI22_X1 U4408 ( .A1(\mem[148][2] ), .A2(n10599), .B1(n26982), .B2(
        data_in[2]), .ZN(n10601) );
  INV_X1 U4409 ( .A(n10602), .ZN(n24919) );
  AOI22_X1 U4410 ( .A1(\mem[148][3] ), .A2(n10599), .B1(n26982), .B2(
        data_in[3]), .ZN(n10602) );
  INV_X1 U4411 ( .A(n10603), .ZN(n24918) );
  AOI22_X1 U4412 ( .A1(\mem[148][4] ), .A2(n10599), .B1(n26982), .B2(
        data_in[4]), .ZN(n10603) );
  INV_X1 U4413 ( .A(n10604), .ZN(n24917) );
  AOI22_X1 U4414 ( .A1(\mem[148][5] ), .A2(n10599), .B1(n26982), .B2(
        data_in[5]), .ZN(n10604) );
  INV_X1 U4415 ( .A(n10605), .ZN(n24916) );
  AOI22_X1 U4416 ( .A1(\mem[148][6] ), .A2(n10599), .B1(n26982), .B2(
        data_in[6]), .ZN(n10605) );
  INV_X1 U4417 ( .A(n10606), .ZN(n24915) );
  AOI22_X1 U4418 ( .A1(\mem[148][7] ), .A2(n10599), .B1(n26982), .B2(
        data_in[7]), .ZN(n10606) );
  INV_X1 U4419 ( .A(n10607), .ZN(n24914) );
  AOI22_X1 U4420 ( .A1(\mem[149][0] ), .A2(n10608), .B1(n26981), .B2(
        data_in[0]), .ZN(n10607) );
  INV_X1 U4421 ( .A(n10609), .ZN(n24913) );
  AOI22_X1 U4422 ( .A1(\mem[149][1] ), .A2(n10608), .B1(n26981), .B2(
        data_in[1]), .ZN(n10609) );
  INV_X1 U4423 ( .A(n10610), .ZN(n24912) );
  AOI22_X1 U4424 ( .A1(\mem[149][2] ), .A2(n10608), .B1(n26981), .B2(
        data_in[2]), .ZN(n10610) );
  INV_X1 U4425 ( .A(n10611), .ZN(n24911) );
  AOI22_X1 U4426 ( .A1(\mem[149][3] ), .A2(n10608), .B1(n26981), .B2(
        data_in[3]), .ZN(n10611) );
  INV_X1 U4427 ( .A(n10612), .ZN(n24910) );
  AOI22_X1 U4428 ( .A1(\mem[149][4] ), .A2(n10608), .B1(n26981), .B2(
        data_in[4]), .ZN(n10612) );
  INV_X1 U4429 ( .A(n10613), .ZN(n24909) );
  AOI22_X1 U4430 ( .A1(\mem[149][5] ), .A2(n10608), .B1(n26981), .B2(
        data_in[5]), .ZN(n10613) );
  INV_X1 U4431 ( .A(n10614), .ZN(n24908) );
  AOI22_X1 U4432 ( .A1(\mem[149][6] ), .A2(n10608), .B1(n26981), .B2(
        data_in[6]), .ZN(n10614) );
  INV_X1 U4433 ( .A(n10615), .ZN(n24907) );
  AOI22_X1 U4434 ( .A1(\mem[149][7] ), .A2(n10608), .B1(n26981), .B2(
        data_in[7]), .ZN(n10615) );
  INV_X1 U4435 ( .A(n10616), .ZN(n24906) );
  AOI22_X1 U4436 ( .A1(\mem[150][0] ), .A2(n10617), .B1(n26980), .B2(
        data_in[0]), .ZN(n10616) );
  INV_X1 U4437 ( .A(n10618), .ZN(n24905) );
  AOI22_X1 U4438 ( .A1(\mem[150][1] ), .A2(n10617), .B1(n26980), .B2(
        data_in[1]), .ZN(n10618) );
  INV_X1 U4439 ( .A(n10619), .ZN(n24904) );
  AOI22_X1 U4440 ( .A1(\mem[150][2] ), .A2(n10617), .B1(n26980), .B2(
        data_in[2]), .ZN(n10619) );
  INV_X1 U4441 ( .A(n10620), .ZN(n24903) );
  AOI22_X1 U4442 ( .A1(\mem[150][3] ), .A2(n10617), .B1(n26980), .B2(
        data_in[3]), .ZN(n10620) );
  INV_X1 U4443 ( .A(n10621), .ZN(n24902) );
  AOI22_X1 U4444 ( .A1(\mem[150][4] ), .A2(n10617), .B1(n26980), .B2(
        data_in[4]), .ZN(n10621) );
  INV_X1 U4445 ( .A(n10622), .ZN(n24901) );
  AOI22_X1 U4446 ( .A1(\mem[150][5] ), .A2(n10617), .B1(n26980), .B2(
        data_in[5]), .ZN(n10622) );
  INV_X1 U4447 ( .A(n10623), .ZN(n24900) );
  AOI22_X1 U4448 ( .A1(\mem[150][6] ), .A2(n10617), .B1(n26980), .B2(
        data_in[6]), .ZN(n10623) );
  INV_X1 U4449 ( .A(n10624), .ZN(n24899) );
  AOI22_X1 U4450 ( .A1(\mem[150][7] ), .A2(n10617), .B1(n26980), .B2(
        data_in[7]), .ZN(n10624) );
  INV_X1 U4451 ( .A(n10625), .ZN(n24898) );
  AOI22_X1 U4452 ( .A1(\mem[151][0] ), .A2(n10626), .B1(n26979), .B2(
        data_in[0]), .ZN(n10625) );
  INV_X1 U4453 ( .A(n10627), .ZN(n24897) );
  AOI22_X1 U4454 ( .A1(\mem[151][1] ), .A2(n10626), .B1(n26979), .B2(
        data_in[1]), .ZN(n10627) );
  INV_X1 U4455 ( .A(n10628), .ZN(n24896) );
  AOI22_X1 U4456 ( .A1(\mem[151][2] ), .A2(n10626), .B1(n26979), .B2(
        data_in[2]), .ZN(n10628) );
  INV_X1 U4457 ( .A(n10629), .ZN(n24895) );
  AOI22_X1 U4458 ( .A1(\mem[151][3] ), .A2(n10626), .B1(n26979), .B2(
        data_in[3]), .ZN(n10629) );
  INV_X1 U4459 ( .A(n10630), .ZN(n24894) );
  AOI22_X1 U4460 ( .A1(\mem[151][4] ), .A2(n10626), .B1(n26979), .B2(
        data_in[4]), .ZN(n10630) );
  INV_X1 U4461 ( .A(n10631), .ZN(n24893) );
  AOI22_X1 U4462 ( .A1(\mem[151][5] ), .A2(n10626), .B1(n26979), .B2(
        data_in[5]), .ZN(n10631) );
  INV_X1 U4463 ( .A(n10632), .ZN(n24892) );
  AOI22_X1 U4464 ( .A1(\mem[151][6] ), .A2(n10626), .B1(n26979), .B2(
        data_in[6]), .ZN(n10632) );
  INV_X1 U4465 ( .A(n10633), .ZN(n24891) );
  AOI22_X1 U4466 ( .A1(\mem[151][7] ), .A2(n10626), .B1(n26979), .B2(
        data_in[7]), .ZN(n10633) );
  INV_X1 U4467 ( .A(n10634), .ZN(n24890) );
  AOI22_X1 U4468 ( .A1(\mem[152][0] ), .A2(n10635), .B1(n26978), .B2(
        data_in[0]), .ZN(n10634) );
  INV_X1 U4469 ( .A(n10636), .ZN(n24889) );
  AOI22_X1 U4470 ( .A1(\mem[152][1] ), .A2(n10635), .B1(n26978), .B2(
        data_in[1]), .ZN(n10636) );
  INV_X1 U4471 ( .A(n10637), .ZN(n24888) );
  AOI22_X1 U4472 ( .A1(\mem[152][2] ), .A2(n10635), .B1(n26978), .B2(
        data_in[2]), .ZN(n10637) );
  INV_X1 U4473 ( .A(n10638), .ZN(n24887) );
  AOI22_X1 U4474 ( .A1(\mem[152][3] ), .A2(n10635), .B1(n26978), .B2(
        data_in[3]), .ZN(n10638) );
  INV_X1 U4475 ( .A(n10639), .ZN(n24886) );
  AOI22_X1 U4476 ( .A1(\mem[152][4] ), .A2(n10635), .B1(n26978), .B2(
        data_in[4]), .ZN(n10639) );
  INV_X1 U4477 ( .A(n10640), .ZN(n24885) );
  AOI22_X1 U4478 ( .A1(\mem[152][5] ), .A2(n10635), .B1(n26978), .B2(
        data_in[5]), .ZN(n10640) );
  INV_X1 U4479 ( .A(n10641), .ZN(n24884) );
  AOI22_X1 U4480 ( .A1(\mem[152][6] ), .A2(n10635), .B1(n26978), .B2(
        data_in[6]), .ZN(n10641) );
  INV_X1 U4481 ( .A(n10642), .ZN(n24883) );
  AOI22_X1 U4482 ( .A1(\mem[152][7] ), .A2(n10635), .B1(n26978), .B2(
        data_in[7]), .ZN(n10642) );
  INV_X1 U4483 ( .A(n10643), .ZN(n24882) );
  AOI22_X1 U4484 ( .A1(\mem[153][0] ), .A2(n10644), .B1(n26977), .B2(
        data_in[0]), .ZN(n10643) );
  INV_X1 U4485 ( .A(n10645), .ZN(n24881) );
  AOI22_X1 U4486 ( .A1(\mem[153][1] ), .A2(n10644), .B1(n26977), .B2(
        data_in[1]), .ZN(n10645) );
  INV_X1 U4487 ( .A(n10646), .ZN(n24880) );
  AOI22_X1 U4488 ( .A1(\mem[153][2] ), .A2(n10644), .B1(n26977), .B2(
        data_in[2]), .ZN(n10646) );
  INV_X1 U4489 ( .A(n10647), .ZN(n24879) );
  AOI22_X1 U4490 ( .A1(\mem[153][3] ), .A2(n10644), .B1(n26977), .B2(
        data_in[3]), .ZN(n10647) );
  INV_X1 U4491 ( .A(n10648), .ZN(n24878) );
  AOI22_X1 U4492 ( .A1(\mem[153][4] ), .A2(n10644), .B1(n26977), .B2(
        data_in[4]), .ZN(n10648) );
  INV_X1 U4493 ( .A(n10649), .ZN(n24877) );
  AOI22_X1 U4494 ( .A1(\mem[153][5] ), .A2(n10644), .B1(n26977), .B2(
        data_in[5]), .ZN(n10649) );
  INV_X1 U4495 ( .A(n10650), .ZN(n24876) );
  AOI22_X1 U4496 ( .A1(\mem[153][6] ), .A2(n10644), .B1(n26977), .B2(
        data_in[6]), .ZN(n10650) );
  INV_X1 U4497 ( .A(n10651), .ZN(n24875) );
  AOI22_X1 U4498 ( .A1(\mem[153][7] ), .A2(n10644), .B1(n26977), .B2(
        data_in[7]), .ZN(n10651) );
  INV_X1 U4499 ( .A(n10652), .ZN(n24874) );
  AOI22_X1 U4500 ( .A1(\mem[154][0] ), .A2(n10653), .B1(n26976), .B2(
        data_in[0]), .ZN(n10652) );
  INV_X1 U4501 ( .A(n10654), .ZN(n24873) );
  AOI22_X1 U4502 ( .A1(\mem[154][1] ), .A2(n10653), .B1(n26976), .B2(
        data_in[1]), .ZN(n10654) );
  INV_X1 U4503 ( .A(n10655), .ZN(n24872) );
  AOI22_X1 U4504 ( .A1(\mem[154][2] ), .A2(n10653), .B1(n26976), .B2(
        data_in[2]), .ZN(n10655) );
  INV_X1 U4505 ( .A(n10656), .ZN(n24871) );
  AOI22_X1 U4506 ( .A1(\mem[154][3] ), .A2(n10653), .B1(n26976), .B2(
        data_in[3]), .ZN(n10656) );
  INV_X1 U4507 ( .A(n10657), .ZN(n24870) );
  AOI22_X1 U4508 ( .A1(\mem[154][4] ), .A2(n10653), .B1(n26976), .B2(
        data_in[4]), .ZN(n10657) );
  INV_X1 U4509 ( .A(n10658), .ZN(n24869) );
  AOI22_X1 U4510 ( .A1(\mem[154][5] ), .A2(n10653), .B1(n26976), .B2(
        data_in[5]), .ZN(n10658) );
  INV_X1 U4511 ( .A(n10659), .ZN(n24868) );
  AOI22_X1 U4512 ( .A1(\mem[154][6] ), .A2(n10653), .B1(n26976), .B2(
        data_in[6]), .ZN(n10659) );
  INV_X1 U4513 ( .A(n10660), .ZN(n24867) );
  AOI22_X1 U4514 ( .A1(\mem[154][7] ), .A2(n10653), .B1(n26976), .B2(
        data_in[7]), .ZN(n10660) );
  INV_X1 U4515 ( .A(n10661), .ZN(n24866) );
  AOI22_X1 U4516 ( .A1(\mem[155][0] ), .A2(n10662), .B1(n26975), .B2(
        data_in[0]), .ZN(n10661) );
  INV_X1 U4517 ( .A(n10663), .ZN(n24865) );
  AOI22_X1 U4518 ( .A1(\mem[155][1] ), .A2(n10662), .B1(n26975), .B2(
        data_in[1]), .ZN(n10663) );
  INV_X1 U4519 ( .A(n10664), .ZN(n24864) );
  AOI22_X1 U4520 ( .A1(\mem[155][2] ), .A2(n10662), .B1(n26975), .B2(
        data_in[2]), .ZN(n10664) );
  INV_X1 U4521 ( .A(n10665), .ZN(n24863) );
  AOI22_X1 U4522 ( .A1(\mem[155][3] ), .A2(n10662), .B1(n26975), .B2(
        data_in[3]), .ZN(n10665) );
  INV_X1 U4523 ( .A(n10666), .ZN(n24862) );
  AOI22_X1 U4524 ( .A1(\mem[155][4] ), .A2(n10662), .B1(n26975), .B2(
        data_in[4]), .ZN(n10666) );
  INV_X1 U4525 ( .A(n10667), .ZN(n24861) );
  AOI22_X1 U4526 ( .A1(\mem[155][5] ), .A2(n10662), .B1(n26975), .B2(
        data_in[5]), .ZN(n10667) );
  INV_X1 U4527 ( .A(n10668), .ZN(n24860) );
  AOI22_X1 U4528 ( .A1(\mem[155][6] ), .A2(n10662), .B1(n26975), .B2(
        data_in[6]), .ZN(n10668) );
  INV_X1 U4529 ( .A(n10669), .ZN(n24859) );
  AOI22_X1 U4530 ( .A1(\mem[155][7] ), .A2(n10662), .B1(n26975), .B2(
        data_in[7]), .ZN(n10669) );
  INV_X1 U4531 ( .A(n10670), .ZN(n24858) );
  AOI22_X1 U4532 ( .A1(\mem[156][0] ), .A2(n10671), .B1(n26974), .B2(
        data_in[0]), .ZN(n10670) );
  INV_X1 U4533 ( .A(n10672), .ZN(n24857) );
  AOI22_X1 U4534 ( .A1(\mem[156][1] ), .A2(n10671), .B1(n26974), .B2(
        data_in[1]), .ZN(n10672) );
  INV_X1 U4535 ( .A(n10673), .ZN(n24856) );
  AOI22_X1 U4536 ( .A1(\mem[156][2] ), .A2(n10671), .B1(n26974), .B2(
        data_in[2]), .ZN(n10673) );
  INV_X1 U4537 ( .A(n10674), .ZN(n24855) );
  AOI22_X1 U4538 ( .A1(\mem[156][3] ), .A2(n10671), .B1(n26974), .B2(
        data_in[3]), .ZN(n10674) );
  INV_X1 U4539 ( .A(n10675), .ZN(n24854) );
  AOI22_X1 U4540 ( .A1(\mem[156][4] ), .A2(n10671), .B1(n26974), .B2(
        data_in[4]), .ZN(n10675) );
  INV_X1 U4541 ( .A(n10676), .ZN(n24853) );
  AOI22_X1 U4542 ( .A1(\mem[156][5] ), .A2(n10671), .B1(n26974), .B2(
        data_in[5]), .ZN(n10676) );
  INV_X1 U4543 ( .A(n10677), .ZN(n24852) );
  AOI22_X1 U4544 ( .A1(\mem[156][6] ), .A2(n10671), .B1(n26974), .B2(
        data_in[6]), .ZN(n10677) );
  INV_X1 U4545 ( .A(n10678), .ZN(n24851) );
  AOI22_X1 U4546 ( .A1(\mem[156][7] ), .A2(n10671), .B1(n26974), .B2(
        data_in[7]), .ZN(n10678) );
  INV_X1 U4547 ( .A(n10679), .ZN(n24850) );
  AOI22_X1 U4548 ( .A1(\mem[157][0] ), .A2(n10680), .B1(n26973), .B2(
        data_in[0]), .ZN(n10679) );
  INV_X1 U4549 ( .A(n10681), .ZN(n24849) );
  AOI22_X1 U4550 ( .A1(\mem[157][1] ), .A2(n10680), .B1(n26973), .B2(
        data_in[1]), .ZN(n10681) );
  INV_X1 U4551 ( .A(n10682), .ZN(n24848) );
  AOI22_X1 U4552 ( .A1(\mem[157][2] ), .A2(n10680), .B1(n26973), .B2(
        data_in[2]), .ZN(n10682) );
  INV_X1 U4553 ( .A(n10683), .ZN(n24847) );
  AOI22_X1 U4554 ( .A1(\mem[157][3] ), .A2(n10680), .B1(n26973), .B2(
        data_in[3]), .ZN(n10683) );
  INV_X1 U4555 ( .A(n10684), .ZN(n24846) );
  AOI22_X1 U4556 ( .A1(\mem[157][4] ), .A2(n10680), .B1(n26973), .B2(
        data_in[4]), .ZN(n10684) );
  INV_X1 U4557 ( .A(n10685), .ZN(n24845) );
  AOI22_X1 U4558 ( .A1(\mem[157][5] ), .A2(n10680), .B1(n26973), .B2(
        data_in[5]), .ZN(n10685) );
  INV_X1 U4559 ( .A(n10686), .ZN(n24844) );
  AOI22_X1 U4560 ( .A1(\mem[157][6] ), .A2(n10680), .B1(n26973), .B2(
        data_in[6]), .ZN(n10686) );
  INV_X1 U4561 ( .A(n10687), .ZN(n24843) );
  AOI22_X1 U4562 ( .A1(\mem[157][7] ), .A2(n10680), .B1(n26973), .B2(
        data_in[7]), .ZN(n10687) );
  INV_X1 U4563 ( .A(n10688), .ZN(n24842) );
  AOI22_X1 U4564 ( .A1(\mem[158][0] ), .A2(n10689), .B1(n26972), .B2(
        data_in[0]), .ZN(n10688) );
  INV_X1 U4565 ( .A(n10690), .ZN(n24841) );
  AOI22_X1 U4566 ( .A1(\mem[158][1] ), .A2(n10689), .B1(n26972), .B2(
        data_in[1]), .ZN(n10690) );
  INV_X1 U4567 ( .A(n10691), .ZN(n24840) );
  AOI22_X1 U4568 ( .A1(\mem[158][2] ), .A2(n10689), .B1(n26972), .B2(
        data_in[2]), .ZN(n10691) );
  INV_X1 U4569 ( .A(n10692), .ZN(n24839) );
  AOI22_X1 U4570 ( .A1(\mem[158][3] ), .A2(n10689), .B1(n26972), .B2(
        data_in[3]), .ZN(n10692) );
  INV_X1 U4571 ( .A(n10693), .ZN(n24838) );
  AOI22_X1 U4572 ( .A1(\mem[158][4] ), .A2(n10689), .B1(n26972), .B2(
        data_in[4]), .ZN(n10693) );
  INV_X1 U4573 ( .A(n10694), .ZN(n24837) );
  AOI22_X1 U4574 ( .A1(\mem[158][5] ), .A2(n10689), .B1(n26972), .B2(
        data_in[5]), .ZN(n10694) );
  INV_X1 U4575 ( .A(n10695), .ZN(n24836) );
  AOI22_X1 U4576 ( .A1(\mem[158][6] ), .A2(n10689), .B1(n26972), .B2(
        data_in[6]), .ZN(n10695) );
  INV_X1 U4577 ( .A(n10696), .ZN(n24835) );
  AOI22_X1 U4578 ( .A1(\mem[158][7] ), .A2(n10689), .B1(n26972), .B2(
        data_in[7]), .ZN(n10696) );
  INV_X1 U4579 ( .A(n10697), .ZN(n24834) );
  AOI22_X1 U4580 ( .A1(\mem[159][0] ), .A2(n10698), .B1(n26971), .B2(
        data_in[0]), .ZN(n10697) );
  INV_X1 U4581 ( .A(n10699), .ZN(n24833) );
  AOI22_X1 U4582 ( .A1(\mem[159][1] ), .A2(n10698), .B1(n26971), .B2(
        data_in[1]), .ZN(n10699) );
  INV_X1 U4583 ( .A(n10700), .ZN(n24832) );
  AOI22_X1 U4584 ( .A1(\mem[159][2] ), .A2(n10698), .B1(n26971), .B2(
        data_in[2]), .ZN(n10700) );
  INV_X1 U4585 ( .A(n10701), .ZN(n24831) );
  AOI22_X1 U4586 ( .A1(\mem[159][3] ), .A2(n10698), .B1(n26971), .B2(
        data_in[3]), .ZN(n10701) );
  INV_X1 U4587 ( .A(n10702), .ZN(n24830) );
  AOI22_X1 U4588 ( .A1(\mem[159][4] ), .A2(n10698), .B1(n26971), .B2(
        data_in[4]), .ZN(n10702) );
  INV_X1 U4589 ( .A(n10703), .ZN(n24829) );
  AOI22_X1 U4590 ( .A1(\mem[159][5] ), .A2(n10698), .B1(n26971), .B2(
        data_in[5]), .ZN(n10703) );
  INV_X1 U4591 ( .A(n10704), .ZN(n24828) );
  AOI22_X1 U4592 ( .A1(\mem[159][6] ), .A2(n10698), .B1(n26971), .B2(
        data_in[6]), .ZN(n10704) );
  INV_X1 U4593 ( .A(n10705), .ZN(n24827) );
  AOI22_X1 U4594 ( .A1(\mem[159][7] ), .A2(n10698), .B1(n26971), .B2(
        data_in[7]), .ZN(n10705) );
  INV_X1 U4595 ( .A(n10780), .ZN(n24762) );
  AOI22_X1 U4596 ( .A1(\mem[168][0] ), .A2(n10781), .B1(n26962), .B2(
        data_in[0]), .ZN(n10780) );
  INV_X1 U4597 ( .A(n10782), .ZN(n24761) );
  AOI22_X1 U4598 ( .A1(\mem[168][1] ), .A2(n10781), .B1(n26962), .B2(
        data_in[1]), .ZN(n10782) );
  INV_X1 U4599 ( .A(n10783), .ZN(n24760) );
  AOI22_X1 U4600 ( .A1(\mem[168][2] ), .A2(n10781), .B1(n26962), .B2(
        data_in[2]), .ZN(n10783) );
  INV_X1 U4601 ( .A(n10784), .ZN(n24759) );
  AOI22_X1 U4602 ( .A1(\mem[168][3] ), .A2(n10781), .B1(n26962), .B2(
        data_in[3]), .ZN(n10784) );
  INV_X1 U4603 ( .A(n10785), .ZN(n24758) );
  AOI22_X1 U4604 ( .A1(\mem[168][4] ), .A2(n10781), .B1(n26962), .B2(
        data_in[4]), .ZN(n10785) );
  INV_X1 U4605 ( .A(n10786), .ZN(n24757) );
  AOI22_X1 U4606 ( .A1(\mem[168][5] ), .A2(n10781), .B1(n26962), .B2(
        data_in[5]), .ZN(n10786) );
  INV_X1 U4607 ( .A(n10787), .ZN(n24756) );
  AOI22_X1 U4608 ( .A1(\mem[168][6] ), .A2(n10781), .B1(n26962), .B2(
        data_in[6]), .ZN(n10787) );
  INV_X1 U4609 ( .A(n10788), .ZN(n24755) );
  AOI22_X1 U4610 ( .A1(\mem[168][7] ), .A2(n10781), .B1(n26962), .B2(
        data_in[7]), .ZN(n10788) );
  INV_X1 U4611 ( .A(n10789), .ZN(n24754) );
  AOI22_X1 U4612 ( .A1(\mem[169][0] ), .A2(n10790), .B1(n26961), .B2(
        data_in[0]), .ZN(n10789) );
  INV_X1 U4613 ( .A(n10791), .ZN(n24753) );
  AOI22_X1 U4614 ( .A1(\mem[169][1] ), .A2(n10790), .B1(n26961), .B2(
        data_in[1]), .ZN(n10791) );
  INV_X1 U4615 ( .A(n10792), .ZN(n24752) );
  AOI22_X1 U4616 ( .A1(\mem[169][2] ), .A2(n10790), .B1(n26961), .B2(
        data_in[2]), .ZN(n10792) );
  INV_X1 U4617 ( .A(n10793), .ZN(n24751) );
  AOI22_X1 U4618 ( .A1(\mem[169][3] ), .A2(n10790), .B1(n26961), .B2(
        data_in[3]), .ZN(n10793) );
  INV_X1 U4619 ( .A(n10794), .ZN(n24750) );
  AOI22_X1 U4620 ( .A1(\mem[169][4] ), .A2(n10790), .B1(n26961), .B2(
        data_in[4]), .ZN(n10794) );
  INV_X1 U4621 ( .A(n10795), .ZN(n24749) );
  AOI22_X1 U4622 ( .A1(\mem[169][5] ), .A2(n10790), .B1(n26961), .B2(
        data_in[5]), .ZN(n10795) );
  INV_X1 U4623 ( .A(n10796), .ZN(n24748) );
  AOI22_X1 U4624 ( .A1(\mem[169][6] ), .A2(n10790), .B1(n26961), .B2(
        data_in[6]), .ZN(n10796) );
  INV_X1 U4625 ( .A(n10797), .ZN(n24747) );
  AOI22_X1 U4626 ( .A1(\mem[169][7] ), .A2(n10790), .B1(n26961), .B2(
        data_in[7]), .ZN(n10797) );
  INV_X1 U4627 ( .A(n10798), .ZN(n24746) );
  AOI22_X1 U4628 ( .A1(\mem[170][0] ), .A2(n10799), .B1(n26960), .B2(
        data_in[0]), .ZN(n10798) );
  INV_X1 U4629 ( .A(n10800), .ZN(n24745) );
  AOI22_X1 U4630 ( .A1(\mem[170][1] ), .A2(n10799), .B1(n26960), .B2(
        data_in[1]), .ZN(n10800) );
  INV_X1 U4631 ( .A(n10801), .ZN(n24744) );
  AOI22_X1 U4632 ( .A1(\mem[170][2] ), .A2(n10799), .B1(n26960), .B2(
        data_in[2]), .ZN(n10801) );
  INV_X1 U4633 ( .A(n10802), .ZN(n24743) );
  AOI22_X1 U4634 ( .A1(\mem[170][3] ), .A2(n10799), .B1(n26960), .B2(
        data_in[3]), .ZN(n10802) );
  INV_X1 U4635 ( .A(n10803), .ZN(n24742) );
  AOI22_X1 U4636 ( .A1(\mem[170][4] ), .A2(n10799), .B1(n26960), .B2(
        data_in[4]), .ZN(n10803) );
  INV_X1 U4637 ( .A(n10804), .ZN(n24741) );
  AOI22_X1 U4638 ( .A1(\mem[170][5] ), .A2(n10799), .B1(n26960), .B2(
        data_in[5]), .ZN(n10804) );
  INV_X1 U4639 ( .A(n10805), .ZN(n24740) );
  AOI22_X1 U4640 ( .A1(\mem[170][6] ), .A2(n10799), .B1(n26960), .B2(
        data_in[6]), .ZN(n10805) );
  INV_X1 U4641 ( .A(n10806), .ZN(n24739) );
  AOI22_X1 U4642 ( .A1(\mem[170][7] ), .A2(n10799), .B1(n26960), .B2(
        data_in[7]), .ZN(n10806) );
  INV_X1 U4643 ( .A(n10807), .ZN(n24738) );
  AOI22_X1 U4644 ( .A1(\mem[171][0] ), .A2(n10808), .B1(n26959), .B2(
        data_in[0]), .ZN(n10807) );
  INV_X1 U4645 ( .A(n10809), .ZN(n24737) );
  AOI22_X1 U4646 ( .A1(\mem[171][1] ), .A2(n10808), .B1(n26959), .B2(
        data_in[1]), .ZN(n10809) );
  INV_X1 U4647 ( .A(n10810), .ZN(n24736) );
  AOI22_X1 U4648 ( .A1(\mem[171][2] ), .A2(n10808), .B1(n26959), .B2(
        data_in[2]), .ZN(n10810) );
  INV_X1 U4649 ( .A(n10811), .ZN(n24735) );
  AOI22_X1 U4650 ( .A1(\mem[171][3] ), .A2(n10808), .B1(n26959), .B2(
        data_in[3]), .ZN(n10811) );
  INV_X1 U4651 ( .A(n10812), .ZN(n24734) );
  AOI22_X1 U4652 ( .A1(\mem[171][4] ), .A2(n10808), .B1(n26959), .B2(
        data_in[4]), .ZN(n10812) );
  INV_X1 U4653 ( .A(n10813), .ZN(n24733) );
  AOI22_X1 U4654 ( .A1(\mem[171][5] ), .A2(n10808), .B1(n26959), .B2(
        data_in[5]), .ZN(n10813) );
  INV_X1 U4655 ( .A(n10814), .ZN(n24732) );
  AOI22_X1 U4656 ( .A1(\mem[171][6] ), .A2(n10808), .B1(n26959), .B2(
        data_in[6]), .ZN(n10814) );
  INV_X1 U4657 ( .A(n10815), .ZN(n24731) );
  AOI22_X1 U4658 ( .A1(\mem[171][7] ), .A2(n10808), .B1(n26959), .B2(
        data_in[7]), .ZN(n10815) );
  INV_X1 U4659 ( .A(n10816), .ZN(n24730) );
  AOI22_X1 U4660 ( .A1(\mem[172][0] ), .A2(n10817), .B1(n26958), .B2(
        data_in[0]), .ZN(n10816) );
  INV_X1 U4661 ( .A(n10818), .ZN(n24729) );
  AOI22_X1 U4662 ( .A1(\mem[172][1] ), .A2(n10817), .B1(n26958), .B2(
        data_in[1]), .ZN(n10818) );
  INV_X1 U4663 ( .A(n10819), .ZN(n24728) );
  AOI22_X1 U4664 ( .A1(\mem[172][2] ), .A2(n10817), .B1(n26958), .B2(
        data_in[2]), .ZN(n10819) );
  INV_X1 U4665 ( .A(n10820), .ZN(n24727) );
  AOI22_X1 U4666 ( .A1(\mem[172][3] ), .A2(n10817), .B1(n26958), .B2(
        data_in[3]), .ZN(n10820) );
  INV_X1 U4667 ( .A(n10821), .ZN(n24726) );
  AOI22_X1 U4668 ( .A1(\mem[172][4] ), .A2(n10817), .B1(n26958), .B2(
        data_in[4]), .ZN(n10821) );
  INV_X1 U4669 ( .A(n10822), .ZN(n24725) );
  AOI22_X1 U4670 ( .A1(\mem[172][5] ), .A2(n10817), .B1(n26958), .B2(
        data_in[5]), .ZN(n10822) );
  INV_X1 U4671 ( .A(n10823), .ZN(n24724) );
  AOI22_X1 U4672 ( .A1(\mem[172][6] ), .A2(n10817), .B1(n26958), .B2(
        data_in[6]), .ZN(n10823) );
  INV_X1 U4673 ( .A(n10824), .ZN(n24723) );
  AOI22_X1 U4674 ( .A1(\mem[172][7] ), .A2(n10817), .B1(n26958), .B2(
        data_in[7]), .ZN(n10824) );
  INV_X1 U4675 ( .A(n10825), .ZN(n24722) );
  AOI22_X1 U4676 ( .A1(\mem[173][0] ), .A2(n10826), .B1(n26957), .B2(
        data_in[0]), .ZN(n10825) );
  INV_X1 U4677 ( .A(n10827), .ZN(n24721) );
  AOI22_X1 U4678 ( .A1(\mem[173][1] ), .A2(n10826), .B1(n26957), .B2(
        data_in[1]), .ZN(n10827) );
  INV_X1 U4679 ( .A(n10828), .ZN(n24720) );
  AOI22_X1 U4680 ( .A1(\mem[173][2] ), .A2(n10826), .B1(n26957), .B2(
        data_in[2]), .ZN(n10828) );
  INV_X1 U4681 ( .A(n10829), .ZN(n24719) );
  AOI22_X1 U4682 ( .A1(\mem[173][3] ), .A2(n10826), .B1(n26957), .B2(
        data_in[3]), .ZN(n10829) );
  INV_X1 U4683 ( .A(n10830), .ZN(n24718) );
  AOI22_X1 U4684 ( .A1(\mem[173][4] ), .A2(n10826), .B1(n26957), .B2(
        data_in[4]), .ZN(n10830) );
  INV_X1 U4685 ( .A(n10831), .ZN(n24717) );
  AOI22_X1 U4686 ( .A1(\mem[173][5] ), .A2(n10826), .B1(n26957), .B2(
        data_in[5]), .ZN(n10831) );
  INV_X1 U4687 ( .A(n10832), .ZN(n24716) );
  AOI22_X1 U4688 ( .A1(\mem[173][6] ), .A2(n10826), .B1(n26957), .B2(
        data_in[6]), .ZN(n10832) );
  INV_X1 U4689 ( .A(n10833), .ZN(n24715) );
  AOI22_X1 U4690 ( .A1(\mem[173][7] ), .A2(n10826), .B1(n26957), .B2(
        data_in[7]), .ZN(n10833) );
  INV_X1 U4691 ( .A(n10834), .ZN(n24714) );
  AOI22_X1 U4692 ( .A1(\mem[174][0] ), .A2(n10835), .B1(n26956), .B2(
        data_in[0]), .ZN(n10834) );
  INV_X1 U4693 ( .A(n10836), .ZN(n24713) );
  AOI22_X1 U4694 ( .A1(\mem[174][1] ), .A2(n10835), .B1(n26956), .B2(
        data_in[1]), .ZN(n10836) );
  INV_X1 U4695 ( .A(n10837), .ZN(n24712) );
  AOI22_X1 U4696 ( .A1(\mem[174][2] ), .A2(n10835), .B1(n26956), .B2(
        data_in[2]), .ZN(n10837) );
  INV_X1 U4697 ( .A(n10838), .ZN(n24711) );
  AOI22_X1 U4698 ( .A1(\mem[174][3] ), .A2(n10835), .B1(n26956), .B2(
        data_in[3]), .ZN(n10838) );
  INV_X1 U4699 ( .A(n10839), .ZN(n24710) );
  AOI22_X1 U4700 ( .A1(\mem[174][4] ), .A2(n10835), .B1(n26956), .B2(
        data_in[4]), .ZN(n10839) );
  INV_X1 U4701 ( .A(n10840), .ZN(n24709) );
  AOI22_X1 U4702 ( .A1(\mem[174][5] ), .A2(n10835), .B1(n26956), .B2(
        data_in[5]), .ZN(n10840) );
  INV_X1 U4703 ( .A(n10841), .ZN(n24708) );
  AOI22_X1 U4704 ( .A1(\mem[174][6] ), .A2(n10835), .B1(n26956), .B2(
        data_in[6]), .ZN(n10841) );
  INV_X1 U4705 ( .A(n10842), .ZN(n24707) );
  AOI22_X1 U4706 ( .A1(\mem[174][7] ), .A2(n10835), .B1(n26956), .B2(
        data_in[7]), .ZN(n10842) );
  INV_X1 U4707 ( .A(n10843), .ZN(n24706) );
  AOI22_X1 U4708 ( .A1(\mem[175][0] ), .A2(n10844), .B1(n26955), .B2(
        data_in[0]), .ZN(n10843) );
  INV_X1 U4709 ( .A(n10845), .ZN(n24705) );
  AOI22_X1 U4710 ( .A1(\mem[175][1] ), .A2(n10844), .B1(n26955), .B2(
        data_in[1]), .ZN(n10845) );
  INV_X1 U4711 ( .A(n10846), .ZN(n24704) );
  AOI22_X1 U4712 ( .A1(\mem[175][2] ), .A2(n10844), .B1(n26955), .B2(
        data_in[2]), .ZN(n10846) );
  INV_X1 U4713 ( .A(n10847), .ZN(n24703) );
  AOI22_X1 U4714 ( .A1(\mem[175][3] ), .A2(n10844), .B1(n26955), .B2(
        data_in[3]), .ZN(n10847) );
  INV_X1 U4715 ( .A(n10848), .ZN(n24702) );
  AOI22_X1 U4716 ( .A1(\mem[175][4] ), .A2(n10844), .B1(n26955), .B2(
        data_in[4]), .ZN(n10848) );
  INV_X1 U4717 ( .A(n10849), .ZN(n24701) );
  AOI22_X1 U4718 ( .A1(\mem[175][5] ), .A2(n10844), .B1(n26955), .B2(
        data_in[5]), .ZN(n10849) );
  INV_X1 U4719 ( .A(n10850), .ZN(n24700) );
  AOI22_X1 U4720 ( .A1(\mem[175][6] ), .A2(n10844), .B1(n26955), .B2(
        data_in[6]), .ZN(n10850) );
  INV_X1 U4721 ( .A(n10851), .ZN(n24699) );
  AOI22_X1 U4722 ( .A1(\mem[175][7] ), .A2(n10844), .B1(n26955), .B2(
        data_in[7]), .ZN(n10851) );
  INV_X1 U4723 ( .A(n10852), .ZN(n24698) );
  AOI22_X1 U4724 ( .A1(\mem[176][0] ), .A2(n10853), .B1(n26954), .B2(
        data_in[0]), .ZN(n10852) );
  INV_X1 U4725 ( .A(n10854), .ZN(n24697) );
  AOI22_X1 U4726 ( .A1(\mem[176][1] ), .A2(n10853), .B1(n26954), .B2(
        data_in[1]), .ZN(n10854) );
  INV_X1 U4727 ( .A(n10855), .ZN(n24696) );
  AOI22_X1 U4728 ( .A1(\mem[176][2] ), .A2(n10853), .B1(n26954), .B2(
        data_in[2]), .ZN(n10855) );
  INV_X1 U4729 ( .A(n10856), .ZN(n24695) );
  AOI22_X1 U4730 ( .A1(\mem[176][3] ), .A2(n10853), .B1(n26954), .B2(
        data_in[3]), .ZN(n10856) );
  INV_X1 U4731 ( .A(n10857), .ZN(n24694) );
  AOI22_X1 U4732 ( .A1(\mem[176][4] ), .A2(n10853), .B1(n26954), .B2(
        data_in[4]), .ZN(n10857) );
  INV_X1 U4733 ( .A(n10858), .ZN(n24693) );
  AOI22_X1 U4734 ( .A1(\mem[176][5] ), .A2(n10853), .B1(n26954), .B2(
        data_in[5]), .ZN(n10858) );
  INV_X1 U4735 ( .A(n10859), .ZN(n24692) );
  AOI22_X1 U4736 ( .A1(\mem[176][6] ), .A2(n10853), .B1(n26954), .B2(
        data_in[6]), .ZN(n10859) );
  INV_X1 U4737 ( .A(n10860), .ZN(n24691) );
  AOI22_X1 U4738 ( .A1(\mem[176][7] ), .A2(n10853), .B1(n26954), .B2(
        data_in[7]), .ZN(n10860) );
  INV_X1 U4739 ( .A(n10861), .ZN(n24690) );
  AOI22_X1 U4740 ( .A1(\mem[177][0] ), .A2(n10862), .B1(n26953), .B2(
        data_in[0]), .ZN(n10861) );
  INV_X1 U4741 ( .A(n10863), .ZN(n24689) );
  AOI22_X1 U4742 ( .A1(\mem[177][1] ), .A2(n10862), .B1(n26953), .B2(
        data_in[1]), .ZN(n10863) );
  INV_X1 U4743 ( .A(n10864), .ZN(n24688) );
  AOI22_X1 U4744 ( .A1(\mem[177][2] ), .A2(n10862), .B1(n26953), .B2(
        data_in[2]), .ZN(n10864) );
  INV_X1 U4745 ( .A(n10865), .ZN(n24687) );
  AOI22_X1 U4746 ( .A1(\mem[177][3] ), .A2(n10862), .B1(n26953), .B2(
        data_in[3]), .ZN(n10865) );
  INV_X1 U4747 ( .A(n10866), .ZN(n24686) );
  AOI22_X1 U4748 ( .A1(\mem[177][4] ), .A2(n10862), .B1(n26953), .B2(
        data_in[4]), .ZN(n10866) );
  INV_X1 U4749 ( .A(n10867), .ZN(n24685) );
  AOI22_X1 U4750 ( .A1(\mem[177][5] ), .A2(n10862), .B1(n26953), .B2(
        data_in[5]), .ZN(n10867) );
  INV_X1 U4751 ( .A(n10868), .ZN(n24684) );
  AOI22_X1 U4752 ( .A1(\mem[177][6] ), .A2(n10862), .B1(n26953), .B2(
        data_in[6]), .ZN(n10868) );
  INV_X1 U4753 ( .A(n10869), .ZN(n24683) );
  AOI22_X1 U4754 ( .A1(\mem[177][7] ), .A2(n10862), .B1(n26953), .B2(
        data_in[7]), .ZN(n10869) );
  INV_X1 U4755 ( .A(n10870), .ZN(n24682) );
  AOI22_X1 U4756 ( .A1(\mem[178][0] ), .A2(n10871), .B1(n26952), .B2(
        data_in[0]), .ZN(n10870) );
  INV_X1 U4757 ( .A(n10872), .ZN(n24681) );
  AOI22_X1 U4758 ( .A1(\mem[178][1] ), .A2(n10871), .B1(n26952), .B2(
        data_in[1]), .ZN(n10872) );
  INV_X1 U4759 ( .A(n10873), .ZN(n24680) );
  AOI22_X1 U4760 ( .A1(\mem[178][2] ), .A2(n10871), .B1(n26952), .B2(
        data_in[2]), .ZN(n10873) );
  INV_X1 U4761 ( .A(n10874), .ZN(n24679) );
  AOI22_X1 U4762 ( .A1(\mem[178][3] ), .A2(n10871), .B1(n26952), .B2(
        data_in[3]), .ZN(n10874) );
  INV_X1 U4763 ( .A(n10875), .ZN(n24678) );
  AOI22_X1 U4764 ( .A1(\mem[178][4] ), .A2(n10871), .B1(n26952), .B2(
        data_in[4]), .ZN(n10875) );
  INV_X1 U4765 ( .A(n10876), .ZN(n24677) );
  AOI22_X1 U4766 ( .A1(\mem[178][5] ), .A2(n10871), .B1(n26952), .B2(
        data_in[5]), .ZN(n10876) );
  INV_X1 U4767 ( .A(n10877), .ZN(n24676) );
  AOI22_X1 U4768 ( .A1(\mem[178][6] ), .A2(n10871), .B1(n26952), .B2(
        data_in[6]), .ZN(n10877) );
  INV_X1 U4769 ( .A(n10878), .ZN(n24675) );
  AOI22_X1 U4770 ( .A1(\mem[178][7] ), .A2(n10871), .B1(n26952), .B2(
        data_in[7]), .ZN(n10878) );
  INV_X1 U4771 ( .A(n10879), .ZN(n24674) );
  AOI22_X1 U4772 ( .A1(\mem[179][0] ), .A2(n10880), .B1(n26951), .B2(
        data_in[0]), .ZN(n10879) );
  INV_X1 U4773 ( .A(n10881), .ZN(n24673) );
  AOI22_X1 U4774 ( .A1(\mem[179][1] ), .A2(n10880), .B1(n26951), .B2(
        data_in[1]), .ZN(n10881) );
  INV_X1 U4775 ( .A(n10882), .ZN(n24672) );
  AOI22_X1 U4776 ( .A1(\mem[179][2] ), .A2(n10880), .B1(n26951), .B2(
        data_in[2]), .ZN(n10882) );
  INV_X1 U4777 ( .A(n10883), .ZN(n24671) );
  AOI22_X1 U4778 ( .A1(\mem[179][3] ), .A2(n10880), .B1(n26951), .B2(
        data_in[3]), .ZN(n10883) );
  INV_X1 U4779 ( .A(n10884), .ZN(n24670) );
  AOI22_X1 U4780 ( .A1(\mem[179][4] ), .A2(n10880), .B1(n26951), .B2(
        data_in[4]), .ZN(n10884) );
  INV_X1 U4781 ( .A(n10885), .ZN(n24669) );
  AOI22_X1 U4782 ( .A1(\mem[179][5] ), .A2(n10880), .B1(n26951), .B2(
        data_in[5]), .ZN(n10885) );
  INV_X1 U4783 ( .A(n10886), .ZN(n24668) );
  AOI22_X1 U4784 ( .A1(\mem[179][6] ), .A2(n10880), .B1(n26951), .B2(
        data_in[6]), .ZN(n10886) );
  INV_X1 U4785 ( .A(n10887), .ZN(n24667) );
  AOI22_X1 U4786 ( .A1(\mem[179][7] ), .A2(n10880), .B1(n26951), .B2(
        data_in[7]), .ZN(n10887) );
  INV_X1 U4787 ( .A(n10888), .ZN(n24666) );
  AOI22_X1 U4788 ( .A1(\mem[180][0] ), .A2(n10889), .B1(n26950), .B2(
        data_in[0]), .ZN(n10888) );
  INV_X1 U4789 ( .A(n10890), .ZN(n24665) );
  AOI22_X1 U4790 ( .A1(\mem[180][1] ), .A2(n10889), .B1(n26950), .B2(
        data_in[1]), .ZN(n10890) );
  INV_X1 U4791 ( .A(n10891), .ZN(n24664) );
  AOI22_X1 U4792 ( .A1(\mem[180][2] ), .A2(n10889), .B1(n26950), .B2(
        data_in[2]), .ZN(n10891) );
  INV_X1 U4793 ( .A(n10892), .ZN(n24663) );
  AOI22_X1 U4794 ( .A1(\mem[180][3] ), .A2(n10889), .B1(n26950), .B2(
        data_in[3]), .ZN(n10892) );
  INV_X1 U4795 ( .A(n10893), .ZN(n24662) );
  AOI22_X1 U4796 ( .A1(\mem[180][4] ), .A2(n10889), .B1(n26950), .B2(
        data_in[4]), .ZN(n10893) );
  INV_X1 U4797 ( .A(n10894), .ZN(n24661) );
  AOI22_X1 U4798 ( .A1(\mem[180][5] ), .A2(n10889), .B1(n26950), .B2(
        data_in[5]), .ZN(n10894) );
  INV_X1 U4799 ( .A(n10895), .ZN(n24660) );
  AOI22_X1 U4800 ( .A1(\mem[180][6] ), .A2(n10889), .B1(n26950), .B2(
        data_in[6]), .ZN(n10895) );
  INV_X1 U4801 ( .A(n10896), .ZN(n24659) );
  AOI22_X1 U4802 ( .A1(\mem[180][7] ), .A2(n10889), .B1(n26950), .B2(
        data_in[7]), .ZN(n10896) );
  INV_X1 U4803 ( .A(n10897), .ZN(n24658) );
  AOI22_X1 U4804 ( .A1(\mem[181][0] ), .A2(n10898), .B1(n26949), .B2(
        data_in[0]), .ZN(n10897) );
  INV_X1 U4805 ( .A(n10899), .ZN(n24657) );
  AOI22_X1 U4806 ( .A1(\mem[181][1] ), .A2(n10898), .B1(n26949), .B2(
        data_in[1]), .ZN(n10899) );
  INV_X1 U4807 ( .A(n10900), .ZN(n24656) );
  AOI22_X1 U4808 ( .A1(\mem[181][2] ), .A2(n10898), .B1(n26949), .B2(
        data_in[2]), .ZN(n10900) );
  INV_X1 U4809 ( .A(n10901), .ZN(n24655) );
  AOI22_X1 U4810 ( .A1(\mem[181][3] ), .A2(n10898), .B1(n26949), .B2(
        data_in[3]), .ZN(n10901) );
  INV_X1 U4811 ( .A(n10902), .ZN(n24654) );
  AOI22_X1 U4812 ( .A1(\mem[181][4] ), .A2(n10898), .B1(n26949), .B2(
        data_in[4]), .ZN(n10902) );
  INV_X1 U4813 ( .A(n10903), .ZN(n24653) );
  AOI22_X1 U4814 ( .A1(\mem[181][5] ), .A2(n10898), .B1(n26949), .B2(
        data_in[5]), .ZN(n10903) );
  INV_X1 U4815 ( .A(n10904), .ZN(n24652) );
  AOI22_X1 U4816 ( .A1(\mem[181][6] ), .A2(n10898), .B1(n26949), .B2(
        data_in[6]), .ZN(n10904) );
  INV_X1 U4817 ( .A(n10905), .ZN(n24651) );
  AOI22_X1 U4818 ( .A1(\mem[181][7] ), .A2(n10898), .B1(n26949), .B2(
        data_in[7]), .ZN(n10905) );
  INV_X1 U4819 ( .A(n10906), .ZN(n24650) );
  AOI22_X1 U4820 ( .A1(\mem[182][0] ), .A2(n10907), .B1(n26948), .B2(
        data_in[0]), .ZN(n10906) );
  INV_X1 U4821 ( .A(n10908), .ZN(n24649) );
  AOI22_X1 U4822 ( .A1(\mem[182][1] ), .A2(n10907), .B1(n26948), .B2(
        data_in[1]), .ZN(n10908) );
  INV_X1 U4823 ( .A(n10909), .ZN(n24648) );
  AOI22_X1 U4824 ( .A1(\mem[182][2] ), .A2(n10907), .B1(n26948), .B2(
        data_in[2]), .ZN(n10909) );
  INV_X1 U4825 ( .A(n10910), .ZN(n24647) );
  AOI22_X1 U4826 ( .A1(\mem[182][3] ), .A2(n10907), .B1(n26948), .B2(
        data_in[3]), .ZN(n10910) );
  INV_X1 U4827 ( .A(n10911), .ZN(n24646) );
  AOI22_X1 U4828 ( .A1(\mem[182][4] ), .A2(n10907), .B1(n26948), .B2(
        data_in[4]), .ZN(n10911) );
  INV_X1 U4829 ( .A(n10912), .ZN(n24645) );
  AOI22_X1 U4830 ( .A1(\mem[182][5] ), .A2(n10907), .B1(n26948), .B2(
        data_in[5]), .ZN(n10912) );
  INV_X1 U4831 ( .A(n10913), .ZN(n24644) );
  AOI22_X1 U4832 ( .A1(\mem[182][6] ), .A2(n10907), .B1(n26948), .B2(
        data_in[6]), .ZN(n10913) );
  INV_X1 U4833 ( .A(n10914), .ZN(n24643) );
  AOI22_X1 U4834 ( .A1(\mem[182][7] ), .A2(n10907), .B1(n26948), .B2(
        data_in[7]), .ZN(n10914) );
  INV_X1 U4835 ( .A(n10915), .ZN(n24642) );
  AOI22_X1 U4836 ( .A1(\mem[183][0] ), .A2(n10916), .B1(n26947), .B2(
        data_in[0]), .ZN(n10915) );
  INV_X1 U4837 ( .A(n10917), .ZN(n24641) );
  AOI22_X1 U4838 ( .A1(\mem[183][1] ), .A2(n10916), .B1(n26947), .B2(
        data_in[1]), .ZN(n10917) );
  INV_X1 U4839 ( .A(n10918), .ZN(n24640) );
  AOI22_X1 U4840 ( .A1(\mem[183][2] ), .A2(n10916), .B1(n26947), .B2(
        data_in[2]), .ZN(n10918) );
  INV_X1 U4841 ( .A(n10919), .ZN(n24639) );
  AOI22_X1 U4842 ( .A1(\mem[183][3] ), .A2(n10916), .B1(n26947), .B2(
        data_in[3]), .ZN(n10919) );
  INV_X1 U4843 ( .A(n10920), .ZN(n24638) );
  AOI22_X1 U4844 ( .A1(\mem[183][4] ), .A2(n10916), .B1(n26947), .B2(
        data_in[4]), .ZN(n10920) );
  INV_X1 U4845 ( .A(n10921), .ZN(n24637) );
  AOI22_X1 U4846 ( .A1(\mem[183][5] ), .A2(n10916), .B1(n26947), .B2(
        data_in[5]), .ZN(n10921) );
  INV_X1 U4847 ( .A(n10922), .ZN(n24636) );
  AOI22_X1 U4848 ( .A1(\mem[183][6] ), .A2(n10916), .B1(n26947), .B2(
        data_in[6]), .ZN(n10922) );
  INV_X1 U4849 ( .A(n10923), .ZN(n24635) );
  AOI22_X1 U4850 ( .A1(\mem[183][7] ), .A2(n10916), .B1(n26947), .B2(
        data_in[7]), .ZN(n10923) );
  INV_X1 U4851 ( .A(n10924), .ZN(n24634) );
  AOI22_X1 U4852 ( .A1(\mem[184][0] ), .A2(n10925), .B1(n26946), .B2(
        data_in[0]), .ZN(n10924) );
  INV_X1 U4853 ( .A(n10926), .ZN(n24633) );
  AOI22_X1 U4854 ( .A1(\mem[184][1] ), .A2(n10925), .B1(n26946), .B2(
        data_in[1]), .ZN(n10926) );
  INV_X1 U4855 ( .A(n10927), .ZN(n24632) );
  AOI22_X1 U4856 ( .A1(\mem[184][2] ), .A2(n10925), .B1(n26946), .B2(
        data_in[2]), .ZN(n10927) );
  INV_X1 U4857 ( .A(n10928), .ZN(n24631) );
  AOI22_X1 U4858 ( .A1(\mem[184][3] ), .A2(n10925), .B1(n26946), .B2(
        data_in[3]), .ZN(n10928) );
  INV_X1 U4859 ( .A(n10929), .ZN(n24630) );
  AOI22_X1 U4860 ( .A1(\mem[184][4] ), .A2(n10925), .B1(n26946), .B2(
        data_in[4]), .ZN(n10929) );
  INV_X1 U4861 ( .A(n10930), .ZN(n24629) );
  AOI22_X1 U4862 ( .A1(\mem[184][5] ), .A2(n10925), .B1(n26946), .B2(
        data_in[5]), .ZN(n10930) );
  INV_X1 U4863 ( .A(n10931), .ZN(n24628) );
  AOI22_X1 U4864 ( .A1(\mem[184][6] ), .A2(n10925), .B1(n26946), .B2(
        data_in[6]), .ZN(n10931) );
  INV_X1 U4865 ( .A(n10932), .ZN(n24627) );
  AOI22_X1 U4866 ( .A1(\mem[184][7] ), .A2(n10925), .B1(n26946), .B2(
        data_in[7]), .ZN(n10932) );
  INV_X1 U4867 ( .A(n10933), .ZN(n24626) );
  AOI22_X1 U4868 ( .A1(\mem[185][0] ), .A2(n10934), .B1(n26945), .B2(
        data_in[0]), .ZN(n10933) );
  INV_X1 U4869 ( .A(n10935), .ZN(n24625) );
  AOI22_X1 U4870 ( .A1(\mem[185][1] ), .A2(n10934), .B1(n26945), .B2(
        data_in[1]), .ZN(n10935) );
  INV_X1 U4871 ( .A(n10936), .ZN(n24624) );
  AOI22_X1 U4872 ( .A1(\mem[185][2] ), .A2(n10934), .B1(n26945), .B2(
        data_in[2]), .ZN(n10936) );
  INV_X1 U4873 ( .A(n10937), .ZN(n24623) );
  AOI22_X1 U4874 ( .A1(\mem[185][3] ), .A2(n10934), .B1(n26945), .B2(
        data_in[3]), .ZN(n10937) );
  INV_X1 U4875 ( .A(n10938), .ZN(n24622) );
  AOI22_X1 U4876 ( .A1(\mem[185][4] ), .A2(n10934), .B1(n26945), .B2(
        data_in[4]), .ZN(n10938) );
  INV_X1 U4877 ( .A(n10939), .ZN(n24621) );
  AOI22_X1 U4878 ( .A1(\mem[185][5] ), .A2(n10934), .B1(n26945), .B2(
        data_in[5]), .ZN(n10939) );
  INV_X1 U4879 ( .A(n10940), .ZN(n24620) );
  AOI22_X1 U4880 ( .A1(\mem[185][6] ), .A2(n10934), .B1(n26945), .B2(
        data_in[6]), .ZN(n10940) );
  INV_X1 U4881 ( .A(n10941), .ZN(n24619) );
  AOI22_X1 U4882 ( .A1(\mem[185][7] ), .A2(n10934), .B1(n26945), .B2(
        data_in[7]), .ZN(n10941) );
  INV_X1 U4883 ( .A(n10942), .ZN(n24618) );
  AOI22_X1 U4884 ( .A1(\mem[186][0] ), .A2(n10943), .B1(n26944), .B2(
        data_in[0]), .ZN(n10942) );
  INV_X1 U4885 ( .A(n10944), .ZN(n24617) );
  AOI22_X1 U4886 ( .A1(\mem[186][1] ), .A2(n10943), .B1(n26944), .B2(
        data_in[1]), .ZN(n10944) );
  INV_X1 U4887 ( .A(n10945), .ZN(n24616) );
  AOI22_X1 U4888 ( .A1(\mem[186][2] ), .A2(n10943), .B1(n26944), .B2(
        data_in[2]), .ZN(n10945) );
  INV_X1 U4889 ( .A(n10946), .ZN(n24615) );
  AOI22_X1 U4890 ( .A1(\mem[186][3] ), .A2(n10943), .B1(n26944), .B2(
        data_in[3]), .ZN(n10946) );
  INV_X1 U4891 ( .A(n10947), .ZN(n24614) );
  AOI22_X1 U4892 ( .A1(\mem[186][4] ), .A2(n10943), .B1(n26944), .B2(
        data_in[4]), .ZN(n10947) );
  INV_X1 U4893 ( .A(n10948), .ZN(n24613) );
  AOI22_X1 U4894 ( .A1(\mem[186][5] ), .A2(n10943), .B1(n26944), .B2(
        data_in[5]), .ZN(n10948) );
  INV_X1 U4895 ( .A(n10949), .ZN(n24612) );
  AOI22_X1 U4896 ( .A1(\mem[186][6] ), .A2(n10943), .B1(n26944), .B2(
        data_in[6]), .ZN(n10949) );
  INV_X1 U4897 ( .A(n10950), .ZN(n24611) );
  AOI22_X1 U4898 ( .A1(\mem[186][7] ), .A2(n10943), .B1(n26944), .B2(
        data_in[7]), .ZN(n10950) );
  INV_X1 U4899 ( .A(n10951), .ZN(n24610) );
  AOI22_X1 U4900 ( .A1(\mem[187][0] ), .A2(n10952), .B1(n26943), .B2(
        data_in[0]), .ZN(n10951) );
  INV_X1 U4901 ( .A(n10953), .ZN(n24609) );
  AOI22_X1 U4902 ( .A1(\mem[187][1] ), .A2(n10952), .B1(n26943), .B2(
        data_in[1]), .ZN(n10953) );
  INV_X1 U4903 ( .A(n10954), .ZN(n24608) );
  AOI22_X1 U4904 ( .A1(\mem[187][2] ), .A2(n10952), .B1(n26943), .B2(
        data_in[2]), .ZN(n10954) );
  INV_X1 U4905 ( .A(n10955), .ZN(n24607) );
  AOI22_X1 U4906 ( .A1(\mem[187][3] ), .A2(n10952), .B1(n26943), .B2(
        data_in[3]), .ZN(n10955) );
  INV_X1 U4907 ( .A(n10956), .ZN(n24606) );
  AOI22_X1 U4908 ( .A1(\mem[187][4] ), .A2(n10952), .B1(n26943), .B2(
        data_in[4]), .ZN(n10956) );
  INV_X1 U4909 ( .A(n10957), .ZN(n24605) );
  AOI22_X1 U4910 ( .A1(\mem[187][5] ), .A2(n10952), .B1(n26943), .B2(
        data_in[5]), .ZN(n10957) );
  INV_X1 U4911 ( .A(n10958), .ZN(n24604) );
  AOI22_X1 U4912 ( .A1(\mem[187][6] ), .A2(n10952), .B1(n26943), .B2(
        data_in[6]), .ZN(n10958) );
  INV_X1 U4913 ( .A(n10959), .ZN(n24603) );
  AOI22_X1 U4914 ( .A1(\mem[187][7] ), .A2(n10952), .B1(n26943), .B2(
        data_in[7]), .ZN(n10959) );
  INV_X1 U4915 ( .A(n10960), .ZN(n24602) );
  AOI22_X1 U4916 ( .A1(\mem[188][0] ), .A2(n10961), .B1(n26942), .B2(
        data_in[0]), .ZN(n10960) );
  INV_X1 U4917 ( .A(n10962), .ZN(n24601) );
  AOI22_X1 U4918 ( .A1(\mem[188][1] ), .A2(n10961), .B1(n26942), .B2(
        data_in[1]), .ZN(n10962) );
  INV_X1 U4919 ( .A(n10963), .ZN(n24600) );
  AOI22_X1 U4920 ( .A1(\mem[188][2] ), .A2(n10961), .B1(n26942), .B2(
        data_in[2]), .ZN(n10963) );
  INV_X1 U4921 ( .A(n10964), .ZN(n24599) );
  AOI22_X1 U4922 ( .A1(\mem[188][3] ), .A2(n10961), .B1(n26942), .B2(
        data_in[3]), .ZN(n10964) );
  INV_X1 U4923 ( .A(n10965), .ZN(n24598) );
  AOI22_X1 U4924 ( .A1(\mem[188][4] ), .A2(n10961), .B1(n26942), .B2(
        data_in[4]), .ZN(n10965) );
  INV_X1 U4925 ( .A(n10966), .ZN(n24597) );
  AOI22_X1 U4926 ( .A1(\mem[188][5] ), .A2(n10961), .B1(n26942), .B2(
        data_in[5]), .ZN(n10966) );
  INV_X1 U4927 ( .A(n10967), .ZN(n24596) );
  AOI22_X1 U4928 ( .A1(\mem[188][6] ), .A2(n10961), .B1(n26942), .B2(
        data_in[6]), .ZN(n10967) );
  INV_X1 U4929 ( .A(n10968), .ZN(n24595) );
  AOI22_X1 U4930 ( .A1(\mem[188][7] ), .A2(n10961), .B1(n26942), .B2(
        data_in[7]), .ZN(n10968) );
  INV_X1 U4931 ( .A(n10969), .ZN(n24594) );
  AOI22_X1 U4932 ( .A1(\mem[189][0] ), .A2(n10970), .B1(n26941), .B2(
        data_in[0]), .ZN(n10969) );
  INV_X1 U4933 ( .A(n10971), .ZN(n24593) );
  AOI22_X1 U4934 ( .A1(\mem[189][1] ), .A2(n10970), .B1(n26941), .B2(
        data_in[1]), .ZN(n10971) );
  INV_X1 U4935 ( .A(n10972), .ZN(n24592) );
  AOI22_X1 U4936 ( .A1(\mem[189][2] ), .A2(n10970), .B1(n26941), .B2(
        data_in[2]), .ZN(n10972) );
  INV_X1 U4937 ( .A(n10973), .ZN(n24591) );
  AOI22_X1 U4938 ( .A1(\mem[189][3] ), .A2(n10970), .B1(n26941), .B2(
        data_in[3]), .ZN(n10973) );
  INV_X1 U4939 ( .A(n10974), .ZN(n24590) );
  AOI22_X1 U4940 ( .A1(\mem[189][4] ), .A2(n10970), .B1(n26941), .B2(
        data_in[4]), .ZN(n10974) );
  INV_X1 U4941 ( .A(n10975), .ZN(n24589) );
  AOI22_X1 U4942 ( .A1(\mem[189][5] ), .A2(n10970), .B1(n26941), .B2(
        data_in[5]), .ZN(n10975) );
  INV_X1 U4943 ( .A(n10976), .ZN(n24588) );
  AOI22_X1 U4944 ( .A1(\mem[189][6] ), .A2(n10970), .B1(n26941), .B2(
        data_in[6]), .ZN(n10976) );
  INV_X1 U4945 ( .A(n10977), .ZN(n24587) );
  AOI22_X1 U4946 ( .A1(\mem[189][7] ), .A2(n10970), .B1(n26941), .B2(
        data_in[7]), .ZN(n10977) );
  INV_X1 U4947 ( .A(n10978), .ZN(n24586) );
  AOI22_X1 U4948 ( .A1(\mem[190][0] ), .A2(n10979), .B1(n26940), .B2(
        data_in[0]), .ZN(n10978) );
  INV_X1 U4949 ( .A(n10980), .ZN(n24585) );
  AOI22_X1 U4950 ( .A1(\mem[190][1] ), .A2(n10979), .B1(n26940), .B2(
        data_in[1]), .ZN(n10980) );
  INV_X1 U4951 ( .A(n10981), .ZN(n24584) );
  AOI22_X1 U4952 ( .A1(\mem[190][2] ), .A2(n10979), .B1(n26940), .B2(
        data_in[2]), .ZN(n10981) );
  INV_X1 U4953 ( .A(n10982), .ZN(n24583) );
  AOI22_X1 U4954 ( .A1(\mem[190][3] ), .A2(n10979), .B1(n26940), .B2(
        data_in[3]), .ZN(n10982) );
  INV_X1 U4955 ( .A(n10983), .ZN(n24582) );
  AOI22_X1 U4956 ( .A1(\mem[190][4] ), .A2(n10979), .B1(n26940), .B2(
        data_in[4]), .ZN(n10983) );
  INV_X1 U4957 ( .A(n10984), .ZN(n24581) );
  AOI22_X1 U4958 ( .A1(\mem[190][5] ), .A2(n10979), .B1(n26940), .B2(
        data_in[5]), .ZN(n10984) );
  INV_X1 U4959 ( .A(n10985), .ZN(n24580) );
  AOI22_X1 U4960 ( .A1(\mem[190][6] ), .A2(n10979), .B1(n26940), .B2(
        data_in[6]), .ZN(n10985) );
  INV_X1 U4961 ( .A(n10986), .ZN(n24579) );
  AOI22_X1 U4962 ( .A1(\mem[190][7] ), .A2(n10979), .B1(n26940), .B2(
        data_in[7]), .ZN(n10986) );
  INV_X1 U4963 ( .A(n10987), .ZN(n24578) );
  AOI22_X1 U4964 ( .A1(\mem[191][0] ), .A2(n10988), .B1(n26939), .B2(
        data_in[0]), .ZN(n10987) );
  INV_X1 U4965 ( .A(n10989), .ZN(n24577) );
  AOI22_X1 U4966 ( .A1(\mem[191][1] ), .A2(n10988), .B1(n26939), .B2(
        data_in[1]), .ZN(n10989) );
  INV_X1 U4967 ( .A(n10990), .ZN(n24576) );
  AOI22_X1 U4968 ( .A1(\mem[191][2] ), .A2(n10988), .B1(n26939), .B2(
        data_in[2]), .ZN(n10990) );
  INV_X1 U4969 ( .A(n10991), .ZN(n24575) );
  AOI22_X1 U4970 ( .A1(\mem[191][3] ), .A2(n10988), .B1(n26939), .B2(
        data_in[3]), .ZN(n10991) );
  INV_X1 U4971 ( .A(n10992), .ZN(n24574) );
  AOI22_X1 U4972 ( .A1(\mem[191][4] ), .A2(n10988), .B1(n26939), .B2(
        data_in[4]), .ZN(n10992) );
  INV_X1 U4973 ( .A(n10993), .ZN(n24573) );
  AOI22_X1 U4974 ( .A1(\mem[191][5] ), .A2(n10988), .B1(n26939), .B2(
        data_in[5]), .ZN(n10993) );
  INV_X1 U4975 ( .A(n10994), .ZN(n24572) );
  AOI22_X1 U4976 ( .A1(\mem[191][6] ), .A2(n10988), .B1(n26939), .B2(
        data_in[6]), .ZN(n10994) );
  INV_X1 U4977 ( .A(n10995), .ZN(n24571) );
  AOI22_X1 U4978 ( .A1(\mem[191][7] ), .A2(n10988), .B1(n26939), .B2(
        data_in[7]), .ZN(n10995) );
  INV_X1 U4979 ( .A(n11070), .ZN(n24506) );
  AOI22_X1 U4980 ( .A1(\mem[200][0] ), .A2(n11071), .B1(n26930), .B2(
        data_in[0]), .ZN(n11070) );
  INV_X1 U4981 ( .A(n11072), .ZN(n24505) );
  AOI22_X1 U4982 ( .A1(\mem[200][1] ), .A2(n11071), .B1(n26930), .B2(
        data_in[1]), .ZN(n11072) );
  INV_X1 U4983 ( .A(n11073), .ZN(n24504) );
  AOI22_X1 U4984 ( .A1(\mem[200][2] ), .A2(n11071), .B1(n26930), .B2(
        data_in[2]), .ZN(n11073) );
  INV_X1 U4985 ( .A(n11074), .ZN(n24503) );
  AOI22_X1 U4986 ( .A1(\mem[200][3] ), .A2(n11071), .B1(n26930), .B2(
        data_in[3]), .ZN(n11074) );
  INV_X1 U4987 ( .A(n11075), .ZN(n24502) );
  AOI22_X1 U4988 ( .A1(\mem[200][4] ), .A2(n11071), .B1(n26930), .B2(
        data_in[4]), .ZN(n11075) );
  INV_X1 U4989 ( .A(n11076), .ZN(n24501) );
  AOI22_X1 U4990 ( .A1(\mem[200][5] ), .A2(n11071), .B1(n26930), .B2(
        data_in[5]), .ZN(n11076) );
  INV_X1 U4991 ( .A(n11077), .ZN(n24500) );
  AOI22_X1 U4992 ( .A1(\mem[200][6] ), .A2(n11071), .B1(n26930), .B2(
        data_in[6]), .ZN(n11077) );
  INV_X1 U4993 ( .A(n11078), .ZN(n24499) );
  AOI22_X1 U4994 ( .A1(\mem[200][7] ), .A2(n11071), .B1(n26930), .B2(
        data_in[7]), .ZN(n11078) );
  INV_X1 U4995 ( .A(n11079), .ZN(n24498) );
  AOI22_X1 U4996 ( .A1(\mem[201][0] ), .A2(n11080), .B1(n26929), .B2(
        data_in[0]), .ZN(n11079) );
  INV_X1 U4997 ( .A(n11081), .ZN(n24497) );
  AOI22_X1 U4998 ( .A1(\mem[201][1] ), .A2(n11080), .B1(n26929), .B2(
        data_in[1]), .ZN(n11081) );
  INV_X1 U4999 ( .A(n11082), .ZN(n24496) );
  AOI22_X1 U5000 ( .A1(\mem[201][2] ), .A2(n11080), .B1(n26929), .B2(
        data_in[2]), .ZN(n11082) );
  INV_X1 U5001 ( .A(n11083), .ZN(n24495) );
  AOI22_X1 U5002 ( .A1(\mem[201][3] ), .A2(n11080), .B1(n26929), .B2(
        data_in[3]), .ZN(n11083) );
  INV_X1 U5003 ( .A(n11084), .ZN(n24494) );
  AOI22_X1 U5004 ( .A1(\mem[201][4] ), .A2(n11080), .B1(n26929), .B2(
        data_in[4]), .ZN(n11084) );
  INV_X1 U5005 ( .A(n11085), .ZN(n24493) );
  AOI22_X1 U5006 ( .A1(\mem[201][5] ), .A2(n11080), .B1(n26929), .B2(
        data_in[5]), .ZN(n11085) );
  INV_X1 U5007 ( .A(n11086), .ZN(n24492) );
  AOI22_X1 U5008 ( .A1(\mem[201][6] ), .A2(n11080), .B1(n26929), .B2(
        data_in[6]), .ZN(n11086) );
  INV_X1 U5009 ( .A(n11087), .ZN(n24491) );
  AOI22_X1 U5010 ( .A1(\mem[201][7] ), .A2(n11080), .B1(n26929), .B2(
        data_in[7]), .ZN(n11087) );
  INV_X1 U5011 ( .A(n11088), .ZN(n24490) );
  AOI22_X1 U5012 ( .A1(\mem[202][0] ), .A2(n11089), .B1(n26928), .B2(
        data_in[0]), .ZN(n11088) );
  INV_X1 U5013 ( .A(n11090), .ZN(n24489) );
  AOI22_X1 U5014 ( .A1(\mem[202][1] ), .A2(n11089), .B1(n26928), .B2(
        data_in[1]), .ZN(n11090) );
  INV_X1 U5015 ( .A(n11091), .ZN(n24488) );
  AOI22_X1 U5016 ( .A1(\mem[202][2] ), .A2(n11089), .B1(n26928), .B2(
        data_in[2]), .ZN(n11091) );
  INV_X1 U5017 ( .A(n11092), .ZN(n24487) );
  AOI22_X1 U5018 ( .A1(\mem[202][3] ), .A2(n11089), .B1(n26928), .B2(
        data_in[3]), .ZN(n11092) );
  INV_X1 U5019 ( .A(n11093), .ZN(n24486) );
  AOI22_X1 U5020 ( .A1(\mem[202][4] ), .A2(n11089), .B1(n26928), .B2(
        data_in[4]), .ZN(n11093) );
  INV_X1 U5021 ( .A(n11094), .ZN(n24485) );
  AOI22_X1 U5022 ( .A1(\mem[202][5] ), .A2(n11089), .B1(n26928), .B2(
        data_in[5]), .ZN(n11094) );
  INV_X1 U5023 ( .A(n11095), .ZN(n24484) );
  AOI22_X1 U5024 ( .A1(\mem[202][6] ), .A2(n11089), .B1(n26928), .B2(
        data_in[6]), .ZN(n11095) );
  INV_X1 U5025 ( .A(n11096), .ZN(n24483) );
  AOI22_X1 U5026 ( .A1(\mem[202][7] ), .A2(n11089), .B1(n26928), .B2(
        data_in[7]), .ZN(n11096) );
  INV_X1 U5027 ( .A(n11097), .ZN(n24482) );
  AOI22_X1 U5028 ( .A1(\mem[203][0] ), .A2(n11098), .B1(n26927), .B2(
        data_in[0]), .ZN(n11097) );
  INV_X1 U5029 ( .A(n11099), .ZN(n24481) );
  AOI22_X1 U5030 ( .A1(\mem[203][1] ), .A2(n11098), .B1(n26927), .B2(
        data_in[1]), .ZN(n11099) );
  INV_X1 U5031 ( .A(n11100), .ZN(n24480) );
  AOI22_X1 U5032 ( .A1(\mem[203][2] ), .A2(n11098), .B1(n26927), .B2(
        data_in[2]), .ZN(n11100) );
  INV_X1 U5033 ( .A(n11101), .ZN(n24479) );
  AOI22_X1 U5034 ( .A1(\mem[203][3] ), .A2(n11098), .B1(n26927), .B2(
        data_in[3]), .ZN(n11101) );
  INV_X1 U5035 ( .A(n11102), .ZN(n24478) );
  AOI22_X1 U5036 ( .A1(\mem[203][4] ), .A2(n11098), .B1(n26927), .B2(
        data_in[4]), .ZN(n11102) );
  INV_X1 U5037 ( .A(n11103), .ZN(n24477) );
  AOI22_X1 U5038 ( .A1(\mem[203][5] ), .A2(n11098), .B1(n26927), .B2(
        data_in[5]), .ZN(n11103) );
  INV_X1 U5039 ( .A(n11104), .ZN(n24476) );
  AOI22_X1 U5040 ( .A1(\mem[203][6] ), .A2(n11098), .B1(n26927), .B2(
        data_in[6]), .ZN(n11104) );
  INV_X1 U5041 ( .A(n11105), .ZN(n24475) );
  AOI22_X1 U5042 ( .A1(\mem[203][7] ), .A2(n11098), .B1(n26927), .B2(
        data_in[7]), .ZN(n11105) );
  INV_X1 U5043 ( .A(n11106), .ZN(n24474) );
  AOI22_X1 U5044 ( .A1(\mem[204][0] ), .A2(n11107), .B1(n26926), .B2(
        data_in[0]), .ZN(n11106) );
  INV_X1 U5045 ( .A(n11108), .ZN(n24473) );
  AOI22_X1 U5046 ( .A1(\mem[204][1] ), .A2(n11107), .B1(n26926), .B2(
        data_in[1]), .ZN(n11108) );
  INV_X1 U5047 ( .A(n11109), .ZN(n24472) );
  AOI22_X1 U5048 ( .A1(\mem[204][2] ), .A2(n11107), .B1(n26926), .B2(
        data_in[2]), .ZN(n11109) );
  INV_X1 U5049 ( .A(n11110), .ZN(n24471) );
  AOI22_X1 U5050 ( .A1(\mem[204][3] ), .A2(n11107), .B1(n26926), .B2(
        data_in[3]), .ZN(n11110) );
  INV_X1 U5051 ( .A(n11111), .ZN(n24470) );
  AOI22_X1 U5052 ( .A1(\mem[204][4] ), .A2(n11107), .B1(n26926), .B2(
        data_in[4]), .ZN(n11111) );
  INV_X1 U5053 ( .A(n11112), .ZN(n24469) );
  AOI22_X1 U5054 ( .A1(\mem[204][5] ), .A2(n11107), .B1(n26926), .B2(
        data_in[5]), .ZN(n11112) );
  INV_X1 U5055 ( .A(n11113), .ZN(n24468) );
  AOI22_X1 U5056 ( .A1(\mem[204][6] ), .A2(n11107), .B1(n26926), .B2(
        data_in[6]), .ZN(n11113) );
  INV_X1 U5057 ( .A(n11114), .ZN(n24467) );
  AOI22_X1 U5058 ( .A1(\mem[204][7] ), .A2(n11107), .B1(n26926), .B2(
        data_in[7]), .ZN(n11114) );
  INV_X1 U5059 ( .A(n11115), .ZN(n24466) );
  AOI22_X1 U5060 ( .A1(\mem[205][0] ), .A2(n11116), .B1(n26925), .B2(
        data_in[0]), .ZN(n11115) );
  INV_X1 U5061 ( .A(n11117), .ZN(n24465) );
  AOI22_X1 U5062 ( .A1(\mem[205][1] ), .A2(n11116), .B1(n26925), .B2(
        data_in[1]), .ZN(n11117) );
  INV_X1 U5063 ( .A(n11118), .ZN(n24464) );
  AOI22_X1 U5064 ( .A1(\mem[205][2] ), .A2(n11116), .B1(n26925), .B2(
        data_in[2]), .ZN(n11118) );
  INV_X1 U5065 ( .A(n11119), .ZN(n24463) );
  AOI22_X1 U5066 ( .A1(\mem[205][3] ), .A2(n11116), .B1(n26925), .B2(
        data_in[3]), .ZN(n11119) );
  INV_X1 U5067 ( .A(n11120), .ZN(n24462) );
  AOI22_X1 U5068 ( .A1(\mem[205][4] ), .A2(n11116), .B1(n26925), .B2(
        data_in[4]), .ZN(n11120) );
  INV_X1 U5069 ( .A(n11121), .ZN(n24461) );
  AOI22_X1 U5070 ( .A1(\mem[205][5] ), .A2(n11116), .B1(n26925), .B2(
        data_in[5]), .ZN(n11121) );
  INV_X1 U5071 ( .A(n11122), .ZN(n24460) );
  AOI22_X1 U5072 ( .A1(\mem[205][6] ), .A2(n11116), .B1(n26925), .B2(
        data_in[6]), .ZN(n11122) );
  INV_X1 U5073 ( .A(n11123), .ZN(n24459) );
  AOI22_X1 U5074 ( .A1(\mem[205][7] ), .A2(n11116), .B1(n26925), .B2(
        data_in[7]), .ZN(n11123) );
  INV_X1 U5075 ( .A(n11124), .ZN(n24458) );
  AOI22_X1 U5076 ( .A1(\mem[206][0] ), .A2(n11125), .B1(n26924), .B2(
        data_in[0]), .ZN(n11124) );
  INV_X1 U5077 ( .A(n11126), .ZN(n24457) );
  AOI22_X1 U5078 ( .A1(\mem[206][1] ), .A2(n11125), .B1(n26924), .B2(
        data_in[1]), .ZN(n11126) );
  INV_X1 U5079 ( .A(n11127), .ZN(n24456) );
  AOI22_X1 U5080 ( .A1(\mem[206][2] ), .A2(n11125), .B1(n26924), .B2(
        data_in[2]), .ZN(n11127) );
  INV_X1 U5081 ( .A(n11128), .ZN(n24455) );
  AOI22_X1 U5082 ( .A1(\mem[206][3] ), .A2(n11125), .B1(n26924), .B2(
        data_in[3]), .ZN(n11128) );
  INV_X1 U5083 ( .A(n11129), .ZN(n24454) );
  AOI22_X1 U5084 ( .A1(\mem[206][4] ), .A2(n11125), .B1(n26924), .B2(
        data_in[4]), .ZN(n11129) );
  INV_X1 U5085 ( .A(n11130), .ZN(n24453) );
  AOI22_X1 U5086 ( .A1(\mem[206][5] ), .A2(n11125), .B1(n26924), .B2(
        data_in[5]), .ZN(n11130) );
  INV_X1 U5087 ( .A(n11131), .ZN(n24452) );
  AOI22_X1 U5088 ( .A1(\mem[206][6] ), .A2(n11125), .B1(n26924), .B2(
        data_in[6]), .ZN(n11131) );
  INV_X1 U5089 ( .A(n11132), .ZN(n24451) );
  AOI22_X1 U5090 ( .A1(\mem[206][7] ), .A2(n11125), .B1(n26924), .B2(
        data_in[7]), .ZN(n11132) );
  INV_X1 U5091 ( .A(n11133), .ZN(n24450) );
  AOI22_X1 U5092 ( .A1(\mem[207][0] ), .A2(n11134), .B1(n26923), .B2(
        data_in[0]), .ZN(n11133) );
  INV_X1 U5093 ( .A(n11135), .ZN(n24449) );
  AOI22_X1 U5094 ( .A1(\mem[207][1] ), .A2(n11134), .B1(n26923), .B2(
        data_in[1]), .ZN(n11135) );
  INV_X1 U5095 ( .A(n11136), .ZN(n24448) );
  AOI22_X1 U5096 ( .A1(\mem[207][2] ), .A2(n11134), .B1(n26923), .B2(
        data_in[2]), .ZN(n11136) );
  INV_X1 U5097 ( .A(n11137), .ZN(n24447) );
  AOI22_X1 U5098 ( .A1(\mem[207][3] ), .A2(n11134), .B1(n26923), .B2(
        data_in[3]), .ZN(n11137) );
  INV_X1 U5099 ( .A(n11138), .ZN(n24446) );
  AOI22_X1 U5100 ( .A1(\mem[207][4] ), .A2(n11134), .B1(n26923), .B2(
        data_in[4]), .ZN(n11138) );
  INV_X1 U5101 ( .A(n11139), .ZN(n24445) );
  AOI22_X1 U5102 ( .A1(\mem[207][5] ), .A2(n11134), .B1(n26923), .B2(
        data_in[5]), .ZN(n11139) );
  INV_X1 U5103 ( .A(n11140), .ZN(n24444) );
  AOI22_X1 U5104 ( .A1(\mem[207][6] ), .A2(n11134), .B1(n26923), .B2(
        data_in[6]), .ZN(n11140) );
  INV_X1 U5105 ( .A(n11141), .ZN(n24443) );
  AOI22_X1 U5106 ( .A1(\mem[207][7] ), .A2(n11134), .B1(n26923), .B2(
        data_in[7]), .ZN(n11141) );
  INV_X1 U5107 ( .A(n11142), .ZN(n24442) );
  AOI22_X1 U5108 ( .A1(\mem[208][0] ), .A2(n11143), .B1(n26922), .B2(
        data_in[0]), .ZN(n11142) );
  INV_X1 U5109 ( .A(n11144), .ZN(n24441) );
  AOI22_X1 U5110 ( .A1(\mem[208][1] ), .A2(n11143), .B1(n26922), .B2(
        data_in[1]), .ZN(n11144) );
  INV_X1 U5111 ( .A(n11145), .ZN(n24440) );
  AOI22_X1 U5112 ( .A1(\mem[208][2] ), .A2(n11143), .B1(n26922), .B2(
        data_in[2]), .ZN(n11145) );
  INV_X1 U5113 ( .A(n11146), .ZN(n24439) );
  AOI22_X1 U5114 ( .A1(\mem[208][3] ), .A2(n11143), .B1(n26922), .B2(
        data_in[3]), .ZN(n11146) );
  INV_X1 U5115 ( .A(n11147), .ZN(n24438) );
  AOI22_X1 U5116 ( .A1(\mem[208][4] ), .A2(n11143), .B1(n26922), .B2(
        data_in[4]), .ZN(n11147) );
  INV_X1 U5117 ( .A(n11148), .ZN(n24437) );
  AOI22_X1 U5118 ( .A1(\mem[208][5] ), .A2(n11143), .B1(n26922), .B2(
        data_in[5]), .ZN(n11148) );
  INV_X1 U5119 ( .A(n11149), .ZN(n24436) );
  AOI22_X1 U5120 ( .A1(\mem[208][6] ), .A2(n11143), .B1(n26922), .B2(
        data_in[6]), .ZN(n11149) );
  INV_X1 U5121 ( .A(n11150), .ZN(n24435) );
  AOI22_X1 U5122 ( .A1(\mem[208][7] ), .A2(n11143), .B1(n26922), .B2(
        data_in[7]), .ZN(n11150) );
  INV_X1 U5123 ( .A(n11151), .ZN(n24434) );
  AOI22_X1 U5124 ( .A1(\mem[209][0] ), .A2(n11152), .B1(n26921), .B2(
        data_in[0]), .ZN(n11151) );
  INV_X1 U5125 ( .A(n11153), .ZN(n24433) );
  AOI22_X1 U5126 ( .A1(\mem[209][1] ), .A2(n11152), .B1(n26921), .B2(
        data_in[1]), .ZN(n11153) );
  INV_X1 U5127 ( .A(n11154), .ZN(n24432) );
  AOI22_X1 U5128 ( .A1(\mem[209][2] ), .A2(n11152), .B1(n26921), .B2(
        data_in[2]), .ZN(n11154) );
  INV_X1 U5129 ( .A(n11155), .ZN(n24431) );
  AOI22_X1 U5130 ( .A1(\mem[209][3] ), .A2(n11152), .B1(n26921), .B2(
        data_in[3]), .ZN(n11155) );
  INV_X1 U5131 ( .A(n11156), .ZN(n24430) );
  AOI22_X1 U5132 ( .A1(\mem[209][4] ), .A2(n11152), .B1(n26921), .B2(
        data_in[4]), .ZN(n11156) );
  INV_X1 U5133 ( .A(n11157), .ZN(n24429) );
  AOI22_X1 U5134 ( .A1(\mem[209][5] ), .A2(n11152), .B1(n26921), .B2(
        data_in[5]), .ZN(n11157) );
  INV_X1 U5135 ( .A(n11158), .ZN(n24428) );
  AOI22_X1 U5136 ( .A1(\mem[209][6] ), .A2(n11152), .B1(n26921), .B2(
        data_in[6]), .ZN(n11158) );
  INV_X1 U5137 ( .A(n11159), .ZN(n24427) );
  AOI22_X1 U5138 ( .A1(\mem[209][7] ), .A2(n11152), .B1(n26921), .B2(
        data_in[7]), .ZN(n11159) );
  INV_X1 U5139 ( .A(n11160), .ZN(n24426) );
  AOI22_X1 U5140 ( .A1(\mem[210][0] ), .A2(n11161), .B1(n26920), .B2(
        data_in[0]), .ZN(n11160) );
  INV_X1 U5141 ( .A(n11162), .ZN(n24425) );
  AOI22_X1 U5142 ( .A1(\mem[210][1] ), .A2(n11161), .B1(n26920), .B2(
        data_in[1]), .ZN(n11162) );
  INV_X1 U5143 ( .A(n11163), .ZN(n24424) );
  AOI22_X1 U5144 ( .A1(\mem[210][2] ), .A2(n11161), .B1(n26920), .B2(
        data_in[2]), .ZN(n11163) );
  INV_X1 U5145 ( .A(n11164), .ZN(n24423) );
  AOI22_X1 U5146 ( .A1(\mem[210][3] ), .A2(n11161), .B1(n26920), .B2(
        data_in[3]), .ZN(n11164) );
  INV_X1 U5147 ( .A(n11165), .ZN(n24422) );
  AOI22_X1 U5148 ( .A1(\mem[210][4] ), .A2(n11161), .B1(n26920), .B2(
        data_in[4]), .ZN(n11165) );
  INV_X1 U5149 ( .A(n11166), .ZN(n24421) );
  AOI22_X1 U5150 ( .A1(\mem[210][5] ), .A2(n11161), .B1(n26920), .B2(
        data_in[5]), .ZN(n11166) );
  INV_X1 U5151 ( .A(n11167), .ZN(n24420) );
  AOI22_X1 U5152 ( .A1(\mem[210][6] ), .A2(n11161), .B1(n26920), .B2(
        data_in[6]), .ZN(n11167) );
  INV_X1 U5153 ( .A(n11168), .ZN(n24419) );
  AOI22_X1 U5154 ( .A1(\mem[210][7] ), .A2(n11161), .B1(n26920), .B2(
        data_in[7]), .ZN(n11168) );
  INV_X1 U5155 ( .A(n11169), .ZN(n24418) );
  AOI22_X1 U5156 ( .A1(\mem[211][0] ), .A2(n11170), .B1(n26919), .B2(
        data_in[0]), .ZN(n11169) );
  INV_X1 U5157 ( .A(n11171), .ZN(n24417) );
  AOI22_X1 U5158 ( .A1(\mem[211][1] ), .A2(n11170), .B1(n26919), .B2(
        data_in[1]), .ZN(n11171) );
  INV_X1 U5159 ( .A(n11172), .ZN(n24416) );
  AOI22_X1 U5160 ( .A1(\mem[211][2] ), .A2(n11170), .B1(n26919), .B2(
        data_in[2]), .ZN(n11172) );
  INV_X1 U5161 ( .A(n11173), .ZN(n24415) );
  AOI22_X1 U5162 ( .A1(\mem[211][3] ), .A2(n11170), .B1(n26919), .B2(
        data_in[3]), .ZN(n11173) );
  INV_X1 U5163 ( .A(n11174), .ZN(n24414) );
  AOI22_X1 U5164 ( .A1(\mem[211][4] ), .A2(n11170), .B1(n26919), .B2(
        data_in[4]), .ZN(n11174) );
  INV_X1 U5165 ( .A(n11175), .ZN(n24413) );
  AOI22_X1 U5166 ( .A1(\mem[211][5] ), .A2(n11170), .B1(n26919), .B2(
        data_in[5]), .ZN(n11175) );
  INV_X1 U5167 ( .A(n11176), .ZN(n24412) );
  AOI22_X1 U5168 ( .A1(\mem[211][6] ), .A2(n11170), .B1(n26919), .B2(
        data_in[6]), .ZN(n11176) );
  INV_X1 U5169 ( .A(n11177), .ZN(n24411) );
  AOI22_X1 U5170 ( .A1(\mem[211][7] ), .A2(n11170), .B1(n26919), .B2(
        data_in[7]), .ZN(n11177) );
  INV_X1 U5171 ( .A(n11178), .ZN(n24410) );
  AOI22_X1 U5172 ( .A1(\mem[212][0] ), .A2(n11179), .B1(n26918), .B2(
        data_in[0]), .ZN(n11178) );
  INV_X1 U5173 ( .A(n11180), .ZN(n24409) );
  AOI22_X1 U5174 ( .A1(\mem[212][1] ), .A2(n11179), .B1(n26918), .B2(
        data_in[1]), .ZN(n11180) );
  INV_X1 U5175 ( .A(n11181), .ZN(n24408) );
  AOI22_X1 U5176 ( .A1(\mem[212][2] ), .A2(n11179), .B1(n26918), .B2(
        data_in[2]), .ZN(n11181) );
  INV_X1 U5177 ( .A(n11182), .ZN(n24407) );
  AOI22_X1 U5178 ( .A1(\mem[212][3] ), .A2(n11179), .B1(n26918), .B2(
        data_in[3]), .ZN(n11182) );
  INV_X1 U5179 ( .A(n11183), .ZN(n24406) );
  AOI22_X1 U5180 ( .A1(\mem[212][4] ), .A2(n11179), .B1(n26918), .B2(
        data_in[4]), .ZN(n11183) );
  INV_X1 U5181 ( .A(n11184), .ZN(n24405) );
  AOI22_X1 U5182 ( .A1(\mem[212][5] ), .A2(n11179), .B1(n26918), .B2(
        data_in[5]), .ZN(n11184) );
  INV_X1 U5183 ( .A(n11185), .ZN(n24404) );
  AOI22_X1 U5184 ( .A1(\mem[212][6] ), .A2(n11179), .B1(n26918), .B2(
        data_in[6]), .ZN(n11185) );
  INV_X1 U5185 ( .A(n11186), .ZN(n24403) );
  AOI22_X1 U5186 ( .A1(\mem[212][7] ), .A2(n11179), .B1(n26918), .B2(
        data_in[7]), .ZN(n11186) );
  INV_X1 U5187 ( .A(n11187), .ZN(n24402) );
  AOI22_X1 U5188 ( .A1(\mem[213][0] ), .A2(n11188), .B1(n26917), .B2(
        data_in[0]), .ZN(n11187) );
  INV_X1 U5189 ( .A(n11189), .ZN(n24401) );
  AOI22_X1 U5190 ( .A1(\mem[213][1] ), .A2(n11188), .B1(n26917), .B2(
        data_in[1]), .ZN(n11189) );
  INV_X1 U5191 ( .A(n11190), .ZN(n24400) );
  AOI22_X1 U5192 ( .A1(\mem[213][2] ), .A2(n11188), .B1(n26917), .B2(
        data_in[2]), .ZN(n11190) );
  INV_X1 U5193 ( .A(n11191), .ZN(n24399) );
  AOI22_X1 U5194 ( .A1(\mem[213][3] ), .A2(n11188), .B1(n26917), .B2(
        data_in[3]), .ZN(n11191) );
  INV_X1 U5195 ( .A(n11192), .ZN(n24398) );
  AOI22_X1 U5196 ( .A1(\mem[213][4] ), .A2(n11188), .B1(n26917), .B2(
        data_in[4]), .ZN(n11192) );
  INV_X1 U5197 ( .A(n11193), .ZN(n24397) );
  AOI22_X1 U5198 ( .A1(\mem[213][5] ), .A2(n11188), .B1(n26917), .B2(
        data_in[5]), .ZN(n11193) );
  INV_X1 U5199 ( .A(n11194), .ZN(n24396) );
  AOI22_X1 U5200 ( .A1(\mem[213][6] ), .A2(n11188), .B1(n26917), .B2(
        data_in[6]), .ZN(n11194) );
  INV_X1 U5201 ( .A(n11195), .ZN(n24395) );
  AOI22_X1 U5202 ( .A1(\mem[213][7] ), .A2(n11188), .B1(n26917), .B2(
        data_in[7]), .ZN(n11195) );
  INV_X1 U5203 ( .A(n11196), .ZN(n24394) );
  AOI22_X1 U5204 ( .A1(\mem[214][0] ), .A2(n11197), .B1(n26916), .B2(
        data_in[0]), .ZN(n11196) );
  INV_X1 U5205 ( .A(n11198), .ZN(n24393) );
  AOI22_X1 U5206 ( .A1(\mem[214][1] ), .A2(n11197), .B1(n26916), .B2(
        data_in[1]), .ZN(n11198) );
  INV_X1 U5207 ( .A(n11199), .ZN(n24392) );
  AOI22_X1 U5208 ( .A1(\mem[214][2] ), .A2(n11197), .B1(n26916), .B2(
        data_in[2]), .ZN(n11199) );
  INV_X1 U5209 ( .A(n11200), .ZN(n24391) );
  AOI22_X1 U5210 ( .A1(\mem[214][3] ), .A2(n11197), .B1(n26916), .B2(
        data_in[3]), .ZN(n11200) );
  INV_X1 U5211 ( .A(n11201), .ZN(n24390) );
  AOI22_X1 U5212 ( .A1(\mem[214][4] ), .A2(n11197), .B1(n26916), .B2(
        data_in[4]), .ZN(n11201) );
  INV_X1 U5213 ( .A(n11202), .ZN(n24389) );
  AOI22_X1 U5214 ( .A1(\mem[214][5] ), .A2(n11197), .B1(n26916), .B2(
        data_in[5]), .ZN(n11202) );
  INV_X1 U5215 ( .A(n11203), .ZN(n24388) );
  AOI22_X1 U5216 ( .A1(\mem[214][6] ), .A2(n11197), .B1(n26916), .B2(
        data_in[6]), .ZN(n11203) );
  INV_X1 U5217 ( .A(n11204), .ZN(n24387) );
  AOI22_X1 U5218 ( .A1(\mem[214][7] ), .A2(n11197), .B1(n26916), .B2(
        data_in[7]), .ZN(n11204) );
  INV_X1 U5219 ( .A(n11205), .ZN(n24386) );
  AOI22_X1 U5220 ( .A1(\mem[215][0] ), .A2(n11206), .B1(n26915), .B2(
        data_in[0]), .ZN(n11205) );
  INV_X1 U5221 ( .A(n11207), .ZN(n24385) );
  AOI22_X1 U5222 ( .A1(\mem[215][1] ), .A2(n11206), .B1(n26915), .B2(
        data_in[1]), .ZN(n11207) );
  INV_X1 U5223 ( .A(n11208), .ZN(n24384) );
  AOI22_X1 U5224 ( .A1(\mem[215][2] ), .A2(n11206), .B1(n26915), .B2(
        data_in[2]), .ZN(n11208) );
  INV_X1 U5225 ( .A(n11209), .ZN(n24383) );
  AOI22_X1 U5226 ( .A1(\mem[215][3] ), .A2(n11206), .B1(n26915), .B2(
        data_in[3]), .ZN(n11209) );
  INV_X1 U5227 ( .A(n11210), .ZN(n24382) );
  AOI22_X1 U5228 ( .A1(\mem[215][4] ), .A2(n11206), .B1(n26915), .B2(
        data_in[4]), .ZN(n11210) );
  INV_X1 U5229 ( .A(n11211), .ZN(n24381) );
  AOI22_X1 U5230 ( .A1(\mem[215][5] ), .A2(n11206), .B1(n26915), .B2(
        data_in[5]), .ZN(n11211) );
  INV_X1 U5231 ( .A(n11212), .ZN(n24380) );
  AOI22_X1 U5232 ( .A1(\mem[215][6] ), .A2(n11206), .B1(n26915), .B2(
        data_in[6]), .ZN(n11212) );
  INV_X1 U5233 ( .A(n11213), .ZN(n24379) );
  AOI22_X1 U5234 ( .A1(\mem[215][7] ), .A2(n11206), .B1(n26915), .B2(
        data_in[7]), .ZN(n11213) );
  INV_X1 U5235 ( .A(n11214), .ZN(n24378) );
  AOI22_X1 U5236 ( .A1(\mem[216][0] ), .A2(n11215), .B1(n26914), .B2(
        data_in[0]), .ZN(n11214) );
  INV_X1 U5237 ( .A(n11216), .ZN(n24377) );
  AOI22_X1 U5238 ( .A1(\mem[216][1] ), .A2(n11215), .B1(n26914), .B2(
        data_in[1]), .ZN(n11216) );
  INV_X1 U5239 ( .A(n11217), .ZN(n24376) );
  AOI22_X1 U5240 ( .A1(\mem[216][2] ), .A2(n11215), .B1(n26914), .B2(
        data_in[2]), .ZN(n11217) );
  INV_X1 U5241 ( .A(n11218), .ZN(n24375) );
  AOI22_X1 U5242 ( .A1(\mem[216][3] ), .A2(n11215), .B1(n26914), .B2(
        data_in[3]), .ZN(n11218) );
  INV_X1 U5243 ( .A(n11219), .ZN(n24374) );
  AOI22_X1 U5244 ( .A1(\mem[216][4] ), .A2(n11215), .B1(n26914), .B2(
        data_in[4]), .ZN(n11219) );
  INV_X1 U5245 ( .A(n11220), .ZN(n24373) );
  AOI22_X1 U5246 ( .A1(\mem[216][5] ), .A2(n11215), .B1(n26914), .B2(
        data_in[5]), .ZN(n11220) );
  INV_X1 U5247 ( .A(n11221), .ZN(n24372) );
  AOI22_X1 U5248 ( .A1(\mem[216][6] ), .A2(n11215), .B1(n26914), .B2(
        data_in[6]), .ZN(n11221) );
  INV_X1 U5249 ( .A(n11222), .ZN(n24371) );
  AOI22_X1 U5250 ( .A1(\mem[216][7] ), .A2(n11215), .B1(n26914), .B2(
        data_in[7]), .ZN(n11222) );
  INV_X1 U5251 ( .A(n11223), .ZN(n24370) );
  AOI22_X1 U5252 ( .A1(\mem[217][0] ), .A2(n11224), .B1(n26913), .B2(
        data_in[0]), .ZN(n11223) );
  INV_X1 U5253 ( .A(n11225), .ZN(n24369) );
  AOI22_X1 U5254 ( .A1(\mem[217][1] ), .A2(n11224), .B1(n26913), .B2(
        data_in[1]), .ZN(n11225) );
  INV_X1 U5255 ( .A(n11226), .ZN(n24368) );
  AOI22_X1 U5256 ( .A1(\mem[217][2] ), .A2(n11224), .B1(n26913), .B2(
        data_in[2]), .ZN(n11226) );
  INV_X1 U5257 ( .A(n11227), .ZN(n24367) );
  AOI22_X1 U5258 ( .A1(\mem[217][3] ), .A2(n11224), .B1(n26913), .B2(
        data_in[3]), .ZN(n11227) );
  INV_X1 U5259 ( .A(n11228), .ZN(n24366) );
  AOI22_X1 U5260 ( .A1(\mem[217][4] ), .A2(n11224), .B1(n26913), .B2(
        data_in[4]), .ZN(n11228) );
  INV_X1 U5261 ( .A(n11229), .ZN(n24365) );
  AOI22_X1 U5262 ( .A1(\mem[217][5] ), .A2(n11224), .B1(n26913), .B2(
        data_in[5]), .ZN(n11229) );
  INV_X1 U5263 ( .A(n11230), .ZN(n24364) );
  AOI22_X1 U5264 ( .A1(\mem[217][6] ), .A2(n11224), .B1(n26913), .B2(
        data_in[6]), .ZN(n11230) );
  INV_X1 U5265 ( .A(n11231), .ZN(n24363) );
  AOI22_X1 U5266 ( .A1(\mem[217][7] ), .A2(n11224), .B1(n26913), .B2(
        data_in[7]), .ZN(n11231) );
  INV_X1 U5267 ( .A(n11232), .ZN(n24362) );
  AOI22_X1 U5268 ( .A1(\mem[218][0] ), .A2(n11233), .B1(n26912), .B2(
        data_in[0]), .ZN(n11232) );
  INV_X1 U5269 ( .A(n11234), .ZN(n24361) );
  AOI22_X1 U5270 ( .A1(\mem[218][1] ), .A2(n11233), .B1(n26912), .B2(
        data_in[1]), .ZN(n11234) );
  INV_X1 U5271 ( .A(n11235), .ZN(n24360) );
  AOI22_X1 U5272 ( .A1(\mem[218][2] ), .A2(n11233), .B1(n26912), .B2(
        data_in[2]), .ZN(n11235) );
  INV_X1 U5273 ( .A(n11236), .ZN(n24359) );
  AOI22_X1 U5274 ( .A1(\mem[218][3] ), .A2(n11233), .B1(n26912), .B2(
        data_in[3]), .ZN(n11236) );
  INV_X1 U5275 ( .A(n11237), .ZN(n24358) );
  AOI22_X1 U5276 ( .A1(\mem[218][4] ), .A2(n11233), .B1(n26912), .B2(
        data_in[4]), .ZN(n11237) );
  INV_X1 U5277 ( .A(n11238), .ZN(n24357) );
  AOI22_X1 U5278 ( .A1(\mem[218][5] ), .A2(n11233), .B1(n26912), .B2(
        data_in[5]), .ZN(n11238) );
  INV_X1 U5279 ( .A(n11239), .ZN(n24356) );
  AOI22_X1 U5280 ( .A1(\mem[218][6] ), .A2(n11233), .B1(n26912), .B2(
        data_in[6]), .ZN(n11239) );
  INV_X1 U5281 ( .A(n11240), .ZN(n24355) );
  AOI22_X1 U5282 ( .A1(\mem[218][7] ), .A2(n11233), .B1(n26912), .B2(
        data_in[7]), .ZN(n11240) );
  INV_X1 U5283 ( .A(n11241), .ZN(n24354) );
  AOI22_X1 U5284 ( .A1(\mem[219][0] ), .A2(n11242), .B1(n26911), .B2(
        data_in[0]), .ZN(n11241) );
  INV_X1 U5285 ( .A(n11243), .ZN(n24353) );
  AOI22_X1 U5286 ( .A1(\mem[219][1] ), .A2(n11242), .B1(n26911), .B2(
        data_in[1]), .ZN(n11243) );
  INV_X1 U5287 ( .A(n11244), .ZN(n24352) );
  AOI22_X1 U5288 ( .A1(\mem[219][2] ), .A2(n11242), .B1(n26911), .B2(
        data_in[2]), .ZN(n11244) );
  INV_X1 U5289 ( .A(n11245), .ZN(n24351) );
  AOI22_X1 U5290 ( .A1(\mem[219][3] ), .A2(n11242), .B1(n26911), .B2(
        data_in[3]), .ZN(n11245) );
  INV_X1 U5291 ( .A(n11246), .ZN(n24350) );
  AOI22_X1 U5292 ( .A1(\mem[219][4] ), .A2(n11242), .B1(n26911), .B2(
        data_in[4]), .ZN(n11246) );
  INV_X1 U5293 ( .A(n11247), .ZN(n24349) );
  AOI22_X1 U5294 ( .A1(\mem[219][5] ), .A2(n11242), .B1(n26911), .B2(
        data_in[5]), .ZN(n11247) );
  INV_X1 U5295 ( .A(n11248), .ZN(n24348) );
  AOI22_X1 U5296 ( .A1(\mem[219][6] ), .A2(n11242), .B1(n26911), .B2(
        data_in[6]), .ZN(n11248) );
  INV_X1 U5297 ( .A(n11249), .ZN(n24347) );
  AOI22_X1 U5298 ( .A1(\mem[219][7] ), .A2(n11242), .B1(n26911), .B2(
        data_in[7]), .ZN(n11249) );
  INV_X1 U5299 ( .A(n11250), .ZN(n24346) );
  AOI22_X1 U5300 ( .A1(\mem[220][0] ), .A2(n11251), .B1(n26910), .B2(
        data_in[0]), .ZN(n11250) );
  INV_X1 U5301 ( .A(n11252), .ZN(n24345) );
  AOI22_X1 U5302 ( .A1(\mem[220][1] ), .A2(n11251), .B1(n26910), .B2(
        data_in[1]), .ZN(n11252) );
  INV_X1 U5303 ( .A(n11253), .ZN(n24344) );
  AOI22_X1 U5304 ( .A1(\mem[220][2] ), .A2(n11251), .B1(n26910), .B2(
        data_in[2]), .ZN(n11253) );
  INV_X1 U5305 ( .A(n11254), .ZN(n24343) );
  AOI22_X1 U5306 ( .A1(\mem[220][3] ), .A2(n11251), .B1(n26910), .B2(
        data_in[3]), .ZN(n11254) );
  INV_X1 U5307 ( .A(n11255), .ZN(n24342) );
  AOI22_X1 U5308 ( .A1(\mem[220][4] ), .A2(n11251), .B1(n26910), .B2(
        data_in[4]), .ZN(n11255) );
  INV_X1 U5309 ( .A(n11256), .ZN(n24341) );
  AOI22_X1 U5310 ( .A1(\mem[220][5] ), .A2(n11251), .B1(n26910), .B2(
        data_in[5]), .ZN(n11256) );
  INV_X1 U5311 ( .A(n11257), .ZN(n24340) );
  AOI22_X1 U5312 ( .A1(\mem[220][6] ), .A2(n11251), .B1(n26910), .B2(
        data_in[6]), .ZN(n11257) );
  INV_X1 U5313 ( .A(n11258), .ZN(n24339) );
  AOI22_X1 U5314 ( .A1(\mem[220][7] ), .A2(n11251), .B1(n26910), .B2(
        data_in[7]), .ZN(n11258) );
  INV_X1 U5315 ( .A(n11259), .ZN(n24338) );
  AOI22_X1 U5316 ( .A1(\mem[221][0] ), .A2(n11260), .B1(n26909), .B2(
        data_in[0]), .ZN(n11259) );
  INV_X1 U5317 ( .A(n11261), .ZN(n24337) );
  AOI22_X1 U5318 ( .A1(\mem[221][1] ), .A2(n11260), .B1(n26909), .B2(
        data_in[1]), .ZN(n11261) );
  INV_X1 U5319 ( .A(n11262), .ZN(n24336) );
  AOI22_X1 U5320 ( .A1(\mem[221][2] ), .A2(n11260), .B1(n26909), .B2(
        data_in[2]), .ZN(n11262) );
  INV_X1 U5321 ( .A(n11263), .ZN(n24335) );
  AOI22_X1 U5322 ( .A1(\mem[221][3] ), .A2(n11260), .B1(n26909), .B2(
        data_in[3]), .ZN(n11263) );
  INV_X1 U5323 ( .A(n11264), .ZN(n24334) );
  AOI22_X1 U5324 ( .A1(\mem[221][4] ), .A2(n11260), .B1(n26909), .B2(
        data_in[4]), .ZN(n11264) );
  INV_X1 U5325 ( .A(n11265), .ZN(n24333) );
  AOI22_X1 U5326 ( .A1(\mem[221][5] ), .A2(n11260), .B1(n26909), .B2(
        data_in[5]), .ZN(n11265) );
  INV_X1 U5327 ( .A(n11266), .ZN(n24332) );
  AOI22_X1 U5328 ( .A1(\mem[221][6] ), .A2(n11260), .B1(n26909), .B2(
        data_in[6]), .ZN(n11266) );
  INV_X1 U5329 ( .A(n11267), .ZN(n24331) );
  AOI22_X1 U5330 ( .A1(\mem[221][7] ), .A2(n11260), .B1(n26909), .B2(
        data_in[7]), .ZN(n11267) );
  INV_X1 U5331 ( .A(n11268), .ZN(n24330) );
  AOI22_X1 U5332 ( .A1(\mem[222][0] ), .A2(n11269), .B1(n26908), .B2(
        data_in[0]), .ZN(n11268) );
  INV_X1 U5333 ( .A(n11270), .ZN(n24329) );
  AOI22_X1 U5334 ( .A1(\mem[222][1] ), .A2(n11269), .B1(n26908), .B2(
        data_in[1]), .ZN(n11270) );
  INV_X1 U5335 ( .A(n11271), .ZN(n24328) );
  AOI22_X1 U5336 ( .A1(\mem[222][2] ), .A2(n11269), .B1(n26908), .B2(
        data_in[2]), .ZN(n11271) );
  INV_X1 U5337 ( .A(n11272), .ZN(n24327) );
  AOI22_X1 U5338 ( .A1(\mem[222][3] ), .A2(n11269), .B1(n26908), .B2(
        data_in[3]), .ZN(n11272) );
  INV_X1 U5339 ( .A(n11273), .ZN(n24326) );
  AOI22_X1 U5340 ( .A1(\mem[222][4] ), .A2(n11269), .B1(n26908), .B2(
        data_in[4]), .ZN(n11273) );
  INV_X1 U5341 ( .A(n11274), .ZN(n24325) );
  AOI22_X1 U5342 ( .A1(\mem[222][5] ), .A2(n11269), .B1(n26908), .B2(
        data_in[5]), .ZN(n11274) );
  INV_X1 U5343 ( .A(n11275), .ZN(n24324) );
  AOI22_X1 U5344 ( .A1(\mem[222][6] ), .A2(n11269), .B1(n26908), .B2(
        data_in[6]), .ZN(n11275) );
  INV_X1 U5345 ( .A(n11276), .ZN(n24323) );
  AOI22_X1 U5346 ( .A1(\mem[222][7] ), .A2(n11269), .B1(n26908), .B2(
        data_in[7]), .ZN(n11276) );
  INV_X1 U5347 ( .A(n11277), .ZN(n24322) );
  AOI22_X1 U5348 ( .A1(\mem[223][0] ), .A2(n11278), .B1(n26907), .B2(
        data_in[0]), .ZN(n11277) );
  INV_X1 U5349 ( .A(n11279), .ZN(n24321) );
  AOI22_X1 U5350 ( .A1(\mem[223][1] ), .A2(n11278), .B1(n26907), .B2(
        data_in[1]), .ZN(n11279) );
  INV_X1 U5351 ( .A(n11280), .ZN(n24320) );
  AOI22_X1 U5352 ( .A1(\mem[223][2] ), .A2(n11278), .B1(n26907), .B2(
        data_in[2]), .ZN(n11280) );
  INV_X1 U5353 ( .A(n11281), .ZN(n24319) );
  AOI22_X1 U5354 ( .A1(\mem[223][3] ), .A2(n11278), .B1(n26907), .B2(
        data_in[3]), .ZN(n11281) );
  INV_X1 U5355 ( .A(n11282), .ZN(n24318) );
  AOI22_X1 U5356 ( .A1(\mem[223][4] ), .A2(n11278), .B1(n26907), .B2(
        data_in[4]), .ZN(n11282) );
  INV_X1 U5357 ( .A(n11283), .ZN(n24317) );
  AOI22_X1 U5358 ( .A1(\mem[223][5] ), .A2(n11278), .B1(n26907), .B2(
        data_in[5]), .ZN(n11283) );
  INV_X1 U5359 ( .A(n11284), .ZN(n24316) );
  AOI22_X1 U5360 ( .A1(\mem[223][6] ), .A2(n11278), .B1(n26907), .B2(
        data_in[6]), .ZN(n11284) );
  INV_X1 U5361 ( .A(n11285), .ZN(n24315) );
  AOI22_X1 U5362 ( .A1(\mem[223][7] ), .A2(n11278), .B1(n26907), .B2(
        data_in[7]), .ZN(n11285) );
  INV_X1 U5363 ( .A(n11360), .ZN(n24250) );
  AOI22_X1 U5364 ( .A1(\mem[232][0] ), .A2(n11361), .B1(n26898), .B2(
        data_in[0]), .ZN(n11360) );
  INV_X1 U5365 ( .A(n11362), .ZN(n24249) );
  AOI22_X1 U5366 ( .A1(\mem[232][1] ), .A2(n11361), .B1(n26898), .B2(
        data_in[1]), .ZN(n11362) );
  INV_X1 U5367 ( .A(n11363), .ZN(n24248) );
  AOI22_X1 U5368 ( .A1(\mem[232][2] ), .A2(n11361), .B1(n26898), .B2(
        data_in[2]), .ZN(n11363) );
  INV_X1 U5369 ( .A(n11364), .ZN(n24247) );
  AOI22_X1 U5370 ( .A1(\mem[232][3] ), .A2(n11361), .B1(n26898), .B2(
        data_in[3]), .ZN(n11364) );
  INV_X1 U5371 ( .A(n11365), .ZN(n24246) );
  AOI22_X1 U5372 ( .A1(\mem[232][4] ), .A2(n11361), .B1(n26898), .B2(
        data_in[4]), .ZN(n11365) );
  INV_X1 U5373 ( .A(n11366), .ZN(n24245) );
  AOI22_X1 U5374 ( .A1(\mem[232][5] ), .A2(n11361), .B1(n26898), .B2(
        data_in[5]), .ZN(n11366) );
  INV_X1 U5375 ( .A(n11367), .ZN(n24244) );
  AOI22_X1 U5376 ( .A1(\mem[232][6] ), .A2(n11361), .B1(n26898), .B2(
        data_in[6]), .ZN(n11367) );
  INV_X1 U5377 ( .A(n11368), .ZN(n24243) );
  AOI22_X1 U5378 ( .A1(\mem[232][7] ), .A2(n11361), .B1(n26898), .B2(
        data_in[7]), .ZN(n11368) );
  INV_X1 U5379 ( .A(n11369), .ZN(n24242) );
  AOI22_X1 U5380 ( .A1(\mem[233][0] ), .A2(n11370), .B1(n26897), .B2(
        data_in[0]), .ZN(n11369) );
  INV_X1 U5381 ( .A(n11371), .ZN(n24241) );
  AOI22_X1 U5382 ( .A1(\mem[233][1] ), .A2(n11370), .B1(n26897), .B2(
        data_in[1]), .ZN(n11371) );
  INV_X1 U5383 ( .A(n11372), .ZN(n24240) );
  AOI22_X1 U5384 ( .A1(\mem[233][2] ), .A2(n11370), .B1(n26897), .B2(
        data_in[2]), .ZN(n11372) );
  INV_X1 U5385 ( .A(n11373), .ZN(n24239) );
  AOI22_X1 U5386 ( .A1(\mem[233][3] ), .A2(n11370), .B1(n26897), .B2(
        data_in[3]), .ZN(n11373) );
  INV_X1 U5387 ( .A(n11374), .ZN(n24238) );
  AOI22_X1 U5388 ( .A1(\mem[233][4] ), .A2(n11370), .B1(n26897), .B2(
        data_in[4]), .ZN(n11374) );
  INV_X1 U5389 ( .A(n11375), .ZN(n24237) );
  AOI22_X1 U5390 ( .A1(\mem[233][5] ), .A2(n11370), .B1(n26897), .B2(
        data_in[5]), .ZN(n11375) );
  INV_X1 U5391 ( .A(n11376), .ZN(n24236) );
  AOI22_X1 U5392 ( .A1(\mem[233][6] ), .A2(n11370), .B1(n26897), .B2(
        data_in[6]), .ZN(n11376) );
  INV_X1 U5393 ( .A(n11377), .ZN(n24235) );
  AOI22_X1 U5394 ( .A1(\mem[233][7] ), .A2(n11370), .B1(n26897), .B2(
        data_in[7]), .ZN(n11377) );
  INV_X1 U5395 ( .A(n11378), .ZN(n24234) );
  AOI22_X1 U5396 ( .A1(\mem[234][0] ), .A2(n11379), .B1(n26896), .B2(
        data_in[0]), .ZN(n11378) );
  INV_X1 U5397 ( .A(n11380), .ZN(n24233) );
  AOI22_X1 U5398 ( .A1(\mem[234][1] ), .A2(n11379), .B1(n26896), .B2(
        data_in[1]), .ZN(n11380) );
  INV_X1 U5399 ( .A(n11381), .ZN(n24232) );
  AOI22_X1 U5400 ( .A1(\mem[234][2] ), .A2(n11379), .B1(n26896), .B2(
        data_in[2]), .ZN(n11381) );
  INV_X1 U5401 ( .A(n11382), .ZN(n24231) );
  AOI22_X1 U5402 ( .A1(\mem[234][3] ), .A2(n11379), .B1(n26896), .B2(
        data_in[3]), .ZN(n11382) );
  INV_X1 U5403 ( .A(n11383), .ZN(n24230) );
  AOI22_X1 U5404 ( .A1(\mem[234][4] ), .A2(n11379), .B1(n26896), .B2(
        data_in[4]), .ZN(n11383) );
  INV_X1 U5405 ( .A(n11384), .ZN(n24229) );
  AOI22_X1 U5406 ( .A1(\mem[234][5] ), .A2(n11379), .B1(n26896), .B2(
        data_in[5]), .ZN(n11384) );
  INV_X1 U5407 ( .A(n11385), .ZN(n24228) );
  AOI22_X1 U5408 ( .A1(\mem[234][6] ), .A2(n11379), .B1(n26896), .B2(
        data_in[6]), .ZN(n11385) );
  INV_X1 U5409 ( .A(n11386), .ZN(n24227) );
  AOI22_X1 U5410 ( .A1(\mem[234][7] ), .A2(n11379), .B1(n26896), .B2(
        data_in[7]), .ZN(n11386) );
  INV_X1 U5411 ( .A(n11387), .ZN(n24226) );
  AOI22_X1 U5412 ( .A1(\mem[235][0] ), .A2(n11388), .B1(n26895), .B2(
        data_in[0]), .ZN(n11387) );
  INV_X1 U5413 ( .A(n11389), .ZN(n24225) );
  AOI22_X1 U5414 ( .A1(\mem[235][1] ), .A2(n11388), .B1(n26895), .B2(
        data_in[1]), .ZN(n11389) );
  INV_X1 U5415 ( .A(n11390), .ZN(n24224) );
  AOI22_X1 U5416 ( .A1(\mem[235][2] ), .A2(n11388), .B1(n26895), .B2(
        data_in[2]), .ZN(n11390) );
  INV_X1 U5417 ( .A(n11391), .ZN(n24223) );
  AOI22_X1 U5418 ( .A1(\mem[235][3] ), .A2(n11388), .B1(n26895), .B2(
        data_in[3]), .ZN(n11391) );
  INV_X1 U5419 ( .A(n11392), .ZN(n24222) );
  AOI22_X1 U5420 ( .A1(\mem[235][4] ), .A2(n11388), .B1(n26895), .B2(
        data_in[4]), .ZN(n11392) );
  INV_X1 U5421 ( .A(n11393), .ZN(n24221) );
  AOI22_X1 U5422 ( .A1(\mem[235][5] ), .A2(n11388), .B1(n26895), .B2(
        data_in[5]), .ZN(n11393) );
  INV_X1 U5423 ( .A(n11394), .ZN(n24220) );
  AOI22_X1 U5424 ( .A1(\mem[235][6] ), .A2(n11388), .B1(n26895), .B2(
        data_in[6]), .ZN(n11394) );
  INV_X1 U5425 ( .A(n11395), .ZN(n24219) );
  AOI22_X1 U5426 ( .A1(\mem[235][7] ), .A2(n11388), .B1(n26895), .B2(
        data_in[7]), .ZN(n11395) );
  INV_X1 U5427 ( .A(n11396), .ZN(n24218) );
  AOI22_X1 U5428 ( .A1(\mem[236][0] ), .A2(n11397), .B1(n26894), .B2(
        data_in[0]), .ZN(n11396) );
  INV_X1 U5429 ( .A(n11398), .ZN(n24217) );
  AOI22_X1 U5430 ( .A1(\mem[236][1] ), .A2(n11397), .B1(n26894), .B2(
        data_in[1]), .ZN(n11398) );
  INV_X1 U5431 ( .A(n11399), .ZN(n24216) );
  AOI22_X1 U5432 ( .A1(\mem[236][2] ), .A2(n11397), .B1(n26894), .B2(
        data_in[2]), .ZN(n11399) );
  INV_X1 U5433 ( .A(n11400), .ZN(n24215) );
  AOI22_X1 U5434 ( .A1(\mem[236][3] ), .A2(n11397), .B1(n26894), .B2(
        data_in[3]), .ZN(n11400) );
  INV_X1 U5435 ( .A(n11401), .ZN(n24214) );
  AOI22_X1 U5436 ( .A1(\mem[236][4] ), .A2(n11397), .B1(n26894), .B2(
        data_in[4]), .ZN(n11401) );
  INV_X1 U5437 ( .A(n11402), .ZN(n24213) );
  AOI22_X1 U5438 ( .A1(\mem[236][5] ), .A2(n11397), .B1(n26894), .B2(
        data_in[5]), .ZN(n11402) );
  INV_X1 U5439 ( .A(n11403), .ZN(n24212) );
  AOI22_X1 U5440 ( .A1(\mem[236][6] ), .A2(n11397), .B1(n26894), .B2(
        data_in[6]), .ZN(n11403) );
  INV_X1 U5441 ( .A(n11404), .ZN(n24211) );
  AOI22_X1 U5442 ( .A1(\mem[236][7] ), .A2(n11397), .B1(n26894), .B2(
        data_in[7]), .ZN(n11404) );
  INV_X1 U5443 ( .A(n11405), .ZN(n24210) );
  AOI22_X1 U5444 ( .A1(\mem[237][0] ), .A2(n11406), .B1(n26893), .B2(
        data_in[0]), .ZN(n11405) );
  INV_X1 U5445 ( .A(n11407), .ZN(n24209) );
  AOI22_X1 U5446 ( .A1(\mem[237][1] ), .A2(n11406), .B1(n26893), .B2(
        data_in[1]), .ZN(n11407) );
  INV_X1 U5447 ( .A(n11408), .ZN(n24208) );
  AOI22_X1 U5448 ( .A1(\mem[237][2] ), .A2(n11406), .B1(n26893), .B2(
        data_in[2]), .ZN(n11408) );
  INV_X1 U5449 ( .A(n11409), .ZN(n24207) );
  AOI22_X1 U5450 ( .A1(\mem[237][3] ), .A2(n11406), .B1(n26893), .B2(
        data_in[3]), .ZN(n11409) );
  INV_X1 U5451 ( .A(n11410), .ZN(n24206) );
  AOI22_X1 U5452 ( .A1(\mem[237][4] ), .A2(n11406), .B1(n26893), .B2(
        data_in[4]), .ZN(n11410) );
  INV_X1 U5453 ( .A(n11411), .ZN(n24205) );
  AOI22_X1 U5454 ( .A1(\mem[237][5] ), .A2(n11406), .B1(n26893), .B2(
        data_in[5]), .ZN(n11411) );
  INV_X1 U5455 ( .A(n11412), .ZN(n24204) );
  AOI22_X1 U5456 ( .A1(\mem[237][6] ), .A2(n11406), .B1(n26893), .B2(
        data_in[6]), .ZN(n11412) );
  INV_X1 U5457 ( .A(n11413), .ZN(n24203) );
  AOI22_X1 U5458 ( .A1(\mem[237][7] ), .A2(n11406), .B1(n26893), .B2(
        data_in[7]), .ZN(n11413) );
  INV_X1 U5459 ( .A(n11414), .ZN(n24202) );
  AOI22_X1 U5460 ( .A1(\mem[238][0] ), .A2(n11415), .B1(n26892), .B2(
        data_in[0]), .ZN(n11414) );
  INV_X1 U5461 ( .A(n11416), .ZN(n24201) );
  AOI22_X1 U5462 ( .A1(\mem[238][1] ), .A2(n11415), .B1(n26892), .B2(
        data_in[1]), .ZN(n11416) );
  INV_X1 U5463 ( .A(n11417), .ZN(n24200) );
  AOI22_X1 U5464 ( .A1(\mem[238][2] ), .A2(n11415), .B1(n26892), .B2(
        data_in[2]), .ZN(n11417) );
  INV_X1 U5465 ( .A(n11418), .ZN(n24199) );
  AOI22_X1 U5466 ( .A1(\mem[238][3] ), .A2(n11415), .B1(n26892), .B2(
        data_in[3]), .ZN(n11418) );
  INV_X1 U5467 ( .A(n11419), .ZN(n24198) );
  AOI22_X1 U5468 ( .A1(\mem[238][4] ), .A2(n11415), .B1(n26892), .B2(
        data_in[4]), .ZN(n11419) );
  INV_X1 U5469 ( .A(n11420), .ZN(n24197) );
  AOI22_X1 U5470 ( .A1(\mem[238][5] ), .A2(n11415), .B1(n26892), .B2(
        data_in[5]), .ZN(n11420) );
  INV_X1 U5471 ( .A(n11421), .ZN(n24196) );
  AOI22_X1 U5472 ( .A1(\mem[238][6] ), .A2(n11415), .B1(n26892), .B2(
        data_in[6]), .ZN(n11421) );
  INV_X1 U5473 ( .A(n11422), .ZN(n24195) );
  AOI22_X1 U5474 ( .A1(\mem[238][7] ), .A2(n11415), .B1(n26892), .B2(
        data_in[7]), .ZN(n11422) );
  INV_X1 U5475 ( .A(n11423), .ZN(n24194) );
  AOI22_X1 U5476 ( .A1(\mem[239][0] ), .A2(n11424), .B1(n26891), .B2(
        data_in[0]), .ZN(n11423) );
  INV_X1 U5477 ( .A(n11425), .ZN(n24193) );
  AOI22_X1 U5478 ( .A1(\mem[239][1] ), .A2(n11424), .B1(n26891), .B2(
        data_in[1]), .ZN(n11425) );
  INV_X1 U5479 ( .A(n11426), .ZN(n24192) );
  AOI22_X1 U5480 ( .A1(\mem[239][2] ), .A2(n11424), .B1(n26891), .B2(
        data_in[2]), .ZN(n11426) );
  INV_X1 U5481 ( .A(n11427), .ZN(n24191) );
  AOI22_X1 U5482 ( .A1(\mem[239][3] ), .A2(n11424), .B1(n26891), .B2(
        data_in[3]), .ZN(n11427) );
  INV_X1 U5483 ( .A(n11428), .ZN(n24190) );
  AOI22_X1 U5484 ( .A1(\mem[239][4] ), .A2(n11424), .B1(n26891), .B2(
        data_in[4]), .ZN(n11428) );
  INV_X1 U5485 ( .A(n11429), .ZN(n24189) );
  AOI22_X1 U5486 ( .A1(\mem[239][5] ), .A2(n11424), .B1(n26891), .B2(
        data_in[5]), .ZN(n11429) );
  INV_X1 U5487 ( .A(n11430), .ZN(n24188) );
  AOI22_X1 U5488 ( .A1(\mem[239][6] ), .A2(n11424), .B1(n26891), .B2(
        data_in[6]), .ZN(n11430) );
  INV_X1 U5489 ( .A(n11431), .ZN(n24187) );
  AOI22_X1 U5490 ( .A1(\mem[239][7] ), .A2(n11424), .B1(n26891), .B2(
        data_in[7]), .ZN(n11431) );
  INV_X1 U5491 ( .A(n11432), .ZN(n24186) );
  AOI22_X1 U5492 ( .A1(\mem[240][0] ), .A2(n11433), .B1(n26890), .B2(
        data_in[0]), .ZN(n11432) );
  INV_X1 U5493 ( .A(n11434), .ZN(n24185) );
  AOI22_X1 U5494 ( .A1(\mem[240][1] ), .A2(n11433), .B1(n26890), .B2(
        data_in[1]), .ZN(n11434) );
  INV_X1 U5495 ( .A(n11435), .ZN(n24184) );
  AOI22_X1 U5496 ( .A1(\mem[240][2] ), .A2(n11433), .B1(n26890), .B2(
        data_in[2]), .ZN(n11435) );
  INV_X1 U5497 ( .A(n11436), .ZN(n24183) );
  AOI22_X1 U5498 ( .A1(\mem[240][3] ), .A2(n11433), .B1(n26890), .B2(
        data_in[3]), .ZN(n11436) );
  INV_X1 U5499 ( .A(n11437), .ZN(n24182) );
  AOI22_X1 U5500 ( .A1(\mem[240][4] ), .A2(n11433), .B1(n26890), .B2(
        data_in[4]), .ZN(n11437) );
  INV_X1 U5501 ( .A(n11438), .ZN(n24181) );
  AOI22_X1 U5502 ( .A1(\mem[240][5] ), .A2(n11433), .B1(n26890), .B2(
        data_in[5]), .ZN(n11438) );
  INV_X1 U5503 ( .A(n11439), .ZN(n24180) );
  AOI22_X1 U5504 ( .A1(\mem[240][6] ), .A2(n11433), .B1(n26890), .B2(
        data_in[6]), .ZN(n11439) );
  INV_X1 U5505 ( .A(n11440), .ZN(n24179) );
  AOI22_X1 U5506 ( .A1(\mem[240][7] ), .A2(n11433), .B1(n26890), .B2(
        data_in[7]), .ZN(n11440) );
  INV_X1 U5507 ( .A(n11441), .ZN(n24178) );
  AOI22_X1 U5508 ( .A1(\mem[241][0] ), .A2(n11442), .B1(n26889), .B2(
        data_in[0]), .ZN(n11441) );
  INV_X1 U5509 ( .A(n11443), .ZN(n24177) );
  AOI22_X1 U5510 ( .A1(\mem[241][1] ), .A2(n11442), .B1(n26889), .B2(
        data_in[1]), .ZN(n11443) );
  INV_X1 U5511 ( .A(n11444), .ZN(n24176) );
  AOI22_X1 U5512 ( .A1(\mem[241][2] ), .A2(n11442), .B1(n26889), .B2(
        data_in[2]), .ZN(n11444) );
  INV_X1 U5513 ( .A(n11445), .ZN(n24175) );
  AOI22_X1 U5514 ( .A1(\mem[241][3] ), .A2(n11442), .B1(n26889), .B2(
        data_in[3]), .ZN(n11445) );
  INV_X1 U5515 ( .A(n11446), .ZN(n24174) );
  AOI22_X1 U5516 ( .A1(\mem[241][4] ), .A2(n11442), .B1(n26889), .B2(
        data_in[4]), .ZN(n11446) );
  INV_X1 U5517 ( .A(n11447), .ZN(n24173) );
  AOI22_X1 U5518 ( .A1(\mem[241][5] ), .A2(n11442), .B1(n26889), .B2(
        data_in[5]), .ZN(n11447) );
  INV_X1 U5519 ( .A(n11448), .ZN(n24172) );
  AOI22_X1 U5520 ( .A1(\mem[241][6] ), .A2(n11442), .B1(n26889), .B2(
        data_in[6]), .ZN(n11448) );
  INV_X1 U5521 ( .A(n11449), .ZN(n24171) );
  AOI22_X1 U5522 ( .A1(\mem[241][7] ), .A2(n11442), .B1(n26889), .B2(
        data_in[7]), .ZN(n11449) );
  INV_X1 U5523 ( .A(n11450), .ZN(n24170) );
  AOI22_X1 U5524 ( .A1(\mem[242][0] ), .A2(n11451), .B1(n26888), .B2(
        data_in[0]), .ZN(n11450) );
  INV_X1 U5525 ( .A(n11452), .ZN(n24169) );
  AOI22_X1 U5526 ( .A1(\mem[242][1] ), .A2(n11451), .B1(n26888), .B2(
        data_in[1]), .ZN(n11452) );
  INV_X1 U5527 ( .A(n11453), .ZN(n24168) );
  AOI22_X1 U5528 ( .A1(\mem[242][2] ), .A2(n11451), .B1(n26888), .B2(
        data_in[2]), .ZN(n11453) );
  INV_X1 U5529 ( .A(n11454), .ZN(n24167) );
  AOI22_X1 U5530 ( .A1(\mem[242][3] ), .A2(n11451), .B1(n26888), .B2(
        data_in[3]), .ZN(n11454) );
  INV_X1 U5531 ( .A(n11455), .ZN(n24166) );
  AOI22_X1 U5532 ( .A1(\mem[242][4] ), .A2(n11451), .B1(n26888), .B2(
        data_in[4]), .ZN(n11455) );
  INV_X1 U5533 ( .A(n11456), .ZN(n24165) );
  AOI22_X1 U5534 ( .A1(\mem[242][5] ), .A2(n11451), .B1(n26888), .B2(
        data_in[5]), .ZN(n11456) );
  INV_X1 U5535 ( .A(n11457), .ZN(n24164) );
  AOI22_X1 U5536 ( .A1(\mem[242][6] ), .A2(n11451), .B1(n26888), .B2(
        data_in[6]), .ZN(n11457) );
  INV_X1 U5537 ( .A(n11458), .ZN(n24163) );
  AOI22_X1 U5538 ( .A1(\mem[242][7] ), .A2(n11451), .B1(n26888), .B2(
        data_in[7]), .ZN(n11458) );
  INV_X1 U5539 ( .A(n11459), .ZN(n24162) );
  AOI22_X1 U5540 ( .A1(\mem[243][0] ), .A2(n11460), .B1(n26887), .B2(
        data_in[0]), .ZN(n11459) );
  INV_X1 U5541 ( .A(n11461), .ZN(n24161) );
  AOI22_X1 U5542 ( .A1(\mem[243][1] ), .A2(n11460), .B1(n26887), .B2(
        data_in[1]), .ZN(n11461) );
  INV_X1 U5543 ( .A(n11462), .ZN(n24160) );
  AOI22_X1 U5544 ( .A1(\mem[243][2] ), .A2(n11460), .B1(n26887), .B2(
        data_in[2]), .ZN(n11462) );
  INV_X1 U5545 ( .A(n11463), .ZN(n24159) );
  AOI22_X1 U5546 ( .A1(\mem[243][3] ), .A2(n11460), .B1(n26887), .B2(
        data_in[3]), .ZN(n11463) );
  INV_X1 U5547 ( .A(n11464), .ZN(n24158) );
  AOI22_X1 U5548 ( .A1(\mem[243][4] ), .A2(n11460), .B1(n26887), .B2(
        data_in[4]), .ZN(n11464) );
  INV_X1 U5549 ( .A(n11465), .ZN(n24157) );
  AOI22_X1 U5550 ( .A1(\mem[243][5] ), .A2(n11460), .B1(n26887), .B2(
        data_in[5]), .ZN(n11465) );
  INV_X1 U5551 ( .A(n11466), .ZN(n24156) );
  AOI22_X1 U5552 ( .A1(\mem[243][6] ), .A2(n11460), .B1(n26887), .B2(
        data_in[6]), .ZN(n11466) );
  INV_X1 U5553 ( .A(n11467), .ZN(n24155) );
  AOI22_X1 U5554 ( .A1(\mem[243][7] ), .A2(n11460), .B1(n26887), .B2(
        data_in[7]), .ZN(n11467) );
  INV_X1 U5555 ( .A(n11468), .ZN(n24154) );
  AOI22_X1 U5556 ( .A1(\mem[244][0] ), .A2(n11469), .B1(n26886), .B2(
        data_in[0]), .ZN(n11468) );
  INV_X1 U5557 ( .A(n11470), .ZN(n24153) );
  AOI22_X1 U5558 ( .A1(\mem[244][1] ), .A2(n11469), .B1(n26886), .B2(
        data_in[1]), .ZN(n11470) );
  INV_X1 U5559 ( .A(n11471), .ZN(n24152) );
  AOI22_X1 U5560 ( .A1(\mem[244][2] ), .A2(n11469), .B1(n26886), .B2(
        data_in[2]), .ZN(n11471) );
  INV_X1 U5561 ( .A(n11472), .ZN(n24151) );
  AOI22_X1 U5562 ( .A1(\mem[244][3] ), .A2(n11469), .B1(n26886), .B2(
        data_in[3]), .ZN(n11472) );
  INV_X1 U5563 ( .A(n11473), .ZN(n24150) );
  AOI22_X1 U5564 ( .A1(\mem[244][4] ), .A2(n11469), .B1(n26886), .B2(
        data_in[4]), .ZN(n11473) );
  INV_X1 U5565 ( .A(n11474), .ZN(n24149) );
  AOI22_X1 U5566 ( .A1(\mem[244][5] ), .A2(n11469), .B1(n26886), .B2(
        data_in[5]), .ZN(n11474) );
  INV_X1 U5567 ( .A(n11475), .ZN(n24148) );
  AOI22_X1 U5568 ( .A1(\mem[244][6] ), .A2(n11469), .B1(n26886), .B2(
        data_in[6]), .ZN(n11475) );
  INV_X1 U5569 ( .A(n11476), .ZN(n24147) );
  AOI22_X1 U5570 ( .A1(\mem[244][7] ), .A2(n11469), .B1(n26886), .B2(
        data_in[7]), .ZN(n11476) );
  INV_X1 U5571 ( .A(n11477), .ZN(n24146) );
  AOI22_X1 U5572 ( .A1(\mem[245][0] ), .A2(n11478), .B1(n26885), .B2(
        data_in[0]), .ZN(n11477) );
  INV_X1 U5573 ( .A(n11479), .ZN(n24145) );
  AOI22_X1 U5574 ( .A1(\mem[245][1] ), .A2(n11478), .B1(n26885), .B2(
        data_in[1]), .ZN(n11479) );
  INV_X1 U5575 ( .A(n11480), .ZN(n24144) );
  AOI22_X1 U5576 ( .A1(\mem[245][2] ), .A2(n11478), .B1(n26885), .B2(
        data_in[2]), .ZN(n11480) );
  INV_X1 U5577 ( .A(n11481), .ZN(n24143) );
  AOI22_X1 U5578 ( .A1(\mem[245][3] ), .A2(n11478), .B1(n26885), .B2(
        data_in[3]), .ZN(n11481) );
  INV_X1 U5579 ( .A(n11482), .ZN(n24142) );
  AOI22_X1 U5580 ( .A1(\mem[245][4] ), .A2(n11478), .B1(n26885), .B2(
        data_in[4]), .ZN(n11482) );
  INV_X1 U5581 ( .A(n11483), .ZN(n24141) );
  AOI22_X1 U5582 ( .A1(\mem[245][5] ), .A2(n11478), .B1(n26885), .B2(
        data_in[5]), .ZN(n11483) );
  INV_X1 U5583 ( .A(n11484), .ZN(n24140) );
  AOI22_X1 U5584 ( .A1(\mem[245][6] ), .A2(n11478), .B1(n26885), .B2(
        data_in[6]), .ZN(n11484) );
  INV_X1 U5585 ( .A(n11485), .ZN(n24139) );
  AOI22_X1 U5586 ( .A1(\mem[245][7] ), .A2(n11478), .B1(n26885), .B2(
        data_in[7]), .ZN(n11485) );
  INV_X1 U5587 ( .A(n11486), .ZN(n24138) );
  AOI22_X1 U5588 ( .A1(\mem[246][0] ), .A2(n11487), .B1(n26884), .B2(
        data_in[0]), .ZN(n11486) );
  INV_X1 U5589 ( .A(n11488), .ZN(n24137) );
  AOI22_X1 U5590 ( .A1(\mem[246][1] ), .A2(n11487), .B1(n26884), .B2(
        data_in[1]), .ZN(n11488) );
  INV_X1 U5591 ( .A(n11489), .ZN(n24136) );
  AOI22_X1 U5592 ( .A1(\mem[246][2] ), .A2(n11487), .B1(n26884), .B2(
        data_in[2]), .ZN(n11489) );
  INV_X1 U5593 ( .A(n11490), .ZN(n24135) );
  AOI22_X1 U5594 ( .A1(\mem[246][3] ), .A2(n11487), .B1(n26884), .B2(
        data_in[3]), .ZN(n11490) );
  INV_X1 U5595 ( .A(n11491), .ZN(n24134) );
  AOI22_X1 U5596 ( .A1(\mem[246][4] ), .A2(n11487), .B1(n26884), .B2(
        data_in[4]), .ZN(n11491) );
  INV_X1 U5597 ( .A(n11492), .ZN(n24133) );
  AOI22_X1 U5598 ( .A1(\mem[246][5] ), .A2(n11487), .B1(n26884), .B2(
        data_in[5]), .ZN(n11492) );
  INV_X1 U5599 ( .A(n11493), .ZN(n24132) );
  AOI22_X1 U5600 ( .A1(\mem[246][6] ), .A2(n11487), .B1(n26884), .B2(
        data_in[6]), .ZN(n11493) );
  INV_X1 U5601 ( .A(n11494), .ZN(n24131) );
  AOI22_X1 U5602 ( .A1(\mem[246][7] ), .A2(n11487), .B1(n26884), .B2(
        data_in[7]), .ZN(n11494) );
  INV_X1 U5603 ( .A(n11495), .ZN(n24130) );
  AOI22_X1 U5604 ( .A1(\mem[247][0] ), .A2(n11496), .B1(n26883), .B2(
        data_in[0]), .ZN(n11495) );
  INV_X1 U5605 ( .A(n11497), .ZN(n24129) );
  AOI22_X1 U5606 ( .A1(\mem[247][1] ), .A2(n11496), .B1(n26883), .B2(
        data_in[1]), .ZN(n11497) );
  INV_X1 U5607 ( .A(n11498), .ZN(n24128) );
  AOI22_X1 U5608 ( .A1(\mem[247][2] ), .A2(n11496), .B1(n26883), .B2(
        data_in[2]), .ZN(n11498) );
  INV_X1 U5609 ( .A(n11499), .ZN(n24127) );
  AOI22_X1 U5610 ( .A1(\mem[247][3] ), .A2(n11496), .B1(n26883), .B2(
        data_in[3]), .ZN(n11499) );
  INV_X1 U5611 ( .A(n11500), .ZN(n24126) );
  AOI22_X1 U5612 ( .A1(\mem[247][4] ), .A2(n11496), .B1(n26883), .B2(
        data_in[4]), .ZN(n11500) );
  INV_X1 U5613 ( .A(n11501), .ZN(n24125) );
  AOI22_X1 U5614 ( .A1(\mem[247][5] ), .A2(n11496), .B1(n26883), .B2(
        data_in[5]), .ZN(n11501) );
  INV_X1 U5615 ( .A(n11502), .ZN(n24124) );
  AOI22_X1 U5616 ( .A1(\mem[247][6] ), .A2(n11496), .B1(n26883), .B2(
        data_in[6]), .ZN(n11502) );
  INV_X1 U5617 ( .A(n11503), .ZN(n24123) );
  AOI22_X1 U5618 ( .A1(\mem[247][7] ), .A2(n11496), .B1(n26883), .B2(
        data_in[7]), .ZN(n11503) );
  INV_X1 U5619 ( .A(n11504), .ZN(n24122) );
  AOI22_X1 U5620 ( .A1(\mem[248][0] ), .A2(n11505), .B1(n26882), .B2(
        data_in[0]), .ZN(n11504) );
  INV_X1 U5621 ( .A(n11506), .ZN(n24121) );
  AOI22_X1 U5622 ( .A1(\mem[248][1] ), .A2(n11505), .B1(n26882), .B2(
        data_in[1]), .ZN(n11506) );
  INV_X1 U5623 ( .A(n11507), .ZN(n24120) );
  AOI22_X1 U5624 ( .A1(\mem[248][2] ), .A2(n11505), .B1(n26882), .B2(
        data_in[2]), .ZN(n11507) );
  INV_X1 U5625 ( .A(n11508), .ZN(n24119) );
  AOI22_X1 U5626 ( .A1(\mem[248][3] ), .A2(n11505), .B1(n26882), .B2(
        data_in[3]), .ZN(n11508) );
  INV_X1 U5627 ( .A(n11509), .ZN(n24118) );
  AOI22_X1 U5628 ( .A1(\mem[248][4] ), .A2(n11505), .B1(n26882), .B2(
        data_in[4]), .ZN(n11509) );
  INV_X1 U5629 ( .A(n11510), .ZN(n24117) );
  AOI22_X1 U5630 ( .A1(\mem[248][5] ), .A2(n11505), .B1(n26882), .B2(
        data_in[5]), .ZN(n11510) );
  INV_X1 U5631 ( .A(n11511), .ZN(n24116) );
  AOI22_X1 U5632 ( .A1(\mem[248][6] ), .A2(n11505), .B1(n26882), .B2(
        data_in[6]), .ZN(n11511) );
  INV_X1 U5633 ( .A(n11512), .ZN(n24115) );
  AOI22_X1 U5634 ( .A1(\mem[248][7] ), .A2(n11505), .B1(n26882), .B2(
        data_in[7]), .ZN(n11512) );
  INV_X1 U5635 ( .A(n11513), .ZN(n24114) );
  AOI22_X1 U5636 ( .A1(\mem[249][0] ), .A2(n11514), .B1(n26881), .B2(
        data_in[0]), .ZN(n11513) );
  INV_X1 U5637 ( .A(n11515), .ZN(n24113) );
  AOI22_X1 U5638 ( .A1(\mem[249][1] ), .A2(n11514), .B1(n26881), .B2(
        data_in[1]), .ZN(n11515) );
  INV_X1 U5639 ( .A(n11516), .ZN(n24112) );
  AOI22_X1 U5640 ( .A1(\mem[249][2] ), .A2(n11514), .B1(n26881), .B2(
        data_in[2]), .ZN(n11516) );
  INV_X1 U5641 ( .A(n11517), .ZN(n24111) );
  AOI22_X1 U5642 ( .A1(\mem[249][3] ), .A2(n11514), .B1(n26881), .B2(
        data_in[3]), .ZN(n11517) );
  INV_X1 U5643 ( .A(n11518), .ZN(n24110) );
  AOI22_X1 U5644 ( .A1(\mem[249][4] ), .A2(n11514), .B1(n26881), .B2(
        data_in[4]), .ZN(n11518) );
  INV_X1 U5645 ( .A(n11519), .ZN(n24109) );
  AOI22_X1 U5646 ( .A1(\mem[249][5] ), .A2(n11514), .B1(n26881), .B2(
        data_in[5]), .ZN(n11519) );
  INV_X1 U5647 ( .A(n11520), .ZN(n24108) );
  AOI22_X1 U5648 ( .A1(\mem[249][6] ), .A2(n11514), .B1(n26881), .B2(
        data_in[6]), .ZN(n11520) );
  INV_X1 U5649 ( .A(n11521), .ZN(n24107) );
  AOI22_X1 U5650 ( .A1(\mem[249][7] ), .A2(n11514), .B1(n26881), .B2(
        data_in[7]), .ZN(n11521) );
  INV_X1 U5651 ( .A(n11522), .ZN(n24106) );
  AOI22_X1 U5652 ( .A1(\mem[250][0] ), .A2(n11523), .B1(n26880), .B2(
        data_in[0]), .ZN(n11522) );
  INV_X1 U5653 ( .A(n11524), .ZN(n24105) );
  AOI22_X1 U5654 ( .A1(\mem[250][1] ), .A2(n11523), .B1(n26880), .B2(
        data_in[1]), .ZN(n11524) );
  INV_X1 U5655 ( .A(n11525), .ZN(n24104) );
  AOI22_X1 U5656 ( .A1(\mem[250][2] ), .A2(n11523), .B1(n26880), .B2(
        data_in[2]), .ZN(n11525) );
  INV_X1 U5657 ( .A(n11526), .ZN(n24103) );
  AOI22_X1 U5658 ( .A1(\mem[250][3] ), .A2(n11523), .B1(n26880), .B2(
        data_in[3]), .ZN(n11526) );
  INV_X1 U5659 ( .A(n11527), .ZN(n24102) );
  AOI22_X1 U5660 ( .A1(\mem[250][4] ), .A2(n11523), .B1(n26880), .B2(
        data_in[4]), .ZN(n11527) );
  INV_X1 U5661 ( .A(n11528), .ZN(n24101) );
  AOI22_X1 U5662 ( .A1(\mem[250][5] ), .A2(n11523), .B1(n26880), .B2(
        data_in[5]), .ZN(n11528) );
  INV_X1 U5663 ( .A(n11529), .ZN(n24100) );
  AOI22_X1 U5664 ( .A1(\mem[250][6] ), .A2(n11523), .B1(n26880), .B2(
        data_in[6]), .ZN(n11529) );
  INV_X1 U5665 ( .A(n11530), .ZN(n24099) );
  AOI22_X1 U5666 ( .A1(\mem[250][7] ), .A2(n11523), .B1(n26880), .B2(
        data_in[7]), .ZN(n11530) );
  INV_X1 U5667 ( .A(n11531), .ZN(n24098) );
  AOI22_X1 U5668 ( .A1(\mem[251][0] ), .A2(n11532), .B1(n26879), .B2(
        data_in[0]), .ZN(n11531) );
  INV_X1 U5669 ( .A(n11533), .ZN(n24097) );
  AOI22_X1 U5670 ( .A1(\mem[251][1] ), .A2(n11532), .B1(n26879), .B2(
        data_in[1]), .ZN(n11533) );
  INV_X1 U5671 ( .A(n11534), .ZN(n24096) );
  AOI22_X1 U5672 ( .A1(\mem[251][2] ), .A2(n11532), .B1(n26879), .B2(
        data_in[2]), .ZN(n11534) );
  INV_X1 U5673 ( .A(n11535), .ZN(n24095) );
  AOI22_X1 U5674 ( .A1(\mem[251][3] ), .A2(n11532), .B1(n26879), .B2(
        data_in[3]), .ZN(n11535) );
  INV_X1 U5675 ( .A(n11536), .ZN(n24094) );
  AOI22_X1 U5676 ( .A1(\mem[251][4] ), .A2(n11532), .B1(n26879), .B2(
        data_in[4]), .ZN(n11536) );
  INV_X1 U5677 ( .A(n11537), .ZN(n24093) );
  AOI22_X1 U5678 ( .A1(\mem[251][5] ), .A2(n11532), .B1(n26879), .B2(
        data_in[5]), .ZN(n11537) );
  INV_X1 U5679 ( .A(n11538), .ZN(n24092) );
  AOI22_X1 U5680 ( .A1(\mem[251][6] ), .A2(n11532), .B1(n26879), .B2(
        data_in[6]), .ZN(n11538) );
  INV_X1 U5681 ( .A(n11539), .ZN(n24091) );
  AOI22_X1 U5682 ( .A1(\mem[251][7] ), .A2(n11532), .B1(n26879), .B2(
        data_in[7]), .ZN(n11539) );
  INV_X1 U5683 ( .A(n11540), .ZN(n24090) );
  AOI22_X1 U5684 ( .A1(\mem[252][0] ), .A2(n11541), .B1(n26878), .B2(
        data_in[0]), .ZN(n11540) );
  INV_X1 U5685 ( .A(n11542), .ZN(n24089) );
  AOI22_X1 U5686 ( .A1(\mem[252][1] ), .A2(n11541), .B1(n26878), .B2(
        data_in[1]), .ZN(n11542) );
  INV_X1 U5687 ( .A(n11543), .ZN(n24088) );
  AOI22_X1 U5688 ( .A1(\mem[252][2] ), .A2(n11541), .B1(n26878), .B2(
        data_in[2]), .ZN(n11543) );
  INV_X1 U5689 ( .A(n11544), .ZN(n24087) );
  AOI22_X1 U5690 ( .A1(\mem[252][3] ), .A2(n11541), .B1(n26878), .B2(
        data_in[3]), .ZN(n11544) );
  INV_X1 U5691 ( .A(n11545), .ZN(n24086) );
  AOI22_X1 U5692 ( .A1(\mem[252][4] ), .A2(n11541), .B1(n26878), .B2(
        data_in[4]), .ZN(n11545) );
  INV_X1 U5693 ( .A(n11546), .ZN(n24085) );
  AOI22_X1 U5694 ( .A1(\mem[252][5] ), .A2(n11541), .B1(n26878), .B2(
        data_in[5]), .ZN(n11546) );
  INV_X1 U5695 ( .A(n11547), .ZN(n24084) );
  AOI22_X1 U5696 ( .A1(\mem[252][6] ), .A2(n11541), .B1(n26878), .B2(
        data_in[6]), .ZN(n11547) );
  INV_X1 U5697 ( .A(n11548), .ZN(n24083) );
  AOI22_X1 U5698 ( .A1(\mem[252][7] ), .A2(n11541), .B1(n26878), .B2(
        data_in[7]), .ZN(n11548) );
  INV_X1 U5699 ( .A(n11549), .ZN(n24082) );
  AOI22_X1 U5700 ( .A1(\mem[253][0] ), .A2(n11550), .B1(n26877), .B2(
        data_in[0]), .ZN(n11549) );
  INV_X1 U5701 ( .A(n11551), .ZN(n24081) );
  AOI22_X1 U5702 ( .A1(\mem[253][1] ), .A2(n11550), .B1(n26877), .B2(
        data_in[1]), .ZN(n11551) );
  INV_X1 U5703 ( .A(n11552), .ZN(n24080) );
  AOI22_X1 U5704 ( .A1(\mem[253][2] ), .A2(n11550), .B1(n26877), .B2(
        data_in[2]), .ZN(n11552) );
  INV_X1 U5705 ( .A(n11553), .ZN(n24079) );
  AOI22_X1 U5706 ( .A1(\mem[253][3] ), .A2(n11550), .B1(n26877), .B2(
        data_in[3]), .ZN(n11553) );
  INV_X1 U5707 ( .A(n11554), .ZN(n24078) );
  AOI22_X1 U5708 ( .A1(\mem[253][4] ), .A2(n11550), .B1(n26877), .B2(
        data_in[4]), .ZN(n11554) );
  INV_X1 U5709 ( .A(n11555), .ZN(n24077) );
  AOI22_X1 U5710 ( .A1(\mem[253][5] ), .A2(n11550), .B1(n26877), .B2(
        data_in[5]), .ZN(n11555) );
  INV_X1 U5711 ( .A(n11556), .ZN(n24076) );
  AOI22_X1 U5712 ( .A1(\mem[253][6] ), .A2(n11550), .B1(n26877), .B2(
        data_in[6]), .ZN(n11556) );
  INV_X1 U5713 ( .A(n11557), .ZN(n24075) );
  AOI22_X1 U5714 ( .A1(\mem[253][7] ), .A2(n11550), .B1(n26877), .B2(
        data_in[7]), .ZN(n11557) );
  INV_X1 U5715 ( .A(n11558), .ZN(n24074) );
  AOI22_X1 U5716 ( .A1(\mem[254][0] ), .A2(n11559), .B1(n26876), .B2(
        data_in[0]), .ZN(n11558) );
  INV_X1 U5717 ( .A(n11560), .ZN(n24073) );
  AOI22_X1 U5718 ( .A1(\mem[254][1] ), .A2(n11559), .B1(n26876), .B2(
        data_in[1]), .ZN(n11560) );
  INV_X1 U5719 ( .A(n11561), .ZN(n24072) );
  AOI22_X1 U5720 ( .A1(\mem[254][2] ), .A2(n11559), .B1(n26876), .B2(
        data_in[2]), .ZN(n11561) );
  INV_X1 U5721 ( .A(n11562), .ZN(n24071) );
  AOI22_X1 U5722 ( .A1(\mem[254][3] ), .A2(n11559), .B1(n26876), .B2(
        data_in[3]), .ZN(n11562) );
  INV_X1 U5723 ( .A(n11563), .ZN(n24070) );
  AOI22_X1 U5724 ( .A1(\mem[254][4] ), .A2(n11559), .B1(n26876), .B2(
        data_in[4]), .ZN(n11563) );
  INV_X1 U5725 ( .A(n11564), .ZN(n24069) );
  AOI22_X1 U5726 ( .A1(\mem[254][5] ), .A2(n11559), .B1(n26876), .B2(
        data_in[5]), .ZN(n11564) );
  INV_X1 U5727 ( .A(n11565), .ZN(n24068) );
  AOI22_X1 U5728 ( .A1(\mem[254][6] ), .A2(n11559), .B1(n26876), .B2(
        data_in[6]), .ZN(n11565) );
  INV_X1 U5729 ( .A(n11566), .ZN(n24067) );
  AOI22_X1 U5730 ( .A1(\mem[254][7] ), .A2(n11559), .B1(n26876), .B2(
        data_in[7]), .ZN(n11566) );
  INV_X1 U5731 ( .A(n11567), .ZN(n24066) );
  AOI22_X1 U5732 ( .A1(\mem[255][0] ), .A2(n11568), .B1(n26875), .B2(
        data_in[0]), .ZN(n11567) );
  INV_X1 U5733 ( .A(n11569), .ZN(n24065) );
  AOI22_X1 U5734 ( .A1(\mem[255][1] ), .A2(n11568), .B1(n26875), .B2(
        data_in[1]), .ZN(n11569) );
  INV_X1 U5735 ( .A(n11570), .ZN(n24064) );
  AOI22_X1 U5736 ( .A1(\mem[255][2] ), .A2(n11568), .B1(n26875), .B2(
        data_in[2]), .ZN(n11570) );
  INV_X1 U5737 ( .A(n11571), .ZN(n24063) );
  AOI22_X1 U5738 ( .A1(\mem[255][3] ), .A2(n11568), .B1(n26875), .B2(
        data_in[3]), .ZN(n11571) );
  INV_X1 U5739 ( .A(n11572), .ZN(n24062) );
  AOI22_X1 U5740 ( .A1(\mem[255][4] ), .A2(n11568), .B1(n26875), .B2(
        data_in[4]), .ZN(n11572) );
  INV_X1 U5741 ( .A(n11573), .ZN(n24061) );
  AOI22_X1 U5742 ( .A1(\mem[255][5] ), .A2(n11568), .B1(n26875), .B2(
        data_in[5]), .ZN(n11573) );
  INV_X1 U5743 ( .A(n11574), .ZN(n24060) );
  AOI22_X1 U5744 ( .A1(\mem[255][6] ), .A2(n11568), .B1(n26875), .B2(
        data_in[6]), .ZN(n11574) );
  INV_X1 U5745 ( .A(n11575), .ZN(n24059) );
  AOI22_X1 U5746 ( .A1(\mem[255][7] ), .A2(n11568), .B1(n26875), .B2(
        data_in[7]), .ZN(n11575) );
  INV_X1 U5747 ( .A(n11650), .ZN(n23994) );
  AOI22_X1 U5748 ( .A1(\mem[264][0] ), .A2(n11651), .B1(n26866), .B2(
        data_in[0]), .ZN(n11650) );
  INV_X1 U5749 ( .A(n11652), .ZN(n23993) );
  AOI22_X1 U5750 ( .A1(\mem[264][1] ), .A2(n11651), .B1(n26866), .B2(
        data_in[1]), .ZN(n11652) );
  INV_X1 U5751 ( .A(n11653), .ZN(n23992) );
  AOI22_X1 U5752 ( .A1(\mem[264][2] ), .A2(n11651), .B1(n26866), .B2(
        data_in[2]), .ZN(n11653) );
  INV_X1 U5753 ( .A(n11654), .ZN(n23991) );
  AOI22_X1 U5754 ( .A1(\mem[264][3] ), .A2(n11651), .B1(n26866), .B2(
        data_in[3]), .ZN(n11654) );
  INV_X1 U5755 ( .A(n11655), .ZN(n23990) );
  AOI22_X1 U5756 ( .A1(\mem[264][4] ), .A2(n11651), .B1(n26866), .B2(
        data_in[4]), .ZN(n11655) );
  INV_X1 U5757 ( .A(n11656), .ZN(n23989) );
  AOI22_X1 U5758 ( .A1(\mem[264][5] ), .A2(n11651), .B1(n26866), .B2(
        data_in[5]), .ZN(n11656) );
  INV_X1 U5759 ( .A(n11657), .ZN(n23988) );
  AOI22_X1 U5760 ( .A1(\mem[264][6] ), .A2(n11651), .B1(n26866), .B2(
        data_in[6]), .ZN(n11657) );
  INV_X1 U5761 ( .A(n11658), .ZN(n23987) );
  AOI22_X1 U5762 ( .A1(\mem[264][7] ), .A2(n11651), .B1(n26866), .B2(
        data_in[7]), .ZN(n11658) );
  INV_X1 U5763 ( .A(n11659), .ZN(n23986) );
  AOI22_X1 U5764 ( .A1(\mem[265][0] ), .A2(n11660), .B1(n26865), .B2(
        data_in[0]), .ZN(n11659) );
  INV_X1 U5765 ( .A(n11661), .ZN(n23985) );
  AOI22_X1 U5766 ( .A1(\mem[265][1] ), .A2(n11660), .B1(n26865), .B2(
        data_in[1]), .ZN(n11661) );
  INV_X1 U5767 ( .A(n11662), .ZN(n23984) );
  AOI22_X1 U5768 ( .A1(\mem[265][2] ), .A2(n11660), .B1(n26865), .B2(
        data_in[2]), .ZN(n11662) );
  INV_X1 U5769 ( .A(n11663), .ZN(n23983) );
  AOI22_X1 U5770 ( .A1(\mem[265][3] ), .A2(n11660), .B1(n26865), .B2(
        data_in[3]), .ZN(n11663) );
  INV_X1 U5771 ( .A(n11664), .ZN(n23982) );
  AOI22_X1 U5772 ( .A1(\mem[265][4] ), .A2(n11660), .B1(n26865), .B2(
        data_in[4]), .ZN(n11664) );
  INV_X1 U5773 ( .A(n11665), .ZN(n23981) );
  AOI22_X1 U5774 ( .A1(\mem[265][5] ), .A2(n11660), .B1(n26865), .B2(
        data_in[5]), .ZN(n11665) );
  INV_X1 U5775 ( .A(n11666), .ZN(n23980) );
  AOI22_X1 U5776 ( .A1(\mem[265][6] ), .A2(n11660), .B1(n26865), .B2(
        data_in[6]), .ZN(n11666) );
  INV_X1 U5777 ( .A(n11667), .ZN(n23979) );
  AOI22_X1 U5778 ( .A1(\mem[265][7] ), .A2(n11660), .B1(n26865), .B2(
        data_in[7]), .ZN(n11667) );
  INV_X1 U5779 ( .A(n11668), .ZN(n23978) );
  AOI22_X1 U5780 ( .A1(\mem[266][0] ), .A2(n11669), .B1(n26864), .B2(
        data_in[0]), .ZN(n11668) );
  INV_X1 U5781 ( .A(n11670), .ZN(n23977) );
  AOI22_X1 U5782 ( .A1(\mem[266][1] ), .A2(n11669), .B1(n26864), .B2(
        data_in[1]), .ZN(n11670) );
  INV_X1 U5783 ( .A(n11671), .ZN(n23976) );
  AOI22_X1 U5784 ( .A1(\mem[266][2] ), .A2(n11669), .B1(n26864), .B2(
        data_in[2]), .ZN(n11671) );
  INV_X1 U5785 ( .A(n11672), .ZN(n23975) );
  AOI22_X1 U5786 ( .A1(\mem[266][3] ), .A2(n11669), .B1(n26864), .B2(
        data_in[3]), .ZN(n11672) );
  INV_X1 U5787 ( .A(n11673), .ZN(n23974) );
  AOI22_X1 U5788 ( .A1(\mem[266][4] ), .A2(n11669), .B1(n26864), .B2(
        data_in[4]), .ZN(n11673) );
  INV_X1 U5789 ( .A(n11674), .ZN(n23973) );
  AOI22_X1 U5790 ( .A1(\mem[266][5] ), .A2(n11669), .B1(n26864), .B2(
        data_in[5]), .ZN(n11674) );
  INV_X1 U5791 ( .A(n11675), .ZN(n23972) );
  AOI22_X1 U5792 ( .A1(\mem[266][6] ), .A2(n11669), .B1(n26864), .B2(
        data_in[6]), .ZN(n11675) );
  INV_X1 U5793 ( .A(n11676), .ZN(n23971) );
  AOI22_X1 U5794 ( .A1(\mem[266][7] ), .A2(n11669), .B1(n26864), .B2(
        data_in[7]), .ZN(n11676) );
  INV_X1 U5795 ( .A(n11677), .ZN(n23970) );
  AOI22_X1 U5796 ( .A1(\mem[267][0] ), .A2(n11678), .B1(n26863), .B2(
        data_in[0]), .ZN(n11677) );
  INV_X1 U5797 ( .A(n11679), .ZN(n23969) );
  AOI22_X1 U5798 ( .A1(\mem[267][1] ), .A2(n11678), .B1(n26863), .B2(
        data_in[1]), .ZN(n11679) );
  INV_X1 U5799 ( .A(n11680), .ZN(n23968) );
  AOI22_X1 U5800 ( .A1(\mem[267][2] ), .A2(n11678), .B1(n26863), .B2(
        data_in[2]), .ZN(n11680) );
  INV_X1 U5801 ( .A(n11681), .ZN(n23967) );
  AOI22_X1 U5802 ( .A1(\mem[267][3] ), .A2(n11678), .B1(n26863), .B2(
        data_in[3]), .ZN(n11681) );
  INV_X1 U5803 ( .A(n11682), .ZN(n23966) );
  AOI22_X1 U5804 ( .A1(\mem[267][4] ), .A2(n11678), .B1(n26863), .B2(
        data_in[4]), .ZN(n11682) );
  INV_X1 U5805 ( .A(n11683), .ZN(n23965) );
  AOI22_X1 U5806 ( .A1(\mem[267][5] ), .A2(n11678), .B1(n26863), .B2(
        data_in[5]), .ZN(n11683) );
  INV_X1 U5807 ( .A(n11684), .ZN(n23964) );
  AOI22_X1 U5808 ( .A1(\mem[267][6] ), .A2(n11678), .B1(n26863), .B2(
        data_in[6]), .ZN(n11684) );
  INV_X1 U5809 ( .A(n11685), .ZN(n23963) );
  AOI22_X1 U5810 ( .A1(\mem[267][7] ), .A2(n11678), .B1(n26863), .B2(
        data_in[7]), .ZN(n11685) );
  INV_X1 U5811 ( .A(n11686), .ZN(n23962) );
  AOI22_X1 U5812 ( .A1(\mem[268][0] ), .A2(n11687), .B1(n26862), .B2(
        data_in[0]), .ZN(n11686) );
  INV_X1 U5813 ( .A(n11688), .ZN(n23961) );
  AOI22_X1 U5814 ( .A1(\mem[268][1] ), .A2(n11687), .B1(n26862), .B2(
        data_in[1]), .ZN(n11688) );
  INV_X1 U5815 ( .A(n11689), .ZN(n23960) );
  AOI22_X1 U5816 ( .A1(\mem[268][2] ), .A2(n11687), .B1(n26862), .B2(
        data_in[2]), .ZN(n11689) );
  INV_X1 U5817 ( .A(n11690), .ZN(n23959) );
  AOI22_X1 U5818 ( .A1(\mem[268][3] ), .A2(n11687), .B1(n26862), .B2(
        data_in[3]), .ZN(n11690) );
  INV_X1 U5819 ( .A(n11691), .ZN(n23958) );
  AOI22_X1 U5820 ( .A1(\mem[268][4] ), .A2(n11687), .B1(n26862), .B2(
        data_in[4]), .ZN(n11691) );
  INV_X1 U5821 ( .A(n11692), .ZN(n23957) );
  AOI22_X1 U5822 ( .A1(\mem[268][5] ), .A2(n11687), .B1(n26862), .B2(
        data_in[5]), .ZN(n11692) );
  INV_X1 U5823 ( .A(n11693), .ZN(n23956) );
  AOI22_X1 U5824 ( .A1(\mem[268][6] ), .A2(n11687), .B1(n26862), .B2(
        data_in[6]), .ZN(n11693) );
  INV_X1 U5825 ( .A(n11694), .ZN(n23955) );
  AOI22_X1 U5826 ( .A1(\mem[268][7] ), .A2(n11687), .B1(n26862), .B2(
        data_in[7]), .ZN(n11694) );
  INV_X1 U5827 ( .A(n11695), .ZN(n23954) );
  AOI22_X1 U5828 ( .A1(\mem[269][0] ), .A2(n11696), .B1(n26861), .B2(
        data_in[0]), .ZN(n11695) );
  INV_X1 U5829 ( .A(n11697), .ZN(n23953) );
  AOI22_X1 U5830 ( .A1(\mem[269][1] ), .A2(n11696), .B1(n26861), .B2(
        data_in[1]), .ZN(n11697) );
  INV_X1 U5831 ( .A(n11698), .ZN(n23952) );
  AOI22_X1 U5832 ( .A1(\mem[269][2] ), .A2(n11696), .B1(n26861), .B2(
        data_in[2]), .ZN(n11698) );
  INV_X1 U5833 ( .A(n11699), .ZN(n23951) );
  AOI22_X1 U5834 ( .A1(\mem[269][3] ), .A2(n11696), .B1(n26861), .B2(
        data_in[3]), .ZN(n11699) );
  INV_X1 U5835 ( .A(n11700), .ZN(n23950) );
  AOI22_X1 U5836 ( .A1(\mem[269][4] ), .A2(n11696), .B1(n26861), .B2(
        data_in[4]), .ZN(n11700) );
  INV_X1 U5837 ( .A(n11701), .ZN(n23949) );
  AOI22_X1 U5838 ( .A1(\mem[269][5] ), .A2(n11696), .B1(n26861), .B2(
        data_in[5]), .ZN(n11701) );
  INV_X1 U5839 ( .A(n11702), .ZN(n23948) );
  AOI22_X1 U5840 ( .A1(\mem[269][6] ), .A2(n11696), .B1(n26861), .B2(
        data_in[6]), .ZN(n11702) );
  INV_X1 U5841 ( .A(n11703), .ZN(n23947) );
  AOI22_X1 U5842 ( .A1(\mem[269][7] ), .A2(n11696), .B1(n26861), .B2(
        data_in[7]), .ZN(n11703) );
  INV_X1 U5843 ( .A(n11704), .ZN(n23946) );
  AOI22_X1 U5844 ( .A1(\mem[270][0] ), .A2(n11705), .B1(n26860), .B2(
        data_in[0]), .ZN(n11704) );
  INV_X1 U5845 ( .A(n11706), .ZN(n23945) );
  AOI22_X1 U5846 ( .A1(\mem[270][1] ), .A2(n11705), .B1(n26860), .B2(
        data_in[1]), .ZN(n11706) );
  INV_X1 U5847 ( .A(n11707), .ZN(n23944) );
  AOI22_X1 U5848 ( .A1(\mem[270][2] ), .A2(n11705), .B1(n26860), .B2(
        data_in[2]), .ZN(n11707) );
  INV_X1 U5849 ( .A(n11708), .ZN(n23943) );
  AOI22_X1 U5850 ( .A1(\mem[270][3] ), .A2(n11705), .B1(n26860), .B2(
        data_in[3]), .ZN(n11708) );
  INV_X1 U5851 ( .A(n11709), .ZN(n23942) );
  AOI22_X1 U5852 ( .A1(\mem[270][4] ), .A2(n11705), .B1(n26860), .B2(
        data_in[4]), .ZN(n11709) );
  INV_X1 U5853 ( .A(n11710), .ZN(n23941) );
  AOI22_X1 U5854 ( .A1(\mem[270][5] ), .A2(n11705), .B1(n26860), .B2(
        data_in[5]), .ZN(n11710) );
  INV_X1 U5855 ( .A(n11711), .ZN(n23940) );
  AOI22_X1 U5856 ( .A1(\mem[270][6] ), .A2(n11705), .B1(n26860), .B2(
        data_in[6]), .ZN(n11711) );
  INV_X1 U5857 ( .A(n11712), .ZN(n23939) );
  AOI22_X1 U5858 ( .A1(\mem[270][7] ), .A2(n11705), .B1(n26860), .B2(
        data_in[7]), .ZN(n11712) );
  INV_X1 U5859 ( .A(n11713), .ZN(n23938) );
  AOI22_X1 U5860 ( .A1(\mem[271][0] ), .A2(n11714), .B1(n26859), .B2(
        data_in[0]), .ZN(n11713) );
  INV_X1 U5861 ( .A(n11715), .ZN(n23937) );
  AOI22_X1 U5862 ( .A1(\mem[271][1] ), .A2(n11714), .B1(n26859), .B2(
        data_in[1]), .ZN(n11715) );
  INV_X1 U5863 ( .A(n11716), .ZN(n23936) );
  AOI22_X1 U5864 ( .A1(\mem[271][2] ), .A2(n11714), .B1(n26859), .B2(
        data_in[2]), .ZN(n11716) );
  INV_X1 U5865 ( .A(n11717), .ZN(n23935) );
  AOI22_X1 U5866 ( .A1(\mem[271][3] ), .A2(n11714), .B1(n26859), .B2(
        data_in[3]), .ZN(n11717) );
  INV_X1 U5867 ( .A(n11718), .ZN(n23934) );
  AOI22_X1 U5868 ( .A1(\mem[271][4] ), .A2(n11714), .B1(n26859), .B2(
        data_in[4]), .ZN(n11718) );
  INV_X1 U5869 ( .A(n11719), .ZN(n23933) );
  AOI22_X1 U5870 ( .A1(\mem[271][5] ), .A2(n11714), .B1(n26859), .B2(
        data_in[5]), .ZN(n11719) );
  INV_X1 U5871 ( .A(n11720), .ZN(n23932) );
  AOI22_X1 U5872 ( .A1(\mem[271][6] ), .A2(n11714), .B1(n26859), .B2(
        data_in[6]), .ZN(n11720) );
  INV_X1 U5873 ( .A(n11721), .ZN(n23931) );
  AOI22_X1 U5874 ( .A1(\mem[271][7] ), .A2(n11714), .B1(n26859), .B2(
        data_in[7]), .ZN(n11721) );
  INV_X1 U5875 ( .A(n11722), .ZN(n23930) );
  AOI22_X1 U5876 ( .A1(\mem[272][0] ), .A2(n11723), .B1(n26858), .B2(
        data_in[0]), .ZN(n11722) );
  INV_X1 U5877 ( .A(n11724), .ZN(n23929) );
  AOI22_X1 U5878 ( .A1(\mem[272][1] ), .A2(n11723), .B1(n26858), .B2(
        data_in[1]), .ZN(n11724) );
  INV_X1 U5879 ( .A(n11725), .ZN(n23928) );
  AOI22_X1 U5880 ( .A1(\mem[272][2] ), .A2(n11723), .B1(n26858), .B2(
        data_in[2]), .ZN(n11725) );
  INV_X1 U5881 ( .A(n11726), .ZN(n23927) );
  AOI22_X1 U5882 ( .A1(\mem[272][3] ), .A2(n11723), .B1(n26858), .B2(
        data_in[3]), .ZN(n11726) );
  INV_X1 U5883 ( .A(n11727), .ZN(n23926) );
  AOI22_X1 U5884 ( .A1(\mem[272][4] ), .A2(n11723), .B1(n26858), .B2(
        data_in[4]), .ZN(n11727) );
  INV_X1 U5885 ( .A(n11728), .ZN(n23925) );
  AOI22_X1 U5886 ( .A1(\mem[272][5] ), .A2(n11723), .B1(n26858), .B2(
        data_in[5]), .ZN(n11728) );
  INV_X1 U5887 ( .A(n11729), .ZN(n23924) );
  AOI22_X1 U5888 ( .A1(\mem[272][6] ), .A2(n11723), .B1(n26858), .B2(
        data_in[6]), .ZN(n11729) );
  INV_X1 U5889 ( .A(n11730), .ZN(n23923) );
  AOI22_X1 U5890 ( .A1(\mem[272][7] ), .A2(n11723), .B1(n26858), .B2(
        data_in[7]), .ZN(n11730) );
  INV_X1 U5891 ( .A(n11731), .ZN(n23922) );
  AOI22_X1 U5892 ( .A1(\mem[273][0] ), .A2(n11732), .B1(n26857), .B2(
        data_in[0]), .ZN(n11731) );
  INV_X1 U5893 ( .A(n11733), .ZN(n23921) );
  AOI22_X1 U5894 ( .A1(\mem[273][1] ), .A2(n11732), .B1(n26857), .B2(
        data_in[1]), .ZN(n11733) );
  INV_X1 U5895 ( .A(n11734), .ZN(n23920) );
  AOI22_X1 U5896 ( .A1(\mem[273][2] ), .A2(n11732), .B1(n26857), .B2(
        data_in[2]), .ZN(n11734) );
  INV_X1 U5897 ( .A(n11735), .ZN(n23919) );
  AOI22_X1 U5898 ( .A1(\mem[273][3] ), .A2(n11732), .B1(n26857), .B2(
        data_in[3]), .ZN(n11735) );
  INV_X1 U5899 ( .A(n11736), .ZN(n23918) );
  AOI22_X1 U5900 ( .A1(\mem[273][4] ), .A2(n11732), .B1(n26857), .B2(
        data_in[4]), .ZN(n11736) );
  INV_X1 U5901 ( .A(n11737), .ZN(n23917) );
  AOI22_X1 U5902 ( .A1(\mem[273][5] ), .A2(n11732), .B1(n26857), .B2(
        data_in[5]), .ZN(n11737) );
  INV_X1 U5903 ( .A(n11738), .ZN(n23916) );
  AOI22_X1 U5904 ( .A1(\mem[273][6] ), .A2(n11732), .B1(n26857), .B2(
        data_in[6]), .ZN(n11738) );
  INV_X1 U5905 ( .A(n11739), .ZN(n23915) );
  AOI22_X1 U5906 ( .A1(\mem[273][7] ), .A2(n11732), .B1(n26857), .B2(
        data_in[7]), .ZN(n11739) );
  INV_X1 U5907 ( .A(n11740), .ZN(n23914) );
  AOI22_X1 U5908 ( .A1(\mem[274][0] ), .A2(n11741), .B1(n26856), .B2(
        data_in[0]), .ZN(n11740) );
  INV_X1 U5909 ( .A(n11742), .ZN(n23913) );
  AOI22_X1 U5910 ( .A1(\mem[274][1] ), .A2(n11741), .B1(n26856), .B2(
        data_in[1]), .ZN(n11742) );
  INV_X1 U5911 ( .A(n11743), .ZN(n23912) );
  AOI22_X1 U5912 ( .A1(\mem[274][2] ), .A2(n11741), .B1(n26856), .B2(
        data_in[2]), .ZN(n11743) );
  INV_X1 U5913 ( .A(n11744), .ZN(n23911) );
  AOI22_X1 U5914 ( .A1(\mem[274][3] ), .A2(n11741), .B1(n26856), .B2(
        data_in[3]), .ZN(n11744) );
  INV_X1 U5915 ( .A(n11745), .ZN(n23910) );
  AOI22_X1 U5916 ( .A1(\mem[274][4] ), .A2(n11741), .B1(n26856), .B2(
        data_in[4]), .ZN(n11745) );
  INV_X1 U5917 ( .A(n11746), .ZN(n23909) );
  AOI22_X1 U5918 ( .A1(\mem[274][5] ), .A2(n11741), .B1(n26856), .B2(
        data_in[5]), .ZN(n11746) );
  INV_X1 U5919 ( .A(n11747), .ZN(n23908) );
  AOI22_X1 U5920 ( .A1(\mem[274][6] ), .A2(n11741), .B1(n26856), .B2(
        data_in[6]), .ZN(n11747) );
  INV_X1 U5921 ( .A(n11748), .ZN(n23907) );
  AOI22_X1 U5922 ( .A1(\mem[274][7] ), .A2(n11741), .B1(n26856), .B2(
        data_in[7]), .ZN(n11748) );
  INV_X1 U5923 ( .A(n11749), .ZN(n23906) );
  AOI22_X1 U5924 ( .A1(\mem[275][0] ), .A2(n11750), .B1(n26855), .B2(
        data_in[0]), .ZN(n11749) );
  INV_X1 U5925 ( .A(n11751), .ZN(n23905) );
  AOI22_X1 U5926 ( .A1(\mem[275][1] ), .A2(n11750), .B1(n26855), .B2(
        data_in[1]), .ZN(n11751) );
  INV_X1 U5927 ( .A(n11752), .ZN(n23904) );
  AOI22_X1 U5928 ( .A1(\mem[275][2] ), .A2(n11750), .B1(n26855), .B2(
        data_in[2]), .ZN(n11752) );
  INV_X1 U5929 ( .A(n11753), .ZN(n23903) );
  AOI22_X1 U5930 ( .A1(\mem[275][3] ), .A2(n11750), .B1(n26855), .B2(
        data_in[3]), .ZN(n11753) );
  INV_X1 U5931 ( .A(n11754), .ZN(n23902) );
  AOI22_X1 U5932 ( .A1(\mem[275][4] ), .A2(n11750), .B1(n26855), .B2(
        data_in[4]), .ZN(n11754) );
  INV_X1 U5933 ( .A(n11755), .ZN(n23901) );
  AOI22_X1 U5934 ( .A1(\mem[275][5] ), .A2(n11750), .B1(n26855), .B2(
        data_in[5]), .ZN(n11755) );
  INV_X1 U5935 ( .A(n11756), .ZN(n23900) );
  AOI22_X1 U5936 ( .A1(\mem[275][6] ), .A2(n11750), .B1(n26855), .B2(
        data_in[6]), .ZN(n11756) );
  INV_X1 U5937 ( .A(n11757), .ZN(n23899) );
  AOI22_X1 U5938 ( .A1(\mem[275][7] ), .A2(n11750), .B1(n26855), .B2(
        data_in[7]), .ZN(n11757) );
  INV_X1 U5939 ( .A(n11758), .ZN(n23898) );
  AOI22_X1 U5940 ( .A1(\mem[276][0] ), .A2(n11759), .B1(n26854), .B2(
        data_in[0]), .ZN(n11758) );
  INV_X1 U5941 ( .A(n11760), .ZN(n23897) );
  AOI22_X1 U5942 ( .A1(\mem[276][1] ), .A2(n11759), .B1(n26854), .B2(
        data_in[1]), .ZN(n11760) );
  INV_X1 U5943 ( .A(n11761), .ZN(n23896) );
  AOI22_X1 U5944 ( .A1(\mem[276][2] ), .A2(n11759), .B1(n26854), .B2(
        data_in[2]), .ZN(n11761) );
  INV_X1 U5945 ( .A(n11762), .ZN(n23895) );
  AOI22_X1 U5946 ( .A1(\mem[276][3] ), .A2(n11759), .B1(n26854), .B2(
        data_in[3]), .ZN(n11762) );
  INV_X1 U5947 ( .A(n11763), .ZN(n23894) );
  AOI22_X1 U5948 ( .A1(\mem[276][4] ), .A2(n11759), .B1(n26854), .B2(
        data_in[4]), .ZN(n11763) );
  INV_X1 U5949 ( .A(n11764), .ZN(n23893) );
  AOI22_X1 U5950 ( .A1(\mem[276][5] ), .A2(n11759), .B1(n26854), .B2(
        data_in[5]), .ZN(n11764) );
  INV_X1 U5951 ( .A(n11765), .ZN(n23892) );
  AOI22_X1 U5952 ( .A1(\mem[276][6] ), .A2(n11759), .B1(n26854), .B2(
        data_in[6]), .ZN(n11765) );
  INV_X1 U5953 ( .A(n11766), .ZN(n23891) );
  AOI22_X1 U5954 ( .A1(\mem[276][7] ), .A2(n11759), .B1(n26854), .B2(
        data_in[7]), .ZN(n11766) );
  INV_X1 U5955 ( .A(n11767), .ZN(n23890) );
  AOI22_X1 U5956 ( .A1(\mem[277][0] ), .A2(n11768), .B1(n26853), .B2(
        data_in[0]), .ZN(n11767) );
  INV_X1 U5957 ( .A(n11769), .ZN(n23889) );
  AOI22_X1 U5958 ( .A1(\mem[277][1] ), .A2(n11768), .B1(n26853), .B2(
        data_in[1]), .ZN(n11769) );
  INV_X1 U5959 ( .A(n11770), .ZN(n23888) );
  AOI22_X1 U5960 ( .A1(\mem[277][2] ), .A2(n11768), .B1(n26853), .B2(
        data_in[2]), .ZN(n11770) );
  INV_X1 U5961 ( .A(n11771), .ZN(n23887) );
  AOI22_X1 U5962 ( .A1(\mem[277][3] ), .A2(n11768), .B1(n26853), .B2(
        data_in[3]), .ZN(n11771) );
  INV_X1 U5963 ( .A(n11772), .ZN(n23886) );
  AOI22_X1 U5964 ( .A1(\mem[277][4] ), .A2(n11768), .B1(n26853), .B2(
        data_in[4]), .ZN(n11772) );
  INV_X1 U5965 ( .A(n11773), .ZN(n23885) );
  AOI22_X1 U5966 ( .A1(\mem[277][5] ), .A2(n11768), .B1(n26853), .B2(
        data_in[5]), .ZN(n11773) );
  INV_X1 U5967 ( .A(n11774), .ZN(n23884) );
  AOI22_X1 U5968 ( .A1(\mem[277][6] ), .A2(n11768), .B1(n26853), .B2(
        data_in[6]), .ZN(n11774) );
  INV_X1 U5969 ( .A(n11775), .ZN(n23883) );
  AOI22_X1 U5970 ( .A1(\mem[277][7] ), .A2(n11768), .B1(n26853), .B2(
        data_in[7]), .ZN(n11775) );
  INV_X1 U5971 ( .A(n11776), .ZN(n23882) );
  AOI22_X1 U5972 ( .A1(\mem[278][0] ), .A2(n11777), .B1(n26852), .B2(
        data_in[0]), .ZN(n11776) );
  INV_X1 U5973 ( .A(n11778), .ZN(n23881) );
  AOI22_X1 U5974 ( .A1(\mem[278][1] ), .A2(n11777), .B1(n26852), .B2(
        data_in[1]), .ZN(n11778) );
  INV_X1 U5975 ( .A(n11779), .ZN(n23880) );
  AOI22_X1 U5976 ( .A1(\mem[278][2] ), .A2(n11777), .B1(n26852), .B2(
        data_in[2]), .ZN(n11779) );
  INV_X1 U5977 ( .A(n11780), .ZN(n23879) );
  AOI22_X1 U5978 ( .A1(\mem[278][3] ), .A2(n11777), .B1(n26852), .B2(
        data_in[3]), .ZN(n11780) );
  INV_X1 U5979 ( .A(n11781), .ZN(n23878) );
  AOI22_X1 U5980 ( .A1(\mem[278][4] ), .A2(n11777), .B1(n26852), .B2(
        data_in[4]), .ZN(n11781) );
  INV_X1 U5981 ( .A(n11782), .ZN(n23877) );
  AOI22_X1 U5982 ( .A1(\mem[278][5] ), .A2(n11777), .B1(n26852), .B2(
        data_in[5]), .ZN(n11782) );
  INV_X1 U5983 ( .A(n11783), .ZN(n23876) );
  AOI22_X1 U5984 ( .A1(\mem[278][6] ), .A2(n11777), .B1(n26852), .B2(
        data_in[6]), .ZN(n11783) );
  INV_X1 U5985 ( .A(n11784), .ZN(n23875) );
  AOI22_X1 U5986 ( .A1(\mem[278][7] ), .A2(n11777), .B1(n26852), .B2(
        data_in[7]), .ZN(n11784) );
  INV_X1 U5987 ( .A(n11785), .ZN(n23874) );
  AOI22_X1 U5988 ( .A1(\mem[279][0] ), .A2(n11786), .B1(n26851), .B2(
        data_in[0]), .ZN(n11785) );
  INV_X1 U5989 ( .A(n11787), .ZN(n23873) );
  AOI22_X1 U5990 ( .A1(\mem[279][1] ), .A2(n11786), .B1(n26851), .B2(
        data_in[1]), .ZN(n11787) );
  INV_X1 U5991 ( .A(n11788), .ZN(n23872) );
  AOI22_X1 U5992 ( .A1(\mem[279][2] ), .A2(n11786), .B1(n26851), .B2(
        data_in[2]), .ZN(n11788) );
  INV_X1 U5993 ( .A(n11789), .ZN(n23871) );
  AOI22_X1 U5994 ( .A1(\mem[279][3] ), .A2(n11786), .B1(n26851), .B2(
        data_in[3]), .ZN(n11789) );
  INV_X1 U5995 ( .A(n11790), .ZN(n23870) );
  AOI22_X1 U5996 ( .A1(\mem[279][4] ), .A2(n11786), .B1(n26851), .B2(
        data_in[4]), .ZN(n11790) );
  INV_X1 U5997 ( .A(n11791), .ZN(n23869) );
  AOI22_X1 U5998 ( .A1(\mem[279][5] ), .A2(n11786), .B1(n26851), .B2(
        data_in[5]), .ZN(n11791) );
  INV_X1 U5999 ( .A(n11792), .ZN(n23868) );
  AOI22_X1 U6000 ( .A1(\mem[279][6] ), .A2(n11786), .B1(n26851), .B2(
        data_in[6]), .ZN(n11792) );
  INV_X1 U6001 ( .A(n11793), .ZN(n23867) );
  AOI22_X1 U6002 ( .A1(\mem[279][7] ), .A2(n11786), .B1(n26851), .B2(
        data_in[7]), .ZN(n11793) );
  INV_X1 U6003 ( .A(n11794), .ZN(n23866) );
  AOI22_X1 U6004 ( .A1(\mem[280][0] ), .A2(n11795), .B1(n26850), .B2(
        data_in[0]), .ZN(n11794) );
  INV_X1 U6005 ( .A(n11796), .ZN(n23865) );
  AOI22_X1 U6006 ( .A1(\mem[280][1] ), .A2(n11795), .B1(n26850), .B2(
        data_in[1]), .ZN(n11796) );
  INV_X1 U6007 ( .A(n11797), .ZN(n23864) );
  AOI22_X1 U6008 ( .A1(\mem[280][2] ), .A2(n11795), .B1(n26850), .B2(
        data_in[2]), .ZN(n11797) );
  INV_X1 U6009 ( .A(n11798), .ZN(n23863) );
  AOI22_X1 U6010 ( .A1(\mem[280][3] ), .A2(n11795), .B1(n26850), .B2(
        data_in[3]), .ZN(n11798) );
  INV_X1 U6011 ( .A(n11799), .ZN(n23862) );
  AOI22_X1 U6012 ( .A1(\mem[280][4] ), .A2(n11795), .B1(n26850), .B2(
        data_in[4]), .ZN(n11799) );
  INV_X1 U6013 ( .A(n11800), .ZN(n23861) );
  AOI22_X1 U6014 ( .A1(\mem[280][5] ), .A2(n11795), .B1(n26850), .B2(
        data_in[5]), .ZN(n11800) );
  INV_X1 U6015 ( .A(n11801), .ZN(n23860) );
  AOI22_X1 U6016 ( .A1(\mem[280][6] ), .A2(n11795), .B1(n26850), .B2(
        data_in[6]), .ZN(n11801) );
  INV_X1 U6017 ( .A(n11802), .ZN(n23859) );
  AOI22_X1 U6018 ( .A1(\mem[280][7] ), .A2(n11795), .B1(n26850), .B2(
        data_in[7]), .ZN(n11802) );
  INV_X1 U6019 ( .A(n11803), .ZN(n23858) );
  AOI22_X1 U6020 ( .A1(\mem[281][0] ), .A2(n11804), .B1(n26849), .B2(
        data_in[0]), .ZN(n11803) );
  INV_X1 U6021 ( .A(n11805), .ZN(n23857) );
  AOI22_X1 U6022 ( .A1(\mem[281][1] ), .A2(n11804), .B1(n26849), .B2(
        data_in[1]), .ZN(n11805) );
  INV_X1 U6023 ( .A(n11806), .ZN(n23856) );
  AOI22_X1 U6024 ( .A1(\mem[281][2] ), .A2(n11804), .B1(n26849), .B2(
        data_in[2]), .ZN(n11806) );
  INV_X1 U6025 ( .A(n11807), .ZN(n23855) );
  AOI22_X1 U6026 ( .A1(\mem[281][3] ), .A2(n11804), .B1(n26849), .B2(
        data_in[3]), .ZN(n11807) );
  INV_X1 U6027 ( .A(n11808), .ZN(n23854) );
  AOI22_X1 U6028 ( .A1(\mem[281][4] ), .A2(n11804), .B1(n26849), .B2(
        data_in[4]), .ZN(n11808) );
  INV_X1 U6029 ( .A(n11809), .ZN(n23853) );
  AOI22_X1 U6030 ( .A1(\mem[281][5] ), .A2(n11804), .B1(n26849), .B2(
        data_in[5]), .ZN(n11809) );
  INV_X1 U6031 ( .A(n11810), .ZN(n23852) );
  AOI22_X1 U6032 ( .A1(\mem[281][6] ), .A2(n11804), .B1(n26849), .B2(
        data_in[6]), .ZN(n11810) );
  INV_X1 U6033 ( .A(n11811), .ZN(n23851) );
  AOI22_X1 U6034 ( .A1(\mem[281][7] ), .A2(n11804), .B1(n26849), .B2(
        data_in[7]), .ZN(n11811) );
  INV_X1 U6035 ( .A(n11812), .ZN(n23850) );
  AOI22_X1 U6036 ( .A1(\mem[282][0] ), .A2(n11813), .B1(n26848), .B2(
        data_in[0]), .ZN(n11812) );
  INV_X1 U6037 ( .A(n11814), .ZN(n23849) );
  AOI22_X1 U6038 ( .A1(\mem[282][1] ), .A2(n11813), .B1(n26848), .B2(
        data_in[1]), .ZN(n11814) );
  INV_X1 U6039 ( .A(n11815), .ZN(n23848) );
  AOI22_X1 U6040 ( .A1(\mem[282][2] ), .A2(n11813), .B1(n26848), .B2(
        data_in[2]), .ZN(n11815) );
  INV_X1 U6041 ( .A(n11816), .ZN(n23847) );
  AOI22_X1 U6042 ( .A1(\mem[282][3] ), .A2(n11813), .B1(n26848), .B2(
        data_in[3]), .ZN(n11816) );
  INV_X1 U6043 ( .A(n11817), .ZN(n23846) );
  AOI22_X1 U6044 ( .A1(\mem[282][4] ), .A2(n11813), .B1(n26848), .B2(
        data_in[4]), .ZN(n11817) );
  INV_X1 U6045 ( .A(n11818), .ZN(n23845) );
  AOI22_X1 U6046 ( .A1(\mem[282][5] ), .A2(n11813), .B1(n26848), .B2(
        data_in[5]), .ZN(n11818) );
  INV_X1 U6047 ( .A(n11819), .ZN(n23844) );
  AOI22_X1 U6048 ( .A1(\mem[282][6] ), .A2(n11813), .B1(n26848), .B2(
        data_in[6]), .ZN(n11819) );
  INV_X1 U6049 ( .A(n11820), .ZN(n23843) );
  AOI22_X1 U6050 ( .A1(\mem[282][7] ), .A2(n11813), .B1(n26848), .B2(
        data_in[7]), .ZN(n11820) );
  INV_X1 U6051 ( .A(n11821), .ZN(n23842) );
  AOI22_X1 U6052 ( .A1(\mem[283][0] ), .A2(n11822), .B1(n26847), .B2(
        data_in[0]), .ZN(n11821) );
  INV_X1 U6053 ( .A(n11823), .ZN(n23841) );
  AOI22_X1 U6054 ( .A1(\mem[283][1] ), .A2(n11822), .B1(n26847), .B2(
        data_in[1]), .ZN(n11823) );
  INV_X1 U6055 ( .A(n11824), .ZN(n23840) );
  AOI22_X1 U6056 ( .A1(\mem[283][2] ), .A2(n11822), .B1(n26847), .B2(
        data_in[2]), .ZN(n11824) );
  INV_X1 U6057 ( .A(n11825), .ZN(n23839) );
  AOI22_X1 U6058 ( .A1(\mem[283][3] ), .A2(n11822), .B1(n26847), .B2(
        data_in[3]), .ZN(n11825) );
  INV_X1 U6059 ( .A(n11826), .ZN(n23838) );
  AOI22_X1 U6060 ( .A1(\mem[283][4] ), .A2(n11822), .B1(n26847), .B2(
        data_in[4]), .ZN(n11826) );
  INV_X1 U6061 ( .A(n11827), .ZN(n23837) );
  AOI22_X1 U6062 ( .A1(\mem[283][5] ), .A2(n11822), .B1(n26847), .B2(
        data_in[5]), .ZN(n11827) );
  INV_X1 U6063 ( .A(n11828), .ZN(n23836) );
  AOI22_X1 U6064 ( .A1(\mem[283][6] ), .A2(n11822), .B1(n26847), .B2(
        data_in[6]), .ZN(n11828) );
  INV_X1 U6065 ( .A(n11829), .ZN(n23835) );
  AOI22_X1 U6066 ( .A1(\mem[283][7] ), .A2(n11822), .B1(n26847), .B2(
        data_in[7]), .ZN(n11829) );
  INV_X1 U6067 ( .A(n11830), .ZN(n23834) );
  AOI22_X1 U6068 ( .A1(\mem[284][0] ), .A2(n11831), .B1(n26846), .B2(
        data_in[0]), .ZN(n11830) );
  INV_X1 U6069 ( .A(n11832), .ZN(n23833) );
  AOI22_X1 U6070 ( .A1(\mem[284][1] ), .A2(n11831), .B1(n26846), .B2(
        data_in[1]), .ZN(n11832) );
  INV_X1 U6071 ( .A(n11833), .ZN(n23832) );
  AOI22_X1 U6072 ( .A1(\mem[284][2] ), .A2(n11831), .B1(n26846), .B2(
        data_in[2]), .ZN(n11833) );
  INV_X1 U6073 ( .A(n11834), .ZN(n23831) );
  AOI22_X1 U6074 ( .A1(\mem[284][3] ), .A2(n11831), .B1(n26846), .B2(
        data_in[3]), .ZN(n11834) );
  INV_X1 U6075 ( .A(n11835), .ZN(n23830) );
  AOI22_X1 U6076 ( .A1(\mem[284][4] ), .A2(n11831), .B1(n26846), .B2(
        data_in[4]), .ZN(n11835) );
  INV_X1 U6077 ( .A(n11836), .ZN(n23829) );
  AOI22_X1 U6078 ( .A1(\mem[284][5] ), .A2(n11831), .B1(n26846), .B2(
        data_in[5]), .ZN(n11836) );
  INV_X1 U6079 ( .A(n11837), .ZN(n23828) );
  AOI22_X1 U6080 ( .A1(\mem[284][6] ), .A2(n11831), .B1(n26846), .B2(
        data_in[6]), .ZN(n11837) );
  INV_X1 U6081 ( .A(n11838), .ZN(n23827) );
  AOI22_X1 U6082 ( .A1(\mem[284][7] ), .A2(n11831), .B1(n26846), .B2(
        data_in[7]), .ZN(n11838) );
  INV_X1 U6083 ( .A(n11839), .ZN(n23826) );
  AOI22_X1 U6084 ( .A1(\mem[285][0] ), .A2(n11840), .B1(n26845), .B2(
        data_in[0]), .ZN(n11839) );
  INV_X1 U6085 ( .A(n11841), .ZN(n23825) );
  AOI22_X1 U6086 ( .A1(\mem[285][1] ), .A2(n11840), .B1(n26845), .B2(
        data_in[1]), .ZN(n11841) );
  INV_X1 U6087 ( .A(n11842), .ZN(n23824) );
  AOI22_X1 U6088 ( .A1(\mem[285][2] ), .A2(n11840), .B1(n26845), .B2(
        data_in[2]), .ZN(n11842) );
  INV_X1 U6089 ( .A(n11843), .ZN(n23823) );
  AOI22_X1 U6090 ( .A1(\mem[285][3] ), .A2(n11840), .B1(n26845), .B2(
        data_in[3]), .ZN(n11843) );
  INV_X1 U6091 ( .A(n11844), .ZN(n23822) );
  AOI22_X1 U6092 ( .A1(\mem[285][4] ), .A2(n11840), .B1(n26845), .B2(
        data_in[4]), .ZN(n11844) );
  INV_X1 U6093 ( .A(n11845), .ZN(n23821) );
  AOI22_X1 U6094 ( .A1(\mem[285][5] ), .A2(n11840), .B1(n26845), .B2(
        data_in[5]), .ZN(n11845) );
  INV_X1 U6095 ( .A(n11846), .ZN(n23820) );
  AOI22_X1 U6096 ( .A1(\mem[285][6] ), .A2(n11840), .B1(n26845), .B2(
        data_in[6]), .ZN(n11846) );
  INV_X1 U6097 ( .A(n11847), .ZN(n23819) );
  AOI22_X1 U6098 ( .A1(\mem[285][7] ), .A2(n11840), .B1(n26845), .B2(
        data_in[7]), .ZN(n11847) );
  INV_X1 U6099 ( .A(n11848), .ZN(n23818) );
  AOI22_X1 U6100 ( .A1(\mem[286][0] ), .A2(n11849), .B1(n26844), .B2(
        data_in[0]), .ZN(n11848) );
  INV_X1 U6101 ( .A(n11850), .ZN(n23817) );
  AOI22_X1 U6102 ( .A1(\mem[286][1] ), .A2(n11849), .B1(n26844), .B2(
        data_in[1]), .ZN(n11850) );
  INV_X1 U6103 ( .A(n11851), .ZN(n23816) );
  AOI22_X1 U6104 ( .A1(\mem[286][2] ), .A2(n11849), .B1(n26844), .B2(
        data_in[2]), .ZN(n11851) );
  INV_X1 U6105 ( .A(n11852), .ZN(n23815) );
  AOI22_X1 U6106 ( .A1(\mem[286][3] ), .A2(n11849), .B1(n26844), .B2(
        data_in[3]), .ZN(n11852) );
  INV_X1 U6107 ( .A(n11853), .ZN(n23814) );
  AOI22_X1 U6108 ( .A1(\mem[286][4] ), .A2(n11849), .B1(n26844), .B2(
        data_in[4]), .ZN(n11853) );
  INV_X1 U6109 ( .A(n11854), .ZN(n23813) );
  AOI22_X1 U6110 ( .A1(\mem[286][5] ), .A2(n11849), .B1(n26844), .B2(
        data_in[5]), .ZN(n11854) );
  INV_X1 U6111 ( .A(n11855), .ZN(n23812) );
  AOI22_X1 U6112 ( .A1(\mem[286][6] ), .A2(n11849), .B1(n26844), .B2(
        data_in[6]), .ZN(n11855) );
  INV_X1 U6113 ( .A(n11856), .ZN(n23811) );
  AOI22_X1 U6114 ( .A1(\mem[286][7] ), .A2(n11849), .B1(n26844), .B2(
        data_in[7]), .ZN(n11856) );
  INV_X1 U6115 ( .A(n11857), .ZN(n23810) );
  AOI22_X1 U6116 ( .A1(\mem[287][0] ), .A2(n11858), .B1(n26843), .B2(
        data_in[0]), .ZN(n11857) );
  INV_X1 U6117 ( .A(n11859), .ZN(n23809) );
  AOI22_X1 U6118 ( .A1(\mem[287][1] ), .A2(n11858), .B1(n26843), .B2(
        data_in[1]), .ZN(n11859) );
  INV_X1 U6119 ( .A(n11860), .ZN(n23808) );
  AOI22_X1 U6120 ( .A1(\mem[287][2] ), .A2(n11858), .B1(n26843), .B2(
        data_in[2]), .ZN(n11860) );
  INV_X1 U6121 ( .A(n11861), .ZN(n23807) );
  AOI22_X1 U6122 ( .A1(\mem[287][3] ), .A2(n11858), .B1(n26843), .B2(
        data_in[3]), .ZN(n11861) );
  INV_X1 U6123 ( .A(n11862), .ZN(n23806) );
  AOI22_X1 U6124 ( .A1(\mem[287][4] ), .A2(n11858), .B1(n26843), .B2(
        data_in[4]), .ZN(n11862) );
  INV_X1 U6125 ( .A(n11863), .ZN(n23805) );
  AOI22_X1 U6126 ( .A1(\mem[287][5] ), .A2(n11858), .B1(n26843), .B2(
        data_in[5]), .ZN(n11863) );
  INV_X1 U6127 ( .A(n11864), .ZN(n23804) );
  AOI22_X1 U6128 ( .A1(\mem[287][6] ), .A2(n11858), .B1(n26843), .B2(
        data_in[6]), .ZN(n11864) );
  INV_X1 U6129 ( .A(n11865), .ZN(n23803) );
  AOI22_X1 U6130 ( .A1(\mem[287][7] ), .A2(n11858), .B1(n26843), .B2(
        data_in[7]), .ZN(n11865) );
  INV_X1 U6131 ( .A(n11940), .ZN(n23738) );
  AOI22_X1 U6132 ( .A1(\mem[296][0] ), .A2(n11941), .B1(n26834), .B2(
        data_in[0]), .ZN(n11940) );
  INV_X1 U6133 ( .A(n11942), .ZN(n23737) );
  AOI22_X1 U6134 ( .A1(\mem[296][1] ), .A2(n11941), .B1(n26834), .B2(
        data_in[1]), .ZN(n11942) );
  INV_X1 U6135 ( .A(n11943), .ZN(n23736) );
  AOI22_X1 U6136 ( .A1(\mem[296][2] ), .A2(n11941), .B1(n26834), .B2(
        data_in[2]), .ZN(n11943) );
  INV_X1 U6137 ( .A(n11944), .ZN(n23735) );
  AOI22_X1 U6138 ( .A1(\mem[296][3] ), .A2(n11941), .B1(n26834), .B2(
        data_in[3]), .ZN(n11944) );
  INV_X1 U6139 ( .A(n11945), .ZN(n23734) );
  AOI22_X1 U6140 ( .A1(\mem[296][4] ), .A2(n11941), .B1(n26834), .B2(
        data_in[4]), .ZN(n11945) );
  INV_X1 U6141 ( .A(n11946), .ZN(n23733) );
  AOI22_X1 U6142 ( .A1(\mem[296][5] ), .A2(n11941), .B1(n26834), .B2(
        data_in[5]), .ZN(n11946) );
  INV_X1 U6143 ( .A(n11947), .ZN(n23732) );
  AOI22_X1 U6144 ( .A1(\mem[296][6] ), .A2(n11941), .B1(n26834), .B2(
        data_in[6]), .ZN(n11947) );
  INV_X1 U6145 ( .A(n11948), .ZN(n23731) );
  AOI22_X1 U6146 ( .A1(\mem[296][7] ), .A2(n11941), .B1(n26834), .B2(
        data_in[7]), .ZN(n11948) );
  INV_X1 U6147 ( .A(n11949), .ZN(n23730) );
  AOI22_X1 U6148 ( .A1(\mem[297][0] ), .A2(n11950), .B1(n26833), .B2(
        data_in[0]), .ZN(n11949) );
  INV_X1 U6149 ( .A(n11951), .ZN(n23729) );
  AOI22_X1 U6150 ( .A1(\mem[297][1] ), .A2(n11950), .B1(n26833), .B2(
        data_in[1]), .ZN(n11951) );
  INV_X1 U6151 ( .A(n11952), .ZN(n23728) );
  AOI22_X1 U6152 ( .A1(\mem[297][2] ), .A2(n11950), .B1(n26833), .B2(
        data_in[2]), .ZN(n11952) );
  INV_X1 U6153 ( .A(n11953), .ZN(n23727) );
  AOI22_X1 U6154 ( .A1(\mem[297][3] ), .A2(n11950), .B1(n26833), .B2(
        data_in[3]), .ZN(n11953) );
  INV_X1 U6155 ( .A(n11954), .ZN(n23726) );
  AOI22_X1 U6156 ( .A1(\mem[297][4] ), .A2(n11950), .B1(n26833), .B2(
        data_in[4]), .ZN(n11954) );
  INV_X1 U6157 ( .A(n11955), .ZN(n23725) );
  AOI22_X1 U6158 ( .A1(\mem[297][5] ), .A2(n11950), .B1(n26833), .B2(
        data_in[5]), .ZN(n11955) );
  INV_X1 U6159 ( .A(n11956), .ZN(n23724) );
  AOI22_X1 U6160 ( .A1(\mem[297][6] ), .A2(n11950), .B1(n26833), .B2(
        data_in[6]), .ZN(n11956) );
  INV_X1 U6161 ( .A(n11957), .ZN(n23723) );
  AOI22_X1 U6162 ( .A1(\mem[297][7] ), .A2(n11950), .B1(n26833), .B2(
        data_in[7]), .ZN(n11957) );
  INV_X1 U6163 ( .A(n11958), .ZN(n23722) );
  AOI22_X1 U6164 ( .A1(\mem[298][0] ), .A2(n11959), .B1(n26832), .B2(
        data_in[0]), .ZN(n11958) );
  INV_X1 U6165 ( .A(n11960), .ZN(n23721) );
  AOI22_X1 U6166 ( .A1(\mem[298][1] ), .A2(n11959), .B1(n26832), .B2(
        data_in[1]), .ZN(n11960) );
  INV_X1 U6167 ( .A(n11961), .ZN(n23720) );
  AOI22_X1 U6168 ( .A1(\mem[298][2] ), .A2(n11959), .B1(n26832), .B2(
        data_in[2]), .ZN(n11961) );
  INV_X1 U6169 ( .A(n11962), .ZN(n23719) );
  AOI22_X1 U6170 ( .A1(\mem[298][3] ), .A2(n11959), .B1(n26832), .B2(
        data_in[3]), .ZN(n11962) );
  INV_X1 U6171 ( .A(n11963), .ZN(n23718) );
  AOI22_X1 U6172 ( .A1(\mem[298][4] ), .A2(n11959), .B1(n26832), .B2(
        data_in[4]), .ZN(n11963) );
  INV_X1 U6173 ( .A(n11964), .ZN(n23717) );
  AOI22_X1 U6174 ( .A1(\mem[298][5] ), .A2(n11959), .B1(n26832), .B2(
        data_in[5]), .ZN(n11964) );
  INV_X1 U6175 ( .A(n11965), .ZN(n23716) );
  AOI22_X1 U6176 ( .A1(\mem[298][6] ), .A2(n11959), .B1(n26832), .B2(
        data_in[6]), .ZN(n11965) );
  INV_X1 U6177 ( .A(n11966), .ZN(n23715) );
  AOI22_X1 U6178 ( .A1(\mem[298][7] ), .A2(n11959), .B1(n26832), .B2(
        data_in[7]), .ZN(n11966) );
  INV_X1 U6179 ( .A(n11967), .ZN(n23714) );
  AOI22_X1 U6180 ( .A1(\mem[299][0] ), .A2(n11968), .B1(n26831), .B2(
        data_in[0]), .ZN(n11967) );
  INV_X1 U6181 ( .A(n11969), .ZN(n23713) );
  AOI22_X1 U6182 ( .A1(\mem[299][1] ), .A2(n11968), .B1(n26831), .B2(
        data_in[1]), .ZN(n11969) );
  INV_X1 U6183 ( .A(n11970), .ZN(n23712) );
  AOI22_X1 U6184 ( .A1(\mem[299][2] ), .A2(n11968), .B1(n26831), .B2(
        data_in[2]), .ZN(n11970) );
  INV_X1 U6185 ( .A(n11971), .ZN(n23711) );
  AOI22_X1 U6186 ( .A1(\mem[299][3] ), .A2(n11968), .B1(n26831), .B2(
        data_in[3]), .ZN(n11971) );
  INV_X1 U6187 ( .A(n11972), .ZN(n23710) );
  AOI22_X1 U6188 ( .A1(\mem[299][4] ), .A2(n11968), .B1(n26831), .B2(
        data_in[4]), .ZN(n11972) );
  INV_X1 U6189 ( .A(n11973), .ZN(n23709) );
  AOI22_X1 U6190 ( .A1(\mem[299][5] ), .A2(n11968), .B1(n26831), .B2(
        data_in[5]), .ZN(n11973) );
  INV_X1 U6191 ( .A(n11974), .ZN(n23708) );
  AOI22_X1 U6192 ( .A1(\mem[299][6] ), .A2(n11968), .B1(n26831), .B2(
        data_in[6]), .ZN(n11974) );
  INV_X1 U6193 ( .A(n11975), .ZN(n23707) );
  AOI22_X1 U6194 ( .A1(\mem[299][7] ), .A2(n11968), .B1(n26831), .B2(
        data_in[7]), .ZN(n11975) );
  INV_X1 U6195 ( .A(n11976), .ZN(n23706) );
  AOI22_X1 U6196 ( .A1(\mem[300][0] ), .A2(n11977), .B1(n26830), .B2(
        data_in[0]), .ZN(n11976) );
  INV_X1 U6197 ( .A(n11978), .ZN(n23705) );
  AOI22_X1 U6198 ( .A1(\mem[300][1] ), .A2(n11977), .B1(n26830), .B2(
        data_in[1]), .ZN(n11978) );
  INV_X1 U6199 ( .A(n11979), .ZN(n23704) );
  AOI22_X1 U6200 ( .A1(\mem[300][2] ), .A2(n11977), .B1(n26830), .B2(
        data_in[2]), .ZN(n11979) );
  INV_X1 U6201 ( .A(n11980), .ZN(n23703) );
  AOI22_X1 U6202 ( .A1(\mem[300][3] ), .A2(n11977), .B1(n26830), .B2(
        data_in[3]), .ZN(n11980) );
  INV_X1 U6203 ( .A(n11981), .ZN(n23702) );
  AOI22_X1 U6204 ( .A1(\mem[300][4] ), .A2(n11977), .B1(n26830), .B2(
        data_in[4]), .ZN(n11981) );
  INV_X1 U6205 ( .A(n11982), .ZN(n23701) );
  AOI22_X1 U6206 ( .A1(\mem[300][5] ), .A2(n11977), .B1(n26830), .B2(
        data_in[5]), .ZN(n11982) );
  INV_X1 U6207 ( .A(n11983), .ZN(n23700) );
  AOI22_X1 U6208 ( .A1(\mem[300][6] ), .A2(n11977), .B1(n26830), .B2(
        data_in[6]), .ZN(n11983) );
  INV_X1 U6209 ( .A(n11984), .ZN(n23699) );
  AOI22_X1 U6210 ( .A1(\mem[300][7] ), .A2(n11977), .B1(n26830), .B2(
        data_in[7]), .ZN(n11984) );
  INV_X1 U6211 ( .A(n11985), .ZN(n23698) );
  AOI22_X1 U6212 ( .A1(\mem[301][0] ), .A2(n11986), .B1(n26829), .B2(
        data_in[0]), .ZN(n11985) );
  INV_X1 U6213 ( .A(n11987), .ZN(n23697) );
  AOI22_X1 U6214 ( .A1(\mem[301][1] ), .A2(n11986), .B1(n26829), .B2(
        data_in[1]), .ZN(n11987) );
  INV_X1 U6215 ( .A(n11988), .ZN(n23696) );
  AOI22_X1 U6216 ( .A1(\mem[301][2] ), .A2(n11986), .B1(n26829), .B2(
        data_in[2]), .ZN(n11988) );
  INV_X1 U6217 ( .A(n11989), .ZN(n23695) );
  AOI22_X1 U6218 ( .A1(\mem[301][3] ), .A2(n11986), .B1(n26829), .B2(
        data_in[3]), .ZN(n11989) );
  INV_X1 U6219 ( .A(n11990), .ZN(n23694) );
  AOI22_X1 U6220 ( .A1(\mem[301][4] ), .A2(n11986), .B1(n26829), .B2(
        data_in[4]), .ZN(n11990) );
  INV_X1 U6221 ( .A(n11991), .ZN(n23693) );
  AOI22_X1 U6222 ( .A1(\mem[301][5] ), .A2(n11986), .B1(n26829), .B2(
        data_in[5]), .ZN(n11991) );
  INV_X1 U6223 ( .A(n11992), .ZN(n23692) );
  AOI22_X1 U6224 ( .A1(\mem[301][6] ), .A2(n11986), .B1(n26829), .B2(
        data_in[6]), .ZN(n11992) );
  INV_X1 U6225 ( .A(n11993), .ZN(n23691) );
  AOI22_X1 U6226 ( .A1(\mem[301][7] ), .A2(n11986), .B1(n26829), .B2(
        data_in[7]), .ZN(n11993) );
  INV_X1 U6227 ( .A(n11994), .ZN(n23690) );
  AOI22_X1 U6228 ( .A1(\mem[302][0] ), .A2(n11995), .B1(n26828), .B2(
        data_in[0]), .ZN(n11994) );
  INV_X1 U6229 ( .A(n11996), .ZN(n23689) );
  AOI22_X1 U6230 ( .A1(\mem[302][1] ), .A2(n11995), .B1(n26828), .B2(
        data_in[1]), .ZN(n11996) );
  INV_X1 U6231 ( .A(n11997), .ZN(n23688) );
  AOI22_X1 U6232 ( .A1(\mem[302][2] ), .A2(n11995), .B1(n26828), .B2(
        data_in[2]), .ZN(n11997) );
  INV_X1 U6233 ( .A(n11998), .ZN(n23687) );
  AOI22_X1 U6234 ( .A1(\mem[302][3] ), .A2(n11995), .B1(n26828), .B2(
        data_in[3]), .ZN(n11998) );
  INV_X1 U6235 ( .A(n11999), .ZN(n23686) );
  AOI22_X1 U6236 ( .A1(\mem[302][4] ), .A2(n11995), .B1(n26828), .B2(
        data_in[4]), .ZN(n11999) );
  INV_X1 U6237 ( .A(n12000), .ZN(n23685) );
  AOI22_X1 U6238 ( .A1(\mem[302][5] ), .A2(n11995), .B1(n26828), .B2(
        data_in[5]), .ZN(n12000) );
  INV_X1 U6239 ( .A(n12001), .ZN(n23684) );
  AOI22_X1 U6240 ( .A1(\mem[302][6] ), .A2(n11995), .B1(n26828), .B2(
        data_in[6]), .ZN(n12001) );
  INV_X1 U6241 ( .A(n12002), .ZN(n23683) );
  AOI22_X1 U6242 ( .A1(\mem[302][7] ), .A2(n11995), .B1(n26828), .B2(
        data_in[7]), .ZN(n12002) );
  INV_X1 U6243 ( .A(n12003), .ZN(n23682) );
  AOI22_X1 U6244 ( .A1(\mem[303][0] ), .A2(n12004), .B1(n26827), .B2(
        data_in[0]), .ZN(n12003) );
  INV_X1 U6245 ( .A(n12005), .ZN(n23681) );
  AOI22_X1 U6246 ( .A1(\mem[303][1] ), .A2(n12004), .B1(n26827), .B2(
        data_in[1]), .ZN(n12005) );
  INV_X1 U6247 ( .A(n12006), .ZN(n23680) );
  AOI22_X1 U6248 ( .A1(\mem[303][2] ), .A2(n12004), .B1(n26827), .B2(
        data_in[2]), .ZN(n12006) );
  INV_X1 U6249 ( .A(n12007), .ZN(n23679) );
  AOI22_X1 U6250 ( .A1(\mem[303][3] ), .A2(n12004), .B1(n26827), .B2(
        data_in[3]), .ZN(n12007) );
  INV_X1 U6251 ( .A(n12008), .ZN(n23678) );
  AOI22_X1 U6252 ( .A1(\mem[303][4] ), .A2(n12004), .B1(n26827), .B2(
        data_in[4]), .ZN(n12008) );
  INV_X1 U6253 ( .A(n12009), .ZN(n23677) );
  AOI22_X1 U6254 ( .A1(\mem[303][5] ), .A2(n12004), .B1(n26827), .B2(
        data_in[5]), .ZN(n12009) );
  INV_X1 U6255 ( .A(n12010), .ZN(n23676) );
  AOI22_X1 U6256 ( .A1(\mem[303][6] ), .A2(n12004), .B1(n26827), .B2(
        data_in[6]), .ZN(n12010) );
  INV_X1 U6257 ( .A(n12011), .ZN(n23675) );
  AOI22_X1 U6258 ( .A1(\mem[303][7] ), .A2(n12004), .B1(n26827), .B2(
        data_in[7]), .ZN(n12011) );
  INV_X1 U6259 ( .A(n12012), .ZN(n23674) );
  AOI22_X1 U6260 ( .A1(\mem[304][0] ), .A2(n12013), .B1(n26826), .B2(
        data_in[0]), .ZN(n12012) );
  INV_X1 U6261 ( .A(n12014), .ZN(n23673) );
  AOI22_X1 U6262 ( .A1(\mem[304][1] ), .A2(n12013), .B1(n26826), .B2(
        data_in[1]), .ZN(n12014) );
  INV_X1 U6263 ( .A(n12015), .ZN(n23672) );
  AOI22_X1 U6264 ( .A1(\mem[304][2] ), .A2(n12013), .B1(n26826), .B2(
        data_in[2]), .ZN(n12015) );
  INV_X1 U6265 ( .A(n12016), .ZN(n23671) );
  AOI22_X1 U6266 ( .A1(\mem[304][3] ), .A2(n12013), .B1(n26826), .B2(
        data_in[3]), .ZN(n12016) );
  INV_X1 U6267 ( .A(n12017), .ZN(n23670) );
  AOI22_X1 U6268 ( .A1(\mem[304][4] ), .A2(n12013), .B1(n26826), .B2(
        data_in[4]), .ZN(n12017) );
  INV_X1 U6269 ( .A(n12018), .ZN(n23669) );
  AOI22_X1 U6270 ( .A1(\mem[304][5] ), .A2(n12013), .B1(n26826), .B2(
        data_in[5]), .ZN(n12018) );
  INV_X1 U6271 ( .A(n12019), .ZN(n23668) );
  AOI22_X1 U6272 ( .A1(\mem[304][6] ), .A2(n12013), .B1(n26826), .B2(
        data_in[6]), .ZN(n12019) );
  INV_X1 U6273 ( .A(n12020), .ZN(n23667) );
  AOI22_X1 U6274 ( .A1(\mem[304][7] ), .A2(n12013), .B1(n26826), .B2(
        data_in[7]), .ZN(n12020) );
  INV_X1 U6275 ( .A(n12021), .ZN(n23666) );
  AOI22_X1 U6276 ( .A1(\mem[305][0] ), .A2(n12022), .B1(n26825), .B2(
        data_in[0]), .ZN(n12021) );
  INV_X1 U6277 ( .A(n12023), .ZN(n23665) );
  AOI22_X1 U6278 ( .A1(\mem[305][1] ), .A2(n12022), .B1(n26825), .B2(
        data_in[1]), .ZN(n12023) );
  INV_X1 U6279 ( .A(n12024), .ZN(n23664) );
  AOI22_X1 U6280 ( .A1(\mem[305][2] ), .A2(n12022), .B1(n26825), .B2(
        data_in[2]), .ZN(n12024) );
  INV_X1 U6281 ( .A(n12025), .ZN(n23663) );
  AOI22_X1 U6282 ( .A1(\mem[305][3] ), .A2(n12022), .B1(n26825), .B2(
        data_in[3]), .ZN(n12025) );
  INV_X1 U6283 ( .A(n12026), .ZN(n23662) );
  AOI22_X1 U6284 ( .A1(\mem[305][4] ), .A2(n12022), .B1(n26825), .B2(
        data_in[4]), .ZN(n12026) );
  INV_X1 U6285 ( .A(n12027), .ZN(n23661) );
  AOI22_X1 U6286 ( .A1(\mem[305][5] ), .A2(n12022), .B1(n26825), .B2(
        data_in[5]), .ZN(n12027) );
  INV_X1 U6287 ( .A(n12028), .ZN(n23660) );
  AOI22_X1 U6288 ( .A1(\mem[305][6] ), .A2(n12022), .B1(n26825), .B2(
        data_in[6]), .ZN(n12028) );
  INV_X1 U6289 ( .A(n12029), .ZN(n23659) );
  AOI22_X1 U6290 ( .A1(\mem[305][7] ), .A2(n12022), .B1(n26825), .B2(
        data_in[7]), .ZN(n12029) );
  INV_X1 U6291 ( .A(n12030), .ZN(n23658) );
  AOI22_X1 U6292 ( .A1(\mem[306][0] ), .A2(n12031), .B1(n26824), .B2(
        data_in[0]), .ZN(n12030) );
  INV_X1 U6293 ( .A(n12032), .ZN(n23657) );
  AOI22_X1 U6294 ( .A1(\mem[306][1] ), .A2(n12031), .B1(n26824), .B2(
        data_in[1]), .ZN(n12032) );
  INV_X1 U6295 ( .A(n12033), .ZN(n23656) );
  AOI22_X1 U6296 ( .A1(\mem[306][2] ), .A2(n12031), .B1(n26824), .B2(
        data_in[2]), .ZN(n12033) );
  INV_X1 U6297 ( .A(n12034), .ZN(n23655) );
  AOI22_X1 U6298 ( .A1(\mem[306][3] ), .A2(n12031), .B1(n26824), .B2(
        data_in[3]), .ZN(n12034) );
  INV_X1 U6299 ( .A(n12035), .ZN(n23654) );
  AOI22_X1 U6300 ( .A1(\mem[306][4] ), .A2(n12031), .B1(n26824), .B2(
        data_in[4]), .ZN(n12035) );
  INV_X1 U6301 ( .A(n12036), .ZN(n23653) );
  AOI22_X1 U6302 ( .A1(\mem[306][5] ), .A2(n12031), .B1(n26824), .B2(
        data_in[5]), .ZN(n12036) );
  INV_X1 U6303 ( .A(n12037), .ZN(n23652) );
  AOI22_X1 U6304 ( .A1(\mem[306][6] ), .A2(n12031), .B1(n26824), .B2(
        data_in[6]), .ZN(n12037) );
  INV_X1 U6305 ( .A(n12038), .ZN(n23651) );
  AOI22_X1 U6306 ( .A1(\mem[306][7] ), .A2(n12031), .B1(n26824), .B2(
        data_in[7]), .ZN(n12038) );
  INV_X1 U6307 ( .A(n12039), .ZN(n23650) );
  AOI22_X1 U6308 ( .A1(\mem[307][0] ), .A2(n12040), .B1(n26823), .B2(
        data_in[0]), .ZN(n12039) );
  INV_X1 U6309 ( .A(n12041), .ZN(n23649) );
  AOI22_X1 U6310 ( .A1(\mem[307][1] ), .A2(n12040), .B1(n26823), .B2(
        data_in[1]), .ZN(n12041) );
  INV_X1 U6311 ( .A(n12042), .ZN(n23648) );
  AOI22_X1 U6312 ( .A1(\mem[307][2] ), .A2(n12040), .B1(n26823), .B2(
        data_in[2]), .ZN(n12042) );
  INV_X1 U6313 ( .A(n12043), .ZN(n23647) );
  AOI22_X1 U6314 ( .A1(\mem[307][3] ), .A2(n12040), .B1(n26823), .B2(
        data_in[3]), .ZN(n12043) );
  INV_X1 U6315 ( .A(n12044), .ZN(n23646) );
  AOI22_X1 U6316 ( .A1(\mem[307][4] ), .A2(n12040), .B1(n26823), .B2(
        data_in[4]), .ZN(n12044) );
  INV_X1 U6317 ( .A(n12045), .ZN(n23645) );
  AOI22_X1 U6318 ( .A1(\mem[307][5] ), .A2(n12040), .B1(n26823), .B2(
        data_in[5]), .ZN(n12045) );
  INV_X1 U6319 ( .A(n12046), .ZN(n23644) );
  AOI22_X1 U6320 ( .A1(\mem[307][6] ), .A2(n12040), .B1(n26823), .B2(
        data_in[6]), .ZN(n12046) );
  INV_X1 U6321 ( .A(n12047), .ZN(n23643) );
  AOI22_X1 U6322 ( .A1(\mem[307][7] ), .A2(n12040), .B1(n26823), .B2(
        data_in[7]), .ZN(n12047) );
  INV_X1 U6323 ( .A(n12048), .ZN(n23642) );
  AOI22_X1 U6324 ( .A1(\mem[308][0] ), .A2(n12049), .B1(n26822), .B2(
        data_in[0]), .ZN(n12048) );
  INV_X1 U6325 ( .A(n12050), .ZN(n23641) );
  AOI22_X1 U6326 ( .A1(\mem[308][1] ), .A2(n12049), .B1(n26822), .B2(
        data_in[1]), .ZN(n12050) );
  INV_X1 U6327 ( .A(n12051), .ZN(n23640) );
  AOI22_X1 U6328 ( .A1(\mem[308][2] ), .A2(n12049), .B1(n26822), .B2(
        data_in[2]), .ZN(n12051) );
  INV_X1 U6329 ( .A(n12052), .ZN(n23639) );
  AOI22_X1 U6330 ( .A1(\mem[308][3] ), .A2(n12049), .B1(n26822), .B2(
        data_in[3]), .ZN(n12052) );
  INV_X1 U6331 ( .A(n12053), .ZN(n23638) );
  AOI22_X1 U6332 ( .A1(\mem[308][4] ), .A2(n12049), .B1(n26822), .B2(
        data_in[4]), .ZN(n12053) );
  INV_X1 U6333 ( .A(n12054), .ZN(n23637) );
  AOI22_X1 U6334 ( .A1(\mem[308][5] ), .A2(n12049), .B1(n26822), .B2(
        data_in[5]), .ZN(n12054) );
  INV_X1 U6335 ( .A(n12055), .ZN(n23636) );
  AOI22_X1 U6336 ( .A1(\mem[308][6] ), .A2(n12049), .B1(n26822), .B2(
        data_in[6]), .ZN(n12055) );
  INV_X1 U6337 ( .A(n12056), .ZN(n23635) );
  AOI22_X1 U6338 ( .A1(\mem[308][7] ), .A2(n12049), .B1(n26822), .B2(
        data_in[7]), .ZN(n12056) );
  INV_X1 U6339 ( .A(n12057), .ZN(n23634) );
  AOI22_X1 U6340 ( .A1(\mem[309][0] ), .A2(n12058), .B1(n26821), .B2(
        data_in[0]), .ZN(n12057) );
  INV_X1 U6341 ( .A(n12059), .ZN(n23633) );
  AOI22_X1 U6342 ( .A1(\mem[309][1] ), .A2(n12058), .B1(n26821), .B2(
        data_in[1]), .ZN(n12059) );
  INV_X1 U6343 ( .A(n12060), .ZN(n23632) );
  AOI22_X1 U6344 ( .A1(\mem[309][2] ), .A2(n12058), .B1(n26821), .B2(
        data_in[2]), .ZN(n12060) );
  INV_X1 U6345 ( .A(n12061), .ZN(n23631) );
  AOI22_X1 U6346 ( .A1(\mem[309][3] ), .A2(n12058), .B1(n26821), .B2(
        data_in[3]), .ZN(n12061) );
  INV_X1 U6347 ( .A(n12062), .ZN(n23630) );
  AOI22_X1 U6348 ( .A1(\mem[309][4] ), .A2(n12058), .B1(n26821), .B2(
        data_in[4]), .ZN(n12062) );
  INV_X1 U6349 ( .A(n12063), .ZN(n23629) );
  AOI22_X1 U6350 ( .A1(\mem[309][5] ), .A2(n12058), .B1(n26821), .B2(
        data_in[5]), .ZN(n12063) );
  INV_X1 U6351 ( .A(n12064), .ZN(n23628) );
  AOI22_X1 U6352 ( .A1(\mem[309][6] ), .A2(n12058), .B1(n26821), .B2(
        data_in[6]), .ZN(n12064) );
  INV_X1 U6353 ( .A(n12065), .ZN(n23627) );
  AOI22_X1 U6354 ( .A1(\mem[309][7] ), .A2(n12058), .B1(n26821), .B2(
        data_in[7]), .ZN(n12065) );
  INV_X1 U6355 ( .A(n12066), .ZN(n23626) );
  AOI22_X1 U6356 ( .A1(\mem[310][0] ), .A2(n12067), .B1(n26820), .B2(
        data_in[0]), .ZN(n12066) );
  INV_X1 U6357 ( .A(n12068), .ZN(n23625) );
  AOI22_X1 U6358 ( .A1(\mem[310][1] ), .A2(n12067), .B1(n26820), .B2(
        data_in[1]), .ZN(n12068) );
  INV_X1 U6359 ( .A(n12069), .ZN(n23624) );
  AOI22_X1 U6360 ( .A1(\mem[310][2] ), .A2(n12067), .B1(n26820), .B2(
        data_in[2]), .ZN(n12069) );
  INV_X1 U6361 ( .A(n12070), .ZN(n23623) );
  AOI22_X1 U6362 ( .A1(\mem[310][3] ), .A2(n12067), .B1(n26820), .B2(
        data_in[3]), .ZN(n12070) );
  INV_X1 U6363 ( .A(n12071), .ZN(n23622) );
  AOI22_X1 U6364 ( .A1(\mem[310][4] ), .A2(n12067), .B1(n26820), .B2(
        data_in[4]), .ZN(n12071) );
  INV_X1 U6365 ( .A(n12072), .ZN(n23621) );
  AOI22_X1 U6366 ( .A1(\mem[310][5] ), .A2(n12067), .B1(n26820), .B2(
        data_in[5]), .ZN(n12072) );
  INV_X1 U6367 ( .A(n12073), .ZN(n23620) );
  AOI22_X1 U6368 ( .A1(\mem[310][6] ), .A2(n12067), .B1(n26820), .B2(
        data_in[6]), .ZN(n12073) );
  INV_X1 U6369 ( .A(n12074), .ZN(n23619) );
  AOI22_X1 U6370 ( .A1(\mem[310][7] ), .A2(n12067), .B1(n26820), .B2(
        data_in[7]), .ZN(n12074) );
  INV_X1 U6371 ( .A(n12075), .ZN(n23618) );
  AOI22_X1 U6372 ( .A1(\mem[311][0] ), .A2(n12076), .B1(n26819), .B2(
        data_in[0]), .ZN(n12075) );
  INV_X1 U6373 ( .A(n12077), .ZN(n23617) );
  AOI22_X1 U6374 ( .A1(\mem[311][1] ), .A2(n12076), .B1(n26819), .B2(
        data_in[1]), .ZN(n12077) );
  INV_X1 U6375 ( .A(n12078), .ZN(n23616) );
  AOI22_X1 U6376 ( .A1(\mem[311][2] ), .A2(n12076), .B1(n26819), .B2(
        data_in[2]), .ZN(n12078) );
  INV_X1 U6377 ( .A(n12079), .ZN(n23615) );
  AOI22_X1 U6378 ( .A1(\mem[311][3] ), .A2(n12076), .B1(n26819), .B2(
        data_in[3]), .ZN(n12079) );
  INV_X1 U6379 ( .A(n12080), .ZN(n23614) );
  AOI22_X1 U6380 ( .A1(\mem[311][4] ), .A2(n12076), .B1(n26819), .B2(
        data_in[4]), .ZN(n12080) );
  INV_X1 U6381 ( .A(n12081), .ZN(n23613) );
  AOI22_X1 U6382 ( .A1(\mem[311][5] ), .A2(n12076), .B1(n26819), .B2(
        data_in[5]), .ZN(n12081) );
  INV_X1 U6383 ( .A(n12082), .ZN(n23612) );
  AOI22_X1 U6384 ( .A1(\mem[311][6] ), .A2(n12076), .B1(n26819), .B2(
        data_in[6]), .ZN(n12082) );
  INV_X1 U6385 ( .A(n12083), .ZN(n23611) );
  AOI22_X1 U6386 ( .A1(\mem[311][7] ), .A2(n12076), .B1(n26819), .B2(
        data_in[7]), .ZN(n12083) );
  INV_X1 U6387 ( .A(n12084), .ZN(n23610) );
  AOI22_X1 U6388 ( .A1(\mem[312][0] ), .A2(n12085), .B1(n26818), .B2(
        data_in[0]), .ZN(n12084) );
  INV_X1 U6389 ( .A(n12086), .ZN(n23609) );
  AOI22_X1 U6390 ( .A1(\mem[312][1] ), .A2(n12085), .B1(n26818), .B2(
        data_in[1]), .ZN(n12086) );
  INV_X1 U6391 ( .A(n12087), .ZN(n23608) );
  AOI22_X1 U6392 ( .A1(\mem[312][2] ), .A2(n12085), .B1(n26818), .B2(
        data_in[2]), .ZN(n12087) );
  INV_X1 U6393 ( .A(n12088), .ZN(n23607) );
  AOI22_X1 U6394 ( .A1(\mem[312][3] ), .A2(n12085), .B1(n26818), .B2(
        data_in[3]), .ZN(n12088) );
  INV_X1 U6395 ( .A(n12089), .ZN(n23606) );
  AOI22_X1 U6396 ( .A1(\mem[312][4] ), .A2(n12085), .B1(n26818), .B2(
        data_in[4]), .ZN(n12089) );
  INV_X1 U6397 ( .A(n12090), .ZN(n23605) );
  AOI22_X1 U6398 ( .A1(\mem[312][5] ), .A2(n12085), .B1(n26818), .B2(
        data_in[5]), .ZN(n12090) );
  INV_X1 U6399 ( .A(n12091), .ZN(n23604) );
  AOI22_X1 U6400 ( .A1(\mem[312][6] ), .A2(n12085), .B1(n26818), .B2(
        data_in[6]), .ZN(n12091) );
  INV_X1 U6401 ( .A(n12092), .ZN(n23603) );
  AOI22_X1 U6402 ( .A1(\mem[312][7] ), .A2(n12085), .B1(n26818), .B2(
        data_in[7]), .ZN(n12092) );
  INV_X1 U6403 ( .A(n12093), .ZN(n23602) );
  AOI22_X1 U6404 ( .A1(\mem[313][0] ), .A2(n12094), .B1(n26817), .B2(
        data_in[0]), .ZN(n12093) );
  INV_X1 U6405 ( .A(n12095), .ZN(n23601) );
  AOI22_X1 U6406 ( .A1(\mem[313][1] ), .A2(n12094), .B1(n26817), .B2(
        data_in[1]), .ZN(n12095) );
  INV_X1 U6407 ( .A(n12096), .ZN(n23600) );
  AOI22_X1 U6408 ( .A1(\mem[313][2] ), .A2(n12094), .B1(n26817), .B2(
        data_in[2]), .ZN(n12096) );
  INV_X1 U6409 ( .A(n12097), .ZN(n23599) );
  AOI22_X1 U6410 ( .A1(\mem[313][3] ), .A2(n12094), .B1(n26817), .B2(
        data_in[3]), .ZN(n12097) );
  INV_X1 U6411 ( .A(n12098), .ZN(n23598) );
  AOI22_X1 U6412 ( .A1(\mem[313][4] ), .A2(n12094), .B1(n26817), .B2(
        data_in[4]), .ZN(n12098) );
  INV_X1 U6413 ( .A(n12099), .ZN(n23597) );
  AOI22_X1 U6414 ( .A1(\mem[313][5] ), .A2(n12094), .B1(n26817), .B2(
        data_in[5]), .ZN(n12099) );
  INV_X1 U6415 ( .A(n12100), .ZN(n23596) );
  AOI22_X1 U6416 ( .A1(\mem[313][6] ), .A2(n12094), .B1(n26817), .B2(
        data_in[6]), .ZN(n12100) );
  INV_X1 U6417 ( .A(n12101), .ZN(n23595) );
  AOI22_X1 U6418 ( .A1(\mem[313][7] ), .A2(n12094), .B1(n26817), .B2(
        data_in[7]), .ZN(n12101) );
  INV_X1 U6419 ( .A(n12102), .ZN(n23594) );
  AOI22_X1 U6420 ( .A1(\mem[314][0] ), .A2(n12103), .B1(n26816), .B2(
        data_in[0]), .ZN(n12102) );
  INV_X1 U6421 ( .A(n12104), .ZN(n23593) );
  AOI22_X1 U6422 ( .A1(\mem[314][1] ), .A2(n12103), .B1(n26816), .B2(
        data_in[1]), .ZN(n12104) );
  INV_X1 U6423 ( .A(n12105), .ZN(n23592) );
  AOI22_X1 U6424 ( .A1(\mem[314][2] ), .A2(n12103), .B1(n26816), .B2(
        data_in[2]), .ZN(n12105) );
  INV_X1 U6425 ( .A(n12106), .ZN(n23591) );
  AOI22_X1 U6426 ( .A1(\mem[314][3] ), .A2(n12103), .B1(n26816), .B2(
        data_in[3]), .ZN(n12106) );
  INV_X1 U6427 ( .A(n12107), .ZN(n23590) );
  AOI22_X1 U6428 ( .A1(\mem[314][4] ), .A2(n12103), .B1(n26816), .B2(
        data_in[4]), .ZN(n12107) );
  INV_X1 U6429 ( .A(n12108), .ZN(n23589) );
  AOI22_X1 U6430 ( .A1(\mem[314][5] ), .A2(n12103), .B1(n26816), .B2(
        data_in[5]), .ZN(n12108) );
  INV_X1 U6431 ( .A(n12109), .ZN(n23588) );
  AOI22_X1 U6432 ( .A1(\mem[314][6] ), .A2(n12103), .B1(n26816), .B2(
        data_in[6]), .ZN(n12109) );
  INV_X1 U6433 ( .A(n12110), .ZN(n23587) );
  AOI22_X1 U6434 ( .A1(\mem[314][7] ), .A2(n12103), .B1(n26816), .B2(
        data_in[7]), .ZN(n12110) );
  INV_X1 U6435 ( .A(n12111), .ZN(n23586) );
  AOI22_X1 U6436 ( .A1(\mem[315][0] ), .A2(n12112), .B1(n26815), .B2(
        data_in[0]), .ZN(n12111) );
  INV_X1 U6437 ( .A(n12113), .ZN(n23585) );
  AOI22_X1 U6438 ( .A1(\mem[315][1] ), .A2(n12112), .B1(n26815), .B2(
        data_in[1]), .ZN(n12113) );
  INV_X1 U6439 ( .A(n12114), .ZN(n23584) );
  AOI22_X1 U6440 ( .A1(\mem[315][2] ), .A2(n12112), .B1(n26815), .B2(
        data_in[2]), .ZN(n12114) );
  INV_X1 U6441 ( .A(n12115), .ZN(n23583) );
  AOI22_X1 U6442 ( .A1(\mem[315][3] ), .A2(n12112), .B1(n26815), .B2(
        data_in[3]), .ZN(n12115) );
  INV_X1 U6443 ( .A(n12116), .ZN(n23582) );
  AOI22_X1 U6444 ( .A1(\mem[315][4] ), .A2(n12112), .B1(n26815), .B2(
        data_in[4]), .ZN(n12116) );
  INV_X1 U6445 ( .A(n12117), .ZN(n23581) );
  AOI22_X1 U6446 ( .A1(\mem[315][5] ), .A2(n12112), .B1(n26815), .B2(
        data_in[5]), .ZN(n12117) );
  INV_X1 U6447 ( .A(n12118), .ZN(n23580) );
  AOI22_X1 U6448 ( .A1(\mem[315][6] ), .A2(n12112), .B1(n26815), .B2(
        data_in[6]), .ZN(n12118) );
  INV_X1 U6449 ( .A(n12119), .ZN(n23579) );
  AOI22_X1 U6450 ( .A1(\mem[315][7] ), .A2(n12112), .B1(n26815), .B2(
        data_in[7]), .ZN(n12119) );
  INV_X1 U6451 ( .A(n12120), .ZN(n23578) );
  AOI22_X1 U6452 ( .A1(\mem[316][0] ), .A2(n12121), .B1(n26814), .B2(
        data_in[0]), .ZN(n12120) );
  INV_X1 U6453 ( .A(n12122), .ZN(n23577) );
  AOI22_X1 U6454 ( .A1(\mem[316][1] ), .A2(n12121), .B1(n26814), .B2(
        data_in[1]), .ZN(n12122) );
  INV_X1 U6455 ( .A(n12123), .ZN(n23576) );
  AOI22_X1 U6456 ( .A1(\mem[316][2] ), .A2(n12121), .B1(n26814), .B2(
        data_in[2]), .ZN(n12123) );
  INV_X1 U6457 ( .A(n12124), .ZN(n23575) );
  AOI22_X1 U6458 ( .A1(\mem[316][3] ), .A2(n12121), .B1(n26814), .B2(
        data_in[3]), .ZN(n12124) );
  INV_X1 U6459 ( .A(n12125), .ZN(n23574) );
  AOI22_X1 U6460 ( .A1(\mem[316][4] ), .A2(n12121), .B1(n26814), .B2(
        data_in[4]), .ZN(n12125) );
  INV_X1 U6461 ( .A(n12126), .ZN(n23573) );
  AOI22_X1 U6462 ( .A1(\mem[316][5] ), .A2(n12121), .B1(n26814), .B2(
        data_in[5]), .ZN(n12126) );
  INV_X1 U6463 ( .A(n12127), .ZN(n23572) );
  AOI22_X1 U6464 ( .A1(\mem[316][6] ), .A2(n12121), .B1(n26814), .B2(
        data_in[6]), .ZN(n12127) );
  INV_X1 U6465 ( .A(n12128), .ZN(n23571) );
  AOI22_X1 U6466 ( .A1(\mem[316][7] ), .A2(n12121), .B1(n26814), .B2(
        data_in[7]), .ZN(n12128) );
  INV_X1 U6467 ( .A(n12129), .ZN(n23570) );
  AOI22_X1 U6468 ( .A1(\mem[317][0] ), .A2(n12130), .B1(n26813), .B2(
        data_in[0]), .ZN(n12129) );
  INV_X1 U6469 ( .A(n12131), .ZN(n23569) );
  AOI22_X1 U6470 ( .A1(\mem[317][1] ), .A2(n12130), .B1(n26813), .B2(
        data_in[1]), .ZN(n12131) );
  INV_X1 U6471 ( .A(n12132), .ZN(n23568) );
  AOI22_X1 U6472 ( .A1(\mem[317][2] ), .A2(n12130), .B1(n26813), .B2(
        data_in[2]), .ZN(n12132) );
  INV_X1 U6473 ( .A(n12133), .ZN(n23567) );
  AOI22_X1 U6474 ( .A1(\mem[317][3] ), .A2(n12130), .B1(n26813), .B2(
        data_in[3]), .ZN(n12133) );
  INV_X1 U6475 ( .A(n12134), .ZN(n23566) );
  AOI22_X1 U6476 ( .A1(\mem[317][4] ), .A2(n12130), .B1(n26813), .B2(
        data_in[4]), .ZN(n12134) );
  INV_X1 U6477 ( .A(n12135), .ZN(n23565) );
  AOI22_X1 U6478 ( .A1(\mem[317][5] ), .A2(n12130), .B1(n26813), .B2(
        data_in[5]), .ZN(n12135) );
  INV_X1 U6479 ( .A(n12136), .ZN(n23564) );
  AOI22_X1 U6480 ( .A1(\mem[317][6] ), .A2(n12130), .B1(n26813), .B2(
        data_in[6]), .ZN(n12136) );
  INV_X1 U6481 ( .A(n12137), .ZN(n23563) );
  AOI22_X1 U6482 ( .A1(\mem[317][7] ), .A2(n12130), .B1(n26813), .B2(
        data_in[7]), .ZN(n12137) );
  INV_X1 U6483 ( .A(n12138), .ZN(n23562) );
  AOI22_X1 U6484 ( .A1(\mem[318][0] ), .A2(n12139), .B1(n26812), .B2(
        data_in[0]), .ZN(n12138) );
  INV_X1 U6485 ( .A(n12140), .ZN(n23561) );
  AOI22_X1 U6486 ( .A1(\mem[318][1] ), .A2(n12139), .B1(n26812), .B2(
        data_in[1]), .ZN(n12140) );
  INV_X1 U6487 ( .A(n12141), .ZN(n23560) );
  AOI22_X1 U6488 ( .A1(\mem[318][2] ), .A2(n12139), .B1(n26812), .B2(
        data_in[2]), .ZN(n12141) );
  INV_X1 U6489 ( .A(n12142), .ZN(n23559) );
  AOI22_X1 U6490 ( .A1(\mem[318][3] ), .A2(n12139), .B1(n26812), .B2(
        data_in[3]), .ZN(n12142) );
  INV_X1 U6491 ( .A(n12143), .ZN(n23558) );
  AOI22_X1 U6492 ( .A1(\mem[318][4] ), .A2(n12139), .B1(n26812), .B2(
        data_in[4]), .ZN(n12143) );
  INV_X1 U6493 ( .A(n12144), .ZN(n23557) );
  AOI22_X1 U6494 ( .A1(\mem[318][5] ), .A2(n12139), .B1(n26812), .B2(
        data_in[5]), .ZN(n12144) );
  INV_X1 U6495 ( .A(n12145), .ZN(n23556) );
  AOI22_X1 U6496 ( .A1(\mem[318][6] ), .A2(n12139), .B1(n26812), .B2(
        data_in[6]), .ZN(n12145) );
  INV_X1 U6497 ( .A(n12146), .ZN(n23555) );
  AOI22_X1 U6498 ( .A1(\mem[318][7] ), .A2(n12139), .B1(n26812), .B2(
        data_in[7]), .ZN(n12146) );
  INV_X1 U6499 ( .A(n12147), .ZN(n23554) );
  AOI22_X1 U6500 ( .A1(\mem[319][0] ), .A2(n12148), .B1(n26811), .B2(
        data_in[0]), .ZN(n12147) );
  INV_X1 U6501 ( .A(n12149), .ZN(n23553) );
  AOI22_X1 U6502 ( .A1(\mem[319][1] ), .A2(n12148), .B1(n26811), .B2(
        data_in[1]), .ZN(n12149) );
  INV_X1 U6503 ( .A(n12150), .ZN(n23552) );
  AOI22_X1 U6504 ( .A1(\mem[319][2] ), .A2(n12148), .B1(n26811), .B2(
        data_in[2]), .ZN(n12150) );
  INV_X1 U6505 ( .A(n12151), .ZN(n23551) );
  AOI22_X1 U6506 ( .A1(\mem[319][3] ), .A2(n12148), .B1(n26811), .B2(
        data_in[3]), .ZN(n12151) );
  INV_X1 U6507 ( .A(n12152), .ZN(n23550) );
  AOI22_X1 U6508 ( .A1(\mem[319][4] ), .A2(n12148), .B1(n26811), .B2(
        data_in[4]), .ZN(n12152) );
  INV_X1 U6509 ( .A(n12153), .ZN(n23549) );
  AOI22_X1 U6510 ( .A1(\mem[319][5] ), .A2(n12148), .B1(n26811), .B2(
        data_in[5]), .ZN(n12153) );
  INV_X1 U6511 ( .A(n12154), .ZN(n23548) );
  AOI22_X1 U6512 ( .A1(\mem[319][6] ), .A2(n12148), .B1(n26811), .B2(
        data_in[6]), .ZN(n12154) );
  INV_X1 U6513 ( .A(n12155), .ZN(n23547) );
  AOI22_X1 U6514 ( .A1(\mem[319][7] ), .A2(n12148), .B1(n26811), .B2(
        data_in[7]), .ZN(n12155) );
  INV_X1 U6515 ( .A(n12229), .ZN(n23482) );
  AOI22_X1 U6516 ( .A1(\mem[328][0] ), .A2(n12230), .B1(n26802), .B2(
        data_in[0]), .ZN(n12229) );
  INV_X1 U6517 ( .A(n12231), .ZN(n23481) );
  AOI22_X1 U6518 ( .A1(\mem[328][1] ), .A2(n12230), .B1(n26802), .B2(
        data_in[1]), .ZN(n12231) );
  INV_X1 U6519 ( .A(n12232), .ZN(n23480) );
  AOI22_X1 U6520 ( .A1(\mem[328][2] ), .A2(n12230), .B1(n26802), .B2(
        data_in[2]), .ZN(n12232) );
  INV_X1 U6521 ( .A(n12233), .ZN(n23479) );
  AOI22_X1 U6522 ( .A1(\mem[328][3] ), .A2(n12230), .B1(n26802), .B2(
        data_in[3]), .ZN(n12233) );
  INV_X1 U6523 ( .A(n12234), .ZN(n23478) );
  AOI22_X1 U6524 ( .A1(\mem[328][4] ), .A2(n12230), .B1(n26802), .B2(
        data_in[4]), .ZN(n12234) );
  INV_X1 U6525 ( .A(n12235), .ZN(n23477) );
  AOI22_X1 U6526 ( .A1(\mem[328][5] ), .A2(n12230), .B1(n26802), .B2(
        data_in[5]), .ZN(n12235) );
  INV_X1 U6527 ( .A(n12236), .ZN(n23476) );
  AOI22_X1 U6528 ( .A1(\mem[328][6] ), .A2(n12230), .B1(n26802), .B2(
        data_in[6]), .ZN(n12236) );
  INV_X1 U6529 ( .A(n12237), .ZN(n23475) );
  AOI22_X1 U6530 ( .A1(\mem[328][7] ), .A2(n12230), .B1(n26802), .B2(
        data_in[7]), .ZN(n12237) );
  INV_X1 U6531 ( .A(n12238), .ZN(n23474) );
  AOI22_X1 U6532 ( .A1(\mem[329][0] ), .A2(n12239), .B1(n26801), .B2(
        data_in[0]), .ZN(n12238) );
  INV_X1 U6533 ( .A(n12240), .ZN(n23473) );
  AOI22_X1 U6534 ( .A1(\mem[329][1] ), .A2(n12239), .B1(n26801), .B2(
        data_in[1]), .ZN(n12240) );
  INV_X1 U6535 ( .A(n12241), .ZN(n23472) );
  AOI22_X1 U6536 ( .A1(\mem[329][2] ), .A2(n12239), .B1(n26801), .B2(
        data_in[2]), .ZN(n12241) );
  INV_X1 U6537 ( .A(n12242), .ZN(n23471) );
  AOI22_X1 U6538 ( .A1(\mem[329][3] ), .A2(n12239), .B1(n26801), .B2(
        data_in[3]), .ZN(n12242) );
  INV_X1 U6539 ( .A(n12243), .ZN(n23470) );
  AOI22_X1 U6540 ( .A1(\mem[329][4] ), .A2(n12239), .B1(n26801), .B2(
        data_in[4]), .ZN(n12243) );
  INV_X1 U6541 ( .A(n12244), .ZN(n23469) );
  AOI22_X1 U6542 ( .A1(\mem[329][5] ), .A2(n12239), .B1(n26801), .B2(
        data_in[5]), .ZN(n12244) );
  INV_X1 U6543 ( .A(n12245), .ZN(n23468) );
  AOI22_X1 U6544 ( .A1(\mem[329][6] ), .A2(n12239), .B1(n26801), .B2(
        data_in[6]), .ZN(n12245) );
  INV_X1 U6545 ( .A(n12246), .ZN(n23467) );
  AOI22_X1 U6546 ( .A1(\mem[329][7] ), .A2(n12239), .B1(n26801), .B2(
        data_in[7]), .ZN(n12246) );
  INV_X1 U6547 ( .A(n12247), .ZN(n23466) );
  AOI22_X1 U6548 ( .A1(\mem[330][0] ), .A2(n12248), .B1(n26800), .B2(
        data_in[0]), .ZN(n12247) );
  INV_X1 U6549 ( .A(n12249), .ZN(n23465) );
  AOI22_X1 U6550 ( .A1(\mem[330][1] ), .A2(n12248), .B1(n26800), .B2(
        data_in[1]), .ZN(n12249) );
  INV_X1 U6551 ( .A(n12250), .ZN(n23464) );
  AOI22_X1 U6552 ( .A1(\mem[330][2] ), .A2(n12248), .B1(n26800), .B2(
        data_in[2]), .ZN(n12250) );
  INV_X1 U6553 ( .A(n12251), .ZN(n23463) );
  AOI22_X1 U6554 ( .A1(\mem[330][3] ), .A2(n12248), .B1(n26800), .B2(
        data_in[3]), .ZN(n12251) );
  INV_X1 U6555 ( .A(n12252), .ZN(n23462) );
  AOI22_X1 U6556 ( .A1(\mem[330][4] ), .A2(n12248), .B1(n26800), .B2(
        data_in[4]), .ZN(n12252) );
  INV_X1 U6557 ( .A(n12253), .ZN(n23461) );
  AOI22_X1 U6558 ( .A1(\mem[330][5] ), .A2(n12248), .B1(n26800), .B2(
        data_in[5]), .ZN(n12253) );
  INV_X1 U6559 ( .A(n12254), .ZN(n23460) );
  AOI22_X1 U6560 ( .A1(\mem[330][6] ), .A2(n12248), .B1(n26800), .B2(
        data_in[6]), .ZN(n12254) );
  INV_X1 U6561 ( .A(n12255), .ZN(n23459) );
  AOI22_X1 U6562 ( .A1(\mem[330][7] ), .A2(n12248), .B1(n26800), .B2(
        data_in[7]), .ZN(n12255) );
  INV_X1 U6563 ( .A(n12256), .ZN(n23458) );
  AOI22_X1 U6564 ( .A1(\mem[331][0] ), .A2(n12257), .B1(n26799), .B2(
        data_in[0]), .ZN(n12256) );
  INV_X1 U6565 ( .A(n12258), .ZN(n23457) );
  AOI22_X1 U6566 ( .A1(\mem[331][1] ), .A2(n12257), .B1(n26799), .B2(
        data_in[1]), .ZN(n12258) );
  INV_X1 U6567 ( .A(n12259), .ZN(n23456) );
  AOI22_X1 U6568 ( .A1(\mem[331][2] ), .A2(n12257), .B1(n26799), .B2(
        data_in[2]), .ZN(n12259) );
  INV_X1 U6569 ( .A(n12260), .ZN(n23455) );
  AOI22_X1 U6570 ( .A1(\mem[331][3] ), .A2(n12257), .B1(n26799), .B2(
        data_in[3]), .ZN(n12260) );
  INV_X1 U6571 ( .A(n12261), .ZN(n23454) );
  AOI22_X1 U6572 ( .A1(\mem[331][4] ), .A2(n12257), .B1(n26799), .B2(
        data_in[4]), .ZN(n12261) );
  INV_X1 U6573 ( .A(n12262), .ZN(n23453) );
  AOI22_X1 U6574 ( .A1(\mem[331][5] ), .A2(n12257), .B1(n26799), .B2(
        data_in[5]), .ZN(n12262) );
  INV_X1 U6575 ( .A(n12263), .ZN(n23452) );
  AOI22_X1 U6576 ( .A1(\mem[331][6] ), .A2(n12257), .B1(n26799), .B2(
        data_in[6]), .ZN(n12263) );
  INV_X1 U6577 ( .A(n12264), .ZN(n23451) );
  AOI22_X1 U6578 ( .A1(\mem[331][7] ), .A2(n12257), .B1(n26799), .B2(
        data_in[7]), .ZN(n12264) );
  INV_X1 U6579 ( .A(n12265), .ZN(n23450) );
  AOI22_X1 U6580 ( .A1(\mem[332][0] ), .A2(n12266), .B1(n26798), .B2(
        data_in[0]), .ZN(n12265) );
  INV_X1 U6581 ( .A(n12267), .ZN(n23449) );
  AOI22_X1 U6582 ( .A1(\mem[332][1] ), .A2(n12266), .B1(n26798), .B2(
        data_in[1]), .ZN(n12267) );
  INV_X1 U6583 ( .A(n12268), .ZN(n23448) );
  AOI22_X1 U6584 ( .A1(\mem[332][2] ), .A2(n12266), .B1(n26798), .B2(
        data_in[2]), .ZN(n12268) );
  INV_X1 U6585 ( .A(n12269), .ZN(n23447) );
  AOI22_X1 U6586 ( .A1(\mem[332][3] ), .A2(n12266), .B1(n26798), .B2(
        data_in[3]), .ZN(n12269) );
  INV_X1 U6587 ( .A(n12270), .ZN(n23446) );
  AOI22_X1 U6588 ( .A1(\mem[332][4] ), .A2(n12266), .B1(n26798), .B2(
        data_in[4]), .ZN(n12270) );
  INV_X1 U6589 ( .A(n12271), .ZN(n23445) );
  AOI22_X1 U6590 ( .A1(\mem[332][5] ), .A2(n12266), .B1(n26798), .B2(
        data_in[5]), .ZN(n12271) );
  INV_X1 U6591 ( .A(n12272), .ZN(n23444) );
  AOI22_X1 U6592 ( .A1(\mem[332][6] ), .A2(n12266), .B1(n26798), .B2(
        data_in[6]), .ZN(n12272) );
  INV_X1 U6593 ( .A(n12273), .ZN(n23443) );
  AOI22_X1 U6594 ( .A1(\mem[332][7] ), .A2(n12266), .B1(n26798), .B2(
        data_in[7]), .ZN(n12273) );
  INV_X1 U6595 ( .A(n12274), .ZN(n23442) );
  AOI22_X1 U6596 ( .A1(\mem[333][0] ), .A2(n12275), .B1(n26797), .B2(
        data_in[0]), .ZN(n12274) );
  INV_X1 U6597 ( .A(n12276), .ZN(n23441) );
  AOI22_X1 U6598 ( .A1(\mem[333][1] ), .A2(n12275), .B1(n26797), .B2(
        data_in[1]), .ZN(n12276) );
  INV_X1 U6599 ( .A(n12277), .ZN(n23440) );
  AOI22_X1 U6600 ( .A1(\mem[333][2] ), .A2(n12275), .B1(n26797), .B2(
        data_in[2]), .ZN(n12277) );
  INV_X1 U6601 ( .A(n12278), .ZN(n23439) );
  AOI22_X1 U6602 ( .A1(\mem[333][3] ), .A2(n12275), .B1(n26797), .B2(
        data_in[3]), .ZN(n12278) );
  INV_X1 U6603 ( .A(n12279), .ZN(n23438) );
  AOI22_X1 U6604 ( .A1(\mem[333][4] ), .A2(n12275), .B1(n26797), .B2(
        data_in[4]), .ZN(n12279) );
  INV_X1 U6605 ( .A(n12280), .ZN(n23437) );
  AOI22_X1 U6606 ( .A1(\mem[333][5] ), .A2(n12275), .B1(n26797), .B2(
        data_in[5]), .ZN(n12280) );
  INV_X1 U6607 ( .A(n12281), .ZN(n23436) );
  AOI22_X1 U6608 ( .A1(\mem[333][6] ), .A2(n12275), .B1(n26797), .B2(
        data_in[6]), .ZN(n12281) );
  INV_X1 U6609 ( .A(n12282), .ZN(n23435) );
  AOI22_X1 U6610 ( .A1(\mem[333][7] ), .A2(n12275), .B1(n26797), .B2(
        data_in[7]), .ZN(n12282) );
  INV_X1 U6611 ( .A(n12283), .ZN(n23434) );
  AOI22_X1 U6612 ( .A1(\mem[334][0] ), .A2(n12284), .B1(n26796), .B2(
        data_in[0]), .ZN(n12283) );
  INV_X1 U6613 ( .A(n12285), .ZN(n23433) );
  AOI22_X1 U6614 ( .A1(\mem[334][1] ), .A2(n12284), .B1(n26796), .B2(
        data_in[1]), .ZN(n12285) );
  INV_X1 U6615 ( .A(n12286), .ZN(n23432) );
  AOI22_X1 U6616 ( .A1(\mem[334][2] ), .A2(n12284), .B1(n26796), .B2(
        data_in[2]), .ZN(n12286) );
  INV_X1 U6617 ( .A(n12287), .ZN(n23431) );
  AOI22_X1 U6618 ( .A1(\mem[334][3] ), .A2(n12284), .B1(n26796), .B2(
        data_in[3]), .ZN(n12287) );
  INV_X1 U6619 ( .A(n12288), .ZN(n23430) );
  AOI22_X1 U6620 ( .A1(\mem[334][4] ), .A2(n12284), .B1(n26796), .B2(
        data_in[4]), .ZN(n12288) );
  INV_X1 U6621 ( .A(n12289), .ZN(n23429) );
  AOI22_X1 U6622 ( .A1(\mem[334][5] ), .A2(n12284), .B1(n26796), .B2(
        data_in[5]), .ZN(n12289) );
  INV_X1 U6623 ( .A(n12290), .ZN(n23428) );
  AOI22_X1 U6624 ( .A1(\mem[334][6] ), .A2(n12284), .B1(n26796), .B2(
        data_in[6]), .ZN(n12290) );
  INV_X1 U6625 ( .A(n12291), .ZN(n23427) );
  AOI22_X1 U6626 ( .A1(\mem[334][7] ), .A2(n12284), .B1(n26796), .B2(
        data_in[7]), .ZN(n12291) );
  INV_X1 U6627 ( .A(n12292), .ZN(n23426) );
  AOI22_X1 U6628 ( .A1(\mem[335][0] ), .A2(n12293), .B1(n26795), .B2(
        data_in[0]), .ZN(n12292) );
  INV_X1 U6629 ( .A(n12294), .ZN(n23425) );
  AOI22_X1 U6630 ( .A1(\mem[335][1] ), .A2(n12293), .B1(n26795), .B2(
        data_in[1]), .ZN(n12294) );
  INV_X1 U6631 ( .A(n12295), .ZN(n23424) );
  AOI22_X1 U6632 ( .A1(\mem[335][2] ), .A2(n12293), .B1(n26795), .B2(
        data_in[2]), .ZN(n12295) );
  INV_X1 U6633 ( .A(n12296), .ZN(n23423) );
  AOI22_X1 U6634 ( .A1(\mem[335][3] ), .A2(n12293), .B1(n26795), .B2(
        data_in[3]), .ZN(n12296) );
  INV_X1 U6635 ( .A(n12297), .ZN(n23422) );
  AOI22_X1 U6636 ( .A1(\mem[335][4] ), .A2(n12293), .B1(n26795), .B2(
        data_in[4]), .ZN(n12297) );
  INV_X1 U6637 ( .A(n12298), .ZN(n23421) );
  AOI22_X1 U6638 ( .A1(\mem[335][5] ), .A2(n12293), .B1(n26795), .B2(
        data_in[5]), .ZN(n12298) );
  INV_X1 U6639 ( .A(n12299), .ZN(n23420) );
  AOI22_X1 U6640 ( .A1(\mem[335][6] ), .A2(n12293), .B1(n26795), .B2(
        data_in[6]), .ZN(n12299) );
  INV_X1 U6641 ( .A(n12300), .ZN(n23419) );
  AOI22_X1 U6642 ( .A1(\mem[335][7] ), .A2(n12293), .B1(n26795), .B2(
        data_in[7]), .ZN(n12300) );
  INV_X1 U6643 ( .A(n12301), .ZN(n23418) );
  AOI22_X1 U6644 ( .A1(\mem[336][0] ), .A2(n12302), .B1(n26794), .B2(
        data_in[0]), .ZN(n12301) );
  INV_X1 U6645 ( .A(n12303), .ZN(n23417) );
  AOI22_X1 U6646 ( .A1(\mem[336][1] ), .A2(n12302), .B1(n26794), .B2(
        data_in[1]), .ZN(n12303) );
  INV_X1 U6647 ( .A(n12304), .ZN(n23416) );
  AOI22_X1 U6648 ( .A1(\mem[336][2] ), .A2(n12302), .B1(n26794), .B2(
        data_in[2]), .ZN(n12304) );
  INV_X1 U6649 ( .A(n12305), .ZN(n23415) );
  AOI22_X1 U6650 ( .A1(\mem[336][3] ), .A2(n12302), .B1(n26794), .B2(
        data_in[3]), .ZN(n12305) );
  INV_X1 U6651 ( .A(n12306), .ZN(n23414) );
  AOI22_X1 U6652 ( .A1(\mem[336][4] ), .A2(n12302), .B1(n26794), .B2(
        data_in[4]), .ZN(n12306) );
  INV_X1 U6653 ( .A(n12307), .ZN(n23413) );
  AOI22_X1 U6654 ( .A1(\mem[336][5] ), .A2(n12302), .B1(n26794), .B2(
        data_in[5]), .ZN(n12307) );
  INV_X1 U6655 ( .A(n12308), .ZN(n23412) );
  AOI22_X1 U6656 ( .A1(\mem[336][6] ), .A2(n12302), .B1(n26794), .B2(
        data_in[6]), .ZN(n12308) );
  INV_X1 U6657 ( .A(n12309), .ZN(n23411) );
  AOI22_X1 U6658 ( .A1(\mem[336][7] ), .A2(n12302), .B1(n26794), .B2(
        data_in[7]), .ZN(n12309) );
  INV_X1 U6659 ( .A(n12310), .ZN(n23410) );
  AOI22_X1 U6660 ( .A1(\mem[337][0] ), .A2(n12311), .B1(n26793), .B2(
        data_in[0]), .ZN(n12310) );
  INV_X1 U6661 ( .A(n12312), .ZN(n23409) );
  AOI22_X1 U6662 ( .A1(\mem[337][1] ), .A2(n12311), .B1(n26793), .B2(
        data_in[1]), .ZN(n12312) );
  INV_X1 U6663 ( .A(n12313), .ZN(n23408) );
  AOI22_X1 U6664 ( .A1(\mem[337][2] ), .A2(n12311), .B1(n26793), .B2(
        data_in[2]), .ZN(n12313) );
  INV_X1 U6665 ( .A(n12314), .ZN(n23407) );
  AOI22_X1 U6666 ( .A1(\mem[337][3] ), .A2(n12311), .B1(n26793), .B2(
        data_in[3]), .ZN(n12314) );
  INV_X1 U6667 ( .A(n12315), .ZN(n23406) );
  AOI22_X1 U6668 ( .A1(\mem[337][4] ), .A2(n12311), .B1(n26793), .B2(
        data_in[4]), .ZN(n12315) );
  INV_X1 U6669 ( .A(n12316), .ZN(n23405) );
  AOI22_X1 U6670 ( .A1(\mem[337][5] ), .A2(n12311), .B1(n26793), .B2(
        data_in[5]), .ZN(n12316) );
  INV_X1 U6671 ( .A(n12317), .ZN(n23404) );
  AOI22_X1 U6672 ( .A1(\mem[337][6] ), .A2(n12311), .B1(n26793), .B2(
        data_in[6]), .ZN(n12317) );
  INV_X1 U6673 ( .A(n12318), .ZN(n23403) );
  AOI22_X1 U6674 ( .A1(\mem[337][7] ), .A2(n12311), .B1(n26793), .B2(
        data_in[7]), .ZN(n12318) );
  INV_X1 U6675 ( .A(n12319), .ZN(n23402) );
  AOI22_X1 U6676 ( .A1(\mem[338][0] ), .A2(n12320), .B1(n26792), .B2(
        data_in[0]), .ZN(n12319) );
  INV_X1 U6677 ( .A(n12321), .ZN(n23401) );
  AOI22_X1 U6678 ( .A1(\mem[338][1] ), .A2(n12320), .B1(n26792), .B2(
        data_in[1]), .ZN(n12321) );
  INV_X1 U6679 ( .A(n12322), .ZN(n23400) );
  AOI22_X1 U6680 ( .A1(\mem[338][2] ), .A2(n12320), .B1(n26792), .B2(
        data_in[2]), .ZN(n12322) );
  INV_X1 U6681 ( .A(n12323), .ZN(n23399) );
  AOI22_X1 U6682 ( .A1(\mem[338][3] ), .A2(n12320), .B1(n26792), .B2(
        data_in[3]), .ZN(n12323) );
  INV_X1 U6683 ( .A(n12324), .ZN(n23398) );
  AOI22_X1 U6684 ( .A1(\mem[338][4] ), .A2(n12320), .B1(n26792), .B2(
        data_in[4]), .ZN(n12324) );
  INV_X1 U6685 ( .A(n12325), .ZN(n23397) );
  AOI22_X1 U6686 ( .A1(\mem[338][5] ), .A2(n12320), .B1(n26792), .B2(
        data_in[5]), .ZN(n12325) );
  INV_X1 U6687 ( .A(n12326), .ZN(n23396) );
  AOI22_X1 U6688 ( .A1(\mem[338][6] ), .A2(n12320), .B1(n26792), .B2(
        data_in[6]), .ZN(n12326) );
  INV_X1 U6689 ( .A(n12327), .ZN(n23395) );
  AOI22_X1 U6690 ( .A1(\mem[338][7] ), .A2(n12320), .B1(n26792), .B2(
        data_in[7]), .ZN(n12327) );
  INV_X1 U6691 ( .A(n12328), .ZN(n23394) );
  AOI22_X1 U6692 ( .A1(\mem[339][0] ), .A2(n12329), .B1(n26791), .B2(
        data_in[0]), .ZN(n12328) );
  INV_X1 U6693 ( .A(n12330), .ZN(n23393) );
  AOI22_X1 U6694 ( .A1(\mem[339][1] ), .A2(n12329), .B1(n26791), .B2(
        data_in[1]), .ZN(n12330) );
  INV_X1 U6695 ( .A(n12331), .ZN(n23392) );
  AOI22_X1 U6696 ( .A1(\mem[339][2] ), .A2(n12329), .B1(n26791), .B2(
        data_in[2]), .ZN(n12331) );
  INV_X1 U6697 ( .A(n12332), .ZN(n23391) );
  AOI22_X1 U6698 ( .A1(\mem[339][3] ), .A2(n12329), .B1(n26791), .B2(
        data_in[3]), .ZN(n12332) );
  INV_X1 U6699 ( .A(n12333), .ZN(n23390) );
  AOI22_X1 U6700 ( .A1(\mem[339][4] ), .A2(n12329), .B1(n26791), .B2(
        data_in[4]), .ZN(n12333) );
  INV_X1 U6701 ( .A(n12334), .ZN(n23389) );
  AOI22_X1 U6702 ( .A1(\mem[339][5] ), .A2(n12329), .B1(n26791), .B2(
        data_in[5]), .ZN(n12334) );
  INV_X1 U6703 ( .A(n12335), .ZN(n23388) );
  AOI22_X1 U6704 ( .A1(\mem[339][6] ), .A2(n12329), .B1(n26791), .B2(
        data_in[6]), .ZN(n12335) );
  INV_X1 U6705 ( .A(n12336), .ZN(n23387) );
  AOI22_X1 U6706 ( .A1(\mem[339][7] ), .A2(n12329), .B1(n26791), .B2(
        data_in[7]), .ZN(n12336) );
  INV_X1 U6707 ( .A(n12337), .ZN(n23386) );
  AOI22_X1 U6708 ( .A1(\mem[340][0] ), .A2(n12338), .B1(n26790), .B2(
        data_in[0]), .ZN(n12337) );
  INV_X1 U6709 ( .A(n12339), .ZN(n23385) );
  AOI22_X1 U6710 ( .A1(\mem[340][1] ), .A2(n12338), .B1(n26790), .B2(
        data_in[1]), .ZN(n12339) );
  INV_X1 U6711 ( .A(n12340), .ZN(n23384) );
  AOI22_X1 U6712 ( .A1(\mem[340][2] ), .A2(n12338), .B1(n26790), .B2(
        data_in[2]), .ZN(n12340) );
  INV_X1 U6713 ( .A(n12341), .ZN(n23383) );
  AOI22_X1 U6714 ( .A1(\mem[340][3] ), .A2(n12338), .B1(n26790), .B2(
        data_in[3]), .ZN(n12341) );
  INV_X1 U6715 ( .A(n12342), .ZN(n23382) );
  AOI22_X1 U6716 ( .A1(\mem[340][4] ), .A2(n12338), .B1(n26790), .B2(
        data_in[4]), .ZN(n12342) );
  INV_X1 U6717 ( .A(n12343), .ZN(n23381) );
  AOI22_X1 U6718 ( .A1(\mem[340][5] ), .A2(n12338), .B1(n26790), .B2(
        data_in[5]), .ZN(n12343) );
  INV_X1 U6719 ( .A(n12344), .ZN(n23380) );
  AOI22_X1 U6720 ( .A1(\mem[340][6] ), .A2(n12338), .B1(n26790), .B2(
        data_in[6]), .ZN(n12344) );
  INV_X1 U6721 ( .A(n12345), .ZN(n23379) );
  AOI22_X1 U6722 ( .A1(\mem[340][7] ), .A2(n12338), .B1(n26790), .B2(
        data_in[7]), .ZN(n12345) );
  INV_X1 U6723 ( .A(n12346), .ZN(n23378) );
  AOI22_X1 U6724 ( .A1(\mem[341][0] ), .A2(n12347), .B1(n26789), .B2(
        data_in[0]), .ZN(n12346) );
  INV_X1 U6725 ( .A(n12348), .ZN(n23377) );
  AOI22_X1 U6726 ( .A1(\mem[341][1] ), .A2(n12347), .B1(n26789), .B2(
        data_in[1]), .ZN(n12348) );
  INV_X1 U6727 ( .A(n12349), .ZN(n23376) );
  AOI22_X1 U6728 ( .A1(\mem[341][2] ), .A2(n12347), .B1(n26789), .B2(
        data_in[2]), .ZN(n12349) );
  INV_X1 U6729 ( .A(n12350), .ZN(n23375) );
  AOI22_X1 U6730 ( .A1(\mem[341][3] ), .A2(n12347), .B1(n26789), .B2(
        data_in[3]), .ZN(n12350) );
  INV_X1 U6731 ( .A(n12351), .ZN(n23374) );
  AOI22_X1 U6732 ( .A1(\mem[341][4] ), .A2(n12347), .B1(n26789), .B2(
        data_in[4]), .ZN(n12351) );
  INV_X1 U6733 ( .A(n12352), .ZN(n23373) );
  AOI22_X1 U6734 ( .A1(\mem[341][5] ), .A2(n12347), .B1(n26789), .B2(
        data_in[5]), .ZN(n12352) );
  INV_X1 U6735 ( .A(n12353), .ZN(n23372) );
  AOI22_X1 U6736 ( .A1(\mem[341][6] ), .A2(n12347), .B1(n26789), .B2(
        data_in[6]), .ZN(n12353) );
  INV_X1 U6737 ( .A(n12354), .ZN(n23371) );
  AOI22_X1 U6738 ( .A1(\mem[341][7] ), .A2(n12347), .B1(n26789), .B2(
        data_in[7]), .ZN(n12354) );
  INV_X1 U6739 ( .A(n12355), .ZN(n23370) );
  AOI22_X1 U6740 ( .A1(\mem[342][0] ), .A2(n12356), .B1(n26788), .B2(
        data_in[0]), .ZN(n12355) );
  INV_X1 U6741 ( .A(n12357), .ZN(n23369) );
  AOI22_X1 U6742 ( .A1(\mem[342][1] ), .A2(n12356), .B1(n26788), .B2(
        data_in[1]), .ZN(n12357) );
  INV_X1 U6743 ( .A(n12358), .ZN(n23368) );
  AOI22_X1 U6744 ( .A1(\mem[342][2] ), .A2(n12356), .B1(n26788), .B2(
        data_in[2]), .ZN(n12358) );
  INV_X1 U6745 ( .A(n12359), .ZN(n23367) );
  AOI22_X1 U6746 ( .A1(\mem[342][3] ), .A2(n12356), .B1(n26788), .B2(
        data_in[3]), .ZN(n12359) );
  INV_X1 U6747 ( .A(n12360), .ZN(n23366) );
  AOI22_X1 U6748 ( .A1(\mem[342][4] ), .A2(n12356), .B1(n26788), .B2(
        data_in[4]), .ZN(n12360) );
  INV_X1 U6749 ( .A(n12361), .ZN(n23365) );
  AOI22_X1 U6750 ( .A1(\mem[342][5] ), .A2(n12356), .B1(n26788), .B2(
        data_in[5]), .ZN(n12361) );
  INV_X1 U6751 ( .A(n12362), .ZN(n23364) );
  AOI22_X1 U6752 ( .A1(\mem[342][6] ), .A2(n12356), .B1(n26788), .B2(
        data_in[6]), .ZN(n12362) );
  INV_X1 U6753 ( .A(n12363), .ZN(n23363) );
  AOI22_X1 U6754 ( .A1(\mem[342][7] ), .A2(n12356), .B1(n26788), .B2(
        data_in[7]), .ZN(n12363) );
  INV_X1 U6755 ( .A(n12364), .ZN(n23362) );
  AOI22_X1 U6756 ( .A1(\mem[343][0] ), .A2(n12365), .B1(n26787), .B2(
        data_in[0]), .ZN(n12364) );
  INV_X1 U6757 ( .A(n12366), .ZN(n23361) );
  AOI22_X1 U6758 ( .A1(\mem[343][1] ), .A2(n12365), .B1(n26787), .B2(
        data_in[1]), .ZN(n12366) );
  INV_X1 U6759 ( .A(n12367), .ZN(n23360) );
  AOI22_X1 U6760 ( .A1(\mem[343][2] ), .A2(n12365), .B1(n26787), .B2(
        data_in[2]), .ZN(n12367) );
  INV_X1 U6761 ( .A(n12368), .ZN(n23359) );
  AOI22_X1 U6762 ( .A1(\mem[343][3] ), .A2(n12365), .B1(n26787), .B2(
        data_in[3]), .ZN(n12368) );
  INV_X1 U6763 ( .A(n12369), .ZN(n23358) );
  AOI22_X1 U6764 ( .A1(\mem[343][4] ), .A2(n12365), .B1(n26787), .B2(
        data_in[4]), .ZN(n12369) );
  INV_X1 U6765 ( .A(n12370), .ZN(n23357) );
  AOI22_X1 U6766 ( .A1(\mem[343][5] ), .A2(n12365), .B1(n26787), .B2(
        data_in[5]), .ZN(n12370) );
  INV_X1 U6767 ( .A(n12371), .ZN(n23356) );
  AOI22_X1 U6768 ( .A1(\mem[343][6] ), .A2(n12365), .B1(n26787), .B2(
        data_in[6]), .ZN(n12371) );
  INV_X1 U6769 ( .A(n12372), .ZN(n23355) );
  AOI22_X1 U6770 ( .A1(\mem[343][7] ), .A2(n12365), .B1(n26787), .B2(
        data_in[7]), .ZN(n12372) );
  INV_X1 U6771 ( .A(n12373), .ZN(n23354) );
  AOI22_X1 U6772 ( .A1(\mem[344][0] ), .A2(n12374), .B1(n26786), .B2(
        data_in[0]), .ZN(n12373) );
  INV_X1 U6773 ( .A(n12375), .ZN(n23353) );
  AOI22_X1 U6774 ( .A1(\mem[344][1] ), .A2(n12374), .B1(n26786), .B2(
        data_in[1]), .ZN(n12375) );
  INV_X1 U6775 ( .A(n12376), .ZN(n23352) );
  AOI22_X1 U6776 ( .A1(\mem[344][2] ), .A2(n12374), .B1(n26786), .B2(
        data_in[2]), .ZN(n12376) );
  INV_X1 U6777 ( .A(n12377), .ZN(n23351) );
  AOI22_X1 U6778 ( .A1(\mem[344][3] ), .A2(n12374), .B1(n26786), .B2(
        data_in[3]), .ZN(n12377) );
  INV_X1 U6779 ( .A(n12378), .ZN(n23350) );
  AOI22_X1 U6780 ( .A1(\mem[344][4] ), .A2(n12374), .B1(n26786), .B2(
        data_in[4]), .ZN(n12378) );
  INV_X1 U6781 ( .A(n12379), .ZN(n23349) );
  AOI22_X1 U6782 ( .A1(\mem[344][5] ), .A2(n12374), .B1(n26786), .B2(
        data_in[5]), .ZN(n12379) );
  INV_X1 U6783 ( .A(n12380), .ZN(n23348) );
  AOI22_X1 U6784 ( .A1(\mem[344][6] ), .A2(n12374), .B1(n26786), .B2(
        data_in[6]), .ZN(n12380) );
  INV_X1 U6785 ( .A(n12381), .ZN(n23347) );
  AOI22_X1 U6786 ( .A1(\mem[344][7] ), .A2(n12374), .B1(n26786), .B2(
        data_in[7]), .ZN(n12381) );
  INV_X1 U6787 ( .A(n12382), .ZN(n23346) );
  AOI22_X1 U6788 ( .A1(\mem[345][0] ), .A2(n12383), .B1(n26785), .B2(
        data_in[0]), .ZN(n12382) );
  INV_X1 U6789 ( .A(n12384), .ZN(n23345) );
  AOI22_X1 U6790 ( .A1(\mem[345][1] ), .A2(n12383), .B1(n26785), .B2(
        data_in[1]), .ZN(n12384) );
  INV_X1 U6791 ( .A(n12385), .ZN(n23344) );
  AOI22_X1 U6792 ( .A1(\mem[345][2] ), .A2(n12383), .B1(n26785), .B2(
        data_in[2]), .ZN(n12385) );
  INV_X1 U6793 ( .A(n12386), .ZN(n23343) );
  AOI22_X1 U6794 ( .A1(\mem[345][3] ), .A2(n12383), .B1(n26785), .B2(
        data_in[3]), .ZN(n12386) );
  INV_X1 U6795 ( .A(n12387), .ZN(n23342) );
  AOI22_X1 U6796 ( .A1(\mem[345][4] ), .A2(n12383), .B1(n26785), .B2(
        data_in[4]), .ZN(n12387) );
  INV_X1 U6797 ( .A(n12388), .ZN(n23341) );
  AOI22_X1 U6798 ( .A1(\mem[345][5] ), .A2(n12383), .B1(n26785), .B2(
        data_in[5]), .ZN(n12388) );
  INV_X1 U6799 ( .A(n12389), .ZN(n23340) );
  AOI22_X1 U6800 ( .A1(\mem[345][6] ), .A2(n12383), .B1(n26785), .B2(
        data_in[6]), .ZN(n12389) );
  INV_X1 U6801 ( .A(n12390), .ZN(n23339) );
  AOI22_X1 U6802 ( .A1(\mem[345][7] ), .A2(n12383), .B1(n26785), .B2(
        data_in[7]), .ZN(n12390) );
  INV_X1 U6803 ( .A(n12391), .ZN(n23338) );
  AOI22_X1 U6804 ( .A1(\mem[346][0] ), .A2(n12392), .B1(n26784), .B2(
        data_in[0]), .ZN(n12391) );
  INV_X1 U6805 ( .A(n12393), .ZN(n23337) );
  AOI22_X1 U6806 ( .A1(\mem[346][1] ), .A2(n12392), .B1(n26784), .B2(
        data_in[1]), .ZN(n12393) );
  INV_X1 U6807 ( .A(n12394), .ZN(n23336) );
  AOI22_X1 U6808 ( .A1(\mem[346][2] ), .A2(n12392), .B1(n26784), .B2(
        data_in[2]), .ZN(n12394) );
  INV_X1 U6809 ( .A(n12395), .ZN(n23335) );
  AOI22_X1 U6810 ( .A1(\mem[346][3] ), .A2(n12392), .B1(n26784), .B2(
        data_in[3]), .ZN(n12395) );
  INV_X1 U6811 ( .A(n12396), .ZN(n23334) );
  AOI22_X1 U6812 ( .A1(\mem[346][4] ), .A2(n12392), .B1(n26784), .B2(
        data_in[4]), .ZN(n12396) );
  INV_X1 U6813 ( .A(n12397), .ZN(n23333) );
  AOI22_X1 U6814 ( .A1(\mem[346][5] ), .A2(n12392), .B1(n26784), .B2(
        data_in[5]), .ZN(n12397) );
  INV_X1 U6815 ( .A(n12398), .ZN(n23332) );
  AOI22_X1 U6816 ( .A1(\mem[346][6] ), .A2(n12392), .B1(n26784), .B2(
        data_in[6]), .ZN(n12398) );
  INV_X1 U6817 ( .A(n12399), .ZN(n23331) );
  AOI22_X1 U6818 ( .A1(\mem[346][7] ), .A2(n12392), .B1(n26784), .B2(
        data_in[7]), .ZN(n12399) );
  INV_X1 U6819 ( .A(n12400), .ZN(n23330) );
  AOI22_X1 U6820 ( .A1(\mem[347][0] ), .A2(n12401), .B1(n26783), .B2(
        data_in[0]), .ZN(n12400) );
  INV_X1 U6821 ( .A(n12402), .ZN(n23329) );
  AOI22_X1 U6822 ( .A1(\mem[347][1] ), .A2(n12401), .B1(n26783), .B2(
        data_in[1]), .ZN(n12402) );
  INV_X1 U6823 ( .A(n12403), .ZN(n23328) );
  AOI22_X1 U6824 ( .A1(\mem[347][2] ), .A2(n12401), .B1(n26783), .B2(
        data_in[2]), .ZN(n12403) );
  INV_X1 U6825 ( .A(n12404), .ZN(n23327) );
  AOI22_X1 U6826 ( .A1(\mem[347][3] ), .A2(n12401), .B1(n26783), .B2(
        data_in[3]), .ZN(n12404) );
  INV_X1 U6827 ( .A(n12405), .ZN(n23326) );
  AOI22_X1 U6828 ( .A1(\mem[347][4] ), .A2(n12401), .B1(n26783), .B2(
        data_in[4]), .ZN(n12405) );
  INV_X1 U6829 ( .A(n12406), .ZN(n23325) );
  AOI22_X1 U6830 ( .A1(\mem[347][5] ), .A2(n12401), .B1(n26783), .B2(
        data_in[5]), .ZN(n12406) );
  INV_X1 U6831 ( .A(n12407), .ZN(n23324) );
  AOI22_X1 U6832 ( .A1(\mem[347][6] ), .A2(n12401), .B1(n26783), .B2(
        data_in[6]), .ZN(n12407) );
  INV_X1 U6833 ( .A(n12408), .ZN(n23323) );
  AOI22_X1 U6834 ( .A1(\mem[347][7] ), .A2(n12401), .B1(n26783), .B2(
        data_in[7]), .ZN(n12408) );
  INV_X1 U6835 ( .A(n12409), .ZN(n23322) );
  AOI22_X1 U6836 ( .A1(\mem[348][0] ), .A2(n12410), .B1(n26782), .B2(
        data_in[0]), .ZN(n12409) );
  INV_X1 U6837 ( .A(n12411), .ZN(n23321) );
  AOI22_X1 U6838 ( .A1(\mem[348][1] ), .A2(n12410), .B1(n26782), .B2(
        data_in[1]), .ZN(n12411) );
  INV_X1 U6839 ( .A(n12412), .ZN(n23320) );
  AOI22_X1 U6840 ( .A1(\mem[348][2] ), .A2(n12410), .B1(n26782), .B2(
        data_in[2]), .ZN(n12412) );
  INV_X1 U6841 ( .A(n12413), .ZN(n23319) );
  AOI22_X1 U6842 ( .A1(\mem[348][3] ), .A2(n12410), .B1(n26782), .B2(
        data_in[3]), .ZN(n12413) );
  INV_X1 U6843 ( .A(n12414), .ZN(n23318) );
  AOI22_X1 U6844 ( .A1(\mem[348][4] ), .A2(n12410), .B1(n26782), .B2(
        data_in[4]), .ZN(n12414) );
  INV_X1 U6845 ( .A(n12415), .ZN(n23317) );
  AOI22_X1 U6846 ( .A1(\mem[348][5] ), .A2(n12410), .B1(n26782), .B2(
        data_in[5]), .ZN(n12415) );
  INV_X1 U6847 ( .A(n12416), .ZN(n23316) );
  AOI22_X1 U6848 ( .A1(\mem[348][6] ), .A2(n12410), .B1(n26782), .B2(
        data_in[6]), .ZN(n12416) );
  INV_X1 U6849 ( .A(n12417), .ZN(n23315) );
  AOI22_X1 U6850 ( .A1(\mem[348][7] ), .A2(n12410), .B1(n26782), .B2(
        data_in[7]), .ZN(n12417) );
  INV_X1 U6851 ( .A(n12418), .ZN(n23314) );
  AOI22_X1 U6852 ( .A1(\mem[349][0] ), .A2(n12419), .B1(n26781), .B2(
        data_in[0]), .ZN(n12418) );
  INV_X1 U6853 ( .A(n12420), .ZN(n23313) );
  AOI22_X1 U6854 ( .A1(\mem[349][1] ), .A2(n12419), .B1(n26781), .B2(
        data_in[1]), .ZN(n12420) );
  INV_X1 U6855 ( .A(n12421), .ZN(n23312) );
  AOI22_X1 U6856 ( .A1(\mem[349][2] ), .A2(n12419), .B1(n26781), .B2(
        data_in[2]), .ZN(n12421) );
  INV_X1 U6857 ( .A(n12422), .ZN(n23311) );
  AOI22_X1 U6858 ( .A1(\mem[349][3] ), .A2(n12419), .B1(n26781), .B2(
        data_in[3]), .ZN(n12422) );
  INV_X1 U6859 ( .A(n12423), .ZN(n23310) );
  AOI22_X1 U6860 ( .A1(\mem[349][4] ), .A2(n12419), .B1(n26781), .B2(
        data_in[4]), .ZN(n12423) );
  INV_X1 U6861 ( .A(n12424), .ZN(n23309) );
  AOI22_X1 U6862 ( .A1(\mem[349][5] ), .A2(n12419), .B1(n26781), .B2(
        data_in[5]), .ZN(n12424) );
  INV_X1 U6863 ( .A(n12425), .ZN(n23308) );
  AOI22_X1 U6864 ( .A1(\mem[349][6] ), .A2(n12419), .B1(n26781), .B2(
        data_in[6]), .ZN(n12425) );
  INV_X1 U6865 ( .A(n12426), .ZN(n23307) );
  AOI22_X1 U6866 ( .A1(\mem[349][7] ), .A2(n12419), .B1(n26781), .B2(
        data_in[7]), .ZN(n12426) );
  INV_X1 U6867 ( .A(n12427), .ZN(n23306) );
  AOI22_X1 U6868 ( .A1(\mem[350][0] ), .A2(n12428), .B1(n26780), .B2(
        data_in[0]), .ZN(n12427) );
  INV_X1 U6869 ( .A(n12429), .ZN(n23305) );
  AOI22_X1 U6870 ( .A1(\mem[350][1] ), .A2(n12428), .B1(n26780), .B2(
        data_in[1]), .ZN(n12429) );
  INV_X1 U6871 ( .A(n12430), .ZN(n23304) );
  AOI22_X1 U6872 ( .A1(\mem[350][2] ), .A2(n12428), .B1(n26780), .B2(
        data_in[2]), .ZN(n12430) );
  INV_X1 U6873 ( .A(n12431), .ZN(n23303) );
  AOI22_X1 U6874 ( .A1(\mem[350][3] ), .A2(n12428), .B1(n26780), .B2(
        data_in[3]), .ZN(n12431) );
  INV_X1 U6875 ( .A(n12432), .ZN(n23302) );
  AOI22_X1 U6876 ( .A1(\mem[350][4] ), .A2(n12428), .B1(n26780), .B2(
        data_in[4]), .ZN(n12432) );
  INV_X1 U6877 ( .A(n12433), .ZN(n23301) );
  AOI22_X1 U6878 ( .A1(\mem[350][5] ), .A2(n12428), .B1(n26780), .B2(
        data_in[5]), .ZN(n12433) );
  INV_X1 U6879 ( .A(n12434), .ZN(n23300) );
  AOI22_X1 U6880 ( .A1(\mem[350][6] ), .A2(n12428), .B1(n26780), .B2(
        data_in[6]), .ZN(n12434) );
  INV_X1 U6881 ( .A(n12435), .ZN(n23299) );
  AOI22_X1 U6882 ( .A1(\mem[350][7] ), .A2(n12428), .B1(n26780), .B2(
        data_in[7]), .ZN(n12435) );
  INV_X1 U6883 ( .A(n12436), .ZN(n23298) );
  AOI22_X1 U6884 ( .A1(\mem[351][0] ), .A2(n12437), .B1(n26779), .B2(
        data_in[0]), .ZN(n12436) );
  INV_X1 U6885 ( .A(n12438), .ZN(n23297) );
  AOI22_X1 U6886 ( .A1(\mem[351][1] ), .A2(n12437), .B1(n26779), .B2(
        data_in[1]), .ZN(n12438) );
  INV_X1 U6887 ( .A(n12439), .ZN(n23296) );
  AOI22_X1 U6888 ( .A1(\mem[351][2] ), .A2(n12437), .B1(n26779), .B2(
        data_in[2]), .ZN(n12439) );
  INV_X1 U6889 ( .A(n12440), .ZN(n23295) );
  AOI22_X1 U6890 ( .A1(\mem[351][3] ), .A2(n12437), .B1(n26779), .B2(
        data_in[3]), .ZN(n12440) );
  INV_X1 U6891 ( .A(n12441), .ZN(n23294) );
  AOI22_X1 U6892 ( .A1(\mem[351][4] ), .A2(n12437), .B1(n26779), .B2(
        data_in[4]), .ZN(n12441) );
  INV_X1 U6893 ( .A(n12442), .ZN(n23293) );
  AOI22_X1 U6894 ( .A1(\mem[351][5] ), .A2(n12437), .B1(n26779), .B2(
        data_in[5]), .ZN(n12442) );
  INV_X1 U6895 ( .A(n12443), .ZN(n23292) );
  AOI22_X1 U6896 ( .A1(\mem[351][6] ), .A2(n12437), .B1(n26779), .B2(
        data_in[6]), .ZN(n12443) );
  INV_X1 U6897 ( .A(n12444), .ZN(n23291) );
  AOI22_X1 U6898 ( .A1(\mem[351][7] ), .A2(n12437), .B1(n26779), .B2(
        data_in[7]), .ZN(n12444) );
  INV_X1 U6899 ( .A(n12518), .ZN(n23226) );
  AOI22_X1 U6900 ( .A1(\mem[360][0] ), .A2(n12519), .B1(n26770), .B2(
        data_in[0]), .ZN(n12518) );
  INV_X1 U6901 ( .A(n12520), .ZN(n23225) );
  AOI22_X1 U6902 ( .A1(\mem[360][1] ), .A2(n12519), .B1(n26770), .B2(
        data_in[1]), .ZN(n12520) );
  INV_X1 U6903 ( .A(n12521), .ZN(n23224) );
  AOI22_X1 U6904 ( .A1(\mem[360][2] ), .A2(n12519), .B1(n26770), .B2(
        data_in[2]), .ZN(n12521) );
  INV_X1 U6905 ( .A(n12522), .ZN(n23223) );
  AOI22_X1 U6906 ( .A1(\mem[360][3] ), .A2(n12519), .B1(n26770), .B2(
        data_in[3]), .ZN(n12522) );
  INV_X1 U6907 ( .A(n12523), .ZN(n23222) );
  AOI22_X1 U6908 ( .A1(\mem[360][4] ), .A2(n12519), .B1(n26770), .B2(
        data_in[4]), .ZN(n12523) );
  INV_X1 U6909 ( .A(n12524), .ZN(n23221) );
  AOI22_X1 U6910 ( .A1(\mem[360][5] ), .A2(n12519), .B1(n26770), .B2(
        data_in[5]), .ZN(n12524) );
  INV_X1 U6911 ( .A(n12525), .ZN(n23220) );
  AOI22_X1 U6912 ( .A1(\mem[360][6] ), .A2(n12519), .B1(n26770), .B2(
        data_in[6]), .ZN(n12525) );
  INV_X1 U6913 ( .A(n12526), .ZN(n23219) );
  AOI22_X1 U6914 ( .A1(\mem[360][7] ), .A2(n12519), .B1(n26770), .B2(
        data_in[7]), .ZN(n12526) );
  INV_X1 U6915 ( .A(n12527), .ZN(n23218) );
  AOI22_X1 U6916 ( .A1(\mem[361][0] ), .A2(n12528), .B1(n26769), .B2(
        data_in[0]), .ZN(n12527) );
  INV_X1 U6917 ( .A(n12529), .ZN(n23217) );
  AOI22_X1 U6918 ( .A1(\mem[361][1] ), .A2(n12528), .B1(n26769), .B2(
        data_in[1]), .ZN(n12529) );
  INV_X1 U6919 ( .A(n12530), .ZN(n23216) );
  AOI22_X1 U6920 ( .A1(\mem[361][2] ), .A2(n12528), .B1(n26769), .B2(
        data_in[2]), .ZN(n12530) );
  INV_X1 U6921 ( .A(n12531), .ZN(n23215) );
  AOI22_X1 U6922 ( .A1(\mem[361][3] ), .A2(n12528), .B1(n26769), .B2(
        data_in[3]), .ZN(n12531) );
  INV_X1 U6923 ( .A(n12532), .ZN(n23214) );
  AOI22_X1 U6924 ( .A1(\mem[361][4] ), .A2(n12528), .B1(n26769), .B2(
        data_in[4]), .ZN(n12532) );
  INV_X1 U6925 ( .A(n12533), .ZN(n23213) );
  AOI22_X1 U6926 ( .A1(\mem[361][5] ), .A2(n12528), .B1(n26769), .B2(
        data_in[5]), .ZN(n12533) );
  INV_X1 U6927 ( .A(n12534), .ZN(n23212) );
  AOI22_X1 U6928 ( .A1(\mem[361][6] ), .A2(n12528), .B1(n26769), .B2(
        data_in[6]), .ZN(n12534) );
  INV_X1 U6929 ( .A(n12535), .ZN(n23211) );
  AOI22_X1 U6930 ( .A1(\mem[361][7] ), .A2(n12528), .B1(n26769), .B2(
        data_in[7]), .ZN(n12535) );
  INV_X1 U6931 ( .A(n12536), .ZN(n23210) );
  AOI22_X1 U6932 ( .A1(\mem[362][0] ), .A2(n12537), .B1(n26768), .B2(
        data_in[0]), .ZN(n12536) );
  INV_X1 U6933 ( .A(n12538), .ZN(n23209) );
  AOI22_X1 U6934 ( .A1(\mem[362][1] ), .A2(n12537), .B1(n26768), .B2(
        data_in[1]), .ZN(n12538) );
  INV_X1 U6935 ( .A(n12539), .ZN(n23208) );
  AOI22_X1 U6936 ( .A1(\mem[362][2] ), .A2(n12537), .B1(n26768), .B2(
        data_in[2]), .ZN(n12539) );
  INV_X1 U6937 ( .A(n12540), .ZN(n23207) );
  AOI22_X1 U6938 ( .A1(\mem[362][3] ), .A2(n12537), .B1(n26768), .B2(
        data_in[3]), .ZN(n12540) );
  INV_X1 U6939 ( .A(n12541), .ZN(n23206) );
  AOI22_X1 U6940 ( .A1(\mem[362][4] ), .A2(n12537), .B1(n26768), .B2(
        data_in[4]), .ZN(n12541) );
  INV_X1 U6941 ( .A(n12542), .ZN(n23205) );
  AOI22_X1 U6942 ( .A1(\mem[362][5] ), .A2(n12537), .B1(n26768), .B2(
        data_in[5]), .ZN(n12542) );
  INV_X1 U6943 ( .A(n12543), .ZN(n23204) );
  AOI22_X1 U6944 ( .A1(\mem[362][6] ), .A2(n12537), .B1(n26768), .B2(
        data_in[6]), .ZN(n12543) );
  INV_X1 U6945 ( .A(n12544), .ZN(n23203) );
  AOI22_X1 U6946 ( .A1(\mem[362][7] ), .A2(n12537), .B1(n26768), .B2(
        data_in[7]), .ZN(n12544) );
  INV_X1 U6947 ( .A(n12545), .ZN(n23202) );
  AOI22_X1 U6948 ( .A1(\mem[363][0] ), .A2(n12546), .B1(n26767), .B2(
        data_in[0]), .ZN(n12545) );
  INV_X1 U6949 ( .A(n12547), .ZN(n23201) );
  AOI22_X1 U6950 ( .A1(\mem[363][1] ), .A2(n12546), .B1(n26767), .B2(
        data_in[1]), .ZN(n12547) );
  INV_X1 U6951 ( .A(n12548), .ZN(n23200) );
  AOI22_X1 U6952 ( .A1(\mem[363][2] ), .A2(n12546), .B1(n26767), .B2(
        data_in[2]), .ZN(n12548) );
  INV_X1 U6953 ( .A(n12549), .ZN(n23199) );
  AOI22_X1 U6954 ( .A1(\mem[363][3] ), .A2(n12546), .B1(n26767), .B2(
        data_in[3]), .ZN(n12549) );
  INV_X1 U6955 ( .A(n12550), .ZN(n23198) );
  AOI22_X1 U6956 ( .A1(\mem[363][4] ), .A2(n12546), .B1(n26767), .B2(
        data_in[4]), .ZN(n12550) );
  INV_X1 U6957 ( .A(n12551), .ZN(n23197) );
  AOI22_X1 U6958 ( .A1(\mem[363][5] ), .A2(n12546), .B1(n26767), .B2(
        data_in[5]), .ZN(n12551) );
  INV_X1 U6959 ( .A(n12552), .ZN(n23196) );
  AOI22_X1 U6960 ( .A1(\mem[363][6] ), .A2(n12546), .B1(n26767), .B2(
        data_in[6]), .ZN(n12552) );
  INV_X1 U6961 ( .A(n12553), .ZN(n23195) );
  AOI22_X1 U6962 ( .A1(\mem[363][7] ), .A2(n12546), .B1(n26767), .B2(
        data_in[7]), .ZN(n12553) );
  INV_X1 U6963 ( .A(n12554), .ZN(n23194) );
  AOI22_X1 U6964 ( .A1(\mem[364][0] ), .A2(n12555), .B1(n26766), .B2(
        data_in[0]), .ZN(n12554) );
  INV_X1 U6965 ( .A(n12556), .ZN(n23193) );
  AOI22_X1 U6966 ( .A1(\mem[364][1] ), .A2(n12555), .B1(n26766), .B2(
        data_in[1]), .ZN(n12556) );
  INV_X1 U6967 ( .A(n12557), .ZN(n23192) );
  AOI22_X1 U6968 ( .A1(\mem[364][2] ), .A2(n12555), .B1(n26766), .B2(
        data_in[2]), .ZN(n12557) );
  INV_X1 U6969 ( .A(n12558), .ZN(n23191) );
  AOI22_X1 U6970 ( .A1(\mem[364][3] ), .A2(n12555), .B1(n26766), .B2(
        data_in[3]), .ZN(n12558) );
  INV_X1 U6971 ( .A(n12559), .ZN(n23190) );
  AOI22_X1 U6972 ( .A1(\mem[364][4] ), .A2(n12555), .B1(n26766), .B2(
        data_in[4]), .ZN(n12559) );
  INV_X1 U6973 ( .A(n12560), .ZN(n23189) );
  AOI22_X1 U6974 ( .A1(\mem[364][5] ), .A2(n12555), .B1(n26766), .B2(
        data_in[5]), .ZN(n12560) );
  INV_X1 U6975 ( .A(n12561), .ZN(n23188) );
  AOI22_X1 U6976 ( .A1(\mem[364][6] ), .A2(n12555), .B1(n26766), .B2(
        data_in[6]), .ZN(n12561) );
  INV_X1 U6977 ( .A(n12562), .ZN(n23187) );
  AOI22_X1 U6978 ( .A1(\mem[364][7] ), .A2(n12555), .B1(n26766), .B2(
        data_in[7]), .ZN(n12562) );
  INV_X1 U6979 ( .A(n12563), .ZN(n23186) );
  AOI22_X1 U6980 ( .A1(\mem[365][0] ), .A2(n12564), .B1(n26765), .B2(
        data_in[0]), .ZN(n12563) );
  INV_X1 U6981 ( .A(n12565), .ZN(n23185) );
  AOI22_X1 U6982 ( .A1(\mem[365][1] ), .A2(n12564), .B1(n26765), .B2(
        data_in[1]), .ZN(n12565) );
  INV_X1 U6983 ( .A(n12566), .ZN(n23184) );
  AOI22_X1 U6984 ( .A1(\mem[365][2] ), .A2(n12564), .B1(n26765), .B2(
        data_in[2]), .ZN(n12566) );
  INV_X1 U6985 ( .A(n12567), .ZN(n23183) );
  AOI22_X1 U6986 ( .A1(\mem[365][3] ), .A2(n12564), .B1(n26765), .B2(
        data_in[3]), .ZN(n12567) );
  INV_X1 U6987 ( .A(n12568), .ZN(n23182) );
  AOI22_X1 U6988 ( .A1(\mem[365][4] ), .A2(n12564), .B1(n26765), .B2(
        data_in[4]), .ZN(n12568) );
  INV_X1 U6989 ( .A(n12569), .ZN(n23181) );
  AOI22_X1 U6990 ( .A1(\mem[365][5] ), .A2(n12564), .B1(n26765), .B2(
        data_in[5]), .ZN(n12569) );
  INV_X1 U6991 ( .A(n12570), .ZN(n23180) );
  AOI22_X1 U6992 ( .A1(\mem[365][6] ), .A2(n12564), .B1(n26765), .B2(
        data_in[6]), .ZN(n12570) );
  INV_X1 U6993 ( .A(n12571), .ZN(n23179) );
  AOI22_X1 U6994 ( .A1(\mem[365][7] ), .A2(n12564), .B1(n26765), .B2(
        data_in[7]), .ZN(n12571) );
  INV_X1 U6995 ( .A(n12572), .ZN(n23178) );
  AOI22_X1 U6996 ( .A1(\mem[366][0] ), .A2(n12573), .B1(n26764), .B2(
        data_in[0]), .ZN(n12572) );
  INV_X1 U6997 ( .A(n12574), .ZN(n23177) );
  AOI22_X1 U6998 ( .A1(\mem[366][1] ), .A2(n12573), .B1(n26764), .B2(
        data_in[1]), .ZN(n12574) );
  INV_X1 U6999 ( .A(n12575), .ZN(n23176) );
  AOI22_X1 U7000 ( .A1(\mem[366][2] ), .A2(n12573), .B1(n26764), .B2(
        data_in[2]), .ZN(n12575) );
  INV_X1 U7001 ( .A(n12576), .ZN(n23175) );
  AOI22_X1 U7002 ( .A1(\mem[366][3] ), .A2(n12573), .B1(n26764), .B2(
        data_in[3]), .ZN(n12576) );
  INV_X1 U7003 ( .A(n12577), .ZN(n23174) );
  AOI22_X1 U7004 ( .A1(\mem[366][4] ), .A2(n12573), .B1(n26764), .B2(
        data_in[4]), .ZN(n12577) );
  INV_X1 U7005 ( .A(n12578), .ZN(n23173) );
  AOI22_X1 U7006 ( .A1(\mem[366][5] ), .A2(n12573), .B1(n26764), .B2(
        data_in[5]), .ZN(n12578) );
  INV_X1 U7007 ( .A(n12579), .ZN(n23172) );
  AOI22_X1 U7008 ( .A1(\mem[366][6] ), .A2(n12573), .B1(n26764), .B2(
        data_in[6]), .ZN(n12579) );
  INV_X1 U7009 ( .A(n12580), .ZN(n23171) );
  AOI22_X1 U7010 ( .A1(\mem[366][7] ), .A2(n12573), .B1(n26764), .B2(
        data_in[7]), .ZN(n12580) );
  INV_X1 U7011 ( .A(n12581), .ZN(n23170) );
  AOI22_X1 U7012 ( .A1(\mem[367][0] ), .A2(n12582), .B1(n26763), .B2(
        data_in[0]), .ZN(n12581) );
  INV_X1 U7013 ( .A(n12583), .ZN(n23169) );
  AOI22_X1 U7014 ( .A1(\mem[367][1] ), .A2(n12582), .B1(n26763), .B2(
        data_in[1]), .ZN(n12583) );
  INV_X1 U7015 ( .A(n12584), .ZN(n23168) );
  AOI22_X1 U7016 ( .A1(\mem[367][2] ), .A2(n12582), .B1(n26763), .B2(
        data_in[2]), .ZN(n12584) );
  INV_X1 U7017 ( .A(n12585), .ZN(n23167) );
  AOI22_X1 U7018 ( .A1(\mem[367][3] ), .A2(n12582), .B1(n26763), .B2(
        data_in[3]), .ZN(n12585) );
  INV_X1 U7019 ( .A(n12586), .ZN(n23166) );
  AOI22_X1 U7020 ( .A1(\mem[367][4] ), .A2(n12582), .B1(n26763), .B2(
        data_in[4]), .ZN(n12586) );
  INV_X1 U7021 ( .A(n12587), .ZN(n23165) );
  AOI22_X1 U7022 ( .A1(\mem[367][5] ), .A2(n12582), .B1(n26763), .B2(
        data_in[5]), .ZN(n12587) );
  INV_X1 U7023 ( .A(n12588), .ZN(n23164) );
  AOI22_X1 U7024 ( .A1(\mem[367][6] ), .A2(n12582), .B1(n26763), .B2(
        data_in[6]), .ZN(n12588) );
  INV_X1 U7025 ( .A(n12589), .ZN(n23163) );
  AOI22_X1 U7026 ( .A1(\mem[367][7] ), .A2(n12582), .B1(n26763), .B2(
        data_in[7]), .ZN(n12589) );
  INV_X1 U7027 ( .A(n12590), .ZN(n23162) );
  AOI22_X1 U7028 ( .A1(\mem[368][0] ), .A2(n12591), .B1(n26762), .B2(
        data_in[0]), .ZN(n12590) );
  INV_X1 U7029 ( .A(n12592), .ZN(n23161) );
  AOI22_X1 U7030 ( .A1(\mem[368][1] ), .A2(n12591), .B1(n26762), .B2(
        data_in[1]), .ZN(n12592) );
  INV_X1 U7031 ( .A(n12593), .ZN(n23160) );
  AOI22_X1 U7032 ( .A1(\mem[368][2] ), .A2(n12591), .B1(n26762), .B2(
        data_in[2]), .ZN(n12593) );
  INV_X1 U7033 ( .A(n12594), .ZN(n23159) );
  AOI22_X1 U7034 ( .A1(\mem[368][3] ), .A2(n12591), .B1(n26762), .B2(
        data_in[3]), .ZN(n12594) );
  INV_X1 U7035 ( .A(n12595), .ZN(n23158) );
  AOI22_X1 U7036 ( .A1(\mem[368][4] ), .A2(n12591), .B1(n26762), .B2(
        data_in[4]), .ZN(n12595) );
  INV_X1 U7037 ( .A(n12596), .ZN(n23157) );
  AOI22_X1 U7038 ( .A1(\mem[368][5] ), .A2(n12591), .B1(n26762), .B2(
        data_in[5]), .ZN(n12596) );
  INV_X1 U7039 ( .A(n12597), .ZN(n23156) );
  AOI22_X1 U7040 ( .A1(\mem[368][6] ), .A2(n12591), .B1(n26762), .B2(
        data_in[6]), .ZN(n12597) );
  INV_X1 U7041 ( .A(n12598), .ZN(n23155) );
  AOI22_X1 U7042 ( .A1(\mem[368][7] ), .A2(n12591), .B1(n26762), .B2(
        data_in[7]), .ZN(n12598) );
  INV_X1 U7043 ( .A(n12599), .ZN(n23154) );
  AOI22_X1 U7044 ( .A1(\mem[369][0] ), .A2(n12600), .B1(n26761), .B2(
        data_in[0]), .ZN(n12599) );
  INV_X1 U7045 ( .A(n12601), .ZN(n23153) );
  AOI22_X1 U7046 ( .A1(\mem[369][1] ), .A2(n12600), .B1(n26761), .B2(
        data_in[1]), .ZN(n12601) );
  INV_X1 U7047 ( .A(n12602), .ZN(n23152) );
  AOI22_X1 U7048 ( .A1(\mem[369][2] ), .A2(n12600), .B1(n26761), .B2(
        data_in[2]), .ZN(n12602) );
  INV_X1 U7049 ( .A(n12603), .ZN(n23151) );
  AOI22_X1 U7050 ( .A1(\mem[369][3] ), .A2(n12600), .B1(n26761), .B2(
        data_in[3]), .ZN(n12603) );
  INV_X1 U7051 ( .A(n12604), .ZN(n23150) );
  AOI22_X1 U7052 ( .A1(\mem[369][4] ), .A2(n12600), .B1(n26761), .B2(
        data_in[4]), .ZN(n12604) );
  INV_X1 U7053 ( .A(n12605), .ZN(n23149) );
  AOI22_X1 U7054 ( .A1(\mem[369][5] ), .A2(n12600), .B1(n26761), .B2(
        data_in[5]), .ZN(n12605) );
  INV_X1 U7055 ( .A(n12606), .ZN(n23148) );
  AOI22_X1 U7056 ( .A1(\mem[369][6] ), .A2(n12600), .B1(n26761), .B2(
        data_in[6]), .ZN(n12606) );
  INV_X1 U7057 ( .A(n12607), .ZN(n23147) );
  AOI22_X1 U7058 ( .A1(\mem[369][7] ), .A2(n12600), .B1(n26761), .B2(
        data_in[7]), .ZN(n12607) );
  INV_X1 U7059 ( .A(n12608), .ZN(n23146) );
  AOI22_X1 U7060 ( .A1(\mem[370][0] ), .A2(n12609), .B1(n26760), .B2(
        data_in[0]), .ZN(n12608) );
  INV_X1 U7061 ( .A(n12610), .ZN(n23145) );
  AOI22_X1 U7062 ( .A1(\mem[370][1] ), .A2(n12609), .B1(n26760), .B2(
        data_in[1]), .ZN(n12610) );
  INV_X1 U7063 ( .A(n12611), .ZN(n23144) );
  AOI22_X1 U7064 ( .A1(\mem[370][2] ), .A2(n12609), .B1(n26760), .B2(
        data_in[2]), .ZN(n12611) );
  INV_X1 U7065 ( .A(n12612), .ZN(n23143) );
  AOI22_X1 U7066 ( .A1(\mem[370][3] ), .A2(n12609), .B1(n26760), .B2(
        data_in[3]), .ZN(n12612) );
  INV_X1 U7067 ( .A(n12613), .ZN(n23142) );
  AOI22_X1 U7068 ( .A1(\mem[370][4] ), .A2(n12609), .B1(n26760), .B2(
        data_in[4]), .ZN(n12613) );
  INV_X1 U7069 ( .A(n12614), .ZN(n23141) );
  AOI22_X1 U7070 ( .A1(\mem[370][5] ), .A2(n12609), .B1(n26760), .B2(
        data_in[5]), .ZN(n12614) );
  INV_X1 U7071 ( .A(n12615), .ZN(n23140) );
  AOI22_X1 U7072 ( .A1(\mem[370][6] ), .A2(n12609), .B1(n26760), .B2(
        data_in[6]), .ZN(n12615) );
  INV_X1 U7073 ( .A(n12616), .ZN(n23139) );
  AOI22_X1 U7074 ( .A1(\mem[370][7] ), .A2(n12609), .B1(n26760), .B2(
        data_in[7]), .ZN(n12616) );
  INV_X1 U7075 ( .A(n12617), .ZN(n23138) );
  AOI22_X1 U7076 ( .A1(\mem[371][0] ), .A2(n12618), .B1(n26759), .B2(
        data_in[0]), .ZN(n12617) );
  INV_X1 U7077 ( .A(n12619), .ZN(n23137) );
  AOI22_X1 U7078 ( .A1(\mem[371][1] ), .A2(n12618), .B1(n26759), .B2(
        data_in[1]), .ZN(n12619) );
  INV_X1 U7079 ( .A(n12620), .ZN(n23136) );
  AOI22_X1 U7080 ( .A1(\mem[371][2] ), .A2(n12618), .B1(n26759), .B2(
        data_in[2]), .ZN(n12620) );
  INV_X1 U7081 ( .A(n12621), .ZN(n23135) );
  AOI22_X1 U7082 ( .A1(\mem[371][3] ), .A2(n12618), .B1(n26759), .B2(
        data_in[3]), .ZN(n12621) );
  INV_X1 U7083 ( .A(n12622), .ZN(n23134) );
  AOI22_X1 U7084 ( .A1(\mem[371][4] ), .A2(n12618), .B1(n26759), .B2(
        data_in[4]), .ZN(n12622) );
  INV_X1 U7085 ( .A(n12623), .ZN(n23133) );
  AOI22_X1 U7086 ( .A1(\mem[371][5] ), .A2(n12618), .B1(n26759), .B2(
        data_in[5]), .ZN(n12623) );
  INV_X1 U7087 ( .A(n12624), .ZN(n23132) );
  AOI22_X1 U7088 ( .A1(\mem[371][6] ), .A2(n12618), .B1(n26759), .B2(
        data_in[6]), .ZN(n12624) );
  INV_X1 U7089 ( .A(n12625), .ZN(n23131) );
  AOI22_X1 U7090 ( .A1(\mem[371][7] ), .A2(n12618), .B1(n26759), .B2(
        data_in[7]), .ZN(n12625) );
  INV_X1 U7091 ( .A(n12626), .ZN(n23130) );
  AOI22_X1 U7092 ( .A1(\mem[372][0] ), .A2(n12627), .B1(n26758), .B2(
        data_in[0]), .ZN(n12626) );
  INV_X1 U7093 ( .A(n12628), .ZN(n23129) );
  AOI22_X1 U7094 ( .A1(\mem[372][1] ), .A2(n12627), .B1(n26758), .B2(
        data_in[1]), .ZN(n12628) );
  INV_X1 U7095 ( .A(n12629), .ZN(n23128) );
  AOI22_X1 U7096 ( .A1(\mem[372][2] ), .A2(n12627), .B1(n26758), .B2(
        data_in[2]), .ZN(n12629) );
  INV_X1 U7097 ( .A(n12630), .ZN(n23127) );
  AOI22_X1 U7098 ( .A1(\mem[372][3] ), .A2(n12627), .B1(n26758), .B2(
        data_in[3]), .ZN(n12630) );
  INV_X1 U7099 ( .A(n12631), .ZN(n23126) );
  AOI22_X1 U7100 ( .A1(\mem[372][4] ), .A2(n12627), .B1(n26758), .B2(
        data_in[4]), .ZN(n12631) );
  INV_X1 U7101 ( .A(n12632), .ZN(n23125) );
  AOI22_X1 U7102 ( .A1(\mem[372][5] ), .A2(n12627), .B1(n26758), .B2(
        data_in[5]), .ZN(n12632) );
  INV_X1 U7103 ( .A(n12633), .ZN(n23124) );
  AOI22_X1 U7104 ( .A1(\mem[372][6] ), .A2(n12627), .B1(n26758), .B2(
        data_in[6]), .ZN(n12633) );
  INV_X1 U7105 ( .A(n12634), .ZN(n23123) );
  AOI22_X1 U7106 ( .A1(\mem[372][7] ), .A2(n12627), .B1(n26758), .B2(
        data_in[7]), .ZN(n12634) );
  INV_X1 U7107 ( .A(n12635), .ZN(n23122) );
  AOI22_X1 U7108 ( .A1(\mem[373][0] ), .A2(n12636), .B1(n26757), .B2(
        data_in[0]), .ZN(n12635) );
  INV_X1 U7109 ( .A(n12637), .ZN(n23121) );
  AOI22_X1 U7110 ( .A1(\mem[373][1] ), .A2(n12636), .B1(n26757), .B2(
        data_in[1]), .ZN(n12637) );
  INV_X1 U7111 ( .A(n12638), .ZN(n23120) );
  AOI22_X1 U7112 ( .A1(\mem[373][2] ), .A2(n12636), .B1(n26757), .B2(
        data_in[2]), .ZN(n12638) );
  INV_X1 U7113 ( .A(n12639), .ZN(n23119) );
  AOI22_X1 U7114 ( .A1(\mem[373][3] ), .A2(n12636), .B1(n26757), .B2(
        data_in[3]), .ZN(n12639) );
  INV_X1 U7115 ( .A(n12640), .ZN(n23118) );
  AOI22_X1 U7116 ( .A1(\mem[373][4] ), .A2(n12636), .B1(n26757), .B2(
        data_in[4]), .ZN(n12640) );
  INV_X1 U7117 ( .A(n12641), .ZN(n23117) );
  AOI22_X1 U7118 ( .A1(\mem[373][5] ), .A2(n12636), .B1(n26757), .B2(
        data_in[5]), .ZN(n12641) );
  INV_X1 U7119 ( .A(n12642), .ZN(n23116) );
  AOI22_X1 U7120 ( .A1(\mem[373][6] ), .A2(n12636), .B1(n26757), .B2(
        data_in[6]), .ZN(n12642) );
  INV_X1 U7121 ( .A(n12643), .ZN(n23115) );
  AOI22_X1 U7122 ( .A1(\mem[373][7] ), .A2(n12636), .B1(n26757), .B2(
        data_in[7]), .ZN(n12643) );
  INV_X1 U7123 ( .A(n12644), .ZN(n23114) );
  AOI22_X1 U7124 ( .A1(\mem[374][0] ), .A2(n12645), .B1(n26756), .B2(
        data_in[0]), .ZN(n12644) );
  INV_X1 U7125 ( .A(n12646), .ZN(n23113) );
  AOI22_X1 U7126 ( .A1(\mem[374][1] ), .A2(n12645), .B1(n26756), .B2(
        data_in[1]), .ZN(n12646) );
  INV_X1 U7127 ( .A(n12647), .ZN(n23112) );
  AOI22_X1 U7128 ( .A1(\mem[374][2] ), .A2(n12645), .B1(n26756), .B2(
        data_in[2]), .ZN(n12647) );
  INV_X1 U7129 ( .A(n12648), .ZN(n23111) );
  AOI22_X1 U7130 ( .A1(\mem[374][3] ), .A2(n12645), .B1(n26756), .B2(
        data_in[3]), .ZN(n12648) );
  INV_X1 U7131 ( .A(n12649), .ZN(n23110) );
  AOI22_X1 U7132 ( .A1(\mem[374][4] ), .A2(n12645), .B1(n26756), .B2(
        data_in[4]), .ZN(n12649) );
  INV_X1 U7133 ( .A(n12650), .ZN(n23109) );
  AOI22_X1 U7134 ( .A1(\mem[374][5] ), .A2(n12645), .B1(n26756), .B2(
        data_in[5]), .ZN(n12650) );
  INV_X1 U7135 ( .A(n12651), .ZN(n23108) );
  AOI22_X1 U7136 ( .A1(\mem[374][6] ), .A2(n12645), .B1(n26756), .B2(
        data_in[6]), .ZN(n12651) );
  INV_X1 U7137 ( .A(n12652), .ZN(n23107) );
  AOI22_X1 U7138 ( .A1(\mem[374][7] ), .A2(n12645), .B1(n26756), .B2(
        data_in[7]), .ZN(n12652) );
  INV_X1 U7139 ( .A(n12653), .ZN(n23106) );
  AOI22_X1 U7140 ( .A1(\mem[375][0] ), .A2(n12654), .B1(n26755), .B2(
        data_in[0]), .ZN(n12653) );
  INV_X1 U7141 ( .A(n12655), .ZN(n23105) );
  AOI22_X1 U7142 ( .A1(\mem[375][1] ), .A2(n12654), .B1(n26755), .B2(
        data_in[1]), .ZN(n12655) );
  INV_X1 U7143 ( .A(n12656), .ZN(n23104) );
  AOI22_X1 U7144 ( .A1(\mem[375][2] ), .A2(n12654), .B1(n26755), .B2(
        data_in[2]), .ZN(n12656) );
  INV_X1 U7145 ( .A(n12657), .ZN(n23103) );
  AOI22_X1 U7146 ( .A1(\mem[375][3] ), .A2(n12654), .B1(n26755), .B2(
        data_in[3]), .ZN(n12657) );
  INV_X1 U7147 ( .A(n12658), .ZN(n23102) );
  AOI22_X1 U7148 ( .A1(\mem[375][4] ), .A2(n12654), .B1(n26755), .B2(
        data_in[4]), .ZN(n12658) );
  INV_X1 U7149 ( .A(n12659), .ZN(n23101) );
  AOI22_X1 U7150 ( .A1(\mem[375][5] ), .A2(n12654), .B1(n26755), .B2(
        data_in[5]), .ZN(n12659) );
  INV_X1 U7151 ( .A(n12660), .ZN(n23100) );
  AOI22_X1 U7152 ( .A1(\mem[375][6] ), .A2(n12654), .B1(n26755), .B2(
        data_in[6]), .ZN(n12660) );
  INV_X1 U7153 ( .A(n12661), .ZN(n23099) );
  AOI22_X1 U7154 ( .A1(\mem[375][7] ), .A2(n12654), .B1(n26755), .B2(
        data_in[7]), .ZN(n12661) );
  INV_X1 U7155 ( .A(n12662), .ZN(n23098) );
  AOI22_X1 U7156 ( .A1(\mem[376][0] ), .A2(n12663), .B1(n26754), .B2(
        data_in[0]), .ZN(n12662) );
  INV_X1 U7157 ( .A(n12664), .ZN(n23097) );
  AOI22_X1 U7158 ( .A1(\mem[376][1] ), .A2(n12663), .B1(n26754), .B2(
        data_in[1]), .ZN(n12664) );
  INV_X1 U7159 ( .A(n12665), .ZN(n23096) );
  AOI22_X1 U7160 ( .A1(\mem[376][2] ), .A2(n12663), .B1(n26754), .B2(
        data_in[2]), .ZN(n12665) );
  INV_X1 U7161 ( .A(n12666), .ZN(n23095) );
  AOI22_X1 U7162 ( .A1(\mem[376][3] ), .A2(n12663), .B1(n26754), .B2(
        data_in[3]), .ZN(n12666) );
  INV_X1 U7163 ( .A(n12667), .ZN(n23094) );
  AOI22_X1 U7164 ( .A1(\mem[376][4] ), .A2(n12663), .B1(n26754), .B2(
        data_in[4]), .ZN(n12667) );
  INV_X1 U7165 ( .A(n12668), .ZN(n23093) );
  AOI22_X1 U7166 ( .A1(\mem[376][5] ), .A2(n12663), .B1(n26754), .B2(
        data_in[5]), .ZN(n12668) );
  INV_X1 U7167 ( .A(n12669), .ZN(n23092) );
  AOI22_X1 U7168 ( .A1(\mem[376][6] ), .A2(n12663), .B1(n26754), .B2(
        data_in[6]), .ZN(n12669) );
  INV_X1 U7169 ( .A(n12670), .ZN(n23091) );
  AOI22_X1 U7170 ( .A1(\mem[376][7] ), .A2(n12663), .B1(n26754), .B2(
        data_in[7]), .ZN(n12670) );
  INV_X1 U7171 ( .A(n12671), .ZN(n23090) );
  AOI22_X1 U7172 ( .A1(\mem[377][0] ), .A2(n12672), .B1(n26753), .B2(
        data_in[0]), .ZN(n12671) );
  INV_X1 U7173 ( .A(n12673), .ZN(n23089) );
  AOI22_X1 U7174 ( .A1(\mem[377][1] ), .A2(n12672), .B1(n26753), .B2(
        data_in[1]), .ZN(n12673) );
  INV_X1 U7175 ( .A(n12674), .ZN(n23088) );
  AOI22_X1 U7176 ( .A1(\mem[377][2] ), .A2(n12672), .B1(n26753), .B2(
        data_in[2]), .ZN(n12674) );
  INV_X1 U7177 ( .A(n12675), .ZN(n23087) );
  AOI22_X1 U7178 ( .A1(\mem[377][3] ), .A2(n12672), .B1(n26753), .B2(
        data_in[3]), .ZN(n12675) );
  INV_X1 U7179 ( .A(n12676), .ZN(n23086) );
  AOI22_X1 U7180 ( .A1(\mem[377][4] ), .A2(n12672), .B1(n26753), .B2(
        data_in[4]), .ZN(n12676) );
  INV_X1 U7181 ( .A(n12677), .ZN(n23085) );
  AOI22_X1 U7182 ( .A1(\mem[377][5] ), .A2(n12672), .B1(n26753), .B2(
        data_in[5]), .ZN(n12677) );
  INV_X1 U7183 ( .A(n12678), .ZN(n23084) );
  AOI22_X1 U7184 ( .A1(\mem[377][6] ), .A2(n12672), .B1(n26753), .B2(
        data_in[6]), .ZN(n12678) );
  INV_X1 U7185 ( .A(n12679), .ZN(n23083) );
  AOI22_X1 U7186 ( .A1(\mem[377][7] ), .A2(n12672), .B1(n26753), .B2(
        data_in[7]), .ZN(n12679) );
  INV_X1 U7187 ( .A(n12680), .ZN(n23082) );
  AOI22_X1 U7188 ( .A1(\mem[378][0] ), .A2(n12681), .B1(n26752), .B2(
        data_in[0]), .ZN(n12680) );
  INV_X1 U7189 ( .A(n12682), .ZN(n23081) );
  AOI22_X1 U7190 ( .A1(\mem[378][1] ), .A2(n12681), .B1(n26752), .B2(
        data_in[1]), .ZN(n12682) );
  INV_X1 U7191 ( .A(n12683), .ZN(n23080) );
  AOI22_X1 U7192 ( .A1(\mem[378][2] ), .A2(n12681), .B1(n26752), .B2(
        data_in[2]), .ZN(n12683) );
  INV_X1 U7193 ( .A(n12684), .ZN(n23079) );
  AOI22_X1 U7194 ( .A1(\mem[378][3] ), .A2(n12681), .B1(n26752), .B2(
        data_in[3]), .ZN(n12684) );
  INV_X1 U7195 ( .A(n12685), .ZN(n23078) );
  AOI22_X1 U7196 ( .A1(\mem[378][4] ), .A2(n12681), .B1(n26752), .B2(
        data_in[4]), .ZN(n12685) );
  INV_X1 U7197 ( .A(n12686), .ZN(n23077) );
  AOI22_X1 U7198 ( .A1(\mem[378][5] ), .A2(n12681), .B1(n26752), .B2(
        data_in[5]), .ZN(n12686) );
  INV_X1 U7199 ( .A(n12687), .ZN(n23076) );
  AOI22_X1 U7200 ( .A1(\mem[378][6] ), .A2(n12681), .B1(n26752), .B2(
        data_in[6]), .ZN(n12687) );
  INV_X1 U7201 ( .A(n12688), .ZN(n23075) );
  AOI22_X1 U7202 ( .A1(\mem[378][7] ), .A2(n12681), .B1(n26752), .B2(
        data_in[7]), .ZN(n12688) );
  INV_X1 U7203 ( .A(n12689), .ZN(n23074) );
  AOI22_X1 U7204 ( .A1(\mem[379][0] ), .A2(n12690), .B1(n26751), .B2(
        data_in[0]), .ZN(n12689) );
  INV_X1 U7205 ( .A(n12691), .ZN(n23073) );
  AOI22_X1 U7206 ( .A1(\mem[379][1] ), .A2(n12690), .B1(n26751), .B2(
        data_in[1]), .ZN(n12691) );
  INV_X1 U7207 ( .A(n12692), .ZN(n23072) );
  AOI22_X1 U7208 ( .A1(\mem[379][2] ), .A2(n12690), .B1(n26751), .B2(
        data_in[2]), .ZN(n12692) );
  INV_X1 U7209 ( .A(n12693), .ZN(n23071) );
  AOI22_X1 U7210 ( .A1(\mem[379][3] ), .A2(n12690), .B1(n26751), .B2(
        data_in[3]), .ZN(n12693) );
  INV_X1 U7211 ( .A(n12694), .ZN(n23070) );
  AOI22_X1 U7212 ( .A1(\mem[379][4] ), .A2(n12690), .B1(n26751), .B2(
        data_in[4]), .ZN(n12694) );
  INV_X1 U7213 ( .A(n12695), .ZN(n23069) );
  AOI22_X1 U7214 ( .A1(\mem[379][5] ), .A2(n12690), .B1(n26751), .B2(
        data_in[5]), .ZN(n12695) );
  INV_X1 U7215 ( .A(n12696), .ZN(n23068) );
  AOI22_X1 U7216 ( .A1(\mem[379][6] ), .A2(n12690), .B1(n26751), .B2(
        data_in[6]), .ZN(n12696) );
  INV_X1 U7217 ( .A(n12697), .ZN(n23067) );
  AOI22_X1 U7218 ( .A1(\mem[379][7] ), .A2(n12690), .B1(n26751), .B2(
        data_in[7]), .ZN(n12697) );
  INV_X1 U7219 ( .A(n12698), .ZN(n23066) );
  AOI22_X1 U7220 ( .A1(\mem[380][0] ), .A2(n12699), .B1(n26750), .B2(
        data_in[0]), .ZN(n12698) );
  INV_X1 U7221 ( .A(n12700), .ZN(n23065) );
  AOI22_X1 U7222 ( .A1(\mem[380][1] ), .A2(n12699), .B1(n26750), .B2(
        data_in[1]), .ZN(n12700) );
  INV_X1 U7223 ( .A(n12701), .ZN(n23064) );
  AOI22_X1 U7224 ( .A1(\mem[380][2] ), .A2(n12699), .B1(n26750), .B2(
        data_in[2]), .ZN(n12701) );
  INV_X1 U7225 ( .A(n12702), .ZN(n23063) );
  AOI22_X1 U7226 ( .A1(\mem[380][3] ), .A2(n12699), .B1(n26750), .B2(
        data_in[3]), .ZN(n12702) );
  INV_X1 U7227 ( .A(n12703), .ZN(n23062) );
  AOI22_X1 U7228 ( .A1(\mem[380][4] ), .A2(n12699), .B1(n26750), .B2(
        data_in[4]), .ZN(n12703) );
  INV_X1 U7229 ( .A(n12704), .ZN(n23061) );
  AOI22_X1 U7230 ( .A1(\mem[380][5] ), .A2(n12699), .B1(n26750), .B2(
        data_in[5]), .ZN(n12704) );
  INV_X1 U7231 ( .A(n12705), .ZN(n23060) );
  AOI22_X1 U7232 ( .A1(\mem[380][6] ), .A2(n12699), .B1(n26750), .B2(
        data_in[6]), .ZN(n12705) );
  INV_X1 U7233 ( .A(n12706), .ZN(n23059) );
  AOI22_X1 U7234 ( .A1(\mem[380][7] ), .A2(n12699), .B1(n26750), .B2(
        data_in[7]), .ZN(n12706) );
  INV_X1 U7235 ( .A(n12707), .ZN(n23058) );
  AOI22_X1 U7236 ( .A1(\mem[381][0] ), .A2(n12708), .B1(n26749), .B2(
        data_in[0]), .ZN(n12707) );
  INV_X1 U7237 ( .A(n12709), .ZN(n23057) );
  AOI22_X1 U7238 ( .A1(\mem[381][1] ), .A2(n12708), .B1(n26749), .B2(
        data_in[1]), .ZN(n12709) );
  INV_X1 U7239 ( .A(n12710), .ZN(n23056) );
  AOI22_X1 U7240 ( .A1(\mem[381][2] ), .A2(n12708), .B1(n26749), .B2(
        data_in[2]), .ZN(n12710) );
  INV_X1 U7241 ( .A(n12711), .ZN(n23055) );
  AOI22_X1 U7242 ( .A1(\mem[381][3] ), .A2(n12708), .B1(n26749), .B2(
        data_in[3]), .ZN(n12711) );
  INV_X1 U7243 ( .A(n12712), .ZN(n23054) );
  AOI22_X1 U7244 ( .A1(\mem[381][4] ), .A2(n12708), .B1(n26749), .B2(
        data_in[4]), .ZN(n12712) );
  INV_X1 U7245 ( .A(n12713), .ZN(n23053) );
  AOI22_X1 U7246 ( .A1(\mem[381][5] ), .A2(n12708), .B1(n26749), .B2(
        data_in[5]), .ZN(n12713) );
  INV_X1 U7247 ( .A(n12714), .ZN(n23052) );
  AOI22_X1 U7248 ( .A1(\mem[381][6] ), .A2(n12708), .B1(n26749), .B2(
        data_in[6]), .ZN(n12714) );
  INV_X1 U7249 ( .A(n12715), .ZN(n23051) );
  AOI22_X1 U7250 ( .A1(\mem[381][7] ), .A2(n12708), .B1(n26749), .B2(
        data_in[7]), .ZN(n12715) );
  INV_X1 U7251 ( .A(n12716), .ZN(n23050) );
  AOI22_X1 U7252 ( .A1(\mem[382][0] ), .A2(n12717), .B1(n26748), .B2(
        data_in[0]), .ZN(n12716) );
  INV_X1 U7253 ( .A(n12718), .ZN(n23049) );
  AOI22_X1 U7254 ( .A1(\mem[382][1] ), .A2(n12717), .B1(n26748), .B2(
        data_in[1]), .ZN(n12718) );
  INV_X1 U7255 ( .A(n12719), .ZN(n23048) );
  AOI22_X1 U7256 ( .A1(\mem[382][2] ), .A2(n12717), .B1(n26748), .B2(
        data_in[2]), .ZN(n12719) );
  INV_X1 U7257 ( .A(n12720), .ZN(n23047) );
  AOI22_X1 U7258 ( .A1(\mem[382][3] ), .A2(n12717), .B1(n26748), .B2(
        data_in[3]), .ZN(n12720) );
  INV_X1 U7259 ( .A(n12721), .ZN(n23046) );
  AOI22_X1 U7260 ( .A1(\mem[382][4] ), .A2(n12717), .B1(n26748), .B2(
        data_in[4]), .ZN(n12721) );
  INV_X1 U7261 ( .A(n12722), .ZN(n23045) );
  AOI22_X1 U7262 ( .A1(\mem[382][5] ), .A2(n12717), .B1(n26748), .B2(
        data_in[5]), .ZN(n12722) );
  INV_X1 U7263 ( .A(n12723), .ZN(n23044) );
  AOI22_X1 U7264 ( .A1(\mem[382][6] ), .A2(n12717), .B1(n26748), .B2(
        data_in[6]), .ZN(n12723) );
  INV_X1 U7265 ( .A(n12724), .ZN(n23043) );
  AOI22_X1 U7266 ( .A1(\mem[382][7] ), .A2(n12717), .B1(n26748), .B2(
        data_in[7]), .ZN(n12724) );
  INV_X1 U7267 ( .A(n12725), .ZN(n23042) );
  AOI22_X1 U7268 ( .A1(\mem[383][0] ), .A2(n12726), .B1(n26747), .B2(
        data_in[0]), .ZN(n12725) );
  INV_X1 U7269 ( .A(n12727), .ZN(n23041) );
  AOI22_X1 U7270 ( .A1(\mem[383][1] ), .A2(n12726), .B1(n26747), .B2(
        data_in[1]), .ZN(n12727) );
  INV_X1 U7271 ( .A(n12728), .ZN(n23040) );
  AOI22_X1 U7272 ( .A1(\mem[383][2] ), .A2(n12726), .B1(n26747), .B2(
        data_in[2]), .ZN(n12728) );
  INV_X1 U7273 ( .A(n12729), .ZN(n23039) );
  AOI22_X1 U7274 ( .A1(\mem[383][3] ), .A2(n12726), .B1(n26747), .B2(
        data_in[3]), .ZN(n12729) );
  INV_X1 U7275 ( .A(n12730), .ZN(n23038) );
  AOI22_X1 U7276 ( .A1(\mem[383][4] ), .A2(n12726), .B1(n26747), .B2(
        data_in[4]), .ZN(n12730) );
  INV_X1 U7277 ( .A(n12731), .ZN(n23037) );
  AOI22_X1 U7278 ( .A1(\mem[383][5] ), .A2(n12726), .B1(n26747), .B2(
        data_in[5]), .ZN(n12731) );
  INV_X1 U7279 ( .A(n12732), .ZN(n23036) );
  AOI22_X1 U7280 ( .A1(\mem[383][6] ), .A2(n12726), .B1(n26747), .B2(
        data_in[6]), .ZN(n12732) );
  INV_X1 U7281 ( .A(n12733), .ZN(n23035) );
  AOI22_X1 U7282 ( .A1(\mem[383][7] ), .A2(n12726), .B1(n26747), .B2(
        data_in[7]), .ZN(n12733) );
  INV_X1 U7283 ( .A(n12807), .ZN(n22970) );
  AOI22_X1 U7284 ( .A1(\mem[392][0] ), .A2(n12808), .B1(n26738), .B2(
        data_in[0]), .ZN(n12807) );
  INV_X1 U7285 ( .A(n12809), .ZN(n22969) );
  AOI22_X1 U7286 ( .A1(\mem[392][1] ), .A2(n12808), .B1(n26738), .B2(
        data_in[1]), .ZN(n12809) );
  INV_X1 U7287 ( .A(n12810), .ZN(n22968) );
  AOI22_X1 U7288 ( .A1(\mem[392][2] ), .A2(n12808), .B1(n26738), .B2(
        data_in[2]), .ZN(n12810) );
  INV_X1 U7289 ( .A(n12811), .ZN(n22967) );
  AOI22_X1 U7290 ( .A1(\mem[392][3] ), .A2(n12808), .B1(n26738), .B2(
        data_in[3]), .ZN(n12811) );
  INV_X1 U7291 ( .A(n12812), .ZN(n22966) );
  AOI22_X1 U7292 ( .A1(\mem[392][4] ), .A2(n12808), .B1(n26738), .B2(
        data_in[4]), .ZN(n12812) );
  INV_X1 U7293 ( .A(n12813), .ZN(n22965) );
  AOI22_X1 U7294 ( .A1(\mem[392][5] ), .A2(n12808), .B1(n26738), .B2(
        data_in[5]), .ZN(n12813) );
  INV_X1 U7295 ( .A(n12814), .ZN(n22964) );
  AOI22_X1 U7296 ( .A1(\mem[392][6] ), .A2(n12808), .B1(n26738), .B2(
        data_in[6]), .ZN(n12814) );
  INV_X1 U7297 ( .A(n12815), .ZN(n22963) );
  AOI22_X1 U7298 ( .A1(\mem[392][7] ), .A2(n12808), .B1(n26738), .B2(
        data_in[7]), .ZN(n12815) );
  INV_X1 U7299 ( .A(n12816), .ZN(n22962) );
  AOI22_X1 U7300 ( .A1(\mem[393][0] ), .A2(n12817), .B1(n26737), .B2(
        data_in[0]), .ZN(n12816) );
  INV_X1 U7301 ( .A(n12818), .ZN(n22961) );
  AOI22_X1 U7302 ( .A1(\mem[393][1] ), .A2(n12817), .B1(n26737), .B2(
        data_in[1]), .ZN(n12818) );
  INV_X1 U7303 ( .A(n12819), .ZN(n22960) );
  AOI22_X1 U7304 ( .A1(\mem[393][2] ), .A2(n12817), .B1(n26737), .B2(
        data_in[2]), .ZN(n12819) );
  INV_X1 U7305 ( .A(n12820), .ZN(n22959) );
  AOI22_X1 U7306 ( .A1(\mem[393][3] ), .A2(n12817), .B1(n26737), .B2(
        data_in[3]), .ZN(n12820) );
  INV_X1 U7307 ( .A(n12821), .ZN(n22958) );
  AOI22_X1 U7308 ( .A1(\mem[393][4] ), .A2(n12817), .B1(n26737), .B2(
        data_in[4]), .ZN(n12821) );
  INV_X1 U7309 ( .A(n12822), .ZN(n22957) );
  AOI22_X1 U7310 ( .A1(\mem[393][5] ), .A2(n12817), .B1(n26737), .B2(
        data_in[5]), .ZN(n12822) );
  INV_X1 U7311 ( .A(n12823), .ZN(n22956) );
  AOI22_X1 U7312 ( .A1(\mem[393][6] ), .A2(n12817), .B1(n26737), .B2(
        data_in[6]), .ZN(n12823) );
  INV_X1 U7313 ( .A(n12824), .ZN(n22955) );
  AOI22_X1 U7314 ( .A1(\mem[393][7] ), .A2(n12817), .B1(n26737), .B2(
        data_in[7]), .ZN(n12824) );
  INV_X1 U7315 ( .A(n12825), .ZN(n22954) );
  AOI22_X1 U7316 ( .A1(\mem[394][0] ), .A2(n12826), .B1(n26736), .B2(
        data_in[0]), .ZN(n12825) );
  INV_X1 U7317 ( .A(n12827), .ZN(n22953) );
  AOI22_X1 U7318 ( .A1(\mem[394][1] ), .A2(n12826), .B1(n26736), .B2(
        data_in[1]), .ZN(n12827) );
  INV_X1 U7319 ( .A(n12828), .ZN(n22952) );
  AOI22_X1 U7320 ( .A1(\mem[394][2] ), .A2(n12826), .B1(n26736), .B2(
        data_in[2]), .ZN(n12828) );
  INV_X1 U7321 ( .A(n12829), .ZN(n22951) );
  AOI22_X1 U7322 ( .A1(\mem[394][3] ), .A2(n12826), .B1(n26736), .B2(
        data_in[3]), .ZN(n12829) );
  INV_X1 U7323 ( .A(n12830), .ZN(n22950) );
  AOI22_X1 U7324 ( .A1(\mem[394][4] ), .A2(n12826), .B1(n26736), .B2(
        data_in[4]), .ZN(n12830) );
  INV_X1 U7325 ( .A(n12831), .ZN(n22949) );
  AOI22_X1 U7326 ( .A1(\mem[394][5] ), .A2(n12826), .B1(n26736), .B2(
        data_in[5]), .ZN(n12831) );
  INV_X1 U7327 ( .A(n12832), .ZN(n22948) );
  AOI22_X1 U7328 ( .A1(\mem[394][6] ), .A2(n12826), .B1(n26736), .B2(
        data_in[6]), .ZN(n12832) );
  INV_X1 U7329 ( .A(n12833), .ZN(n22947) );
  AOI22_X1 U7330 ( .A1(\mem[394][7] ), .A2(n12826), .B1(n26736), .B2(
        data_in[7]), .ZN(n12833) );
  INV_X1 U7331 ( .A(n12834), .ZN(n22946) );
  AOI22_X1 U7332 ( .A1(\mem[395][0] ), .A2(n12835), .B1(n26735), .B2(
        data_in[0]), .ZN(n12834) );
  INV_X1 U7333 ( .A(n12836), .ZN(n22945) );
  AOI22_X1 U7334 ( .A1(\mem[395][1] ), .A2(n12835), .B1(n26735), .B2(
        data_in[1]), .ZN(n12836) );
  INV_X1 U7335 ( .A(n12837), .ZN(n22944) );
  AOI22_X1 U7336 ( .A1(\mem[395][2] ), .A2(n12835), .B1(n26735), .B2(
        data_in[2]), .ZN(n12837) );
  INV_X1 U7337 ( .A(n12838), .ZN(n22943) );
  AOI22_X1 U7338 ( .A1(\mem[395][3] ), .A2(n12835), .B1(n26735), .B2(
        data_in[3]), .ZN(n12838) );
  INV_X1 U7339 ( .A(n12839), .ZN(n22942) );
  AOI22_X1 U7340 ( .A1(\mem[395][4] ), .A2(n12835), .B1(n26735), .B2(
        data_in[4]), .ZN(n12839) );
  INV_X1 U7341 ( .A(n12840), .ZN(n22941) );
  AOI22_X1 U7342 ( .A1(\mem[395][5] ), .A2(n12835), .B1(n26735), .B2(
        data_in[5]), .ZN(n12840) );
  INV_X1 U7343 ( .A(n12841), .ZN(n22940) );
  AOI22_X1 U7344 ( .A1(\mem[395][6] ), .A2(n12835), .B1(n26735), .B2(
        data_in[6]), .ZN(n12841) );
  INV_X1 U7345 ( .A(n12842), .ZN(n22939) );
  AOI22_X1 U7346 ( .A1(\mem[395][7] ), .A2(n12835), .B1(n26735), .B2(
        data_in[7]), .ZN(n12842) );
  INV_X1 U7347 ( .A(n12843), .ZN(n22938) );
  AOI22_X1 U7348 ( .A1(\mem[396][0] ), .A2(n12844), .B1(n26734), .B2(
        data_in[0]), .ZN(n12843) );
  INV_X1 U7349 ( .A(n12845), .ZN(n22937) );
  AOI22_X1 U7350 ( .A1(\mem[396][1] ), .A2(n12844), .B1(n26734), .B2(
        data_in[1]), .ZN(n12845) );
  INV_X1 U7351 ( .A(n12846), .ZN(n22936) );
  AOI22_X1 U7352 ( .A1(\mem[396][2] ), .A2(n12844), .B1(n26734), .B2(
        data_in[2]), .ZN(n12846) );
  INV_X1 U7353 ( .A(n12847), .ZN(n22935) );
  AOI22_X1 U7354 ( .A1(\mem[396][3] ), .A2(n12844), .B1(n26734), .B2(
        data_in[3]), .ZN(n12847) );
  INV_X1 U7355 ( .A(n12848), .ZN(n22934) );
  AOI22_X1 U7356 ( .A1(\mem[396][4] ), .A2(n12844), .B1(n26734), .B2(
        data_in[4]), .ZN(n12848) );
  INV_X1 U7357 ( .A(n12849), .ZN(n22933) );
  AOI22_X1 U7358 ( .A1(\mem[396][5] ), .A2(n12844), .B1(n26734), .B2(
        data_in[5]), .ZN(n12849) );
  INV_X1 U7359 ( .A(n12850), .ZN(n22932) );
  AOI22_X1 U7360 ( .A1(\mem[396][6] ), .A2(n12844), .B1(n26734), .B2(
        data_in[6]), .ZN(n12850) );
  INV_X1 U7361 ( .A(n12851), .ZN(n22931) );
  AOI22_X1 U7362 ( .A1(\mem[396][7] ), .A2(n12844), .B1(n26734), .B2(
        data_in[7]), .ZN(n12851) );
  INV_X1 U7363 ( .A(n12852), .ZN(n22930) );
  AOI22_X1 U7364 ( .A1(\mem[397][0] ), .A2(n12853), .B1(n26733), .B2(
        data_in[0]), .ZN(n12852) );
  INV_X1 U7365 ( .A(n12854), .ZN(n22929) );
  AOI22_X1 U7366 ( .A1(\mem[397][1] ), .A2(n12853), .B1(n26733), .B2(
        data_in[1]), .ZN(n12854) );
  INV_X1 U7367 ( .A(n12855), .ZN(n22928) );
  AOI22_X1 U7368 ( .A1(\mem[397][2] ), .A2(n12853), .B1(n26733), .B2(
        data_in[2]), .ZN(n12855) );
  INV_X1 U7369 ( .A(n12856), .ZN(n22927) );
  AOI22_X1 U7370 ( .A1(\mem[397][3] ), .A2(n12853), .B1(n26733), .B2(
        data_in[3]), .ZN(n12856) );
  INV_X1 U7371 ( .A(n12857), .ZN(n22926) );
  AOI22_X1 U7372 ( .A1(\mem[397][4] ), .A2(n12853), .B1(n26733), .B2(
        data_in[4]), .ZN(n12857) );
  INV_X1 U7373 ( .A(n12858), .ZN(n22925) );
  AOI22_X1 U7374 ( .A1(\mem[397][5] ), .A2(n12853), .B1(n26733), .B2(
        data_in[5]), .ZN(n12858) );
  INV_X1 U7375 ( .A(n12859), .ZN(n22924) );
  AOI22_X1 U7376 ( .A1(\mem[397][6] ), .A2(n12853), .B1(n26733), .B2(
        data_in[6]), .ZN(n12859) );
  INV_X1 U7377 ( .A(n12860), .ZN(n22923) );
  AOI22_X1 U7378 ( .A1(\mem[397][7] ), .A2(n12853), .B1(n26733), .B2(
        data_in[7]), .ZN(n12860) );
  INV_X1 U7379 ( .A(n12861), .ZN(n22922) );
  AOI22_X1 U7380 ( .A1(\mem[398][0] ), .A2(n12862), .B1(n26732), .B2(
        data_in[0]), .ZN(n12861) );
  INV_X1 U7381 ( .A(n12863), .ZN(n22921) );
  AOI22_X1 U7382 ( .A1(\mem[398][1] ), .A2(n12862), .B1(n26732), .B2(
        data_in[1]), .ZN(n12863) );
  INV_X1 U7383 ( .A(n12864), .ZN(n22920) );
  AOI22_X1 U7384 ( .A1(\mem[398][2] ), .A2(n12862), .B1(n26732), .B2(
        data_in[2]), .ZN(n12864) );
  INV_X1 U7385 ( .A(n12865), .ZN(n22919) );
  AOI22_X1 U7386 ( .A1(\mem[398][3] ), .A2(n12862), .B1(n26732), .B2(
        data_in[3]), .ZN(n12865) );
  INV_X1 U7387 ( .A(n12866), .ZN(n22918) );
  AOI22_X1 U7388 ( .A1(\mem[398][4] ), .A2(n12862), .B1(n26732), .B2(
        data_in[4]), .ZN(n12866) );
  INV_X1 U7389 ( .A(n12867), .ZN(n22917) );
  AOI22_X1 U7390 ( .A1(\mem[398][5] ), .A2(n12862), .B1(n26732), .B2(
        data_in[5]), .ZN(n12867) );
  INV_X1 U7391 ( .A(n12868), .ZN(n22916) );
  AOI22_X1 U7392 ( .A1(\mem[398][6] ), .A2(n12862), .B1(n26732), .B2(
        data_in[6]), .ZN(n12868) );
  INV_X1 U7393 ( .A(n12869), .ZN(n22915) );
  AOI22_X1 U7394 ( .A1(\mem[398][7] ), .A2(n12862), .B1(n26732), .B2(
        data_in[7]), .ZN(n12869) );
  INV_X1 U7395 ( .A(n12870), .ZN(n22914) );
  AOI22_X1 U7396 ( .A1(\mem[399][0] ), .A2(n12871), .B1(n26731), .B2(
        data_in[0]), .ZN(n12870) );
  INV_X1 U7397 ( .A(n12872), .ZN(n22913) );
  AOI22_X1 U7398 ( .A1(\mem[399][1] ), .A2(n12871), .B1(n26731), .B2(
        data_in[1]), .ZN(n12872) );
  INV_X1 U7399 ( .A(n12873), .ZN(n22912) );
  AOI22_X1 U7400 ( .A1(\mem[399][2] ), .A2(n12871), .B1(n26731), .B2(
        data_in[2]), .ZN(n12873) );
  INV_X1 U7401 ( .A(n12874), .ZN(n22911) );
  AOI22_X1 U7402 ( .A1(\mem[399][3] ), .A2(n12871), .B1(n26731), .B2(
        data_in[3]), .ZN(n12874) );
  INV_X1 U7403 ( .A(n12875), .ZN(n22910) );
  AOI22_X1 U7404 ( .A1(\mem[399][4] ), .A2(n12871), .B1(n26731), .B2(
        data_in[4]), .ZN(n12875) );
  INV_X1 U7405 ( .A(n12876), .ZN(n22909) );
  AOI22_X1 U7406 ( .A1(\mem[399][5] ), .A2(n12871), .B1(n26731), .B2(
        data_in[5]), .ZN(n12876) );
  INV_X1 U7407 ( .A(n12877), .ZN(n22908) );
  AOI22_X1 U7408 ( .A1(\mem[399][6] ), .A2(n12871), .B1(n26731), .B2(
        data_in[6]), .ZN(n12877) );
  INV_X1 U7409 ( .A(n12878), .ZN(n22907) );
  AOI22_X1 U7410 ( .A1(\mem[399][7] ), .A2(n12871), .B1(n26731), .B2(
        data_in[7]), .ZN(n12878) );
  INV_X1 U7411 ( .A(n12879), .ZN(n22906) );
  AOI22_X1 U7412 ( .A1(\mem[400][0] ), .A2(n12880), .B1(n26730), .B2(
        data_in[0]), .ZN(n12879) );
  INV_X1 U7413 ( .A(n12881), .ZN(n22905) );
  AOI22_X1 U7414 ( .A1(\mem[400][1] ), .A2(n12880), .B1(n26730), .B2(
        data_in[1]), .ZN(n12881) );
  INV_X1 U7415 ( .A(n12882), .ZN(n22904) );
  AOI22_X1 U7416 ( .A1(\mem[400][2] ), .A2(n12880), .B1(n26730), .B2(
        data_in[2]), .ZN(n12882) );
  INV_X1 U7417 ( .A(n12883), .ZN(n22903) );
  AOI22_X1 U7418 ( .A1(\mem[400][3] ), .A2(n12880), .B1(n26730), .B2(
        data_in[3]), .ZN(n12883) );
  INV_X1 U7419 ( .A(n12884), .ZN(n22902) );
  AOI22_X1 U7420 ( .A1(\mem[400][4] ), .A2(n12880), .B1(n26730), .B2(
        data_in[4]), .ZN(n12884) );
  INV_X1 U7421 ( .A(n12885), .ZN(n22901) );
  AOI22_X1 U7422 ( .A1(\mem[400][5] ), .A2(n12880), .B1(n26730), .B2(
        data_in[5]), .ZN(n12885) );
  INV_X1 U7423 ( .A(n12886), .ZN(n22900) );
  AOI22_X1 U7424 ( .A1(\mem[400][6] ), .A2(n12880), .B1(n26730), .B2(
        data_in[6]), .ZN(n12886) );
  INV_X1 U7425 ( .A(n12887), .ZN(n22899) );
  AOI22_X1 U7426 ( .A1(\mem[400][7] ), .A2(n12880), .B1(n26730), .B2(
        data_in[7]), .ZN(n12887) );
  INV_X1 U7427 ( .A(n12888), .ZN(n22898) );
  AOI22_X1 U7428 ( .A1(\mem[401][0] ), .A2(n12889), .B1(n26729), .B2(
        data_in[0]), .ZN(n12888) );
  INV_X1 U7429 ( .A(n12890), .ZN(n22897) );
  AOI22_X1 U7430 ( .A1(\mem[401][1] ), .A2(n12889), .B1(n26729), .B2(
        data_in[1]), .ZN(n12890) );
  INV_X1 U7431 ( .A(n12891), .ZN(n22896) );
  AOI22_X1 U7432 ( .A1(\mem[401][2] ), .A2(n12889), .B1(n26729), .B2(
        data_in[2]), .ZN(n12891) );
  INV_X1 U7433 ( .A(n12892), .ZN(n22895) );
  AOI22_X1 U7434 ( .A1(\mem[401][3] ), .A2(n12889), .B1(n26729), .B2(
        data_in[3]), .ZN(n12892) );
  INV_X1 U7435 ( .A(n12893), .ZN(n22894) );
  AOI22_X1 U7436 ( .A1(\mem[401][4] ), .A2(n12889), .B1(n26729), .B2(
        data_in[4]), .ZN(n12893) );
  INV_X1 U7437 ( .A(n12894), .ZN(n22893) );
  AOI22_X1 U7438 ( .A1(\mem[401][5] ), .A2(n12889), .B1(n26729), .B2(
        data_in[5]), .ZN(n12894) );
  INV_X1 U7439 ( .A(n12895), .ZN(n22892) );
  AOI22_X1 U7440 ( .A1(\mem[401][6] ), .A2(n12889), .B1(n26729), .B2(
        data_in[6]), .ZN(n12895) );
  INV_X1 U7441 ( .A(n12896), .ZN(n22891) );
  AOI22_X1 U7442 ( .A1(\mem[401][7] ), .A2(n12889), .B1(n26729), .B2(
        data_in[7]), .ZN(n12896) );
  INV_X1 U7443 ( .A(n12897), .ZN(n22890) );
  AOI22_X1 U7444 ( .A1(\mem[402][0] ), .A2(n12898), .B1(n26728), .B2(
        data_in[0]), .ZN(n12897) );
  INV_X1 U7445 ( .A(n12899), .ZN(n22889) );
  AOI22_X1 U7446 ( .A1(\mem[402][1] ), .A2(n12898), .B1(n26728), .B2(
        data_in[1]), .ZN(n12899) );
  INV_X1 U7447 ( .A(n12900), .ZN(n22888) );
  AOI22_X1 U7448 ( .A1(\mem[402][2] ), .A2(n12898), .B1(n26728), .B2(
        data_in[2]), .ZN(n12900) );
  INV_X1 U7449 ( .A(n12901), .ZN(n22887) );
  AOI22_X1 U7450 ( .A1(\mem[402][3] ), .A2(n12898), .B1(n26728), .B2(
        data_in[3]), .ZN(n12901) );
  INV_X1 U7451 ( .A(n12902), .ZN(n22886) );
  AOI22_X1 U7452 ( .A1(\mem[402][4] ), .A2(n12898), .B1(n26728), .B2(
        data_in[4]), .ZN(n12902) );
  INV_X1 U7453 ( .A(n12903), .ZN(n22885) );
  AOI22_X1 U7454 ( .A1(\mem[402][5] ), .A2(n12898), .B1(n26728), .B2(
        data_in[5]), .ZN(n12903) );
  INV_X1 U7455 ( .A(n12904), .ZN(n22884) );
  AOI22_X1 U7456 ( .A1(\mem[402][6] ), .A2(n12898), .B1(n26728), .B2(
        data_in[6]), .ZN(n12904) );
  INV_X1 U7457 ( .A(n12905), .ZN(n22883) );
  AOI22_X1 U7458 ( .A1(\mem[402][7] ), .A2(n12898), .B1(n26728), .B2(
        data_in[7]), .ZN(n12905) );
  INV_X1 U7459 ( .A(n12906), .ZN(n22882) );
  AOI22_X1 U7460 ( .A1(\mem[403][0] ), .A2(n12907), .B1(n26727), .B2(
        data_in[0]), .ZN(n12906) );
  INV_X1 U7461 ( .A(n12908), .ZN(n22881) );
  AOI22_X1 U7462 ( .A1(\mem[403][1] ), .A2(n12907), .B1(n26727), .B2(
        data_in[1]), .ZN(n12908) );
  INV_X1 U7463 ( .A(n12909), .ZN(n22880) );
  AOI22_X1 U7464 ( .A1(\mem[403][2] ), .A2(n12907), .B1(n26727), .B2(
        data_in[2]), .ZN(n12909) );
  INV_X1 U7465 ( .A(n12910), .ZN(n22879) );
  AOI22_X1 U7466 ( .A1(\mem[403][3] ), .A2(n12907), .B1(n26727), .B2(
        data_in[3]), .ZN(n12910) );
  INV_X1 U7467 ( .A(n12911), .ZN(n22878) );
  AOI22_X1 U7468 ( .A1(\mem[403][4] ), .A2(n12907), .B1(n26727), .B2(
        data_in[4]), .ZN(n12911) );
  INV_X1 U7469 ( .A(n12912), .ZN(n22877) );
  AOI22_X1 U7470 ( .A1(\mem[403][5] ), .A2(n12907), .B1(n26727), .B2(
        data_in[5]), .ZN(n12912) );
  INV_X1 U7471 ( .A(n12913), .ZN(n22876) );
  AOI22_X1 U7472 ( .A1(\mem[403][6] ), .A2(n12907), .B1(n26727), .B2(
        data_in[6]), .ZN(n12913) );
  INV_X1 U7473 ( .A(n12914), .ZN(n22875) );
  AOI22_X1 U7474 ( .A1(\mem[403][7] ), .A2(n12907), .B1(n26727), .B2(
        data_in[7]), .ZN(n12914) );
  INV_X1 U7475 ( .A(n12915), .ZN(n22874) );
  AOI22_X1 U7476 ( .A1(\mem[404][0] ), .A2(n12916), .B1(n26726), .B2(
        data_in[0]), .ZN(n12915) );
  INV_X1 U7477 ( .A(n12917), .ZN(n22873) );
  AOI22_X1 U7478 ( .A1(\mem[404][1] ), .A2(n12916), .B1(n26726), .B2(
        data_in[1]), .ZN(n12917) );
  INV_X1 U7479 ( .A(n12918), .ZN(n22872) );
  AOI22_X1 U7480 ( .A1(\mem[404][2] ), .A2(n12916), .B1(n26726), .B2(
        data_in[2]), .ZN(n12918) );
  INV_X1 U7481 ( .A(n12919), .ZN(n22871) );
  AOI22_X1 U7482 ( .A1(\mem[404][3] ), .A2(n12916), .B1(n26726), .B2(
        data_in[3]), .ZN(n12919) );
  INV_X1 U7483 ( .A(n12920), .ZN(n22870) );
  AOI22_X1 U7484 ( .A1(\mem[404][4] ), .A2(n12916), .B1(n26726), .B2(
        data_in[4]), .ZN(n12920) );
  INV_X1 U7485 ( .A(n12921), .ZN(n22869) );
  AOI22_X1 U7486 ( .A1(\mem[404][5] ), .A2(n12916), .B1(n26726), .B2(
        data_in[5]), .ZN(n12921) );
  INV_X1 U7487 ( .A(n12922), .ZN(n22868) );
  AOI22_X1 U7488 ( .A1(\mem[404][6] ), .A2(n12916), .B1(n26726), .B2(
        data_in[6]), .ZN(n12922) );
  INV_X1 U7489 ( .A(n12923), .ZN(n22867) );
  AOI22_X1 U7490 ( .A1(\mem[404][7] ), .A2(n12916), .B1(n26726), .B2(
        data_in[7]), .ZN(n12923) );
  INV_X1 U7491 ( .A(n12924), .ZN(n22866) );
  AOI22_X1 U7492 ( .A1(\mem[405][0] ), .A2(n12925), .B1(n26725), .B2(
        data_in[0]), .ZN(n12924) );
  INV_X1 U7493 ( .A(n12926), .ZN(n22865) );
  AOI22_X1 U7494 ( .A1(\mem[405][1] ), .A2(n12925), .B1(n26725), .B2(
        data_in[1]), .ZN(n12926) );
  INV_X1 U7495 ( .A(n12927), .ZN(n22864) );
  AOI22_X1 U7496 ( .A1(\mem[405][2] ), .A2(n12925), .B1(n26725), .B2(
        data_in[2]), .ZN(n12927) );
  INV_X1 U7497 ( .A(n12928), .ZN(n22863) );
  AOI22_X1 U7498 ( .A1(\mem[405][3] ), .A2(n12925), .B1(n26725), .B2(
        data_in[3]), .ZN(n12928) );
  INV_X1 U7499 ( .A(n12929), .ZN(n22862) );
  AOI22_X1 U7500 ( .A1(\mem[405][4] ), .A2(n12925), .B1(n26725), .B2(
        data_in[4]), .ZN(n12929) );
  INV_X1 U7501 ( .A(n12930), .ZN(n22861) );
  AOI22_X1 U7502 ( .A1(\mem[405][5] ), .A2(n12925), .B1(n26725), .B2(
        data_in[5]), .ZN(n12930) );
  INV_X1 U7503 ( .A(n12931), .ZN(n22860) );
  AOI22_X1 U7504 ( .A1(\mem[405][6] ), .A2(n12925), .B1(n26725), .B2(
        data_in[6]), .ZN(n12931) );
  INV_X1 U7505 ( .A(n12932), .ZN(n22859) );
  AOI22_X1 U7506 ( .A1(\mem[405][7] ), .A2(n12925), .B1(n26725), .B2(
        data_in[7]), .ZN(n12932) );
  INV_X1 U7507 ( .A(n12933), .ZN(n22858) );
  AOI22_X1 U7508 ( .A1(\mem[406][0] ), .A2(n12934), .B1(n26724), .B2(
        data_in[0]), .ZN(n12933) );
  INV_X1 U7509 ( .A(n12935), .ZN(n22857) );
  AOI22_X1 U7510 ( .A1(\mem[406][1] ), .A2(n12934), .B1(n26724), .B2(
        data_in[1]), .ZN(n12935) );
  INV_X1 U7511 ( .A(n12936), .ZN(n22856) );
  AOI22_X1 U7512 ( .A1(\mem[406][2] ), .A2(n12934), .B1(n26724), .B2(
        data_in[2]), .ZN(n12936) );
  INV_X1 U7513 ( .A(n12937), .ZN(n22855) );
  AOI22_X1 U7514 ( .A1(\mem[406][3] ), .A2(n12934), .B1(n26724), .B2(
        data_in[3]), .ZN(n12937) );
  INV_X1 U7515 ( .A(n12938), .ZN(n22854) );
  AOI22_X1 U7516 ( .A1(\mem[406][4] ), .A2(n12934), .B1(n26724), .B2(
        data_in[4]), .ZN(n12938) );
  INV_X1 U7517 ( .A(n12939), .ZN(n22853) );
  AOI22_X1 U7518 ( .A1(\mem[406][5] ), .A2(n12934), .B1(n26724), .B2(
        data_in[5]), .ZN(n12939) );
  INV_X1 U7519 ( .A(n12940), .ZN(n22852) );
  AOI22_X1 U7520 ( .A1(\mem[406][6] ), .A2(n12934), .B1(n26724), .B2(
        data_in[6]), .ZN(n12940) );
  INV_X1 U7521 ( .A(n12941), .ZN(n22851) );
  AOI22_X1 U7522 ( .A1(\mem[406][7] ), .A2(n12934), .B1(n26724), .B2(
        data_in[7]), .ZN(n12941) );
  INV_X1 U7523 ( .A(n12942), .ZN(n22850) );
  AOI22_X1 U7524 ( .A1(\mem[407][0] ), .A2(n12943), .B1(n26723), .B2(
        data_in[0]), .ZN(n12942) );
  INV_X1 U7525 ( .A(n12944), .ZN(n22849) );
  AOI22_X1 U7526 ( .A1(\mem[407][1] ), .A2(n12943), .B1(n26723), .B2(
        data_in[1]), .ZN(n12944) );
  INV_X1 U7527 ( .A(n12945), .ZN(n22848) );
  AOI22_X1 U7528 ( .A1(\mem[407][2] ), .A2(n12943), .B1(n26723), .B2(
        data_in[2]), .ZN(n12945) );
  INV_X1 U7529 ( .A(n12946), .ZN(n22847) );
  AOI22_X1 U7530 ( .A1(\mem[407][3] ), .A2(n12943), .B1(n26723), .B2(
        data_in[3]), .ZN(n12946) );
  INV_X1 U7531 ( .A(n12947), .ZN(n22846) );
  AOI22_X1 U7532 ( .A1(\mem[407][4] ), .A2(n12943), .B1(n26723), .B2(
        data_in[4]), .ZN(n12947) );
  INV_X1 U7533 ( .A(n12948), .ZN(n22845) );
  AOI22_X1 U7534 ( .A1(\mem[407][5] ), .A2(n12943), .B1(n26723), .B2(
        data_in[5]), .ZN(n12948) );
  INV_X1 U7535 ( .A(n12949), .ZN(n22844) );
  AOI22_X1 U7536 ( .A1(\mem[407][6] ), .A2(n12943), .B1(n26723), .B2(
        data_in[6]), .ZN(n12949) );
  INV_X1 U7537 ( .A(n12950), .ZN(n22843) );
  AOI22_X1 U7538 ( .A1(\mem[407][7] ), .A2(n12943), .B1(n26723), .B2(
        data_in[7]), .ZN(n12950) );
  INV_X1 U7539 ( .A(n12951), .ZN(n22842) );
  AOI22_X1 U7540 ( .A1(\mem[408][0] ), .A2(n12952), .B1(n26722), .B2(
        data_in[0]), .ZN(n12951) );
  INV_X1 U7541 ( .A(n12953), .ZN(n22841) );
  AOI22_X1 U7542 ( .A1(\mem[408][1] ), .A2(n12952), .B1(n26722), .B2(
        data_in[1]), .ZN(n12953) );
  INV_X1 U7543 ( .A(n12954), .ZN(n22840) );
  AOI22_X1 U7544 ( .A1(\mem[408][2] ), .A2(n12952), .B1(n26722), .B2(
        data_in[2]), .ZN(n12954) );
  INV_X1 U7545 ( .A(n12955), .ZN(n22839) );
  AOI22_X1 U7546 ( .A1(\mem[408][3] ), .A2(n12952), .B1(n26722), .B2(
        data_in[3]), .ZN(n12955) );
  INV_X1 U7547 ( .A(n12956), .ZN(n22838) );
  AOI22_X1 U7548 ( .A1(\mem[408][4] ), .A2(n12952), .B1(n26722), .B2(
        data_in[4]), .ZN(n12956) );
  INV_X1 U7549 ( .A(n12957), .ZN(n22837) );
  AOI22_X1 U7550 ( .A1(\mem[408][5] ), .A2(n12952), .B1(n26722), .B2(
        data_in[5]), .ZN(n12957) );
  INV_X1 U7551 ( .A(n12958), .ZN(n22836) );
  AOI22_X1 U7552 ( .A1(\mem[408][6] ), .A2(n12952), .B1(n26722), .B2(
        data_in[6]), .ZN(n12958) );
  INV_X1 U7553 ( .A(n12959), .ZN(n22835) );
  AOI22_X1 U7554 ( .A1(\mem[408][7] ), .A2(n12952), .B1(n26722), .B2(
        data_in[7]), .ZN(n12959) );
  INV_X1 U7555 ( .A(n12960), .ZN(n22834) );
  AOI22_X1 U7556 ( .A1(\mem[409][0] ), .A2(n12961), .B1(n26721), .B2(
        data_in[0]), .ZN(n12960) );
  INV_X1 U7557 ( .A(n12962), .ZN(n22833) );
  AOI22_X1 U7558 ( .A1(\mem[409][1] ), .A2(n12961), .B1(n26721), .B2(
        data_in[1]), .ZN(n12962) );
  INV_X1 U7559 ( .A(n12963), .ZN(n22832) );
  AOI22_X1 U7560 ( .A1(\mem[409][2] ), .A2(n12961), .B1(n26721), .B2(
        data_in[2]), .ZN(n12963) );
  INV_X1 U7561 ( .A(n12964), .ZN(n22831) );
  AOI22_X1 U7562 ( .A1(\mem[409][3] ), .A2(n12961), .B1(n26721), .B2(
        data_in[3]), .ZN(n12964) );
  INV_X1 U7563 ( .A(n12965), .ZN(n22830) );
  AOI22_X1 U7564 ( .A1(\mem[409][4] ), .A2(n12961), .B1(n26721), .B2(
        data_in[4]), .ZN(n12965) );
  INV_X1 U7565 ( .A(n12966), .ZN(n22829) );
  AOI22_X1 U7566 ( .A1(\mem[409][5] ), .A2(n12961), .B1(n26721), .B2(
        data_in[5]), .ZN(n12966) );
  INV_X1 U7567 ( .A(n12967), .ZN(n22828) );
  AOI22_X1 U7568 ( .A1(\mem[409][6] ), .A2(n12961), .B1(n26721), .B2(
        data_in[6]), .ZN(n12967) );
  INV_X1 U7569 ( .A(n12968), .ZN(n22827) );
  AOI22_X1 U7570 ( .A1(\mem[409][7] ), .A2(n12961), .B1(n26721), .B2(
        data_in[7]), .ZN(n12968) );
  INV_X1 U7571 ( .A(n12969), .ZN(n22826) );
  AOI22_X1 U7572 ( .A1(\mem[410][0] ), .A2(n12970), .B1(n26720), .B2(
        data_in[0]), .ZN(n12969) );
  INV_X1 U7573 ( .A(n12971), .ZN(n22825) );
  AOI22_X1 U7574 ( .A1(\mem[410][1] ), .A2(n12970), .B1(n26720), .B2(
        data_in[1]), .ZN(n12971) );
  INV_X1 U7575 ( .A(n12972), .ZN(n22824) );
  AOI22_X1 U7576 ( .A1(\mem[410][2] ), .A2(n12970), .B1(n26720), .B2(
        data_in[2]), .ZN(n12972) );
  INV_X1 U7577 ( .A(n12973), .ZN(n22823) );
  AOI22_X1 U7578 ( .A1(\mem[410][3] ), .A2(n12970), .B1(n26720), .B2(
        data_in[3]), .ZN(n12973) );
  INV_X1 U7579 ( .A(n12974), .ZN(n22822) );
  AOI22_X1 U7580 ( .A1(\mem[410][4] ), .A2(n12970), .B1(n26720), .B2(
        data_in[4]), .ZN(n12974) );
  INV_X1 U7581 ( .A(n12975), .ZN(n22821) );
  AOI22_X1 U7582 ( .A1(\mem[410][5] ), .A2(n12970), .B1(n26720), .B2(
        data_in[5]), .ZN(n12975) );
  INV_X1 U7583 ( .A(n12976), .ZN(n22820) );
  AOI22_X1 U7584 ( .A1(\mem[410][6] ), .A2(n12970), .B1(n26720), .B2(
        data_in[6]), .ZN(n12976) );
  INV_X1 U7585 ( .A(n12977), .ZN(n22819) );
  AOI22_X1 U7586 ( .A1(\mem[410][7] ), .A2(n12970), .B1(n26720), .B2(
        data_in[7]), .ZN(n12977) );
  INV_X1 U7587 ( .A(n12978), .ZN(n22818) );
  AOI22_X1 U7588 ( .A1(\mem[411][0] ), .A2(n12979), .B1(n26719), .B2(
        data_in[0]), .ZN(n12978) );
  INV_X1 U7589 ( .A(n12980), .ZN(n22817) );
  AOI22_X1 U7590 ( .A1(\mem[411][1] ), .A2(n12979), .B1(n26719), .B2(
        data_in[1]), .ZN(n12980) );
  INV_X1 U7591 ( .A(n12981), .ZN(n22816) );
  AOI22_X1 U7592 ( .A1(\mem[411][2] ), .A2(n12979), .B1(n26719), .B2(
        data_in[2]), .ZN(n12981) );
  INV_X1 U7593 ( .A(n12982), .ZN(n22815) );
  AOI22_X1 U7594 ( .A1(\mem[411][3] ), .A2(n12979), .B1(n26719), .B2(
        data_in[3]), .ZN(n12982) );
  INV_X1 U7595 ( .A(n12983), .ZN(n22814) );
  AOI22_X1 U7596 ( .A1(\mem[411][4] ), .A2(n12979), .B1(n26719), .B2(
        data_in[4]), .ZN(n12983) );
  INV_X1 U7597 ( .A(n12984), .ZN(n22813) );
  AOI22_X1 U7598 ( .A1(\mem[411][5] ), .A2(n12979), .B1(n26719), .B2(
        data_in[5]), .ZN(n12984) );
  INV_X1 U7599 ( .A(n12985), .ZN(n22812) );
  AOI22_X1 U7600 ( .A1(\mem[411][6] ), .A2(n12979), .B1(n26719), .B2(
        data_in[6]), .ZN(n12985) );
  INV_X1 U7601 ( .A(n12986), .ZN(n22811) );
  AOI22_X1 U7602 ( .A1(\mem[411][7] ), .A2(n12979), .B1(n26719), .B2(
        data_in[7]), .ZN(n12986) );
  INV_X1 U7603 ( .A(n12987), .ZN(n22810) );
  AOI22_X1 U7604 ( .A1(\mem[412][0] ), .A2(n12988), .B1(n26718), .B2(
        data_in[0]), .ZN(n12987) );
  INV_X1 U7605 ( .A(n12989), .ZN(n22809) );
  AOI22_X1 U7606 ( .A1(\mem[412][1] ), .A2(n12988), .B1(n26718), .B2(
        data_in[1]), .ZN(n12989) );
  INV_X1 U7607 ( .A(n12990), .ZN(n22808) );
  AOI22_X1 U7608 ( .A1(\mem[412][2] ), .A2(n12988), .B1(n26718), .B2(
        data_in[2]), .ZN(n12990) );
  INV_X1 U7609 ( .A(n12991), .ZN(n22807) );
  AOI22_X1 U7610 ( .A1(\mem[412][3] ), .A2(n12988), .B1(n26718), .B2(
        data_in[3]), .ZN(n12991) );
  INV_X1 U7611 ( .A(n12992), .ZN(n22806) );
  AOI22_X1 U7612 ( .A1(\mem[412][4] ), .A2(n12988), .B1(n26718), .B2(
        data_in[4]), .ZN(n12992) );
  INV_X1 U7613 ( .A(n12993), .ZN(n22805) );
  AOI22_X1 U7614 ( .A1(\mem[412][5] ), .A2(n12988), .B1(n26718), .B2(
        data_in[5]), .ZN(n12993) );
  INV_X1 U7615 ( .A(n12994), .ZN(n22804) );
  AOI22_X1 U7616 ( .A1(\mem[412][6] ), .A2(n12988), .B1(n26718), .B2(
        data_in[6]), .ZN(n12994) );
  INV_X1 U7617 ( .A(n12995), .ZN(n22803) );
  AOI22_X1 U7618 ( .A1(\mem[412][7] ), .A2(n12988), .B1(n26718), .B2(
        data_in[7]), .ZN(n12995) );
  INV_X1 U7619 ( .A(n12996), .ZN(n22802) );
  AOI22_X1 U7620 ( .A1(\mem[413][0] ), .A2(n12997), .B1(n26717), .B2(
        data_in[0]), .ZN(n12996) );
  INV_X1 U7621 ( .A(n12998), .ZN(n22801) );
  AOI22_X1 U7622 ( .A1(\mem[413][1] ), .A2(n12997), .B1(n26717), .B2(
        data_in[1]), .ZN(n12998) );
  INV_X1 U7623 ( .A(n12999), .ZN(n22800) );
  AOI22_X1 U7624 ( .A1(\mem[413][2] ), .A2(n12997), .B1(n26717), .B2(
        data_in[2]), .ZN(n12999) );
  INV_X1 U7625 ( .A(n13000), .ZN(n22799) );
  AOI22_X1 U7626 ( .A1(\mem[413][3] ), .A2(n12997), .B1(n26717), .B2(
        data_in[3]), .ZN(n13000) );
  INV_X1 U7627 ( .A(n13001), .ZN(n22798) );
  AOI22_X1 U7628 ( .A1(\mem[413][4] ), .A2(n12997), .B1(n26717), .B2(
        data_in[4]), .ZN(n13001) );
  INV_X1 U7629 ( .A(n13002), .ZN(n22797) );
  AOI22_X1 U7630 ( .A1(\mem[413][5] ), .A2(n12997), .B1(n26717), .B2(
        data_in[5]), .ZN(n13002) );
  INV_X1 U7631 ( .A(n13003), .ZN(n22796) );
  AOI22_X1 U7632 ( .A1(\mem[413][6] ), .A2(n12997), .B1(n26717), .B2(
        data_in[6]), .ZN(n13003) );
  INV_X1 U7633 ( .A(n13004), .ZN(n22795) );
  AOI22_X1 U7634 ( .A1(\mem[413][7] ), .A2(n12997), .B1(n26717), .B2(
        data_in[7]), .ZN(n13004) );
  INV_X1 U7635 ( .A(n13005), .ZN(n22794) );
  AOI22_X1 U7636 ( .A1(\mem[414][0] ), .A2(n13006), .B1(n26716), .B2(
        data_in[0]), .ZN(n13005) );
  INV_X1 U7637 ( .A(n13007), .ZN(n22793) );
  AOI22_X1 U7638 ( .A1(\mem[414][1] ), .A2(n13006), .B1(n26716), .B2(
        data_in[1]), .ZN(n13007) );
  INV_X1 U7639 ( .A(n13008), .ZN(n22792) );
  AOI22_X1 U7640 ( .A1(\mem[414][2] ), .A2(n13006), .B1(n26716), .B2(
        data_in[2]), .ZN(n13008) );
  INV_X1 U7641 ( .A(n13009), .ZN(n22791) );
  AOI22_X1 U7642 ( .A1(\mem[414][3] ), .A2(n13006), .B1(n26716), .B2(
        data_in[3]), .ZN(n13009) );
  INV_X1 U7643 ( .A(n13010), .ZN(n22790) );
  AOI22_X1 U7644 ( .A1(\mem[414][4] ), .A2(n13006), .B1(n26716), .B2(
        data_in[4]), .ZN(n13010) );
  INV_X1 U7645 ( .A(n13011), .ZN(n22789) );
  AOI22_X1 U7646 ( .A1(\mem[414][5] ), .A2(n13006), .B1(n26716), .B2(
        data_in[5]), .ZN(n13011) );
  INV_X1 U7647 ( .A(n13012), .ZN(n22788) );
  AOI22_X1 U7648 ( .A1(\mem[414][6] ), .A2(n13006), .B1(n26716), .B2(
        data_in[6]), .ZN(n13012) );
  INV_X1 U7649 ( .A(n13013), .ZN(n22787) );
  AOI22_X1 U7650 ( .A1(\mem[414][7] ), .A2(n13006), .B1(n26716), .B2(
        data_in[7]), .ZN(n13013) );
  INV_X1 U7651 ( .A(n13014), .ZN(n22786) );
  AOI22_X1 U7652 ( .A1(\mem[415][0] ), .A2(n13015), .B1(n26715), .B2(
        data_in[0]), .ZN(n13014) );
  INV_X1 U7653 ( .A(n13016), .ZN(n22785) );
  AOI22_X1 U7654 ( .A1(\mem[415][1] ), .A2(n13015), .B1(n26715), .B2(
        data_in[1]), .ZN(n13016) );
  INV_X1 U7655 ( .A(n13017), .ZN(n22784) );
  AOI22_X1 U7656 ( .A1(\mem[415][2] ), .A2(n13015), .B1(n26715), .B2(
        data_in[2]), .ZN(n13017) );
  INV_X1 U7657 ( .A(n13018), .ZN(n22783) );
  AOI22_X1 U7658 ( .A1(\mem[415][3] ), .A2(n13015), .B1(n26715), .B2(
        data_in[3]), .ZN(n13018) );
  INV_X1 U7659 ( .A(n13019), .ZN(n22782) );
  AOI22_X1 U7660 ( .A1(\mem[415][4] ), .A2(n13015), .B1(n26715), .B2(
        data_in[4]), .ZN(n13019) );
  INV_X1 U7661 ( .A(n13020), .ZN(n22781) );
  AOI22_X1 U7662 ( .A1(\mem[415][5] ), .A2(n13015), .B1(n26715), .B2(
        data_in[5]), .ZN(n13020) );
  INV_X1 U7663 ( .A(n13021), .ZN(n22780) );
  AOI22_X1 U7664 ( .A1(\mem[415][6] ), .A2(n13015), .B1(n26715), .B2(
        data_in[6]), .ZN(n13021) );
  INV_X1 U7665 ( .A(n13022), .ZN(n22779) );
  AOI22_X1 U7666 ( .A1(\mem[415][7] ), .A2(n13015), .B1(n26715), .B2(
        data_in[7]), .ZN(n13022) );
  INV_X1 U7667 ( .A(n13096), .ZN(n22714) );
  AOI22_X1 U7668 ( .A1(\mem[424][0] ), .A2(n13097), .B1(n26706), .B2(
        data_in[0]), .ZN(n13096) );
  INV_X1 U7669 ( .A(n13098), .ZN(n22713) );
  AOI22_X1 U7670 ( .A1(\mem[424][1] ), .A2(n13097), .B1(n26706), .B2(
        data_in[1]), .ZN(n13098) );
  INV_X1 U7671 ( .A(n13099), .ZN(n22712) );
  AOI22_X1 U7672 ( .A1(\mem[424][2] ), .A2(n13097), .B1(n26706), .B2(
        data_in[2]), .ZN(n13099) );
  INV_X1 U7673 ( .A(n13100), .ZN(n22711) );
  AOI22_X1 U7674 ( .A1(\mem[424][3] ), .A2(n13097), .B1(n26706), .B2(
        data_in[3]), .ZN(n13100) );
  INV_X1 U7675 ( .A(n13101), .ZN(n22710) );
  AOI22_X1 U7676 ( .A1(\mem[424][4] ), .A2(n13097), .B1(n26706), .B2(
        data_in[4]), .ZN(n13101) );
  INV_X1 U7677 ( .A(n13102), .ZN(n22709) );
  AOI22_X1 U7678 ( .A1(\mem[424][5] ), .A2(n13097), .B1(n26706), .B2(
        data_in[5]), .ZN(n13102) );
  INV_X1 U7679 ( .A(n13103), .ZN(n22708) );
  AOI22_X1 U7680 ( .A1(\mem[424][6] ), .A2(n13097), .B1(n26706), .B2(
        data_in[6]), .ZN(n13103) );
  INV_X1 U7681 ( .A(n13104), .ZN(n22707) );
  AOI22_X1 U7682 ( .A1(\mem[424][7] ), .A2(n13097), .B1(n26706), .B2(
        data_in[7]), .ZN(n13104) );
  INV_X1 U7683 ( .A(n13105), .ZN(n22706) );
  AOI22_X1 U7684 ( .A1(\mem[425][0] ), .A2(n13106), .B1(n26705), .B2(
        data_in[0]), .ZN(n13105) );
  INV_X1 U7685 ( .A(n13107), .ZN(n22705) );
  AOI22_X1 U7686 ( .A1(\mem[425][1] ), .A2(n13106), .B1(n26705), .B2(
        data_in[1]), .ZN(n13107) );
  INV_X1 U7687 ( .A(n13108), .ZN(n22704) );
  AOI22_X1 U7688 ( .A1(\mem[425][2] ), .A2(n13106), .B1(n26705), .B2(
        data_in[2]), .ZN(n13108) );
  INV_X1 U7689 ( .A(n13109), .ZN(n22703) );
  AOI22_X1 U7690 ( .A1(\mem[425][3] ), .A2(n13106), .B1(n26705), .B2(
        data_in[3]), .ZN(n13109) );
  INV_X1 U7691 ( .A(n13110), .ZN(n22702) );
  AOI22_X1 U7692 ( .A1(\mem[425][4] ), .A2(n13106), .B1(n26705), .B2(
        data_in[4]), .ZN(n13110) );
  INV_X1 U7693 ( .A(n13111), .ZN(n22701) );
  AOI22_X1 U7694 ( .A1(\mem[425][5] ), .A2(n13106), .B1(n26705), .B2(
        data_in[5]), .ZN(n13111) );
  INV_X1 U7695 ( .A(n13112), .ZN(n22700) );
  AOI22_X1 U7696 ( .A1(\mem[425][6] ), .A2(n13106), .B1(n26705), .B2(
        data_in[6]), .ZN(n13112) );
  INV_X1 U7697 ( .A(n13113), .ZN(n22699) );
  AOI22_X1 U7698 ( .A1(\mem[425][7] ), .A2(n13106), .B1(n26705), .B2(
        data_in[7]), .ZN(n13113) );
  INV_X1 U7699 ( .A(n13114), .ZN(n22698) );
  AOI22_X1 U7700 ( .A1(\mem[426][0] ), .A2(n13115), .B1(n26704), .B2(
        data_in[0]), .ZN(n13114) );
  INV_X1 U7701 ( .A(n13116), .ZN(n22697) );
  AOI22_X1 U7702 ( .A1(\mem[426][1] ), .A2(n13115), .B1(n26704), .B2(
        data_in[1]), .ZN(n13116) );
  INV_X1 U7703 ( .A(n13117), .ZN(n22696) );
  AOI22_X1 U7704 ( .A1(\mem[426][2] ), .A2(n13115), .B1(n26704), .B2(
        data_in[2]), .ZN(n13117) );
  INV_X1 U7705 ( .A(n13118), .ZN(n22695) );
  AOI22_X1 U7706 ( .A1(\mem[426][3] ), .A2(n13115), .B1(n26704), .B2(
        data_in[3]), .ZN(n13118) );
  INV_X1 U7707 ( .A(n13119), .ZN(n22694) );
  AOI22_X1 U7708 ( .A1(\mem[426][4] ), .A2(n13115), .B1(n26704), .B2(
        data_in[4]), .ZN(n13119) );
  INV_X1 U7709 ( .A(n13120), .ZN(n22693) );
  AOI22_X1 U7710 ( .A1(\mem[426][5] ), .A2(n13115), .B1(n26704), .B2(
        data_in[5]), .ZN(n13120) );
  INV_X1 U7711 ( .A(n13121), .ZN(n22692) );
  AOI22_X1 U7712 ( .A1(\mem[426][6] ), .A2(n13115), .B1(n26704), .B2(
        data_in[6]), .ZN(n13121) );
  INV_X1 U7713 ( .A(n13122), .ZN(n22691) );
  AOI22_X1 U7714 ( .A1(\mem[426][7] ), .A2(n13115), .B1(n26704), .B2(
        data_in[7]), .ZN(n13122) );
  INV_X1 U7715 ( .A(n13123), .ZN(n22690) );
  AOI22_X1 U7716 ( .A1(\mem[427][0] ), .A2(n13124), .B1(n26703), .B2(
        data_in[0]), .ZN(n13123) );
  INV_X1 U7717 ( .A(n13125), .ZN(n22689) );
  AOI22_X1 U7718 ( .A1(\mem[427][1] ), .A2(n13124), .B1(n26703), .B2(
        data_in[1]), .ZN(n13125) );
  INV_X1 U7719 ( .A(n13126), .ZN(n22688) );
  AOI22_X1 U7720 ( .A1(\mem[427][2] ), .A2(n13124), .B1(n26703), .B2(
        data_in[2]), .ZN(n13126) );
  INV_X1 U7721 ( .A(n13127), .ZN(n22687) );
  AOI22_X1 U7722 ( .A1(\mem[427][3] ), .A2(n13124), .B1(n26703), .B2(
        data_in[3]), .ZN(n13127) );
  INV_X1 U7723 ( .A(n13128), .ZN(n22686) );
  AOI22_X1 U7724 ( .A1(\mem[427][4] ), .A2(n13124), .B1(n26703), .B2(
        data_in[4]), .ZN(n13128) );
  INV_X1 U7725 ( .A(n13129), .ZN(n22685) );
  AOI22_X1 U7726 ( .A1(\mem[427][5] ), .A2(n13124), .B1(n26703), .B2(
        data_in[5]), .ZN(n13129) );
  INV_X1 U7727 ( .A(n13130), .ZN(n22684) );
  AOI22_X1 U7728 ( .A1(\mem[427][6] ), .A2(n13124), .B1(n26703), .B2(
        data_in[6]), .ZN(n13130) );
  INV_X1 U7729 ( .A(n13131), .ZN(n22683) );
  AOI22_X1 U7730 ( .A1(\mem[427][7] ), .A2(n13124), .B1(n26703), .B2(
        data_in[7]), .ZN(n13131) );
  INV_X1 U7731 ( .A(n13132), .ZN(n22682) );
  AOI22_X1 U7732 ( .A1(\mem[428][0] ), .A2(n13133), .B1(n26702), .B2(
        data_in[0]), .ZN(n13132) );
  INV_X1 U7733 ( .A(n13134), .ZN(n22681) );
  AOI22_X1 U7734 ( .A1(\mem[428][1] ), .A2(n13133), .B1(n26702), .B2(
        data_in[1]), .ZN(n13134) );
  INV_X1 U7735 ( .A(n13135), .ZN(n22680) );
  AOI22_X1 U7736 ( .A1(\mem[428][2] ), .A2(n13133), .B1(n26702), .B2(
        data_in[2]), .ZN(n13135) );
  INV_X1 U7737 ( .A(n13136), .ZN(n22679) );
  AOI22_X1 U7738 ( .A1(\mem[428][3] ), .A2(n13133), .B1(n26702), .B2(
        data_in[3]), .ZN(n13136) );
  INV_X1 U7739 ( .A(n13137), .ZN(n22678) );
  AOI22_X1 U7740 ( .A1(\mem[428][4] ), .A2(n13133), .B1(n26702), .B2(
        data_in[4]), .ZN(n13137) );
  INV_X1 U7741 ( .A(n13138), .ZN(n22677) );
  AOI22_X1 U7742 ( .A1(\mem[428][5] ), .A2(n13133), .B1(n26702), .B2(
        data_in[5]), .ZN(n13138) );
  INV_X1 U7743 ( .A(n13139), .ZN(n22676) );
  AOI22_X1 U7744 ( .A1(\mem[428][6] ), .A2(n13133), .B1(n26702), .B2(
        data_in[6]), .ZN(n13139) );
  INV_X1 U7745 ( .A(n13140), .ZN(n22675) );
  AOI22_X1 U7746 ( .A1(\mem[428][7] ), .A2(n13133), .B1(n26702), .B2(
        data_in[7]), .ZN(n13140) );
  INV_X1 U7747 ( .A(n13141), .ZN(n22674) );
  AOI22_X1 U7748 ( .A1(\mem[429][0] ), .A2(n13142), .B1(n26701), .B2(
        data_in[0]), .ZN(n13141) );
  INV_X1 U7749 ( .A(n13143), .ZN(n22673) );
  AOI22_X1 U7750 ( .A1(\mem[429][1] ), .A2(n13142), .B1(n26701), .B2(
        data_in[1]), .ZN(n13143) );
  INV_X1 U7751 ( .A(n13144), .ZN(n22672) );
  AOI22_X1 U7752 ( .A1(\mem[429][2] ), .A2(n13142), .B1(n26701), .B2(
        data_in[2]), .ZN(n13144) );
  INV_X1 U7753 ( .A(n13145), .ZN(n22671) );
  AOI22_X1 U7754 ( .A1(\mem[429][3] ), .A2(n13142), .B1(n26701), .B2(
        data_in[3]), .ZN(n13145) );
  INV_X1 U7755 ( .A(n13146), .ZN(n22670) );
  AOI22_X1 U7756 ( .A1(\mem[429][4] ), .A2(n13142), .B1(n26701), .B2(
        data_in[4]), .ZN(n13146) );
  INV_X1 U7757 ( .A(n13147), .ZN(n22669) );
  AOI22_X1 U7758 ( .A1(\mem[429][5] ), .A2(n13142), .B1(n26701), .B2(
        data_in[5]), .ZN(n13147) );
  INV_X1 U7759 ( .A(n13148), .ZN(n22668) );
  AOI22_X1 U7760 ( .A1(\mem[429][6] ), .A2(n13142), .B1(n26701), .B2(
        data_in[6]), .ZN(n13148) );
  INV_X1 U7761 ( .A(n13149), .ZN(n22667) );
  AOI22_X1 U7762 ( .A1(\mem[429][7] ), .A2(n13142), .B1(n26701), .B2(
        data_in[7]), .ZN(n13149) );
  INV_X1 U7763 ( .A(n13150), .ZN(n22666) );
  AOI22_X1 U7764 ( .A1(\mem[430][0] ), .A2(n13151), .B1(n26700), .B2(
        data_in[0]), .ZN(n13150) );
  INV_X1 U7765 ( .A(n13152), .ZN(n22665) );
  AOI22_X1 U7766 ( .A1(\mem[430][1] ), .A2(n13151), .B1(n26700), .B2(
        data_in[1]), .ZN(n13152) );
  INV_X1 U7767 ( .A(n13153), .ZN(n22664) );
  AOI22_X1 U7768 ( .A1(\mem[430][2] ), .A2(n13151), .B1(n26700), .B2(
        data_in[2]), .ZN(n13153) );
  INV_X1 U7769 ( .A(n13154), .ZN(n22663) );
  AOI22_X1 U7770 ( .A1(\mem[430][3] ), .A2(n13151), .B1(n26700), .B2(
        data_in[3]), .ZN(n13154) );
  INV_X1 U7771 ( .A(n13155), .ZN(n22662) );
  AOI22_X1 U7772 ( .A1(\mem[430][4] ), .A2(n13151), .B1(n26700), .B2(
        data_in[4]), .ZN(n13155) );
  INV_X1 U7773 ( .A(n13156), .ZN(n22661) );
  AOI22_X1 U7774 ( .A1(\mem[430][5] ), .A2(n13151), .B1(n26700), .B2(
        data_in[5]), .ZN(n13156) );
  INV_X1 U7775 ( .A(n13157), .ZN(n22660) );
  AOI22_X1 U7776 ( .A1(\mem[430][6] ), .A2(n13151), .B1(n26700), .B2(
        data_in[6]), .ZN(n13157) );
  INV_X1 U7777 ( .A(n13158), .ZN(n22659) );
  AOI22_X1 U7778 ( .A1(\mem[430][7] ), .A2(n13151), .B1(n26700), .B2(
        data_in[7]), .ZN(n13158) );
  INV_X1 U7779 ( .A(n13159), .ZN(n22658) );
  AOI22_X1 U7780 ( .A1(\mem[431][0] ), .A2(n13160), .B1(n26699), .B2(
        data_in[0]), .ZN(n13159) );
  INV_X1 U7781 ( .A(n13161), .ZN(n22657) );
  AOI22_X1 U7782 ( .A1(\mem[431][1] ), .A2(n13160), .B1(n26699), .B2(
        data_in[1]), .ZN(n13161) );
  INV_X1 U7783 ( .A(n13162), .ZN(n22656) );
  AOI22_X1 U7784 ( .A1(\mem[431][2] ), .A2(n13160), .B1(n26699), .B2(
        data_in[2]), .ZN(n13162) );
  INV_X1 U7785 ( .A(n13163), .ZN(n22655) );
  AOI22_X1 U7786 ( .A1(\mem[431][3] ), .A2(n13160), .B1(n26699), .B2(
        data_in[3]), .ZN(n13163) );
  INV_X1 U7787 ( .A(n13164), .ZN(n22654) );
  AOI22_X1 U7788 ( .A1(\mem[431][4] ), .A2(n13160), .B1(n26699), .B2(
        data_in[4]), .ZN(n13164) );
  INV_X1 U7789 ( .A(n13165), .ZN(n22653) );
  AOI22_X1 U7790 ( .A1(\mem[431][5] ), .A2(n13160), .B1(n26699), .B2(
        data_in[5]), .ZN(n13165) );
  INV_X1 U7791 ( .A(n13166), .ZN(n22652) );
  AOI22_X1 U7792 ( .A1(\mem[431][6] ), .A2(n13160), .B1(n26699), .B2(
        data_in[6]), .ZN(n13166) );
  INV_X1 U7793 ( .A(n13167), .ZN(n22651) );
  AOI22_X1 U7794 ( .A1(\mem[431][7] ), .A2(n13160), .B1(n26699), .B2(
        data_in[7]), .ZN(n13167) );
  INV_X1 U7795 ( .A(n13168), .ZN(n22650) );
  AOI22_X1 U7796 ( .A1(\mem[432][0] ), .A2(n13169), .B1(n26698), .B2(
        data_in[0]), .ZN(n13168) );
  INV_X1 U7797 ( .A(n13170), .ZN(n22649) );
  AOI22_X1 U7798 ( .A1(\mem[432][1] ), .A2(n13169), .B1(n26698), .B2(
        data_in[1]), .ZN(n13170) );
  INV_X1 U7799 ( .A(n13171), .ZN(n22648) );
  AOI22_X1 U7800 ( .A1(\mem[432][2] ), .A2(n13169), .B1(n26698), .B2(
        data_in[2]), .ZN(n13171) );
  INV_X1 U7801 ( .A(n13172), .ZN(n22647) );
  AOI22_X1 U7802 ( .A1(\mem[432][3] ), .A2(n13169), .B1(n26698), .B2(
        data_in[3]), .ZN(n13172) );
  INV_X1 U7803 ( .A(n13173), .ZN(n22646) );
  AOI22_X1 U7804 ( .A1(\mem[432][4] ), .A2(n13169), .B1(n26698), .B2(
        data_in[4]), .ZN(n13173) );
  INV_X1 U7805 ( .A(n13174), .ZN(n22645) );
  AOI22_X1 U7806 ( .A1(\mem[432][5] ), .A2(n13169), .B1(n26698), .B2(
        data_in[5]), .ZN(n13174) );
  INV_X1 U7807 ( .A(n13175), .ZN(n22644) );
  AOI22_X1 U7808 ( .A1(\mem[432][6] ), .A2(n13169), .B1(n26698), .B2(
        data_in[6]), .ZN(n13175) );
  INV_X1 U7809 ( .A(n13176), .ZN(n22643) );
  AOI22_X1 U7810 ( .A1(\mem[432][7] ), .A2(n13169), .B1(n26698), .B2(
        data_in[7]), .ZN(n13176) );
  INV_X1 U7811 ( .A(n13177), .ZN(n22642) );
  AOI22_X1 U7812 ( .A1(\mem[433][0] ), .A2(n13178), .B1(n26697), .B2(
        data_in[0]), .ZN(n13177) );
  INV_X1 U7813 ( .A(n13179), .ZN(n22641) );
  AOI22_X1 U7814 ( .A1(\mem[433][1] ), .A2(n13178), .B1(n26697), .B2(
        data_in[1]), .ZN(n13179) );
  INV_X1 U7815 ( .A(n13180), .ZN(n22640) );
  AOI22_X1 U7816 ( .A1(\mem[433][2] ), .A2(n13178), .B1(n26697), .B2(
        data_in[2]), .ZN(n13180) );
  INV_X1 U7817 ( .A(n13181), .ZN(n22639) );
  AOI22_X1 U7818 ( .A1(\mem[433][3] ), .A2(n13178), .B1(n26697), .B2(
        data_in[3]), .ZN(n13181) );
  INV_X1 U7819 ( .A(n13182), .ZN(n22638) );
  AOI22_X1 U7820 ( .A1(\mem[433][4] ), .A2(n13178), .B1(n26697), .B2(
        data_in[4]), .ZN(n13182) );
  INV_X1 U7821 ( .A(n13183), .ZN(n22637) );
  AOI22_X1 U7822 ( .A1(\mem[433][5] ), .A2(n13178), .B1(n26697), .B2(
        data_in[5]), .ZN(n13183) );
  INV_X1 U7823 ( .A(n13184), .ZN(n22636) );
  AOI22_X1 U7824 ( .A1(\mem[433][6] ), .A2(n13178), .B1(n26697), .B2(
        data_in[6]), .ZN(n13184) );
  INV_X1 U7825 ( .A(n13185), .ZN(n22635) );
  AOI22_X1 U7826 ( .A1(\mem[433][7] ), .A2(n13178), .B1(n26697), .B2(
        data_in[7]), .ZN(n13185) );
  INV_X1 U7827 ( .A(n13186), .ZN(n22634) );
  AOI22_X1 U7828 ( .A1(\mem[434][0] ), .A2(n13187), .B1(n26696), .B2(
        data_in[0]), .ZN(n13186) );
  INV_X1 U7829 ( .A(n13188), .ZN(n22633) );
  AOI22_X1 U7830 ( .A1(\mem[434][1] ), .A2(n13187), .B1(n26696), .B2(
        data_in[1]), .ZN(n13188) );
  INV_X1 U7831 ( .A(n13189), .ZN(n22632) );
  AOI22_X1 U7832 ( .A1(\mem[434][2] ), .A2(n13187), .B1(n26696), .B2(
        data_in[2]), .ZN(n13189) );
  INV_X1 U7833 ( .A(n13190), .ZN(n22631) );
  AOI22_X1 U7834 ( .A1(\mem[434][3] ), .A2(n13187), .B1(n26696), .B2(
        data_in[3]), .ZN(n13190) );
  INV_X1 U7835 ( .A(n13191), .ZN(n22630) );
  AOI22_X1 U7836 ( .A1(\mem[434][4] ), .A2(n13187), .B1(n26696), .B2(
        data_in[4]), .ZN(n13191) );
  INV_X1 U7837 ( .A(n13192), .ZN(n22629) );
  AOI22_X1 U7838 ( .A1(\mem[434][5] ), .A2(n13187), .B1(n26696), .B2(
        data_in[5]), .ZN(n13192) );
  INV_X1 U7839 ( .A(n13193), .ZN(n22628) );
  AOI22_X1 U7840 ( .A1(\mem[434][6] ), .A2(n13187), .B1(n26696), .B2(
        data_in[6]), .ZN(n13193) );
  INV_X1 U7841 ( .A(n13194), .ZN(n22627) );
  AOI22_X1 U7842 ( .A1(\mem[434][7] ), .A2(n13187), .B1(n26696), .B2(
        data_in[7]), .ZN(n13194) );
  INV_X1 U7843 ( .A(n13195), .ZN(n22626) );
  AOI22_X1 U7844 ( .A1(\mem[435][0] ), .A2(n13196), .B1(n26695), .B2(
        data_in[0]), .ZN(n13195) );
  INV_X1 U7845 ( .A(n13197), .ZN(n22625) );
  AOI22_X1 U7846 ( .A1(\mem[435][1] ), .A2(n13196), .B1(n26695), .B2(
        data_in[1]), .ZN(n13197) );
  INV_X1 U7847 ( .A(n13198), .ZN(n22624) );
  AOI22_X1 U7848 ( .A1(\mem[435][2] ), .A2(n13196), .B1(n26695), .B2(
        data_in[2]), .ZN(n13198) );
  INV_X1 U7849 ( .A(n13199), .ZN(n22623) );
  AOI22_X1 U7850 ( .A1(\mem[435][3] ), .A2(n13196), .B1(n26695), .B2(
        data_in[3]), .ZN(n13199) );
  INV_X1 U7851 ( .A(n13200), .ZN(n22622) );
  AOI22_X1 U7852 ( .A1(\mem[435][4] ), .A2(n13196), .B1(n26695), .B2(
        data_in[4]), .ZN(n13200) );
  INV_X1 U7853 ( .A(n13201), .ZN(n22621) );
  AOI22_X1 U7854 ( .A1(\mem[435][5] ), .A2(n13196), .B1(n26695), .B2(
        data_in[5]), .ZN(n13201) );
  INV_X1 U7855 ( .A(n13202), .ZN(n22620) );
  AOI22_X1 U7856 ( .A1(\mem[435][6] ), .A2(n13196), .B1(n26695), .B2(
        data_in[6]), .ZN(n13202) );
  INV_X1 U7857 ( .A(n13203), .ZN(n22619) );
  AOI22_X1 U7858 ( .A1(\mem[435][7] ), .A2(n13196), .B1(n26695), .B2(
        data_in[7]), .ZN(n13203) );
  INV_X1 U7859 ( .A(n13204), .ZN(n22618) );
  AOI22_X1 U7860 ( .A1(\mem[436][0] ), .A2(n13205), .B1(n26694), .B2(
        data_in[0]), .ZN(n13204) );
  INV_X1 U7861 ( .A(n13206), .ZN(n22617) );
  AOI22_X1 U7862 ( .A1(\mem[436][1] ), .A2(n13205), .B1(n26694), .B2(
        data_in[1]), .ZN(n13206) );
  INV_X1 U7863 ( .A(n13207), .ZN(n22616) );
  AOI22_X1 U7864 ( .A1(\mem[436][2] ), .A2(n13205), .B1(n26694), .B2(
        data_in[2]), .ZN(n13207) );
  INV_X1 U7865 ( .A(n13208), .ZN(n22615) );
  AOI22_X1 U7866 ( .A1(\mem[436][3] ), .A2(n13205), .B1(n26694), .B2(
        data_in[3]), .ZN(n13208) );
  INV_X1 U7867 ( .A(n13209), .ZN(n22614) );
  AOI22_X1 U7868 ( .A1(\mem[436][4] ), .A2(n13205), .B1(n26694), .B2(
        data_in[4]), .ZN(n13209) );
  INV_X1 U7869 ( .A(n13210), .ZN(n22613) );
  AOI22_X1 U7870 ( .A1(\mem[436][5] ), .A2(n13205), .B1(n26694), .B2(
        data_in[5]), .ZN(n13210) );
  INV_X1 U7871 ( .A(n13211), .ZN(n22612) );
  AOI22_X1 U7872 ( .A1(\mem[436][6] ), .A2(n13205), .B1(n26694), .B2(
        data_in[6]), .ZN(n13211) );
  INV_X1 U7873 ( .A(n13212), .ZN(n22611) );
  AOI22_X1 U7874 ( .A1(\mem[436][7] ), .A2(n13205), .B1(n26694), .B2(
        data_in[7]), .ZN(n13212) );
  INV_X1 U7875 ( .A(n13213), .ZN(n22610) );
  AOI22_X1 U7876 ( .A1(\mem[437][0] ), .A2(n13214), .B1(n26693), .B2(
        data_in[0]), .ZN(n13213) );
  INV_X1 U7877 ( .A(n13215), .ZN(n22609) );
  AOI22_X1 U7878 ( .A1(\mem[437][1] ), .A2(n13214), .B1(n26693), .B2(
        data_in[1]), .ZN(n13215) );
  INV_X1 U7879 ( .A(n13216), .ZN(n22608) );
  AOI22_X1 U7880 ( .A1(\mem[437][2] ), .A2(n13214), .B1(n26693), .B2(
        data_in[2]), .ZN(n13216) );
  INV_X1 U7881 ( .A(n13217), .ZN(n22607) );
  AOI22_X1 U7882 ( .A1(\mem[437][3] ), .A2(n13214), .B1(n26693), .B2(
        data_in[3]), .ZN(n13217) );
  INV_X1 U7883 ( .A(n13218), .ZN(n22606) );
  AOI22_X1 U7884 ( .A1(\mem[437][4] ), .A2(n13214), .B1(n26693), .B2(
        data_in[4]), .ZN(n13218) );
  INV_X1 U7885 ( .A(n13219), .ZN(n22605) );
  AOI22_X1 U7886 ( .A1(\mem[437][5] ), .A2(n13214), .B1(n26693), .B2(
        data_in[5]), .ZN(n13219) );
  INV_X1 U7887 ( .A(n13220), .ZN(n22604) );
  AOI22_X1 U7888 ( .A1(\mem[437][6] ), .A2(n13214), .B1(n26693), .B2(
        data_in[6]), .ZN(n13220) );
  INV_X1 U7889 ( .A(n13221), .ZN(n22603) );
  AOI22_X1 U7890 ( .A1(\mem[437][7] ), .A2(n13214), .B1(n26693), .B2(
        data_in[7]), .ZN(n13221) );
  INV_X1 U7891 ( .A(n13222), .ZN(n22602) );
  AOI22_X1 U7892 ( .A1(\mem[438][0] ), .A2(n13223), .B1(n26692), .B2(
        data_in[0]), .ZN(n13222) );
  INV_X1 U7893 ( .A(n13224), .ZN(n22601) );
  AOI22_X1 U7894 ( .A1(\mem[438][1] ), .A2(n13223), .B1(n26692), .B2(
        data_in[1]), .ZN(n13224) );
  INV_X1 U7895 ( .A(n13225), .ZN(n22600) );
  AOI22_X1 U7896 ( .A1(\mem[438][2] ), .A2(n13223), .B1(n26692), .B2(
        data_in[2]), .ZN(n13225) );
  INV_X1 U7897 ( .A(n13226), .ZN(n22599) );
  AOI22_X1 U7898 ( .A1(\mem[438][3] ), .A2(n13223), .B1(n26692), .B2(
        data_in[3]), .ZN(n13226) );
  INV_X1 U7899 ( .A(n13227), .ZN(n22598) );
  AOI22_X1 U7900 ( .A1(\mem[438][4] ), .A2(n13223), .B1(n26692), .B2(
        data_in[4]), .ZN(n13227) );
  INV_X1 U7901 ( .A(n13228), .ZN(n22597) );
  AOI22_X1 U7902 ( .A1(\mem[438][5] ), .A2(n13223), .B1(n26692), .B2(
        data_in[5]), .ZN(n13228) );
  INV_X1 U7903 ( .A(n13229), .ZN(n22596) );
  AOI22_X1 U7904 ( .A1(\mem[438][6] ), .A2(n13223), .B1(n26692), .B2(
        data_in[6]), .ZN(n13229) );
  INV_X1 U7905 ( .A(n13230), .ZN(n22595) );
  AOI22_X1 U7906 ( .A1(\mem[438][7] ), .A2(n13223), .B1(n26692), .B2(
        data_in[7]), .ZN(n13230) );
  INV_X1 U7907 ( .A(n13231), .ZN(n22594) );
  AOI22_X1 U7908 ( .A1(\mem[439][0] ), .A2(n13232), .B1(n26691), .B2(
        data_in[0]), .ZN(n13231) );
  INV_X1 U7909 ( .A(n13233), .ZN(n22593) );
  AOI22_X1 U7910 ( .A1(\mem[439][1] ), .A2(n13232), .B1(n26691), .B2(
        data_in[1]), .ZN(n13233) );
  INV_X1 U7911 ( .A(n13234), .ZN(n22592) );
  AOI22_X1 U7912 ( .A1(\mem[439][2] ), .A2(n13232), .B1(n26691), .B2(
        data_in[2]), .ZN(n13234) );
  INV_X1 U7913 ( .A(n13235), .ZN(n22591) );
  AOI22_X1 U7914 ( .A1(\mem[439][3] ), .A2(n13232), .B1(n26691), .B2(
        data_in[3]), .ZN(n13235) );
  INV_X1 U7915 ( .A(n13236), .ZN(n22590) );
  AOI22_X1 U7916 ( .A1(\mem[439][4] ), .A2(n13232), .B1(n26691), .B2(
        data_in[4]), .ZN(n13236) );
  INV_X1 U7917 ( .A(n13237), .ZN(n22589) );
  AOI22_X1 U7918 ( .A1(\mem[439][5] ), .A2(n13232), .B1(n26691), .B2(
        data_in[5]), .ZN(n13237) );
  INV_X1 U7919 ( .A(n13238), .ZN(n22588) );
  AOI22_X1 U7920 ( .A1(\mem[439][6] ), .A2(n13232), .B1(n26691), .B2(
        data_in[6]), .ZN(n13238) );
  INV_X1 U7921 ( .A(n13239), .ZN(n22587) );
  AOI22_X1 U7922 ( .A1(\mem[439][7] ), .A2(n13232), .B1(n26691), .B2(
        data_in[7]), .ZN(n13239) );
  INV_X1 U7923 ( .A(n13240), .ZN(n22586) );
  AOI22_X1 U7924 ( .A1(\mem[440][0] ), .A2(n13241), .B1(n26690), .B2(
        data_in[0]), .ZN(n13240) );
  INV_X1 U7925 ( .A(n13242), .ZN(n22585) );
  AOI22_X1 U7926 ( .A1(\mem[440][1] ), .A2(n13241), .B1(n26690), .B2(
        data_in[1]), .ZN(n13242) );
  INV_X1 U7927 ( .A(n13243), .ZN(n22584) );
  AOI22_X1 U7928 ( .A1(\mem[440][2] ), .A2(n13241), .B1(n26690), .B2(
        data_in[2]), .ZN(n13243) );
  INV_X1 U7929 ( .A(n13244), .ZN(n22583) );
  AOI22_X1 U7930 ( .A1(\mem[440][3] ), .A2(n13241), .B1(n26690), .B2(
        data_in[3]), .ZN(n13244) );
  INV_X1 U7931 ( .A(n13245), .ZN(n22582) );
  AOI22_X1 U7932 ( .A1(\mem[440][4] ), .A2(n13241), .B1(n26690), .B2(
        data_in[4]), .ZN(n13245) );
  INV_X1 U7933 ( .A(n13246), .ZN(n22581) );
  AOI22_X1 U7934 ( .A1(\mem[440][5] ), .A2(n13241), .B1(n26690), .B2(
        data_in[5]), .ZN(n13246) );
  INV_X1 U7935 ( .A(n13247), .ZN(n22580) );
  AOI22_X1 U7936 ( .A1(\mem[440][6] ), .A2(n13241), .B1(n26690), .B2(
        data_in[6]), .ZN(n13247) );
  INV_X1 U7937 ( .A(n13248), .ZN(n22579) );
  AOI22_X1 U7938 ( .A1(\mem[440][7] ), .A2(n13241), .B1(n26690), .B2(
        data_in[7]), .ZN(n13248) );
  INV_X1 U7939 ( .A(n13249), .ZN(n22578) );
  AOI22_X1 U7940 ( .A1(\mem[441][0] ), .A2(n13250), .B1(n26689), .B2(
        data_in[0]), .ZN(n13249) );
  INV_X1 U7941 ( .A(n13251), .ZN(n22577) );
  AOI22_X1 U7942 ( .A1(\mem[441][1] ), .A2(n13250), .B1(n26689), .B2(
        data_in[1]), .ZN(n13251) );
  INV_X1 U7943 ( .A(n13252), .ZN(n22576) );
  AOI22_X1 U7944 ( .A1(\mem[441][2] ), .A2(n13250), .B1(n26689), .B2(
        data_in[2]), .ZN(n13252) );
  INV_X1 U7945 ( .A(n13253), .ZN(n22575) );
  AOI22_X1 U7946 ( .A1(\mem[441][3] ), .A2(n13250), .B1(n26689), .B2(
        data_in[3]), .ZN(n13253) );
  INV_X1 U7947 ( .A(n13254), .ZN(n22574) );
  AOI22_X1 U7948 ( .A1(\mem[441][4] ), .A2(n13250), .B1(n26689), .B2(
        data_in[4]), .ZN(n13254) );
  INV_X1 U7949 ( .A(n13255), .ZN(n22573) );
  AOI22_X1 U7950 ( .A1(\mem[441][5] ), .A2(n13250), .B1(n26689), .B2(
        data_in[5]), .ZN(n13255) );
  INV_X1 U7951 ( .A(n13256), .ZN(n22572) );
  AOI22_X1 U7952 ( .A1(\mem[441][6] ), .A2(n13250), .B1(n26689), .B2(
        data_in[6]), .ZN(n13256) );
  INV_X1 U7953 ( .A(n13257), .ZN(n22571) );
  AOI22_X1 U7954 ( .A1(\mem[441][7] ), .A2(n13250), .B1(n26689), .B2(
        data_in[7]), .ZN(n13257) );
  INV_X1 U7955 ( .A(n13258), .ZN(n22570) );
  AOI22_X1 U7956 ( .A1(\mem[442][0] ), .A2(n13259), .B1(n26688), .B2(
        data_in[0]), .ZN(n13258) );
  INV_X1 U7957 ( .A(n13260), .ZN(n22569) );
  AOI22_X1 U7958 ( .A1(\mem[442][1] ), .A2(n13259), .B1(n26688), .B2(
        data_in[1]), .ZN(n13260) );
  INV_X1 U7959 ( .A(n13261), .ZN(n22568) );
  AOI22_X1 U7960 ( .A1(\mem[442][2] ), .A2(n13259), .B1(n26688), .B2(
        data_in[2]), .ZN(n13261) );
  INV_X1 U7961 ( .A(n13262), .ZN(n22567) );
  AOI22_X1 U7962 ( .A1(\mem[442][3] ), .A2(n13259), .B1(n26688), .B2(
        data_in[3]), .ZN(n13262) );
  INV_X1 U7963 ( .A(n13263), .ZN(n22566) );
  AOI22_X1 U7964 ( .A1(\mem[442][4] ), .A2(n13259), .B1(n26688), .B2(
        data_in[4]), .ZN(n13263) );
  INV_X1 U7965 ( .A(n13264), .ZN(n22565) );
  AOI22_X1 U7966 ( .A1(\mem[442][5] ), .A2(n13259), .B1(n26688), .B2(
        data_in[5]), .ZN(n13264) );
  INV_X1 U7967 ( .A(n13265), .ZN(n22564) );
  AOI22_X1 U7968 ( .A1(\mem[442][6] ), .A2(n13259), .B1(n26688), .B2(
        data_in[6]), .ZN(n13265) );
  INV_X1 U7969 ( .A(n13266), .ZN(n22563) );
  AOI22_X1 U7970 ( .A1(\mem[442][7] ), .A2(n13259), .B1(n26688), .B2(
        data_in[7]), .ZN(n13266) );
  INV_X1 U7971 ( .A(n13267), .ZN(n22562) );
  AOI22_X1 U7972 ( .A1(\mem[443][0] ), .A2(n13268), .B1(n26687), .B2(
        data_in[0]), .ZN(n13267) );
  INV_X1 U7973 ( .A(n13269), .ZN(n22561) );
  AOI22_X1 U7974 ( .A1(\mem[443][1] ), .A2(n13268), .B1(n26687), .B2(
        data_in[1]), .ZN(n13269) );
  INV_X1 U7975 ( .A(n13270), .ZN(n22560) );
  AOI22_X1 U7976 ( .A1(\mem[443][2] ), .A2(n13268), .B1(n26687), .B2(
        data_in[2]), .ZN(n13270) );
  INV_X1 U7977 ( .A(n13271), .ZN(n22559) );
  AOI22_X1 U7978 ( .A1(\mem[443][3] ), .A2(n13268), .B1(n26687), .B2(
        data_in[3]), .ZN(n13271) );
  INV_X1 U7979 ( .A(n13272), .ZN(n22558) );
  AOI22_X1 U7980 ( .A1(\mem[443][4] ), .A2(n13268), .B1(n26687), .B2(
        data_in[4]), .ZN(n13272) );
  INV_X1 U7981 ( .A(n13273), .ZN(n22557) );
  AOI22_X1 U7982 ( .A1(\mem[443][5] ), .A2(n13268), .B1(n26687), .B2(
        data_in[5]), .ZN(n13273) );
  INV_X1 U7983 ( .A(n13274), .ZN(n22556) );
  AOI22_X1 U7984 ( .A1(\mem[443][6] ), .A2(n13268), .B1(n26687), .B2(
        data_in[6]), .ZN(n13274) );
  INV_X1 U7985 ( .A(n13275), .ZN(n22555) );
  AOI22_X1 U7986 ( .A1(\mem[443][7] ), .A2(n13268), .B1(n26687), .B2(
        data_in[7]), .ZN(n13275) );
  INV_X1 U7987 ( .A(n13276), .ZN(n22554) );
  AOI22_X1 U7988 ( .A1(\mem[444][0] ), .A2(n13277), .B1(n26686), .B2(
        data_in[0]), .ZN(n13276) );
  INV_X1 U7989 ( .A(n13278), .ZN(n22553) );
  AOI22_X1 U7990 ( .A1(\mem[444][1] ), .A2(n13277), .B1(n26686), .B2(
        data_in[1]), .ZN(n13278) );
  INV_X1 U7991 ( .A(n13279), .ZN(n22552) );
  AOI22_X1 U7992 ( .A1(\mem[444][2] ), .A2(n13277), .B1(n26686), .B2(
        data_in[2]), .ZN(n13279) );
  INV_X1 U7993 ( .A(n13280), .ZN(n22551) );
  AOI22_X1 U7994 ( .A1(\mem[444][3] ), .A2(n13277), .B1(n26686), .B2(
        data_in[3]), .ZN(n13280) );
  INV_X1 U7995 ( .A(n13281), .ZN(n22550) );
  AOI22_X1 U7996 ( .A1(\mem[444][4] ), .A2(n13277), .B1(n26686), .B2(
        data_in[4]), .ZN(n13281) );
  INV_X1 U7997 ( .A(n13282), .ZN(n22549) );
  AOI22_X1 U7998 ( .A1(\mem[444][5] ), .A2(n13277), .B1(n26686), .B2(
        data_in[5]), .ZN(n13282) );
  INV_X1 U7999 ( .A(n13283), .ZN(n22548) );
  AOI22_X1 U8000 ( .A1(\mem[444][6] ), .A2(n13277), .B1(n26686), .B2(
        data_in[6]), .ZN(n13283) );
  INV_X1 U8001 ( .A(n13284), .ZN(n22547) );
  AOI22_X1 U8002 ( .A1(\mem[444][7] ), .A2(n13277), .B1(n26686), .B2(
        data_in[7]), .ZN(n13284) );
  INV_X1 U8003 ( .A(n13285), .ZN(n22546) );
  AOI22_X1 U8004 ( .A1(\mem[445][0] ), .A2(n13286), .B1(n26685), .B2(
        data_in[0]), .ZN(n13285) );
  INV_X1 U8005 ( .A(n13287), .ZN(n22545) );
  AOI22_X1 U8006 ( .A1(\mem[445][1] ), .A2(n13286), .B1(n26685), .B2(
        data_in[1]), .ZN(n13287) );
  INV_X1 U8007 ( .A(n13288), .ZN(n22544) );
  AOI22_X1 U8008 ( .A1(\mem[445][2] ), .A2(n13286), .B1(n26685), .B2(
        data_in[2]), .ZN(n13288) );
  INV_X1 U8009 ( .A(n13289), .ZN(n22543) );
  AOI22_X1 U8010 ( .A1(\mem[445][3] ), .A2(n13286), .B1(n26685), .B2(
        data_in[3]), .ZN(n13289) );
  INV_X1 U8011 ( .A(n13290), .ZN(n22542) );
  AOI22_X1 U8012 ( .A1(\mem[445][4] ), .A2(n13286), .B1(n26685), .B2(
        data_in[4]), .ZN(n13290) );
  INV_X1 U8013 ( .A(n13291), .ZN(n22541) );
  AOI22_X1 U8014 ( .A1(\mem[445][5] ), .A2(n13286), .B1(n26685), .B2(
        data_in[5]), .ZN(n13291) );
  INV_X1 U8015 ( .A(n13292), .ZN(n22540) );
  AOI22_X1 U8016 ( .A1(\mem[445][6] ), .A2(n13286), .B1(n26685), .B2(
        data_in[6]), .ZN(n13292) );
  INV_X1 U8017 ( .A(n13293), .ZN(n22539) );
  AOI22_X1 U8018 ( .A1(\mem[445][7] ), .A2(n13286), .B1(n26685), .B2(
        data_in[7]), .ZN(n13293) );
  INV_X1 U8019 ( .A(n13294), .ZN(n22538) );
  AOI22_X1 U8020 ( .A1(\mem[446][0] ), .A2(n13295), .B1(n26684), .B2(
        data_in[0]), .ZN(n13294) );
  INV_X1 U8021 ( .A(n13296), .ZN(n22537) );
  AOI22_X1 U8022 ( .A1(\mem[446][1] ), .A2(n13295), .B1(n26684), .B2(
        data_in[1]), .ZN(n13296) );
  INV_X1 U8023 ( .A(n13297), .ZN(n22536) );
  AOI22_X1 U8024 ( .A1(\mem[446][2] ), .A2(n13295), .B1(n26684), .B2(
        data_in[2]), .ZN(n13297) );
  INV_X1 U8025 ( .A(n13298), .ZN(n22535) );
  AOI22_X1 U8026 ( .A1(\mem[446][3] ), .A2(n13295), .B1(n26684), .B2(
        data_in[3]), .ZN(n13298) );
  INV_X1 U8027 ( .A(n13299), .ZN(n22534) );
  AOI22_X1 U8028 ( .A1(\mem[446][4] ), .A2(n13295), .B1(n26684), .B2(
        data_in[4]), .ZN(n13299) );
  INV_X1 U8029 ( .A(n13300), .ZN(n22533) );
  AOI22_X1 U8030 ( .A1(\mem[446][5] ), .A2(n13295), .B1(n26684), .B2(
        data_in[5]), .ZN(n13300) );
  INV_X1 U8031 ( .A(n13301), .ZN(n22532) );
  AOI22_X1 U8032 ( .A1(\mem[446][6] ), .A2(n13295), .B1(n26684), .B2(
        data_in[6]), .ZN(n13301) );
  INV_X1 U8033 ( .A(n13302), .ZN(n22531) );
  AOI22_X1 U8034 ( .A1(\mem[446][7] ), .A2(n13295), .B1(n26684), .B2(
        data_in[7]), .ZN(n13302) );
  INV_X1 U8035 ( .A(n13303), .ZN(n22530) );
  AOI22_X1 U8036 ( .A1(\mem[447][0] ), .A2(n13304), .B1(n26683), .B2(
        data_in[0]), .ZN(n13303) );
  INV_X1 U8037 ( .A(n13305), .ZN(n22529) );
  AOI22_X1 U8038 ( .A1(\mem[447][1] ), .A2(n13304), .B1(n26683), .B2(
        data_in[1]), .ZN(n13305) );
  INV_X1 U8039 ( .A(n13306), .ZN(n22528) );
  AOI22_X1 U8040 ( .A1(\mem[447][2] ), .A2(n13304), .B1(n26683), .B2(
        data_in[2]), .ZN(n13306) );
  INV_X1 U8041 ( .A(n13307), .ZN(n22527) );
  AOI22_X1 U8042 ( .A1(\mem[447][3] ), .A2(n13304), .B1(n26683), .B2(
        data_in[3]), .ZN(n13307) );
  INV_X1 U8043 ( .A(n13308), .ZN(n22526) );
  AOI22_X1 U8044 ( .A1(\mem[447][4] ), .A2(n13304), .B1(n26683), .B2(
        data_in[4]), .ZN(n13308) );
  INV_X1 U8045 ( .A(n13309), .ZN(n22525) );
  AOI22_X1 U8046 ( .A1(\mem[447][5] ), .A2(n13304), .B1(n26683), .B2(
        data_in[5]), .ZN(n13309) );
  INV_X1 U8047 ( .A(n13310), .ZN(n22524) );
  AOI22_X1 U8048 ( .A1(\mem[447][6] ), .A2(n13304), .B1(n26683), .B2(
        data_in[6]), .ZN(n13310) );
  INV_X1 U8049 ( .A(n13311), .ZN(n22523) );
  AOI22_X1 U8050 ( .A1(\mem[447][7] ), .A2(n13304), .B1(n26683), .B2(
        data_in[7]), .ZN(n13311) );
  INV_X1 U8051 ( .A(n13385), .ZN(n22458) );
  AOI22_X1 U8052 ( .A1(\mem[456][0] ), .A2(n13386), .B1(n26674), .B2(
        data_in[0]), .ZN(n13385) );
  INV_X1 U8053 ( .A(n13387), .ZN(n22457) );
  AOI22_X1 U8054 ( .A1(\mem[456][1] ), .A2(n13386), .B1(n26674), .B2(
        data_in[1]), .ZN(n13387) );
  INV_X1 U8055 ( .A(n13388), .ZN(n22456) );
  AOI22_X1 U8056 ( .A1(\mem[456][2] ), .A2(n13386), .B1(n26674), .B2(
        data_in[2]), .ZN(n13388) );
  INV_X1 U8057 ( .A(n13389), .ZN(n22455) );
  AOI22_X1 U8058 ( .A1(\mem[456][3] ), .A2(n13386), .B1(n26674), .B2(
        data_in[3]), .ZN(n13389) );
  INV_X1 U8059 ( .A(n13390), .ZN(n22454) );
  AOI22_X1 U8060 ( .A1(\mem[456][4] ), .A2(n13386), .B1(n26674), .B2(
        data_in[4]), .ZN(n13390) );
  INV_X1 U8061 ( .A(n13391), .ZN(n22453) );
  AOI22_X1 U8062 ( .A1(\mem[456][5] ), .A2(n13386), .B1(n26674), .B2(
        data_in[5]), .ZN(n13391) );
  INV_X1 U8063 ( .A(n13392), .ZN(n22452) );
  AOI22_X1 U8064 ( .A1(\mem[456][6] ), .A2(n13386), .B1(n26674), .B2(
        data_in[6]), .ZN(n13392) );
  INV_X1 U8065 ( .A(n13393), .ZN(n22451) );
  AOI22_X1 U8066 ( .A1(\mem[456][7] ), .A2(n13386), .B1(n26674), .B2(
        data_in[7]), .ZN(n13393) );
  INV_X1 U8067 ( .A(n13394), .ZN(n22450) );
  AOI22_X1 U8068 ( .A1(\mem[457][0] ), .A2(n13395), .B1(n26673), .B2(
        data_in[0]), .ZN(n13394) );
  INV_X1 U8069 ( .A(n13396), .ZN(n22449) );
  AOI22_X1 U8070 ( .A1(\mem[457][1] ), .A2(n13395), .B1(n26673), .B2(
        data_in[1]), .ZN(n13396) );
  INV_X1 U8071 ( .A(n13397), .ZN(n22448) );
  AOI22_X1 U8072 ( .A1(\mem[457][2] ), .A2(n13395), .B1(n26673), .B2(
        data_in[2]), .ZN(n13397) );
  INV_X1 U8073 ( .A(n13398), .ZN(n22447) );
  AOI22_X1 U8074 ( .A1(\mem[457][3] ), .A2(n13395), .B1(n26673), .B2(
        data_in[3]), .ZN(n13398) );
  INV_X1 U8075 ( .A(n13399), .ZN(n22446) );
  AOI22_X1 U8076 ( .A1(\mem[457][4] ), .A2(n13395), .B1(n26673), .B2(
        data_in[4]), .ZN(n13399) );
  INV_X1 U8077 ( .A(n13400), .ZN(n22445) );
  AOI22_X1 U8078 ( .A1(\mem[457][5] ), .A2(n13395), .B1(n26673), .B2(
        data_in[5]), .ZN(n13400) );
  INV_X1 U8079 ( .A(n13401), .ZN(n22444) );
  AOI22_X1 U8080 ( .A1(\mem[457][6] ), .A2(n13395), .B1(n26673), .B2(
        data_in[6]), .ZN(n13401) );
  INV_X1 U8081 ( .A(n13402), .ZN(n22443) );
  AOI22_X1 U8082 ( .A1(\mem[457][7] ), .A2(n13395), .B1(n26673), .B2(
        data_in[7]), .ZN(n13402) );
  INV_X1 U8083 ( .A(n13403), .ZN(n22442) );
  AOI22_X1 U8084 ( .A1(\mem[458][0] ), .A2(n13404), .B1(n26672), .B2(
        data_in[0]), .ZN(n13403) );
  INV_X1 U8085 ( .A(n13405), .ZN(n22441) );
  AOI22_X1 U8086 ( .A1(\mem[458][1] ), .A2(n13404), .B1(n26672), .B2(
        data_in[1]), .ZN(n13405) );
  INV_X1 U8087 ( .A(n13406), .ZN(n22440) );
  AOI22_X1 U8088 ( .A1(\mem[458][2] ), .A2(n13404), .B1(n26672), .B2(
        data_in[2]), .ZN(n13406) );
  INV_X1 U8089 ( .A(n13407), .ZN(n22439) );
  AOI22_X1 U8090 ( .A1(\mem[458][3] ), .A2(n13404), .B1(n26672), .B2(
        data_in[3]), .ZN(n13407) );
  INV_X1 U8091 ( .A(n13408), .ZN(n22438) );
  AOI22_X1 U8092 ( .A1(\mem[458][4] ), .A2(n13404), .B1(n26672), .B2(
        data_in[4]), .ZN(n13408) );
  INV_X1 U8093 ( .A(n13409), .ZN(n22437) );
  AOI22_X1 U8094 ( .A1(\mem[458][5] ), .A2(n13404), .B1(n26672), .B2(
        data_in[5]), .ZN(n13409) );
  INV_X1 U8095 ( .A(n13410), .ZN(n22436) );
  AOI22_X1 U8096 ( .A1(\mem[458][6] ), .A2(n13404), .B1(n26672), .B2(
        data_in[6]), .ZN(n13410) );
  INV_X1 U8097 ( .A(n13411), .ZN(n22435) );
  AOI22_X1 U8098 ( .A1(\mem[458][7] ), .A2(n13404), .B1(n26672), .B2(
        data_in[7]), .ZN(n13411) );
  INV_X1 U8099 ( .A(n13412), .ZN(n22434) );
  AOI22_X1 U8100 ( .A1(\mem[459][0] ), .A2(n13413), .B1(n26671), .B2(
        data_in[0]), .ZN(n13412) );
  INV_X1 U8101 ( .A(n13414), .ZN(n22433) );
  AOI22_X1 U8102 ( .A1(\mem[459][1] ), .A2(n13413), .B1(n26671), .B2(
        data_in[1]), .ZN(n13414) );
  INV_X1 U8103 ( .A(n13415), .ZN(n22432) );
  AOI22_X1 U8104 ( .A1(\mem[459][2] ), .A2(n13413), .B1(n26671), .B2(
        data_in[2]), .ZN(n13415) );
  INV_X1 U8105 ( .A(n13416), .ZN(n22431) );
  AOI22_X1 U8106 ( .A1(\mem[459][3] ), .A2(n13413), .B1(n26671), .B2(
        data_in[3]), .ZN(n13416) );
  INV_X1 U8107 ( .A(n13417), .ZN(n22430) );
  AOI22_X1 U8108 ( .A1(\mem[459][4] ), .A2(n13413), .B1(n26671), .B2(
        data_in[4]), .ZN(n13417) );
  INV_X1 U8109 ( .A(n13418), .ZN(n22429) );
  AOI22_X1 U8110 ( .A1(\mem[459][5] ), .A2(n13413), .B1(n26671), .B2(
        data_in[5]), .ZN(n13418) );
  INV_X1 U8111 ( .A(n13419), .ZN(n22428) );
  AOI22_X1 U8112 ( .A1(\mem[459][6] ), .A2(n13413), .B1(n26671), .B2(
        data_in[6]), .ZN(n13419) );
  INV_X1 U8113 ( .A(n13420), .ZN(n22427) );
  AOI22_X1 U8114 ( .A1(\mem[459][7] ), .A2(n13413), .B1(n26671), .B2(
        data_in[7]), .ZN(n13420) );
  INV_X1 U8115 ( .A(n13421), .ZN(n22426) );
  AOI22_X1 U8116 ( .A1(\mem[460][0] ), .A2(n13422), .B1(n26670), .B2(
        data_in[0]), .ZN(n13421) );
  INV_X1 U8117 ( .A(n13423), .ZN(n22425) );
  AOI22_X1 U8118 ( .A1(\mem[460][1] ), .A2(n13422), .B1(n26670), .B2(
        data_in[1]), .ZN(n13423) );
  INV_X1 U8119 ( .A(n13424), .ZN(n22424) );
  AOI22_X1 U8120 ( .A1(\mem[460][2] ), .A2(n13422), .B1(n26670), .B2(
        data_in[2]), .ZN(n13424) );
  INV_X1 U8121 ( .A(n13425), .ZN(n22423) );
  AOI22_X1 U8122 ( .A1(\mem[460][3] ), .A2(n13422), .B1(n26670), .B2(
        data_in[3]), .ZN(n13425) );
  INV_X1 U8123 ( .A(n13426), .ZN(n22422) );
  AOI22_X1 U8124 ( .A1(\mem[460][4] ), .A2(n13422), .B1(n26670), .B2(
        data_in[4]), .ZN(n13426) );
  INV_X1 U8125 ( .A(n13427), .ZN(n22421) );
  AOI22_X1 U8126 ( .A1(\mem[460][5] ), .A2(n13422), .B1(n26670), .B2(
        data_in[5]), .ZN(n13427) );
  INV_X1 U8127 ( .A(n13428), .ZN(n22420) );
  AOI22_X1 U8128 ( .A1(\mem[460][6] ), .A2(n13422), .B1(n26670), .B2(
        data_in[6]), .ZN(n13428) );
  INV_X1 U8129 ( .A(n13429), .ZN(n22419) );
  AOI22_X1 U8130 ( .A1(\mem[460][7] ), .A2(n13422), .B1(n26670), .B2(
        data_in[7]), .ZN(n13429) );
  INV_X1 U8131 ( .A(n13430), .ZN(n22418) );
  AOI22_X1 U8132 ( .A1(\mem[461][0] ), .A2(n13431), .B1(n26669), .B2(
        data_in[0]), .ZN(n13430) );
  INV_X1 U8133 ( .A(n13432), .ZN(n22417) );
  AOI22_X1 U8134 ( .A1(\mem[461][1] ), .A2(n13431), .B1(n26669), .B2(
        data_in[1]), .ZN(n13432) );
  INV_X1 U8135 ( .A(n13433), .ZN(n22416) );
  AOI22_X1 U8136 ( .A1(\mem[461][2] ), .A2(n13431), .B1(n26669), .B2(
        data_in[2]), .ZN(n13433) );
  INV_X1 U8137 ( .A(n13434), .ZN(n22415) );
  AOI22_X1 U8138 ( .A1(\mem[461][3] ), .A2(n13431), .B1(n26669), .B2(
        data_in[3]), .ZN(n13434) );
  INV_X1 U8139 ( .A(n13435), .ZN(n22414) );
  AOI22_X1 U8140 ( .A1(\mem[461][4] ), .A2(n13431), .B1(n26669), .B2(
        data_in[4]), .ZN(n13435) );
  INV_X1 U8141 ( .A(n13436), .ZN(n22413) );
  AOI22_X1 U8142 ( .A1(\mem[461][5] ), .A2(n13431), .B1(n26669), .B2(
        data_in[5]), .ZN(n13436) );
  INV_X1 U8143 ( .A(n13437), .ZN(n22412) );
  AOI22_X1 U8144 ( .A1(\mem[461][6] ), .A2(n13431), .B1(n26669), .B2(
        data_in[6]), .ZN(n13437) );
  INV_X1 U8145 ( .A(n13438), .ZN(n22411) );
  AOI22_X1 U8146 ( .A1(\mem[461][7] ), .A2(n13431), .B1(n26669), .B2(
        data_in[7]), .ZN(n13438) );
  INV_X1 U8147 ( .A(n13439), .ZN(n22410) );
  AOI22_X1 U8148 ( .A1(\mem[462][0] ), .A2(n13440), .B1(n26668), .B2(
        data_in[0]), .ZN(n13439) );
  INV_X1 U8149 ( .A(n13441), .ZN(n22409) );
  AOI22_X1 U8150 ( .A1(\mem[462][1] ), .A2(n13440), .B1(n26668), .B2(
        data_in[1]), .ZN(n13441) );
  INV_X1 U8151 ( .A(n13442), .ZN(n22408) );
  AOI22_X1 U8152 ( .A1(\mem[462][2] ), .A2(n13440), .B1(n26668), .B2(
        data_in[2]), .ZN(n13442) );
  INV_X1 U8153 ( .A(n13443), .ZN(n22407) );
  AOI22_X1 U8154 ( .A1(\mem[462][3] ), .A2(n13440), .B1(n26668), .B2(
        data_in[3]), .ZN(n13443) );
  INV_X1 U8155 ( .A(n13444), .ZN(n22406) );
  AOI22_X1 U8156 ( .A1(\mem[462][4] ), .A2(n13440), .B1(n26668), .B2(
        data_in[4]), .ZN(n13444) );
  INV_X1 U8157 ( .A(n13445), .ZN(n22405) );
  AOI22_X1 U8158 ( .A1(\mem[462][5] ), .A2(n13440), .B1(n26668), .B2(
        data_in[5]), .ZN(n13445) );
  INV_X1 U8159 ( .A(n13446), .ZN(n22404) );
  AOI22_X1 U8160 ( .A1(\mem[462][6] ), .A2(n13440), .B1(n26668), .B2(
        data_in[6]), .ZN(n13446) );
  INV_X1 U8161 ( .A(n13447), .ZN(n22403) );
  AOI22_X1 U8162 ( .A1(\mem[462][7] ), .A2(n13440), .B1(n26668), .B2(
        data_in[7]), .ZN(n13447) );
  INV_X1 U8163 ( .A(n13448), .ZN(n22402) );
  AOI22_X1 U8164 ( .A1(\mem[463][0] ), .A2(n13449), .B1(n26667), .B2(
        data_in[0]), .ZN(n13448) );
  INV_X1 U8165 ( .A(n13450), .ZN(n22401) );
  AOI22_X1 U8166 ( .A1(\mem[463][1] ), .A2(n13449), .B1(n26667), .B2(
        data_in[1]), .ZN(n13450) );
  INV_X1 U8167 ( .A(n13451), .ZN(n22400) );
  AOI22_X1 U8168 ( .A1(\mem[463][2] ), .A2(n13449), .B1(n26667), .B2(
        data_in[2]), .ZN(n13451) );
  INV_X1 U8169 ( .A(n13452), .ZN(n22399) );
  AOI22_X1 U8170 ( .A1(\mem[463][3] ), .A2(n13449), .B1(n26667), .B2(
        data_in[3]), .ZN(n13452) );
  INV_X1 U8171 ( .A(n13453), .ZN(n22398) );
  AOI22_X1 U8172 ( .A1(\mem[463][4] ), .A2(n13449), .B1(n26667), .B2(
        data_in[4]), .ZN(n13453) );
  INV_X1 U8173 ( .A(n13454), .ZN(n22397) );
  AOI22_X1 U8174 ( .A1(\mem[463][5] ), .A2(n13449), .B1(n26667), .B2(
        data_in[5]), .ZN(n13454) );
  INV_X1 U8175 ( .A(n13455), .ZN(n22396) );
  AOI22_X1 U8176 ( .A1(\mem[463][6] ), .A2(n13449), .B1(n26667), .B2(
        data_in[6]), .ZN(n13455) );
  INV_X1 U8177 ( .A(n13456), .ZN(n22395) );
  AOI22_X1 U8178 ( .A1(\mem[463][7] ), .A2(n13449), .B1(n26667), .B2(
        data_in[7]), .ZN(n13456) );
  INV_X1 U8179 ( .A(n13457), .ZN(n22394) );
  AOI22_X1 U8180 ( .A1(\mem[464][0] ), .A2(n13458), .B1(n26666), .B2(
        data_in[0]), .ZN(n13457) );
  INV_X1 U8181 ( .A(n13459), .ZN(n22393) );
  AOI22_X1 U8182 ( .A1(\mem[464][1] ), .A2(n13458), .B1(n26666), .B2(
        data_in[1]), .ZN(n13459) );
  INV_X1 U8183 ( .A(n13460), .ZN(n22392) );
  AOI22_X1 U8184 ( .A1(\mem[464][2] ), .A2(n13458), .B1(n26666), .B2(
        data_in[2]), .ZN(n13460) );
  INV_X1 U8185 ( .A(n13461), .ZN(n22391) );
  AOI22_X1 U8186 ( .A1(\mem[464][3] ), .A2(n13458), .B1(n26666), .B2(
        data_in[3]), .ZN(n13461) );
  INV_X1 U8187 ( .A(n13462), .ZN(n22390) );
  AOI22_X1 U8188 ( .A1(\mem[464][4] ), .A2(n13458), .B1(n26666), .B2(
        data_in[4]), .ZN(n13462) );
  INV_X1 U8189 ( .A(n13463), .ZN(n22389) );
  AOI22_X1 U8190 ( .A1(\mem[464][5] ), .A2(n13458), .B1(n26666), .B2(
        data_in[5]), .ZN(n13463) );
  INV_X1 U8191 ( .A(n13464), .ZN(n22388) );
  AOI22_X1 U8192 ( .A1(\mem[464][6] ), .A2(n13458), .B1(n26666), .B2(
        data_in[6]), .ZN(n13464) );
  INV_X1 U8193 ( .A(n13465), .ZN(n22387) );
  AOI22_X1 U8194 ( .A1(\mem[464][7] ), .A2(n13458), .B1(n26666), .B2(
        data_in[7]), .ZN(n13465) );
  INV_X1 U8195 ( .A(n13466), .ZN(n22386) );
  AOI22_X1 U8196 ( .A1(\mem[465][0] ), .A2(n13467), .B1(n26665), .B2(
        data_in[0]), .ZN(n13466) );
  INV_X1 U8197 ( .A(n13468), .ZN(n22385) );
  AOI22_X1 U8198 ( .A1(\mem[465][1] ), .A2(n13467), .B1(n26665), .B2(
        data_in[1]), .ZN(n13468) );
  INV_X1 U8199 ( .A(n13469), .ZN(n22384) );
  AOI22_X1 U8200 ( .A1(\mem[465][2] ), .A2(n13467), .B1(n26665), .B2(
        data_in[2]), .ZN(n13469) );
  INV_X1 U8201 ( .A(n13470), .ZN(n22383) );
  AOI22_X1 U8202 ( .A1(\mem[465][3] ), .A2(n13467), .B1(n26665), .B2(
        data_in[3]), .ZN(n13470) );
  INV_X1 U8203 ( .A(n13471), .ZN(n22382) );
  AOI22_X1 U8204 ( .A1(\mem[465][4] ), .A2(n13467), .B1(n26665), .B2(
        data_in[4]), .ZN(n13471) );
  INV_X1 U8205 ( .A(n13472), .ZN(n22381) );
  AOI22_X1 U8206 ( .A1(\mem[465][5] ), .A2(n13467), .B1(n26665), .B2(
        data_in[5]), .ZN(n13472) );
  INV_X1 U8207 ( .A(n13473), .ZN(n22380) );
  AOI22_X1 U8208 ( .A1(\mem[465][6] ), .A2(n13467), .B1(n26665), .B2(
        data_in[6]), .ZN(n13473) );
  INV_X1 U8209 ( .A(n13474), .ZN(n22379) );
  AOI22_X1 U8210 ( .A1(\mem[465][7] ), .A2(n13467), .B1(n26665), .B2(
        data_in[7]), .ZN(n13474) );
  INV_X1 U8211 ( .A(n13475), .ZN(n22378) );
  AOI22_X1 U8212 ( .A1(\mem[466][0] ), .A2(n13476), .B1(n26664), .B2(
        data_in[0]), .ZN(n13475) );
  INV_X1 U8213 ( .A(n13477), .ZN(n22377) );
  AOI22_X1 U8214 ( .A1(\mem[466][1] ), .A2(n13476), .B1(n26664), .B2(
        data_in[1]), .ZN(n13477) );
  INV_X1 U8215 ( .A(n13478), .ZN(n22376) );
  AOI22_X1 U8216 ( .A1(\mem[466][2] ), .A2(n13476), .B1(n26664), .B2(
        data_in[2]), .ZN(n13478) );
  INV_X1 U8217 ( .A(n13479), .ZN(n22375) );
  AOI22_X1 U8218 ( .A1(\mem[466][3] ), .A2(n13476), .B1(n26664), .B2(
        data_in[3]), .ZN(n13479) );
  INV_X1 U8219 ( .A(n13480), .ZN(n22374) );
  AOI22_X1 U8220 ( .A1(\mem[466][4] ), .A2(n13476), .B1(n26664), .B2(
        data_in[4]), .ZN(n13480) );
  INV_X1 U8221 ( .A(n13481), .ZN(n22373) );
  AOI22_X1 U8222 ( .A1(\mem[466][5] ), .A2(n13476), .B1(n26664), .B2(
        data_in[5]), .ZN(n13481) );
  INV_X1 U8223 ( .A(n13482), .ZN(n22372) );
  AOI22_X1 U8224 ( .A1(\mem[466][6] ), .A2(n13476), .B1(n26664), .B2(
        data_in[6]), .ZN(n13482) );
  INV_X1 U8225 ( .A(n13483), .ZN(n22371) );
  AOI22_X1 U8226 ( .A1(\mem[466][7] ), .A2(n13476), .B1(n26664), .B2(
        data_in[7]), .ZN(n13483) );
  INV_X1 U8227 ( .A(n13484), .ZN(n22370) );
  AOI22_X1 U8228 ( .A1(\mem[467][0] ), .A2(n13485), .B1(n26663), .B2(
        data_in[0]), .ZN(n13484) );
  INV_X1 U8229 ( .A(n13486), .ZN(n22369) );
  AOI22_X1 U8230 ( .A1(\mem[467][1] ), .A2(n13485), .B1(n26663), .B2(
        data_in[1]), .ZN(n13486) );
  INV_X1 U8231 ( .A(n13487), .ZN(n22368) );
  AOI22_X1 U8232 ( .A1(\mem[467][2] ), .A2(n13485), .B1(n26663), .B2(
        data_in[2]), .ZN(n13487) );
  INV_X1 U8233 ( .A(n13488), .ZN(n22367) );
  AOI22_X1 U8234 ( .A1(\mem[467][3] ), .A2(n13485), .B1(n26663), .B2(
        data_in[3]), .ZN(n13488) );
  INV_X1 U8235 ( .A(n13489), .ZN(n22366) );
  AOI22_X1 U8236 ( .A1(\mem[467][4] ), .A2(n13485), .B1(n26663), .B2(
        data_in[4]), .ZN(n13489) );
  INV_X1 U8237 ( .A(n13490), .ZN(n22365) );
  AOI22_X1 U8238 ( .A1(\mem[467][5] ), .A2(n13485), .B1(n26663), .B2(
        data_in[5]), .ZN(n13490) );
  INV_X1 U8239 ( .A(n13491), .ZN(n22364) );
  AOI22_X1 U8240 ( .A1(\mem[467][6] ), .A2(n13485), .B1(n26663), .B2(
        data_in[6]), .ZN(n13491) );
  INV_X1 U8241 ( .A(n13492), .ZN(n22363) );
  AOI22_X1 U8242 ( .A1(\mem[467][7] ), .A2(n13485), .B1(n26663), .B2(
        data_in[7]), .ZN(n13492) );
  INV_X1 U8243 ( .A(n13493), .ZN(n22362) );
  AOI22_X1 U8244 ( .A1(\mem[468][0] ), .A2(n13494), .B1(n26662), .B2(
        data_in[0]), .ZN(n13493) );
  INV_X1 U8245 ( .A(n13495), .ZN(n22361) );
  AOI22_X1 U8246 ( .A1(\mem[468][1] ), .A2(n13494), .B1(n26662), .B2(
        data_in[1]), .ZN(n13495) );
  INV_X1 U8247 ( .A(n13496), .ZN(n22360) );
  AOI22_X1 U8248 ( .A1(\mem[468][2] ), .A2(n13494), .B1(n26662), .B2(
        data_in[2]), .ZN(n13496) );
  INV_X1 U8249 ( .A(n13497), .ZN(n22359) );
  AOI22_X1 U8250 ( .A1(\mem[468][3] ), .A2(n13494), .B1(n26662), .B2(
        data_in[3]), .ZN(n13497) );
  INV_X1 U8251 ( .A(n13498), .ZN(n22358) );
  AOI22_X1 U8252 ( .A1(\mem[468][4] ), .A2(n13494), .B1(n26662), .B2(
        data_in[4]), .ZN(n13498) );
  INV_X1 U8253 ( .A(n13499), .ZN(n22357) );
  AOI22_X1 U8254 ( .A1(\mem[468][5] ), .A2(n13494), .B1(n26662), .B2(
        data_in[5]), .ZN(n13499) );
  INV_X1 U8255 ( .A(n13500), .ZN(n22356) );
  AOI22_X1 U8256 ( .A1(\mem[468][6] ), .A2(n13494), .B1(n26662), .B2(
        data_in[6]), .ZN(n13500) );
  INV_X1 U8257 ( .A(n13501), .ZN(n22355) );
  AOI22_X1 U8258 ( .A1(\mem[468][7] ), .A2(n13494), .B1(n26662), .B2(
        data_in[7]), .ZN(n13501) );
  INV_X1 U8259 ( .A(n13502), .ZN(n22354) );
  AOI22_X1 U8260 ( .A1(\mem[469][0] ), .A2(n13503), .B1(n26661), .B2(
        data_in[0]), .ZN(n13502) );
  INV_X1 U8261 ( .A(n13504), .ZN(n22353) );
  AOI22_X1 U8262 ( .A1(\mem[469][1] ), .A2(n13503), .B1(n26661), .B2(
        data_in[1]), .ZN(n13504) );
  INV_X1 U8263 ( .A(n13505), .ZN(n22352) );
  AOI22_X1 U8264 ( .A1(\mem[469][2] ), .A2(n13503), .B1(n26661), .B2(
        data_in[2]), .ZN(n13505) );
  INV_X1 U8265 ( .A(n13506), .ZN(n22351) );
  AOI22_X1 U8266 ( .A1(\mem[469][3] ), .A2(n13503), .B1(n26661), .B2(
        data_in[3]), .ZN(n13506) );
  INV_X1 U8267 ( .A(n13507), .ZN(n22350) );
  AOI22_X1 U8268 ( .A1(\mem[469][4] ), .A2(n13503), .B1(n26661), .B2(
        data_in[4]), .ZN(n13507) );
  INV_X1 U8269 ( .A(n13508), .ZN(n22349) );
  AOI22_X1 U8270 ( .A1(\mem[469][5] ), .A2(n13503), .B1(n26661), .B2(
        data_in[5]), .ZN(n13508) );
  INV_X1 U8271 ( .A(n13509), .ZN(n22348) );
  AOI22_X1 U8272 ( .A1(\mem[469][6] ), .A2(n13503), .B1(n26661), .B2(
        data_in[6]), .ZN(n13509) );
  INV_X1 U8273 ( .A(n13510), .ZN(n22347) );
  AOI22_X1 U8274 ( .A1(\mem[469][7] ), .A2(n13503), .B1(n26661), .B2(
        data_in[7]), .ZN(n13510) );
  INV_X1 U8275 ( .A(n13511), .ZN(n22346) );
  AOI22_X1 U8276 ( .A1(\mem[470][0] ), .A2(n13512), .B1(n26660), .B2(
        data_in[0]), .ZN(n13511) );
  INV_X1 U8277 ( .A(n13513), .ZN(n22345) );
  AOI22_X1 U8278 ( .A1(\mem[470][1] ), .A2(n13512), .B1(n26660), .B2(
        data_in[1]), .ZN(n13513) );
  INV_X1 U8279 ( .A(n13514), .ZN(n22344) );
  AOI22_X1 U8280 ( .A1(\mem[470][2] ), .A2(n13512), .B1(n26660), .B2(
        data_in[2]), .ZN(n13514) );
  INV_X1 U8281 ( .A(n13515), .ZN(n22343) );
  AOI22_X1 U8282 ( .A1(\mem[470][3] ), .A2(n13512), .B1(n26660), .B2(
        data_in[3]), .ZN(n13515) );
  INV_X1 U8283 ( .A(n13516), .ZN(n22342) );
  AOI22_X1 U8284 ( .A1(\mem[470][4] ), .A2(n13512), .B1(n26660), .B2(
        data_in[4]), .ZN(n13516) );
  INV_X1 U8285 ( .A(n13517), .ZN(n22341) );
  AOI22_X1 U8286 ( .A1(\mem[470][5] ), .A2(n13512), .B1(n26660), .B2(
        data_in[5]), .ZN(n13517) );
  INV_X1 U8287 ( .A(n13518), .ZN(n22340) );
  AOI22_X1 U8288 ( .A1(\mem[470][6] ), .A2(n13512), .B1(n26660), .B2(
        data_in[6]), .ZN(n13518) );
  INV_X1 U8289 ( .A(n13519), .ZN(n22339) );
  AOI22_X1 U8290 ( .A1(\mem[470][7] ), .A2(n13512), .B1(n26660), .B2(
        data_in[7]), .ZN(n13519) );
  INV_X1 U8291 ( .A(n13520), .ZN(n22338) );
  AOI22_X1 U8292 ( .A1(\mem[471][0] ), .A2(n13521), .B1(n26659), .B2(
        data_in[0]), .ZN(n13520) );
  INV_X1 U8293 ( .A(n13522), .ZN(n22337) );
  AOI22_X1 U8294 ( .A1(\mem[471][1] ), .A2(n13521), .B1(n26659), .B2(
        data_in[1]), .ZN(n13522) );
  INV_X1 U8295 ( .A(n13523), .ZN(n22336) );
  AOI22_X1 U8296 ( .A1(\mem[471][2] ), .A2(n13521), .B1(n26659), .B2(
        data_in[2]), .ZN(n13523) );
  INV_X1 U8297 ( .A(n13524), .ZN(n22335) );
  AOI22_X1 U8298 ( .A1(\mem[471][3] ), .A2(n13521), .B1(n26659), .B2(
        data_in[3]), .ZN(n13524) );
  INV_X1 U8299 ( .A(n13525), .ZN(n22334) );
  AOI22_X1 U8300 ( .A1(\mem[471][4] ), .A2(n13521), .B1(n26659), .B2(
        data_in[4]), .ZN(n13525) );
  INV_X1 U8301 ( .A(n13526), .ZN(n22333) );
  AOI22_X1 U8302 ( .A1(\mem[471][5] ), .A2(n13521), .B1(n26659), .B2(
        data_in[5]), .ZN(n13526) );
  INV_X1 U8303 ( .A(n13527), .ZN(n22332) );
  AOI22_X1 U8304 ( .A1(\mem[471][6] ), .A2(n13521), .B1(n26659), .B2(
        data_in[6]), .ZN(n13527) );
  INV_X1 U8305 ( .A(n13528), .ZN(n22331) );
  AOI22_X1 U8306 ( .A1(\mem[471][7] ), .A2(n13521), .B1(n26659), .B2(
        data_in[7]), .ZN(n13528) );
  INV_X1 U8307 ( .A(n13529), .ZN(n22330) );
  AOI22_X1 U8308 ( .A1(\mem[472][0] ), .A2(n13530), .B1(n26658), .B2(
        data_in[0]), .ZN(n13529) );
  INV_X1 U8309 ( .A(n13531), .ZN(n22329) );
  AOI22_X1 U8310 ( .A1(\mem[472][1] ), .A2(n13530), .B1(n26658), .B2(
        data_in[1]), .ZN(n13531) );
  INV_X1 U8311 ( .A(n13532), .ZN(n22328) );
  AOI22_X1 U8312 ( .A1(\mem[472][2] ), .A2(n13530), .B1(n26658), .B2(
        data_in[2]), .ZN(n13532) );
  INV_X1 U8313 ( .A(n13533), .ZN(n22327) );
  AOI22_X1 U8314 ( .A1(\mem[472][3] ), .A2(n13530), .B1(n26658), .B2(
        data_in[3]), .ZN(n13533) );
  INV_X1 U8315 ( .A(n13534), .ZN(n22326) );
  AOI22_X1 U8316 ( .A1(\mem[472][4] ), .A2(n13530), .B1(n26658), .B2(
        data_in[4]), .ZN(n13534) );
  INV_X1 U8317 ( .A(n13535), .ZN(n22325) );
  AOI22_X1 U8318 ( .A1(\mem[472][5] ), .A2(n13530), .B1(n26658), .B2(
        data_in[5]), .ZN(n13535) );
  INV_X1 U8319 ( .A(n13536), .ZN(n22324) );
  AOI22_X1 U8320 ( .A1(\mem[472][6] ), .A2(n13530), .B1(n26658), .B2(
        data_in[6]), .ZN(n13536) );
  INV_X1 U8321 ( .A(n13537), .ZN(n22323) );
  AOI22_X1 U8322 ( .A1(\mem[472][7] ), .A2(n13530), .B1(n26658), .B2(
        data_in[7]), .ZN(n13537) );
  INV_X1 U8323 ( .A(n13538), .ZN(n22322) );
  AOI22_X1 U8324 ( .A1(\mem[473][0] ), .A2(n13539), .B1(n26657), .B2(
        data_in[0]), .ZN(n13538) );
  INV_X1 U8325 ( .A(n13540), .ZN(n22321) );
  AOI22_X1 U8326 ( .A1(\mem[473][1] ), .A2(n13539), .B1(n26657), .B2(
        data_in[1]), .ZN(n13540) );
  INV_X1 U8327 ( .A(n13541), .ZN(n22320) );
  AOI22_X1 U8328 ( .A1(\mem[473][2] ), .A2(n13539), .B1(n26657), .B2(
        data_in[2]), .ZN(n13541) );
  INV_X1 U8329 ( .A(n13542), .ZN(n22319) );
  AOI22_X1 U8330 ( .A1(\mem[473][3] ), .A2(n13539), .B1(n26657), .B2(
        data_in[3]), .ZN(n13542) );
  INV_X1 U8331 ( .A(n13543), .ZN(n22318) );
  AOI22_X1 U8332 ( .A1(\mem[473][4] ), .A2(n13539), .B1(n26657), .B2(
        data_in[4]), .ZN(n13543) );
  INV_X1 U8333 ( .A(n13544), .ZN(n22317) );
  AOI22_X1 U8334 ( .A1(\mem[473][5] ), .A2(n13539), .B1(n26657), .B2(
        data_in[5]), .ZN(n13544) );
  INV_X1 U8335 ( .A(n13545), .ZN(n22316) );
  AOI22_X1 U8336 ( .A1(\mem[473][6] ), .A2(n13539), .B1(n26657), .B2(
        data_in[6]), .ZN(n13545) );
  INV_X1 U8337 ( .A(n13546), .ZN(n22315) );
  AOI22_X1 U8338 ( .A1(\mem[473][7] ), .A2(n13539), .B1(n26657), .B2(
        data_in[7]), .ZN(n13546) );
  INV_X1 U8339 ( .A(n13547), .ZN(n22314) );
  AOI22_X1 U8340 ( .A1(\mem[474][0] ), .A2(n13548), .B1(n26656), .B2(
        data_in[0]), .ZN(n13547) );
  INV_X1 U8341 ( .A(n13549), .ZN(n22313) );
  AOI22_X1 U8342 ( .A1(\mem[474][1] ), .A2(n13548), .B1(n26656), .B2(
        data_in[1]), .ZN(n13549) );
  INV_X1 U8343 ( .A(n13550), .ZN(n22312) );
  AOI22_X1 U8344 ( .A1(\mem[474][2] ), .A2(n13548), .B1(n26656), .B2(
        data_in[2]), .ZN(n13550) );
  INV_X1 U8345 ( .A(n13551), .ZN(n22311) );
  AOI22_X1 U8346 ( .A1(\mem[474][3] ), .A2(n13548), .B1(n26656), .B2(
        data_in[3]), .ZN(n13551) );
  INV_X1 U8347 ( .A(n13552), .ZN(n22310) );
  AOI22_X1 U8348 ( .A1(\mem[474][4] ), .A2(n13548), .B1(n26656), .B2(
        data_in[4]), .ZN(n13552) );
  INV_X1 U8349 ( .A(n13553), .ZN(n22309) );
  AOI22_X1 U8350 ( .A1(\mem[474][5] ), .A2(n13548), .B1(n26656), .B2(
        data_in[5]), .ZN(n13553) );
  INV_X1 U8351 ( .A(n13554), .ZN(n22308) );
  AOI22_X1 U8352 ( .A1(\mem[474][6] ), .A2(n13548), .B1(n26656), .B2(
        data_in[6]), .ZN(n13554) );
  INV_X1 U8353 ( .A(n13555), .ZN(n22307) );
  AOI22_X1 U8354 ( .A1(\mem[474][7] ), .A2(n13548), .B1(n26656), .B2(
        data_in[7]), .ZN(n13555) );
  INV_X1 U8355 ( .A(n13556), .ZN(n22306) );
  AOI22_X1 U8356 ( .A1(\mem[475][0] ), .A2(n13557), .B1(n26655), .B2(
        data_in[0]), .ZN(n13556) );
  INV_X1 U8357 ( .A(n13558), .ZN(n22305) );
  AOI22_X1 U8358 ( .A1(\mem[475][1] ), .A2(n13557), .B1(n26655), .B2(
        data_in[1]), .ZN(n13558) );
  INV_X1 U8359 ( .A(n13559), .ZN(n22304) );
  AOI22_X1 U8360 ( .A1(\mem[475][2] ), .A2(n13557), .B1(n26655), .B2(
        data_in[2]), .ZN(n13559) );
  INV_X1 U8361 ( .A(n13560), .ZN(n22303) );
  AOI22_X1 U8362 ( .A1(\mem[475][3] ), .A2(n13557), .B1(n26655), .B2(
        data_in[3]), .ZN(n13560) );
  INV_X1 U8363 ( .A(n13561), .ZN(n22302) );
  AOI22_X1 U8364 ( .A1(\mem[475][4] ), .A2(n13557), .B1(n26655), .B2(
        data_in[4]), .ZN(n13561) );
  INV_X1 U8365 ( .A(n13562), .ZN(n22301) );
  AOI22_X1 U8366 ( .A1(\mem[475][5] ), .A2(n13557), .B1(n26655), .B2(
        data_in[5]), .ZN(n13562) );
  INV_X1 U8367 ( .A(n13563), .ZN(n22300) );
  AOI22_X1 U8368 ( .A1(\mem[475][6] ), .A2(n13557), .B1(n26655), .B2(
        data_in[6]), .ZN(n13563) );
  INV_X1 U8369 ( .A(n13564), .ZN(n22299) );
  AOI22_X1 U8370 ( .A1(\mem[475][7] ), .A2(n13557), .B1(n26655), .B2(
        data_in[7]), .ZN(n13564) );
  INV_X1 U8371 ( .A(n13565), .ZN(n22298) );
  AOI22_X1 U8372 ( .A1(\mem[476][0] ), .A2(n13566), .B1(n26654), .B2(
        data_in[0]), .ZN(n13565) );
  INV_X1 U8373 ( .A(n13567), .ZN(n22297) );
  AOI22_X1 U8374 ( .A1(\mem[476][1] ), .A2(n13566), .B1(n26654), .B2(
        data_in[1]), .ZN(n13567) );
  INV_X1 U8375 ( .A(n13568), .ZN(n22296) );
  AOI22_X1 U8376 ( .A1(\mem[476][2] ), .A2(n13566), .B1(n26654), .B2(
        data_in[2]), .ZN(n13568) );
  INV_X1 U8377 ( .A(n13569), .ZN(n22295) );
  AOI22_X1 U8378 ( .A1(\mem[476][3] ), .A2(n13566), .B1(n26654), .B2(
        data_in[3]), .ZN(n13569) );
  INV_X1 U8379 ( .A(n13570), .ZN(n22294) );
  AOI22_X1 U8380 ( .A1(\mem[476][4] ), .A2(n13566), .B1(n26654), .B2(
        data_in[4]), .ZN(n13570) );
  INV_X1 U8381 ( .A(n13571), .ZN(n22293) );
  AOI22_X1 U8382 ( .A1(\mem[476][5] ), .A2(n13566), .B1(n26654), .B2(
        data_in[5]), .ZN(n13571) );
  INV_X1 U8383 ( .A(n13572), .ZN(n22292) );
  AOI22_X1 U8384 ( .A1(\mem[476][6] ), .A2(n13566), .B1(n26654), .B2(
        data_in[6]), .ZN(n13572) );
  INV_X1 U8385 ( .A(n13573), .ZN(n22291) );
  AOI22_X1 U8386 ( .A1(\mem[476][7] ), .A2(n13566), .B1(n26654), .B2(
        data_in[7]), .ZN(n13573) );
  INV_X1 U8387 ( .A(n13574), .ZN(n22290) );
  AOI22_X1 U8388 ( .A1(\mem[477][0] ), .A2(n13575), .B1(n26653), .B2(
        data_in[0]), .ZN(n13574) );
  INV_X1 U8389 ( .A(n13576), .ZN(n22289) );
  AOI22_X1 U8390 ( .A1(\mem[477][1] ), .A2(n13575), .B1(n26653), .B2(
        data_in[1]), .ZN(n13576) );
  INV_X1 U8391 ( .A(n13577), .ZN(n22288) );
  AOI22_X1 U8392 ( .A1(\mem[477][2] ), .A2(n13575), .B1(n26653), .B2(
        data_in[2]), .ZN(n13577) );
  INV_X1 U8393 ( .A(n13578), .ZN(n22287) );
  AOI22_X1 U8394 ( .A1(\mem[477][3] ), .A2(n13575), .B1(n26653), .B2(
        data_in[3]), .ZN(n13578) );
  INV_X1 U8395 ( .A(n13579), .ZN(n22286) );
  AOI22_X1 U8396 ( .A1(\mem[477][4] ), .A2(n13575), .B1(n26653), .B2(
        data_in[4]), .ZN(n13579) );
  INV_X1 U8397 ( .A(n13580), .ZN(n22285) );
  AOI22_X1 U8398 ( .A1(\mem[477][5] ), .A2(n13575), .B1(n26653), .B2(
        data_in[5]), .ZN(n13580) );
  INV_X1 U8399 ( .A(n13581), .ZN(n22284) );
  AOI22_X1 U8400 ( .A1(\mem[477][6] ), .A2(n13575), .B1(n26653), .B2(
        data_in[6]), .ZN(n13581) );
  INV_X1 U8401 ( .A(n13582), .ZN(n22283) );
  AOI22_X1 U8402 ( .A1(\mem[477][7] ), .A2(n13575), .B1(n26653), .B2(
        data_in[7]), .ZN(n13582) );
  INV_X1 U8403 ( .A(n13583), .ZN(n22282) );
  AOI22_X1 U8404 ( .A1(\mem[478][0] ), .A2(n13584), .B1(n26652), .B2(
        data_in[0]), .ZN(n13583) );
  INV_X1 U8405 ( .A(n13585), .ZN(n22281) );
  AOI22_X1 U8406 ( .A1(\mem[478][1] ), .A2(n13584), .B1(n26652), .B2(
        data_in[1]), .ZN(n13585) );
  INV_X1 U8407 ( .A(n13586), .ZN(n22280) );
  AOI22_X1 U8408 ( .A1(\mem[478][2] ), .A2(n13584), .B1(n26652), .B2(
        data_in[2]), .ZN(n13586) );
  INV_X1 U8409 ( .A(n13587), .ZN(n22279) );
  AOI22_X1 U8410 ( .A1(\mem[478][3] ), .A2(n13584), .B1(n26652), .B2(
        data_in[3]), .ZN(n13587) );
  INV_X1 U8411 ( .A(n13588), .ZN(n22278) );
  AOI22_X1 U8412 ( .A1(\mem[478][4] ), .A2(n13584), .B1(n26652), .B2(
        data_in[4]), .ZN(n13588) );
  INV_X1 U8413 ( .A(n13589), .ZN(n22277) );
  AOI22_X1 U8414 ( .A1(\mem[478][5] ), .A2(n13584), .B1(n26652), .B2(
        data_in[5]), .ZN(n13589) );
  INV_X1 U8415 ( .A(n13590), .ZN(n22276) );
  AOI22_X1 U8416 ( .A1(\mem[478][6] ), .A2(n13584), .B1(n26652), .B2(
        data_in[6]), .ZN(n13590) );
  INV_X1 U8417 ( .A(n13591), .ZN(n22275) );
  AOI22_X1 U8418 ( .A1(\mem[478][7] ), .A2(n13584), .B1(n26652), .B2(
        data_in[7]), .ZN(n13591) );
  INV_X1 U8419 ( .A(n13592), .ZN(n22274) );
  AOI22_X1 U8420 ( .A1(\mem[479][0] ), .A2(n13593), .B1(n26651), .B2(
        data_in[0]), .ZN(n13592) );
  INV_X1 U8421 ( .A(n13594), .ZN(n22273) );
  AOI22_X1 U8422 ( .A1(\mem[479][1] ), .A2(n13593), .B1(n26651), .B2(
        data_in[1]), .ZN(n13594) );
  INV_X1 U8423 ( .A(n13595), .ZN(n22272) );
  AOI22_X1 U8424 ( .A1(\mem[479][2] ), .A2(n13593), .B1(n26651), .B2(
        data_in[2]), .ZN(n13595) );
  INV_X1 U8425 ( .A(n13596), .ZN(n22271) );
  AOI22_X1 U8426 ( .A1(\mem[479][3] ), .A2(n13593), .B1(n26651), .B2(
        data_in[3]), .ZN(n13596) );
  INV_X1 U8427 ( .A(n13597), .ZN(n22270) );
  AOI22_X1 U8428 ( .A1(\mem[479][4] ), .A2(n13593), .B1(n26651), .B2(
        data_in[4]), .ZN(n13597) );
  INV_X1 U8429 ( .A(n13598), .ZN(n22269) );
  AOI22_X1 U8430 ( .A1(\mem[479][5] ), .A2(n13593), .B1(n26651), .B2(
        data_in[5]), .ZN(n13598) );
  INV_X1 U8431 ( .A(n13599), .ZN(n22268) );
  AOI22_X1 U8432 ( .A1(\mem[479][6] ), .A2(n13593), .B1(n26651), .B2(
        data_in[6]), .ZN(n13599) );
  INV_X1 U8433 ( .A(n13600), .ZN(n22267) );
  AOI22_X1 U8434 ( .A1(\mem[479][7] ), .A2(n13593), .B1(n26651), .B2(
        data_in[7]), .ZN(n13600) );
  INV_X1 U8435 ( .A(n13674), .ZN(n22202) );
  AOI22_X1 U8436 ( .A1(\mem[488][0] ), .A2(n13675), .B1(n26642), .B2(
        data_in[0]), .ZN(n13674) );
  INV_X1 U8437 ( .A(n13676), .ZN(n22201) );
  AOI22_X1 U8438 ( .A1(\mem[488][1] ), .A2(n13675), .B1(n26642), .B2(
        data_in[1]), .ZN(n13676) );
  INV_X1 U8439 ( .A(n13677), .ZN(n22200) );
  AOI22_X1 U8440 ( .A1(\mem[488][2] ), .A2(n13675), .B1(n26642), .B2(
        data_in[2]), .ZN(n13677) );
  INV_X1 U8441 ( .A(n13678), .ZN(n22199) );
  AOI22_X1 U8442 ( .A1(\mem[488][3] ), .A2(n13675), .B1(n26642), .B2(
        data_in[3]), .ZN(n13678) );
  INV_X1 U8443 ( .A(n13679), .ZN(n22198) );
  AOI22_X1 U8444 ( .A1(\mem[488][4] ), .A2(n13675), .B1(n26642), .B2(
        data_in[4]), .ZN(n13679) );
  INV_X1 U8445 ( .A(n13680), .ZN(n22197) );
  AOI22_X1 U8446 ( .A1(\mem[488][5] ), .A2(n13675), .B1(n26642), .B2(
        data_in[5]), .ZN(n13680) );
  INV_X1 U8447 ( .A(n13681), .ZN(n22196) );
  AOI22_X1 U8448 ( .A1(\mem[488][6] ), .A2(n13675), .B1(n26642), .B2(
        data_in[6]), .ZN(n13681) );
  INV_X1 U8449 ( .A(n13682), .ZN(n22195) );
  AOI22_X1 U8450 ( .A1(\mem[488][7] ), .A2(n13675), .B1(n26642), .B2(
        data_in[7]), .ZN(n13682) );
  INV_X1 U8451 ( .A(n13683), .ZN(n22194) );
  AOI22_X1 U8452 ( .A1(\mem[489][0] ), .A2(n13684), .B1(n26641), .B2(
        data_in[0]), .ZN(n13683) );
  INV_X1 U8453 ( .A(n13685), .ZN(n22193) );
  AOI22_X1 U8454 ( .A1(\mem[489][1] ), .A2(n13684), .B1(n26641), .B2(
        data_in[1]), .ZN(n13685) );
  INV_X1 U8455 ( .A(n13686), .ZN(n22192) );
  AOI22_X1 U8456 ( .A1(\mem[489][2] ), .A2(n13684), .B1(n26641), .B2(
        data_in[2]), .ZN(n13686) );
  INV_X1 U8457 ( .A(n13687), .ZN(n22191) );
  AOI22_X1 U8458 ( .A1(\mem[489][3] ), .A2(n13684), .B1(n26641), .B2(
        data_in[3]), .ZN(n13687) );
  INV_X1 U8459 ( .A(n13688), .ZN(n22190) );
  AOI22_X1 U8460 ( .A1(\mem[489][4] ), .A2(n13684), .B1(n26641), .B2(
        data_in[4]), .ZN(n13688) );
  INV_X1 U8461 ( .A(n13689), .ZN(n22189) );
  AOI22_X1 U8462 ( .A1(\mem[489][5] ), .A2(n13684), .B1(n26641), .B2(
        data_in[5]), .ZN(n13689) );
  INV_X1 U8463 ( .A(n13690), .ZN(n22188) );
  AOI22_X1 U8464 ( .A1(\mem[489][6] ), .A2(n13684), .B1(n26641), .B2(
        data_in[6]), .ZN(n13690) );
  INV_X1 U8465 ( .A(n13691), .ZN(n22187) );
  AOI22_X1 U8466 ( .A1(\mem[489][7] ), .A2(n13684), .B1(n26641), .B2(
        data_in[7]), .ZN(n13691) );
  INV_X1 U8467 ( .A(n13692), .ZN(n22186) );
  AOI22_X1 U8468 ( .A1(\mem[490][0] ), .A2(n13693), .B1(n26640), .B2(
        data_in[0]), .ZN(n13692) );
  INV_X1 U8469 ( .A(n13694), .ZN(n22185) );
  AOI22_X1 U8470 ( .A1(\mem[490][1] ), .A2(n13693), .B1(n26640), .B2(
        data_in[1]), .ZN(n13694) );
  INV_X1 U8471 ( .A(n13695), .ZN(n22184) );
  AOI22_X1 U8472 ( .A1(\mem[490][2] ), .A2(n13693), .B1(n26640), .B2(
        data_in[2]), .ZN(n13695) );
  INV_X1 U8473 ( .A(n13696), .ZN(n22183) );
  AOI22_X1 U8474 ( .A1(\mem[490][3] ), .A2(n13693), .B1(n26640), .B2(
        data_in[3]), .ZN(n13696) );
  INV_X1 U8475 ( .A(n13697), .ZN(n22182) );
  AOI22_X1 U8476 ( .A1(\mem[490][4] ), .A2(n13693), .B1(n26640), .B2(
        data_in[4]), .ZN(n13697) );
  INV_X1 U8477 ( .A(n13698), .ZN(n22181) );
  AOI22_X1 U8478 ( .A1(\mem[490][5] ), .A2(n13693), .B1(n26640), .B2(
        data_in[5]), .ZN(n13698) );
  INV_X1 U8479 ( .A(n13699), .ZN(n22180) );
  AOI22_X1 U8480 ( .A1(\mem[490][6] ), .A2(n13693), .B1(n26640), .B2(
        data_in[6]), .ZN(n13699) );
  INV_X1 U8481 ( .A(n13700), .ZN(n22179) );
  AOI22_X1 U8482 ( .A1(\mem[490][7] ), .A2(n13693), .B1(n26640), .B2(
        data_in[7]), .ZN(n13700) );
  INV_X1 U8483 ( .A(n13701), .ZN(n22178) );
  AOI22_X1 U8484 ( .A1(\mem[491][0] ), .A2(n13702), .B1(n26639), .B2(
        data_in[0]), .ZN(n13701) );
  INV_X1 U8485 ( .A(n13703), .ZN(n22177) );
  AOI22_X1 U8486 ( .A1(\mem[491][1] ), .A2(n13702), .B1(n26639), .B2(
        data_in[1]), .ZN(n13703) );
  INV_X1 U8487 ( .A(n13704), .ZN(n22176) );
  AOI22_X1 U8488 ( .A1(\mem[491][2] ), .A2(n13702), .B1(n26639), .B2(
        data_in[2]), .ZN(n13704) );
  INV_X1 U8489 ( .A(n13705), .ZN(n22175) );
  AOI22_X1 U8490 ( .A1(\mem[491][3] ), .A2(n13702), .B1(n26639), .B2(
        data_in[3]), .ZN(n13705) );
  INV_X1 U8491 ( .A(n13706), .ZN(n22174) );
  AOI22_X1 U8492 ( .A1(\mem[491][4] ), .A2(n13702), .B1(n26639), .B2(
        data_in[4]), .ZN(n13706) );
  INV_X1 U8493 ( .A(n13707), .ZN(n22173) );
  AOI22_X1 U8494 ( .A1(\mem[491][5] ), .A2(n13702), .B1(n26639), .B2(
        data_in[5]), .ZN(n13707) );
  INV_X1 U8495 ( .A(n13708), .ZN(n22172) );
  AOI22_X1 U8496 ( .A1(\mem[491][6] ), .A2(n13702), .B1(n26639), .B2(
        data_in[6]), .ZN(n13708) );
  INV_X1 U8497 ( .A(n13709), .ZN(n22171) );
  AOI22_X1 U8498 ( .A1(\mem[491][7] ), .A2(n13702), .B1(n26639), .B2(
        data_in[7]), .ZN(n13709) );
  INV_X1 U8499 ( .A(n13710), .ZN(n22170) );
  AOI22_X1 U8500 ( .A1(\mem[492][0] ), .A2(n13711), .B1(n26638), .B2(
        data_in[0]), .ZN(n13710) );
  INV_X1 U8501 ( .A(n13712), .ZN(n22169) );
  AOI22_X1 U8502 ( .A1(\mem[492][1] ), .A2(n13711), .B1(n26638), .B2(
        data_in[1]), .ZN(n13712) );
  INV_X1 U8503 ( .A(n13713), .ZN(n22168) );
  AOI22_X1 U8504 ( .A1(\mem[492][2] ), .A2(n13711), .B1(n26638), .B2(
        data_in[2]), .ZN(n13713) );
  INV_X1 U8505 ( .A(n13714), .ZN(n22167) );
  AOI22_X1 U8506 ( .A1(\mem[492][3] ), .A2(n13711), .B1(n26638), .B2(
        data_in[3]), .ZN(n13714) );
  INV_X1 U8507 ( .A(n13715), .ZN(n22166) );
  AOI22_X1 U8508 ( .A1(\mem[492][4] ), .A2(n13711), .B1(n26638), .B2(
        data_in[4]), .ZN(n13715) );
  INV_X1 U8509 ( .A(n13716), .ZN(n22165) );
  AOI22_X1 U8510 ( .A1(\mem[492][5] ), .A2(n13711), .B1(n26638), .B2(
        data_in[5]), .ZN(n13716) );
  INV_X1 U8511 ( .A(n13717), .ZN(n22164) );
  AOI22_X1 U8512 ( .A1(\mem[492][6] ), .A2(n13711), .B1(n26638), .B2(
        data_in[6]), .ZN(n13717) );
  INV_X1 U8513 ( .A(n13718), .ZN(n22163) );
  AOI22_X1 U8514 ( .A1(\mem[492][7] ), .A2(n13711), .B1(n26638), .B2(
        data_in[7]), .ZN(n13718) );
  INV_X1 U8515 ( .A(n13719), .ZN(n22162) );
  AOI22_X1 U8516 ( .A1(\mem[493][0] ), .A2(n13720), .B1(n26637), .B2(
        data_in[0]), .ZN(n13719) );
  INV_X1 U8517 ( .A(n13721), .ZN(n22161) );
  AOI22_X1 U8518 ( .A1(\mem[493][1] ), .A2(n13720), .B1(n26637), .B2(
        data_in[1]), .ZN(n13721) );
  INV_X1 U8519 ( .A(n13722), .ZN(n22160) );
  AOI22_X1 U8520 ( .A1(\mem[493][2] ), .A2(n13720), .B1(n26637), .B2(
        data_in[2]), .ZN(n13722) );
  INV_X1 U8521 ( .A(n13723), .ZN(n22159) );
  AOI22_X1 U8522 ( .A1(\mem[493][3] ), .A2(n13720), .B1(n26637), .B2(
        data_in[3]), .ZN(n13723) );
  INV_X1 U8523 ( .A(n13724), .ZN(n22158) );
  AOI22_X1 U8524 ( .A1(\mem[493][4] ), .A2(n13720), .B1(n26637), .B2(
        data_in[4]), .ZN(n13724) );
  INV_X1 U8525 ( .A(n13725), .ZN(n22157) );
  AOI22_X1 U8526 ( .A1(\mem[493][5] ), .A2(n13720), .B1(n26637), .B2(
        data_in[5]), .ZN(n13725) );
  INV_X1 U8527 ( .A(n13726), .ZN(n22156) );
  AOI22_X1 U8528 ( .A1(\mem[493][6] ), .A2(n13720), .B1(n26637), .B2(
        data_in[6]), .ZN(n13726) );
  INV_X1 U8529 ( .A(n13727), .ZN(n22155) );
  AOI22_X1 U8530 ( .A1(\mem[493][7] ), .A2(n13720), .B1(n26637), .B2(
        data_in[7]), .ZN(n13727) );
  INV_X1 U8531 ( .A(n13728), .ZN(n22154) );
  AOI22_X1 U8532 ( .A1(\mem[494][0] ), .A2(n13729), .B1(n26636), .B2(
        data_in[0]), .ZN(n13728) );
  INV_X1 U8533 ( .A(n13730), .ZN(n22153) );
  AOI22_X1 U8534 ( .A1(\mem[494][1] ), .A2(n13729), .B1(n26636), .B2(
        data_in[1]), .ZN(n13730) );
  INV_X1 U8535 ( .A(n13731), .ZN(n22152) );
  AOI22_X1 U8536 ( .A1(\mem[494][2] ), .A2(n13729), .B1(n26636), .B2(
        data_in[2]), .ZN(n13731) );
  INV_X1 U8537 ( .A(n13732), .ZN(n22151) );
  AOI22_X1 U8538 ( .A1(\mem[494][3] ), .A2(n13729), .B1(n26636), .B2(
        data_in[3]), .ZN(n13732) );
  INV_X1 U8539 ( .A(n13733), .ZN(n22150) );
  AOI22_X1 U8540 ( .A1(\mem[494][4] ), .A2(n13729), .B1(n26636), .B2(
        data_in[4]), .ZN(n13733) );
  INV_X1 U8541 ( .A(n13734), .ZN(n22149) );
  AOI22_X1 U8542 ( .A1(\mem[494][5] ), .A2(n13729), .B1(n26636), .B2(
        data_in[5]), .ZN(n13734) );
  INV_X1 U8543 ( .A(n13735), .ZN(n22148) );
  AOI22_X1 U8544 ( .A1(\mem[494][6] ), .A2(n13729), .B1(n26636), .B2(
        data_in[6]), .ZN(n13735) );
  INV_X1 U8545 ( .A(n13736), .ZN(n22147) );
  AOI22_X1 U8546 ( .A1(\mem[494][7] ), .A2(n13729), .B1(n26636), .B2(
        data_in[7]), .ZN(n13736) );
  INV_X1 U8547 ( .A(n13737), .ZN(n22146) );
  AOI22_X1 U8548 ( .A1(\mem[495][0] ), .A2(n13738), .B1(n26635), .B2(
        data_in[0]), .ZN(n13737) );
  INV_X1 U8549 ( .A(n13739), .ZN(n22145) );
  AOI22_X1 U8550 ( .A1(\mem[495][1] ), .A2(n13738), .B1(n26635), .B2(
        data_in[1]), .ZN(n13739) );
  INV_X1 U8551 ( .A(n13740), .ZN(n22144) );
  AOI22_X1 U8552 ( .A1(\mem[495][2] ), .A2(n13738), .B1(n26635), .B2(
        data_in[2]), .ZN(n13740) );
  INV_X1 U8553 ( .A(n13741), .ZN(n22143) );
  AOI22_X1 U8554 ( .A1(\mem[495][3] ), .A2(n13738), .B1(n26635), .B2(
        data_in[3]), .ZN(n13741) );
  INV_X1 U8555 ( .A(n13742), .ZN(n22142) );
  AOI22_X1 U8556 ( .A1(\mem[495][4] ), .A2(n13738), .B1(n26635), .B2(
        data_in[4]), .ZN(n13742) );
  INV_X1 U8557 ( .A(n13743), .ZN(n22141) );
  AOI22_X1 U8558 ( .A1(\mem[495][5] ), .A2(n13738), .B1(n26635), .B2(
        data_in[5]), .ZN(n13743) );
  INV_X1 U8559 ( .A(n13744), .ZN(n22140) );
  AOI22_X1 U8560 ( .A1(\mem[495][6] ), .A2(n13738), .B1(n26635), .B2(
        data_in[6]), .ZN(n13744) );
  INV_X1 U8561 ( .A(n13745), .ZN(n22139) );
  AOI22_X1 U8562 ( .A1(\mem[495][7] ), .A2(n13738), .B1(n26635), .B2(
        data_in[7]), .ZN(n13745) );
  INV_X1 U8563 ( .A(n13746), .ZN(n22138) );
  AOI22_X1 U8564 ( .A1(\mem[496][0] ), .A2(n13747), .B1(n26634), .B2(
        data_in[0]), .ZN(n13746) );
  INV_X1 U8565 ( .A(n13748), .ZN(n22137) );
  AOI22_X1 U8566 ( .A1(\mem[496][1] ), .A2(n13747), .B1(n26634), .B2(
        data_in[1]), .ZN(n13748) );
  INV_X1 U8567 ( .A(n13749), .ZN(n22136) );
  AOI22_X1 U8568 ( .A1(\mem[496][2] ), .A2(n13747), .B1(n26634), .B2(
        data_in[2]), .ZN(n13749) );
  INV_X1 U8569 ( .A(n13750), .ZN(n22135) );
  AOI22_X1 U8570 ( .A1(\mem[496][3] ), .A2(n13747), .B1(n26634), .B2(
        data_in[3]), .ZN(n13750) );
  INV_X1 U8571 ( .A(n13751), .ZN(n22134) );
  AOI22_X1 U8572 ( .A1(\mem[496][4] ), .A2(n13747), .B1(n26634), .B2(
        data_in[4]), .ZN(n13751) );
  INV_X1 U8573 ( .A(n13752), .ZN(n22133) );
  AOI22_X1 U8574 ( .A1(\mem[496][5] ), .A2(n13747), .B1(n26634), .B2(
        data_in[5]), .ZN(n13752) );
  INV_X1 U8575 ( .A(n13753), .ZN(n22132) );
  AOI22_X1 U8576 ( .A1(\mem[496][6] ), .A2(n13747), .B1(n26634), .B2(
        data_in[6]), .ZN(n13753) );
  INV_X1 U8577 ( .A(n13754), .ZN(n22131) );
  AOI22_X1 U8578 ( .A1(\mem[496][7] ), .A2(n13747), .B1(n26634), .B2(
        data_in[7]), .ZN(n13754) );
  INV_X1 U8579 ( .A(n13755), .ZN(n22130) );
  AOI22_X1 U8580 ( .A1(\mem[497][0] ), .A2(n13756), .B1(n26633), .B2(
        data_in[0]), .ZN(n13755) );
  INV_X1 U8581 ( .A(n13757), .ZN(n22129) );
  AOI22_X1 U8582 ( .A1(\mem[497][1] ), .A2(n13756), .B1(n26633), .B2(
        data_in[1]), .ZN(n13757) );
  INV_X1 U8583 ( .A(n13758), .ZN(n22128) );
  AOI22_X1 U8584 ( .A1(\mem[497][2] ), .A2(n13756), .B1(n26633), .B2(
        data_in[2]), .ZN(n13758) );
  INV_X1 U8585 ( .A(n13759), .ZN(n22127) );
  AOI22_X1 U8586 ( .A1(\mem[497][3] ), .A2(n13756), .B1(n26633), .B2(
        data_in[3]), .ZN(n13759) );
  INV_X1 U8587 ( .A(n13760), .ZN(n22126) );
  AOI22_X1 U8588 ( .A1(\mem[497][4] ), .A2(n13756), .B1(n26633), .B2(
        data_in[4]), .ZN(n13760) );
  INV_X1 U8589 ( .A(n13761), .ZN(n22125) );
  AOI22_X1 U8590 ( .A1(\mem[497][5] ), .A2(n13756), .B1(n26633), .B2(
        data_in[5]), .ZN(n13761) );
  INV_X1 U8591 ( .A(n13762), .ZN(n22124) );
  AOI22_X1 U8592 ( .A1(\mem[497][6] ), .A2(n13756), .B1(n26633), .B2(
        data_in[6]), .ZN(n13762) );
  INV_X1 U8593 ( .A(n13763), .ZN(n22123) );
  AOI22_X1 U8594 ( .A1(\mem[497][7] ), .A2(n13756), .B1(n26633), .B2(
        data_in[7]), .ZN(n13763) );
  INV_X1 U8595 ( .A(n13764), .ZN(n22122) );
  AOI22_X1 U8596 ( .A1(\mem[498][0] ), .A2(n13765), .B1(n26632), .B2(
        data_in[0]), .ZN(n13764) );
  INV_X1 U8597 ( .A(n13766), .ZN(n22121) );
  AOI22_X1 U8598 ( .A1(\mem[498][1] ), .A2(n13765), .B1(n26632), .B2(
        data_in[1]), .ZN(n13766) );
  INV_X1 U8599 ( .A(n13767), .ZN(n22120) );
  AOI22_X1 U8600 ( .A1(\mem[498][2] ), .A2(n13765), .B1(n26632), .B2(
        data_in[2]), .ZN(n13767) );
  INV_X1 U8601 ( .A(n13768), .ZN(n22119) );
  AOI22_X1 U8602 ( .A1(\mem[498][3] ), .A2(n13765), .B1(n26632), .B2(
        data_in[3]), .ZN(n13768) );
  INV_X1 U8603 ( .A(n13769), .ZN(n22118) );
  AOI22_X1 U8604 ( .A1(\mem[498][4] ), .A2(n13765), .B1(n26632), .B2(
        data_in[4]), .ZN(n13769) );
  INV_X1 U8605 ( .A(n13770), .ZN(n22117) );
  AOI22_X1 U8606 ( .A1(\mem[498][5] ), .A2(n13765), .B1(n26632), .B2(
        data_in[5]), .ZN(n13770) );
  INV_X1 U8607 ( .A(n13771), .ZN(n22116) );
  AOI22_X1 U8608 ( .A1(\mem[498][6] ), .A2(n13765), .B1(n26632), .B2(
        data_in[6]), .ZN(n13771) );
  INV_X1 U8609 ( .A(n13772), .ZN(n22115) );
  AOI22_X1 U8610 ( .A1(\mem[498][7] ), .A2(n13765), .B1(n26632), .B2(
        data_in[7]), .ZN(n13772) );
  INV_X1 U8611 ( .A(n13773), .ZN(n22114) );
  AOI22_X1 U8612 ( .A1(\mem[499][0] ), .A2(n13774), .B1(n26631), .B2(
        data_in[0]), .ZN(n13773) );
  INV_X1 U8613 ( .A(n13775), .ZN(n22113) );
  AOI22_X1 U8614 ( .A1(\mem[499][1] ), .A2(n13774), .B1(n26631), .B2(
        data_in[1]), .ZN(n13775) );
  INV_X1 U8615 ( .A(n13776), .ZN(n22112) );
  AOI22_X1 U8616 ( .A1(\mem[499][2] ), .A2(n13774), .B1(n26631), .B2(
        data_in[2]), .ZN(n13776) );
  INV_X1 U8617 ( .A(n13777), .ZN(n22111) );
  AOI22_X1 U8618 ( .A1(\mem[499][3] ), .A2(n13774), .B1(n26631), .B2(
        data_in[3]), .ZN(n13777) );
  INV_X1 U8619 ( .A(n13778), .ZN(n22110) );
  AOI22_X1 U8620 ( .A1(\mem[499][4] ), .A2(n13774), .B1(n26631), .B2(
        data_in[4]), .ZN(n13778) );
  INV_X1 U8621 ( .A(n13779), .ZN(n22109) );
  AOI22_X1 U8622 ( .A1(\mem[499][5] ), .A2(n13774), .B1(n26631), .B2(
        data_in[5]), .ZN(n13779) );
  INV_X1 U8623 ( .A(n13780), .ZN(n22108) );
  AOI22_X1 U8624 ( .A1(\mem[499][6] ), .A2(n13774), .B1(n26631), .B2(
        data_in[6]), .ZN(n13780) );
  INV_X1 U8625 ( .A(n13781), .ZN(n22107) );
  AOI22_X1 U8626 ( .A1(\mem[499][7] ), .A2(n13774), .B1(n26631), .B2(
        data_in[7]), .ZN(n13781) );
  INV_X1 U8627 ( .A(n13782), .ZN(n22106) );
  AOI22_X1 U8628 ( .A1(\mem[500][0] ), .A2(n13783), .B1(n26630), .B2(
        data_in[0]), .ZN(n13782) );
  INV_X1 U8629 ( .A(n13784), .ZN(n22105) );
  AOI22_X1 U8630 ( .A1(\mem[500][1] ), .A2(n13783), .B1(n26630), .B2(
        data_in[1]), .ZN(n13784) );
  INV_X1 U8631 ( .A(n13785), .ZN(n22104) );
  AOI22_X1 U8632 ( .A1(\mem[500][2] ), .A2(n13783), .B1(n26630), .B2(
        data_in[2]), .ZN(n13785) );
  INV_X1 U8633 ( .A(n13786), .ZN(n22103) );
  AOI22_X1 U8634 ( .A1(\mem[500][3] ), .A2(n13783), .B1(n26630), .B2(
        data_in[3]), .ZN(n13786) );
  INV_X1 U8635 ( .A(n13787), .ZN(n22102) );
  AOI22_X1 U8636 ( .A1(\mem[500][4] ), .A2(n13783), .B1(n26630), .B2(
        data_in[4]), .ZN(n13787) );
  INV_X1 U8637 ( .A(n13788), .ZN(n22101) );
  AOI22_X1 U8638 ( .A1(\mem[500][5] ), .A2(n13783), .B1(n26630), .B2(
        data_in[5]), .ZN(n13788) );
  INV_X1 U8639 ( .A(n13789), .ZN(n22100) );
  AOI22_X1 U8640 ( .A1(\mem[500][6] ), .A2(n13783), .B1(n26630), .B2(
        data_in[6]), .ZN(n13789) );
  INV_X1 U8641 ( .A(n13790), .ZN(n22099) );
  AOI22_X1 U8642 ( .A1(\mem[500][7] ), .A2(n13783), .B1(n26630), .B2(
        data_in[7]), .ZN(n13790) );
  INV_X1 U8643 ( .A(n13791), .ZN(n22098) );
  AOI22_X1 U8644 ( .A1(\mem[501][0] ), .A2(n13792), .B1(n26629), .B2(
        data_in[0]), .ZN(n13791) );
  INV_X1 U8645 ( .A(n13793), .ZN(n22097) );
  AOI22_X1 U8646 ( .A1(\mem[501][1] ), .A2(n13792), .B1(n26629), .B2(
        data_in[1]), .ZN(n13793) );
  INV_X1 U8647 ( .A(n13794), .ZN(n22096) );
  AOI22_X1 U8648 ( .A1(\mem[501][2] ), .A2(n13792), .B1(n26629), .B2(
        data_in[2]), .ZN(n13794) );
  INV_X1 U8649 ( .A(n13795), .ZN(n22095) );
  AOI22_X1 U8650 ( .A1(\mem[501][3] ), .A2(n13792), .B1(n26629), .B2(
        data_in[3]), .ZN(n13795) );
  INV_X1 U8651 ( .A(n13796), .ZN(n22094) );
  AOI22_X1 U8652 ( .A1(\mem[501][4] ), .A2(n13792), .B1(n26629), .B2(
        data_in[4]), .ZN(n13796) );
  INV_X1 U8653 ( .A(n13797), .ZN(n22093) );
  AOI22_X1 U8654 ( .A1(\mem[501][5] ), .A2(n13792), .B1(n26629), .B2(
        data_in[5]), .ZN(n13797) );
  INV_X1 U8655 ( .A(n13798), .ZN(n22092) );
  AOI22_X1 U8656 ( .A1(\mem[501][6] ), .A2(n13792), .B1(n26629), .B2(
        data_in[6]), .ZN(n13798) );
  INV_X1 U8657 ( .A(n13799), .ZN(n22091) );
  AOI22_X1 U8658 ( .A1(\mem[501][7] ), .A2(n13792), .B1(n26629), .B2(
        data_in[7]), .ZN(n13799) );
  INV_X1 U8659 ( .A(n13800), .ZN(n22090) );
  AOI22_X1 U8660 ( .A1(\mem[502][0] ), .A2(n13801), .B1(n26628), .B2(
        data_in[0]), .ZN(n13800) );
  INV_X1 U8661 ( .A(n13802), .ZN(n22089) );
  AOI22_X1 U8662 ( .A1(\mem[502][1] ), .A2(n13801), .B1(n26628), .B2(
        data_in[1]), .ZN(n13802) );
  INV_X1 U8663 ( .A(n13803), .ZN(n22088) );
  AOI22_X1 U8664 ( .A1(\mem[502][2] ), .A2(n13801), .B1(n26628), .B2(
        data_in[2]), .ZN(n13803) );
  INV_X1 U8665 ( .A(n13804), .ZN(n22087) );
  AOI22_X1 U8666 ( .A1(\mem[502][3] ), .A2(n13801), .B1(n26628), .B2(
        data_in[3]), .ZN(n13804) );
  INV_X1 U8667 ( .A(n13805), .ZN(n22086) );
  AOI22_X1 U8668 ( .A1(\mem[502][4] ), .A2(n13801), .B1(n26628), .B2(
        data_in[4]), .ZN(n13805) );
  INV_X1 U8669 ( .A(n13806), .ZN(n22085) );
  AOI22_X1 U8670 ( .A1(\mem[502][5] ), .A2(n13801), .B1(n26628), .B2(
        data_in[5]), .ZN(n13806) );
  INV_X1 U8671 ( .A(n13807), .ZN(n22084) );
  AOI22_X1 U8672 ( .A1(\mem[502][6] ), .A2(n13801), .B1(n26628), .B2(
        data_in[6]), .ZN(n13807) );
  INV_X1 U8673 ( .A(n13808), .ZN(n22083) );
  AOI22_X1 U8674 ( .A1(\mem[502][7] ), .A2(n13801), .B1(n26628), .B2(
        data_in[7]), .ZN(n13808) );
  INV_X1 U8675 ( .A(n13809), .ZN(n22082) );
  AOI22_X1 U8676 ( .A1(\mem[503][0] ), .A2(n13810), .B1(n26627), .B2(
        data_in[0]), .ZN(n13809) );
  INV_X1 U8677 ( .A(n13811), .ZN(n22081) );
  AOI22_X1 U8678 ( .A1(\mem[503][1] ), .A2(n13810), .B1(n26627), .B2(
        data_in[1]), .ZN(n13811) );
  INV_X1 U8679 ( .A(n13812), .ZN(n22080) );
  AOI22_X1 U8680 ( .A1(\mem[503][2] ), .A2(n13810), .B1(n26627), .B2(
        data_in[2]), .ZN(n13812) );
  INV_X1 U8681 ( .A(n13813), .ZN(n22079) );
  AOI22_X1 U8682 ( .A1(\mem[503][3] ), .A2(n13810), .B1(n26627), .B2(
        data_in[3]), .ZN(n13813) );
  INV_X1 U8683 ( .A(n13814), .ZN(n22078) );
  AOI22_X1 U8684 ( .A1(\mem[503][4] ), .A2(n13810), .B1(n26627), .B2(
        data_in[4]), .ZN(n13814) );
  INV_X1 U8685 ( .A(n13815), .ZN(n22077) );
  AOI22_X1 U8686 ( .A1(\mem[503][5] ), .A2(n13810), .B1(n26627), .B2(
        data_in[5]), .ZN(n13815) );
  INV_X1 U8687 ( .A(n13816), .ZN(n22076) );
  AOI22_X1 U8688 ( .A1(\mem[503][6] ), .A2(n13810), .B1(n26627), .B2(
        data_in[6]), .ZN(n13816) );
  INV_X1 U8689 ( .A(n13817), .ZN(n22075) );
  AOI22_X1 U8690 ( .A1(\mem[503][7] ), .A2(n13810), .B1(n26627), .B2(
        data_in[7]), .ZN(n13817) );
  INV_X1 U8691 ( .A(n13818), .ZN(n22074) );
  AOI22_X1 U8692 ( .A1(\mem[504][0] ), .A2(n13819), .B1(n26626), .B2(
        data_in[0]), .ZN(n13818) );
  INV_X1 U8693 ( .A(n13820), .ZN(n22073) );
  AOI22_X1 U8694 ( .A1(\mem[504][1] ), .A2(n13819), .B1(n26626), .B2(
        data_in[1]), .ZN(n13820) );
  INV_X1 U8695 ( .A(n13821), .ZN(n22072) );
  AOI22_X1 U8696 ( .A1(\mem[504][2] ), .A2(n13819), .B1(n26626), .B2(
        data_in[2]), .ZN(n13821) );
  INV_X1 U8697 ( .A(n13822), .ZN(n22071) );
  AOI22_X1 U8698 ( .A1(\mem[504][3] ), .A2(n13819), .B1(n26626), .B2(
        data_in[3]), .ZN(n13822) );
  INV_X1 U8699 ( .A(n13823), .ZN(n22070) );
  AOI22_X1 U8700 ( .A1(\mem[504][4] ), .A2(n13819), .B1(n26626), .B2(
        data_in[4]), .ZN(n13823) );
  INV_X1 U8701 ( .A(n13824), .ZN(n22069) );
  AOI22_X1 U8702 ( .A1(\mem[504][5] ), .A2(n13819), .B1(n26626), .B2(
        data_in[5]), .ZN(n13824) );
  INV_X1 U8703 ( .A(n13825), .ZN(n22068) );
  AOI22_X1 U8704 ( .A1(\mem[504][6] ), .A2(n13819), .B1(n26626), .B2(
        data_in[6]), .ZN(n13825) );
  INV_X1 U8705 ( .A(n13826), .ZN(n22067) );
  AOI22_X1 U8706 ( .A1(\mem[504][7] ), .A2(n13819), .B1(n26626), .B2(
        data_in[7]), .ZN(n13826) );
  INV_X1 U8707 ( .A(n13827), .ZN(n22066) );
  AOI22_X1 U8708 ( .A1(\mem[505][0] ), .A2(n13828), .B1(n26625), .B2(
        data_in[0]), .ZN(n13827) );
  INV_X1 U8709 ( .A(n13829), .ZN(n22065) );
  AOI22_X1 U8710 ( .A1(\mem[505][1] ), .A2(n13828), .B1(n26625), .B2(
        data_in[1]), .ZN(n13829) );
  INV_X1 U8711 ( .A(n13830), .ZN(n22064) );
  AOI22_X1 U8712 ( .A1(\mem[505][2] ), .A2(n13828), .B1(n26625), .B2(
        data_in[2]), .ZN(n13830) );
  INV_X1 U8713 ( .A(n13831), .ZN(n22063) );
  AOI22_X1 U8714 ( .A1(\mem[505][3] ), .A2(n13828), .B1(n26625), .B2(
        data_in[3]), .ZN(n13831) );
  INV_X1 U8715 ( .A(n13832), .ZN(n22062) );
  AOI22_X1 U8716 ( .A1(\mem[505][4] ), .A2(n13828), .B1(n26625), .B2(
        data_in[4]), .ZN(n13832) );
  INV_X1 U8717 ( .A(n13833), .ZN(n22061) );
  AOI22_X1 U8718 ( .A1(\mem[505][5] ), .A2(n13828), .B1(n26625), .B2(
        data_in[5]), .ZN(n13833) );
  INV_X1 U8719 ( .A(n13834), .ZN(n22060) );
  AOI22_X1 U8720 ( .A1(\mem[505][6] ), .A2(n13828), .B1(n26625), .B2(
        data_in[6]), .ZN(n13834) );
  INV_X1 U8721 ( .A(n13835), .ZN(n22059) );
  AOI22_X1 U8722 ( .A1(\mem[505][7] ), .A2(n13828), .B1(n26625), .B2(
        data_in[7]), .ZN(n13835) );
  INV_X1 U8723 ( .A(n13836), .ZN(n22058) );
  AOI22_X1 U8724 ( .A1(\mem[506][0] ), .A2(n13837), .B1(n26624), .B2(
        data_in[0]), .ZN(n13836) );
  INV_X1 U8725 ( .A(n13838), .ZN(n22057) );
  AOI22_X1 U8726 ( .A1(\mem[506][1] ), .A2(n13837), .B1(n26624), .B2(
        data_in[1]), .ZN(n13838) );
  INV_X1 U8727 ( .A(n13839), .ZN(n22056) );
  AOI22_X1 U8728 ( .A1(\mem[506][2] ), .A2(n13837), .B1(n26624), .B2(
        data_in[2]), .ZN(n13839) );
  INV_X1 U8729 ( .A(n13840), .ZN(n22055) );
  AOI22_X1 U8730 ( .A1(\mem[506][3] ), .A2(n13837), .B1(n26624), .B2(
        data_in[3]), .ZN(n13840) );
  INV_X1 U8731 ( .A(n13841), .ZN(n22054) );
  AOI22_X1 U8732 ( .A1(\mem[506][4] ), .A2(n13837), .B1(n26624), .B2(
        data_in[4]), .ZN(n13841) );
  INV_X1 U8733 ( .A(n13842), .ZN(n22053) );
  AOI22_X1 U8734 ( .A1(\mem[506][5] ), .A2(n13837), .B1(n26624), .B2(
        data_in[5]), .ZN(n13842) );
  INV_X1 U8735 ( .A(n13843), .ZN(n22052) );
  AOI22_X1 U8736 ( .A1(\mem[506][6] ), .A2(n13837), .B1(n26624), .B2(
        data_in[6]), .ZN(n13843) );
  INV_X1 U8737 ( .A(n13844), .ZN(n22051) );
  AOI22_X1 U8738 ( .A1(\mem[506][7] ), .A2(n13837), .B1(n26624), .B2(
        data_in[7]), .ZN(n13844) );
  INV_X1 U8739 ( .A(n13845), .ZN(n22050) );
  AOI22_X1 U8740 ( .A1(\mem[507][0] ), .A2(n13846), .B1(n26623), .B2(
        data_in[0]), .ZN(n13845) );
  INV_X1 U8741 ( .A(n13847), .ZN(n22049) );
  AOI22_X1 U8742 ( .A1(\mem[507][1] ), .A2(n13846), .B1(n26623), .B2(
        data_in[1]), .ZN(n13847) );
  INV_X1 U8743 ( .A(n13848), .ZN(n22048) );
  AOI22_X1 U8744 ( .A1(\mem[507][2] ), .A2(n13846), .B1(n26623), .B2(
        data_in[2]), .ZN(n13848) );
  INV_X1 U8745 ( .A(n13849), .ZN(n22047) );
  AOI22_X1 U8746 ( .A1(\mem[507][3] ), .A2(n13846), .B1(n26623), .B2(
        data_in[3]), .ZN(n13849) );
  INV_X1 U8747 ( .A(n13850), .ZN(n22046) );
  AOI22_X1 U8748 ( .A1(\mem[507][4] ), .A2(n13846), .B1(n26623), .B2(
        data_in[4]), .ZN(n13850) );
  INV_X1 U8749 ( .A(n13851), .ZN(n22045) );
  AOI22_X1 U8750 ( .A1(\mem[507][5] ), .A2(n13846), .B1(n26623), .B2(
        data_in[5]), .ZN(n13851) );
  INV_X1 U8751 ( .A(n13852), .ZN(n22044) );
  AOI22_X1 U8752 ( .A1(\mem[507][6] ), .A2(n13846), .B1(n26623), .B2(
        data_in[6]), .ZN(n13852) );
  INV_X1 U8753 ( .A(n13853), .ZN(n22043) );
  AOI22_X1 U8754 ( .A1(\mem[507][7] ), .A2(n13846), .B1(n26623), .B2(
        data_in[7]), .ZN(n13853) );
  INV_X1 U8755 ( .A(n13854), .ZN(n22042) );
  AOI22_X1 U8756 ( .A1(\mem[508][0] ), .A2(n13855), .B1(n26622), .B2(
        data_in[0]), .ZN(n13854) );
  INV_X1 U8757 ( .A(n13856), .ZN(n22041) );
  AOI22_X1 U8758 ( .A1(\mem[508][1] ), .A2(n13855), .B1(n26622), .B2(
        data_in[1]), .ZN(n13856) );
  INV_X1 U8759 ( .A(n13857), .ZN(n22040) );
  AOI22_X1 U8760 ( .A1(\mem[508][2] ), .A2(n13855), .B1(n26622), .B2(
        data_in[2]), .ZN(n13857) );
  INV_X1 U8761 ( .A(n13858), .ZN(n22039) );
  AOI22_X1 U8762 ( .A1(\mem[508][3] ), .A2(n13855), .B1(n26622), .B2(
        data_in[3]), .ZN(n13858) );
  INV_X1 U8763 ( .A(n13859), .ZN(n22038) );
  AOI22_X1 U8764 ( .A1(\mem[508][4] ), .A2(n13855), .B1(n26622), .B2(
        data_in[4]), .ZN(n13859) );
  INV_X1 U8765 ( .A(n13860), .ZN(n22037) );
  AOI22_X1 U8766 ( .A1(\mem[508][5] ), .A2(n13855), .B1(n26622), .B2(
        data_in[5]), .ZN(n13860) );
  INV_X1 U8767 ( .A(n13861), .ZN(n22036) );
  AOI22_X1 U8768 ( .A1(\mem[508][6] ), .A2(n13855), .B1(n26622), .B2(
        data_in[6]), .ZN(n13861) );
  INV_X1 U8769 ( .A(n13862), .ZN(n22035) );
  AOI22_X1 U8770 ( .A1(\mem[508][7] ), .A2(n13855), .B1(n26622), .B2(
        data_in[7]), .ZN(n13862) );
  INV_X1 U8771 ( .A(n13863), .ZN(n22034) );
  AOI22_X1 U8772 ( .A1(\mem[509][0] ), .A2(n13864), .B1(n26621), .B2(
        data_in[0]), .ZN(n13863) );
  INV_X1 U8773 ( .A(n13865), .ZN(n22033) );
  AOI22_X1 U8774 ( .A1(\mem[509][1] ), .A2(n13864), .B1(n26621), .B2(
        data_in[1]), .ZN(n13865) );
  INV_X1 U8775 ( .A(n13866), .ZN(n22032) );
  AOI22_X1 U8776 ( .A1(\mem[509][2] ), .A2(n13864), .B1(n26621), .B2(
        data_in[2]), .ZN(n13866) );
  INV_X1 U8777 ( .A(n13867), .ZN(n22031) );
  AOI22_X1 U8778 ( .A1(\mem[509][3] ), .A2(n13864), .B1(n26621), .B2(
        data_in[3]), .ZN(n13867) );
  INV_X1 U8779 ( .A(n13868), .ZN(n22030) );
  AOI22_X1 U8780 ( .A1(\mem[509][4] ), .A2(n13864), .B1(n26621), .B2(
        data_in[4]), .ZN(n13868) );
  INV_X1 U8781 ( .A(n13869), .ZN(n22029) );
  AOI22_X1 U8782 ( .A1(\mem[509][5] ), .A2(n13864), .B1(n26621), .B2(
        data_in[5]), .ZN(n13869) );
  INV_X1 U8783 ( .A(n13870), .ZN(n22028) );
  AOI22_X1 U8784 ( .A1(\mem[509][6] ), .A2(n13864), .B1(n26621), .B2(
        data_in[6]), .ZN(n13870) );
  INV_X1 U8785 ( .A(n13871), .ZN(n22027) );
  AOI22_X1 U8786 ( .A1(\mem[509][7] ), .A2(n13864), .B1(n26621), .B2(
        data_in[7]), .ZN(n13871) );
  INV_X1 U8787 ( .A(n13872), .ZN(n22026) );
  AOI22_X1 U8788 ( .A1(\mem[510][0] ), .A2(n13873), .B1(n26620), .B2(
        data_in[0]), .ZN(n13872) );
  INV_X1 U8789 ( .A(n13874), .ZN(n22025) );
  AOI22_X1 U8790 ( .A1(\mem[510][1] ), .A2(n13873), .B1(n26620), .B2(
        data_in[1]), .ZN(n13874) );
  INV_X1 U8791 ( .A(n13875), .ZN(n22024) );
  AOI22_X1 U8792 ( .A1(\mem[510][2] ), .A2(n13873), .B1(n26620), .B2(
        data_in[2]), .ZN(n13875) );
  INV_X1 U8793 ( .A(n13876), .ZN(n22023) );
  AOI22_X1 U8794 ( .A1(\mem[510][3] ), .A2(n13873), .B1(n26620), .B2(
        data_in[3]), .ZN(n13876) );
  INV_X1 U8795 ( .A(n13877), .ZN(n22022) );
  AOI22_X1 U8796 ( .A1(\mem[510][4] ), .A2(n13873), .B1(n26620), .B2(
        data_in[4]), .ZN(n13877) );
  INV_X1 U8797 ( .A(n13878), .ZN(n22021) );
  AOI22_X1 U8798 ( .A1(\mem[510][5] ), .A2(n13873), .B1(n26620), .B2(
        data_in[5]), .ZN(n13878) );
  INV_X1 U8799 ( .A(n13879), .ZN(n22020) );
  AOI22_X1 U8800 ( .A1(\mem[510][6] ), .A2(n13873), .B1(n26620), .B2(
        data_in[6]), .ZN(n13879) );
  INV_X1 U8801 ( .A(n13880), .ZN(n22019) );
  AOI22_X1 U8802 ( .A1(\mem[510][7] ), .A2(n13873), .B1(n26620), .B2(
        data_in[7]), .ZN(n13880) );
  INV_X1 U8803 ( .A(n13881), .ZN(n22018) );
  AOI22_X1 U8804 ( .A1(\mem[511][0] ), .A2(n13882), .B1(n26619), .B2(
        data_in[0]), .ZN(n13881) );
  INV_X1 U8805 ( .A(n13883), .ZN(n22017) );
  AOI22_X1 U8806 ( .A1(\mem[511][1] ), .A2(n13882), .B1(n26619), .B2(
        data_in[1]), .ZN(n13883) );
  INV_X1 U8807 ( .A(n13884), .ZN(n22016) );
  AOI22_X1 U8808 ( .A1(\mem[511][2] ), .A2(n13882), .B1(n26619), .B2(
        data_in[2]), .ZN(n13884) );
  INV_X1 U8809 ( .A(n13885), .ZN(n22015) );
  AOI22_X1 U8810 ( .A1(\mem[511][3] ), .A2(n13882), .B1(n26619), .B2(
        data_in[3]), .ZN(n13885) );
  INV_X1 U8811 ( .A(n13886), .ZN(n22014) );
  AOI22_X1 U8812 ( .A1(\mem[511][4] ), .A2(n13882), .B1(n26619), .B2(
        data_in[4]), .ZN(n13886) );
  INV_X1 U8813 ( .A(n13887), .ZN(n22013) );
  AOI22_X1 U8814 ( .A1(\mem[511][5] ), .A2(n13882), .B1(n26619), .B2(
        data_in[5]), .ZN(n13887) );
  INV_X1 U8815 ( .A(n13888), .ZN(n22012) );
  AOI22_X1 U8816 ( .A1(\mem[511][6] ), .A2(n13882), .B1(n26619), .B2(
        data_in[6]), .ZN(n13888) );
  INV_X1 U8817 ( .A(n13889), .ZN(n22011) );
  AOI22_X1 U8818 ( .A1(\mem[511][7] ), .A2(n13882), .B1(n26619), .B2(
        data_in[7]), .ZN(n13889) );
  INV_X1 U8819 ( .A(n13963), .ZN(n21946) );
  AOI22_X1 U8820 ( .A1(\mem[520][0] ), .A2(n13964), .B1(n26610), .B2(
        data_in[0]), .ZN(n13963) );
  INV_X1 U8821 ( .A(n13965), .ZN(n21945) );
  AOI22_X1 U8822 ( .A1(\mem[520][1] ), .A2(n13964), .B1(n26610), .B2(
        data_in[1]), .ZN(n13965) );
  INV_X1 U8823 ( .A(n13966), .ZN(n21944) );
  AOI22_X1 U8824 ( .A1(\mem[520][2] ), .A2(n13964), .B1(n26610), .B2(
        data_in[2]), .ZN(n13966) );
  INV_X1 U8825 ( .A(n13967), .ZN(n21943) );
  AOI22_X1 U8826 ( .A1(\mem[520][3] ), .A2(n13964), .B1(n26610), .B2(
        data_in[3]), .ZN(n13967) );
  INV_X1 U8827 ( .A(n13968), .ZN(n21942) );
  AOI22_X1 U8828 ( .A1(\mem[520][4] ), .A2(n13964), .B1(n26610), .B2(
        data_in[4]), .ZN(n13968) );
  INV_X1 U8829 ( .A(n13969), .ZN(n21941) );
  AOI22_X1 U8830 ( .A1(\mem[520][5] ), .A2(n13964), .B1(n26610), .B2(
        data_in[5]), .ZN(n13969) );
  INV_X1 U8831 ( .A(n13970), .ZN(n21940) );
  AOI22_X1 U8832 ( .A1(\mem[520][6] ), .A2(n13964), .B1(n26610), .B2(
        data_in[6]), .ZN(n13970) );
  INV_X1 U8833 ( .A(n13971), .ZN(n21939) );
  AOI22_X1 U8834 ( .A1(\mem[520][7] ), .A2(n13964), .B1(n26610), .B2(
        data_in[7]), .ZN(n13971) );
  INV_X1 U8835 ( .A(n13972), .ZN(n21938) );
  AOI22_X1 U8836 ( .A1(\mem[521][0] ), .A2(n13973), .B1(n26609), .B2(
        data_in[0]), .ZN(n13972) );
  INV_X1 U8837 ( .A(n13974), .ZN(n21937) );
  AOI22_X1 U8838 ( .A1(\mem[521][1] ), .A2(n13973), .B1(n26609), .B2(
        data_in[1]), .ZN(n13974) );
  INV_X1 U8839 ( .A(n13975), .ZN(n21936) );
  AOI22_X1 U8840 ( .A1(\mem[521][2] ), .A2(n13973), .B1(n26609), .B2(
        data_in[2]), .ZN(n13975) );
  INV_X1 U8841 ( .A(n13976), .ZN(n21935) );
  AOI22_X1 U8842 ( .A1(\mem[521][3] ), .A2(n13973), .B1(n26609), .B2(
        data_in[3]), .ZN(n13976) );
  INV_X1 U8843 ( .A(n13977), .ZN(n21934) );
  AOI22_X1 U8844 ( .A1(\mem[521][4] ), .A2(n13973), .B1(n26609), .B2(
        data_in[4]), .ZN(n13977) );
  INV_X1 U8845 ( .A(n13978), .ZN(n21933) );
  AOI22_X1 U8846 ( .A1(\mem[521][5] ), .A2(n13973), .B1(n26609), .B2(
        data_in[5]), .ZN(n13978) );
  INV_X1 U8847 ( .A(n13979), .ZN(n21932) );
  AOI22_X1 U8848 ( .A1(\mem[521][6] ), .A2(n13973), .B1(n26609), .B2(
        data_in[6]), .ZN(n13979) );
  INV_X1 U8849 ( .A(n13980), .ZN(n21931) );
  AOI22_X1 U8850 ( .A1(\mem[521][7] ), .A2(n13973), .B1(n26609), .B2(
        data_in[7]), .ZN(n13980) );
  INV_X1 U8851 ( .A(n13981), .ZN(n21930) );
  AOI22_X1 U8852 ( .A1(\mem[522][0] ), .A2(n13982), .B1(n26608), .B2(
        data_in[0]), .ZN(n13981) );
  INV_X1 U8853 ( .A(n13983), .ZN(n21929) );
  AOI22_X1 U8854 ( .A1(\mem[522][1] ), .A2(n13982), .B1(n26608), .B2(
        data_in[1]), .ZN(n13983) );
  INV_X1 U8855 ( .A(n13984), .ZN(n21928) );
  AOI22_X1 U8856 ( .A1(\mem[522][2] ), .A2(n13982), .B1(n26608), .B2(
        data_in[2]), .ZN(n13984) );
  INV_X1 U8857 ( .A(n13985), .ZN(n21927) );
  AOI22_X1 U8858 ( .A1(\mem[522][3] ), .A2(n13982), .B1(n26608), .B2(
        data_in[3]), .ZN(n13985) );
  INV_X1 U8859 ( .A(n13986), .ZN(n21926) );
  AOI22_X1 U8860 ( .A1(\mem[522][4] ), .A2(n13982), .B1(n26608), .B2(
        data_in[4]), .ZN(n13986) );
  INV_X1 U8861 ( .A(n13987), .ZN(n21925) );
  AOI22_X1 U8862 ( .A1(\mem[522][5] ), .A2(n13982), .B1(n26608), .B2(
        data_in[5]), .ZN(n13987) );
  INV_X1 U8863 ( .A(n13988), .ZN(n21924) );
  AOI22_X1 U8864 ( .A1(\mem[522][6] ), .A2(n13982), .B1(n26608), .B2(
        data_in[6]), .ZN(n13988) );
  INV_X1 U8865 ( .A(n13989), .ZN(n21923) );
  AOI22_X1 U8866 ( .A1(\mem[522][7] ), .A2(n13982), .B1(n26608), .B2(
        data_in[7]), .ZN(n13989) );
  INV_X1 U8867 ( .A(n13990), .ZN(n21922) );
  AOI22_X1 U8868 ( .A1(\mem[523][0] ), .A2(n13991), .B1(n26607), .B2(
        data_in[0]), .ZN(n13990) );
  INV_X1 U8869 ( .A(n13992), .ZN(n21921) );
  AOI22_X1 U8870 ( .A1(\mem[523][1] ), .A2(n13991), .B1(n26607), .B2(
        data_in[1]), .ZN(n13992) );
  INV_X1 U8871 ( .A(n13993), .ZN(n21920) );
  AOI22_X1 U8872 ( .A1(\mem[523][2] ), .A2(n13991), .B1(n26607), .B2(
        data_in[2]), .ZN(n13993) );
  INV_X1 U8873 ( .A(n13994), .ZN(n21919) );
  AOI22_X1 U8874 ( .A1(\mem[523][3] ), .A2(n13991), .B1(n26607), .B2(
        data_in[3]), .ZN(n13994) );
  INV_X1 U8875 ( .A(n13995), .ZN(n21918) );
  AOI22_X1 U8876 ( .A1(\mem[523][4] ), .A2(n13991), .B1(n26607), .B2(
        data_in[4]), .ZN(n13995) );
  INV_X1 U8877 ( .A(n13996), .ZN(n21917) );
  AOI22_X1 U8878 ( .A1(\mem[523][5] ), .A2(n13991), .B1(n26607), .B2(
        data_in[5]), .ZN(n13996) );
  INV_X1 U8879 ( .A(n13997), .ZN(n21916) );
  AOI22_X1 U8880 ( .A1(\mem[523][6] ), .A2(n13991), .B1(n26607), .B2(
        data_in[6]), .ZN(n13997) );
  INV_X1 U8881 ( .A(n13998), .ZN(n21915) );
  AOI22_X1 U8882 ( .A1(\mem[523][7] ), .A2(n13991), .B1(n26607), .B2(
        data_in[7]), .ZN(n13998) );
  INV_X1 U8883 ( .A(n13999), .ZN(n21914) );
  AOI22_X1 U8884 ( .A1(\mem[524][0] ), .A2(n14000), .B1(n26606), .B2(
        data_in[0]), .ZN(n13999) );
  INV_X1 U8885 ( .A(n14001), .ZN(n21913) );
  AOI22_X1 U8886 ( .A1(\mem[524][1] ), .A2(n14000), .B1(n26606), .B2(
        data_in[1]), .ZN(n14001) );
  INV_X1 U8887 ( .A(n14002), .ZN(n21912) );
  AOI22_X1 U8888 ( .A1(\mem[524][2] ), .A2(n14000), .B1(n26606), .B2(
        data_in[2]), .ZN(n14002) );
  INV_X1 U8889 ( .A(n14003), .ZN(n21911) );
  AOI22_X1 U8890 ( .A1(\mem[524][3] ), .A2(n14000), .B1(n26606), .B2(
        data_in[3]), .ZN(n14003) );
  INV_X1 U8891 ( .A(n14004), .ZN(n21910) );
  AOI22_X1 U8892 ( .A1(\mem[524][4] ), .A2(n14000), .B1(n26606), .B2(
        data_in[4]), .ZN(n14004) );
  INV_X1 U8893 ( .A(n14005), .ZN(n21909) );
  AOI22_X1 U8894 ( .A1(\mem[524][5] ), .A2(n14000), .B1(n26606), .B2(
        data_in[5]), .ZN(n14005) );
  INV_X1 U8895 ( .A(n14006), .ZN(n21908) );
  AOI22_X1 U8896 ( .A1(\mem[524][6] ), .A2(n14000), .B1(n26606), .B2(
        data_in[6]), .ZN(n14006) );
  INV_X1 U8897 ( .A(n14007), .ZN(n21907) );
  AOI22_X1 U8898 ( .A1(\mem[524][7] ), .A2(n14000), .B1(n26606), .B2(
        data_in[7]), .ZN(n14007) );
  INV_X1 U8899 ( .A(n14008), .ZN(n21906) );
  AOI22_X1 U8900 ( .A1(\mem[525][0] ), .A2(n14009), .B1(n26605), .B2(
        data_in[0]), .ZN(n14008) );
  INV_X1 U8901 ( .A(n14010), .ZN(n21905) );
  AOI22_X1 U8902 ( .A1(\mem[525][1] ), .A2(n14009), .B1(n26605), .B2(
        data_in[1]), .ZN(n14010) );
  INV_X1 U8903 ( .A(n14011), .ZN(n21904) );
  AOI22_X1 U8904 ( .A1(\mem[525][2] ), .A2(n14009), .B1(n26605), .B2(
        data_in[2]), .ZN(n14011) );
  INV_X1 U8905 ( .A(n14012), .ZN(n21903) );
  AOI22_X1 U8906 ( .A1(\mem[525][3] ), .A2(n14009), .B1(n26605), .B2(
        data_in[3]), .ZN(n14012) );
  INV_X1 U8907 ( .A(n14013), .ZN(n21902) );
  AOI22_X1 U8908 ( .A1(\mem[525][4] ), .A2(n14009), .B1(n26605), .B2(
        data_in[4]), .ZN(n14013) );
  INV_X1 U8909 ( .A(n14014), .ZN(n21901) );
  AOI22_X1 U8910 ( .A1(\mem[525][5] ), .A2(n14009), .B1(n26605), .B2(
        data_in[5]), .ZN(n14014) );
  INV_X1 U8911 ( .A(n14015), .ZN(n21900) );
  AOI22_X1 U8912 ( .A1(\mem[525][6] ), .A2(n14009), .B1(n26605), .B2(
        data_in[6]), .ZN(n14015) );
  INV_X1 U8913 ( .A(n14016), .ZN(n21899) );
  AOI22_X1 U8914 ( .A1(\mem[525][7] ), .A2(n14009), .B1(n26605), .B2(
        data_in[7]), .ZN(n14016) );
  INV_X1 U8915 ( .A(n14017), .ZN(n21898) );
  AOI22_X1 U8916 ( .A1(\mem[526][0] ), .A2(n14018), .B1(n26604), .B2(
        data_in[0]), .ZN(n14017) );
  INV_X1 U8917 ( .A(n14019), .ZN(n21897) );
  AOI22_X1 U8918 ( .A1(\mem[526][1] ), .A2(n14018), .B1(n26604), .B2(
        data_in[1]), .ZN(n14019) );
  INV_X1 U8919 ( .A(n14020), .ZN(n21896) );
  AOI22_X1 U8920 ( .A1(\mem[526][2] ), .A2(n14018), .B1(n26604), .B2(
        data_in[2]), .ZN(n14020) );
  INV_X1 U8921 ( .A(n14021), .ZN(n21895) );
  AOI22_X1 U8922 ( .A1(\mem[526][3] ), .A2(n14018), .B1(n26604), .B2(
        data_in[3]), .ZN(n14021) );
  INV_X1 U8923 ( .A(n14022), .ZN(n21894) );
  AOI22_X1 U8924 ( .A1(\mem[526][4] ), .A2(n14018), .B1(n26604), .B2(
        data_in[4]), .ZN(n14022) );
  INV_X1 U8925 ( .A(n14023), .ZN(n21893) );
  AOI22_X1 U8926 ( .A1(\mem[526][5] ), .A2(n14018), .B1(n26604), .B2(
        data_in[5]), .ZN(n14023) );
  INV_X1 U8927 ( .A(n14024), .ZN(n21892) );
  AOI22_X1 U8928 ( .A1(\mem[526][6] ), .A2(n14018), .B1(n26604), .B2(
        data_in[6]), .ZN(n14024) );
  INV_X1 U8929 ( .A(n14025), .ZN(n21891) );
  AOI22_X1 U8930 ( .A1(\mem[526][7] ), .A2(n14018), .B1(n26604), .B2(
        data_in[7]), .ZN(n14025) );
  INV_X1 U8931 ( .A(n14026), .ZN(n21890) );
  AOI22_X1 U8932 ( .A1(\mem[527][0] ), .A2(n14027), .B1(n26603), .B2(
        data_in[0]), .ZN(n14026) );
  INV_X1 U8933 ( .A(n14028), .ZN(n21889) );
  AOI22_X1 U8934 ( .A1(\mem[527][1] ), .A2(n14027), .B1(n26603), .B2(
        data_in[1]), .ZN(n14028) );
  INV_X1 U8935 ( .A(n14029), .ZN(n21888) );
  AOI22_X1 U8936 ( .A1(\mem[527][2] ), .A2(n14027), .B1(n26603), .B2(
        data_in[2]), .ZN(n14029) );
  INV_X1 U8937 ( .A(n14030), .ZN(n21887) );
  AOI22_X1 U8938 ( .A1(\mem[527][3] ), .A2(n14027), .B1(n26603), .B2(
        data_in[3]), .ZN(n14030) );
  INV_X1 U8939 ( .A(n14031), .ZN(n21886) );
  AOI22_X1 U8940 ( .A1(\mem[527][4] ), .A2(n14027), .B1(n26603), .B2(
        data_in[4]), .ZN(n14031) );
  INV_X1 U8941 ( .A(n14032), .ZN(n21885) );
  AOI22_X1 U8942 ( .A1(\mem[527][5] ), .A2(n14027), .B1(n26603), .B2(
        data_in[5]), .ZN(n14032) );
  INV_X1 U8943 ( .A(n14033), .ZN(n21884) );
  AOI22_X1 U8944 ( .A1(\mem[527][6] ), .A2(n14027), .B1(n26603), .B2(
        data_in[6]), .ZN(n14033) );
  INV_X1 U8945 ( .A(n14034), .ZN(n21883) );
  AOI22_X1 U8946 ( .A1(\mem[527][7] ), .A2(n14027), .B1(n26603), .B2(
        data_in[7]), .ZN(n14034) );
  INV_X1 U8947 ( .A(n14035), .ZN(n21882) );
  AOI22_X1 U8948 ( .A1(\mem[528][0] ), .A2(n14036), .B1(n26602), .B2(
        data_in[0]), .ZN(n14035) );
  INV_X1 U8949 ( .A(n14037), .ZN(n21881) );
  AOI22_X1 U8950 ( .A1(\mem[528][1] ), .A2(n14036), .B1(n26602), .B2(
        data_in[1]), .ZN(n14037) );
  INV_X1 U8951 ( .A(n14038), .ZN(n21880) );
  AOI22_X1 U8952 ( .A1(\mem[528][2] ), .A2(n14036), .B1(n26602), .B2(
        data_in[2]), .ZN(n14038) );
  INV_X1 U8953 ( .A(n14039), .ZN(n21879) );
  AOI22_X1 U8954 ( .A1(\mem[528][3] ), .A2(n14036), .B1(n26602), .B2(
        data_in[3]), .ZN(n14039) );
  INV_X1 U8955 ( .A(n14040), .ZN(n21878) );
  AOI22_X1 U8956 ( .A1(\mem[528][4] ), .A2(n14036), .B1(n26602), .B2(
        data_in[4]), .ZN(n14040) );
  INV_X1 U8957 ( .A(n14041), .ZN(n21877) );
  AOI22_X1 U8958 ( .A1(\mem[528][5] ), .A2(n14036), .B1(n26602), .B2(
        data_in[5]), .ZN(n14041) );
  INV_X1 U8959 ( .A(n14042), .ZN(n21876) );
  AOI22_X1 U8960 ( .A1(\mem[528][6] ), .A2(n14036), .B1(n26602), .B2(
        data_in[6]), .ZN(n14042) );
  INV_X1 U8961 ( .A(n14043), .ZN(n21875) );
  AOI22_X1 U8962 ( .A1(\mem[528][7] ), .A2(n14036), .B1(n26602), .B2(
        data_in[7]), .ZN(n14043) );
  INV_X1 U8963 ( .A(n14044), .ZN(n21874) );
  AOI22_X1 U8964 ( .A1(\mem[529][0] ), .A2(n14045), .B1(n26601), .B2(
        data_in[0]), .ZN(n14044) );
  INV_X1 U8965 ( .A(n14046), .ZN(n21873) );
  AOI22_X1 U8966 ( .A1(\mem[529][1] ), .A2(n14045), .B1(n26601), .B2(
        data_in[1]), .ZN(n14046) );
  INV_X1 U8967 ( .A(n14047), .ZN(n21872) );
  AOI22_X1 U8968 ( .A1(\mem[529][2] ), .A2(n14045), .B1(n26601), .B2(
        data_in[2]), .ZN(n14047) );
  INV_X1 U8969 ( .A(n14048), .ZN(n21871) );
  AOI22_X1 U8970 ( .A1(\mem[529][3] ), .A2(n14045), .B1(n26601), .B2(
        data_in[3]), .ZN(n14048) );
  INV_X1 U8971 ( .A(n14049), .ZN(n21870) );
  AOI22_X1 U8972 ( .A1(\mem[529][4] ), .A2(n14045), .B1(n26601), .B2(
        data_in[4]), .ZN(n14049) );
  INV_X1 U8973 ( .A(n14050), .ZN(n21869) );
  AOI22_X1 U8974 ( .A1(\mem[529][5] ), .A2(n14045), .B1(n26601), .B2(
        data_in[5]), .ZN(n14050) );
  INV_X1 U8975 ( .A(n14051), .ZN(n21868) );
  AOI22_X1 U8976 ( .A1(\mem[529][6] ), .A2(n14045), .B1(n26601), .B2(
        data_in[6]), .ZN(n14051) );
  INV_X1 U8977 ( .A(n14052), .ZN(n21867) );
  AOI22_X1 U8978 ( .A1(\mem[529][7] ), .A2(n14045), .B1(n26601), .B2(
        data_in[7]), .ZN(n14052) );
  INV_X1 U8979 ( .A(n14053), .ZN(n21866) );
  AOI22_X1 U8980 ( .A1(\mem[530][0] ), .A2(n14054), .B1(n26600), .B2(
        data_in[0]), .ZN(n14053) );
  INV_X1 U8981 ( .A(n14055), .ZN(n21865) );
  AOI22_X1 U8982 ( .A1(\mem[530][1] ), .A2(n14054), .B1(n26600), .B2(
        data_in[1]), .ZN(n14055) );
  INV_X1 U8983 ( .A(n14056), .ZN(n21864) );
  AOI22_X1 U8984 ( .A1(\mem[530][2] ), .A2(n14054), .B1(n26600), .B2(
        data_in[2]), .ZN(n14056) );
  INV_X1 U8985 ( .A(n14057), .ZN(n21863) );
  AOI22_X1 U8986 ( .A1(\mem[530][3] ), .A2(n14054), .B1(n26600), .B2(
        data_in[3]), .ZN(n14057) );
  INV_X1 U8987 ( .A(n14058), .ZN(n21862) );
  AOI22_X1 U8988 ( .A1(\mem[530][4] ), .A2(n14054), .B1(n26600), .B2(
        data_in[4]), .ZN(n14058) );
  INV_X1 U8989 ( .A(n14059), .ZN(n21861) );
  AOI22_X1 U8990 ( .A1(\mem[530][5] ), .A2(n14054), .B1(n26600), .B2(
        data_in[5]), .ZN(n14059) );
  INV_X1 U8991 ( .A(n14060), .ZN(n21860) );
  AOI22_X1 U8992 ( .A1(\mem[530][6] ), .A2(n14054), .B1(n26600), .B2(
        data_in[6]), .ZN(n14060) );
  INV_X1 U8993 ( .A(n14061), .ZN(n21859) );
  AOI22_X1 U8994 ( .A1(\mem[530][7] ), .A2(n14054), .B1(n26600), .B2(
        data_in[7]), .ZN(n14061) );
  INV_X1 U8995 ( .A(n14062), .ZN(n21858) );
  AOI22_X1 U8996 ( .A1(\mem[531][0] ), .A2(n14063), .B1(n26599), .B2(
        data_in[0]), .ZN(n14062) );
  INV_X1 U8997 ( .A(n14064), .ZN(n21857) );
  AOI22_X1 U8998 ( .A1(\mem[531][1] ), .A2(n14063), .B1(n26599), .B2(
        data_in[1]), .ZN(n14064) );
  INV_X1 U8999 ( .A(n14065), .ZN(n21856) );
  AOI22_X1 U9000 ( .A1(\mem[531][2] ), .A2(n14063), .B1(n26599), .B2(
        data_in[2]), .ZN(n14065) );
  INV_X1 U9001 ( .A(n14066), .ZN(n21855) );
  AOI22_X1 U9002 ( .A1(\mem[531][3] ), .A2(n14063), .B1(n26599), .B2(
        data_in[3]), .ZN(n14066) );
  INV_X1 U9003 ( .A(n14067), .ZN(n21854) );
  AOI22_X1 U9004 ( .A1(\mem[531][4] ), .A2(n14063), .B1(n26599), .B2(
        data_in[4]), .ZN(n14067) );
  INV_X1 U9005 ( .A(n14068), .ZN(n21853) );
  AOI22_X1 U9006 ( .A1(\mem[531][5] ), .A2(n14063), .B1(n26599), .B2(
        data_in[5]), .ZN(n14068) );
  INV_X1 U9007 ( .A(n14069), .ZN(n21852) );
  AOI22_X1 U9008 ( .A1(\mem[531][6] ), .A2(n14063), .B1(n26599), .B2(
        data_in[6]), .ZN(n14069) );
  INV_X1 U9009 ( .A(n14070), .ZN(n21851) );
  AOI22_X1 U9010 ( .A1(\mem[531][7] ), .A2(n14063), .B1(n26599), .B2(
        data_in[7]), .ZN(n14070) );
  INV_X1 U9011 ( .A(n14071), .ZN(n21850) );
  AOI22_X1 U9012 ( .A1(\mem[532][0] ), .A2(n14072), .B1(n26598), .B2(
        data_in[0]), .ZN(n14071) );
  INV_X1 U9013 ( .A(n14073), .ZN(n21849) );
  AOI22_X1 U9014 ( .A1(\mem[532][1] ), .A2(n14072), .B1(n26598), .B2(
        data_in[1]), .ZN(n14073) );
  INV_X1 U9015 ( .A(n14074), .ZN(n21848) );
  AOI22_X1 U9016 ( .A1(\mem[532][2] ), .A2(n14072), .B1(n26598), .B2(
        data_in[2]), .ZN(n14074) );
  INV_X1 U9017 ( .A(n14075), .ZN(n21847) );
  AOI22_X1 U9018 ( .A1(\mem[532][3] ), .A2(n14072), .B1(n26598), .B2(
        data_in[3]), .ZN(n14075) );
  INV_X1 U9019 ( .A(n14076), .ZN(n21846) );
  AOI22_X1 U9020 ( .A1(\mem[532][4] ), .A2(n14072), .B1(n26598), .B2(
        data_in[4]), .ZN(n14076) );
  INV_X1 U9021 ( .A(n14077), .ZN(n21845) );
  AOI22_X1 U9022 ( .A1(\mem[532][5] ), .A2(n14072), .B1(n26598), .B2(
        data_in[5]), .ZN(n14077) );
  INV_X1 U9023 ( .A(n14078), .ZN(n21844) );
  AOI22_X1 U9024 ( .A1(\mem[532][6] ), .A2(n14072), .B1(n26598), .B2(
        data_in[6]), .ZN(n14078) );
  INV_X1 U9025 ( .A(n14079), .ZN(n21843) );
  AOI22_X1 U9026 ( .A1(\mem[532][7] ), .A2(n14072), .B1(n26598), .B2(
        data_in[7]), .ZN(n14079) );
  INV_X1 U9027 ( .A(n14080), .ZN(n21842) );
  AOI22_X1 U9028 ( .A1(\mem[533][0] ), .A2(n14081), .B1(n26597), .B2(
        data_in[0]), .ZN(n14080) );
  INV_X1 U9029 ( .A(n14082), .ZN(n21841) );
  AOI22_X1 U9030 ( .A1(\mem[533][1] ), .A2(n14081), .B1(n26597), .B2(
        data_in[1]), .ZN(n14082) );
  INV_X1 U9031 ( .A(n14083), .ZN(n21840) );
  AOI22_X1 U9032 ( .A1(\mem[533][2] ), .A2(n14081), .B1(n26597), .B2(
        data_in[2]), .ZN(n14083) );
  INV_X1 U9033 ( .A(n14084), .ZN(n21839) );
  AOI22_X1 U9034 ( .A1(\mem[533][3] ), .A2(n14081), .B1(n26597), .B2(
        data_in[3]), .ZN(n14084) );
  INV_X1 U9035 ( .A(n14085), .ZN(n21838) );
  AOI22_X1 U9036 ( .A1(\mem[533][4] ), .A2(n14081), .B1(n26597), .B2(
        data_in[4]), .ZN(n14085) );
  INV_X1 U9037 ( .A(n14086), .ZN(n21837) );
  AOI22_X1 U9038 ( .A1(\mem[533][5] ), .A2(n14081), .B1(n26597), .B2(
        data_in[5]), .ZN(n14086) );
  INV_X1 U9039 ( .A(n14087), .ZN(n21836) );
  AOI22_X1 U9040 ( .A1(\mem[533][6] ), .A2(n14081), .B1(n26597), .B2(
        data_in[6]), .ZN(n14087) );
  INV_X1 U9041 ( .A(n14088), .ZN(n21835) );
  AOI22_X1 U9042 ( .A1(\mem[533][7] ), .A2(n14081), .B1(n26597), .B2(
        data_in[7]), .ZN(n14088) );
  INV_X1 U9043 ( .A(n14089), .ZN(n21834) );
  AOI22_X1 U9044 ( .A1(\mem[534][0] ), .A2(n14090), .B1(n26596), .B2(
        data_in[0]), .ZN(n14089) );
  INV_X1 U9045 ( .A(n14091), .ZN(n21833) );
  AOI22_X1 U9046 ( .A1(\mem[534][1] ), .A2(n14090), .B1(n26596), .B2(
        data_in[1]), .ZN(n14091) );
  INV_X1 U9047 ( .A(n14092), .ZN(n21832) );
  AOI22_X1 U9048 ( .A1(\mem[534][2] ), .A2(n14090), .B1(n26596), .B2(
        data_in[2]), .ZN(n14092) );
  INV_X1 U9049 ( .A(n14093), .ZN(n21831) );
  AOI22_X1 U9050 ( .A1(\mem[534][3] ), .A2(n14090), .B1(n26596), .B2(
        data_in[3]), .ZN(n14093) );
  INV_X1 U9051 ( .A(n14094), .ZN(n21830) );
  AOI22_X1 U9052 ( .A1(\mem[534][4] ), .A2(n14090), .B1(n26596), .B2(
        data_in[4]), .ZN(n14094) );
  INV_X1 U9053 ( .A(n14095), .ZN(n21829) );
  AOI22_X1 U9054 ( .A1(\mem[534][5] ), .A2(n14090), .B1(n26596), .B2(
        data_in[5]), .ZN(n14095) );
  INV_X1 U9055 ( .A(n14096), .ZN(n21828) );
  AOI22_X1 U9056 ( .A1(\mem[534][6] ), .A2(n14090), .B1(n26596), .B2(
        data_in[6]), .ZN(n14096) );
  INV_X1 U9057 ( .A(n14097), .ZN(n21827) );
  AOI22_X1 U9058 ( .A1(\mem[534][7] ), .A2(n14090), .B1(n26596), .B2(
        data_in[7]), .ZN(n14097) );
  INV_X1 U9059 ( .A(n14098), .ZN(n21826) );
  AOI22_X1 U9060 ( .A1(\mem[535][0] ), .A2(n14099), .B1(n26595), .B2(
        data_in[0]), .ZN(n14098) );
  INV_X1 U9061 ( .A(n14100), .ZN(n21825) );
  AOI22_X1 U9062 ( .A1(\mem[535][1] ), .A2(n14099), .B1(n26595), .B2(
        data_in[1]), .ZN(n14100) );
  INV_X1 U9063 ( .A(n14101), .ZN(n21824) );
  AOI22_X1 U9064 ( .A1(\mem[535][2] ), .A2(n14099), .B1(n26595), .B2(
        data_in[2]), .ZN(n14101) );
  INV_X1 U9065 ( .A(n14102), .ZN(n21823) );
  AOI22_X1 U9066 ( .A1(\mem[535][3] ), .A2(n14099), .B1(n26595), .B2(
        data_in[3]), .ZN(n14102) );
  INV_X1 U9067 ( .A(n14103), .ZN(n21822) );
  AOI22_X1 U9068 ( .A1(\mem[535][4] ), .A2(n14099), .B1(n26595), .B2(
        data_in[4]), .ZN(n14103) );
  INV_X1 U9069 ( .A(n14104), .ZN(n21821) );
  AOI22_X1 U9070 ( .A1(\mem[535][5] ), .A2(n14099), .B1(n26595), .B2(
        data_in[5]), .ZN(n14104) );
  INV_X1 U9071 ( .A(n14105), .ZN(n21820) );
  AOI22_X1 U9072 ( .A1(\mem[535][6] ), .A2(n14099), .B1(n26595), .B2(
        data_in[6]), .ZN(n14105) );
  INV_X1 U9073 ( .A(n14106), .ZN(n21819) );
  AOI22_X1 U9074 ( .A1(\mem[535][7] ), .A2(n14099), .B1(n26595), .B2(
        data_in[7]), .ZN(n14106) );
  INV_X1 U9075 ( .A(n14107), .ZN(n21818) );
  AOI22_X1 U9076 ( .A1(\mem[536][0] ), .A2(n14108), .B1(n26594), .B2(
        data_in[0]), .ZN(n14107) );
  INV_X1 U9077 ( .A(n14109), .ZN(n21817) );
  AOI22_X1 U9078 ( .A1(\mem[536][1] ), .A2(n14108), .B1(n26594), .B2(
        data_in[1]), .ZN(n14109) );
  INV_X1 U9079 ( .A(n14110), .ZN(n21816) );
  AOI22_X1 U9080 ( .A1(\mem[536][2] ), .A2(n14108), .B1(n26594), .B2(
        data_in[2]), .ZN(n14110) );
  INV_X1 U9081 ( .A(n14111), .ZN(n21815) );
  AOI22_X1 U9082 ( .A1(\mem[536][3] ), .A2(n14108), .B1(n26594), .B2(
        data_in[3]), .ZN(n14111) );
  INV_X1 U9083 ( .A(n14112), .ZN(n21814) );
  AOI22_X1 U9084 ( .A1(\mem[536][4] ), .A2(n14108), .B1(n26594), .B2(
        data_in[4]), .ZN(n14112) );
  INV_X1 U9085 ( .A(n14113), .ZN(n21813) );
  AOI22_X1 U9086 ( .A1(\mem[536][5] ), .A2(n14108), .B1(n26594), .B2(
        data_in[5]), .ZN(n14113) );
  INV_X1 U9087 ( .A(n14114), .ZN(n21812) );
  AOI22_X1 U9088 ( .A1(\mem[536][6] ), .A2(n14108), .B1(n26594), .B2(
        data_in[6]), .ZN(n14114) );
  INV_X1 U9089 ( .A(n14115), .ZN(n21811) );
  AOI22_X1 U9090 ( .A1(\mem[536][7] ), .A2(n14108), .B1(n26594), .B2(
        data_in[7]), .ZN(n14115) );
  INV_X1 U9091 ( .A(n14116), .ZN(n21810) );
  AOI22_X1 U9092 ( .A1(\mem[537][0] ), .A2(n14117), .B1(n26593), .B2(
        data_in[0]), .ZN(n14116) );
  INV_X1 U9093 ( .A(n14118), .ZN(n21809) );
  AOI22_X1 U9094 ( .A1(\mem[537][1] ), .A2(n14117), .B1(n26593), .B2(
        data_in[1]), .ZN(n14118) );
  INV_X1 U9095 ( .A(n14119), .ZN(n21808) );
  AOI22_X1 U9096 ( .A1(\mem[537][2] ), .A2(n14117), .B1(n26593), .B2(
        data_in[2]), .ZN(n14119) );
  INV_X1 U9097 ( .A(n14120), .ZN(n21807) );
  AOI22_X1 U9098 ( .A1(\mem[537][3] ), .A2(n14117), .B1(n26593), .B2(
        data_in[3]), .ZN(n14120) );
  INV_X1 U9099 ( .A(n14121), .ZN(n21806) );
  AOI22_X1 U9100 ( .A1(\mem[537][4] ), .A2(n14117), .B1(n26593), .B2(
        data_in[4]), .ZN(n14121) );
  INV_X1 U9101 ( .A(n14122), .ZN(n21805) );
  AOI22_X1 U9102 ( .A1(\mem[537][5] ), .A2(n14117), .B1(n26593), .B2(
        data_in[5]), .ZN(n14122) );
  INV_X1 U9103 ( .A(n14123), .ZN(n21804) );
  AOI22_X1 U9104 ( .A1(\mem[537][6] ), .A2(n14117), .B1(n26593), .B2(
        data_in[6]), .ZN(n14123) );
  INV_X1 U9105 ( .A(n14124), .ZN(n21803) );
  AOI22_X1 U9106 ( .A1(\mem[537][7] ), .A2(n14117), .B1(n26593), .B2(
        data_in[7]), .ZN(n14124) );
  INV_X1 U9107 ( .A(n14125), .ZN(n21802) );
  AOI22_X1 U9108 ( .A1(\mem[538][0] ), .A2(n14126), .B1(n26592), .B2(
        data_in[0]), .ZN(n14125) );
  INV_X1 U9109 ( .A(n14127), .ZN(n21801) );
  AOI22_X1 U9110 ( .A1(\mem[538][1] ), .A2(n14126), .B1(n26592), .B2(
        data_in[1]), .ZN(n14127) );
  INV_X1 U9111 ( .A(n14128), .ZN(n21800) );
  AOI22_X1 U9112 ( .A1(\mem[538][2] ), .A2(n14126), .B1(n26592), .B2(
        data_in[2]), .ZN(n14128) );
  INV_X1 U9113 ( .A(n14129), .ZN(n21799) );
  AOI22_X1 U9114 ( .A1(\mem[538][3] ), .A2(n14126), .B1(n26592), .B2(
        data_in[3]), .ZN(n14129) );
  INV_X1 U9115 ( .A(n14130), .ZN(n21798) );
  AOI22_X1 U9116 ( .A1(\mem[538][4] ), .A2(n14126), .B1(n26592), .B2(
        data_in[4]), .ZN(n14130) );
  INV_X1 U9117 ( .A(n14131), .ZN(n21797) );
  AOI22_X1 U9118 ( .A1(\mem[538][5] ), .A2(n14126), .B1(n26592), .B2(
        data_in[5]), .ZN(n14131) );
  INV_X1 U9119 ( .A(n14132), .ZN(n21796) );
  AOI22_X1 U9120 ( .A1(\mem[538][6] ), .A2(n14126), .B1(n26592), .B2(
        data_in[6]), .ZN(n14132) );
  INV_X1 U9121 ( .A(n14133), .ZN(n21795) );
  AOI22_X1 U9122 ( .A1(\mem[538][7] ), .A2(n14126), .B1(n26592), .B2(
        data_in[7]), .ZN(n14133) );
  INV_X1 U9123 ( .A(n14134), .ZN(n21794) );
  AOI22_X1 U9124 ( .A1(\mem[539][0] ), .A2(n14135), .B1(n26591), .B2(
        data_in[0]), .ZN(n14134) );
  INV_X1 U9125 ( .A(n14136), .ZN(n21793) );
  AOI22_X1 U9126 ( .A1(\mem[539][1] ), .A2(n14135), .B1(n26591), .B2(
        data_in[1]), .ZN(n14136) );
  INV_X1 U9127 ( .A(n14137), .ZN(n21792) );
  AOI22_X1 U9128 ( .A1(\mem[539][2] ), .A2(n14135), .B1(n26591), .B2(
        data_in[2]), .ZN(n14137) );
  INV_X1 U9129 ( .A(n14138), .ZN(n21791) );
  AOI22_X1 U9130 ( .A1(\mem[539][3] ), .A2(n14135), .B1(n26591), .B2(
        data_in[3]), .ZN(n14138) );
  INV_X1 U9131 ( .A(n14139), .ZN(n21790) );
  AOI22_X1 U9132 ( .A1(\mem[539][4] ), .A2(n14135), .B1(n26591), .B2(
        data_in[4]), .ZN(n14139) );
  INV_X1 U9133 ( .A(n14140), .ZN(n21789) );
  AOI22_X1 U9134 ( .A1(\mem[539][5] ), .A2(n14135), .B1(n26591), .B2(
        data_in[5]), .ZN(n14140) );
  INV_X1 U9135 ( .A(n14141), .ZN(n21788) );
  AOI22_X1 U9136 ( .A1(\mem[539][6] ), .A2(n14135), .B1(n26591), .B2(
        data_in[6]), .ZN(n14141) );
  INV_X1 U9137 ( .A(n14142), .ZN(n21787) );
  AOI22_X1 U9138 ( .A1(\mem[539][7] ), .A2(n14135), .B1(n26591), .B2(
        data_in[7]), .ZN(n14142) );
  INV_X1 U9139 ( .A(n14143), .ZN(n21786) );
  AOI22_X1 U9140 ( .A1(\mem[540][0] ), .A2(n14144), .B1(n26590), .B2(
        data_in[0]), .ZN(n14143) );
  INV_X1 U9141 ( .A(n14145), .ZN(n21785) );
  AOI22_X1 U9142 ( .A1(\mem[540][1] ), .A2(n14144), .B1(n26590), .B2(
        data_in[1]), .ZN(n14145) );
  INV_X1 U9143 ( .A(n14146), .ZN(n21784) );
  AOI22_X1 U9144 ( .A1(\mem[540][2] ), .A2(n14144), .B1(n26590), .B2(
        data_in[2]), .ZN(n14146) );
  INV_X1 U9145 ( .A(n14147), .ZN(n21783) );
  AOI22_X1 U9146 ( .A1(\mem[540][3] ), .A2(n14144), .B1(n26590), .B2(
        data_in[3]), .ZN(n14147) );
  INV_X1 U9147 ( .A(n14148), .ZN(n21782) );
  AOI22_X1 U9148 ( .A1(\mem[540][4] ), .A2(n14144), .B1(n26590), .B2(
        data_in[4]), .ZN(n14148) );
  INV_X1 U9149 ( .A(n14149), .ZN(n21781) );
  AOI22_X1 U9150 ( .A1(\mem[540][5] ), .A2(n14144), .B1(n26590), .B2(
        data_in[5]), .ZN(n14149) );
  INV_X1 U9151 ( .A(n14150), .ZN(n21780) );
  AOI22_X1 U9152 ( .A1(\mem[540][6] ), .A2(n14144), .B1(n26590), .B2(
        data_in[6]), .ZN(n14150) );
  INV_X1 U9153 ( .A(n14151), .ZN(n21779) );
  AOI22_X1 U9154 ( .A1(\mem[540][7] ), .A2(n14144), .B1(n26590), .B2(
        data_in[7]), .ZN(n14151) );
  INV_X1 U9155 ( .A(n14152), .ZN(n21778) );
  AOI22_X1 U9156 ( .A1(\mem[541][0] ), .A2(n14153), .B1(n26589), .B2(
        data_in[0]), .ZN(n14152) );
  INV_X1 U9157 ( .A(n14154), .ZN(n21777) );
  AOI22_X1 U9158 ( .A1(\mem[541][1] ), .A2(n14153), .B1(n26589), .B2(
        data_in[1]), .ZN(n14154) );
  INV_X1 U9159 ( .A(n14155), .ZN(n21776) );
  AOI22_X1 U9160 ( .A1(\mem[541][2] ), .A2(n14153), .B1(n26589), .B2(
        data_in[2]), .ZN(n14155) );
  INV_X1 U9161 ( .A(n14156), .ZN(n21775) );
  AOI22_X1 U9162 ( .A1(\mem[541][3] ), .A2(n14153), .B1(n26589), .B2(
        data_in[3]), .ZN(n14156) );
  INV_X1 U9163 ( .A(n14157), .ZN(n21774) );
  AOI22_X1 U9164 ( .A1(\mem[541][4] ), .A2(n14153), .B1(n26589), .B2(
        data_in[4]), .ZN(n14157) );
  INV_X1 U9165 ( .A(n14158), .ZN(n21773) );
  AOI22_X1 U9166 ( .A1(\mem[541][5] ), .A2(n14153), .B1(n26589), .B2(
        data_in[5]), .ZN(n14158) );
  INV_X1 U9167 ( .A(n14159), .ZN(n21772) );
  AOI22_X1 U9168 ( .A1(\mem[541][6] ), .A2(n14153), .B1(n26589), .B2(
        data_in[6]), .ZN(n14159) );
  INV_X1 U9169 ( .A(n14160), .ZN(n21771) );
  AOI22_X1 U9170 ( .A1(\mem[541][7] ), .A2(n14153), .B1(n26589), .B2(
        data_in[7]), .ZN(n14160) );
  INV_X1 U9171 ( .A(n14161), .ZN(n21770) );
  AOI22_X1 U9172 ( .A1(\mem[542][0] ), .A2(n14162), .B1(n26588), .B2(
        data_in[0]), .ZN(n14161) );
  INV_X1 U9173 ( .A(n14163), .ZN(n21769) );
  AOI22_X1 U9174 ( .A1(\mem[542][1] ), .A2(n14162), .B1(n26588), .B2(
        data_in[1]), .ZN(n14163) );
  INV_X1 U9175 ( .A(n14164), .ZN(n21768) );
  AOI22_X1 U9176 ( .A1(\mem[542][2] ), .A2(n14162), .B1(n26588), .B2(
        data_in[2]), .ZN(n14164) );
  INV_X1 U9177 ( .A(n14165), .ZN(n21767) );
  AOI22_X1 U9178 ( .A1(\mem[542][3] ), .A2(n14162), .B1(n26588), .B2(
        data_in[3]), .ZN(n14165) );
  INV_X1 U9179 ( .A(n14166), .ZN(n21766) );
  AOI22_X1 U9180 ( .A1(\mem[542][4] ), .A2(n14162), .B1(n26588), .B2(
        data_in[4]), .ZN(n14166) );
  INV_X1 U9181 ( .A(n14167), .ZN(n21765) );
  AOI22_X1 U9182 ( .A1(\mem[542][5] ), .A2(n14162), .B1(n26588), .B2(
        data_in[5]), .ZN(n14167) );
  INV_X1 U9183 ( .A(n14168), .ZN(n21764) );
  AOI22_X1 U9184 ( .A1(\mem[542][6] ), .A2(n14162), .B1(n26588), .B2(
        data_in[6]), .ZN(n14168) );
  INV_X1 U9185 ( .A(n14169), .ZN(n21763) );
  AOI22_X1 U9186 ( .A1(\mem[542][7] ), .A2(n14162), .B1(n26588), .B2(
        data_in[7]), .ZN(n14169) );
  INV_X1 U9187 ( .A(n14170), .ZN(n21762) );
  AOI22_X1 U9188 ( .A1(\mem[543][0] ), .A2(n14171), .B1(n26587), .B2(
        data_in[0]), .ZN(n14170) );
  INV_X1 U9189 ( .A(n14172), .ZN(n21761) );
  AOI22_X1 U9190 ( .A1(\mem[543][1] ), .A2(n14171), .B1(n26587), .B2(
        data_in[1]), .ZN(n14172) );
  INV_X1 U9191 ( .A(n14173), .ZN(n21760) );
  AOI22_X1 U9192 ( .A1(\mem[543][2] ), .A2(n14171), .B1(n26587), .B2(
        data_in[2]), .ZN(n14173) );
  INV_X1 U9193 ( .A(n14174), .ZN(n21759) );
  AOI22_X1 U9194 ( .A1(\mem[543][3] ), .A2(n14171), .B1(n26587), .B2(
        data_in[3]), .ZN(n14174) );
  INV_X1 U9195 ( .A(n14175), .ZN(n21758) );
  AOI22_X1 U9196 ( .A1(\mem[543][4] ), .A2(n14171), .B1(n26587), .B2(
        data_in[4]), .ZN(n14175) );
  INV_X1 U9197 ( .A(n14176), .ZN(n21757) );
  AOI22_X1 U9198 ( .A1(\mem[543][5] ), .A2(n14171), .B1(n26587), .B2(
        data_in[5]), .ZN(n14176) );
  INV_X1 U9199 ( .A(n14177), .ZN(n21756) );
  AOI22_X1 U9200 ( .A1(\mem[543][6] ), .A2(n14171), .B1(n26587), .B2(
        data_in[6]), .ZN(n14177) );
  INV_X1 U9201 ( .A(n14178), .ZN(n21755) );
  AOI22_X1 U9202 ( .A1(\mem[543][7] ), .A2(n14171), .B1(n26587), .B2(
        data_in[7]), .ZN(n14178) );
  INV_X1 U9203 ( .A(n14253), .ZN(n21690) );
  AOI22_X1 U9204 ( .A1(\mem[552][0] ), .A2(n14254), .B1(n26578), .B2(
        data_in[0]), .ZN(n14253) );
  INV_X1 U9205 ( .A(n14255), .ZN(n21689) );
  AOI22_X1 U9206 ( .A1(\mem[552][1] ), .A2(n14254), .B1(n26578), .B2(
        data_in[1]), .ZN(n14255) );
  INV_X1 U9207 ( .A(n14256), .ZN(n21688) );
  AOI22_X1 U9208 ( .A1(\mem[552][2] ), .A2(n14254), .B1(n26578), .B2(
        data_in[2]), .ZN(n14256) );
  INV_X1 U9209 ( .A(n14257), .ZN(n21687) );
  AOI22_X1 U9210 ( .A1(\mem[552][3] ), .A2(n14254), .B1(n26578), .B2(
        data_in[3]), .ZN(n14257) );
  INV_X1 U9211 ( .A(n14258), .ZN(n21686) );
  AOI22_X1 U9212 ( .A1(\mem[552][4] ), .A2(n14254), .B1(n26578), .B2(
        data_in[4]), .ZN(n14258) );
  INV_X1 U9213 ( .A(n14259), .ZN(n21685) );
  AOI22_X1 U9214 ( .A1(\mem[552][5] ), .A2(n14254), .B1(n26578), .B2(
        data_in[5]), .ZN(n14259) );
  INV_X1 U9215 ( .A(n14260), .ZN(n21684) );
  AOI22_X1 U9216 ( .A1(\mem[552][6] ), .A2(n14254), .B1(n26578), .B2(
        data_in[6]), .ZN(n14260) );
  INV_X1 U9217 ( .A(n14261), .ZN(n21683) );
  AOI22_X1 U9218 ( .A1(\mem[552][7] ), .A2(n14254), .B1(n26578), .B2(
        data_in[7]), .ZN(n14261) );
  INV_X1 U9219 ( .A(n14262), .ZN(n21682) );
  AOI22_X1 U9220 ( .A1(\mem[553][0] ), .A2(n14263), .B1(n26577), .B2(
        data_in[0]), .ZN(n14262) );
  INV_X1 U9221 ( .A(n14264), .ZN(n21681) );
  AOI22_X1 U9222 ( .A1(\mem[553][1] ), .A2(n14263), .B1(n26577), .B2(
        data_in[1]), .ZN(n14264) );
  INV_X1 U9223 ( .A(n14265), .ZN(n21680) );
  AOI22_X1 U9224 ( .A1(\mem[553][2] ), .A2(n14263), .B1(n26577), .B2(
        data_in[2]), .ZN(n14265) );
  INV_X1 U9225 ( .A(n14266), .ZN(n21679) );
  AOI22_X1 U9226 ( .A1(\mem[553][3] ), .A2(n14263), .B1(n26577), .B2(
        data_in[3]), .ZN(n14266) );
  INV_X1 U9227 ( .A(n14267), .ZN(n21678) );
  AOI22_X1 U9228 ( .A1(\mem[553][4] ), .A2(n14263), .B1(n26577), .B2(
        data_in[4]), .ZN(n14267) );
  INV_X1 U9229 ( .A(n14268), .ZN(n21677) );
  AOI22_X1 U9230 ( .A1(\mem[553][5] ), .A2(n14263), .B1(n26577), .B2(
        data_in[5]), .ZN(n14268) );
  INV_X1 U9231 ( .A(n14269), .ZN(n21676) );
  AOI22_X1 U9232 ( .A1(\mem[553][6] ), .A2(n14263), .B1(n26577), .B2(
        data_in[6]), .ZN(n14269) );
  INV_X1 U9233 ( .A(n14270), .ZN(n21675) );
  AOI22_X1 U9234 ( .A1(\mem[553][7] ), .A2(n14263), .B1(n26577), .B2(
        data_in[7]), .ZN(n14270) );
  INV_X1 U9235 ( .A(n14271), .ZN(n21674) );
  AOI22_X1 U9236 ( .A1(\mem[554][0] ), .A2(n14272), .B1(n26576), .B2(
        data_in[0]), .ZN(n14271) );
  INV_X1 U9237 ( .A(n14273), .ZN(n21673) );
  AOI22_X1 U9238 ( .A1(\mem[554][1] ), .A2(n14272), .B1(n26576), .B2(
        data_in[1]), .ZN(n14273) );
  INV_X1 U9239 ( .A(n14274), .ZN(n21672) );
  AOI22_X1 U9240 ( .A1(\mem[554][2] ), .A2(n14272), .B1(n26576), .B2(
        data_in[2]), .ZN(n14274) );
  INV_X1 U9241 ( .A(n14275), .ZN(n21671) );
  AOI22_X1 U9242 ( .A1(\mem[554][3] ), .A2(n14272), .B1(n26576), .B2(
        data_in[3]), .ZN(n14275) );
  INV_X1 U9243 ( .A(n14276), .ZN(n21670) );
  AOI22_X1 U9244 ( .A1(\mem[554][4] ), .A2(n14272), .B1(n26576), .B2(
        data_in[4]), .ZN(n14276) );
  INV_X1 U9245 ( .A(n14277), .ZN(n21669) );
  AOI22_X1 U9246 ( .A1(\mem[554][5] ), .A2(n14272), .B1(n26576), .B2(
        data_in[5]), .ZN(n14277) );
  INV_X1 U9247 ( .A(n14278), .ZN(n21668) );
  AOI22_X1 U9248 ( .A1(\mem[554][6] ), .A2(n14272), .B1(n26576), .B2(
        data_in[6]), .ZN(n14278) );
  INV_X1 U9249 ( .A(n14279), .ZN(n21667) );
  AOI22_X1 U9250 ( .A1(\mem[554][7] ), .A2(n14272), .B1(n26576), .B2(
        data_in[7]), .ZN(n14279) );
  INV_X1 U9251 ( .A(n14280), .ZN(n21666) );
  AOI22_X1 U9252 ( .A1(\mem[555][0] ), .A2(n14281), .B1(n26575), .B2(
        data_in[0]), .ZN(n14280) );
  INV_X1 U9253 ( .A(n14282), .ZN(n21665) );
  AOI22_X1 U9254 ( .A1(\mem[555][1] ), .A2(n14281), .B1(n26575), .B2(
        data_in[1]), .ZN(n14282) );
  INV_X1 U9255 ( .A(n14283), .ZN(n21664) );
  AOI22_X1 U9256 ( .A1(\mem[555][2] ), .A2(n14281), .B1(n26575), .B2(
        data_in[2]), .ZN(n14283) );
  INV_X1 U9257 ( .A(n14284), .ZN(n21663) );
  AOI22_X1 U9258 ( .A1(\mem[555][3] ), .A2(n14281), .B1(n26575), .B2(
        data_in[3]), .ZN(n14284) );
  INV_X1 U9259 ( .A(n14285), .ZN(n21662) );
  AOI22_X1 U9260 ( .A1(\mem[555][4] ), .A2(n14281), .B1(n26575), .B2(
        data_in[4]), .ZN(n14285) );
  INV_X1 U9261 ( .A(n14286), .ZN(n21661) );
  AOI22_X1 U9262 ( .A1(\mem[555][5] ), .A2(n14281), .B1(n26575), .B2(
        data_in[5]), .ZN(n14286) );
  INV_X1 U9263 ( .A(n14287), .ZN(n21660) );
  AOI22_X1 U9264 ( .A1(\mem[555][6] ), .A2(n14281), .B1(n26575), .B2(
        data_in[6]), .ZN(n14287) );
  INV_X1 U9265 ( .A(n14288), .ZN(n21659) );
  AOI22_X1 U9266 ( .A1(\mem[555][7] ), .A2(n14281), .B1(n26575), .B2(
        data_in[7]), .ZN(n14288) );
  INV_X1 U9267 ( .A(n14289), .ZN(n21658) );
  AOI22_X1 U9268 ( .A1(\mem[556][0] ), .A2(n14290), .B1(n26574), .B2(
        data_in[0]), .ZN(n14289) );
  INV_X1 U9269 ( .A(n14291), .ZN(n21657) );
  AOI22_X1 U9270 ( .A1(\mem[556][1] ), .A2(n14290), .B1(n26574), .B2(
        data_in[1]), .ZN(n14291) );
  INV_X1 U9271 ( .A(n14292), .ZN(n21656) );
  AOI22_X1 U9272 ( .A1(\mem[556][2] ), .A2(n14290), .B1(n26574), .B2(
        data_in[2]), .ZN(n14292) );
  INV_X1 U9273 ( .A(n14293), .ZN(n21655) );
  AOI22_X1 U9274 ( .A1(\mem[556][3] ), .A2(n14290), .B1(n26574), .B2(
        data_in[3]), .ZN(n14293) );
  INV_X1 U9275 ( .A(n14294), .ZN(n21654) );
  AOI22_X1 U9276 ( .A1(\mem[556][4] ), .A2(n14290), .B1(n26574), .B2(
        data_in[4]), .ZN(n14294) );
  INV_X1 U9277 ( .A(n14295), .ZN(n21653) );
  AOI22_X1 U9278 ( .A1(\mem[556][5] ), .A2(n14290), .B1(n26574), .B2(
        data_in[5]), .ZN(n14295) );
  INV_X1 U9279 ( .A(n14296), .ZN(n21652) );
  AOI22_X1 U9280 ( .A1(\mem[556][6] ), .A2(n14290), .B1(n26574), .B2(
        data_in[6]), .ZN(n14296) );
  INV_X1 U9281 ( .A(n14297), .ZN(n21651) );
  AOI22_X1 U9282 ( .A1(\mem[556][7] ), .A2(n14290), .B1(n26574), .B2(
        data_in[7]), .ZN(n14297) );
  INV_X1 U9283 ( .A(n14298), .ZN(n21650) );
  AOI22_X1 U9284 ( .A1(\mem[557][0] ), .A2(n14299), .B1(n26573), .B2(
        data_in[0]), .ZN(n14298) );
  INV_X1 U9285 ( .A(n14300), .ZN(n21649) );
  AOI22_X1 U9286 ( .A1(\mem[557][1] ), .A2(n14299), .B1(n26573), .B2(
        data_in[1]), .ZN(n14300) );
  INV_X1 U9287 ( .A(n14301), .ZN(n21648) );
  AOI22_X1 U9288 ( .A1(\mem[557][2] ), .A2(n14299), .B1(n26573), .B2(
        data_in[2]), .ZN(n14301) );
  INV_X1 U9289 ( .A(n14302), .ZN(n21647) );
  AOI22_X1 U9290 ( .A1(\mem[557][3] ), .A2(n14299), .B1(n26573), .B2(
        data_in[3]), .ZN(n14302) );
  INV_X1 U9291 ( .A(n14303), .ZN(n21646) );
  AOI22_X1 U9292 ( .A1(\mem[557][4] ), .A2(n14299), .B1(n26573), .B2(
        data_in[4]), .ZN(n14303) );
  INV_X1 U9293 ( .A(n14304), .ZN(n21645) );
  AOI22_X1 U9294 ( .A1(\mem[557][5] ), .A2(n14299), .B1(n26573), .B2(
        data_in[5]), .ZN(n14304) );
  INV_X1 U9295 ( .A(n14305), .ZN(n21644) );
  AOI22_X1 U9296 ( .A1(\mem[557][6] ), .A2(n14299), .B1(n26573), .B2(
        data_in[6]), .ZN(n14305) );
  INV_X1 U9297 ( .A(n14306), .ZN(n21643) );
  AOI22_X1 U9298 ( .A1(\mem[557][7] ), .A2(n14299), .B1(n26573), .B2(
        data_in[7]), .ZN(n14306) );
  INV_X1 U9299 ( .A(n14307), .ZN(n21642) );
  AOI22_X1 U9300 ( .A1(\mem[558][0] ), .A2(n14308), .B1(n26572), .B2(
        data_in[0]), .ZN(n14307) );
  INV_X1 U9301 ( .A(n14309), .ZN(n21641) );
  AOI22_X1 U9302 ( .A1(\mem[558][1] ), .A2(n14308), .B1(n26572), .B2(
        data_in[1]), .ZN(n14309) );
  INV_X1 U9303 ( .A(n14310), .ZN(n21640) );
  AOI22_X1 U9304 ( .A1(\mem[558][2] ), .A2(n14308), .B1(n26572), .B2(
        data_in[2]), .ZN(n14310) );
  INV_X1 U9305 ( .A(n14311), .ZN(n21639) );
  AOI22_X1 U9306 ( .A1(\mem[558][3] ), .A2(n14308), .B1(n26572), .B2(
        data_in[3]), .ZN(n14311) );
  INV_X1 U9307 ( .A(n14312), .ZN(n21638) );
  AOI22_X1 U9308 ( .A1(\mem[558][4] ), .A2(n14308), .B1(n26572), .B2(
        data_in[4]), .ZN(n14312) );
  INV_X1 U9309 ( .A(n14313), .ZN(n21637) );
  AOI22_X1 U9310 ( .A1(\mem[558][5] ), .A2(n14308), .B1(n26572), .B2(
        data_in[5]), .ZN(n14313) );
  INV_X1 U9311 ( .A(n14314), .ZN(n21636) );
  AOI22_X1 U9312 ( .A1(\mem[558][6] ), .A2(n14308), .B1(n26572), .B2(
        data_in[6]), .ZN(n14314) );
  INV_X1 U9313 ( .A(n14315), .ZN(n21635) );
  AOI22_X1 U9314 ( .A1(\mem[558][7] ), .A2(n14308), .B1(n26572), .B2(
        data_in[7]), .ZN(n14315) );
  INV_X1 U9315 ( .A(n14316), .ZN(n21634) );
  AOI22_X1 U9316 ( .A1(\mem[559][0] ), .A2(n14317), .B1(n26571), .B2(
        data_in[0]), .ZN(n14316) );
  INV_X1 U9317 ( .A(n14318), .ZN(n21633) );
  AOI22_X1 U9318 ( .A1(\mem[559][1] ), .A2(n14317), .B1(n26571), .B2(
        data_in[1]), .ZN(n14318) );
  INV_X1 U9319 ( .A(n14319), .ZN(n21632) );
  AOI22_X1 U9320 ( .A1(\mem[559][2] ), .A2(n14317), .B1(n26571), .B2(
        data_in[2]), .ZN(n14319) );
  INV_X1 U9321 ( .A(n14320), .ZN(n21631) );
  AOI22_X1 U9322 ( .A1(\mem[559][3] ), .A2(n14317), .B1(n26571), .B2(
        data_in[3]), .ZN(n14320) );
  INV_X1 U9323 ( .A(n14321), .ZN(n21630) );
  AOI22_X1 U9324 ( .A1(\mem[559][4] ), .A2(n14317), .B1(n26571), .B2(
        data_in[4]), .ZN(n14321) );
  INV_X1 U9325 ( .A(n14322), .ZN(n21629) );
  AOI22_X1 U9326 ( .A1(\mem[559][5] ), .A2(n14317), .B1(n26571), .B2(
        data_in[5]), .ZN(n14322) );
  INV_X1 U9327 ( .A(n14323), .ZN(n21628) );
  AOI22_X1 U9328 ( .A1(\mem[559][6] ), .A2(n14317), .B1(n26571), .B2(
        data_in[6]), .ZN(n14323) );
  INV_X1 U9329 ( .A(n14324), .ZN(n21627) );
  AOI22_X1 U9330 ( .A1(\mem[559][7] ), .A2(n14317), .B1(n26571), .B2(
        data_in[7]), .ZN(n14324) );
  INV_X1 U9331 ( .A(n14325), .ZN(n21626) );
  AOI22_X1 U9332 ( .A1(\mem[560][0] ), .A2(n14326), .B1(n26570), .B2(
        data_in[0]), .ZN(n14325) );
  INV_X1 U9333 ( .A(n14327), .ZN(n21625) );
  AOI22_X1 U9334 ( .A1(\mem[560][1] ), .A2(n14326), .B1(n26570), .B2(
        data_in[1]), .ZN(n14327) );
  INV_X1 U9335 ( .A(n14328), .ZN(n21624) );
  AOI22_X1 U9336 ( .A1(\mem[560][2] ), .A2(n14326), .B1(n26570), .B2(
        data_in[2]), .ZN(n14328) );
  INV_X1 U9337 ( .A(n14329), .ZN(n21623) );
  AOI22_X1 U9338 ( .A1(\mem[560][3] ), .A2(n14326), .B1(n26570), .B2(
        data_in[3]), .ZN(n14329) );
  INV_X1 U9339 ( .A(n14330), .ZN(n21622) );
  AOI22_X1 U9340 ( .A1(\mem[560][4] ), .A2(n14326), .B1(n26570), .B2(
        data_in[4]), .ZN(n14330) );
  INV_X1 U9341 ( .A(n14331), .ZN(n21621) );
  AOI22_X1 U9342 ( .A1(\mem[560][5] ), .A2(n14326), .B1(n26570), .B2(
        data_in[5]), .ZN(n14331) );
  INV_X1 U9343 ( .A(n14332), .ZN(n21620) );
  AOI22_X1 U9344 ( .A1(\mem[560][6] ), .A2(n14326), .B1(n26570), .B2(
        data_in[6]), .ZN(n14332) );
  INV_X1 U9345 ( .A(n14333), .ZN(n21619) );
  AOI22_X1 U9346 ( .A1(\mem[560][7] ), .A2(n14326), .B1(n26570), .B2(
        data_in[7]), .ZN(n14333) );
  INV_X1 U9347 ( .A(n14334), .ZN(n21618) );
  AOI22_X1 U9348 ( .A1(\mem[561][0] ), .A2(n14335), .B1(n26569), .B2(
        data_in[0]), .ZN(n14334) );
  INV_X1 U9349 ( .A(n14336), .ZN(n21617) );
  AOI22_X1 U9350 ( .A1(\mem[561][1] ), .A2(n14335), .B1(n26569), .B2(
        data_in[1]), .ZN(n14336) );
  INV_X1 U9351 ( .A(n14337), .ZN(n21616) );
  AOI22_X1 U9352 ( .A1(\mem[561][2] ), .A2(n14335), .B1(n26569), .B2(
        data_in[2]), .ZN(n14337) );
  INV_X1 U9353 ( .A(n14338), .ZN(n21615) );
  AOI22_X1 U9354 ( .A1(\mem[561][3] ), .A2(n14335), .B1(n26569), .B2(
        data_in[3]), .ZN(n14338) );
  INV_X1 U9355 ( .A(n14339), .ZN(n21614) );
  AOI22_X1 U9356 ( .A1(\mem[561][4] ), .A2(n14335), .B1(n26569), .B2(
        data_in[4]), .ZN(n14339) );
  INV_X1 U9357 ( .A(n14340), .ZN(n21613) );
  AOI22_X1 U9358 ( .A1(\mem[561][5] ), .A2(n14335), .B1(n26569), .B2(
        data_in[5]), .ZN(n14340) );
  INV_X1 U9359 ( .A(n14341), .ZN(n21612) );
  AOI22_X1 U9360 ( .A1(\mem[561][6] ), .A2(n14335), .B1(n26569), .B2(
        data_in[6]), .ZN(n14341) );
  INV_X1 U9361 ( .A(n14342), .ZN(n21611) );
  AOI22_X1 U9362 ( .A1(\mem[561][7] ), .A2(n14335), .B1(n26569), .B2(
        data_in[7]), .ZN(n14342) );
  INV_X1 U9363 ( .A(n14343), .ZN(n21610) );
  AOI22_X1 U9364 ( .A1(\mem[562][0] ), .A2(n14344), .B1(n26568), .B2(
        data_in[0]), .ZN(n14343) );
  INV_X1 U9365 ( .A(n14345), .ZN(n21609) );
  AOI22_X1 U9366 ( .A1(\mem[562][1] ), .A2(n14344), .B1(n26568), .B2(
        data_in[1]), .ZN(n14345) );
  INV_X1 U9367 ( .A(n14346), .ZN(n21608) );
  AOI22_X1 U9368 ( .A1(\mem[562][2] ), .A2(n14344), .B1(n26568), .B2(
        data_in[2]), .ZN(n14346) );
  INV_X1 U9369 ( .A(n14347), .ZN(n21607) );
  AOI22_X1 U9370 ( .A1(\mem[562][3] ), .A2(n14344), .B1(n26568), .B2(
        data_in[3]), .ZN(n14347) );
  INV_X1 U9371 ( .A(n14348), .ZN(n21606) );
  AOI22_X1 U9372 ( .A1(\mem[562][4] ), .A2(n14344), .B1(n26568), .B2(
        data_in[4]), .ZN(n14348) );
  INV_X1 U9373 ( .A(n14349), .ZN(n21605) );
  AOI22_X1 U9374 ( .A1(\mem[562][5] ), .A2(n14344), .B1(n26568), .B2(
        data_in[5]), .ZN(n14349) );
  INV_X1 U9375 ( .A(n14350), .ZN(n21604) );
  AOI22_X1 U9376 ( .A1(\mem[562][6] ), .A2(n14344), .B1(n26568), .B2(
        data_in[6]), .ZN(n14350) );
  INV_X1 U9377 ( .A(n14351), .ZN(n21603) );
  AOI22_X1 U9378 ( .A1(\mem[562][7] ), .A2(n14344), .B1(n26568), .B2(
        data_in[7]), .ZN(n14351) );
  INV_X1 U9379 ( .A(n14352), .ZN(n21602) );
  AOI22_X1 U9380 ( .A1(\mem[563][0] ), .A2(n14353), .B1(n26567), .B2(
        data_in[0]), .ZN(n14352) );
  INV_X1 U9381 ( .A(n14354), .ZN(n21601) );
  AOI22_X1 U9382 ( .A1(\mem[563][1] ), .A2(n14353), .B1(n26567), .B2(
        data_in[1]), .ZN(n14354) );
  INV_X1 U9383 ( .A(n14355), .ZN(n21600) );
  AOI22_X1 U9384 ( .A1(\mem[563][2] ), .A2(n14353), .B1(n26567), .B2(
        data_in[2]), .ZN(n14355) );
  INV_X1 U9385 ( .A(n14356), .ZN(n21599) );
  AOI22_X1 U9386 ( .A1(\mem[563][3] ), .A2(n14353), .B1(n26567), .B2(
        data_in[3]), .ZN(n14356) );
  INV_X1 U9387 ( .A(n14357), .ZN(n21598) );
  AOI22_X1 U9388 ( .A1(\mem[563][4] ), .A2(n14353), .B1(n26567), .B2(
        data_in[4]), .ZN(n14357) );
  INV_X1 U9389 ( .A(n14358), .ZN(n21597) );
  AOI22_X1 U9390 ( .A1(\mem[563][5] ), .A2(n14353), .B1(n26567), .B2(
        data_in[5]), .ZN(n14358) );
  INV_X1 U9391 ( .A(n14359), .ZN(n21596) );
  AOI22_X1 U9392 ( .A1(\mem[563][6] ), .A2(n14353), .B1(n26567), .B2(
        data_in[6]), .ZN(n14359) );
  INV_X1 U9393 ( .A(n14360), .ZN(n21595) );
  AOI22_X1 U9394 ( .A1(\mem[563][7] ), .A2(n14353), .B1(n26567), .B2(
        data_in[7]), .ZN(n14360) );
  INV_X1 U9395 ( .A(n14361), .ZN(n21594) );
  AOI22_X1 U9396 ( .A1(\mem[564][0] ), .A2(n14362), .B1(n26566), .B2(
        data_in[0]), .ZN(n14361) );
  INV_X1 U9397 ( .A(n14363), .ZN(n21593) );
  AOI22_X1 U9398 ( .A1(\mem[564][1] ), .A2(n14362), .B1(n26566), .B2(
        data_in[1]), .ZN(n14363) );
  INV_X1 U9399 ( .A(n14364), .ZN(n21592) );
  AOI22_X1 U9400 ( .A1(\mem[564][2] ), .A2(n14362), .B1(n26566), .B2(
        data_in[2]), .ZN(n14364) );
  INV_X1 U9401 ( .A(n14365), .ZN(n21591) );
  AOI22_X1 U9402 ( .A1(\mem[564][3] ), .A2(n14362), .B1(n26566), .B2(
        data_in[3]), .ZN(n14365) );
  INV_X1 U9403 ( .A(n14366), .ZN(n21590) );
  AOI22_X1 U9404 ( .A1(\mem[564][4] ), .A2(n14362), .B1(n26566), .B2(
        data_in[4]), .ZN(n14366) );
  INV_X1 U9405 ( .A(n14367), .ZN(n21589) );
  AOI22_X1 U9406 ( .A1(\mem[564][5] ), .A2(n14362), .B1(n26566), .B2(
        data_in[5]), .ZN(n14367) );
  INV_X1 U9407 ( .A(n14368), .ZN(n21588) );
  AOI22_X1 U9408 ( .A1(\mem[564][6] ), .A2(n14362), .B1(n26566), .B2(
        data_in[6]), .ZN(n14368) );
  INV_X1 U9409 ( .A(n14369), .ZN(n21587) );
  AOI22_X1 U9410 ( .A1(\mem[564][7] ), .A2(n14362), .B1(n26566), .B2(
        data_in[7]), .ZN(n14369) );
  INV_X1 U9411 ( .A(n14370), .ZN(n21586) );
  AOI22_X1 U9412 ( .A1(\mem[565][0] ), .A2(n14371), .B1(n26565), .B2(
        data_in[0]), .ZN(n14370) );
  INV_X1 U9413 ( .A(n14372), .ZN(n21585) );
  AOI22_X1 U9414 ( .A1(\mem[565][1] ), .A2(n14371), .B1(n26565), .B2(
        data_in[1]), .ZN(n14372) );
  INV_X1 U9415 ( .A(n14373), .ZN(n21584) );
  AOI22_X1 U9416 ( .A1(\mem[565][2] ), .A2(n14371), .B1(n26565), .B2(
        data_in[2]), .ZN(n14373) );
  INV_X1 U9417 ( .A(n14374), .ZN(n21583) );
  AOI22_X1 U9418 ( .A1(\mem[565][3] ), .A2(n14371), .B1(n26565), .B2(
        data_in[3]), .ZN(n14374) );
  INV_X1 U9419 ( .A(n14375), .ZN(n21582) );
  AOI22_X1 U9420 ( .A1(\mem[565][4] ), .A2(n14371), .B1(n26565), .B2(
        data_in[4]), .ZN(n14375) );
  INV_X1 U9421 ( .A(n14376), .ZN(n21581) );
  AOI22_X1 U9422 ( .A1(\mem[565][5] ), .A2(n14371), .B1(n26565), .B2(
        data_in[5]), .ZN(n14376) );
  INV_X1 U9423 ( .A(n14377), .ZN(n21580) );
  AOI22_X1 U9424 ( .A1(\mem[565][6] ), .A2(n14371), .B1(n26565), .B2(
        data_in[6]), .ZN(n14377) );
  INV_X1 U9425 ( .A(n14378), .ZN(n21579) );
  AOI22_X1 U9426 ( .A1(\mem[565][7] ), .A2(n14371), .B1(n26565), .B2(
        data_in[7]), .ZN(n14378) );
  INV_X1 U9427 ( .A(n14379), .ZN(n21578) );
  AOI22_X1 U9428 ( .A1(\mem[566][0] ), .A2(n14380), .B1(n26564), .B2(
        data_in[0]), .ZN(n14379) );
  INV_X1 U9429 ( .A(n14381), .ZN(n21577) );
  AOI22_X1 U9430 ( .A1(\mem[566][1] ), .A2(n14380), .B1(n26564), .B2(
        data_in[1]), .ZN(n14381) );
  INV_X1 U9431 ( .A(n14382), .ZN(n21576) );
  AOI22_X1 U9432 ( .A1(\mem[566][2] ), .A2(n14380), .B1(n26564), .B2(
        data_in[2]), .ZN(n14382) );
  INV_X1 U9433 ( .A(n14383), .ZN(n21575) );
  AOI22_X1 U9434 ( .A1(\mem[566][3] ), .A2(n14380), .B1(n26564), .B2(
        data_in[3]), .ZN(n14383) );
  INV_X1 U9435 ( .A(n14384), .ZN(n21574) );
  AOI22_X1 U9436 ( .A1(\mem[566][4] ), .A2(n14380), .B1(n26564), .B2(
        data_in[4]), .ZN(n14384) );
  INV_X1 U9437 ( .A(n14385), .ZN(n21573) );
  AOI22_X1 U9438 ( .A1(\mem[566][5] ), .A2(n14380), .B1(n26564), .B2(
        data_in[5]), .ZN(n14385) );
  INV_X1 U9439 ( .A(n14386), .ZN(n21572) );
  AOI22_X1 U9440 ( .A1(\mem[566][6] ), .A2(n14380), .B1(n26564), .B2(
        data_in[6]), .ZN(n14386) );
  INV_X1 U9441 ( .A(n14387), .ZN(n21571) );
  AOI22_X1 U9442 ( .A1(\mem[566][7] ), .A2(n14380), .B1(n26564), .B2(
        data_in[7]), .ZN(n14387) );
  INV_X1 U9443 ( .A(n14388), .ZN(n21570) );
  AOI22_X1 U9444 ( .A1(\mem[567][0] ), .A2(n14389), .B1(n26563), .B2(
        data_in[0]), .ZN(n14388) );
  INV_X1 U9445 ( .A(n14390), .ZN(n21569) );
  AOI22_X1 U9446 ( .A1(\mem[567][1] ), .A2(n14389), .B1(n26563), .B2(
        data_in[1]), .ZN(n14390) );
  INV_X1 U9447 ( .A(n14391), .ZN(n21568) );
  AOI22_X1 U9448 ( .A1(\mem[567][2] ), .A2(n14389), .B1(n26563), .B2(
        data_in[2]), .ZN(n14391) );
  INV_X1 U9449 ( .A(n14392), .ZN(n21567) );
  AOI22_X1 U9450 ( .A1(\mem[567][3] ), .A2(n14389), .B1(n26563), .B2(
        data_in[3]), .ZN(n14392) );
  INV_X1 U9451 ( .A(n14393), .ZN(n21566) );
  AOI22_X1 U9452 ( .A1(\mem[567][4] ), .A2(n14389), .B1(n26563), .B2(
        data_in[4]), .ZN(n14393) );
  INV_X1 U9453 ( .A(n14394), .ZN(n21565) );
  AOI22_X1 U9454 ( .A1(\mem[567][5] ), .A2(n14389), .B1(n26563), .B2(
        data_in[5]), .ZN(n14394) );
  INV_X1 U9455 ( .A(n14395), .ZN(n21564) );
  AOI22_X1 U9456 ( .A1(\mem[567][6] ), .A2(n14389), .B1(n26563), .B2(
        data_in[6]), .ZN(n14395) );
  INV_X1 U9457 ( .A(n14396), .ZN(n21563) );
  AOI22_X1 U9458 ( .A1(\mem[567][7] ), .A2(n14389), .B1(n26563), .B2(
        data_in[7]), .ZN(n14396) );
  INV_X1 U9459 ( .A(n14397), .ZN(n21562) );
  AOI22_X1 U9460 ( .A1(\mem[568][0] ), .A2(n14398), .B1(n26562), .B2(
        data_in[0]), .ZN(n14397) );
  INV_X1 U9461 ( .A(n14399), .ZN(n21561) );
  AOI22_X1 U9462 ( .A1(\mem[568][1] ), .A2(n14398), .B1(n26562), .B2(
        data_in[1]), .ZN(n14399) );
  INV_X1 U9463 ( .A(n14400), .ZN(n21560) );
  AOI22_X1 U9464 ( .A1(\mem[568][2] ), .A2(n14398), .B1(n26562), .B2(
        data_in[2]), .ZN(n14400) );
  INV_X1 U9465 ( .A(n14401), .ZN(n21559) );
  AOI22_X1 U9466 ( .A1(\mem[568][3] ), .A2(n14398), .B1(n26562), .B2(
        data_in[3]), .ZN(n14401) );
  INV_X1 U9467 ( .A(n14402), .ZN(n21558) );
  AOI22_X1 U9468 ( .A1(\mem[568][4] ), .A2(n14398), .B1(n26562), .B2(
        data_in[4]), .ZN(n14402) );
  INV_X1 U9469 ( .A(n14403), .ZN(n21557) );
  AOI22_X1 U9470 ( .A1(\mem[568][5] ), .A2(n14398), .B1(n26562), .B2(
        data_in[5]), .ZN(n14403) );
  INV_X1 U9471 ( .A(n14404), .ZN(n21556) );
  AOI22_X1 U9472 ( .A1(\mem[568][6] ), .A2(n14398), .B1(n26562), .B2(
        data_in[6]), .ZN(n14404) );
  INV_X1 U9473 ( .A(n14405), .ZN(n21555) );
  AOI22_X1 U9474 ( .A1(\mem[568][7] ), .A2(n14398), .B1(n26562), .B2(
        data_in[7]), .ZN(n14405) );
  INV_X1 U9475 ( .A(n14406), .ZN(n21554) );
  AOI22_X1 U9476 ( .A1(\mem[569][0] ), .A2(n14407), .B1(n26561), .B2(
        data_in[0]), .ZN(n14406) );
  INV_X1 U9477 ( .A(n14408), .ZN(n21553) );
  AOI22_X1 U9478 ( .A1(\mem[569][1] ), .A2(n14407), .B1(n26561), .B2(
        data_in[1]), .ZN(n14408) );
  INV_X1 U9479 ( .A(n14409), .ZN(n21552) );
  AOI22_X1 U9480 ( .A1(\mem[569][2] ), .A2(n14407), .B1(n26561), .B2(
        data_in[2]), .ZN(n14409) );
  INV_X1 U9481 ( .A(n14410), .ZN(n21551) );
  AOI22_X1 U9482 ( .A1(\mem[569][3] ), .A2(n14407), .B1(n26561), .B2(
        data_in[3]), .ZN(n14410) );
  INV_X1 U9483 ( .A(n14411), .ZN(n21550) );
  AOI22_X1 U9484 ( .A1(\mem[569][4] ), .A2(n14407), .B1(n26561), .B2(
        data_in[4]), .ZN(n14411) );
  INV_X1 U9485 ( .A(n14412), .ZN(n21549) );
  AOI22_X1 U9486 ( .A1(\mem[569][5] ), .A2(n14407), .B1(n26561), .B2(
        data_in[5]), .ZN(n14412) );
  INV_X1 U9487 ( .A(n14413), .ZN(n21548) );
  AOI22_X1 U9488 ( .A1(\mem[569][6] ), .A2(n14407), .B1(n26561), .B2(
        data_in[6]), .ZN(n14413) );
  INV_X1 U9489 ( .A(n14414), .ZN(n21547) );
  AOI22_X1 U9490 ( .A1(\mem[569][7] ), .A2(n14407), .B1(n26561), .B2(
        data_in[7]), .ZN(n14414) );
  INV_X1 U9491 ( .A(n14415), .ZN(n21546) );
  AOI22_X1 U9492 ( .A1(\mem[570][0] ), .A2(n14416), .B1(n26560), .B2(
        data_in[0]), .ZN(n14415) );
  INV_X1 U9493 ( .A(n14417), .ZN(n21545) );
  AOI22_X1 U9494 ( .A1(\mem[570][1] ), .A2(n14416), .B1(n26560), .B2(
        data_in[1]), .ZN(n14417) );
  INV_X1 U9495 ( .A(n14418), .ZN(n21544) );
  AOI22_X1 U9496 ( .A1(\mem[570][2] ), .A2(n14416), .B1(n26560), .B2(
        data_in[2]), .ZN(n14418) );
  INV_X1 U9497 ( .A(n14419), .ZN(n21543) );
  AOI22_X1 U9498 ( .A1(\mem[570][3] ), .A2(n14416), .B1(n26560), .B2(
        data_in[3]), .ZN(n14419) );
  INV_X1 U9499 ( .A(n14420), .ZN(n21542) );
  AOI22_X1 U9500 ( .A1(\mem[570][4] ), .A2(n14416), .B1(n26560), .B2(
        data_in[4]), .ZN(n14420) );
  INV_X1 U9501 ( .A(n14421), .ZN(n21541) );
  AOI22_X1 U9502 ( .A1(\mem[570][5] ), .A2(n14416), .B1(n26560), .B2(
        data_in[5]), .ZN(n14421) );
  INV_X1 U9503 ( .A(n14422), .ZN(n21540) );
  AOI22_X1 U9504 ( .A1(\mem[570][6] ), .A2(n14416), .B1(n26560), .B2(
        data_in[6]), .ZN(n14422) );
  INV_X1 U9505 ( .A(n14423), .ZN(n21539) );
  AOI22_X1 U9506 ( .A1(\mem[570][7] ), .A2(n14416), .B1(n26560), .B2(
        data_in[7]), .ZN(n14423) );
  INV_X1 U9507 ( .A(n14424), .ZN(n21538) );
  AOI22_X1 U9508 ( .A1(\mem[571][0] ), .A2(n14425), .B1(n26559), .B2(
        data_in[0]), .ZN(n14424) );
  INV_X1 U9509 ( .A(n14426), .ZN(n21537) );
  AOI22_X1 U9510 ( .A1(\mem[571][1] ), .A2(n14425), .B1(n26559), .B2(
        data_in[1]), .ZN(n14426) );
  INV_X1 U9511 ( .A(n14427), .ZN(n21536) );
  AOI22_X1 U9512 ( .A1(\mem[571][2] ), .A2(n14425), .B1(n26559), .B2(
        data_in[2]), .ZN(n14427) );
  INV_X1 U9513 ( .A(n14428), .ZN(n21535) );
  AOI22_X1 U9514 ( .A1(\mem[571][3] ), .A2(n14425), .B1(n26559), .B2(
        data_in[3]), .ZN(n14428) );
  INV_X1 U9515 ( .A(n14429), .ZN(n21534) );
  AOI22_X1 U9516 ( .A1(\mem[571][4] ), .A2(n14425), .B1(n26559), .B2(
        data_in[4]), .ZN(n14429) );
  INV_X1 U9517 ( .A(n14430), .ZN(n21533) );
  AOI22_X1 U9518 ( .A1(\mem[571][5] ), .A2(n14425), .B1(n26559), .B2(
        data_in[5]), .ZN(n14430) );
  INV_X1 U9519 ( .A(n14431), .ZN(n21532) );
  AOI22_X1 U9520 ( .A1(\mem[571][6] ), .A2(n14425), .B1(n26559), .B2(
        data_in[6]), .ZN(n14431) );
  INV_X1 U9521 ( .A(n14432), .ZN(n21531) );
  AOI22_X1 U9522 ( .A1(\mem[571][7] ), .A2(n14425), .B1(n26559), .B2(
        data_in[7]), .ZN(n14432) );
  INV_X1 U9523 ( .A(n14433), .ZN(n21530) );
  AOI22_X1 U9524 ( .A1(\mem[572][0] ), .A2(n14434), .B1(n26558), .B2(
        data_in[0]), .ZN(n14433) );
  INV_X1 U9525 ( .A(n14435), .ZN(n21529) );
  AOI22_X1 U9526 ( .A1(\mem[572][1] ), .A2(n14434), .B1(n26558), .B2(
        data_in[1]), .ZN(n14435) );
  INV_X1 U9527 ( .A(n14436), .ZN(n21528) );
  AOI22_X1 U9528 ( .A1(\mem[572][2] ), .A2(n14434), .B1(n26558), .B2(
        data_in[2]), .ZN(n14436) );
  INV_X1 U9529 ( .A(n14437), .ZN(n21527) );
  AOI22_X1 U9530 ( .A1(\mem[572][3] ), .A2(n14434), .B1(n26558), .B2(
        data_in[3]), .ZN(n14437) );
  INV_X1 U9531 ( .A(n14438), .ZN(n21526) );
  AOI22_X1 U9532 ( .A1(\mem[572][4] ), .A2(n14434), .B1(n26558), .B2(
        data_in[4]), .ZN(n14438) );
  INV_X1 U9533 ( .A(n14439), .ZN(n21525) );
  AOI22_X1 U9534 ( .A1(\mem[572][5] ), .A2(n14434), .B1(n26558), .B2(
        data_in[5]), .ZN(n14439) );
  INV_X1 U9535 ( .A(n14440), .ZN(n21524) );
  AOI22_X1 U9536 ( .A1(\mem[572][6] ), .A2(n14434), .B1(n26558), .B2(
        data_in[6]), .ZN(n14440) );
  INV_X1 U9537 ( .A(n14441), .ZN(n21523) );
  AOI22_X1 U9538 ( .A1(\mem[572][7] ), .A2(n14434), .B1(n26558), .B2(
        data_in[7]), .ZN(n14441) );
  INV_X1 U9539 ( .A(n14442), .ZN(n21522) );
  AOI22_X1 U9540 ( .A1(\mem[573][0] ), .A2(n14443), .B1(n26557), .B2(
        data_in[0]), .ZN(n14442) );
  INV_X1 U9541 ( .A(n14444), .ZN(n21521) );
  AOI22_X1 U9542 ( .A1(\mem[573][1] ), .A2(n14443), .B1(n26557), .B2(
        data_in[1]), .ZN(n14444) );
  INV_X1 U9543 ( .A(n14445), .ZN(n21520) );
  AOI22_X1 U9544 ( .A1(\mem[573][2] ), .A2(n14443), .B1(n26557), .B2(
        data_in[2]), .ZN(n14445) );
  INV_X1 U9545 ( .A(n14446), .ZN(n21519) );
  AOI22_X1 U9546 ( .A1(\mem[573][3] ), .A2(n14443), .B1(n26557), .B2(
        data_in[3]), .ZN(n14446) );
  INV_X1 U9547 ( .A(n14447), .ZN(n21518) );
  AOI22_X1 U9548 ( .A1(\mem[573][4] ), .A2(n14443), .B1(n26557), .B2(
        data_in[4]), .ZN(n14447) );
  INV_X1 U9549 ( .A(n14448), .ZN(n21517) );
  AOI22_X1 U9550 ( .A1(\mem[573][5] ), .A2(n14443), .B1(n26557), .B2(
        data_in[5]), .ZN(n14448) );
  INV_X1 U9551 ( .A(n14449), .ZN(n21516) );
  AOI22_X1 U9552 ( .A1(\mem[573][6] ), .A2(n14443), .B1(n26557), .B2(
        data_in[6]), .ZN(n14449) );
  INV_X1 U9553 ( .A(n14450), .ZN(n21515) );
  AOI22_X1 U9554 ( .A1(\mem[573][7] ), .A2(n14443), .B1(n26557), .B2(
        data_in[7]), .ZN(n14450) );
  INV_X1 U9555 ( .A(n14451), .ZN(n21514) );
  AOI22_X1 U9556 ( .A1(\mem[574][0] ), .A2(n14452), .B1(n26556), .B2(
        data_in[0]), .ZN(n14451) );
  INV_X1 U9557 ( .A(n14453), .ZN(n21513) );
  AOI22_X1 U9558 ( .A1(\mem[574][1] ), .A2(n14452), .B1(n26556), .B2(
        data_in[1]), .ZN(n14453) );
  INV_X1 U9559 ( .A(n14454), .ZN(n21512) );
  AOI22_X1 U9560 ( .A1(\mem[574][2] ), .A2(n14452), .B1(n26556), .B2(
        data_in[2]), .ZN(n14454) );
  INV_X1 U9561 ( .A(n14455), .ZN(n21511) );
  AOI22_X1 U9562 ( .A1(\mem[574][3] ), .A2(n14452), .B1(n26556), .B2(
        data_in[3]), .ZN(n14455) );
  INV_X1 U9563 ( .A(n14456), .ZN(n21510) );
  AOI22_X1 U9564 ( .A1(\mem[574][4] ), .A2(n14452), .B1(n26556), .B2(
        data_in[4]), .ZN(n14456) );
  INV_X1 U9565 ( .A(n14457), .ZN(n21509) );
  AOI22_X1 U9566 ( .A1(\mem[574][5] ), .A2(n14452), .B1(n26556), .B2(
        data_in[5]), .ZN(n14457) );
  INV_X1 U9567 ( .A(n14458), .ZN(n21508) );
  AOI22_X1 U9568 ( .A1(\mem[574][6] ), .A2(n14452), .B1(n26556), .B2(
        data_in[6]), .ZN(n14458) );
  INV_X1 U9569 ( .A(n14459), .ZN(n21507) );
  AOI22_X1 U9570 ( .A1(\mem[574][7] ), .A2(n14452), .B1(n26556), .B2(
        data_in[7]), .ZN(n14459) );
  INV_X1 U9571 ( .A(n14460), .ZN(n21506) );
  AOI22_X1 U9572 ( .A1(\mem[575][0] ), .A2(n14461), .B1(n26555), .B2(
        data_in[0]), .ZN(n14460) );
  INV_X1 U9573 ( .A(n14462), .ZN(n21505) );
  AOI22_X1 U9574 ( .A1(\mem[575][1] ), .A2(n14461), .B1(n26555), .B2(
        data_in[1]), .ZN(n14462) );
  INV_X1 U9575 ( .A(n14463), .ZN(n21504) );
  AOI22_X1 U9576 ( .A1(\mem[575][2] ), .A2(n14461), .B1(n26555), .B2(
        data_in[2]), .ZN(n14463) );
  INV_X1 U9577 ( .A(n14464), .ZN(n21503) );
  AOI22_X1 U9578 ( .A1(\mem[575][3] ), .A2(n14461), .B1(n26555), .B2(
        data_in[3]), .ZN(n14464) );
  INV_X1 U9579 ( .A(n14465), .ZN(n21502) );
  AOI22_X1 U9580 ( .A1(\mem[575][4] ), .A2(n14461), .B1(n26555), .B2(
        data_in[4]), .ZN(n14465) );
  INV_X1 U9581 ( .A(n14466), .ZN(n21501) );
  AOI22_X1 U9582 ( .A1(\mem[575][5] ), .A2(n14461), .B1(n26555), .B2(
        data_in[5]), .ZN(n14466) );
  INV_X1 U9583 ( .A(n14467), .ZN(n21500) );
  AOI22_X1 U9584 ( .A1(\mem[575][6] ), .A2(n14461), .B1(n26555), .B2(
        data_in[6]), .ZN(n14467) );
  INV_X1 U9585 ( .A(n14468), .ZN(n21499) );
  AOI22_X1 U9586 ( .A1(\mem[575][7] ), .A2(n14461), .B1(n26555), .B2(
        data_in[7]), .ZN(n14468) );
  INV_X1 U9587 ( .A(n14542), .ZN(n21434) );
  AOI22_X1 U9588 ( .A1(\mem[584][0] ), .A2(n14543), .B1(n26546), .B2(
        data_in[0]), .ZN(n14542) );
  INV_X1 U9589 ( .A(n14544), .ZN(n21433) );
  AOI22_X1 U9590 ( .A1(\mem[584][1] ), .A2(n14543), .B1(n26546), .B2(
        data_in[1]), .ZN(n14544) );
  INV_X1 U9591 ( .A(n14545), .ZN(n21432) );
  AOI22_X1 U9592 ( .A1(\mem[584][2] ), .A2(n14543), .B1(n26546), .B2(
        data_in[2]), .ZN(n14545) );
  INV_X1 U9593 ( .A(n14546), .ZN(n21431) );
  AOI22_X1 U9594 ( .A1(\mem[584][3] ), .A2(n14543), .B1(n26546), .B2(
        data_in[3]), .ZN(n14546) );
  INV_X1 U9595 ( .A(n14547), .ZN(n21430) );
  AOI22_X1 U9596 ( .A1(\mem[584][4] ), .A2(n14543), .B1(n26546), .B2(
        data_in[4]), .ZN(n14547) );
  INV_X1 U9597 ( .A(n14548), .ZN(n21429) );
  AOI22_X1 U9598 ( .A1(\mem[584][5] ), .A2(n14543), .B1(n26546), .B2(
        data_in[5]), .ZN(n14548) );
  INV_X1 U9599 ( .A(n14549), .ZN(n21428) );
  AOI22_X1 U9600 ( .A1(\mem[584][6] ), .A2(n14543), .B1(n26546), .B2(
        data_in[6]), .ZN(n14549) );
  INV_X1 U9601 ( .A(n14550), .ZN(n21427) );
  AOI22_X1 U9602 ( .A1(\mem[584][7] ), .A2(n14543), .B1(n26546), .B2(
        data_in[7]), .ZN(n14550) );
  INV_X1 U9603 ( .A(n14551), .ZN(n21426) );
  AOI22_X1 U9604 ( .A1(\mem[585][0] ), .A2(n14552), .B1(n26545), .B2(
        data_in[0]), .ZN(n14551) );
  INV_X1 U9605 ( .A(n14553), .ZN(n21425) );
  AOI22_X1 U9606 ( .A1(\mem[585][1] ), .A2(n14552), .B1(n26545), .B2(
        data_in[1]), .ZN(n14553) );
  INV_X1 U9607 ( .A(n14554), .ZN(n21424) );
  AOI22_X1 U9608 ( .A1(\mem[585][2] ), .A2(n14552), .B1(n26545), .B2(
        data_in[2]), .ZN(n14554) );
  INV_X1 U9609 ( .A(n14555), .ZN(n21423) );
  AOI22_X1 U9610 ( .A1(\mem[585][3] ), .A2(n14552), .B1(n26545), .B2(
        data_in[3]), .ZN(n14555) );
  INV_X1 U9611 ( .A(n14556), .ZN(n21422) );
  AOI22_X1 U9612 ( .A1(\mem[585][4] ), .A2(n14552), .B1(n26545), .B2(
        data_in[4]), .ZN(n14556) );
  INV_X1 U9613 ( .A(n14557), .ZN(n21421) );
  AOI22_X1 U9614 ( .A1(\mem[585][5] ), .A2(n14552), .B1(n26545), .B2(
        data_in[5]), .ZN(n14557) );
  INV_X1 U9615 ( .A(n14558), .ZN(n21420) );
  AOI22_X1 U9616 ( .A1(\mem[585][6] ), .A2(n14552), .B1(n26545), .B2(
        data_in[6]), .ZN(n14558) );
  INV_X1 U9617 ( .A(n14559), .ZN(n21419) );
  AOI22_X1 U9618 ( .A1(\mem[585][7] ), .A2(n14552), .B1(n26545), .B2(
        data_in[7]), .ZN(n14559) );
  INV_X1 U9619 ( .A(n14560), .ZN(n21418) );
  AOI22_X1 U9620 ( .A1(\mem[586][0] ), .A2(n14561), .B1(n26544), .B2(
        data_in[0]), .ZN(n14560) );
  INV_X1 U9621 ( .A(n14562), .ZN(n21417) );
  AOI22_X1 U9622 ( .A1(\mem[586][1] ), .A2(n14561), .B1(n26544), .B2(
        data_in[1]), .ZN(n14562) );
  INV_X1 U9623 ( .A(n14563), .ZN(n21416) );
  AOI22_X1 U9624 ( .A1(\mem[586][2] ), .A2(n14561), .B1(n26544), .B2(
        data_in[2]), .ZN(n14563) );
  INV_X1 U9625 ( .A(n14564), .ZN(n21415) );
  AOI22_X1 U9626 ( .A1(\mem[586][3] ), .A2(n14561), .B1(n26544), .B2(
        data_in[3]), .ZN(n14564) );
  INV_X1 U9627 ( .A(n14565), .ZN(n21414) );
  AOI22_X1 U9628 ( .A1(\mem[586][4] ), .A2(n14561), .B1(n26544), .B2(
        data_in[4]), .ZN(n14565) );
  INV_X1 U9629 ( .A(n14566), .ZN(n21413) );
  AOI22_X1 U9630 ( .A1(\mem[586][5] ), .A2(n14561), .B1(n26544), .B2(
        data_in[5]), .ZN(n14566) );
  INV_X1 U9631 ( .A(n14567), .ZN(n21412) );
  AOI22_X1 U9632 ( .A1(\mem[586][6] ), .A2(n14561), .B1(n26544), .B2(
        data_in[6]), .ZN(n14567) );
  INV_X1 U9633 ( .A(n14568), .ZN(n21411) );
  AOI22_X1 U9634 ( .A1(\mem[586][7] ), .A2(n14561), .B1(n26544), .B2(
        data_in[7]), .ZN(n14568) );
  INV_X1 U9635 ( .A(n14569), .ZN(n21410) );
  AOI22_X1 U9636 ( .A1(\mem[587][0] ), .A2(n14570), .B1(n26543), .B2(
        data_in[0]), .ZN(n14569) );
  INV_X1 U9637 ( .A(n14571), .ZN(n21409) );
  AOI22_X1 U9638 ( .A1(\mem[587][1] ), .A2(n14570), .B1(n26543), .B2(
        data_in[1]), .ZN(n14571) );
  INV_X1 U9639 ( .A(n14572), .ZN(n21408) );
  AOI22_X1 U9640 ( .A1(\mem[587][2] ), .A2(n14570), .B1(n26543), .B2(
        data_in[2]), .ZN(n14572) );
  INV_X1 U9641 ( .A(n14573), .ZN(n21407) );
  AOI22_X1 U9642 ( .A1(\mem[587][3] ), .A2(n14570), .B1(n26543), .B2(
        data_in[3]), .ZN(n14573) );
  INV_X1 U9643 ( .A(n14574), .ZN(n21406) );
  AOI22_X1 U9644 ( .A1(\mem[587][4] ), .A2(n14570), .B1(n26543), .B2(
        data_in[4]), .ZN(n14574) );
  INV_X1 U9645 ( .A(n14575), .ZN(n21405) );
  AOI22_X1 U9646 ( .A1(\mem[587][5] ), .A2(n14570), .B1(n26543), .B2(
        data_in[5]), .ZN(n14575) );
  INV_X1 U9647 ( .A(n14576), .ZN(n21404) );
  AOI22_X1 U9648 ( .A1(\mem[587][6] ), .A2(n14570), .B1(n26543), .B2(
        data_in[6]), .ZN(n14576) );
  INV_X1 U9649 ( .A(n14577), .ZN(n21403) );
  AOI22_X1 U9650 ( .A1(\mem[587][7] ), .A2(n14570), .B1(n26543), .B2(
        data_in[7]), .ZN(n14577) );
  INV_X1 U9651 ( .A(n14578), .ZN(n21402) );
  AOI22_X1 U9652 ( .A1(\mem[588][0] ), .A2(n14579), .B1(n26542), .B2(
        data_in[0]), .ZN(n14578) );
  INV_X1 U9653 ( .A(n14580), .ZN(n21401) );
  AOI22_X1 U9654 ( .A1(\mem[588][1] ), .A2(n14579), .B1(n26542), .B2(
        data_in[1]), .ZN(n14580) );
  INV_X1 U9655 ( .A(n14581), .ZN(n21400) );
  AOI22_X1 U9656 ( .A1(\mem[588][2] ), .A2(n14579), .B1(n26542), .B2(
        data_in[2]), .ZN(n14581) );
  INV_X1 U9657 ( .A(n14582), .ZN(n21399) );
  AOI22_X1 U9658 ( .A1(\mem[588][3] ), .A2(n14579), .B1(n26542), .B2(
        data_in[3]), .ZN(n14582) );
  INV_X1 U9659 ( .A(n14583), .ZN(n21398) );
  AOI22_X1 U9660 ( .A1(\mem[588][4] ), .A2(n14579), .B1(n26542), .B2(
        data_in[4]), .ZN(n14583) );
  INV_X1 U9661 ( .A(n14584), .ZN(n21397) );
  AOI22_X1 U9662 ( .A1(\mem[588][5] ), .A2(n14579), .B1(n26542), .B2(
        data_in[5]), .ZN(n14584) );
  INV_X1 U9663 ( .A(n14585), .ZN(n21396) );
  AOI22_X1 U9664 ( .A1(\mem[588][6] ), .A2(n14579), .B1(n26542), .B2(
        data_in[6]), .ZN(n14585) );
  INV_X1 U9665 ( .A(n14586), .ZN(n21395) );
  AOI22_X1 U9666 ( .A1(\mem[588][7] ), .A2(n14579), .B1(n26542), .B2(
        data_in[7]), .ZN(n14586) );
  INV_X1 U9667 ( .A(n14587), .ZN(n21394) );
  AOI22_X1 U9668 ( .A1(\mem[589][0] ), .A2(n14588), .B1(n26541), .B2(
        data_in[0]), .ZN(n14587) );
  INV_X1 U9669 ( .A(n14589), .ZN(n21393) );
  AOI22_X1 U9670 ( .A1(\mem[589][1] ), .A2(n14588), .B1(n26541), .B2(
        data_in[1]), .ZN(n14589) );
  INV_X1 U9671 ( .A(n14590), .ZN(n21392) );
  AOI22_X1 U9672 ( .A1(\mem[589][2] ), .A2(n14588), .B1(n26541), .B2(
        data_in[2]), .ZN(n14590) );
  INV_X1 U9673 ( .A(n14591), .ZN(n21391) );
  AOI22_X1 U9674 ( .A1(\mem[589][3] ), .A2(n14588), .B1(n26541), .B2(
        data_in[3]), .ZN(n14591) );
  INV_X1 U9675 ( .A(n14592), .ZN(n21390) );
  AOI22_X1 U9676 ( .A1(\mem[589][4] ), .A2(n14588), .B1(n26541), .B2(
        data_in[4]), .ZN(n14592) );
  INV_X1 U9677 ( .A(n14593), .ZN(n21389) );
  AOI22_X1 U9678 ( .A1(\mem[589][5] ), .A2(n14588), .B1(n26541), .B2(
        data_in[5]), .ZN(n14593) );
  INV_X1 U9679 ( .A(n14594), .ZN(n21388) );
  AOI22_X1 U9680 ( .A1(\mem[589][6] ), .A2(n14588), .B1(n26541), .B2(
        data_in[6]), .ZN(n14594) );
  INV_X1 U9681 ( .A(n14595), .ZN(n21387) );
  AOI22_X1 U9682 ( .A1(\mem[589][7] ), .A2(n14588), .B1(n26541), .B2(
        data_in[7]), .ZN(n14595) );
  INV_X1 U9683 ( .A(n14596), .ZN(n21386) );
  AOI22_X1 U9684 ( .A1(\mem[590][0] ), .A2(n14597), .B1(n26540), .B2(
        data_in[0]), .ZN(n14596) );
  INV_X1 U9685 ( .A(n14598), .ZN(n21385) );
  AOI22_X1 U9686 ( .A1(\mem[590][1] ), .A2(n14597), .B1(n26540), .B2(
        data_in[1]), .ZN(n14598) );
  INV_X1 U9687 ( .A(n14599), .ZN(n21384) );
  AOI22_X1 U9688 ( .A1(\mem[590][2] ), .A2(n14597), .B1(n26540), .B2(
        data_in[2]), .ZN(n14599) );
  INV_X1 U9689 ( .A(n14600), .ZN(n21383) );
  AOI22_X1 U9690 ( .A1(\mem[590][3] ), .A2(n14597), .B1(n26540), .B2(
        data_in[3]), .ZN(n14600) );
  INV_X1 U9691 ( .A(n14601), .ZN(n21382) );
  AOI22_X1 U9692 ( .A1(\mem[590][4] ), .A2(n14597), .B1(n26540), .B2(
        data_in[4]), .ZN(n14601) );
  INV_X1 U9693 ( .A(n14602), .ZN(n21381) );
  AOI22_X1 U9694 ( .A1(\mem[590][5] ), .A2(n14597), .B1(n26540), .B2(
        data_in[5]), .ZN(n14602) );
  INV_X1 U9695 ( .A(n14603), .ZN(n21380) );
  AOI22_X1 U9696 ( .A1(\mem[590][6] ), .A2(n14597), .B1(n26540), .B2(
        data_in[6]), .ZN(n14603) );
  INV_X1 U9697 ( .A(n14604), .ZN(n21379) );
  AOI22_X1 U9698 ( .A1(\mem[590][7] ), .A2(n14597), .B1(n26540), .B2(
        data_in[7]), .ZN(n14604) );
  INV_X1 U9699 ( .A(n14605), .ZN(n21378) );
  AOI22_X1 U9700 ( .A1(\mem[591][0] ), .A2(n14606), .B1(n26539), .B2(
        data_in[0]), .ZN(n14605) );
  INV_X1 U9701 ( .A(n14607), .ZN(n21377) );
  AOI22_X1 U9702 ( .A1(\mem[591][1] ), .A2(n14606), .B1(n26539), .B2(
        data_in[1]), .ZN(n14607) );
  INV_X1 U9703 ( .A(n14608), .ZN(n21376) );
  AOI22_X1 U9704 ( .A1(\mem[591][2] ), .A2(n14606), .B1(n26539), .B2(
        data_in[2]), .ZN(n14608) );
  INV_X1 U9705 ( .A(n14609), .ZN(n21375) );
  AOI22_X1 U9706 ( .A1(\mem[591][3] ), .A2(n14606), .B1(n26539), .B2(
        data_in[3]), .ZN(n14609) );
  INV_X1 U9707 ( .A(n14610), .ZN(n21374) );
  AOI22_X1 U9708 ( .A1(\mem[591][4] ), .A2(n14606), .B1(n26539), .B2(
        data_in[4]), .ZN(n14610) );
  INV_X1 U9709 ( .A(n14611), .ZN(n21373) );
  AOI22_X1 U9710 ( .A1(\mem[591][5] ), .A2(n14606), .B1(n26539), .B2(
        data_in[5]), .ZN(n14611) );
  INV_X1 U9711 ( .A(n14612), .ZN(n21372) );
  AOI22_X1 U9712 ( .A1(\mem[591][6] ), .A2(n14606), .B1(n26539), .B2(
        data_in[6]), .ZN(n14612) );
  INV_X1 U9713 ( .A(n14613), .ZN(n21371) );
  AOI22_X1 U9714 ( .A1(\mem[591][7] ), .A2(n14606), .B1(n26539), .B2(
        data_in[7]), .ZN(n14613) );
  INV_X1 U9715 ( .A(n14614), .ZN(n21370) );
  AOI22_X1 U9716 ( .A1(\mem[592][0] ), .A2(n14615), .B1(n26538), .B2(
        data_in[0]), .ZN(n14614) );
  INV_X1 U9717 ( .A(n14616), .ZN(n21369) );
  AOI22_X1 U9718 ( .A1(\mem[592][1] ), .A2(n14615), .B1(n26538), .B2(
        data_in[1]), .ZN(n14616) );
  INV_X1 U9719 ( .A(n14617), .ZN(n21368) );
  AOI22_X1 U9720 ( .A1(\mem[592][2] ), .A2(n14615), .B1(n26538), .B2(
        data_in[2]), .ZN(n14617) );
  INV_X1 U9721 ( .A(n14618), .ZN(n21367) );
  AOI22_X1 U9722 ( .A1(\mem[592][3] ), .A2(n14615), .B1(n26538), .B2(
        data_in[3]), .ZN(n14618) );
  INV_X1 U9723 ( .A(n14619), .ZN(n21366) );
  AOI22_X1 U9724 ( .A1(\mem[592][4] ), .A2(n14615), .B1(n26538), .B2(
        data_in[4]), .ZN(n14619) );
  INV_X1 U9725 ( .A(n14620), .ZN(n21365) );
  AOI22_X1 U9726 ( .A1(\mem[592][5] ), .A2(n14615), .B1(n26538), .B2(
        data_in[5]), .ZN(n14620) );
  INV_X1 U9727 ( .A(n14621), .ZN(n21364) );
  AOI22_X1 U9728 ( .A1(\mem[592][6] ), .A2(n14615), .B1(n26538), .B2(
        data_in[6]), .ZN(n14621) );
  INV_X1 U9729 ( .A(n14622), .ZN(n21363) );
  AOI22_X1 U9730 ( .A1(\mem[592][7] ), .A2(n14615), .B1(n26538), .B2(
        data_in[7]), .ZN(n14622) );
  INV_X1 U9731 ( .A(n14623), .ZN(n21362) );
  AOI22_X1 U9732 ( .A1(\mem[593][0] ), .A2(n14624), .B1(n26537), .B2(
        data_in[0]), .ZN(n14623) );
  INV_X1 U9733 ( .A(n14625), .ZN(n21361) );
  AOI22_X1 U9734 ( .A1(\mem[593][1] ), .A2(n14624), .B1(n26537), .B2(
        data_in[1]), .ZN(n14625) );
  INV_X1 U9735 ( .A(n14626), .ZN(n21360) );
  AOI22_X1 U9736 ( .A1(\mem[593][2] ), .A2(n14624), .B1(n26537), .B2(
        data_in[2]), .ZN(n14626) );
  INV_X1 U9737 ( .A(n14627), .ZN(n21359) );
  AOI22_X1 U9738 ( .A1(\mem[593][3] ), .A2(n14624), .B1(n26537), .B2(
        data_in[3]), .ZN(n14627) );
  INV_X1 U9739 ( .A(n14628), .ZN(n21358) );
  AOI22_X1 U9740 ( .A1(\mem[593][4] ), .A2(n14624), .B1(n26537), .B2(
        data_in[4]), .ZN(n14628) );
  INV_X1 U9741 ( .A(n14629), .ZN(n21357) );
  AOI22_X1 U9742 ( .A1(\mem[593][5] ), .A2(n14624), .B1(n26537), .B2(
        data_in[5]), .ZN(n14629) );
  INV_X1 U9743 ( .A(n14630), .ZN(n21356) );
  AOI22_X1 U9744 ( .A1(\mem[593][6] ), .A2(n14624), .B1(n26537), .B2(
        data_in[6]), .ZN(n14630) );
  INV_X1 U9745 ( .A(n14631), .ZN(n21355) );
  AOI22_X1 U9746 ( .A1(\mem[593][7] ), .A2(n14624), .B1(n26537), .B2(
        data_in[7]), .ZN(n14631) );
  INV_X1 U9747 ( .A(n14632), .ZN(n21354) );
  AOI22_X1 U9748 ( .A1(\mem[594][0] ), .A2(n14633), .B1(n26536), .B2(
        data_in[0]), .ZN(n14632) );
  INV_X1 U9749 ( .A(n14634), .ZN(n21353) );
  AOI22_X1 U9750 ( .A1(\mem[594][1] ), .A2(n14633), .B1(n26536), .B2(
        data_in[1]), .ZN(n14634) );
  INV_X1 U9751 ( .A(n14635), .ZN(n21352) );
  AOI22_X1 U9752 ( .A1(\mem[594][2] ), .A2(n14633), .B1(n26536), .B2(
        data_in[2]), .ZN(n14635) );
  INV_X1 U9753 ( .A(n14636), .ZN(n21351) );
  AOI22_X1 U9754 ( .A1(\mem[594][3] ), .A2(n14633), .B1(n26536), .B2(
        data_in[3]), .ZN(n14636) );
  INV_X1 U9755 ( .A(n14637), .ZN(n21350) );
  AOI22_X1 U9756 ( .A1(\mem[594][4] ), .A2(n14633), .B1(n26536), .B2(
        data_in[4]), .ZN(n14637) );
  INV_X1 U9757 ( .A(n14638), .ZN(n21349) );
  AOI22_X1 U9758 ( .A1(\mem[594][5] ), .A2(n14633), .B1(n26536), .B2(
        data_in[5]), .ZN(n14638) );
  INV_X1 U9759 ( .A(n14639), .ZN(n21348) );
  AOI22_X1 U9760 ( .A1(\mem[594][6] ), .A2(n14633), .B1(n26536), .B2(
        data_in[6]), .ZN(n14639) );
  INV_X1 U9761 ( .A(n14640), .ZN(n21347) );
  AOI22_X1 U9762 ( .A1(\mem[594][7] ), .A2(n14633), .B1(n26536), .B2(
        data_in[7]), .ZN(n14640) );
  INV_X1 U9763 ( .A(n14641), .ZN(n21346) );
  AOI22_X1 U9764 ( .A1(\mem[595][0] ), .A2(n14642), .B1(n26535), .B2(
        data_in[0]), .ZN(n14641) );
  INV_X1 U9765 ( .A(n14643), .ZN(n21345) );
  AOI22_X1 U9766 ( .A1(\mem[595][1] ), .A2(n14642), .B1(n26535), .B2(
        data_in[1]), .ZN(n14643) );
  INV_X1 U9767 ( .A(n14644), .ZN(n21344) );
  AOI22_X1 U9768 ( .A1(\mem[595][2] ), .A2(n14642), .B1(n26535), .B2(
        data_in[2]), .ZN(n14644) );
  INV_X1 U9769 ( .A(n14645), .ZN(n21343) );
  AOI22_X1 U9770 ( .A1(\mem[595][3] ), .A2(n14642), .B1(n26535), .B2(
        data_in[3]), .ZN(n14645) );
  INV_X1 U9771 ( .A(n14646), .ZN(n21342) );
  AOI22_X1 U9772 ( .A1(\mem[595][4] ), .A2(n14642), .B1(n26535), .B2(
        data_in[4]), .ZN(n14646) );
  INV_X1 U9773 ( .A(n14647), .ZN(n21341) );
  AOI22_X1 U9774 ( .A1(\mem[595][5] ), .A2(n14642), .B1(n26535), .B2(
        data_in[5]), .ZN(n14647) );
  INV_X1 U9775 ( .A(n14648), .ZN(n21340) );
  AOI22_X1 U9776 ( .A1(\mem[595][6] ), .A2(n14642), .B1(n26535), .B2(
        data_in[6]), .ZN(n14648) );
  INV_X1 U9777 ( .A(n14649), .ZN(n21339) );
  AOI22_X1 U9778 ( .A1(\mem[595][7] ), .A2(n14642), .B1(n26535), .B2(
        data_in[7]), .ZN(n14649) );
  INV_X1 U9779 ( .A(n14650), .ZN(n21338) );
  AOI22_X1 U9780 ( .A1(\mem[596][0] ), .A2(n14651), .B1(n26534), .B2(
        data_in[0]), .ZN(n14650) );
  INV_X1 U9781 ( .A(n14652), .ZN(n21337) );
  AOI22_X1 U9782 ( .A1(\mem[596][1] ), .A2(n14651), .B1(n26534), .B2(
        data_in[1]), .ZN(n14652) );
  INV_X1 U9783 ( .A(n14653), .ZN(n21336) );
  AOI22_X1 U9784 ( .A1(\mem[596][2] ), .A2(n14651), .B1(n26534), .B2(
        data_in[2]), .ZN(n14653) );
  INV_X1 U9785 ( .A(n14654), .ZN(n21335) );
  AOI22_X1 U9786 ( .A1(\mem[596][3] ), .A2(n14651), .B1(n26534), .B2(
        data_in[3]), .ZN(n14654) );
  INV_X1 U9787 ( .A(n14655), .ZN(n21334) );
  AOI22_X1 U9788 ( .A1(\mem[596][4] ), .A2(n14651), .B1(n26534), .B2(
        data_in[4]), .ZN(n14655) );
  INV_X1 U9789 ( .A(n14656), .ZN(n21333) );
  AOI22_X1 U9790 ( .A1(\mem[596][5] ), .A2(n14651), .B1(n26534), .B2(
        data_in[5]), .ZN(n14656) );
  INV_X1 U9791 ( .A(n14657), .ZN(n21332) );
  AOI22_X1 U9792 ( .A1(\mem[596][6] ), .A2(n14651), .B1(n26534), .B2(
        data_in[6]), .ZN(n14657) );
  INV_X1 U9793 ( .A(n14658), .ZN(n21331) );
  AOI22_X1 U9794 ( .A1(\mem[596][7] ), .A2(n14651), .B1(n26534), .B2(
        data_in[7]), .ZN(n14658) );
  INV_X1 U9795 ( .A(n14659), .ZN(n21330) );
  AOI22_X1 U9796 ( .A1(\mem[597][0] ), .A2(n14660), .B1(n26533), .B2(
        data_in[0]), .ZN(n14659) );
  INV_X1 U9797 ( .A(n14661), .ZN(n21329) );
  AOI22_X1 U9798 ( .A1(\mem[597][1] ), .A2(n14660), .B1(n26533), .B2(
        data_in[1]), .ZN(n14661) );
  INV_X1 U9799 ( .A(n14662), .ZN(n21328) );
  AOI22_X1 U9800 ( .A1(\mem[597][2] ), .A2(n14660), .B1(n26533), .B2(
        data_in[2]), .ZN(n14662) );
  INV_X1 U9801 ( .A(n14663), .ZN(n21327) );
  AOI22_X1 U9802 ( .A1(\mem[597][3] ), .A2(n14660), .B1(n26533), .B2(
        data_in[3]), .ZN(n14663) );
  INV_X1 U9803 ( .A(n14664), .ZN(n21326) );
  AOI22_X1 U9804 ( .A1(\mem[597][4] ), .A2(n14660), .B1(n26533), .B2(
        data_in[4]), .ZN(n14664) );
  INV_X1 U9805 ( .A(n14665), .ZN(n21325) );
  AOI22_X1 U9806 ( .A1(\mem[597][5] ), .A2(n14660), .B1(n26533), .B2(
        data_in[5]), .ZN(n14665) );
  INV_X1 U9807 ( .A(n14666), .ZN(n21324) );
  AOI22_X1 U9808 ( .A1(\mem[597][6] ), .A2(n14660), .B1(n26533), .B2(
        data_in[6]), .ZN(n14666) );
  INV_X1 U9809 ( .A(n14667), .ZN(n21323) );
  AOI22_X1 U9810 ( .A1(\mem[597][7] ), .A2(n14660), .B1(n26533), .B2(
        data_in[7]), .ZN(n14667) );
  INV_X1 U9811 ( .A(n14668), .ZN(n21322) );
  AOI22_X1 U9812 ( .A1(\mem[598][0] ), .A2(n14669), .B1(n26532), .B2(
        data_in[0]), .ZN(n14668) );
  INV_X1 U9813 ( .A(n14670), .ZN(n21321) );
  AOI22_X1 U9814 ( .A1(\mem[598][1] ), .A2(n14669), .B1(n26532), .B2(
        data_in[1]), .ZN(n14670) );
  INV_X1 U9815 ( .A(n14671), .ZN(n21320) );
  AOI22_X1 U9816 ( .A1(\mem[598][2] ), .A2(n14669), .B1(n26532), .B2(
        data_in[2]), .ZN(n14671) );
  INV_X1 U9817 ( .A(n14672), .ZN(n21319) );
  AOI22_X1 U9818 ( .A1(\mem[598][3] ), .A2(n14669), .B1(n26532), .B2(
        data_in[3]), .ZN(n14672) );
  INV_X1 U9819 ( .A(n14673), .ZN(n21318) );
  AOI22_X1 U9820 ( .A1(\mem[598][4] ), .A2(n14669), .B1(n26532), .B2(
        data_in[4]), .ZN(n14673) );
  INV_X1 U9821 ( .A(n14674), .ZN(n21317) );
  AOI22_X1 U9822 ( .A1(\mem[598][5] ), .A2(n14669), .B1(n26532), .B2(
        data_in[5]), .ZN(n14674) );
  INV_X1 U9823 ( .A(n14675), .ZN(n21316) );
  AOI22_X1 U9824 ( .A1(\mem[598][6] ), .A2(n14669), .B1(n26532), .B2(
        data_in[6]), .ZN(n14675) );
  INV_X1 U9825 ( .A(n14676), .ZN(n21315) );
  AOI22_X1 U9826 ( .A1(\mem[598][7] ), .A2(n14669), .B1(n26532), .B2(
        data_in[7]), .ZN(n14676) );
  INV_X1 U9827 ( .A(n14677), .ZN(n21314) );
  AOI22_X1 U9828 ( .A1(\mem[599][0] ), .A2(n14678), .B1(n26531), .B2(
        data_in[0]), .ZN(n14677) );
  INV_X1 U9829 ( .A(n14679), .ZN(n21313) );
  AOI22_X1 U9830 ( .A1(\mem[599][1] ), .A2(n14678), .B1(n26531), .B2(
        data_in[1]), .ZN(n14679) );
  INV_X1 U9831 ( .A(n14680), .ZN(n21312) );
  AOI22_X1 U9832 ( .A1(\mem[599][2] ), .A2(n14678), .B1(n26531), .B2(
        data_in[2]), .ZN(n14680) );
  INV_X1 U9833 ( .A(n14681), .ZN(n21311) );
  AOI22_X1 U9834 ( .A1(\mem[599][3] ), .A2(n14678), .B1(n26531), .B2(
        data_in[3]), .ZN(n14681) );
  INV_X1 U9835 ( .A(n14682), .ZN(n21310) );
  AOI22_X1 U9836 ( .A1(\mem[599][4] ), .A2(n14678), .B1(n26531), .B2(
        data_in[4]), .ZN(n14682) );
  INV_X1 U9837 ( .A(n14683), .ZN(n21309) );
  AOI22_X1 U9838 ( .A1(\mem[599][5] ), .A2(n14678), .B1(n26531), .B2(
        data_in[5]), .ZN(n14683) );
  INV_X1 U9839 ( .A(n14684), .ZN(n21308) );
  AOI22_X1 U9840 ( .A1(\mem[599][6] ), .A2(n14678), .B1(n26531), .B2(
        data_in[6]), .ZN(n14684) );
  INV_X1 U9841 ( .A(n14685), .ZN(n21307) );
  AOI22_X1 U9842 ( .A1(\mem[599][7] ), .A2(n14678), .B1(n26531), .B2(
        data_in[7]), .ZN(n14685) );
  INV_X1 U9843 ( .A(n14686), .ZN(n21306) );
  AOI22_X1 U9844 ( .A1(\mem[600][0] ), .A2(n14687), .B1(n26530), .B2(
        data_in[0]), .ZN(n14686) );
  INV_X1 U9845 ( .A(n14688), .ZN(n21305) );
  AOI22_X1 U9846 ( .A1(\mem[600][1] ), .A2(n14687), .B1(n26530), .B2(
        data_in[1]), .ZN(n14688) );
  INV_X1 U9847 ( .A(n14689), .ZN(n21304) );
  AOI22_X1 U9848 ( .A1(\mem[600][2] ), .A2(n14687), .B1(n26530), .B2(
        data_in[2]), .ZN(n14689) );
  INV_X1 U9849 ( .A(n14690), .ZN(n21303) );
  AOI22_X1 U9850 ( .A1(\mem[600][3] ), .A2(n14687), .B1(n26530), .B2(
        data_in[3]), .ZN(n14690) );
  INV_X1 U9851 ( .A(n14691), .ZN(n21302) );
  AOI22_X1 U9852 ( .A1(\mem[600][4] ), .A2(n14687), .B1(n26530), .B2(
        data_in[4]), .ZN(n14691) );
  INV_X1 U9853 ( .A(n14692), .ZN(n21301) );
  AOI22_X1 U9854 ( .A1(\mem[600][5] ), .A2(n14687), .B1(n26530), .B2(
        data_in[5]), .ZN(n14692) );
  INV_X1 U9855 ( .A(n14693), .ZN(n21300) );
  AOI22_X1 U9856 ( .A1(\mem[600][6] ), .A2(n14687), .B1(n26530), .B2(
        data_in[6]), .ZN(n14693) );
  INV_X1 U9857 ( .A(n14694), .ZN(n21299) );
  AOI22_X1 U9858 ( .A1(\mem[600][7] ), .A2(n14687), .B1(n26530), .B2(
        data_in[7]), .ZN(n14694) );
  INV_X1 U9859 ( .A(n14695), .ZN(n21298) );
  AOI22_X1 U9860 ( .A1(\mem[601][0] ), .A2(n14696), .B1(n26529), .B2(
        data_in[0]), .ZN(n14695) );
  INV_X1 U9861 ( .A(n14697), .ZN(n21297) );
  AOI22_X1 U9862 ( .A1(\mem[601][1] ), .A2(n14696), .B1(n26529), .B2(
        data_in[1]), .ZN(n14697) );
  INV_X1 U9863 ( .A(n14698), .ZN(n21296) );
  AOI22_X1 U9864 ( .A1(\mem[601][2] ), .A2(n14696), .B1(n26529), .B2(
        data_in[2]), .ZN(n14698) );
  INV_X1 U9865 ( .A(n14699), .ZN(n21295) );
  AOI22_X1 U9866 ( .A1(\mem[601][3] ), .A2(n14696), .B1(n26529), .B2(
        data_in[3]), .ZN(n14699) );
  INV_X1 U9867 ( .A(n14700), .ZN(n21294) );
  AOI22_X1 U9868 ( .A1(\mem[601][4] ), .A2(n14696), .B1(n26529), .B2(
        data_in[4]), .ZN(n14700) );
  INV_X1 U9869 ( .A(n14701), .ZN(n21293) );
  AOI22_X1 U9870 ( .A1(\mem[601][5] ), .A2(n14696), .B1(n26529), .B2(
        data_in[5]), .ZN(n14701) );
  INV_X1 U9871 ( .A(n14702), .ZN(n21292) );
  AOI22_X1 U9872 ( .A1(\mem[601][6] ), .A2(n14696), .B1(n26529), .B2(
        data_in[6]), .ZN(n14702) );
  INV_X1 U9873 ( .A(n14703), .ZN(n21291) );
  AOI22_X1 U9874 ( .A1(\mem[601][7] ), .A2(n14696), .B1(n26529), .B2(
        data_in[7]), .ZN(n14703) );
  INV_X1 U9875 ( .A(n14704), .ZN(n21290) );
  AOI22_X1 U9876 ( .A1(\mem[602][0] ), .A2(n14705), .B1(n26528), .B2(
        data_in[0]), .ZN(n14704) );
  INV_X1 U9877 ( .A(n14706), .ZN(n21289) );
  AOI22_X1 U9878 ( .A1(\mem[602][1] ), .A2(n14705), .B1(n26528), .B2(
        data_in[1]), .ZN(n14706) );
  INV_X1 U9879 ( .A(n14707), .ZN(n21288) );
  AOI22_X1 U9880 ( .A1(\mem[602][2] ), .A2(n14705), .B1(n26528), .B2(
        data_in[2]), .ZN(n14707) );
  INV_X1 U9881 ( .A(n14708), .ZN(n21287) );
  AOI22_X1 U9882 ( .A1(\mem[602][3] ), .A2(n14705), .B1(n26528), .B2(
        data_in[3]), .ZN(n14708) );
  INV_X1 U9883 ( .A(n14709), .ZN(n21286) );
  AOI22_X1 U9884 ( .A1(\mem[602][4] ), .A2(n14705), .B1(n26528), .B2(
        data_in[4]), .ZN(n14709) );
  INV_X1 U9885 ( .A(n14710), .ZN(n21285) );
  AOI22_X1 U9886 ( .A1(\mem[602][5] ), .A2(n14705), .B1(n26528), .B2(
        data_in[5]), .ZN(n14710) );
  INV_X1 U9887 ( .A(n14711), .ZN(n21284) );
  AOI22_X1 U9888 ( .A1(\mem[602][6] ), .A2(n14705), .B1(n26528), .B2(
        data_in[6]), .ZN(n14711) );
  INV_X1 U9889 ( .A(n14712), .ZN(n21283) );
  AOI22_X1 U9890 ( .A1(\mem[602][7] ), .A2(n14705), .B1(n26528), .B2(
        data_in[7]), .ZN(n14712) );
  INV_X1 U9891 ( .A(n14713), .ZN(n21282) );
  AOI22_X1 U9892 ( .A1(\mem[603][0] ), .A2(n14714), .B1(n26527), .B2(
        data_in[0]), .ZN(n14713) );
  INV_X1 U9893 ( .A(n14715), .ZN(n21281) );
  AOI22_X1 U9894 ( .A1(\mem[603][1] ), .A2(n14714), .B1(n26527), .B2(
        data_in[1]), .ZN(n14715) );
  INV_X1 U9895 ( .A(n14716), .ZN(n21280) );
  AOI22_X1 U9896 ( .A1(\mem[603][2] ), .A2(n14714), .B1(n26527), .B2(
        data_in[2]), .ZN(n14716) );
  INV_X1 U9897 ( .A(n14717), .ZN(n21279) );
  AOI22_X1 U9898 ( .A1(\mem[603][3] ), .A2(n14714), .B1(n26527), .B2(
        data_in[3]), .ZN(n14717) );
  INV_X1 U9899 ( .A(n14718), .ZN(n21278) );
  AOI22_X1 U9900 ( .A1(\mem[603][4] ), .A2(n14714), .B1(n26527), .B2(
        data_in[4]), .ZN(n14718) );
  INV_X1 U9901 ( .A(n14719), .ZN(n21277) );
  AOI22_X1 U9902 ( .A1(\mem[603][5] ), .A2(n14714), .B1(n26527), .B2(
        data_in[5]), .ZN(n14719) );
  INV_X1 U9903 ( .A(n14720), .ZN(n21276) );
  AOI22_X1 U9904 ( .A1(\mem[603][6] ), .A2(n14714), .B1(n26527), .B2(
        data_in[6]), .ZN(n14720) );
  INV_X1 U9905 ( .A(n14721), .ZN(n21275) );
  AOI22_X1 U9906 ( .A1(\mem[603][7] ), .A2(n14714), .B1(n26527), .B2(
        data_in[7]), .ZN(n14721) );
  INV_X1 U9907 ( .A(n14722), .ZN(n21274) );
  AOI22_X1 U9908 ( .A1(\mem[604][0] ), .A2(n14723), .B1(n26526), .B2(
        data_in[0]), .ZN(n14722) );
  INV_X1 U9909 ( .A(n14724), .ZN(n21273) );
  AOI22_X1 U9910 ( .A1(\mem[604][1] ), .A2(n14723), .B1(n26526), .B2(
        data_in[1]), .ZN(n14724) );
  INV_X1 U9911 ( .A(n14725), .ZN(n21272) );
  AOI22_X1 U9912 ( .A1(\mem[604][2] ), .A2(n14723), .B1(n26526), .B2(
        data_in[2]), .ZN(n14725) );
  INV_X1 U9913 ( .A(n14726), .ZN(n21271) );
  AOI22_X1 U9914 ( .A1(\mem[604][3] ), .A2(n14723), .B1(n26526), .B2(
        data_in[3]), .ZN(n14726) );
  INV_X1 U9915 ( .A(n14727), .ZN(n21270) );
  AOI22_X1 U9916 ( .A1(\mem[604][4] ), .A2(n14723), .B1(n26526), .B2(
        data_in[4]), .ZN(n14727) );
  INV_X1 U9917 ( .A(n14728), .ZN(n21269) );
  AOI22_X1 U9918 ( .A1(\mem[604][5] ), .A2(n14723), .B1(n26526), .B2(
        data_in[5]), .ZN(n14728) );
  INV_X1 U9919 ( .A(n14729), .ZN(n21268) );
  AOI22_X1 U9920 ( .A1(\mem[604][6] ), .A2(n14723), .B1(n26526), .B2(
        data_in[6]), .ZN(n14729) );
  INV_X1 U9921 ( .A(n14730), .ZN(n21267) );
  AOI22_X1 U9922 ( .A1(\mem[604][7] ), .A2(n14723), .B1(n26526), .B2(
        data_in[7]), .ZN(n14730) );
  INV_X1 U9923 ( .A(n14731), .ZN(n21266) );
  AOI22_X1 U9924 ( .A1(\mem[605][0] ), .A2(n14732), .B1(n26525), .B2(
        data_in[0]), .ZN(n14731) );
  INV_X1 U9925 ( .A(n14733), .ZN(n21265) );
  AOI22_X1 U9926 ( .A1(\mem[605][1] ), .A2(n14732), .B1(n26525), .B2(
        data_in[1]), .ZN(n14733) );
  INV_X1 U9927 ( .A(n14734), .ZN(n21264) );
  AOI22_X1 U9928 ( .A1(\mem[605][2] ), .A2(n14732), .B1(n26525), .B2(
        data_in[2]), .ZN(n14734) );
  INV_X1 U9929 ( .A(n14735), .ZN(n21263) );
  AOI22_X1 U9930 ( .A1(\mem[605][3] ), .A2(n14732), .B1(n26525), .B2(
        data_in[3]), .ZN(n14735) );
  INV_X1 U9931 ( .A(n14736), .ZN(n21262) );
  AOI22_X1 U9932 ( .A1(\mem[605][4] ), .A2(n14732), .B1(n26525), .B2(
        data_in[4]), .ZN(n14736) );
  INV_X1 U9933 ( .A(n14737), .ZN(n21261) );
  AOI22_X1 U9934 ( .A1(\mem[605][5] ), .A2(n14732), .B1(n26525), .B2(
        data_in[5]), .ZN(n14737) );
  INV_X1 U9935 ( .A(n14738), .ZN(n21260) );
  AOI22_X1 U9936 ( .A1(\mem[605][6] ), .A2(n14732), .B1(n26525), .B2(
        data_in[6]), .ZN(n14738) );
  INV_X1 U9937 ( .A(n14739), .ZN(n21259) );
  AOI22_X1 U9938 ( .A1(\mem[605][7] ), .A2(n14732), .B1(n26525), .B2(
        data_in[7]), .ZN(n14739) );
  INV_X1 U9939 ( .A(n14740), .ZN(n21258) );
  AOI22_X1 U9940 ( .A1(\mem[606][0] ), .A2(n14741), .B1(n26524), .B2(
        data_in[0]), .ZN(n14740) );
  INV_X1 U9941 ( .A(n14742), .ZN(n21257) );
  AOI22_X1 U9942 ( .A1(\mem[606][1] ), .A2(n14741), .B1(n26524), .B2(
        data_in[1]), .ZN(n14742) );
  INV_X1 U9943 ( .A(n14743), .ZN(n21256) );
  AOI22_X1 U9944 ( .A1(\mem[606][2] ), .A2(n14741), .B1(n26524), .B2(
        data_in[2]), .ZN(n14743) );
  INV_X1 U9945 ( .A(n14744), .ZN(n21255) );
  AOI22_X1 U9946 ( .A1(\mem[606][3] ), .A2(n14741), .B1(n26524), .B2(
        data_in[3]), .ZN(n14744) );
  INV_X1 U9947 ( .A(n14745), .ZN(n21254) );
  AOI22_X1 U9948 ( .A1(\mem[606][4] ), .A2(n14741), .B1(n26524), .B2(
        data_in[4]), .ZN(n14745) );
  INV_X1 U9949 ( .A(n14746), .ZN(n21253) );
  AOI22_X1 U9950 ( .A1(\mem[606][5] ), .A2(n14741), .B1(n26524), .B2(
        data_in[5]), .ZN(n14746) );
  INV_X1 U9951 ( .A(n14747), .ZN(n21252) );
  AOI22_X1 U9952 ( .A1(\mem[606][6] ), .A2(n14741), .B1(n26524), .B2(
        data_in[6]), .ZN(n14747) );
  INV_X1 U9953 ( .A(n14748), .ZN(n21251) );
  AOI22_X1 U9954 ( .A1(\mem[606][7] ), .A2(n14741), .B1(n26524), .B2(
        data_in[7]), .ZN(n14748) );
  INV_X1 U9955 ( .A(n14749), .ZN(n21250) );
  AOI22_X1 U9956 ( .A1(\mem[607][0] ), .A2(n14750), .B1(n26523), .B2(
        data_in[0]), .ZN(n14749) );
  INV_X1 U9957 ( .A(n14751), .ZN(n21249) );
  AOI22_X1 U9958 ( .A1(\mem[607][1] ), .A2(n14750), .B1(n26523), .B2(
        data_in[1]), .ZN(n14751) );
  INV_X1 U9959 ( .A(n14752), .ZN(n21248) );
  AOI22_X1 U9960 ( .A1(\mem[607][2] ), .A2(n14750), .B1(n26523), .B2(
        data_in[2]), .ZN(n14752) );
  INV_X1 U9961 ( .A(n14753), .ZN(n21247) );
  AOI22_X1 U9962 ( .A1(\mem[607][3] ), .A2(n14750), .B1(n26523), .B2(
        data_in[3]), .ZN(n14753) );
  INV_X1 U9963 ( .A(n14754), .ZN(n21246) );
  AOI22_X1 U9964 ( .A1(\mem[607][4] ), .A2(n14750), .B1(n26523), .B2(
        data_in[4]), .ZN(n14754) );
  INV_X1 U9965 ( .A(n14755), .ZN(n21245) );
  AOI22_X1 U9966 ( .A1(\mem[607][5] ), .A2(n14750), .B1(n26523), .B2(
        data_in[5]), .ZN(n14755) );
  INV_X1 U9967 ( .A(n14756), .ZN(n21244) );
  AOI22_X1 U9968 ( .A1(\mem[607][6] ), .A2(n14750), .B1(n26523), .B2(
        data_in[6]), .ZN(n14756) );
  INV_X1 U9969 ( .A(n14757), .ZN(n21243) );
  AOI22_X1 U9970 ( .A1(\mem[607][7] ), .A2(n14750), .B1(n26523), .B2(
        data_in[7]), .ZN(n14757) );
  INV_X1 U9971 ( .A(n14831), .ZN(n21178) );
  AOI22_X1 U9972 ( .A1(\mem[616][0] ), .A2(n14832), .B1(n26514), .B2(
        data_in[0]), .ZN(n14831) );
  INV_X1 U9973 ( .A(n14833), .ZN(n21177) );
  AOI22_X1 U9974 ( .A1(\mem[616][1] ), .A2(n14832), .B1(n26514), .B2(
        data_in[1]), .ZN(n14833) );
  INV_X1 U9975 ( .A(n14834), .ZN(n21176) );
  AOI22_X1 U9976 ( .A1(\mem[616][2] ), .A2(n14832), .B1(n26514), .B2(
        data_in[2]), .ZN(n14834) );
  INV_X1 U9977 ( .A(n14835), .ZN(n21175) );
  AOI22_X1 U9978 ( .A1(\mem[616][3] ), .A2(n14832), .B1(n26514), .B2(
        data_in[3]), .ZN(n14835) );
  INV_X1 U9979 ( .A(n14836), .ZN(n21174) );
  AOI22_X1 U9980 ( .A1(\mem[616][4] ), .A2(n14832), .B1(n26514), .B2(
        data_in[4]), .ZN(n14836) );
  INV_X1 U9981 ( .A(n14837), .ZN(n21173) );
  AOI22_X1 U9982 ( .A1(\mem[616][5] ), .A2(n14832), .B1(n26514), .B2(
        data_in[5]), .ZN(n14837) );
  INV_X1 U9983 ( .A(n14838), .ZN(n21172) );
  AOI22_X1 U9984 ( .A1(\mem[616][6] ), .A2(n14832), .B1(n26514), .B2(
        data_in[6]), .ZN(n14838) );
  INV_X1 U9985 ( .A(n14839), .ZN(n21171) );
  AOI22_X1 U9986 ( .A1(\mem[616][7] ), .A2(n14832), .B1(n26514), .B2(
        data_in[7]), .ZN(n14839) );
  INV_X1 U9987 ( .A(n14840), .ZN(n21170) );
  AOI22_X1 U9988 ( .A1(\mem[617][0] ), .A2(n14841), .B1(n26513), .B2(
        data_in[0]), .ZN(n14840) );
  INV_X1 U9989 ( .A(n14842), .ZN(n21169) );
  AOI22_X1 U9990 ( .A1(\mem[617][1] ), .A2(n14841), .B1(n26513), .B2(
        data_in[1]), .ZN(n14842) );
  INV_X1 U9991 ( .A(n14843), .ZN(n21168) );
  AOI22_X1 U9992 ( .A1(\mem[617][2] ), .A2(n14841), .B1(n26513), .B2(
        data_in[2]), .ZN(n14843) );
  INV_X1 U9993 ( .A(n14844), .ZN(n21167) );
  AOI22_X1 U9994 ( .A1(\mem[617][3] ), .A2(n14841), .B1(n26513), .B2(
        data_in[3]), .ZN(n14844) );
  INV_X1 U9995 ( .A(n14845), .ZN(n21166) );
  AOI22_X1 U9996 ( .A1(\mem[617][4] ), .A2(n14841), .B1(n26513), .B2(
        data_in[4]), .ZN(n14845) );
  INV_X1 U9997 ( .A(n14846), .ZN(n21165) );
  AOI22_X1 U9998 ( .A1(\mem[617][5] ), .A2(n14841), .B1(n26513), .B2(
        data_in[5]), .ZN(n14846) );
  INV_X1 U9999 ( .A(n14847), .ZN(n21164) );
  AOI22_X1 U10000 ( .A1(\mem[617][6] ), .A2(n14841), .B1(n26513), .B2(
        data_in[6]), .ZN(n14847) );
  INV_X1 U10001 ( .A(n14848), .ZN(n21163) );
  AOI22_X1 U10002 ( .A1(\mem[617][7] ), .A2(n14841), .B1(n26513), .B2(
        data_in[7]), .ZN(n14848) );
  INV_X1 U10003 ( .A(n14849), .ZN(n21162) );
  AOI22_X1 U10004 ( .A1(\mem[618][0] ), .A2(n14850), .B1(n26512), .B2(
        data_in[0]), .ZN(n14849) );
  INV_X1 U10005 ( .A(n14851), .ZN(n21161) );
  AOI22_X1 U10006 ( .A1(\mem[618][1] ), .A2(n14850), .B1(n26512), .B2(
        data_in[1]), .ZN(n14851) );
  INV_X1 U10007 ( .A(n14852), .ZN(n21160) );
  AOI22_X1 U10008 ( .A1(\mem[618][2] ), .A2(n14850), .B1(n26512), .B2(
        data_in[2]), .ZN(n14852) );
  INV_X1 U10009 ( .A(n14853), .ZN(n21159) );
  AOI22_X1 U10010 ( .A1(\mem[618][3] ), .A2(n14850), .B1(n26512), .B2(
        data_in[3]), .ZN(n14853) );
  INV_X1 U10011 ( .A(n14854), .ZN(n21158) );
  AOI22_X1 U10012 ( .A1(\mem[618][4] ), .A2(n14850), .B1(n26512), .B2(
        data_in[4]), .ZN(n14854) );
  INV_X1 U10013 ( .A(n14855), .ZN(n21157) );
  AOI22_X1 U10014 ( .A1(\mem[618][5] ), .A2(n14850), .B1(n26512), .B2(
        data_in[5]), .ZN(n14855) );
  INV_X1 U10015 ( .A(n14856), .ZN(n21156) );
  AOI22_X1 U10016 ( .A1(\mem[618][6] ), .A2(n14850), .B1(n26512), .B2(
        data_in[6]), .ZN(n14856) );
  INV_X1 U10017 ( .A(n14857), .ZN(n21155) );
  AOI22_X1 U10018 ( .A1(\mem[618][7] ), .A2(n14850), .B1(n26512), .B2(
        data_in[7]), .ZN(n14857) );
  INV_X1 U10019 ( .A(n14858), .ZN(n21154) );
  AOI22_X1 U10020 ( .A1(\mem[619][0] ), .A2(n14859), .B1(n26511), .B2(
        data_in[0]), .ZN(n14858) );
  INV_X1 U10021 ( .A(n14860), .ZN(n21153) );
  AOI22_X1 U10022 ( .A1(\mem[619][1] ), .A2(n14859), .B1(n26511), .B2(
        data_in[1]), .ZN(n14860) );
  INV_X1 U10023 ( .A(n14861), .ZN(n21152) );
  AOI22_X1 U10024 ( .A1(\mem[619][2] ), .A2(n14859), .B1(n26511), .B2(
        data_in[2]), .ZN(n14861) );
  INV_X1 U10025 ( .A(n14862), .ZN(n21151) );
  AOI22_X1 U10026 ( .A1(\mem[619][3] ), .A2(n14859), .B1(n26511), .B2(
        data_in[3]), .ZN(n14862) );
  INV_X1 U10027 ( .A(n14863), .ZN(n21150) );
  AOI22_X1 U10028 ( .A1(\mem[619][4] ), .A2(n14859), .B1(n26511), .B2(
        data_in[4]), .ZN(n14863) );
  INV_X1 U10029 ( .A(n14864), .ZN(n21149) );
  AOI22_X1 U10030 ( .A1(\mem[619][5] ), .A2(n14859), .B1(n26511), .B2(
        data_in[5]), .ZN(n14864) );
  INV_X1 U10031 ( .A(n14865), .ZN(n21148) );
  AOI22_X1 U10032 ( .A1(\mem[619][6] ), .A2(n14859), .B1(n26511), .B2(
        data_in[6]), .ZN(n14865) );
  INV_X1 U10033 ( .A(n14866), .ZN(n21147) );
  AOI22_X1 U10034 ( .A1(\mem[619][7] ), .A2(n14859), .B1(n26511), .B2(
        data_in[7]), .ZN(n14866) );
  INV_X1 U10035 ( .A(n14867), .ZN(n21146) );
  AOI22_X1 U10036 ( .A1(\mem[620][0] ), .A2(n14868), .B1(n26510), .B2(
        data_in[0]), .ZN(n14867) );
  INV_X1 U10037 ( .A(n14869), .ZN(n21145) );
  AOI22_X1 U10038 ( .A1(\mem[620][1] ), .A2(n14868), .B1(n26510), .B2(
        data_in[1]), .ZN(n14869) );
  INV_X1 U10039 ( .A(n14870), .ZN(n21144) );
  AOI22_X1 U10040 ( .A1(\mem[620][2] ), .A2(n14868), .B1(n26510), .B2(
        data_in[2]), .ZN(n14870) );
  INV_X1 U10041 ( .A(n14871), .ZN(n21143) );
  AOI22_X1 U10042 ( .A1(\mem[620][3] ), .A2(n14868), .B1(n26510), .B2(
        data_in[3]), .ZN(n14871) );
  INV_X1 U10043 ( .A(n14872), .ZN(n21142) );
  AOI22_X1 U10044 ( .A1(\mem[620][4] ), .A2(n14868), .B1(n26510), .B2(
        data_in[4]), .ZN(n14872) );
  INV_X1 U10045 ( .A(n14873), .ZN(n21141) );
  AOI22_X1 U10046 ( .A1(\mem[620][5] ), .A2(n14868), .B1(n26510), .B2(
        data_in[5]), .ZN(n14873) );
  INV_X1 U10047 ( .A(n14874), .ZN(n21140) );
  AOI22_X1 U10048 ( .A1(\mem[620][6] ), .A2(n14868), .B1(n26510), .B2(
        data_in[6]), .ZN(n14874) );
  INV_X1 U10049 ( .A(n14875), .ZN(n21139) );
  AOI22_X1 U10050 ( .A1(\mem[620][7] ), .A2(n14868), .B1(n26510), .B2(
        data_in[7]), .ZN(n14875) );
  INV_X1 U10051 ( .A(n14876), .ZN(n21138) );
  AOI22_X1 U10052 ( .A1(\mem[621][0] ), .A2(n14877), .B1(n26509), .B2(
        data_in[0]), .ZN(n14876) );
  INV_X1 U10053 ( .A(n14878), .ZN(n21137) );
  AOI22_X1 U10054 ( .A1(\mem[621][1] ), .A2(n14877), .B1(n26509), .B2(
        data_in[1]), .ZN(n14878) );
  INV_X1 U10055 ( .A(n14879), .ZN(n21136) );
  AOI22_X1 U10056 ( .A1(\mem[621][2] ), .A2(n14877), .B1(n26509), .B2(
        data_in[2]), .ZN(n14879) );
  INV_X1 U10057 ( .A(n14880), .ZN(n21135) );
  AOI22_X1 U10058 ( .A1(\mem[621][3] ), .A2(n14877), .B1(n26509), .B2(
        data_in[3]), .ZN(n14880) );
  INV_X1 U10059 ( .A(n14881), .ZN(n21134) );
  AOI22_X1 U10060 ( .A1(\mem[621][4] ), .A2(n14877), .B1(n26509), .B2(
        data_in[4]), .ZN(n14881) );
  INV_X1 U10061 ( .A(n14882), .ZN(n21133) );
  AOI22_X1 U10062 ( .A1(\mem[621][5] ), .A2(n14877), .B1(n26509), .B2(
        data_in[5]), .ZN(n14882) );
  INV_X1 U10063 ( .A(n14883), .ZN(n21132) );
  AOI22_X1 U10064 ( .A1(\mem[621][6] ), .A2(n14877), .B1(n26509), .B2(
        data_in[6]), .ZN(n14883) );
  INV_X1 U10065 ( .A(n14884), .ZN(n21131) );
  AOI22_X1 U10066 ( .A1(\mem[621][7] ), .A2(n14877), .B1(n26509), .B2(
        data_in[7]), .ZN(n14884) );
  INV_X1 U10067 ( .A(n14885), .ZN(n21130) );
  AOI22_X1 U10068 ( .A1(\mem[622][0] ), .A2(n14886), .B1(n26508), .B2(
        data_in[0]), .ZN(n14885) );
  INV_X1 U10069 ( .A(n14887), .ZN(n21129) );
  AOI22_X1 U10070 ( .A1(\mem[622][1] ), .A2(n14886), .B1(n26508), .B2(
        data_in[1]), .ZN(n14887) );
  INV_X1 U10071 ( .A(n14888), .ZN(n21128) );
  AOI22_X1 U10072 ( .A1(\mem[622][2] ), .A2(n14886), .B1(n26508), .B2(
        data_in[2]), .ZN(n14888) );
  INV_X1 U10073 ( .A(n14889), .ZN(n21127) );
  AOI22_X1 U10074 ( .A1(\mem[622][3] ), .A2(n14886), .B1(n26508), .B2(
        data_in[3]), .ZN(n14889) );
  INV_X1 U10075 ( .A(n14890), .ZN(n21126) );
  AOI22_X1 U10076 ( .A1(\mem[622][4] ), .A2(n14886), .B1(n26508), .B2(
        data_in[4]), .ZN(n14890) );
  INV_X1 U10077 ( .A(n14891), .ZN(n21125) );
  AOI22_X1 U10078 ( .A1(\mem[622][5] ), .A2(n14886), .B1(n26508), .B2(
        data_in[5]), .ZN(n14891) );
  INV_X1 U10079 ( .A(n14892), .ZN(n21124) );
  AOI22_X1 U10080 ( .A1(\mem[622][6] ), .A2(n14886), .B1(n26508), .B2(
        data_in[6]), .ZN(n14892) );
  INV_X1 U10081 ( .A(n14893), .ZN(n21123) );
  AOI22_X1 U10082 ( .A1(\mem[622][7] ), .A2(n14886), .B1(n26508), .B2(
        data_in[7]), .ZN(n14893) );
  INV_X1 U10083 ( .A(n14894), .ZN(n21122) );
  AOI22_X1 U10084 ( .A1(\mem[623][0] ), .A2(n14895), .B1(n26507), .B2(
        data_in[0]), .ZN(n14894) );
  INV_X1 U10085 ( .A(n14896), .ZN(n21121) );
  AOI22_X1 U10086 ( .A1(\mem[623][1] ), .A2(n14895), .B1(n26507), .B2(
        data_in[1]), .ZN(n14896) );
  INV_X1 U10087 ( .A(n14897), .ZN(n21120) );
  AOI22_X1 U10088 ( .A1(\mem[623][2] ), .A2(n14895), .B1(n26507), .B2(
        data_in[2]), .ZN(n14897) );
  INV_X1 U10089 ( .A(n14898), .ZN(n21119) );
  AOI22_X1 U10090 ( .A1(\mem[623][3] ), .A2(n14895), .B1(n26507), .B2(
        data_in[3]), .ZN(n14898) );
  INV_X1 U10091 ( .A(n14899), .ZN(n21118) );
  AOI22_X1 U10092 ( .A1(\mem[623][4] ), .A2(n14895), .B1(n26507), .B2(
        data_in[4]), .ZN(n14899) );
  INV_X1 U10093 ( .A(n14900), .ZN(n21117) );
  AOI22_X1 U10094 ( .A1(\mem[623][5] ), .A2(n14895), .B1(n26507), .B2(
        data_in[5]), .ZN(n14900) );
  INV_X1 U10095 ( .A(n14901), .ZN(n21116) );
  AOI22_X1 U10096 ( .A1(\mem[623][6] ), .A2(n14895), .B1(n26507), .B2(
        data_in[6]), .ZN(n14901) );
  INV_X1 U10097 ( .A(n14902), .ZN(n21115) );
  AOI22_X1 U10098 ( .A1(\mem[623][7] ), .A2(n14895), .B1(n26507), .B2(
        data_in[7]), .ZN(n14902) );
  INV_X1 U10099 ( .A(n14903), .ZN(n21114) );
  AOI22_X1 U10100 ( .A1(\mem[624][0] ), .A2(n14904), .B1(n26506), .B2(
        data_in[0]), .ZN(n14903) );
  INV_X1 U10101 ( .A(n14905), .ZN(n21113) );
  AOI22_X1 U10102 ( .A1(\mem[624][1] ), .A2(n14904), .B1(n26506), .B2(
        data_in[1]), .ZN(n14905) );
  INV_X1 U10103 ( .A(n14906), .ZN(n21112) );
  AOI22_X1 U10104 ( .A1(\mem[624][2] ), .A2(n14904), .B1(n26506), .B2(
        data_in[2]), .ZN(n14906) );
  INV_X1 U10105 ( .A(n14907), .ZN(n21111) );
  AOI22_X1 U10106 ( .A1(\mem[624][3] ), .A2(n14904), .B1(n26506), .B2(
        data_in[3]), .ZN(n14907) );
  INV_X1 U10107 ( .A(n14908), .ZN(n21110) );
  AOI22_X1 U10108 ( .A1(\mem[624][4] ), .A2(n14904), .B1(n26506), .B2(
        data_in[4]), .ZN(n14908) );
  INV_X1 U10109 ( .A(n14909), .ZN(n21109) );
  AOI22_X1 U10110 ( .A1(\mem[624][5] ), .A2(n14904), .B1(n26506), .B2(
        data_in[5]), .ZN(n14909) );
  INV_X1 U10111 ( .A(n14910), .ZN(n21108) );
  AOI22_X1 U10112 ( .A1(\mem[624][6] ), .A2(n14904), .B1(n26506), .B2(
        data_in[6]), .ZN(n14910) );
  INV_X1 U10113 ( .A(n14911), .ZN(n21107) );
  AOI22_X1 U10114 ( .A1(\mem[624][7] ), .A2(n14904), .B1(n26506), .B2(
        data_in[7]), .ZN(n14911) );
  INV_X1 U10115 ( .A(n14912), .ZN(n21106) );
  AOI22_X1 U10116 ( .A1(\mem[625][0] ), .A2(n14913), .B1(n26505), .B2(
        data_in[0]), .ZN(n14912) );
  INV_X1 U10117 ( .A(n14914), .ZN(n21105) );
  AOI22_X1 U10118 ( .A1(\mem[625][1] ), .A2(n14913), .B1(n26505), .B2(
        data_in[1]), .ZN(n14914) );
  INV_X1 U10119 ( .A(n14915), .ZN(n21104) );
  AOI22_X1 U10120 ( .A1(\mem[625][2] ), .A2(n14913), .B1(n26505), .B2(
        data_in[2]), .ZN(n14915) );
  INV_X1 U10121 ( .A(n14916), .ZN(n21103) );
  AOI22_X1 U10122 ( .A1(\mem[625][3] ), .A2(n14913), .B1(n26505), .B2(
        data_in[3]), .ZN(n14916) );
  INV_X1 U10123 ( .A(n14917), .ZN(n21102) );
  AOI22_X1 U10124 ( .A1(\mem[625][4] ), .A2(n14913), .B1(n26505), .B2(
        data_in[4]), .ZN(n14917) );
  INV_X1 U10125 ( .A(n14918), .ZN(n21101) );
  AOI22_X1 U10126 ( .A1(\mem[625][5] ), .A2(n14913), .B1(n26505), .B2(
        data_in[5]), .ZN(n14918) );
  INV_X1 U10127 ( .A(n14919), .ZN(n21100) );
  AOI22_X1 U10128 ( .A1(\mem[625][6] ), .A2(n14913), .B1(n26505), .B2(
        data_in[6]), .ZN(n14919) );
  INV_X1 U10129 ( .A(n14920), .ZN(n21099) );
  AOI22_X1 U10130 ( .A1(\mem[625][7] ), .A2(n14913), .B1(n26505), .B2(
        data_in[7]), .ZN(n14920) );
  INV_X1 U10131 ( .A(n14921), .ZN(n21098) );
  AOI22_X1 U10132 ( .A1(\mem[626][0] ), .A2(n14922), .B1(n26504), .B2(
        data_in[0]), .ZN(n14921) );
  INV_X1 U10133 ( .A(n14923), .ZN(n21097) );
  AOI22_X1 U10134 ( .A1(\mem[626][1] ), .A2(n14922), .B1(n26504), .B2(
        data_in[1]), .ZN(n14923) );
  INV_X1 U10135 ( .A(n14924), .ZN(n21096) );
  AOI22_X1 U10136 ( .A1(\mem[626][2] ), .A2(n14922), .B1(n26504), .B2(
        data_in[2]), .ZN(n14924) );
  INV_X1 U10137 ( .A(n14925), .ZN(n21095) );
  AOI22_X1 U10138 ( .A1(\mem[626][3] ), .A2(n14922), .B1(n26504), .B2(
        data_in[3]), .ZN(n14925) );
  INV_X1 U10139 ( .A(n14926), .ZN(n21094) );
  AOI22_X1 U10140 ( .A1(\mem[626][4] ), .A2(n14922), .B1(n26504), .B2(
        data_in[4]), .ZN(n14926) );
  INV_X1 U10141 ( .A(n14927), .ZN(n21093) );
  AOI22_X1 U10142 ( .A1(\mem[626][5] ), .A2(n14922), .B1(n26504), .B2(
        data_in[5]), .ZN(n14927) );
  INV_X1 U10143 ( .A(n14928), .ZN(n21092) );
  AOI22_X1 U10144 ( .A1(\mem[626][6] ), .A2(n14922), .B1(n26504), .B2(
        data_in[6]), .ZN(n14928) );
  INV_X1 U10145 ( .A(n14929), .ZN(n21091) );
  AOI22_X1 U10146 ( .A1(\mem[626][7] ), .A2(n14922), .B1(n26504), .B2(
        data_in[7]), .ZN(n14929) );
  INV_X1 U10147 ( .A(n14930), .ZN(n21090) );
  AOI22_X1 U10148 ( .A1(\mem[627][0] ), .A2(n14931), .B1(n26503), .B2(
        data_in[0]), .ZN(n14930) );
  INV_X1 U10149 ( .A(n14932), .ZN(n21089) );
  AOI22_X1 U10150 ( .A1(\mem[627][1] ), .A2(n14931), .B1(n26503), .B2(
        data_in[1]), .ZN(n14932) );
  INV_X1 U10151 ( .A(n14933), .ZN(n21088) );
  AOI22_X1 U10152 ( .A1(\mem[627][2] ), .A2(n14931), .B1(n26503), .B2(
        data_in[2]), .ZN(n14933) );
  INV_X1 U10153 ( .A(n14934), .ZN(n21087) );
  AOI22_X1 U10154 ( .A1(\mem[627][3] ), .A2(n14931), .B1(n26503), .B2(
        data_in[3]), .ZN(n14934) );
  INV_X1 U10155 ( .A(n14935), .ZN(n21086) );
  AOI22_X1 U10156 ( .A1(\mem[627][4] ), .A2(n14931), .B1(n26503), .B2(
        data_in[4]), .ZN(n14935) );
  INV_X1 U10157 ( .A(n14936), .ZN(n21085) );
  AOI22_X1 U10158 ( .A1(\mem[627][5] ), .A2(n14931), .B1(n26503), .B2(
        data_in[5]), .ZN(n14936) );
  INV_X1 U10159 ( .A(n14937), .ZN(n21084) );
  AOI22_X1 U10160 ( .A1(\mem[627][6] ), .A2(n14931), .B1(n26503), .B2(
        data_in[6]), .ZN(n14937) );
  INV_X1 U10161 ( .A(n14938), .ZN(n21083) );
  AOI22_X1 U10162 ( .A1(\mem[627][7] ), .A2(n14931), .B1(n26503), .B2(
        data_in[7]), .ZN(n14938) );
  INV_X1 U10163 ( .A(n14939), .ZN(n21082) );
  AOI22_X1 U10164 ( .A1(\mem[628][0] ), .A2(n14940), .B1(n26502), .B2(
        data_in[0]), .ZN(n14939) );
  INV_X1 U10165 ( .A(n14941), .ZN(n21081) );
  AOI22_X1 U10166 ( .A1(\mem[628][1] ), .A2(n14940), .B1(n26502), .B2(
        data_in[1]), .ZN(n14941) );
  INV_X1 U10167 ( .A(n14942), .ZN(n21080) );
  AOI22_X1 U10168 ( .A1(\mem[628][2] ), .A2(n14940), .B1(n26502), .B2(
        data_in[2]), .ZN(n14942) );
  INV_X1 U10169 ( .A(n14943), .ZN(n21079) );
  AOI22_X1 U10170 ( .A1(\mem[628][3] ), .A2(n14940), .B1(n26502), .B2(
        data_in[3]), .ZN(n14943) );
  INV_X1 U10171 ( .A(n14944), .ZN(n21078) );
  AOI22_X1 U10172 ( .A1(\mem[628][4] ), .A2(n14940), .B1(n26502), .B2(
        data_in[4]), .ZN(n14944) );
  INV_X1 U10173 ( .A(n14945), .ZN(n21077) );
  AOI22_X1 U10174 ( .A1(\mem[628][5] ), .A2(n14940), .B1(n26502), .B2(
        data_in[5]), .ZN(n14945) );
  INV_X1 U10175 ( .A(n14946), .ZN(n21076) );
  AOI22_X1 U10176 ( .A1(\mem[628][6] ), .A2(n14940), .B1(n26502), .B2(
        data_in[6]), .ZN(n14946) );
  INV_X1 U10177 ( .A(n14947), .ZN(n21075) );
  AOI22_X1 U10178 ( .A1(\mem[628][7] ), .A2(n14940), .B1(n26502), .B2(
        data_in[7]), .ZN(n14947) );
  INV_X1 U10179 ( .A(n14948), .ZN(n21074) );
  AOI22_X1 U10180 ( .A1(\mem[629][0] ), .A2(n14949), .B1(n26501), .B2(
        data_in[0]), .ZN(n14948) );
  INV_X1 U10181 ( .A(n14950), .ZN(n21073) );
  AOI22_X1 U10182 ( .A1(\mem[629][1] ), .A2(n14949), .B1(n26501), .B2(
        data_in[1]), .ZN(n14950) );
  INV_X1 U10183 ( .A(n14951), .ZN(n21072) );
  AOI22_X1 U10184 ( .A1(\mem[629][2] ), .A2(n14949), .B1(n26501), .B2(
        data_in[2]), .ZN(n14951) );
  INV_X1 U10185 ( .A(n14952), .ZN(n21071) );
  AOI22_X1 U10186 ( .A1(\mem[629][3] ), .A2(n14949), .B1(n26501), .B2(
        data_in[3]), .ZN(n14952) );
  INV_X1 U10187 ( .A(n14953), .ZN(n21070) );
  AOI22_X1 U10188 ( .A1(\mem[629][4] ), .A2(n14949), .B1(n26501), .B2(
        data_in[4]), .ZN(n14953) );
  INV_X1 U10189 ( .A(n14954), .ZN(n21069) );
  AOI22_X1 U10190 ( .A1(\mem[629][5] ), .A2(n14949), .B1(n26501), .B2(
        data_in[5]), .ZN(n14954) );
  INV_X1 U10191 ( .A(n14955), .ZN(n21068) );
  AOI22_X1 U10192 ( .A1(\mem[629][6] ), .A2(n14949), .B1(n26501), .B2(
        data_in[6]), .ZN(n14955) );
  INV_X1 U10193 ( .A(n14956), .ZN(n21067) );
  AOI22_X1 U10194 ( .A1(\mem[629][7] ), .A2(n14949), .B1(n26501), .B2(
        data_in[7]), .ZN(n14956) );
  INV_X1 U10195 ( .A(n14957), .ZN(n21066) );
  AOI22_X1 U10196 ( .A1(\mem[630][0] ), .A2(n14958), .B1(n26500), .B2(
        data_in[0]), .ZN(n14957) );
  INV_X1 U10197 ( .A(n14959), .ZN(n21065) );
  AOI22_X1 U10198 ( .A1(\mem[630][1] ), .A2(n14958), .B1(n26500), .B2(
        data_in[1]), .ZN(n14959) );
  INV_X1 U10199 ( .A(n14960), .ZN(n21064) );
  AOI22_X1 U10200 ( .A1(\mem[630][2] ), .A2(n14958), .B1(n26500), .B2(
        data_in[2]), .ZN(n14960) );
  INV_X1 U10201 ( .A(n14961), .ZN(n21063) );
  AOI22_X1 U10202 ( .A1(\mem[630][3] ), .A2(n14958), .B1(n26500), .B2(
        data_in[3]), .ZN(n14961) );
  INV_X1 U10203 ( .A(n14962), .ZN(n21062) );
  AOI22_X1 U10204 ( .A1(\mem[630][4] ), .A2(n14958), .B1(n26500), .B2(
        data_in[4]), .ZN(n14962) );
  INV_X1 U10205 ( .A(n14963), .ZN(n21061) );
  AOI22_X1 U10206 ( .A1(\mem[630][5] ), .A2(n14958), .B1(n26500), .B2(
        data_in[5]), .ZN(n14963) );
  INV_X1 U10207 ( .A(n14964), .ZN(n21060) );
  AOI22_X1 U10208 ( .A1(\mem[630][6] ), .A2(n14958), .B1(n26500), .B2(
        data_in[6]), .ZN(n14964) );
  INV_X1 U10209 ( .A(n14965), .ZN(n21059) );
  AOI22_X1 U10210 ( .A1(\mem[630][7] ), .A2(n14958), .B1(n26500), .B2(
        data_in[7]), .ZN(n14965) );
  INV_X1 U10211 ( .A(n14966), .ZN(n21058) );
  AOI22_X1 U10212 ( .A1(\mem[631][0] ), .A2(n14967), .B1(n26499), .B2(
        data_in[0]), .ZN(n14966) );
  INV_X1 U10213 ( .A(n14968), .ZN(n21057) );
  AOI22_X1 U10214 ( .A1(\mem[631][1] ), .A2(n14967), .B1(n26499), .B2(
        data_in[1]), .ZN(n14968) );
  INV_X1 U10215 ( .A(n14969), .ZN(n21056) );
  AOI22_X1 U10216 ( .A1(\mem[631][2] ), .A2(n14967), .B1(n26499), .B2(
        data_in[2]), .ZN(n14969) );
  INV_X1 U10217 ( .A(n14970), .ZN(n21055) );
  AOI22_X1 U10218 ( .A1(\mem[631][3] ), .A2(n14967), .B1(n26499), .B2(
        data_in[3]), .ZN(n14970) );
  INV_X1 U10219 ( .A(n14971), .ZN(n21054) );
  AOI22_X1 U10220 ( .A1(\mem[631][4] ), .A2(n14967), .B1(n26499), .B2(
        data_in[4]), .ZN(n14971) );
  INV_X1 U10221 ( .A(n14972), .ZN(n21053) );
  AOI22_X1 U10222 ( .A1(\mem[631][5] ), .A2(n14967), .B1(n26499), .B2(
        data_in[5]), .ZN(n14972) );
  INV_X1 U10223 ( .A(n14973), .ZN(n21052) );
  AOI22_X1 U10224 ( .A1(\mem[631][6] ), .A2(n14967), .B1(n26499), .B2(
        data_in[6]), .ZN(n14973) );
  INV_X1 U10225 ( .A(n14974), .ZN(n21051) );
  AOI22_X1 U10226 ( .A1(\mem[631][7] ), .A2(n14967), .B1(n26499), .B2(
        data_in[7]), .ZN(n14974) );
  INV_X1 U10227 ( .A(n14975), .ZN(n21050) );
  AOI22_X1 U10228 ( .A1(\mem[632][0] ), .A2(n14976), .B1(n26498), .B2(
        data_in[0]), .ZN(n14975) );
  INV_X1 U10229 ( .A(n14977), .ZN(n21049) );
  AOI22_X1 U10230 ( .A1(\mem[632][1] ), .A2(n14976), .B1(n26498), .B2(
        data_in[1]), .ZN(n14977) );
  INV_X1 U10231 ( .A(n14978), .ZN(n21048) );
  AOI22_X1 U10232 ( .A1(\mem[632][2] ), .A2(n14976), .B1(n26498), .B2(
        data_in[2]), .ZN(n14978) );
  INV_X1 U10233 ( .A(n14979), .ZN(n21047) );
  AOI22_X1 U10234 ( .A1(\mem[632][3] ), .A2(n14976), .B1(n26498), .B2(
        data_in[3]), .ZN(n14979) );
  INV_X1 U10235 ( .A(n14980), .ZN(n21046) );
  AOI22_X1 U10236 ( .A1(\mem[632][4] ), .A2(n14976), .B1(n26498), .B2(
        data_in[4]), .ZN(n14980) );
  INV_X1 U10237 ( .A(n14981), .ZN(n21045) );
  AOI22_X1 U10238 ( .A1(\mem[632][5] ), .A2(n14976), .B1(n26498), .B2(
        data_in[5]), .ZN(n14981) );
  INV_X1 U10239 ( .A(n14982), .ZN(n21044) );
  AOI22_X1 U10240 ( .A1(\mem[632][6] ), .A2(n14976), .B1(n26498), .B2(
        data_in[6]), .ZN(n14982) );
  INV_X1 U10241 ( .A(n14983), .ZN(n21043) );
  AOI22_X1 U10242 ( .A1(\mem[632][7] ), .A2(n14976), .B1(n26498), .B2(
        data_in[7]), .ZN(n14983) );
  INV_X1 U10243 ( .A(n14984), .ZN(n21042) );
  AOI22_X1 U10244 ( .A1(\mem[633][0] ), .A2(n14985), .B1(n26497), .B2(
        data_in[0]), .ZN(n14984) );
  INV_X1 U10245 ( .A(n14986), .ZN(n21041) );
  AOI22_X1 U10246 ( .A1(\mem[633][1] ), .A2(n14985), .B1(n26497), .B2(
        data_in[1]), .ZN(n14986) );
  INV_X1 U10247 ( .A(n14987), .ZN(n21040) );
  AOI22_X1 U10248 ( .A1(\mem[633][2] ), .A2(n14985), .B1(n26497), .B2(
        data_in[2]), .ZN(n14987) );
  INV_X1 U10249 ( .A(n14988), .ZN(n21039) );
  AOI22_X1 U10250 ( .A1(\mem[633][3] ), .A2(n14985), .B1(n26497), .B2(
        data_in[3]), .ZN(n14988) );
  INV_X1 U10251 ( .A(n14989), .ZN(n21038) );
  AOI22_X1 U10252 ( .A1(\mem[633][4] ), .A2(n14985), .B1(n26497), .B2(
        data_in[4]), .ZN(n14989) );
  INV_X1 U10253 ( .A(n14990), .ZN(n21037) );
  AOI22_X1 U10254 ( .A1(\mem[633][5] ), .A2(n14985), .B1(n26497), .B2(
        data_in[5]), .ZN(n14990) );
  INV_X1 U10255 ( .A(n14991), .ZN(n21036) );
  AOI22_X1 U10256 ( .A1(\mem[633][6] ), .A2(n14985), .B1(n26497), .B2(
        data_in[6]), .ZN(n14991) );
  INV_X1 U10257 ( .A(n14992), .ZN(n21035) );
  AOI22_X1 U10258 ( .A1(\mem[633][7] ), .A2(n14985), .B1(n26497), .B2(
        data_in[7]), .ZN(n14992) );
  INV_X1 U10259 ( .A(n14993), .ZN(n21034) );
  AOI22_X1 U10260 ( .A1(\mem[634][0] ), .A2(n14994), .B1(n26496), .B2(
        data_in[0]), .ZN(n14993) );
  INV_X1 U10261 ( .A(n14995), .ZN(n21033) );
  AOI22_X1 U10262 ( .A1(\mem[634][1] ), .A2(n14994), .B1(n26496), .B2(
        data_in[1]), .ZN(n14995) );
  INV_X1 U10263 ( .A(n14996), .ZN(n21032) );
  AOI22_X1 U10264 ( .A1(\mem[634][2] ), .A2(n14994), .B1(n26496), .B2(
        data_in[2]), .ZN(n14996) );
  INV_X1 U10265 ( .A(n14997), .ZN(n21031) );
  AOI22_X1 U10266 ( .A1(\mem[634][3] ), .A2(n14994), .B1(n26496), .B2(
        data_in[3]), .ZN(n14997) );
  INV_X1 U10267 ( .A(n14998), .ZN(n21030) );
  AOI22_X1 U10268 ( .A1(\mem[634][4] ), .A2(n14994), .B1(n26496), .B2(
        data_in[4]), .ZN(n14998) );
  INV_X1 U10269 ( .A(n14999), .ZN(n21029) );
  AOI22_X1 U10270 ( .A1(\mem[634][5] ), .A2(n14994), .B1(n26496), .B2(
        data_in[5]), .ZN(n14999) );
  INV_X1 U10271 ( .A(n15000), .ZN(n21028) );
  AOI22_X1 U10272 ( .A1(\mem[634][6] ), .A2(n14994), .B1(n26496), .B2(
        data_in[6]), .ZN(n15000) );
  INV_X1 U10273 ( .A(n15001), .ZN(n21027) );
  AOI22_X1 U10274 ( .A1(\mem[634][7] ), .A2(n14994), .B1(n26496), .B2(
        data_in[7]), .ZN(n15001) );
  INV_X1 U10275 ( .A(n15002), .ZN(n21026) );
  AOI22_X1 U10276 ( .A1(\mem[635][0] ), .A2(n15003), .B1(n26495), .B2(
        data_in[0]), .ZN(n15002) );
  INV_X1 U10277 ( .A(n15004), .ZN(n21025) );
  AOI22_X1 U10278 ( .A1(\mem[635][1] ), .A2(n15003), .B1(n26495), .B2(
        data_in[1]), .ZN(n15004) );
  INV_X1 U10279 ( .A(n15005), .ZN(n21024) );
  AOI22_X1 U10280 ( .A1(\mem[635][2] ), .A2(n15003), .B1(n26495), .B2(
        data_in[2]), .ZN(n15005) );
  INV_X1 U10281 ( .A(n15006), .ZN(n21023) );
  AOI22_X1 U10282 ( .A1(\mem[635][3] ), .A2(n15003), .B1(n26495), .B2(
        data_in[3]), .ZN(n15006) );
  INV_X1 U10283 ( .A(n15007), .ZN(n21022) );
  AOI22_X1 U10284 ( .A1(\mem[635][4] ), .A2(n15003), .B1(n26495), .B2(
        data_in[4]), .ZN(n15007) );
  INV_X1 U10285 ( .A(n15008), .ZN(n21021) );
  AOI22_X1 U10286 ( .A1(\mem[635][5] ), .A2(n15003), .B1(n26495), .B2(
        data_in[5]), .ZN(n15008) );
  INV_X1 U10287 ( .A(n15009), .ZN(n21020) );
  AOI22_X1 U10288 ( .A1(\mem[635][6] ), .A2(n15003), .B1(n26495), .B2(
        data_in[6]), .ZN(n15009) );
  INV_X1 U10289 ( .A(n15010), .ZN(n21019) );
  AOI22_X1 U10290 ( .A1(\mem[635][7] ), .A2(n15003), .B1(n26495), .B2(
        data_in[7]), .ZN(n15010) );
  INV_X1 U10291 ( .A(n15011), .ZN(n21018) );
  AOI22_X1 U10292 ( .A1(\mem[636][0] ), .A2(n15012), .B1(n26494), .B2(
        data_in[0]), .ZN(n15011) );
  INV_X1 U10293 ( .A(n15013), .ZN(n21017) );
  AOI22_X1 U10294 ( .A1(\mem[636][1] ), .A2(n15012), .B1(n26494), .B2(
        data_in[1]), .ZN(n15013) );
  INV_X1 U10295 ( .A(n15014), .ZN(n21016) );
  AOI22_X1 U10296 ( .A1(\mem[636][2] ), .A2(n15012), .B1(n26494), .B2(
        data_in[2]), .ZN(n15014) );
  INV_X1 U10297 ( .A(n15015), .ZN(n21015) );
  AOI22_X1 U10298 ( .A1(\mem[636][3] ), .A2(n15012), .B1(n26494), .B2(
        data_in[3]), .ZN(n15015) );
  INV_X1 U10299 ( .A(n15016), .ZN(n21014) );
  AOI22_X1 U10300 ( .A1(\mem[636][4] ), .A2(n15012), .B1(n26494), .B2(
        data_in[4]), .ZN(n15016) );
  INV_X1 U10301 ( .A(n15017), .ZN(n21013) );
  AOI22_X1 U10302 ( .A1(\mem[636][5] ), .A2(n15012), .B1(n26494), .B2(
        data_in[5]), .ZN(n15017) );
  INV_X1 U10303 ( .A(n15018), .ZN(n21012) );
  AOI22_X1 U10304 ( .A1(\mem[636][6] ), .A2(n15012), .B1(n26494), .B2(
        data_in[6]), .ZN(n15018) );
  INV_X1 U10305 ( .A(n15019), .ZN(n21011) );
  AOI22_X1 U10306 ( .A1(\mem[636][7] ), .A2(n15012), .B1(n26494), .B2(
        data_in[7]), .ZN(n15019) );
  INV_X1 U10307 ( .A(n15020), .ZN(n21010) );
  AOI22_X1 U10308 ( .A1(\mem[637][0] ), .A2(n15021), .B1(n26493), .B2(
        data_in[0]), .ZN(n15020) );
  INV_X1 U10309 ( .A(n15022), .ZN(n21009) );
  AOI22_X1 U10310 ( .A1(\mem[637][1] ), .A2(n15021), .B1(n26493), .B2(
        data_in[1]), .ZN(n15022) );
  INV_X1 U10311 ( .A(n15023), .ZN(n21008) );
  AOI22_X1 U10312 ( .A1(\mem[637][2] ), .A2(n15021), .B1(n26493), .B2(
        data_in[2]), .ZN(n15023) );
  INV_X1 U10313 ( .A(n15024), .ZN(n21007) );
  AOI22_X1 U10314 ( .A1(\mem[637][3] ), .A2(n15021), .B1(n26493), .B2(
        data_in[3]), .ZN(n15024) );
  INV_X1 U10315 ( .A(n15025), .ZN(n21006) );
  AOI22_X1 U10316 ( .A1(\mem[637][4] ), .A2(n15021), .B1(n26493), .B2(
        data_in[4]), .ZN(n15025) );
  INV_X1 U10317 ( .A(n15026), .ZN(n21005) );
  AOI22_X1 U10318 ( .A1(\mem[637][5] ), .A2(n15021), .B1(n26493), .B2(
        data_in[5]), .ZN(n15026) );
  INV_X1 U10319 ( .A(n15027), .ZN(n21004) );
  AOI22_X1 U10320 ( .A1(\mem[637][6] ), .A2(n15021), .B1(n26493), .B2(
        data_in[6]), .ZN(n15027) );
  INV_X1 U10321 ( .A(n15028), .ZN(n21003) );
  AOI22_X1 U10322 ( .A1(\mem[637][7] ), .A2(n15021), .B1(n26493), .B2(
        data_in[7]), .ZN(n15028) );
  INV_X1 U10323 ( .A(n15029), .ZN(n21002) );
  AOI22_X1 U10324 ( .A1(\mem[638][0] ), .A2(n15030), .B1(n26492), .B2(
        data_in[0]), .ZN(n15029) );
  INV_X1 U10325 ( .A(n15031), .ZN(n21001) );
  AOI22_X1 U10326 ( .A1(\mem[638][1] ), .A2(n15030), .B1(n26492), .B2(
        data_in[1]), .ZN(n15031) );
  INV_X1 U10327 ( .A(n15032), .ZN(n21000) );
  AOI22_X1 U10328 ( .A1(\mem[638][2] ), .A2(n15030), .B1(n26492), .B2(
        data_in[2]), .ZN(n15032) );
  INV_X1 U10329 ( .A(n15033), .ZN(n20999) );
  AOI22_X1 U10330 ( .A1(\mem[638][3] ), .A2(n15030), .B1(n26492), .B2(
        data_in[3]), .ZN(n15033) );
  INV_X1 U10331 ( .A(n15034), .ZN(n20998) );
  AOI22_X1 U10332 ( .A1(\mem[638][4] ), .A2(n15030), .B1(n26492), .B2(
        data_in[4]), .ZN(n15034) );
  INV_X1 U10333 ( .A(n15035), .ZN(n20997) );
  AOI22_X1 U10334 ( .A1(\mem[638][5] ), .A2(n15030), .B1(n26492), .B2(
        data_in[5]), .ZN(n15035) );
  INV_X1 U10335 ( .A(n15036), .ZN(n20996) );
  AOI22_X1 U10336 ( .A1(\mem[638][6] ), .A2(n15030), .B1(n26492), .B2(
        data_in[6]), .ZN(n15036) );
  INV_X1 U10337 ( .A(n15037), .ZN(n20995) );
  AOI22_X1 U10338 ( .A1(\mem[638][7] ), .A2(n15030), .B1(n26492), .B2(
        data_in[7]), .ZN(n15037) );
  INV_X1 U10339 ( .A(n15038), .ZN(n20994) );
  AOI22_X1 U10340 ( .A1(\mem[639][0] ), .A2(n15039), .B1(n26491), .B2(
        data_in[0]), .ZN(n15038) );
  INV_X1 U10341 ( .A(n15040), .ZN(n20993) );
  AOI22_X1 U10342 ( .A1(\mem[639][1] ), .A2(n15039), .B1(n26491), .B2(
        data_in[1]), .ZN(n15040) );
  INV_X1 U10343 ( .A(n15041), .ZN(n20992) );
  AOI22_X1 U10344 ( .A1(\mem[639][2] ), .A2(n15039), .B1(n26491), .B2(
        data_in[2]), .ZN(n15041) );
  INV_X1 U10345 ( .A(n15042), .ZN(n20991) );
  AOI22_X1 U10346 ( .A1(\mem[639][3] ), .A2(n15039), .B1(n26491), .B2(
        data_in[3]), .ZN(n15042) );
  INV_X1 U10347 ( .A(n15043), .ZN(n20990) );
  AOI22_X1 U10348 ( .A1(\mem[639][4] ), .A2(n15039), .B1(n26491), .B2(
        data_in[4]), .ZN(n15043) );
  INV_X1 U10349 ( .A(n15044), .ZN(n20989) );
  AOI22_X1 U10350 ( .A1(\mem[639][5] ), .A2(n15039), .B1(n26491), .B2(
        data_in[5]), .ZN(n15044) );
  INV_X1 U10351 ( .A(n15045), .ZN(n20988) );
  AOI22_X1 U10352 ( .A1(\mem[639][6] ), .A2(n15039), .B1(n26491), .B2(
        data_in[6]), .ZN(n15045) );
  INV_X1 U10353 ( .A(n15046), .ZN(n20987) );
  AOI22_X1 U10354 ( .A1(\mem[639][7] ), .A2(n15039), .B1(n26491), .B2(
        data_in[7]), .ZN(n15046) );
  INV_X1 U10355 ( .A(n15120), .ZN(n20922) );
  AOI22_X1 U10356 ( .A1(\mem[648][0] ), .A2(n15121), .B1(n26482), .B2(
        data_in[0]), .ZN(n15120) );
  INV_X1 U10357 ( .A(n15122), .ZN(n20921) );
  AOI22_X1 U10358 ( .A1(\mem[648][1] ), .A2(n15121), .B1(n26482), .B2(
        data_in[1]), .ZN(n15122) );
  INV_X1 U10359 ( .A(n15123), .ZN(n20920) );
  AOI22_X1 U10360 ( .A1(\mem[648][2] ), .A2(n15121), .B1(n26482), .B2(
        data_in[2]), .ZN(n15123) );
  INV_X1 U10361 ( .A(n15124), .ZN(n20919) );
  AOI22_X1 U10362 ( .A1(\mem[648][3] ), .A2(n15121), .B1(n26482), .B2(
        data_in[3]), .ZN(n15124) );
  INV_X1 U10363 ( .A(n15125), .ZN(n20918) );
  AOI22_X1 U10364 ( .A1(\mem[648][4] ), .A2(n15121), .B1(n26482), .B2(
        data_in[4]), .ZN(n15125) );
  INV_X1 U10365 ( .A(n15126), .ZN(n20917) );
  AOI22_X1 U10366 ( .A1(\mem[648][5] ), .A2(n15121), .B1(n26482), .B2(
        data_in[5]), .ZN(n15126) );
  INV_X1 U10367 ( .A(n15127), .ZN(n20916) );
  AOI22_X1 U10368 ( .A1(\mem[648][6] ), .A2(n15121), .B1(n26482), .B2(
        data_in[6]), .ZN(n15127) );
  INV_X1 U10369 ( .A(n15128), .ZN(n20915) );
  AOI22_X1 U10370 ( .A1(\mem[648][7] ), .A2(n15121), .B1(n26482), .B2(
        data_in[7]), .ZN(n15128) );
  INV_X1 U10371 ( .A(n15129), .ZN(n20914) );
  AOI22_X1 U10372 ( .A1(\mem[649][0] ), .A2(n15130), .B1(n26481), .B2(
        data_in[0]), .ZN(n15129) );
  INV_X1 U10373 ( .A(n15131), .ZN(n20913) );
  AOI22_X1 U10374 ( .A1(\mem[649][1] ), .A2(n15130), .B1(n26481), .B2(
        data_in[1]), .ZN(n15131) );
  INV_X1 U10375 ( .A(n15132), .ZN(n20912) );
  AOI22_X1 U10376 ( .A1(\mem[649][2] ), .A2(n15130), .B1(n26481), .B2(
        data_in[2]), .ZN(n15132) );
  INV_X1 U10377 ( .A(n15133), .ZN(n20911) );
  AOI22_X1 U10378 ( .A1(\mem[649][3] ), .A2(n15130), .B1(n26481), .B2(
        data_in[3]), .ZN(n15133) );
  INV_X1 U10379 ( .A(n15134), .ZN(n20910) );
  AOI22_X1 U10380 ( .A1(\mem[649][4] ), .A2(n15130), .B1(n26481), .B2(
        data_in[4]), .ZN(n15134) );
  INV_X1 U10381 ( .A(n15135), .ZN(n20909) );
  AOI22_X1 U10382 ( .A1(\mem[649][5] ), .A2(n15130), .B1(n26481), .B2(
        data_in[5]), .ZN(n15135) );
  INV_X1 U10383 ( .A(n15136), .ZN(n20908) );
  AOI22_X1 U10384 ( .A1(\mem[649][6] ), .A2(n15130), .B1(n26481), .B2(
        data_in[6]), .ZN(n15136) );
  INV_X1 U10385 ( .A(n15137), .ZN(n20907) );
  AOI22_X1 U10386 ( .A1(\mem[649][7] ), .A2(n15130), .B1(n26481), .B2(
        data_in[7]), .ZN(n15137) );
  INV_X1 U10387 ( .A(n15138), .ZN(n20906) );
  AOI22_X1 U10388 ( .A1(\mem[650][0] ), .A2(n15139), .B1(n26480), .B2(
        data_in[0]), .ZN(n15138) );
  INV_X1 U10389 ( .A(n15140), .ZN(n20905) );
  AOI22_X1 U10390 ( .A1(\mem[650][1] ), .A2(n15139), .B1(n26480), .B2(
        data_in[1]), .ZN(n15140) );
  INV_X1 U10391 ( .A(n15141), .ZN(n20904) );
  AOI22_X1 U10392 ( .A1(\mem[650][2] ), .A2(n15139), .B1(n26480), .B2(
        data_in[2]), .ZN(n15141) );
  INV_X1 U10393 ( .A(n15142), .ZN(n20903) );
  AOI22_X1 U10394 ( .A1(\mem[650][3] ), .A2(n15139), .B1(n26480), .B2(
        data_in[3]), .ZN(n15142) );
  INV_X1 U10395 ( .A(n15143), .ZN(n20902) );
  AOI22_X1 U10396 ( .A1(\mem[650][4] ), .A2(n15139), .B1(n26480), .B2(
        data_in[4]), .ZN(n15143) );
  INV_X1 U10397 ( .A(n15144), .ZN(n20901) );
  AOI22_X1 U10398 ( .A1(\mem[650][5] ), .A2(n15139), .B1(n26480), .B2(
        data_in[5]), .ZN(n15144) );
  INV_X1 U10399 ( .A(n15145), .ZN(n20900) );
  AOI22_X1 U10400 ( .A1(\mem[650][6] ), .A2(n15139), .B1(n26480), .B2(
        data_in[6]), .ZN(n15145) );
  INV_X1 U10401 ( .A(n15146), .ZN(n20899) );
  AOI22_X1 U10402 ( .A1(\mem[650][7] ), .A2(n15139), .B1(n26480), .B2(
        data_in[7]), .ZN(n15146) );
  INV_X1 U10403 ( .A(n15147), .ZN(n20898) );
  AOI22_X1 U10404 ( .A1(\mem[651][0] ), .A2(n15148), .B1(n26479), .B2(
        data_in[0]), .ZN(n15147) );
  INV_X1 U10405 ( .A(n15149), .ZN(n20897) );
  AOI22_X1 U10406 ( .A1(\mem[651][1] ), .A2(n15148), .B1(n26479), .B2(
        data_in[1]), .ZN(n15149) );
  INV_X1 U10407 ( .A(n15150), .ZN(n20896) );
  AOI22_X1 U10408 ( .A1(\mem[651][2] ), .A2(n15148), .B1(n26479), .B2(
        data_in[2]), .ZN(n15150) );
  INV_X1 U10409 ( .A(n15151), .ZN(n20895) );
  AOI22_X1 U10410 ( .A1(\mem[651][3] ), .A2(n15148), .B1(n26479), .B2(
        data_in[3]), .ZN(n15151) );
  INV_X1 U10411 ( .A(n15152), .ZN(n20894) );
  AOI22_X1 U10412 ( .A1(\mem[651][4] ), .A2(n15148), .B1(n26479), .B2(
        data_in[4]), .ZN(n15152) );
  INV_X1 U10413 ( .A(n15153), .ZN(n20893) );
  AOI22_X1 U10414 ( .A1(\mem[651][5] ), .A2(n15148), .B1(n26479), .B2(
        data_in[5]), .ZN(n15153) );
  INV_X1 U10415 ( .A(n15154), .ZN(n20892) );
  AOI22_X1 U10416 ( .A1(\mem[651][6] ), .A2(n15148), .B1(n26479), .B2(
        data_in[6]), .ZN(n15154) );
  INV_X1 U10417 ( .A(n15155), .ZN(n20891) );
  AOI22_X1 U10418 ( .A1(\mem[651][7] ), .A2(n15148), .B1(n26479), .B2(
        data_in[7]), .ZN(n15155) );
  INV_X1 U10419 ( .A(n15156), .ZN(n20890) );
  AOI22_X1 U10420 ( .A1(\mem[652][0] ), .A2(n15157), .B1(n26478), .B2(
        data_in[0]), .ZN(n15156) );
  INV_X1 U10421 ( .A(n15158), .ZN(n20889) );
  AOI22_X1 U10422 ( .A1(\mem[652][1] ), .A2(n15157), .B1(n26478), .B2(
        data_in[1]), .ZN(n15158) );
  INV_X1 U10423 ( .A(n15159), .ZN(n20888) );
  AOI22_X1 U10424 ( .A1(\mem[652][2] ), .A2(n15157), .B1(n26478), .B2(
        data_in[2]), .ZN(n15159) );
  INV_X1 U10425 ( .A(n15160), .ZN(n20887) );
  AOI22_X1 U10426 ( .A1(\mem[652][3] ), .A2(n15157), .B1(n26478), .B2(
        data_in[3]), .ZN(n15160) );
  INV_X1 U10427 ( .A(n15161), .ZN(n20886) );
  AOI22_X1 U10428 ( .A1(\mem[652][4] ), .A2(n15157), .B1(n26478), .B2(
        data_in[4]), .ZN(n15161) );
  INV_X1 U10429 ( .A(n15162), .ZN(n20885) );
  AOI22_X1 U10430 ( .A1(\mem[652][5] ), .A2(n15157), .B1(n26478), .B2(
        data_in[5]), .ZN(n15162) );
  INV_X1 U10431 ( .A(n15163), .ZN(n20884) );
  AOI22_X1 U10432 ( .A1(\mem[652][6] ), .A2(n15157), .B1(n26478), .B2(
        data_in[6]), .ZN(n15163) );
  INV_X1 U10433 ( .A(n15164), .ZN(n20883) );
  AOI22_X1 U10434 ( .A1(\mem[652][7] ), .A2(n15157), .B1(n26478), .B2(
        data_in[7]), .ZN(n15164) );
  INV_X1 U10435 ( .A(n15165), .ZN(n20882) );
  AOI22_X1 U10436 ( .A1(\mem[653][0] ), .A2(n15166), .B1(n26477), .B2(
        data_in[0]), .ZN(n15165) );
  INV_X1 U10437 ( .A(n15167), .ZN(n20881) );
  AOI22_X1 U10438 ( .A1(\mem[653][1] ), .A2(n15166), .B1(n26477), .B2(
        data_in[1]), .ZN(n15167) );
  INV_X1 U10439 ( .A(n15168), .ZN(n20880) );
  AOI22_X1 U10440 ( .A1(\mem[653][2] ), .A2(n15166), .B1(n26477), .B2(
        data_in[2]), .ZN(n15168) );
  INV_X1 U10441 ( .A(n15169), .ZN(n20879) );
  AOI22_X1 U10442 ( .A1(\mem[653][3] ), .A2(n15166), .B1(n26477), .B2(
        data_in[3]), .ZN(n15169) );
  INV_X1 U10443 ( .A(n15170), .ZN(n20878) );
  AOI22_X1 U10444 ( .A1(\mem[653][4] ), .A2(n15166), .B1(n26477), .B2(
        data_in[4]), .ZN(n15170) );
  INV_X1 U10445 ( .A(n15171), .ZN(n20877) );
  AOI22_X1 U10446 ( .A1(\mem[653][5] ), .A2(n15166), .B1(n26477), .B2(
        data_in[5]), .ZN(n15171) );
  INV_X1 U10447 ( .A(n15172), .ZN(n20876) );
  AOI22_X1 U10448 ( .A1(\mem[653][6] ), .A2(n15166), .B1(n26477), .B2(
        data_in[6]), .ZN(n15172) );
  INV_X1 U10449 ( .A(n15173), .ZN(n20875) );
  AOI22_X1 U10450 ( .A1(\mem[653][7] ), .A2(n15166), .B1(n26477), .B2(
        data_in[7]), .ZN(n15173) );
  INV_X1 U10451 ( .A(n15174), .ZN(n20874) );
  AOI22_X1 U10452 ( .A1(\mem[654][0] ), .A2(n15175), .B1(n26476), .B2(
        data_in[0]), .ZN(n15174) );
  INV_X1 U10453 ( .A(n15176), .ZN(n20873) );
  AOI22_X1 U10454 ( .A1(\mem[654][1] ), .A2(n15175), .B1(n26476), .B2(
        data_in[1]), .ZN(n15176) );
  INV_X1 U10455 ( .A(n15177), .ZN(n20872) );
  AOI22_X1 U10456 ( .A1(\mem[654][2] ), .A2(n15175), .B1(n26476), .B2(
        data_in[2]), .ZN(n15177) );
  INV_X1 U10457 ( .A(n15178), .ZN(n20871) );
  AOI22_X1 U10458 ( .A1(\mem[654][3] ), .A2(n15175), .B1(n26476), .B2(
        data_in[3]), .ZN(n15178) );
  INV_X1 U10459 ( .A(n15179), .ZN(n20870) );
  AOI22_X1 U10460 ( .A1(\mem[654][4] ), .A2(n15175), .B1(n26476), .B2(
        data_in[4]), .ZN(n15179) );
  INV_X1 U10461 ( .A(n15180), .ZN(n20869) );
  AOI22_X1 U10462 ( .A1(\mem[654][5] ), .A2(n15175), .B1(n26476), .B2(
        data_in[5]), .ZN(n15180) );
  INV_X1 U10463 ( .A(n15181), .ZN(n20868) );
  AOI22_X1 U10464 ( .A1(\mem[654][6] ), .A2(n15175), .B1(n26476), .B2(
        data_in[6]), .ZN(n15181) );
  INV_X1 U10465 ( .A(n15182), .ZN(n20867) );
  AOI22_X1 U10466 ( .A1(\mem[654][7] ), .A2(n15175), .B1(n26476), .B2(
        data_in[7]), .ZN(n15182) );
  INV_X1 U10467 ( .A(n15183), .ZN(n20866) );
  AOI22_X1 U10468 ( .A1(\mem[655][0] ), .A2(n15184), .B1(n26475), .B2(
        data_in[0]), .ZN(n15183) );
  INV_X1 U10469 ( .A(n15185), .ZN(n20865) );
  AOI22_X1 U10470 ( .A1(\mem[655][1] ), .A2(n15184), .B1(n26475), .B2(
        data_in[1]), .ZN(n15185) );
  INV_X1 U10471 ( .A(n15186), .ZN(n20864) );
  AOI22_X1 U10472 ( .A1(\mem[655][2] ), .A2(n15184), .B1(n26475), .B2(
        data_in[2]), .ZN(n15186) );
  INV_X1 U10473 ( .A(n15187), .ZN(n20863) );
  AOI22_X1 U10474 ( .A1(\mem[655][3] ), .A2(n15184), .B1(n26475), .B2(
        data_in[3]), .ZN(n15187) );
  INV_X1 U10475 ( .A(n15188), .ZN(n20862) );
  AOI22_X1 U10476 ( .A1(\mem[655][4] ), .A2(n15184), .B1(n26475), .B2(
        data_in[4]), .ZN(n15188) );
  INV_X1 U10477 ( .A(n15189), .ZN(n20861) );
  AOI22_X1 U10478 ( .A1(\mem[655][5] ), .A2(n15184), .B1(n26475), .B2(
        data_in[5]), .ZN(n15189) );
  INV_X1 U10479 ( .A(n15190), .ZN(n20860) );
  AOI22_X1 U10480 ( .A1(\mem[655][6] ), .A2(n15184), .B1(n26475), .B2(
        data_in[6]), .ZN(n15190) );
  INV_X1 U10481 ( .A(n15191), .ZN(n20859) );
  AOI22_X1 U10482 ( .A1(\mem[655][7] ), .A2(n15184), .B1(n26475), .B2(
        data_in[7]), .ZN(n15191) );
  INV_X1 U10483 ( .A(n15192), .ZN(n20858) );
  AOI22_X1 U10484 ( .A1(\mem[656][0] ), .A2(n15193), .B1(n26474), .B2(
        data_in[0]), .ZN(n15192) );
  INV_X1 U10485 ( .A(n15194), .ZN(n20857) );
  AOI22_X1 U10486 ( .A1(\mem[656][1] ), .A2(n15193), .B1(n26474), .B2(
        data_in[1]), .ZN(n15194) );
  INV_X1 U10487 ( .A(n15195), .ZN(n20856) );
  AOI22_X1 U10488 ( .A1(\mem[656][2] ), .A2(n15193), .B1(n26474), .B2(
        data_in[2]), .ZN(n15195) );
  INV_X1 U10489 ( .A(n15196), .ZN(n20855) );
  AOI22_X1 U10490 ( .A1(\mem[656][3] ), .A2(n15193), .B1(n26474), .B2(
        data_in[3]), .ZN(n15196) );
  INV_X1 U10491 ( .A(n15197), .ZN(n20854) );
  AOI22_X1 U10492 ( .A1(\mem[656][4] ), .A2(n15193), .B1(n26474), .B2(
        data_in[4]), .ZN(n15197) );
  INV_X1 U10493 ( .A(n15198), .ZN(n20853) );
  AOI22_X1 U10494 ( .A1(\mem[656][5] ), .A2(n15193), .B1(n26474), .B2(
        data_in[5]), .ZN(n15198) );
  INV_X1 U10495 ( .A(n15199), .ZN(n20852) );
  AOI22_X1 U10496 ( .A1(\mem[656][6] ), .A2(n15193), .B1(n26474), .B2(
        data_in[6]), .ZN(n15199) );
  INV_X1 U10497 ( .A(n15200), .ZN(n20851) );
  AOI22_X1 U10498 ( .A1(\mem[656][7] ), .A2(n15193), .B1(n26474), .B2(
        data_in[7]), .ZN(n15200) );
  INV_X1 U10499 ( .A(n15201), .ZN(n20850) );
  AOI22_X1 U10500 ( .A1(\mem[657][0] ), .A2(n15202), .B1(n26473), .B2(
        data_in[0]), .ZN(n15201) );
  INV_X1 U10501 ( .A(n15203), .ZN(n20849) );
  AOI22_X1 U10502 ( .A1(\mem[657][1] ), .A2(n15202), .B1(n26473), .B2(
        data_in[1]), .ZN(n15203) );
  INV_X1 U10503 ( .A(n15204), .ZN(n20848) );
  AOI22_X1 U10504 ( .A1(\mem[657][2] ), .A2(n15202), .B1(n26473), .B2(
        data_in[2]), .ZN(n15204) );
  INV_X1 U10505 ( .A(n15205), .ZN(n20847) );
  AOI22_X1 U10506 ( .A1(\mem[657][3] ), .A2(n15202), .B1(n26473), .B2(
        data_in[3]), .ZN(n15205) );
  INV_X1 U10507 ( .A(n15206), .ZN(n20846) );
  AOI22_X1 U10508 ( .A1(\mem[657][4] ), .A2(n15202), .B1(n26473), .B2(
        data_in[4]), .ZN(n15206) );
  INV_X1 U10509 ( .A(n15207), .ZN(n20845) );
  AOI22_X1 U10510 ( .A1(\mem[657][5] ), .A2(n15202), .B1(n26473), .B2(
        data_in[5]), .ZN(n15207) );
  INV_X1 U10511 ( .A(n15208), .ZN(n20844) );
  AOI22_X1 U10512 ( .A1(\mem[657][6] ), .A2(n15202), .B1(n26473), .B2(
        data_in[6]), .ZN(n15208) );
  INV_X1 U10513 ( .A(n15209), .ZN(n20843) );
  AOI22_X1 U10514 ( .A1(\mem[657][7] ), .A2(n15202), .B1(n26473), .B2(
        data_in[7]), .ZN(n15209) );
  INV_X1 U10515 ( .A(n15210), .ZN(n20842) );
  AOI22_X1 U10516 ( .A1(\mem[658][0] ), .A2(n15211), .B1(n26472), .B2(
        data_in[0]), .ZN(n15210) );
  INV_X1 U10517 ( .A(n15212), .ZN(n20841) );
  AOI22_X1 U10518 ( .A1(\mem[658][1] ), .A2(n15211), .B1(n26472), .B2(
        data_in[1]), .ZN(n15212) );
  INV_X1 U10519 ( .A(n15213), .ZN(n20840) );
  AOI22_X1 U10520 ( .A1(\mem[658][2] ), .A2(n15211), .B1(n26472), .B2(
        data_in[2]), .ZN(n15213) );
  INV_X1 U10521 ( .A(n15214), .ZN(n20839) );
  AOI22_X1 U10522 ( .A1(\mem[658][3] ), .A2(n15211), .B1(n26472), .B2(
        data_in[3]), .ZN(n15214) );
  INV_X1 U10523 ( .A(n15215), .ZN(n20838) );
  AOI22_X1 U10524 ( .A1(\mem[658][4] ), .A2(n15211), .B1(n26472), .B2(
        data_in[4]), .ZN(n15215) );
  INV_X1 U10525 ( .A(n15216), .ZN(n20837) );
  AOI22_X1 U10526 ( .A1(\mem[658][5] ), .A2(n15211), .B1(n26472), .B2(
        data_in[5]), .ZN(n15216) );
  INV_X1 U10527 ( .A(n15217), .ZN(n20836) );
  AOI22_X1 U10528 ( .A1(\mem[658][6] ), .A2(n15211), .B1(n26472), .B2(
        data_in[6]), .ZN(n15217) );
  INV_X1 U10529 ( .A(n15218), .ZN(n20835) );
  AOI22_X1 U10530 ( .A1(\mem[658][7] ), .A2(n15211), .B1(n26472), .B2(
        data_in[7]), .ZN(n15218) );
  INV_X1 U10531 ( .A(n15219), .ZN(n20834) );
  AOI22_X1 U10532 ( .A1(\mem[659][0] ), .A2(n15220), .B1(n26471), .B2(
        data_in[0]), .ZN(n15219) );
  INV_X1 U10533 ( .A(n15221), .ZN(n20833) );
  AOI22_X1 U10534 ( .A1(\mem[659][1] ), .A2(n15220), .B1(n26471), .B2(
        data_in[1]), .ZN(n15221) );
  INV_X1 U10535 ( .A(n15222), .ZN(n20832) );
  AOI22_X1 U10536 ( .A1(\mem[659][2] ), .A2(n15220), .B1(n26471), .B2(
        data_in[2]), .ZN(n15222) );
  INV_X1 U10537 ( .A(n15223), .ZN(n20831) );
  AOI22_X1 U10538 ( .A1(\mem[659][3] ), .A2(n15220), .B1(n26471), .B2(
        data_in[3]), .ZN(n15223) );
  INV_X1 U10539 ( .A(n15224), .ZN(n20830) );
  AOI22_X1 U10540 ( .A1(\mem[659][4] ), .A2(n15220), .B1(n26471), .B2(
        data_in[4]), .ZN(n15224) );
  INV_X1 U10541 ( .A(n15225), .ZN(n20829) );
  AOI22_X1 U10542 ( .A1(\mem[659][5] ), .A2(n15220), .B1(n26471), .B2(
        data_in[5]), .ZN(n15225) );
  INV_X1 U10543 ( .A(n15226), .ZN(n20828) );
  AOI22_X1 U10544 ( .A1(\mem[659][6] ), .A2(n15220), .B1(n26471), .B2(
        data_in[6]), .ZN(n15226) );
  INV_X1 U10545 ( .A(n15227), .ZN(n20827) );
  AOI22_X1 U10546 ( .A1(\mem[659][7] ), .A2(n15220), .B1(n26471), .B2(
        data_in[7]), .ZN(n15227) );
  INV_X1 U10547 ( .A(n15228), .ZN(n20826) );
  AOI22_X1 U10548 ( .A1(\mem[660][0] ), .A2(n15229), .B1(n26470), .B2(
        data_in[0]), .ZN(n15228) );
  INV_X1 U10549 ( .A(n15230), .ZN(n20825) );
  AOI22_X1 U10550 ( .A1(\mem[660][1] ), .A2(n15229), .B1(n26470), .B2(
        data_in[1]), .ZN(n15230) );
  INV_X1 U10551 ( .A(n15231), .ZN(n20824) );
  AOI22_X1 U10552 ( .A1(\mem[660][2] ), .A2(n15229), .B1(n26470), .B2(
        data_in[2]), .ZN(n15231) );
  INV_X1 U10553 ( .A(n15232), .ZN(n20823) );
  AOI22_X1 U10554 ( .A1(\mem[660][3] ), .A2(n15229), .B1(n26470), .B2(
        data_in[3]), .ZN(n15232) );
  INV_X1 U10555 ( .A(n15233), .ZN(n20822) );
  AOI22_X1 U10556 ( .A1(\mem[660][4] ), .A2(n15229), .B1(n26470), .B2(
        data_in[4]), .ZN(n15233) );
  INV_X1 U10557 ( .A(n15234), .ZN(n20821) );
  AOI22_X1 U10558 ( .A1(\mem[660][5] ), .A2(n15229), .B1(n26470), .B2(
        data_in[5]), .ZN(n15234) );
  INV_X1 U10559 ( .A(n15235), .ZN(n20820) );
  AOI22_X1 U10560 ( .A1(\mem[660][6] ), .A2(n15229), .B1(n26470), .B2(
        data_in[6]), .ZN(n15235) );
  INV_X1 U10561 ( .A(n15236), .ZN(n20819) );
  AOI22_X1 U10562 ( .A1(\mem[660][7] ), .A2(n15229), .B1(n26470), .B2(
        data_in[7]), .ZN(n15236) );
  INV_X1 U10563 ( .A(n15237), .ZN(n20818) );
  AOI22_X1 U10564 ( .A1(\mem[661][0] ), .A2(n15238), .B1(n26469), .B2(
        data_in[0]), .ZN(n15237) );
  INV_X1 U10565 ( .A(n15239), .ZN(n20817) );
  AOI22_X1 U10566 ( .A1(\mem[661][1] ), .A2(n15238), .B1(n26469), .B2(
        data_in[1]), .ZN(n15239) );
  INV_X1 U10567 ( .A(n15240), .ZN(n20816) );
  AOI22_X1 U10568 ( .A1(\mem[661][2] ), .A2(n15238), .B1(n26469), .B2(
        data_in[2]), .ZN(n15240) );
  INV_X1 U10569 ( .A(n15241), .ZN(n20815) );
  AOI22_X1 U10570 ( .A1(\mem[661][3] ), .A2(n15238), .B1(n26469), .B2(
        data_in[3]), .ZN(n15241) );
  INV_X1 U10571 ( .A(n15242), .ZN(n20814) );
  AOI22_X1 U10572 ( .A1(\mem[661][4] ), .A2(n15238), .B1(n26469), .B2(
        data_in[4]), .ZN(n15242) );
  INV_X1 U10573 ( .A(n15243), .ZN(n20813) );
  AOI22_X1 U10574 ( .A1(\mem[661][5] ), .A2(n15238), .B1(n26469), .B2(
        data_in[5]), .ZN(n15243) );
  INV_X1 U10575 ( .A(n15244), .ZN(n20812) );
  AOI22_X1 U10576 ( .A1(\mem[661][6] ), .A2(n15238), .B1(n26469), .B2(
        data_in[6]), .ZN(n15244) );
  INV_X1 U10577 ( .A(n15245), .ZN(n20811) );
  AOI22_X1 U10578 ( .A1(\mem[661][7] ), .A2(n15238), .B1(n26469), .B2(
        data_in[7]), .ZN(n15245) );
  INV_X1 U10579 ( .A(n15246), .ZN(n20810) );
  AOI22_X1 U10580 ( .A1(\mem[662][0] ), .A2(n15247), .B1(n26468), .B2(
        data_in[0]), .ZN(n15246) );
  INV_X1 U10581 ( .A(n15248), .ZN(n20809) );
  AOI22_X1 U10582 ( .A1(\mem[662][1] ), .A2(n15247), .B1(n26468), .B2(
        data_in[1]), .ZN(n15248) );
  INV_X1 U10583 ( .A(n15249), .ZN(n20808) );
  AOI22_X1 U10584 ( .A1(\mem[662][2] ), .A2(n15247), .B1(n26468), .B2(
        data_in[2]), .ZN(n15249) );
  INV_X1 U10585 ( .A(n15250), .ZN(n20807) );
  AOI22_X1 U10586 ( .A1(\mem[662][3] ), .A2(n15247), .B1(n26468), .B2(
        data_in[3]), .ZN(n15250) );
  INV_X1 U10587 ( .A(n15251), .ZN(n20806) );
  AOI22_X1 U10588 ( .A1(\mem[662][4] ), .A2(n15247), .B1(n26468), .B2(
        data_in[4]), .ZN(n15251) );
  INV_X1 U10589 ( .A(n15252), .ZN(n20805) );
  AOI22_X1 U10590 ( .A1(\mem[662][5] ), .A2(n15247), .B1(n26468), .B2(
        data_in[5]), .ZN(n15252) );
  INV_X1 U10591 ( .A(n15253), .ZN(n20804) );
  AOI22_X1 U10592 ( .A1(\mem[662][6] ), .A2(n15247), .B1(n26468), .B2(
        data_in[6]), .ZN(n15253) );
  INV_X1 U10593 ( .A(n15254), .ZN(n20803) );
  AOI22_X1 U10594 ( .A1(\mem[662][7] ), .A2(n15247), .B1(n26468), .B2(
        data_in[7]), .ZN(n15254) );
  INV_X1 U10595 ( .A(n15255), .ZN(n20802) );
  AOI22_X1 U10596 ( .A1(\mem[663][0] ), .A2(n15256), .B1(n26467), .B2(
        data_in[0]), .ZN(n15255) );
  INV_X1 U10597 ( .A(n15257), .ZN(n20801) );
  AOI22_X1 U10598 ( .A1(\mem[663][1] ), .A2(n15256), .B1(n26467), .B2(
        data_in[1]), .ZN(n15257) );
  INV_X1 U10599 ( .A(n15258), .ZN(n20800) );
  AOI22_X1 U10600 ( .A1(\mem[663][2] ), .A2(n15256), .B1(n26467), .B2(
        data_in[2]), .ZN(n15258) );
  INV_X1 U10601 ( .A(n15259), .ZN(n20799) );
  AOI22_X1 U10602 ( .A1(\mem[663][3] ), .A2(n15256), .B1(n26467), .B2(
        data_in[3]), .ZN(n15259) );
  INV_X1 U10603 ( .A(n15260), .ZN(n20798) );
  AOI22_X1 U10604 ( .A1(\mem[663][4] ), .A2(n15256), .B1(n26467), .B2(
        data_in[4]), .ZN(n15260) );
  INV_X1 U10605 ( .A(n15261), .ZN(n20797) );
  AOI22_X1 U10606 ( .A1(\mem[663][5] ), .A2(n15256), .B1(n26467), .B2(
        data_in[5]), .ZN(n15261) );
  INV_X1 U10607 ( .A(n15262), .ZN(n20796) );
  AOI22_X1 U10608 ( .A1(\mem[663][6] ), .A2(n15256), .B1(n26467), .B2(
        data_in[6]), .ZN(n15262) );
  INV_X1 U10609 ( .A(n15263), .ZN(n20795) );
  AOI22_X1 U10610 ( .A1(\mem[663][7] ), .A2(n15256), .B1(n26467), .B2(
        data_in[7]), .ZN(n15263) );
  INV_X1 U10611 ( .A(n15264), .ZN(n20794) );
  AOI22_X1 U10612 ( .A1(\mem[664][0] ), .A2(n15265), .B1(n26466), .B2(
        data_in[0]), .ZN(n15264) );
  INV_X1 U10613 ( .A(n15266), .ZN(n20793) );
  AOI22_X1 U10614 ( .A1(\mem[664][1] ), .A2(n15265), .B1(n26466), .B2(
        data_in[1]), .ZN(n15266) );
  INV_X1 U10615 ( .A(n15267), .ZN(n20792) );
  AOI22_X1 U10616 ( .A1(\mem[664][2] ), .A2(n15265), .B1(n26466), .B2(
        data_in[2]), .ZN(n15267) );
  INV_X1 U10617 ( .A(n15268), .ZN(n20791) );
  AOI22_X1 U10618 ( .A1(\mem[664][3] ), .A2(n15265), .B1(n26466), .B2(
        data_in[3]), .ZN(n15268) );
  INV_X1 U10619 ( .A(n15269), .ZN(n20790) );
  AOI22_X1 U10620 ( .A1(\mem[664][4] ), .A2(n15265), .B1(n26466), .B2(
        data_in[4]), .ZN(n15269) );
  INV_X1 U10621 ( .A(n15270), .ZN(n20789) );
  AOI22_X1 U10622 ( .A1(\mem[664][5] ), .A2(n15265), .B1(n26466), .B2(
        data_in[5]), .ZN(n15270) );
  INV_X1 U10623 ( .A(n15271), .ZN(n20788) );
  AOI22_X1 U10624 ( .A1(\mem[664][6] ), .A2(n15265), .B1(n26466), .B2(
        data_in[6]), .ZN(n15271) );
  INV_X1 U10625 ( .A(n15272), .ZN(n20787) );
  AOI22_X1 U10626 ( .A1(\mem[664][7] ), .A2(n15265), .B1(n26466), .B2(
        data_in[7]), .ZN(n15272) );
  INV_X1 U10627 ( .A(n15273), .ZN(n20786) );
  AOI22_X1 U10628 ( .A1(\mem[665][0] ), .A2(n15274), .B1(n26465), .B2(
        data_in[0]), .ZN(n15273) );
  INV_X1 U10629 ( .A(n15275), .ZN(n20785) );
  AOI22_X1 U10630 ( .A1(\mem[665][1] ), .A2(n15274), .B1(n26465), .B2(
        data_in[1]), .ZN(n15275) );
  INV_X1 U10631 ( .A(n15276), .ZN(n20784) );
  AOI22_X1 U10632 ( .A1(\mem[665][2] ), .A2(n15274), .B1(n26465), .B2(
        data_in[2]), .ZN(n15276) );
  INV_X1 U10633 ( .A(n15277), .ZN(n20783) );
  AOI22_X1 U10634 ( .A1(\mem[665][3] ), .A2(n15274), .B1(n26465), .B2(
        data_in[3]), .ZN(n15277) );
  INV_X1 U10635 ( .A(n15278), .ZN(n20782) );
  AOI22_X1 U10636 ( .A1(\mem[665][4] ), .A2(n15274), .B1(n26465), .B2(
        data_in[4]), .ZN(n15278) );
  INV_X1 U10637 ( .A(n15279), .ZN(n20781) );
  AOI22_X1 U10638 ( .A1(\mem[665][5] ), .A2(n15274), .B1(n26465), .B2(
        data_in[5]), .ZN(n15279) );
  INV_X1 U10639 ( .A(n15280), .ZN(n20780) );
  AOI22_X1 U10640 ( .A1(\mem[665][6] ), .A2(n15274), .B1(n26465), .B2(
        data_in[6]), .ZN(n15280) );
  INV_X1 U10641 ( .A(n15281), .ZN(n20779) );
  AOI22_X1 U10642 ( .A1(\mem[665][7] ), .A2(n15274), .B1(n26465), .B2(
        data_in[7]), .ZN(n15281) );
  INV_X1 U10643 ( .A(n15282), .ZN(n20778) );
  AOI22_X1 U10644 ( .A1(\mem[666][0] ), .A2(n15283), .B1(n26464), .B2(
        data_in[0]), .ZN(n15282) );
  INV_X1 U10645 ( .A(n15284), .ZN(n20777) );
  AOI22_X1 U10646 ( .A1(\mem[666][1] ), .A2(n15283), .B1(n26464), .B2(
        data_in[1]), .ZN(n15284) );
  INV_X1 U10647 ( .A(n15285), .ZN(n20776) );
  AOI22_X1 U10648 ( .A1(\mem[666][2] ), .A2(n15283), .B1(n26464), .B2(
        data_in[2]), .ZN(n15285) );
  INV_X1 U10649 ( .A(n15286), .ZN(n20775) );
  AOI22_X1 U10650 ( .A1(\mem[666][3] ), .A2(n15283), .B1(n26464), .B2(
        data_in[3]), .ZN(n15286) );
  INV_X1 U10651 ( .A(n15287), .ZN(n20774) );
  AOI22_X1 U10652 ( .A1(\mem[666][4] ), .A2(n15283), .B1(n26464), .B2(
        data_in[4]), .ZN(n15287) );
  INV_X1 U10653 ( .A(n15288), .ZN(n20773) );
  AOI22_X1 U10654 ( .A1(\mem[666][5] ), .A2(n15283), .B1(n26464), .B2(
        data_in[5]), .ZN(n15288) );
  INV_X1 U10655 ( .A(n15289), .ZN(n20772) );
  AOI22_X1 U10656 ( .A1(\mem[666][6] ), .A2(n15283), .B1(n26464), .B2(
        data_in[6]), .ZN(n15289) );
  INV_X1 U10657 ( .A(n15290), .ZN(n20771) );
  AOI22_X1 U10658 ( .A1(\mem[666][7] ), .A2(n15283), .B1(n26464), .B2(
        data_in[7]), .ZN(n15290) );
  INV_X1 U10659 ( .A(n15291), .ZN(n20770) );
  AOI22_X1 U10660 ( .A1(\mem[667][0] ), .A2(n15292), .B1(n26463), .B2(
        data_in[0]), .ZN(n15291) );
  INV_X1 U10661 ( .A(n15293), .ZN(n20769) );
  AOI22_X1 U10662 ( .A1(\mem[667][1] ), .A2(n15292), .B1(n26463), .B2(
        data_in[1]), .ZN(n15293) );
  INV_X1 U10663 ( .A(n15294), .ZN(n20768) );
  AOI22_X1 U10664 ( .A1(\mem[667][2] ), .A2(n15292), .B1(n26463), .B2(
        data_in[2]), .ZN(n15294) );
  INV_X1 U10665 ( .A(n15295), .ZN(n20767) );
  AOI22_X1 U10666 ( .A1(\mem[667][3] ), .A2(n15292), .B1(n26463), .B2(
        data_in[3]), .ZN(n15295) );
  INV_X1 U10667 ( .A(n15296), .ZN(n20766) );
  AOI22_X1 U10668 ( .A1(\mem[667][4] ), .A2(n15292), .B1(n26463), .B2(
        data_in[4]), .ZN(n15296) );
  INV_X1 U10669 ( .A(n15297), .ZN(n20765) );
  AOI22_X1 U10670 ( .A1(\mem[667][5] ), .A2(n15292), .B1(n26463), .B2(
        data_in[5]), .ZN(n15297) );
  INV_X1 U10671 ( .A(n15298), .ZN(n20764) );
  AOI22_X1 U10672 ( .A1(\mem[667][6] ), .A2(n15292), .B1(n26463), .B2(
        data_in[6]), .ZN(n15298) );
  INV_X1 U10673 ( .A(n15299), .ZN(n20763) );
  AOI22_X1 U10674 ( .A1(\mem[667][7] ), .A2(n15292), .B1(n26463), .B2(
        data_in[7]), .ZN(n15299) );
  INV_X1 U10675 ( .A(n15300), .ZN(n20762) );
  AOI22_X1 U10676 ( .A1(\mem[668][0] ), .A2(n15301), .B1(n26462), .B2(
        data_in[0]), .ZN(n15300) );
  INV_X1 U10677 ( .A(n15302), .ZN(n20761) );
  AOI22_X1 U10678 ( .A1(\mem[668][1] ), .A2(n15301), .B1(n26462), .B2(
        data_in[1]), .ZN(n15302) );
  INV_X1 U10679 ( .A(n15303), .ZN(n20760) );
  AOI22_X1 U10680 ( .A1(\mem[668][2] ), .A2(n15301), .B1(n26462), .B2(
        data_in[2]), .ZN(n15303) );
  INV_X1 U10681 ( .A(n15304), .ZN(n20759) );
  AOI22_X1 U10682 ( .A1(\mem[668][3] ), .A2(n15301), .B1(n26462), .B2(
        data_in[3]), .ZN(n15304) );
  INV_X1 U10683 ( .A(n15305), .ZN(n20758) );
  AOI22_X1 U10684 ( .A1(\mem[668][4] ), .A2(n15301), .B1(n26462), .B2(
        data_in[4]), .ZN(n15305) );
  INV_X1 U10685 ( .A(n15306), .ZN(n20757) );
  AOI22_X1 U10686 ( .A1(\mem[668][5] ), .A2(n15301), .B1(n26462), .B2(
        data_in[5]), .ZN(n15306) );
  INV_X1 U10687 ( .A(n15307), .ZN(n20756) );
  AOI22_X1 U10688 ( .A1(\mem[668][6] ), .A2(n15301), .B1(n26462), .B2(
        data_in[6]), .ZN(n15307) );
  INV_X1 U10689 ( .A(n15308), .ZN(n20755) );
  AOI22_X1 U10690 ( .A1(\mem[668][7] ), .A2(n15301), .B1(n26462), .B2(
        data_in[7]), .ZN(n15308) );
  INV_X1 U10691 ( .A(n15309), .ZN(n20754) );
  AOI22_X1 U10692 ( .A1(\mem[669][0] ), .A2(n15310), .B1(n26461), .B2(
        data_in[0]), .ZN(n15309) );
  INV_X1 U10693 ( .A(n15311), .ZN(n20753) );
  AOI22_X1 U10694 ( .A1(\mem[669][1] ), .A2(n15310), .B1(n26461), .B2(
        data_in[1]), .ZN(n15311) );
  INV_X1 U10695 ( .A(n15312), .ZN(n20752) );
  AOI22_X1 U10696 ( .A1(\mem[669][2] ), .A2(n15310), .B1(n26461), .B2(
        data_in[2]), .ZN(n15312) );
  INV_X1 U10697 ( .A(n15313), .ZN(n20751) );
  AOI22_X1 U10698 ( .A1(\mem[669][3] ), .A2(n15310), .B1(n26461), .B2(
        data_in[3]), .ZN(n15313) );
  INV_X1 U10699 ( .A(n15314), .ZN(n20750) );
  AOI22_X1 U10700 ( .A1(\mem[669][4] ), .A2(n15310), .B1(n26461), .B2(
        data_in[4]), .ZN(n15314) );
  INV_X1 U10701 ( .A(n15315), .ZN(n20749) );
  AOI22_X1 U10702 ( .A1(\mem[669][5] ), .A2(n15310), .B1(n26461), .B2(
        data_in[5]), .ZN(n15315) );
  INV_X1 U10703 ( .A(n15316), .ZN(n20748) );
  AOI22_X1 U10704 ( .A1(\mem[669][6] ), .A2(n15310), .B1(n26461), .B2(
        data_in[6]), .ZN(n15316) );
  INV_X1 U10705 ( .A(n15317), .ZN(n20747) );
  AOI22_X1 U10706 ( .A1(\mem[669][7] ), .A2(n15310), .B1(n26461), .B2(
        data_in[7]), .ZN(n15317) );
  INV_X1 U10707 ( .A(n15318), .ZN(n20746) );
  AOI22_X1 U10708 ( .A1(\mem[670][0] ), .A2(n15319), .B1(n26460), .B2(
        data_in[0]), .ZN(n15318) );
  INV_X1 U10709 ( .A(n15320), .ZN(n20745) );
  AOI22_X1 U10710 ( .A1(\mem[670][1] ), .A2(n15319), .B1(n26460), .B2(
        data_in[1]), .ZN(n15320) );
  INV_X1 U10711 ( .A(n15321), .ZN(n20744) );
  AOI22_X1 U10712 ( .A1(\mem[670][2] ), .A2(n15319), .B1(n26460), .B2(
        data_in[2]), .ZN(n15321) );
  INV_X1 U10713 ( .A(n15322), .ZN(n20743) );
  AOI22_X1 U10714 ( .A1(\mem[670][3] ), .A2(n15319), .B1(n26460), .B2(
        data_in[3]), .ZN(n15322) );
  INV_X1 U10715 ( .A(n15323), .ZN(n20742) );
  AOI22_X1 U10716 ( .A1(\mem[670][4] ), .A2(n15319), .B1(n26460), .B2(
        data_in[4]), .ZN(n15323) );
  INV_X1 U10717 ( .A(n15324), .ZN(n20741) );
  AOI22_X1 U10718 ( .A1(\mem[670][5] ), .A2(n15319), .B1(n26460), .B2(
        data_in[5]), .ZN(n15324) );
  INV_X1 U10719 ( .A(n15325), .ZN(n20740) );
  AOI22_X1 U10720 ( .A1(\mem[670][6] ), .A2(n15319), .B1(n26460), .B2(
        data_in[6]), .ZN(n15325) );
  INV_X1 U10721 ( .A(n15326), .ZN(n20739) );
  AOI22_X1 U10722 ( .A1(\mem[670][7] ), .A2(n15319), .B1(n26460), .B2(
        data_in[7]), .ZN(n15326) );
  INV_X1 U10723 ( .A(n15327), .ZN(n20738) );
  AOI22_X1 U10724 ( .A1(\mem[671][0] ), .A2(n15328), .B1(n26459), .B2(
        data_in[0]), .ZN(n15327) );
  INV_X1 U10725 ( .A(n15329), .ZN(n20737) );
  AOI22_X1 U10726 ( .A1(\mem[671][1] ), .A2(n15328), .B1(n26459), .B2(
        data_in[1]), .ZN(n15329) );
  INV_X1 U10727 ( .A(n15330), .ZN(n20736) );
  AOI22_X1 U10728 ( .A1(\mem[671][2] ), .A2(n15328), .B1(n26459), .B2(
        data_in[2]), .ZN(n15330) );
  INV_X1 U10729 ( .A(n15331), .ZN(n20735) );
  AOI22_X1 U10730 ( .A1(\mem[671][3] ), .A2(n15328), .B1(n26459), .B2(
        data_in[3]), .ZN(n15331) );
  INV_X1 U10731 ( .A(n15332), .ZN(n20734) );
  AOI22_X1 U10732 ( .A1(\mem[671][4] ), .A2(n15328), .B1(n26459), .B2(
        data_in[4]), .ZN(n15332) );
  INV_X1 U10733 ( .A(n15333), .ZN(n20733) );
  AOI22_X1 U10734 ( .A1(\mem[671][5] ), .A2(n15328), .B1(n26459), .B2(
        data_in[5]), .ZN(n15333) );
  INV_X1 U10735 ( .A(n15334), .ZN(n20732) );
  AOI22_X1 U10736 ( .A1(\mem[671][6] ), .A2(n15328), .B1(n26459), .B2(
        data_in[6]), .ZN(n15334) );
  INV_X1 U10737 ( .A(n15335), .ZN(n20731) );
  AOI22_X1 U10738 ( .A1(\mem[671][7] ), .A2(n15328), .B1(n26459), .B2(
        data_in[7]), .ZN(n15335) );
  INV_X1 U10739 ( .A(n15409), .ZN(n20666) );
  AOI22_X1 U10740 ( .A1(\mem[680][0] ), .A2(n15410), .B1(n26450), .B2(
        data_in[0]), .ZN(n15409) );
  INV_X1 U10741 ( .A(n15411), .ZN(n20665) );
  AOI22_X1 U10742 ( .A1(\mem[680][1] ), .A2(n15410), .B1(n26450), .B2(
        data_in[1]), .ZN(n15411) );
  INV_X1 U10743 ( .A(n15412), .ZN(n20664) );
  AOI22_X1 U10744 ( .A1(\mem[680][2] ), .A2(n15410), .B1(n26450), .B2(
        data_in[2]), .ZN(n15412) );
  INV_X1 U10745 ( .A(n15413), .ZN(n20663) );
  AOI22_X1 U10746 ( .A1(\mem[680][3] ), .A2(n15410), .B1(n26450), .B2(
        data_in[3]), .ZN(n15413) );
  INV_X1 U10747 ( .A(n15414), .ZN(n20662) );
  AOI22_X1 U10748 ( .A1(\mem[680][4] ), .A2(n15410), .B1(n26450), .B2(
        data_in[4]), .ZN(n15414) );
  INV_X1 U10749 ( .A(n15415), .ZN(n20661) );
  AOI22_X1 U10750 ( .A1(\mem[680][5] ), .A2(n15410), .B1(n26450), .B2(
        data_in[5]), .ZN(n15415) );
  INV_X1 U10751 ( .A(n15416), .ZN(n20660) );
  AOI22_X1 U10752 ( .A1(\mem[680][6] ), .A2(n15410), .B1(n26450), .B2(
        data_in[6]), .ZN(n15416) );
  INV_X1 U10753 ( .A(n15417), .ZN(n20659) );
  AOI22_X1 U10754 ( .A1(\mem[680][7] ), .A2(n15410), .B1(n26450), .B2(
        data_in[7]), .ZN(n15417) );
  INV_X1 U10755 ( .A(n15418), .ZN(n20658) );
  AOI22_X1 U10756 ( .A1(\mem[681][0] ), .A2(n15419), .B1(n26449), .B2(
        data_in[0]), .ZN(n15418) );
  INV_X1 U10757 ( .A(n15420), .ZN(n20657) );
  AOI22_X1 U10758 ( .A1(\mem[681][1] ), .A2(n15419), .B1(n26449), .B2(
        data_in[1]), .ZN(n15420) );
  INV_X1 U10759 ( .A(n15421), .ZN(n20656) );
  AOI22_X1 U10760 ( .A1(\mem[681][2] ), .A2(n15419), .B1(n26449), .B2(
        data_in[2]), .ZN(n15421) );
  INV_X1 U10761 ( .A(n15422), .ZN(n20655) );
  AOI22_X1 U10762 ( .A1(\mem[681][3] ), .A2(n15419), .B1(n26449), .B2(
        data_in[3]), .ZN(n15422) );
  INV_X1 U10763 ( .A(n15423), .ZN(n20654) );
  AOI22_X1 U10764 ( .A1(\mem[681][4] ), .A2(n15419), .B1(n26449), .B2(
        data_in[4]), .ZN(n15423) );
  INV_X1 U10765 ( .A(n15424), .ZN(n20653) );
  AOI22_X1 U10766 ( .A1(\mem[681][5] ), .A2(n15419), .B1(n26449), .B2(
        data_in[5]), .ZN(n15424) );
  INV_X1 U10767 ( .A(n15425), .ZN(n20652) );
  AOI22_X1 U10768 ( .A1(\mem[681][6] ), .A2(n15419), .B1(n26449), .B2(
        data_in[6]), .ZN(n15425) );
  INV_X1 U10769 ( .A(n15426), .ZN(n20651) );
  AOI22_X1 U10770 ( .A1(\mem[681][7] ), .A2(n15419), .B1(n26449), .B2(
        data_in[7]), .ZN(n15426) );
  INV_X1 U10771 ( .A(n15427), .ZN(n20650) );
  AOI22_X1 U10772 ( .A1(\mem[682][0] ), .A2(n15428), .B1(n26448), .B2(
        data_in[0]), .ZN(n15427) );
  INV_X1 U10773 ( .A(n15429), .ZN(n20649) );
  AOI22_X1 U10774 ( .A1(\mem[682][1] ), .A2(n15428), .B1(n26448), .B2(
        data_in[1]), .ZN(n15429) );
  INV_X1 U10775 ( .A(n15430), .ZN(n20648) );
  AOI22_X1 U10776 ( .A1(\mem[682][2] ), .A2(n15428), .B1(n26448), .B2(
        data_in[2]), .ZN(n15430) );
  INV_X1 U10777 ( .A(n15431), .ZN(n20647) );
  AOI22_X1 U10778 ( .A1(\mem[682][3] ), .A2(n15428), .B1(n26448), .B2(
        data_in[3]), .ZN(n15431) );
  INV_X1 U10779 ( .A(n15432), .ZN(n20646) );
  AOI22_X1 U10780 ( .A1(\mem[682][4] ), .A2(n15428), .B1(n26448), .B2(
        data_in[4]), .ZN(n15432) );
  INV_X1 U10781 ( .A(n15433), .ZN(n20645) );
  AOI22_X1 U10782 ( .A1(\mem[682][5] ), .A2(n15428), .B1(n26448), .B2(
        data_in[5]), .ZN(n15433) );
  INV_X1 U10783 ( .A(n15434), .ZN(n20644) );
  AOI22_X1 U10784 ( .A1(\mem[682][6] ), .A2(n15428), .B1(n26448), .B2(
        data_in[6]), .ZN(n15434) );
  INV_X1 U10785 ( .A(n15435), .ZN(n20643) );
  AOI22_X1 U10786 ( .A1(\mem[682][7] ), .A2(n15428), .B1(n26448), .B2(
        data_in[7]), .ZN(n15435) );
  INV_X1 U10787 ( .A(n15436), .ZN(n20642) );
  AOI22_X1 U10788 ( .A1(\mem[683][0] ), .A2(n15437), .B1(n26447), .B2(
        data_in[0]), .ZN(n15436) );
  INV_X1 U10789 ( .A(n15438), .ZN(n20641) );
  AOI22_X1 U10790 ( .A1(\mem[683][1] ), .A2(n15437), .B1(n26447), .B2(
        data_in[1]), .ZN(n15438) );
  INV_X1 U10791 ( .A(n15439), .ZN(n20640) );
  AOI22_X1 U10792 ( .A1(\mem[683][2] ), .A2(n15437), .B1(n26447), .B2(
        data_in[2]), .ZN(n15439) );
  INV_X1 U10793 ( .A(n15440), .ZN(n20639) );
  AOI22_X1 U10794 ( .A1(\mem[683][3] ), .A2(n15437), .B1(n26447), .B2(
        data_in[3]), .ZN(n15440) );
  INV_X1 U10795 ( .A(n15441), .ZN(n20638) );
  AOI22_X1 U10796 ( .A1(\mem[683][4] ), .A2(n15437), .B1(n26447), .B2(
        data_in[4]), .ZN(n15441) );
  INV_X1 U10797 ( .A(n15442), .ZN(n20637) );
  AOI22_X1 U10798 ( .A1(\mem[683][5] ), .A2(n15437), .B1(n26447), .B2(
        data_in[5]), .ZN(n15442) );
  INV_X1 U10799 ( .A(n15443), .ZN(n20636) );
  AOI22_X1 U10800 ( .A1(\mem[683][6] ), .A2(n15437), .B1(n26447), .B2(
        data_in[6]), .ZN(n15443) );
  INV_X1 U10801 ( .A(n15444), .ZN(n20635) );
  AOI22_X1 U10802 ( .A1(\mem[683][7] ), .A2(n15437), .B1(n26447), .B2(
        data_in[7]), .ZN(n15444) );
  INV_X1 U10803 ( .A(n15445), .ZN(n20634) );
  AOI22_X1 U10804 ( .A1(\mem[684][0] ), .A2(n15446), .B1(n26446), .B2(
        data_in[0]), .ZN(n15445) );
  INV_X1 U10805 ( .A(n15447), .ZN(n20633) );
  AOI22_X1 U10806 ( .A1(\mem[684][1] ), .A2(n15446), .B1(n26446), .B2(
        data_in[1]), .ZN(n15447) );
  INV_X1 U10807 ( .A(n15448), .ZN(n20632) );
  AOI22_X1 U10808 ( .A1(\mem[684][2] ), .A2(n15446), .B1(n26446), .B2(
        data_in[2]), .ZN(n15448) );
  INV_X1 U10809 ( .A(n15449), .ZN(n20631) );
  AOI22_X1 U10810 ( .A1(\mem[684][3] ), .A2(n15446), .B1(n26446), .B2(
        data_in[3]), .ZN(n15449) );
  INV_X1 U10811 ( .A(n15450), .ZN(n20630) );
  AOI22_X1 U10812 ( .A1(\mem[684][4] ), .A2(n15446), .B1(n26446), .B2(
        data_in[4]), .ZN(n15450) );
  INV_X1 U10813 ( .A(n15451), .ZN(n20629) );
  AOI22_X1 U10814 ( .A1(\mem[684][5] ), .A2(n15446), .B1(n26446), .B2(
        data_in[5]), .ZN(n15451) );
  INV_X1 U10815 ( .A(n15452), .ZN(n20628) );
  AOI22_X1 U10816 ( .A1(\mem[684][6] ), .A2(n15446), .B1(n26446), .B2(
        data_in[6]), .ZN(n15452) );
  INV_X1 U10817 ( .A(n15453), .ZN(n20627) );
  AOI22_X1 U10818 ( .A1(\mem[684][7] ), .A2(n15446), .B1(n26446), .B2(
        data_in[7]), .ZN(n15453) );
  INV_X1 U10819 ( .A(n15454), .ZN(n20626) );
  AOI22_X1 U10820 ( .A1(\mem[685][0] ), .A2(n15455), .B1(n26445), .B2(
        data_in[0]), .ZN(n15454) );
  INV_X1 U10821 ( .A(n15456), .ZN(n20625) );
  AOI22_X1 U10822 ( .A1(\mem[685][1] ), .A2(n15455), .B1(n26445), .B2(
        data_in[1]), .ZN(n15456) );
  INV_X1 U10823 ( .A(n15457), .ZN(n20624) );
  AOI22_X1 U10824 ( .A1(\mem[685][2] ), .A2(n15455), .B1(n26445), .B2(
        data_in[2]), .ZN(n15457) );
  INV_X1 U10825 ( .A(n15458), .ZN(n20623) );
  AOI22_X1 U10826 ( .A1(\mem[685][3] ), .A2(n15455), .B1(n26445), .B2(
        data_in[3]), .ZN(n15458) );
  INV_X1 U10827 ( .A(n15459), .ZN(n20622) );
  AOI22_X1 U10828 ( .A1(\mem[685][4] ), .A2(n15455), .B1(n26445), .B2(
        data_in[4]), .ZN(n15459) );
  INV_X1 U10829 ( .A(n15460), .ZN(n20621) );
  AOI22_X1 U10830 ( .A1(\mem[685][5] ), .A2(n15455), .B1(n26445), .B2(
        data_in[5]), .ZN(n15460) );
  INV_X1 U10831 ( .A(n15461), .ZN(n20620) );
  AOI22_X1 U10832 ( .A1(\mem[685][6] ), .A2(n15455), .B1(n26445), .B2(
        data_in[6]), .ZN(n15461) );
  INV_X1 U10833 ( .A(n15462), .ZN(n20619) );
  AOI22_X1 U10834 ( .A1(\mem[685][7] ), .A2(n15455), .B1(n26445), .B2(
        data_in[7]), .ZN(n15462) );
  INV_X1 U10835 ( .A(n15463), .ZN(n20618) );
  AOI22_X1 U10836 ( .A1(\mem[686][0] ), .A2(n15464), .B1(n26444), .B2(
        data_in[0]), .ZN(n15463) );
  INV_X1 U10837 ( .A(n15465), .ZN(n20617) );
  AOI22_X1 U10838 ( .A1(\mem[686][1] ), .A2(n15464), .B1(n26444), .B2(
        data_in[1]), .ZN(n15465) );
  INV_X1 U10839 ( .A(n15466), .ZN(n20616) );
  AOI22_X1 U10840 ( .A1(\mem[686][2] ), .A2(n15464), .B1(n26444), .B2(
        data_in[2]), .ZN(n15466) );
  INV_X1 U10841 ( .A(n15467), .ZN(n20615) );
  AOI22_X1 U10842 ( .A1(\mem[686][3] ), .A2(n15464), .B1(n26444), .B2(
        data_in[3]), .ZN(n15467) );
  INV_X1 U10843 ( .A(n15468), .ZN(n20614) );
  AOI22_X1 U10844 ( .A1(\mem[686][4] ), .A2(n15464), .B1(n26444), .B2(
        data_in[4]), .ZN(n15468) );
  INV_X1 U10845 ( .A(n15469), .ZN(n20613) );
  AOI22_X1 U10846 ( .A1(\mem[686][5] ), .A2(n15464), .B1(n26444), .B2(
        data_in[5]), .ZN(n15469) );
  INV_X1 U10847 ( .A(n15470), .ZN(n20612) );
  AOI22_X1 U10848 ( .A1(\mem[686][6] ), .A2(n15464), .B1(n26444), .B2(
        data_in[6]), .ZN(n15470) );
  INV_X1 U10849 ( .A(n15471), .ZN(n20611) );
  AOI22_X1 U10850 ( .A1(\mem[686][7] ), .A2(n15464), .B1(n26444), .B2(
        data_in[7]), .ZN(n15471) );
  INV_X1 U10851 ( .A(n15472), .ZN(n20610) );
  AOI22_X1 U10852 ( .A1(\mem[687][0] ), .A2(n15473), .B1(n26443), .B2(
        data_in[0]), .ZN(n15472) );
  INV_X1 U10853 ( .A(n15474), .ZN(n20609) );
  AOI22_X1 U10854 ( .A1(\mem[687][1] ), .A2(n15473), .B1(n26443), .B2(
        data_in[1]), .ZN(n15474) );
  INV_X1 U10855 ( .A(n15475), .ZN(n20608) );
  AOI22_X1 U10856 ( .A1(\mem[687][2] ), .A2(n15473), .B1(n26443), .B2(
        data_in[2]), .ZN(n15475) );
  INV_X1 U10857 ( .A(n15476), .ZN(n20607) );
  AOI22_X1 U10858 ( .A1(\mem[687][3] ), .A2(n15473), .B1(n26443), .B2(
        data_in[3]), .ZN(n15476) );
  INV_X1 U10859 ( .A(n15477), .ZN(n20606) );
  AOI22_X1 U10860 ( .A1(\mem[687][4] ), .A2(n15473), .B1(n26443), .B2(
        data_in[4]), .ZN(n15477) );
  INV_X1 U10861 ( .A(n15478), .ZN(n20605) );
  AOI22_X1 U10862 ( .A1(\mem[687][5] ), .A2(n15473), .B1(n26443), .B2(
        data_in[5]), .ZN(n15478) );
  INV_X1 U10863 ( .A(n15479), .ZN(n20604) );
  AOI22_X1 U10864 ( .A1(\mem[687][6] ), .A2(n15473), .B1(n26443), .B2(
        data_in[6]), .ZN(n15479) );
  INV_X1 U10865 ( .A(n15480), .ZN(n20603) );
  AOI22_X1 U10866 ( .A1(\mem[687][7] ), .A2(n15473), .B1(n26443), .B2(
        data_in[7]), .ZN(n15480) );
  INV_X1 U10867 ( .A(n15481), .ZN(n20602) );
  AOI22_X1 U10868 ( .A1(\mem[688][0] ), .A2(n15482), .B1(n26442), .B2(
        data_in[0]), .ZN(n15481) );
  INV_X1 U10869 ( .A(n15483), .ZN(n20601) );
  AOI22_X1 U10870 ( .A1(\mem[688][1] ), .A2(n15482), .B1(n26442), .B2(
        data_in[1]), .ZN(n15483) );
  INV_X1 U10871 ( .A(n15484), .ZN(n20600) );
  AOI22_X1 U10872 ( .A1(\mem[688][2] ), .A2(n15482), .B1(n26442), .B2(
        data_in[2]), .ZN(n15484) );
  INV_X1 U10873 ( .A(n15485), .ZN(n20599) );
  AOI22_X1 U10874 ( .A1(\mem[688][3] ), .A2(n15482), .B1(n26442), .B2(
        data_in[3]), .ZN(n15485) );
  INV_X1 U10875 ( .A(n15486), .ZN(n20598) );
  AOI22_X1 U10876 ( .A1(\mem[688][4] ), .A2(n15482), .B1(n26442), .B2(
        data_in[4]), .ZN(n15486) );
  INV_X1 U10877 ( .A(n15487), .ZN(n20597) );
  AOI22_X1 U10878 ( .A1(\mem[688][5] ), .A2(n15482), .B1(n26442), .B2(
        data_in[5]), .ZN(n15487) );
  INV_X1 U10879 ( .A(n15488), .ZN(n20596) );
  AOI22_X1 U10880 ( .A1(\mem[688][6] ), .A2(n15482), .B1(n26442), .B2(
        data_in[6]), .ZN(n15488) );
  INV_X1 U10881 ( .A(n15489), .ZN(n20595) );
  AOI22_X1 U10882 ( .A1(\mem[688][7] ), .A2(n15482), .B1(n26442), .B2(
        data_in[7]), .ZN(n15489) );
  INV_X1 U10883 ( .A(n15490), .ZN(n20594) );
  AOI22_X1 U10884 ( .A1(\mem[689][0] ), .A2(n15491), .B1(n26441), .B2(
        data_in[0]), .ZN(n15490) );
  INV_X1 U10885 ( .A(n15492), .ZN(n20593) );
  AOI22_X1 U10886 ( .A1(\mem[689][1] ), .A2(n15491), .B1(n26441), .B2(
        data_in[1]), .ZN(n15492) );
  INV_X1 U10887 ( .A(n15493), .ZN(n20592) );
  AOI22_X1 U10888 ( .A1(\mem[689][2] ), .A2(n15491), .B1(n26441), .B2(
        data_in[2]), .ZN(n15493) );
  INV_X1 U10889 ( .A(n15494), .ZN(n20591) );
  AOI22_X1 U10890 ( .A1(\mem[689][3] ), .A2(n15491), .B1(n26441), .B2(
        data_in[3]), .ZN(n15494) );
  INV_X1 U10891 ( .A(n15495), .ZN(n20590) );
  AOI22_X1 U10892 ( .A1(\mem[689][4] ), .A2(n15491), .B1(n26441), .B2(
        data_in[4]), .ZN(n15495) );
  INV_X1 U10893 ( .A(n15496), .ZN(n20589) );
  AOI22_X1 U10894 ( .A1(\mem[689][5] ), .A2(n15491), .B1(n26441), .B2(
        data_in[5]), .ZN(n15496) );
  INV_X1 U10895 ( .A(n15497), .ZN(n20588) );
  AOI22_X1 U10896 ( .A1(\mem[689][6] ), .A2(n15491), .B1(n26441), .B2(
        data_in[6]), .ZN(n15497) );
  INV_X1 U10897 ( .A(n15498), .ZN(n20587) );
  AOI22_X1 U10898 ( .A1(\mem[689][7] ), .A2(n15491), .B1(n26441), .B2(
        data_in[7]), .ZN(n15498) );
  INV_X1 U10899 ( .A(n15499), .ZN(n20586) );
  AOI22_X1 U10900 ( .A1(\mem[690][0] ), .A2(n15500), .B1(n26440), .B2(
        data_in[0]), .ZN(n15499) );
  INV_X1 U10901 ( .A(n15501), .ZN(n20585) );
  AOI22_X1 U10902 ( .A1(\mem[690][1] ), .A2(n15500), .B1(n26440), .B2(
        data_in[1]), .ZN(n15501) );
  INV_X1 U10903 ( .A(n15502), .ZN(n20584) );
  AOI22_X1 U10904 ( .A1(\mem[690][2] ), .A2(n15500), .B1(n26440), .B2(
        data_in[2]), .ZN(n15502) );
  INV_X1 U10905 ( .A(n15503), .ZN(n20583) );
  AOI22_X1 U10906 ( .A1(\mem[690][3] ), .A2(n15500), .B1(n26440), .B2(
        data_in[3]), .ZN(n15503) );
  INV_X1 U10907 ( .A(n15504), .ZN(n20582) );
  AOI22_X1 U10908 ( .A1(\mem[690][4] ), .A2(n15500), .B1(n26440), .B2(
        data_in[4]), .ZN(n15504) );
  INV_X1 U10909 ( .A(n15505), .ZN(n20581) );
  AOI22_X1 U10910 ( .A1(\mem[690][5] ), .A2(n15500), .B1(n26440), .B2(
        data_in[5]), .ZN(n15505) );
  INV_X1 U10911 ( .A(n15506), .ZN(n20580) );
  AOI22_X1 U10912 ( .A1(\mem[690][6] ), .A2(n15500), .B1(n26440), .B2(
        data_in[6]), .ZN(n15506) );
  INV_X1 U10913 ( .A(n15507), .ZN(n20579) );
  AOI22_X1 U10914 ( .A1(\mem[690][7] ), .A2(n15500), .B1(n26440), .B2(
        data_in[7]), .ZN(n15507) );
  INV_X1 U10915 ( .A(n15508), .ZN(n20578) );
  AOI22_X1 U10916 ( .A1(\mem[691][0] ), .A2(n15509), .B1(n26439), .B2(
        data_in[0]), .ZN(n15508) );
  INV_X1 U10917 ( .A(n15510), .ZN(n20577) );
  AOI22_X1 U10918 ( .A1(\mem[691][1] ), .A2(n15509), .B1(n26439), .B2(
        data_in[1]), .ZN(n15510) );
  INV_X1 U10919 ( .A(n15511), .ZN(n20576) );
  AOI22_X1 U10920 ( .A1(\mem[691][2] ), .A2(n15509), .B1(n26439), .B2(
        data_in[2]), .ZN(n15511) );
  INV_X1 U10921 ( .A(n15512), .ZN(n20575) );
  AOI22_X1 U10922 ( .A1(\mem[691][3] ), .A2(n15509), .B1(n26439), .B2(
        data_in[3]), .ZN(n15512) );
  INV_X1 U10923 ( .A(n15513), .ZN(n20574) );
  AOI22_X1 U10924 ( .A1(\mem[691][4] ), .A2(n15509), .B1(n26439), .B2(
        data_in[4]), .ZN(n15513) );
  INV_X1 U10925 ( .A(n15514), .ZN(n20573) );
  AOI22_X1 U10926 ( .A1(\mem[691][5] ), .A2(n15509), .B1(n26439), .B2(
        data_in[5]), .ZN(n15514) );
  INV_X1 U10927 ( .A(n15515), .ZN(n20572) );
  AOI22_X1 U10928 ( .A1(\mem[691][6] ), .A2(n15509), .B1(n26439), .B2(
        data_in[6]), .ZN(n15515) );
  INV_X1 U10929 ( .A(n15516), .ZN(n20571) );
  AOI22_X1 U10930 ( .A1(\mem[691][7] ), .A2(n15509), .B1(n26439), .B2(
        data_in[7]), .ZN(n15516) );
  INV_X1 U10931 ( .A(n15517), .ZN(n20570) );
  AOI22_X1 U10932 ( .A1(\mem[692][0] ), .A2(n15518), .B1(n26438), .B2(
        data_in[0]), .ZN(n15517) );
  INV_X1 U10933 ( .A(n15519), .ZN(n20569) );
  AOI22_X1 U10934 ( .A1(\mem[692][1] ), .A2(n15518), .B1(n26438), .B2(
        data_in[1]), .ZN(n15519) );
  INV_X1 U10935 ( .A(n15520), .ZN(n20568) );
  AOI22_X1 U10936 ( .A1(\mem[692][2] ), .A2(n15518), .B1(n26438), .B2(
        data_in[2]), .ZN(n15520) );
  INV_X1 U10937 ( .A(n15521), .ZN(n20567) );
  AOI22_X1 U10938 ( .A1(\mem[692][3] ), .A2(n15518), .B1(n26438), .B2(
        data_in[3]), .ZN(n15521) );
  INV_X1 U10939 ( .A(n15522), .ZN(n20566) );
  AOI22_X1 U10940 ( .A1(\mem[692][4] ), .A2(n15518), .B1(n26438), .B2(
        data_in[4]), .ZN(n15522) );
  INV_X1 U10941 ( .A(n15523), .ZN(n20565) );
  AOI22_X1 U10942 ( .A1(\mem[692][5] ), .A2(n15518), .B1(n26438), .B2(
        data_in[5]), .ZN(n15523) );
  INV_X1 U10943 ( .A(n15524), .ZN(n20564) );
  AOI22_X1 U10944 ( .A1(\mem[692][6] ), .A2(n15518), .B1(n26438), .B2(
        data_in[6]), .ZN(n15524) );
  INV_X1 U10945 ( .A(n15525), .ZN(n20563) );
  AOI22_X1 U10946 ( .A1(\mem[692][7] ), .A2(n15518), .B1(n26438), .B2(
        data_in[7]), .ZN(n15525) );
  INV_X1 U10947 ( .A(n15526), .ZN(n20562) );
  AOI22_X1 U10948 ( .A1(\mem[693][0] ), .A2(n15527), .B1(n26437), .B2(
        data_in[0]), .ZN(n15526) );
  INV_X1 U10949 ( .A(n15528), .ZN(n20561) );
  AOI22_X1 U10950 ( .A1(\mem[693][1] ), .A2(n15527), .B1(n26437), .B2(
        data_in[1]), .ZN(n15528) );
  INV_X1 U10951 ( .A(n15529), .ZN(n20560) );
  AOI22_X1 U10952 ( .A1(\mem[693][2] ), .A2(n15527), .B1(n26437), .B2(
        data_in[2]), .ZN(n15529) );
  INV_X1 U10953 ( .A(n15530), .ZN(n20559) );
  AOI22_X1 U10954 ( .A1(\mem[693][3] ), .A2(n15527), .B1(n26437), .B2(
        data_in[3]), .ZN(n15530) );
  INV_X1 U10955 ( .A(n15531), .ZN(n20558) );
  AOI22_X1 U10956 ( .A1(\mem[693][4] ), .A2(n15527), .B1(n26437), .B2(
        data_in[4]), .ZN(n15531) );
  INV_X1 U10957 ( .A(n15532), .ZN(n20557) );
  AOI22_X1 U10958 ( .A1(\mem[693][5] ), .A2(n15527), .B1(n26437), .B2(
        data_in[5]), .ZN(n15532) );
  INV_X1 U10959 ( .A(n15533), .ZN(n20556) );
  AOI22_X1 U10960 ( .A1(\mem[693][6] ), .A2(n15527), .B1(n26437), .B2(
        data_in[6]), .ZN(n15533) );
  INV_X1 U10961 ( .A(n15534), .ZN(n20555) );
  AOI22_X1 U10962 ( .A1(\mem[693][7] ), .A2(n15527), .B1(n26437), .B2(
        data_in[7]), .ZN(n15534) );
  INV_X1 U10963 ( .A(n15535), .ZN(n20554) );
  AOI22_X1 U10964 ( .A1(\mem[694][0] ), .A2(n15536), .B1(n26436), .B2(
        data_in[0]), .ZN(n15535) );
  INV_X1 U10965 ( .A(n15537), .ZN(n20553) );
  AOI22_X1 U10966 ( .A1(\mem[694][1] ), .A2(n15536), .B1(n26436), .B2(
        data_in[1]), .ZN(n15537) );
  INV_X1 U10967 ( .A(n15538), .ZN(n20552) );
  AOI22_X1 U10968 ( .A1(\mem[694][2] ), .A2(n15536), .B1(n26436), .B2(
        data_in[2]), .ZN(n15538) );
  INV_X1 U10969 ( .A(n15539), .ZN(n20551) );
  AOI22_X1 U10970 ( .A1(\mem[694][3] ), .A2(n15536), .B1(n26436), .B2(
        data_in[3]), .ZN(n15539) );
  INV_X1 U10971 ( .A(n15540), .ZN(n20550) );
  AOI22_X1 U10972 ( .A1(\mem[694][4] ), .A2(n15536), .B1(n26436), .B2(
        data_in[4]), .ZN(n15540) );
  INV_X1 U10973 ( .A(n15541), .ZN(n20549) );
  AOI22_X1 U10974 ( .A1(\mem[694][5] ), .A2(n15536), .B1(n26436), .B2(
        data_in[5]), .ZN(n15541) );
  INV_X1 U10975 ( .A(n15542), .ZN(n20548) );
  AOI22_X1 U10976 ( .A1(\mem[694][6] ), .A2(n15536), .B1(n26436), .B2(
        data_in[6]), .ZN(n15542) );
  INV_X1 U10977 ( .A(n15543), .ZN(n20547) );
  AOI22_X1 U10978 ( .A1(\mem[694][7] ), .A2(n15536), .B1(n26436), .B2(
        data_in[7]), .ZN(n15543) );
  INV_X1 U10979 ( .A(n15544), .ZN(n20546) );
  AOI22_X1 U10980 ( .A1(\mem[695][0] ), .A2(n15545), .B1(n26435), .B2(
        data_in[0]), .ZN(n15544) );
  INV_X1 U10981 ( .A(n15546), .ZN(n20545) );
  AOI22_X1 U10982 ( .A1(\mem[695][1] ), .A2(n15545), .B1(n26435), .B2(
        data_in[1]), .ZN(n15546) );
  INV_X1 U10983 ( .A(n15547), .ZN(n20544) );
  AOI22_X1 U10984 ( .A1(\mem[695][2] ), .A2(n15545), .B1(n26435), .B2(
        data_in[2]), .ZN(n15547) );
  INV_X1 U10985 ( .A(n15548), .ZN(n20543) );
  AOI22_X1 U10986 ( .A1(\mem[695][3] ), .A2(n15545), .B1(n26435), .B2(
        data_in[3]), .ZN(n15548) );
  INV_X1 U10987 ( .A(n15549), .ZN(n20542) );
  AOI22_X1 U10988 ( .A1(\mem[695][4] ), .A2(n15545), .B1(n26435), .B2(
        data_in[4]), .ZN(n15549) );
  INV_X1 U10989 ( .A(n15550), .ZN(n20541) );
  AOI22_X1 U10990 ( .A1(\mem[695][5] ), .A2(n15545), .B1(n26435), .B2(
        data_in[5]), .ZN(n15550) );
  INV_X1 U10991 ( .A(n15551), .ZN(n20540) );
  AOI22_X1 U10992 ( .A1(\mem[695][6] ), .A2(n15545), .B1(n26435), .B2(
        data_in[6]), .ZN(n15551) );
  INV_X1 U10993 ( .A(n15552), .ZN(n20539) );
  AOI22_X1 U10994 ( .A1(\mem[695][7] ), .A2(n15545), .B1(n26435), .B2(
        data_in[7]), .ZN(n15552) );
  INV_X1 U10995 ( .A(n15553), .ZN(n20538) );
  AOI22_X1 U10996 ( .A1(\mem[696][0] ), .A2(n15554), .B1(n26434), .B2(
        data_in[0]), .ZN(n15553) );
  INV_X1 U10997 ( .A(n15555), .ZN(n20537) );
  AOI22_X1 U10998 ( .A1(\mem[696][1] ), .A2(n15554), .B1(n26434), .B2(
        data_in[1]), .ZN(n15555) );
  INV_X1 U10999 ( .A(n15556), .ZN(n20536) );
  AOI22_X1 U11000 ( .A1(\mem[696][2] ), .A2(n15554), .B1(n26434), .B2(
        data_in[2]), .ZN(n15556) );
  INV_X1 U11001 ( .A(n15557), .ZN(n20535) );
  AOI22_X1 U11002 ( .A1(\mem[696][3] ), .A2(n15554), .B1(n26434), .B2(
        data_in[3]), .ZN(n15557) );
  INV_X1 U11003 ( .A(n15558), .ZN(n20534) );
  AOI22_X1 U11004 ( .A1(\mem[696][4] ), .A2(n15554), .B1(n26434), .B2(
        data_in[4]), .ZN(n15558) );
  INV_X1 U11005 ( .A(n15559), .ZN(n20533) );
  AOI22_X1 U11006 ( .A1(\mem[696][5] ), .A2(n15554), .B1(n26434), .B2(
        data_in[5]), .ZN(n15559) );
  INV_X1 U11007 ( .A(n15560), .ZN(n20532) );
  AOI22_X1 U11008 ( .A1(\mem[696][6] ), .A2(n15554), .B1(n26434), .B2(
        data_in[6]), .ZN(n15560) );
  INV_X1 U11009 ( .A(n15561), .ZN(n20531) );
  AOI22_X1 U11010 ( .A1(\mem[696][7] ), .A2(n15554), .B1(n26434), .B2(
        data_in[7]), .ZN(n15561) );
  INV_X1 U11011 ( .A(n15562), .ZN(n20530) );
  AOI22_X1 U11012 ( .A1(\mem[697][0] ), .A2(n15563), .B1(n26433), .B2(
        data_in[0]), .ZN(n15562) );
  INV_X1 U11013 ( .A(n15564), .ZN(n20529) );
  AOI22_X1 U11014 ( .A1(\mem[697][1] ), .A2(n15563), .B1(n26433), .B2(
        data_in[1]), .ZN(n15564) );
  INV_X1 U11015 ( .A(n15565), .ZN(n20528) );
  AOI22_X1 U11016 ( .A1(\mem[697][2] ), .A2(n15563), .B1(n26433), .B2(
        data_in[2]), .ZN(n15565) );
  INV_X1 U11017 ( .A(n15566), .ZN(n20527) );
  AOI22_X1 U11018 ( .A1(\mem[697][3] ), .A2(n15563), .B1(n26433), .B2(
        data_in[3]), .ZN(n15566) );
  INV_X1 U11019 ( .A(n15567), .ZN(n20526) );
  AOI22_X1 U11020 ( .A1(\mem[697][4] ), .A2(n15563), .B1(n26433), .B2(
        data_in[4]), .ZN(n15567) );
  INV_X1 U11021 ( .A(n15568), .ZN(n20525) );
  AOI22_X1 U11022 ( .A1(\mem[697][5] ), .A2(n15563), .B1(n26433), .B2(
        data_in[5]), .ZN(n15568) );
  INV_X1 U11023 ( .A(n15569), .ZN(n20524) );
  AOI22_X1 U11024 ( .A1(\mem[697][6] ), .A2(n15563), .B1(n26433), .B2(
        data_in[6]), .ZN(n15569) );
  INV_X1 U11025 ( .A(n15570), .ZN(n20523) );
  AOI22_X1 U11026 ( .A1(\mem[697][7] ), .A2(n15563), .B1(n26433), .B2(
        data_in[7]), .ZN(n15570) );
  INV_X1 U11027 ( .A(n15571), .ZN(n20522) );
  AOI22_X1 U11028 ( .A1(\mem[698][0] ), .A2(n15572), .B1(n26432), .B2(
        data_in[0]), .ZN(n15571) );
  INV_X1 U11029 ( .A(n15573), .ZN(n20521) );
  AOI22_X1 U11030 ( .A1(\mem[698][1] ), .A2(n15572), .B1(n26432), .B2(
        data_in[1]), .ZN(n15573) );
  INV_X1 U11031 ( .A(n15574), .ZN(n20520) );
  AOI22_X1 U11032 ( .A1(\mem[698][2] ), .A2(n15572), .B1(n26432), .B2(
        data_in[2]), .ZN(n15574) );
  INV_X1 U11033 ( .A(n15575), .ZN(n20519) );
  AOI22_X1 U11034 ( .A1(\mem[698][3] ), .A2(n15572), .B1(n26432), .B2(
        data_in[3]), .ZN(n15575) );
  INV_X1 U11035 ( .A(n15576), .ZN(n20518) );
  AOI22_X1 U11036 ( .A1(\mem[698][4] ), .A2(n15572), .B1(n26432), .B2(
        data_in[4]), .ZN(n15576) );
  INV_X1 U11037 ( .A(n15577), .ZN(n20517) );
  AOI22_X1 U11038 ( .A1(\mem[698][5] ), .A2(n15572), .B1(n26432), .B2(
        data_in[5]), .ZN(n15577) );
  INV_X1 U11039 ( .A(n15578), .ZN(n20516) );
  AOI22_X1 U11040 ( .A1(\mem[698][6] ), .A2(n15572), .B1(n26432), .B2(
        data_in[6]), .ZN(n15578) );
  INV_X1 U11041 ( .A(n15579), .ZN(n20515) );
  AOI22_X1 U11042 ( .A1(\mem[698][7] ), .A2(n15572), .B1(n26432), .B2(
        data_in[7]), .ZN(n15579) );
  INV_X1 U11043 ( .A(n15580), .ZN(n20514) );
  AOI22_X1 U11044 ( .A1(\mem[699][0] ), .A2(n15581), .B1(n26431), .B2(
        data_in[0]), .ZN(n15580) );
  INV_X1 U11045 ( .A(n15582), .ZN(n20513) );
  AOI22_X1 U11046 ( .A1(\mem[699][1] ), .A2(n15581), .B1(n26431), .B2(
        data_in[1]), .ZN(n15582) );
  INV_X1 U11047 ( .A(n15583), .ZN(n20512) );
  AOI22_X1 U11048 ( .A1(\mem[699][2] ), .A2(n15581), .B1(n26431), .B2(
        data_in[2]), .ZN(n15583) );
  INV_X1 U11049 ( .A(n15584), .ZN(n20511) );
  AOI22_X1 U11050 ( .A1(\mem[699][3] ), .A2(n15581), .B1(n26431), .B2(
        data_in[3]), .ZN(n15584) );
  INV_X1 U11051 ( .A(n15585), .ZN(n20510) );
  AOI22_X1 U11052 ( .A1(\mem[699][4] ), .A2(n15581), .B1(n26431), .B2(
        data_in[4]), .ZN(n15585) );
  INV_X1 U11053 ( .A(n15586), .ZN(n20509) );
  AOI22_X1 U11054 ( .A1(\mem[699][5] ), .A2(n15581), .B1(n26431), .B2(
        data_in[5]), .ZN(n15586) );
  INV_X1 U11055 ( .A(n15587), .ZN(n20508) );
  AOI22_X1 U11056 ( .A1(\mem[699][6] ), .A2(n15581), .B1(n26431), .B2(
        data_in[6]), .ZN(n15587) );
  INV_X1 U11057 ( .A(n15588), .ZN(n20507) );
  AOI22_X1 U11058 ( .A1(\mem[699][7] ), .A2(n15581), .B1(n26431), .B2(
        data_in[7]), .ZN(n15588) );
  INV_X1 U11059 ( .A(n15589), .ZN(n20506) );
  AOI22_X1 U11060 ( .A1(\mem[700][0] ), .A2(n15590), .B1(n26430), .B2(
        data_in[0]), .ZN(n15589) );
  INV_X1 U11061 ( .A(n15591), .ZN(n20505) );
  AOI22_X1 U11062 ( .A1(\mem[700][1] ), .A2(n15590), .B1(n26430), .B2(
        data_in[1]), .ZN(n15591) );
  INV_X1 U11063 ( .A(n15592), .ZN(n20504) );
  AOI22_X1 U11064 ( .A1(\mem[700][2] ), .A2(n15590), .B1(n26430), .B2(
        data_in[2]), .ZN(n15592) );
  INV_X1 U11065 ( .A(n15593), .ZN(n20503) );
  AOI22_X1 U11066 ( .A1(\mem[700][3] ), .A2(n15590), .B1(n26430), .B2(
        data_in[3]), .ZN(n15593) );
  INV_X1 U11067 ( .A(n15594), .ZN(n20502) );
  AOI22_X1 U11068 ( .A1(\mem[700][4] ), .A2(n15590), .B1(n26430), .B2(
        data_in[4]), .ZN(n15594) );
  INV_X1 U11069 ( .A(n15595), .ZN(n20501) );
  AOI22_X1 U11070 ( .A1(\mem[700][5] ), .A2(n15590), .B1(n26430), .B2(
        data_in[5]), .ZN(n15595) );
  INV_X1 U11071 ( .A(n15596), .ZN(n20500) );
  AOI22_X1 U11072 ( .A1(\mem[700][6] ), .A2(n15590), .B1(n26430), .B2(
        data_in[6]), .ZN(n15596) );
  INV_X1 U11073 ( .A(n15597), .ZN(n20499) );
  AOI22_X1 U11074 ( .A1(\mem[700][7] ), .A2(n15590), .B1(n26430), .B2(
        data_in[7]), .ZN(n15597) );
  INV_X1 U11075 ( .A(n15598), .ZN(n20498) );
  AOI22_X1 U11076 ( .A1(\mem[701][0] ), .A2(n15599), .B1(n26429), .B2(
        data_in[0]), .ZN(n15598) );
  INV_X1 U11077 ( .A(n15600), .ZN(n20497) );
  AOI22_X1 U11078 ( .A1(\mem[701][1] ), .A2(n15599), .B1(n26429), .B2(
        data_in[1]), .ZN(n15600) );
  INV_X1 U11079 ( .A(n15601), .ZN(n20496) );
  AOI22_X1 U11080 ( .A1(\mem[701][2] ), .A2(n15599), .B1(n26429), .B2(
        data_in[2]), .ZN(n15601) );
  INV_X1 U11081 ( .A(n15602), .ZN(n20495) );
  AOI22_X1 U11082 ( .A1(\mem[701][3] ), .A2(n15599), .B1(n26429), .B2(
        data_in[3]), .ZN(n15602) );
  INV_X1 U11083 ( .A(n15603), .ZN(n20494) );
  AOI22_X1 U11084 ( .A1(\mem[701][4] ), .A2(n15599), .B1(n26429), .B2(
        data_in[4]), .ZN(n15603) );
  INV_X1 U11085 ( .A(n15604), .ZN(n20493) );
  AOI22_X1 U11086 ( .A1(\mem[701][5] ), .A2(n15599), .B1(n26429), .B2(
        data_in[5]), .ZN(n15604) );
  INV_X1 U11087 ( .A(n15605), .ZN(n20492) );
  AOI22_X1 U11088 ( .A1(\mem[701][6] ), .A2(n15599), .B1(n26429), .B2(
        data_in[6]), .ZN(n15605) );
  INV_X1 U11089 ( .A(n15606), .ZN(n20491) );
  AOI22_X1 U11090 ( .A1(\mem[701][7] ), .A2(n15599), .B1(n26429), .B2(
        data_in[7]), .ZN(n15606) );
  INV_X1 U11091 ( .A(n15607), .ZN(n20490) );
  AOI22_X1 U11092 ( .A1(\mem[702][0] ), .A2(n15608), .B1(n26428), .B2(
        data_in[0]), .ZN(n15607) );
  INV_X1 U11093 ( .A(n15609), .ZN(n20489) );
  AOI22_X1 U11094 ( .A1(\mem[702][1] ), .A2(n15608), .B1(n26428), .B2(
        data_in[1]), .ZN(n15609) );
  INV_X1 U11095 ( .A(n15610), .ZN(n20488) );
  AOI22_X1 U11096 ( .A1(\mem[702][2] ), .A2(n15608), .B1(n26428), .B2(
        data_in[2]), .ZN(n15610) );
  INV_X1 U11097 ( .A(n15611), .ZN(n20487) );
  AOI22_X1 U11098 ( .A1(\mem[702][3] ), .A2(n15608), .B1(n26428), .B2(
        data_in[3]), .ZN(n15611) );
  INV_X1 U11099 ( .A(n15612), .ZN(n20486) );
  AOI22_X1 U11100 ( .A1(\mem[702][4] ), .A2(n15608), .B1(n26428), .B2(
        data_in[4]), .ZN(n15612) );
  INV_X1 U11101 ( .A(n15613), .ZN(n20485) );
  AOI22_X1 U11102 ( .A1(\mem[702][5] ), .A2(n15608), .B1(n26428), .B2(
        data_in[5]), .ZN(n15613) );
  INV_X1 U11103 ( .A(n15614), .ZN(n20484) );
  AOI22_X1 U11104 ( .A1(\mem[702][6] ), .A2(n15608), .B1(n26428), .B2(
        data_in[6]), .ZN(n15614) );
  INV_X1 U11105 ( .A(n15615), .ZN(n20483) );
  AOI22_X1 U11106 ( .A1(\mem[702][7] ), .A2(n15608), .B1(n26428), .B2(
        data_in[7]), .ZN(n15615) );
  INV_X1 U11107 ( .A(n15616), .ZN(n20482) );
  AOI22_X1 U11108 ( .A1(\mem[703][0] ), .A2(n15617), .B1(n26427), .B2(
        data_in[0]), .ZN(n15616) );
  INV_X1 U11109 ( .A(n15618), .ZN(n20481) );
  AOI22_X1 U11110 ( .A1(\mem[703][1] ), .A2(n15617), .B1(n26427), .B2(
        data_in[1]), .ZN(n15618) );
  INV_X1 U11111 ( .A(n15619), .ZN(n20480) );
  AOI22_X1 U11112 ( .A1(\mem[703][2] ), .A2(n15617), .B1(n26427), .B2(
        data_in[2]), .ZN(n15619) );
  INV_X1 U11113 ( .A(n15620), .ZN(n20479) );
  AOI22_X1 U11114 ( .A1(\mem[703][3] ), .A2(n15617), .B1(n26427), .B2(
        data_in[3]), .ZN(n15620) );
  INV_X1 U11115 ( .A(n15621), .ZN(n20478) );
  AOI22_X1 U11116 ( .A1(\mem[703][4] ), .A2(n15617), .B1(n26427), .B2(
        data_in[4]), .ZN(n15621) );
  INV_X1 U11117 ( .A(n15622), .ZN(n20477) );
  AOI22_X1 U11118 ( .A1(\mem[703][5] ), .A2(n15617), .B1(n26427), .B2(
        data_in[5]), .ZN(n15622) );
  INV_X1 U11119 ( .A(n15623), .ZN(n20476) );
  AOI22_X1 U11120 ( .A1(\mem[703][6] ), .A2(n15617), .B1(n26427), .B2(
        data_in[6]), .ZN(n15623) );
  INV_X1 U11121 ( .A(n15624), .ZN(n20475) );
  AOI22_X1 U11122 ( .A1(\mem[703][7] ), .A2(n15617), .B1(n26427), .B2(
        data_in[7]), .ZN(n15624) );
  INV_X1 U11123 ( .A(n15698), .ZN(n20410) );
  AOI22_X1 U11124 ( .A1(\mem[712][0] ), .A2(n15699), .B1(n26418), .B2(
        data_in[0]), .ZN(n15698) );
  INV_X1 U11125 ( .A(n15700), .ZN(n20409) );
  AOI22_X1 U11126 ( .A1(\mem[712][1] ), .A2(n15699), .B1(n26418), .B2(
        data_in[1]), .ZN(n15700) );
  INV_X1 U11127 ( .A(n15701), .ZN(n20408) );
  AOI22_X1 U11128 ( .A1(\mem[712][2] ), .A2(n15699), .B1(n26418), .B2(
        data_in[2]), .ZN(n15701) );
  INV_X1 U11129 ( .A(n15702), .ZN(n20407) );
  AOI22_X1 U11130 ( .A1(\mem[712][3] ), .A2(n15699), .B1(n26418), .B2(
        data_in[3]), .ZN(n15702) );
  INV_X1 U11131 ( .A(n15703), .ZN(n20406) );
  AOI22_X1 U11132 ( .A1(\mem[712][4] ), .A2(n15699), .B1(n26418), .B2(
        data_in[4]), .ZN(n15703) );
  INV_X1 U11133 ( .A(n15704), .ZN(n20405) );
  AOI22_X1 U11134 ( .A1(\mem[712][5] ), .A2(n15699), .B1(n26418), .B2(
        data_in[5]), .ZN(n15704) );
  INV_X1 U11135 ( .A(n15705), .ZN(n20404) );
  AOI22_X1 U11136 ( .A1(\mem[712][6] ), .A2(n15699), .B1(n26418), .B2(
        data_in[6]), .ZN(n15705) );
  INV_X1 U11137 ( .A(n15706), .ZN(n20403) );
  AOI22_X1 U11138 ( .A1(\mem[712][7] ), .A2(n15699), .B1(n26418), .B2(
        data_in[7]), .ZN(n15706) );
  INV_X1 U11139 ( .A(n15707), .ZN(n20402) );
  AOI22_X1 U11140 ( .A1(\mem[713][0] ), .A2(n15708), .B1(n26417), .B2(
        data_in[0]), .ZN(n15707) );
  INV_X1 U11141 ( .A(n15709), .ZN(n20401) );
  AOI22_X1 U11142 ( .A1(\mem[713][1] ), .A2(n15708), .B1(n26417), .B2(
        data_in[1]), .ZN(n15709) );
  INV_X1 U11143 ( .A(n15710), .ZN(n20400) );
  AOI22_X1 U11144 ( .A1(\mem[713][2] ), .A2(n15708), .B1(n26417), .B2(
        data_in[2]), .ZN(n15710) );
  INV_X1 U11145 ( .A(n15711), .ZN(n20399) );
  AOI22_X1 U11146 ( .A1(\mem[713][3] ), .A2(n15708), .B1(n26417), .B2(
        data_in[3]), .ZN(n15711) );
  INV_X1 U11147 ( .A(n15712), .ZN(n20398) );
  AOI22_X1 U11148 ( .A1(\mem[713][4] ), .A2(n15708), .B1(n26417), .B2(
        data_in[4]), .ZN(n15712) );
  INV_X1 U11149 ( .A(n15713), .ZN(n20397) );
  AOI22_X1 U11150 ( .A1(\mem[713][5] ), .A2(n15708), .B1(n26417), .B2(
        data_in[5]), .ZN(n15713) );
  INV_X1 U11151 ( .A(n15714), .ZN(n20396) );
  AOI22_X1 U11152 ( .A1(\mem[713][6] ), .A2(n15708), .B1(n26417), .B2(
        data_in[6]), .ZN(n15714) );
  INV_X1 U11153 ( .A(n15715), .ZN(n20395) );
  AOI22_X1 U11154 ( .A1(\mem[713][7] ), .A2(n15708), .B1(n26417), .B2(
        data_in[7]), .ZN(n15715) );
  INV_X1 U11155 ( .A(n15716), .ZN(n20394) );
  AOI22_X1 U11156 ( .A1(\mem[714][0] ), .A2(n15717), .B1(n26416), .B2(
        data_in[0]), .ZN(n15716) );
  INV_X1 U11157 ( .A(n15718), .ZN(n20393) );
  AOI22_X1 U11158 ( .A1(\mem[714][1] ), .A2(n15717), .B1(n26416), .B2(
        data_in[1]), .ZN(n15718) );
  INV_X1 U11159 ( .A(n15719), .ZN(n20392) );
  AOI22_X1 U11160 ( .A1(\mem[714][2] ), .A2(n15717), .B1(n26416), .B2(
        data_in[2]), .ZN(n15719) );
  INV_X1 U11161 ( .A(n15720), .ZN(n20391) );
  AOI22_X1 U11162 ( .A1(\mem[714][3] ), .A2(n15717), .B1(n26416), .B2(
        data_in[3]), .ZN(n15720) );
  INV_X1 U11163 ( .A(n15721), .ZN(n20390) );
  AOI22_X1 U11164 ( .A1(\mem[714][4] ), .A2(n15717), .B1(n26416), .B2(
        data_in[4]), .ZN(n15721) );
  INV_X1 U11165 ( .A(n15722), .ZN(n20389) );
  AOI22_X1 U11166 ( .A1(\mem[714][5] ), .A2(n15717), .B1(n26416), .B2(
        data_in[5]), .ZN(n15722) );
  INV_X1 U11167 ( .A(n15723), .ZN(n20388) );
  AOI22_X1 U11168 ( .A1(\mem[714][6] ), .A2(n15717), .B1(n26416), .B2(
        data_in[6]), .ZN(n15723) );
  INV_X1 U11169 ( .A(n15724), .ZN(n20387) );
  AOI22_X1 U11170 ( .A1(\mem[714][7] ), .A2(n15717), .B1(n26416), .B2(
        data_in[7]), .ZN(n15724) );
  INV_X1 U11171 ( .A(n15725), .ZN(n20386) );
  AOI22_X1 U11172 ( .A1(\mem[715][0] ), .A2(n15726), .B1(n26415), .B2(
        data_in[0]), .ZN(n15725) );
  INV_X1 U11173 ( .A(n15727), .ZN(n20385) );
  AOI22_X1 U11174 ( .A1(\mem[715][1] ), .A2(n15726), .B1(n26415), .B2(
        data_in[1]), .ZN(n15727) );
  INV_X1 U11175 ( .A(n15728), .ZN(n20384) );
  AOI22_X1 U11176 ( .A1(\mem[715][2] ), .A2(n15726), .B1(n26415), .B2(
        data_in[2]), .ZN(n15728) );
  INV_X1 U11177 ( .A(n15729), .ZN(n20383) );
  AOI22_X1 U11178 ( .A1(\mem[715][3] ), .A2(n15726), .B1(n26415), .B2(
        data_in[3]), .ZN(n15729) );
  INV_X1 U11179 ( .A(n15730), .ZN(n20382) );
  AOI22_X1 U11180 ( .A1(\mem[715][4] ), .A2(n15726), .B1(n26415), .B2(
        data_in[4]), .ZN(n15730) );
  INV_X1 U11181 ( .A(n15731), .ZN(n20381) );
  AOI22_X1 U11182 ( .A1(\mem[715][5] ), .A2(n15726), .B1(n26415), .B2(
        data_in[5]), .ZN(n15731) );
  INV_X1 U11183 ( .A(n15732), .ZN(n20380) );
  AOI22_X1 U11184 ( .A1(\mem[715][6] ), .A2(n15726), .B1(n26415), .B2(
        data_in[6]), .ZN(n15732) );
  INV_X1 U11185 ( .A(n15733), .ZN(n20379) );
  AOI22_X1 U11186 ( .A1(\mem[715][7] ), .A2(n15726), .B1(n26415), .B2(
        data_in[7]), .ZN(n15733) );
  INV_X1 U11187 ( .A(n15734), .ZN(n20378) );
  AOI22_X1 U11188 ( .A1(\mem[716][0] ), .A2(n15735), .B1(n26414), .B2(
        data_in[0]), .ZN(n15734) );
  INV_X1 U11189 ( .A(n15736), .ZN(n20377) );
  AOI22_X1 U11190 ( .A1(\mem[716][1] ), .A2(n15735), .B1(n26414), .B2(
        data_in[1]), .ZN(n15736) );
  INV_X1 U11191 ( .A(n15737), .ZN(n20376) );
  AOI22_X1 U11192 ( .A1(\mem[716][2] ), .A2(n15735), .B1(n26414), .B2(
        data_in[2]), .ZN(n15737) );
  INV_X1 U11193 ( .A(n15738), .ZN(n20375) );
  AOI22_X1 U11194 ( .A1(\mem[716][3] ), .A2(n15735), .B1(n26414), .B2(
        data_in[3]), .ZN(n15738) );
  INV_X1 U11195 ( .A(n15739), .ZN(n20374) );
  AOI22_X1 U11196 ( .A1(\mem[716][4] ), .A2(n15735), .B1(n26414), .B2(
        data_in[4]), .ZN(n15739) );
  INV_X1 U11197 ( .A(n15740), .ZN(n20373) );
  AOI22_X1 U11198 ( .A1(\mem[716][5] ), .A2(n15735), .B1(n26414), .B2(
        data_in[5]), .ZN(n15740) );
  INV_X1 U11199 ( .A(n15741), .ZN(n20372) );
  AOI22_X1 U11200 ( .A1(\mem[716][6] ), .A2(n15735), .B1(n26414), .B2(
        data_in[6]), .ZN(n15741) );
  INV_X1 U11201 ( .A(n15742), .ZN(n20371) );
  AOI22_X1 U11202 ( .A1(\mem[716][7] ), .A2(n15735), .B1(n26414), .B2(
        data_in[7]), .ZN(n15742) );
  INV_X1 U11203 ( .A(n15743), .ZN(n20370) );
  AOI22_X1 U11204 ( .A1(\mem[717][0] ), .A2(n15744), .B1(n26413), .B2(
        data_in[0]), .ZN(n15743) );
  INV_X1 U11205 ( .A(n15745), .ZN(n20369) );
  AOI22_X1 U11206 ( .A1(\mem[717][1] ), .A2(n15744), .B1(n26413), .B2(
        data_in[1]), .ZN(n15745) );
  INV_X1 U11207 ( .A(n15746), .ZN(n20368) );
  AOI22_X1 U11208 ( .A1(\mem[717][2] ), .A2(n15744), .B1(n26413), .B2(
        data_in[2]), .ZN(n15746) );
  INV_X1 U11209 ( .A(n15747), .ZN(n20367) );
  AOI22_X1 U11210 ( .A1(\mem[717][3] ), .A2(n15744), .B1(n26413), .B2(
        data_in[3]), .ZN(n15747) );
  INV_X1 U11211 ( .A(n15748), .ZN(n20366) );
  AOI22_X1 U11212 ( .A1(\mem[717][4] ), .A2(n15744), .B1(n26413), .B2(
        data_in[4]), .ZN(n15748) );
  INV_X1 U11213 ( .A(n15749), .ZN(n20365) );
  AOI22_X1 U11214 ( .A1(\mem[717][5] ), .A2(n15744), .B1(n26413), .B2(
        data_in[5]), .ZN(n15749) );
  INV_X1 U11215 ( .A(n15750), .ZN(n20364) );
  AOI22_X1 U11216 ( .A1(\mem[717][6] ), .A2(n15744), .B1(n26413), .B2(
        data_in[6]), .ZN(n15750) );
  INV_X1 U11217 ( .A(n15751), .ZN(n20363) );
  AOI22_X1 U11218 ( .A1(\mem[717][7] ), .A2(n15744), .B1(n26413), .B2(
        data_in[7]), .ZN(n15751) );
  INV_X1 U11219 ( .A(n15752), .ZN(n20362) );
  AOI22_X1 U11220 ( .A1(\mem[718][0] ), .A2(n15753), .B1(n26412), .B2(
        data_in[0]), .ZN(n15752) );
  INV_X1 U11221 ( .A(n15754), .ZN(n20361) );
  AOI22_X1 U11222 ( .A1(\mem[718][1] ), .A2(n15753), .B1(n26412), .B2(
        data_in[1]), .ZN(n15754) );
  INV_X1 U11223 ( .A(n15755), .ZN(n20360) );
  AOI22_X1 U11224 ( .A1(\mem[718][2] ), .A2(n15753), .B1(n26412), .B2(
        data_in[2]), .ZN(n15755) );
  INV_X1 U11225 ( .A(n15756), .ZN(n20359) );
  AOI22_X1 U11226 ( .A1(\mem[718][3] ), .A2(n15753), .B1(n26412), .B2(
        data_in[3]), .ZN(n15756) );
  INV_X1 U11227 ( .A(n15757), .ZN(n20358) );
  AOI22_X1 U11228 ( .A1(\mem[718][4] ), .A2(n15753), .B1(n26412), .B2(
        data_in[4]), .ZN(n15757) );
  INV_X1 U11229 ( .A(n15758), .ZN(n20357) );
  AOI22_X1 U11230 ( .A1(\mem[718][5] ), .A2(n15753), .B1(n26412), .B2(
        data_in[5]), .ZN(n15758) );
  INV_X1 U11231 ( .A(n15759), .ZN(n20356) );
  AOI22_X1 U11232 ( .A1(\mem[718][6] ), .A2(n15753), .B1(n26412), .B2(
        data_in[6]), .ZN(n15759) );
  INV_X1 U11233 ( .A(n15760), .ZN(n20355) );
  AOI22_X1 U11234 ( .A1(\mem[718][7] ), .A2(n15753), .B1(n26412), .B2(
        data_in[7]), .ZN(n15760) );
  INV_X1 U11235 ( .A(n15761), .ZN(n20354) );
  AOI22_X1 U11236 ( .A1(\mem[719][0] ), .A2(n15762), .B1(n26411), .B2(
        data_in[0]), .ZN(n15761) );
  INV_X1 U11237 ( .A(n15763), .ZN(n20353) );
  AOI22_X1 U11238 ( .A1(\mem[719][1] ), .A2(n15762), .B1(n26411), .B2(
        data_in[1]), .ZN(n15763) );
  INV_X1 U11239 ( .A(n15764), .ZN(n20352) );
  AOI22_X1 U11240 ( .A1(\mem[719][2] ), .A2(n15762), .B1(n26411), .B2(
        data_in[2]), .ZN(n15764) );
  INV_X1 U11241 ( .A(n15765), .ZN(n20351) );
  AOI22_X1 U11242 ( .A1(\mem[719][3] ), .A2(n15762), .B1(n26411), .B2(
        data_in[3]), .ZN(n15765) );
  INV_X1 U11243 ( .A(n15766), .ZN(n20350) );
  AOI22_X1 U11244 ( .A1(\mem[719][4] ), .A2(n15762), .B1(n26411), .B2(
        data_in[4]), .ZN(n15766) );
  INV_X1 U11245 ( .A(n15767), .ZN(n20349) );
  AOI22_X1 U11246 ( .A1(\mem[719][5] ), .A2(n15762), .B1(n26411), .B2(
        data_in[5]), .ZN(n15767) );
  INV_X1 U11247 ( .A(n15768), .ZN(n20348) );
  AOI22_X1 U11248 ( .A1(\mem[719][6] ), .A2(n15762), .B1(n26411), .B2(
        data_in[6]), .ZN(n15768) );
  INV_X1 U11249 ( .A(n15769), .ZN(n20347) );
  AOI22_X1 U11250 ( .A1(\mem[719][7] ), .A2(n15762), .B1(n26411), .B2(
        data_in[7]), .ZN(n15769) );
  INV_X1 U11251 ( .A(n15770), .ZN(n20346) );
  AOI22_X1 U11252 ( .A1(\mem[720][0] ), .A2(n15771), .B1(n26410), .B2(
        data_in[0]), .ZN(n15770) );
  INV_X1 U11253 ( .A(n15772), .ZN(n20345) );
  AOI22_X1 U11254 ( .A1(\mem[720][1] ), .A2(n15771), .B1(n26410), .B2(
        data_in[1]), .ZN(n15772) );
  INV_X1 U11255 ( .A(n15773), .ZN(n20344) );
  AOI22_X1 U11256 ( .A1(\mem[720][2] ), .A2(n15771), .B1(n26410), .B2(
        data_in[2]), .ZN(n15773) );
  INV_X1 U11257 ( .A(n15774), .ZN(n20343) );
  AOI22_X1 U11258 ( .A1(\mem[720][3] ), .A2(n15771), .B1(n26410), .B2(
        data_in[3]), .ZN(n15774) );
  INV_X1 U11259 ( .A(n15775), .ZN(n20342) );
  AOI22_X1 U11260 ( .A1(\mem[720][4] ), .A2(n15771), .B1(n26410), .B2(
        data_in[4]), .ZN(n15775) );
  INV_X1 U11261 ( .A(n15776), .ZN(n20341) );
  AOI22_X1 U11262 ( .A1(\mem[720][5] ), .A2(n15771), .B1(n26410), .B2(
        data_in[5]), .ZN(n15776) );
  INV_X1 U11263 ( .A(n15777), .ZN(n20340) );
  AOI22_X1 U11264 ( .A1(\mem[720][6] ), .A2(n15771), .B1(n26410), .B2(
        data_in[6]), .ZN(n15777) );
  INV_X1 U11265 ( .A(n15778), .ZN(n20339) );
  AOI22_X1 U11266 ( .A1(\mem[720][7] ), .A2(n15771), .B1(n26410), .B2(
        data_in[7]), .ZN(n15778) );
  INV_X1 U11267 ( .A(n15779), .ZN(n20338) );
  AOI22_X1 U11268 ( .A1(\mem[721][0] ), .A2(n15780), .B1(n26409), .B2(
        data_in[0]), .ZN(n15779) );
  INV_X1 U11269 ( .A(n15781), .ZN(n20337) );
  AOI22_X1 U11270 ( .A1(\mem[721][1] ), .A2(n15780), .B1(n26409), .B2(
        data_in[1]), .ZN(n15781) );
  INV_X1 U11271 ( .A(n15782), .ZN(n20336) );
  AOI22_X1 U11272 ( .A1(\mem[721][2] ), .A2(n15780), .B1(n26409), .B2(
        data_in[2]), .ZN(n15782) );
  INV_X1 U11273 ( .A(n15783), .ZN(n20335) );
  AOI22_X1 U11274 ( .A1(\mem[721][3] ), .A2(n15780), .B1(n26409), .B2(
        data_in[3]), .ZN(n15783) );
  INV_X1 U11275 ( .A(n15784), .ZN(n20334) );
  AOI22_X1 U11276 ( .A1(\mem[721][4] ), .A2(n15780), .B1(n26409), .B2(
        data_in[4]), .ZN(n15784) );
  INV_X1 U11277 ( .A(n15785), .ZN(n20333) );
  AOI22_X1 U11278 ( .A1(\mem[721][5] ), .A2(n15780), .B1(n26409), .B2(
        data_in[5]), .ZN(n15785) );
  INV_X1 U11279 ( .A(n15786), .ZN(n20332) );
  AOI22_X1 U11280 ( .A1(\mem[721][6] ), .A2(n15780), .B1(n26409), .B2(
        data_in[6]), .ZN(n15786) );
  INV_X1 U11281 ( .A(n15787), .ZN(n20331) );
  AOI22_X1 U11282 ( .A1(\mem[721][7] ), .A2(n15780), .B1(n26409), .B2(
        data_in[7]), .ZN(n15787) );
  INV_X1 U11283 ( .A(n15788), .ZN(n20330) );
  AOI22_X1 U11284 ( .A1(\mem[722][0] ), .A2(n15789), .B1(n26408), .B2(
        data_in[0]), .ZN(n15788) );
  INV_X1 U11285 ( .A(n15790), .ZN(n20329) );
  AOI22_X1 U11286 ( .A1(\mem[722][1] ), .A2(n15789), .B1(n26408), .B2(
        data_in[1]), .ZN(n15790) );
  INV_X1 U11287 ( .A(n15791), .ZN(n20328) );
  AOI22_X1 U11288 ( .A1(\mem[722][2] ), .A2(n15789), .B1(n26408), .B2(
        data_in[2]), .ZN(n15791) );
  INV_X1 U11289 ( .A(n15792), .ZN(n20327) );
  AOI22_X1 U11290 ( .A1(\mem[722][3] ), .A2(n15789), .B1(n26408), .B2(
        data_in[3]), .ZN(n15792) );
  INV_X1 U11291 ( .A(n15793), .ZN(n20326) );
  AOI22_X1 U11292 ( .A1(\mem[722][4] ), .A2(n15789), .B1(n26408), .B2(
        data_in[4]), .ZN(n15793) );
  INV_X1 U11293 ( .A(n15794), .ZN(n20325) );
  AOI22_X1 U11294 ( .A1(\mem[722][5] ), .A2(n15789), .B1(n26408), .B2(
        data_in[5]), .ZN(n15794) );
  INV_X1 U11295 ( .A(n15795), .ZN(n20324) );
  AOI22_X1 U11296 ( .A1(\mem[722][6] ), .A2(n15789), .B1(n26408), .B2(
        data_in[6]), .ZN(n15795) );
  INV_X1 U11297 ( .A(n15796), .ZN(n20323) );
  AOI22_X1 U11298 ( .A1(\mem[722][7] ), .A2(n15789), .B1(n26408), .B2(
        data_in[7]), .ZN(n15796) );
  INV_X1 U11299 ( .A(n15797), .ZN(n20322) );
  AOI22_X1 U11300 ( .A1(\mem[723][0] ), .A2(n15798), .B1(n26407), .B2(
        data_in[0]), .ZN(n15797) );
  INV_X1 U11301 ( .A(n15799), .ZN(n20321) );
  AOI22_X1 U11302 ( .A1(\mem[723][1] ), .A2(n15798), .B1(n26407), .B2(
        data_in[1]), .ZN(n15799) );
  INV_X1 U11303 ( .A(n15800), .ZN(n20320) );
  AOI22_X1 U11304 ( .A1(\mem[723][2] ), .A2(n15798), .B1(n26407), .B2(
        data_in[2]), .ZN(n15800) );
  INV_X1 U11305 ( .A(n15801), .ZN(n20319) );
  AOI22_X1 U11306 ( .A1(\mem[723][3] ), .A2(n15798), .B1(n26407), .B2(
        data_in[3]), .ZN(n15801) );
  INV_X1 U11307 ( .A(n15802), .ZN(n20318) );
  AOI22_X1 U11308 ( .A1(\mem[723][4] ), .A2(n15798), .B1(n26407), .B2(
        data_in[4]), .ZN(n15802) );
  INV_X1 U11309 ( .A(n15803), .ZN(n20317) );
  AOI22_X1 U11310 ( .A1(\mem[723][5] ), .A2(n15798), .B1(n26407), .B2(
        data_in[5]), .ZN(n15803) );
  INV_X1 U11311 ( .A(n15804), .ZN(n20316) );
  AOI22_X1 U11312 ( .A1(\mem[723][6] ), .A2(n15798), .B1(n26407), .B2(
        data_in[6]), .ZN(n15804) );
  INV_X1 U11313 ( .A(n15805), .ZN(n20315) );
  AOI22_X1 U11314 ( .A1(\mem[723][7] ), .A2(n15798), .B1(n26407), .B2(
        data_in[7]), .ZN(n15805) );
  INV_X1 U11315 ( .A(n15806), .ZN(n20314) );
  AOI22_X1 U11316 ( .A1(\mem[724][0] ), .A2(n15807), .B1(n26406), .B2(
        data_in[0]), .ZN(n15806) );
  INV_X1 U11317 ( .A(n15808), .ZN(n20313) );
  AOI22_X1 U11318 ( .A1(\mem[724][1] ), .A2(n15807), .B1(n26406), .B2(
        data_in[1]), .ZN(n15808) );
  INV_X1 U11319 ( .A(n15809), .ZN(n20312) );
  AOI22_X1 U11320 ( .A1(\mem[724][2] ), .A2(n15807), .B1(n26406), .B2(
        data_in[2]), .ZN(n15809) );
  INV_X1 U11321 ( .A(n15810), .ZN(n20311) );
  AOI22_X1 U11322 ( .A1(\mem[724][3] ), .A2(n15807), .B1(n26406), .B2(
        data_in[3]), .ZN(n15810) );
  INV_X1 U11323 ( .A(n15811), .ZN(n20310) );
  AOI22_X1 U11324 ( .A1(\mem[724][4] ), .A2(n15807), .B1(n26406), .B2(
        data_in[4]), .ZN(n15811) );
  INV_X1 U11325 ( .A(n15812), .ZN(n20309) );
  AOI22_X1 U11326 ( .A1(\mem[724][5] ), .A2(n15807), .B1(n26406), .B2(
        data_in[5]), .ZN(n15812) );
  INV_X1 U11327 ( .A(n15813), .ZN(n20308) );
  AOI22_X1 U11328 ( .A1(\mem[724][6] ), .A2(n15807), .B1(n26406), .B2(
        data_in[6]), .ZN(n15813) );
  INV_X1 U11329 ( .A(n15814), .ZN(n20307) );
  AOI22_X1 U11330 ( .A1(\mem[724][7] ), .A2(n15807), .B1(n26406), .B2(
        data_in[7]), .ZN(n15814) );
  INV_X1 U11331 ( .A(n15815), .ZN(n20306) );
  AOI22_X1 U11332 ( .A1(\mem[725][0] ), .A2(n15816), .B1(n26405), .B2(
        data_in[0]), .ZN(n15815) );
  INV_X1 U11333 ( .A(n15817), .ZN(n20305) );
  AOI22_X1 U11334 ( .A1(\mem[725][1] ), .A2(n15816), .B1(n26405), .B2(
        data_in[1]), .ZN(n15817) );
  INV_X1 U11335 ( .A(n15818), .ZN(n20304) );
  AOI22_X1 U11336 ( .A1(\mem[725][2] ), .A2(n15816), .B1(n26405), .B2(
        data_in[2]), .ZN(n15818) );
  INV_X1 U11337 ( .A(n15819), .ZN(n20303) );
  AOI22_X1 U11338 ( .A1(\mem[725][3] ), .A2(n15816), .B1(n26405), .B2(
        data_in[3]), .ZN(n15819) );
  INV_X1 U11339 ( .A(n15820), .ZN(n20302) );
  AOI22_X1 U11340 ( .A1(\mem[725][4] ), .A2(n15816), .B1(n26405), .B2(
        data_in[4]), .ZN(n15820) );
  INV_X1 U11341 ( .A(n15821), .ZN(n20301) );
  AOI22_X1 U11342 ( .A1(\mem[725][5] ), .A2(n15816), .B1(n26405), .B2(
        data_in[5]), .ZN(n15821) );
  INV_X1 U11343 ( .A(n15822), .ZN(n20300) );
  AOI22_X1 U11344 ( .A1(\mem[725][6] ), .A2(n15816), .B1(n26405), .B2(
        data_in[6]), .ZN(n15822) );
  INV_X1 U11345 ( .A(n15823), .ZN(n20299) );
  AOI22_X1 U11346 ( .A1(\mem[725][7] ), .A2(n15816), .B1(n26405), .B2(
        data_in[7]), .ZN(n15823) );
  INV_X1 U11347 ( .A(n15824), .ZN(n20298) );
  AOI22_X1 U11348 ( .A1(\mem[726][0] ), .A2(n15825), .B1(n26404), .B2(
        data_in[0]), .ZN(n15824) );
  INV_X1 U11349 ( .A(n15826), .ZN(n20297) );
  AOI22_X1 U11350 ( .A1(\mem[726][1] ), .A2(n15825), .B1(n26404), .B2(
        data_in[1]), .ZN(n15826) );
  INV_X1 U11351 ( .A(n15827), .ZN(n20296) );
  AOI22_X1 U11352 ( .A1(\mem[726][2] ), .A2(n15825), .B1(n26404), .B2(
        data_in[2]), .ZN(n15827) );
  INV_X1 U11353 ( .A(n15828), .ZN(n20295) );
  AOI22_X1 U11354 ( .A1(\mem[726][3] ), .A2(n15825), .B1(n26404), .B2(
        data_in[3]), .ZN(n15828) );
  INV_X1 U11355 ( .A(n15829), .ZN(n20294) );
  AOI22_X1 U11356 ( .A1(\mem[726][4] ), .A2(n15825), .B1(n26404), .B2(
        data_in[4]), .ZN(n15829) );
  INV_X1 U11357 ( .A(n15830), .ZN(n20293) );
  AOI22_X1 U11358 ( .A1(\mem[726][5] ), .A2(n15825), .B1(n26404), .B2(
        data_in[5]), .ZN(n15830) );
  INV_X1 U11359 ( .A(n15831), .ZN(n20292) );
  AOI22_X1 U11360 ( .A1(\mem[726][6] ), .A2(n15825), .B1(n26404), .B2(
        data_in[6]), .ZN(n15831) );
  INV_X1 U11361 ( .A(n15832), .ZN(n20291) );
  AOI22_X1 U11362 ( .A1(\mem[726][7] ), .A2(n15825), .B1(n26404), .B2(
        data_in[7]), .ZN(n15832) );
  INV_X1 U11363 ( .A(n15833), .ZN(n20290) );
  AOI22_X1 U11364 ( .A1(\mem[727][0] ), .A2(n15834), .B1(n26403), .B2(
        data_in[0]), .ZN(n15833) );
  INV_X1 U11365 ( .A(n15835), .ZN(n20289) );
  AOI22_X1 U11366 ( .A1(\mem[727][1] ), .A2(n15834), .B1(n26403), .B2(
        data_in[1]), .ZN(n15835) );
  INV_X1 U11367 ( .A(n15836), .ZN(n20288) );
  AOI22_X1 U11368 ( .A1(\mem[727][2] ), .A2(n15834), .B1(n26403), .B2(
        data_in[2]), .ZN(n15836) );
  INV_X1 U11369 ( .A(n15837), .ZN(n20287) );
  AOI22_X1 U11370 ( .A1(\mem[727][3] ), .A2(n15834), .B1(n26403), .B2(
        data_in[3]), .ZN(n15837) );
  INV_X1 U11371 ( .A(n15838), .ZN(n20286) );
  AOI22_X1 U11372 ( .A1(\mem[727][4] ), .A2(n15834), .B1(n26403), .B2(
        data_in[4]), .ZN(n15838) );
  INV_X1 U11373 ( .A(n15839), .ZN(n20285) );
  AOI22_X1 U11374 ( .A1(\mem[727][5] ), .A2(n15834), .B1(n26403), .B2(
        data_in[5]), .ZN(n15839) );
  INV_X1 U11375 ( .A(n15840), .ZN(n20284) );
  AOI22_X1 U11376 ( .A1(\mem[727][6] ), .A2(n15834), .B1(n26403), .B2(
        data_in[6]), .ZN(n15840) );
  INV_X1 U11377 ( .A(n15841), .ZN(n20283) );
  AOI22_X1 U11378 ( .A1(\mem[727][7] ), .A2(n15834), .B1(n26403), .B2(
        data_in[7]), .ZN(n15841) );
  INV_X1 U11379 ( .A(n15842), .ZN(n20282) );
  AOI22_X1 U11380 ( .A1(\mem[728][0] ), .A2(n15843), .B1(n26402), .B2(
        data_in[0]), .ZN(n15842) );
  INV_X1 U11381 ( .A(n15844), .ZN(n20281) );
  AOI22_X1 U11382 ( .A1(\mem[728][1] ), .A2(n15843), .B1(n26402), .B2(
        data_in[1]), .ZN(n15844) );
  INV_X1 U11383 ( .A(n15845), .ZN(n20280) );
  AOI22_X1 U11384 ( .A1(\mem[728][2] ), .A2(n15843), .B1(n26402), .B2(
        data_in[2]), .ZN(n15845) );
  INV_X1 U11385 ( .A(n15846), .ZN(n20279) );
  AOI22_X1 U11386 ( .A1(\mem[728][3] ), .A2(n15843), .B1(n26402), .B2(
        data_in[3]), .ZN(n15846) );
  INV_X1 U11387 ( .A(n15847), .ZN(n20278) );
  AOI22_X1 U11388 ( .A1(\mem[728][4] ), .A2(n15843), .B1(n26402), .B2(
        data_in[4]), .ZN(n15847) );
  INV_X1 U11389 ( .A(n15848), .ZN(n20277) );
  AOI22_X1 U11390 ( .A1(\mem[728][5] ), .A2(n15843), .B1(n26402), .B2(
        data_in[5]), .ZN(n15848) );
  INV_X1 U11391 ( .A(n15849), .ZN(n20276) );
  AOI22_X1 U11392 ( .A1(\mem[728][6] ), .A2(n15843), .B1(n26402), .B2(
        data_in[6]), .ZN(n15849) );
  INV_X1 U11393 ( .A(n15850), .ZN(n20275) );
  AOI22_X1 U11394 ( .A1(\mem[728][7] ), .A2(n15843), .B1(n26402), .B2(
        data_in[7]), .ZN(n15850) );
  INV_X1 U11395 ( .A(n15851), .ZN(n20274) );
  AOI22_X1 U11396 ( .A1(\mem[729][0] ), .A2(n15852), .B1(n26401), .B2(
        data_in[0]), .ZN(n15851) );
  INV_X1 U11397 ( .A(n15853), .ZN(n20273) );
  AOI22_X1 U11398 ( .A1(\mem[729][1] ), .A2(n15852), .B1(n26401), .B2(
        data_in[1]), .ZN(n15853) );
  INV_X1 U11399 ( .A(n15854), .ZN(n20272) );
  AOI22_X1 U11400 ( .A1(\mem[729][2] ), .A2(n15852), .B1(n26401), .B2(
        data_in[2]), .ZN(n15854) );
  INV_X1 U11401 ( .A(n15855), .ZN(n20271) );
  AOI22_X1 U11402 ( .A1(\mem[729][3] ), .A2(n15852), .B1(n26401), .B2(
        data_in[3]), .ZN(n15855) );
  INV_X1 U11403 ( .A(n15856), .ZN(n20270) );
  AOI22_X1 U11404 ( .A1(\mem[729][4] ), .A2(n15852), .B1(n26401), .B2(
        data_in[4]), .ZN(n15856) );
  INV_X1 U11405 ( .A(n15857), .ZN(n20269) );
  AOI22_X1 U11406 ( .A1(\mem[729][5] ), .A2(n15852), .B1(n26401), .B2(
        data_in[5]), .ZN(n15857) );
  INV_X1 U11407 ( .A(n15858), .ZN(n20268) );
  AOI22_X1 U11408 ( .A1(\mem[729][6] ), .A2(n15852), .B1(n26401), .B2(
        data_in[6]), .ZN(n15858) );
  INV_X1 U11409 ( .A(n15859), .ZN(n20267) );
  AOI22_X1 U11410 ( .A1(\mem[729][7] ), .A2(n15852), .B1(n26401), .B2(
        data_in[7]), .ZN(n15859) );
  INV_X1 U11411 ( .A(n15860), .ZN(n20266) );
  AOI22_X1 U11412 ( .A1(\mem[730][0] ), .A2(n15861), .B1(n26400), .B2(
        data_in[0]), .ZN(n15860) );
  INV_X1 U11413 ( .A(n15862), .ZN(n20265) );
  AOI22_X1 U11414 ( .A1(\mem[730][1] ), .A2(n15861), .B1(n26400), .B2(
        data_in[1]), .ZN(n15862) );
  INV_X1 U11415 ( .A(n15863), .ZN(n20264) );
  AOI22_X1 U11416 ( .A1(\mem[730][2] ), .A2(n15861), .B1(n26400), .B2(
        data_in[2]), .ZN(n15863) );
  INV_X1 U11417 ( .A(n15864), .ZN(n20263) );
  AOI22_X1 U11418 ( .A1(\mem[730][3] ), .A2(n15861), .B1(n26400), .B2(
        data_in[3]), .ZN(n15864) );
  INV_X1 U11419 ( .A(n15865), .ZN(n20262) );
  AOI22_X1 U11420 ( .A1(\mem[730][4] ), .A2(n15861), .B1(n26400), .B2(
        data_in[4]), .ZN(n15865) );
  INV_X1 U11421 ( .A(n15866), .ZN(n20261) );
  AOI22_X1 U11422 ( .A1(\mem[730][5] ), .A2(n15861), .B1(n26400), .B2(
        data_in[5]), .ZN(n15866) );
  INV_X1 U11423 ( .A(n15867), .ZN(n20260) );
  AOI22_X1 U11424 ( .A1(\mem[730][6] ), .A2(n15861), .B1(n26400), .B2(
        data_in[6]), .ZN(n15867) );
  INV_X1 U11425 ( .A(n15868), .ZN(n20259) );
  AOI22_X1 U11426 ( .A1(\mem[730][7] ), .A2(n15861), .B1(n26400), .B2(
        data_in[7]), .ZN(n15868) );
  INV_X1 U11427 ( .A(n15869), .ZN(n20258) );
  AOI22_X1 U11428 ( .A1(\mem[731][0] ), .A2(n15870), .B1(n26399), .B2(
        data_in[0]), .ZN(n15869) );
  INV_X1 U11429 ( .A(n15871), .ZN(n20257) );
  AOI22_X1 U11430 ( .A1(\mem[731][1] ), .A2(n15870), .B1(n26399), .B2(
        data_in[1]), .ZN(n15871) );
  INV_X1 U11431 ( .A(n15872), .ZN(n20256) );
  AOI22_X1 U11432 ( .A1(\mem[731][2] ), .A2(n15870), .B1(n26399), .B2(
        data_in[2]), .ZN(n15872) );
  INV_X1 U11433 ( .A(n15873), .ZN(n20255) );
  AOI22_X1 U11434 ( .A1(\mem[731][3] ), .A2(n15870), .B1(n26399), .B2(
        data_in[3]), .ZN(n15873) );
  INV_X1 U11435 ( .A(n15874), .ZN(n20254) );
  AOI22_X1 U11436 ( .A1(\mem[731][4] ), .A2(n15870), .B1(n26399), .B2(
        data_in[4]), .ZN(n15874) );
  INV_X1 U11437 ( .A(n15875), .ZN(n20253) );
  AOI22_X1 U11438 ( .A1(\mem[731][5] ), .A2(n15870), .B1(n26399), .B2(
        data_in[5]), .ZN(n15875) );
  INV_X1 U11439 ( .A(n15876), .ZN(n20252) );
  AOI22_X1 U11440 ( .A1(\mem[731][6] ), .A2(n15870), .B1(n26399), .B2(
        data_in[6]), .ZN(n15876) );
  INV_X1 U11441 ( .A(n15877), .ZN(n20251) );
  AOI22_X1 U11442 ( .A1(\mem[731][7] ), .A2(n15870), .B1(n26399), .B2(
        data_in[7]), .ZN(n15877) );
  INV_X1 U11443 ( .A(n15878), .ZN(n20250) );
  AOI22_X1 U11444 ( .A1(\mem[732][0] ), .A2(n15879), .B1(n26398), .B2(
        data_in[0]), .ZN(n15878) );
  INV_X1 U11445 ( .A(n15880), .ZN(n20249) );
  AOI22_X1 U11446 ( .A1(\mem[732][1] ), .A2(n15879), .B1(n26398), .B2(
        data_in[1]), .ZN(n15880) );
  INV_X1 U11447 ( .A(n15881), .ZN(n20248) );
  AOI22_X1 U11448 ( .A1(\mem[732][2] ), .A2(n15879), .B1(n26398), .B2(
        data_in[2]), .ZN(n15881) );
  INV_X1 U11449 ( .A(n15882), .ZN(n20247) );
  AOI22_X1 U11450 ( .A1(\mem[732][3] ), .A2(n15879), .B1(n26398), .B2(
        data_in[3]), .ZN(n15882) );
  INV_X1 U11451 ( .A(n15883), .ZN(n20246) );
  AOI22_X1 U11452 ( .A1(\mem[732][4] ), .A2(n15879), .B1(n26398), .B2(
        data_in[4]), .ZN(n15883) );
  INV_X1 U11453 ( .A(n15884), .ZN(n20245) );
  AOI22_X1 U11454 ( .A1(\mem[732][5] ), .A2(n15879), .B1(n26398), .B2(
        data_in[5]), .ZN(n15884) );
  INV_X1 U11455 ( .A(n15885), .ZN(n20244) );
  AOI22_X1 U11456 ( .A1(\mem[732][6] ), .A2(n15879), .B1(n26398), .B2(
        data_in[6]), .ZN(n15885) );
  INV_X1 U11457 ( .A(n15886), .ZN(n20243) );
  AOI22_X1 U11458 ( .A1(\mem[732][7] ), .A2(n15879), .B1(n26398), .B2(
        data_in[7]), .ZN(n15886) );
  INV_X1 U11459 ( .A(n15887), .ZN(n20242) );
  AOI22_X1 U11460 ( .A1(\mem[733][0] ), .A2(n15888), .B1(n26397), .B2(
        data_in[0]), .ZN(n15887) );
  INV_X1 U11461 ( .A(n15889), .ZN(n20241) );
  AOI22_X1 U11462 ( .A1(\mem[733][1] ), .A2(n15888), .B1(n26397), .B2(
        data_in[1]), .ZN(n15889) );
  INV_X1 U11463 ( .A(n15890), .ZN(n20240) );
  AOI22_X1 U11464 ( .A1(\mem[733][2] ), .A2(n15888), .B1(n26397), .B2(
        data_in[2]), .ZN(n15890) );
  INV_X1 U11465 ( .A(n15891), .ZN(n20239) );
  AOI22_X1 U11466 ( .A1(\mem[733][3] ), .A2(n15888), .B1(n26397), .B2(
        data_in[3]), .ZN(n15891) );
  INV_X1 U11467 ( .A(n15892), .ZN(n20238) );
  AOI22_X1 U11468 ( .A1(\mem[733][4] ), .A2(n15888), .B1(n26397), .B2(
        data_in[4]), .ZN(n15892) );
  INV_X1 U11469 ( .A(n15893), .ZN(n20237) );
  AOI22_X1 U11470 ( .A1(\mem[733][5] ), .A2(n15888), .B1(n26397), .B2(
        data_in[5]), .ZN(n15893) );
  INV_X1 U11471 ( .A(n15894), .ZN(n20236) );
  AOI22_X1 U11472 ( .A1(\mem[733][6] ), .A2(n15888), .B1(n26397), .B2(
        data_in[6]), .ZN(n15894) );
  INV_X1 U11473 ( .A(n15895), .ZN(n20235) );
  AOI22_X1 U11474 ( .A1(\mem[733][7] ), .A2(n15888), .B1(n26397), .B2(
        data_in[7]), .ZN(n15895) );
  INV_X1 U11475 ( .A(n15896), .ZN(n20234) );
  AOI22_X1 U11476 ( .A1(\mem[734][0] ), .A2(n15897), .B1(n26396), .B2(
        data_in[0]), .ZN(n15896) );
  INV_X1 U11477 ( .A(n15898), .ZN(n20233) );
  AOI22_X1 U11478 ( .A1(\mem[734][1] ), .A2(n15897), .B1(n26396), .B2(
        data_in[1]), .ZN(n15898) );
  INV_X1 U11479 ( .A(n15899), .ZN(n20232) );
  AOI22_X1 U11480 ( .A1(\mem[734][2] ), .A2(n15897), .B1(n26396), .B2(
        data_in[2]), .ZN(n15899) );
  INV_X1 U11481 ( .A(n15900), .ZN(n20231) );
  AOI22_X1 U11482 ( .A1(\mem[734][3] ), .A2(n15897), .B1(n26396), .B2(
        data_in[3]), .ZN(n15900) );
  INV_X1 U11483 ( .A(n15901), .ZN(n20230) );
  AOI22_X1 U11484 ( .A1(\mem[734][4] ), .A2(n15897), .B1(n26396), .B2(
        data_in[4]), .ZN(n15901) );
  INV_X1 U11485 ( .A(n15902), .ZN(n20229) );
  AOI22_X1 U11486 ( .A1(\mem[734][5] ), .A2(n15897), .B1(n26396), .B2(
        data_in[5]), .ZN(n15902) );
  INV_X1 U11487 ( .A(n15903), .ZN(n20228) );
  AOI22_X1 U11488 ( .A1(\mem[734][6] ), .A2(n15897), .B1(n26396), .B2(
        data_in[6]), .ZN(n15903) );
  INV_X1 U11489 ( .A(n15904), .ZN(n20227) );
  AOI22_X1 U11490 ( .A1(\mem[734][7] ), .A2(n15897), .B1(n26396), .B2(
        data_in[7]), .ZN(n15904) );
  INV_X1 U11491 ( .A(n15905), .ZN(n20226) );
  AOI22_X1 U11492 ( .A1(\mem[735][0] ), .A2(n15906), .B1(n26395), .B2(
        data_in[0]), .ZN(n15905) );
  INV_X1 U11493 ( .A(n15907), .ZN(n20225) );
  AOI22_X1 U11494 ( .A1(\mem[735][1] ), .A2(n15906), .B1(n26395), .B2(
        data_in[1]), .ZN(n15907) );
  INV_X1 U11495 ( .A(n15908), .ZN(n20224) );
  AOI22_X1 U11496 ( .A1(\mem[735][2] ), .A2(n15906), .B1(n26395), .B2(
        data_in[2]), .ZN(n15908) );
  INV_X1 U11497 ( .A(n15909), .ZN(n20223) );
  AOI22_X1 U11498 ( .A1(\mem[735][3] ), .A2(n15906), .B1(n26395), .B2(
        data_in[3]), .ZN(n15909) );
  INV_X1 U11499 ( .A(n15910), .ZN(n20222) );
  AOI22_X1 U11500 ( .A1(\mem[735][4] ), .A2(n15906), .B1(n26395), .B2(
        data_in[4]), .ZN(n15910) );
  INV_X1 U11501 ( .A(n15911), .ZN(n20221) );
  AOI22_X1 U11502 ( .A1(\mem[735][5] ), .A2(n15906), .B1(n26395), .B2(
        data_in[5]), .ZN(n15911) );
  INV_X1 U11503 ( .A(n15912), .ZN(n20220) );
  AOI22_X1 U11504 ( .A1(\mem[735][6] ), .A2(n15906), .B1(n26395), .B2(
        data_in[6]), .ZN(n15912) );
  INV_X1 U11505 ( .A(n15913), .ZN(n20219) );
  AOI22_X1 U11506 ( .A1(\mem[735][7] ), .A2(n15906), .B1(n26395), .B2(
        data_in[7]), .ZN(n15913) );
  INV_X1 U11507 ( .A(n15987), .ZN(n20154) );
  AOI22_X1 U11508 ( .A1(\mem[744][0] ), .A2(n15988), .B1(n26386), .B2(
        data_in[0]), .ZN(n15987) );
  INV_X1 U11509 ( .A(n15989), .ZN(n20153) );
  AOI22_X1 U11510 ( .A1(\mem[744][1] ), .A2(n15988), .B1(n26386), .B2(
        data_in[1]), .ZN(n15989) );
  INV_X1 U11511 ( .A(n15990), .ZN(n20152) );
  AOI22_X1 U11512 ( .A1(\mem[744][2] ), .A2(n15988), .B1(n26386), .B2(
        data_in[2]), .ZN(n15990) );
  INV_X1 U11513 ( .A(n15991), .ZN(n20151) );
  AOI22_X1 U11514 ( .A1(\mem[744][3] ), .A2(n15988), .B1(n26386), .B2(
        data_in[3]), .ZN(n15991) );
  INV_X1 U11515 ( .A(n15992), .ZN(n20150) );
  AOI22_X1 U11516 ( .A1(\mem[744][4] ), .A2(n15988), .B1(n26386), .B2(
        data_in[4]), .ZN(n15992) );
  INV_X1 U11517 ( .A(n15993), .ZN(n20149) );
  AOI22_X1 U11518 ( .A1(\mem[744][5] ), .A2(n15988), .B1(n26386), .B2(
        data_in[5]), .ZN(n15993) );
  INV_X1 U11519 ( .A(n15994), .ZN(n20148) );
  AOI22_X1 U11520 ( .A1(\mem[744][6] ), .A2(n15988), .B1(n26386), .B2(
        data_in[6]), .ZN(n15994) );
  INV_X1 U11521 ( .A(n15995), .ZN(n20147) );
  AOI22_X1 U11522 ( .A1(\mem[744][7] ), .A2(n15988), .B1(n26386), .B2(
        data_in[7]), .ZN(n15995) );
  INV_X1 U11523 ( .A(n15996), .ZN(n20146) );
  AOI22_X1 U11524 ( .A1(\mem[745][0] ), .A2(n15997), .B1(n26385), .B2(
        data_in[0]), .ZN(n15996) );
  INV_X1 U11525 ( .A(n15998), .ZN(n20145) );
  AOI22_X1 U11526 ( .A1(\mem[745][1] ), .A2(n15997), .B1(n26385), .B2(
        data_in[1]), .ZN(n15998) );
  INV_X1 U11527 ( .A(n15999), .ZN(n20144) );
  AOI22_X1 U11528 ( .A1(\mem[745][2] ), .A2(n15997), .B1(n26385), .B2(
        data_in[2]), .ZN(n15999) );
  INV_X1 U11529 ( .A(n16000), .ZN(n20143) );
  AOI22_X1 U11530 ( .A1(\mem[745][3] ), .A2(n15997), .B1(n26385), .B2(
        data_in[3]), .ZN(n16000) );
  INV_X1 U11531 ( .A(n16001), .ZN(n20142) );
  AOI22_X1 U11532 ( .A1(\mem[745][4] ), .A2(n15997), .B1(n26385), .B2(
        data_in[4]), .ZN(n16001) );
  INV_X1 U11533 ( .A(n16002), .ZN(n20141) );
  AOI22_X1 U11534 ( .A1(\mem[745][5] ), .A2(n15997), .B1(n26385), .B2(
        data_in[5]), .ZN(n16002) );
  INV_X1 U11535 ( .A(n16003), .ZN(n20140) );
  AOI22_X1 U11536 ( .A1(\mem[745][6] ), .A2(n15997), .B1(n26385), .B2(
        data_in[6]), .ZN(n16003) );
  INV_X1 U11537 ( .A(n16004), .ZN(n20139) );
  AOI22_X1 U11538 ( .A1(\mem[745][7] ), .A2(n15997), .B1(n26385), .B2(
        data_in[7]), .ZN(n16004) );
  INV_X1 U11539 ( .A(n16005), .ZN(n20138) );
  AOI22_X1 U11540 ( .A1(\mem[746][0] ), .A2(n16006), .B1(n26384), .B2(
        data_in[0]), .ZN(n16005) );
  INV_X1 U11541 ( .A(n16007), .ZN(n20137) );
  AOI22_X1 U11542 ( .A1(\mem[746][1] ), .A2(n16006), .B1(n26384), .B2(
        data_in[1]), .ZN(n16007) );
  INV_X1 U11543 ( .A(n16008), .ZN(n20136) );
  AOI22_X1 U11544 ( .A1(\mem[746][2] ), .A2(n16006), .B1(n26384), .B2(
        data_in[2]), .ZN(n16008) );
  INV_X1 U11545 ( .A(n16009), .ZN(n20135) );
  AOI22_X1 U11546 ( .A1(\mem[746][3] ), .A2(n16006), .B1(n26384), .B2(
        data_in[3]), .ZN(n16009) );
  INV_X1 U11547 ( .A(n16010), .ZN(n20134) );
  AOI22_X1 U11548 ( .A1(\mem[746][4] ), .A2(n16006), .B1(n26384), .B2(
        data_in[4]), .ZN(n16010) );
  INV_X1 U11549 ( .A(n16011), .ZN(n20133) );
  AOI22_X1 U11550 ( .A1(\mem[746][5] ), .A2(n16006), .B1(n26384), .B2(
        data_in[5]), .ZN(n16011) );
  INV_X1 U11551 ( .A(n16012), .ZN(n20132) );
  AOI22_X1 U11552 ( .A1(\mem[746][6] ), .A2(n16006), .B1(n26384), .B2(
        data_in[6]), .ZN(n16012) );
  INV_X1 U11553 ( .A(n16013), .ZN(n20131) );
  AOI22_X1 U11554 ( .A1(\mem[746][7] ), .A2(n16006), .B1(n26384), .B2(
        data_in[7]), .ZN(n16013) );
  INV_X1 U11555 ( .A(n16014), .ZN(n20130) );
  AOI22_X1 U11556 ( .A1(\mem[747][0] ), .A2(n16015), .B1(n26383), .B2(
        data_in[0]), .ZN(n16014) );
  INV_X1 U11557 ( .A(n16016), .ZN(n20129) );
  AOI22_X1 U11558 ( .A1(\mem[747][1] ), .A2(n16015), .B1(n26383), .B2(
        data_in[1]), .ZN(n16016) );
  INV_X1 U11559 ( .A(n16017), .ZN(n20128) );
  AOI22_X1 U11560 ( .A1(\mem[747][2] ), .A2(n16015), .B1(n26383), .B2(
        data_in[2]), .ZN(n16017) );
  INV_X1 U11561 ( .A(n16018), .ZN(n20127) );
  AOI22_X1 U11562 ( .A1(\mem[747][3] ), .A2(n16015), .B1(n26383), .B2(
        data_in[3]), .ZN(n16018) );
  INV_X1 U11563 ( .A(n16019), .ZN(n20126) );
  AOI22_X1 U11564 ( .A1(\mem[747][4] ), .A2(n16015), .B1(n26383), .B2(
        data_in[4]), .ZN(n16019) );
  INV_X1 U11565 ( .A(n16020), .ZN(n20125) );
  AOI22_X1 U11566 ( .A1(\mem[747][5] ), .A2(n16015), .B1(n26383), .B2(
        data_in[5]), .ZN(n16020) );
  INV_X1 U11567 ( .A(n16021), .ZN(n20124) );
  AOI22_X1 U11568 ( .A1(\mem[747][6] ), .A2(n16015), .B1(n26383), .B2(
        data_in[6]), .ZN(n16021) );
  INV_X1 U11569 ( .A(n16022), .ZN(n20123) );
  AOI22_X1 U11570 ( .A1(\mem[747][7] ), .A2(n16015), .B1(n26383), .B2(
        data_in[7]), .ZN(n16022) );
  INV_X1 U11571 ( .A(n16023), .ZN(n20122) );
  AOI22_X1 U11572 ( .A1(\mem[748][0] ), .A2(n16024), .B1(n26382), .B2(
        data_in[0]), .ZN(n16023) );
  INV_X1 U11573 ( .A(n16025), .ZN(n20121) );
  AOI22_X1 U11574 ( .A1(\mem[748][1] ), .A2(n16024), .B1(n26382), .B2(
        data_in[1]), .ZN(n16025) );
  INV_X1 U11575 ( .A(n16026), .ZN(n20120) );
  AOI22_X1 U11576 ( .A1(\mem[748][2] ), .A2(n16024), .B1(n26382), .B2(
        data_in[2]), .ZN(n16026) );
  INV_X1 U11577 ( .A(n16027), .ZN(n20119) );
  AOI22_X1 U11578 ( .A1(\mem[748][3] ), .A2(n16024), .B1(n26382), .B2(
        data_in[3]), .ZN(n16027) );
  INV_X1 U11579 ( .A(n16028), .ZN(n20118) );
  AOI22_X1 U11580 ( .A1(\mem[748][4] ), .A2(n16024), .B1(n26382), .B2(
        data_in[4]), .ZN(n16028) );
  INV_X1 U11581 ( .A(n16029), .ZN(n20117) );
  AOI22_X1 U11582 ( .A1(\mem[748][5] ), .A2(n16024), .B1(n26382), .B2(
        data_in[5]), .ZN(n16029) );
  INV_X1 U11583 ( .A(n16030), .ZN(n20116) );
  AOI22_X1 U11584 ( .A1(\mem[748][6] ), .A2(n16024), .B1(n26382), .B2(
        data_in[6]), .ZN(n16030) );
  INV_X1 U11585 ( .A(n16031), .ZN(n20115) );
  AOI22_X1 U11586 ( .A1(\mem[748][7] ), .A2(n16024), .B1(n26382), .B2(
        data_in[7]), .ZN(n16031) );
  INV_X1 U11587 ( .A(n16032), .ZN(n20114) );
  AOI22_X1 U11588 ( .A1(\mem[749][0] ), .A2(n16033), .B1(n26381), .B2(
        data_in[0]), .ZN(n16032) );
  INV_X1 U11589 ( .A(n16034), .ZN(n20113) );
  AOI22_X1 U11590 ( .A1(\mem[749][1] ), .A2(n16033), .B1(n26381), .B2(
        data_in[1]), .ZN(n16034) );
  INV_X1 U11591 ( .A(n16035), .ZN(n20112) );
  AOI22_X1 U11592 ( .A1(\mem[749][2] ), .A2(n16033), .B1(n26381), .B2(
        data_in[2]), .ZN(n16035) );
  INV_X1 U11593 ( .A(n16036), .ZN(n20111) );
  AOI22_X1 U11594 ( .A1(\mem[749][3] ), .A2(n16033), .B1(n26381), .B2(
        data_in[3]), .ZN(n16036) );
  INV_X1 U11595 ( .A(n16037), .ZN(n20110) );
  AOI22_X1 U11596 ( .A1(\mem[749][4] ), .A2(n16033), .B1(n26381), .B2(
        data_in[4]), .ZN(n16037) );
  INV_X1 U11597 ( .A(n16038), .ZN(n20109) );
  AOI22_X1 U11598 ( .A1(\mem[749][5] ), .A2(n16033), .B1(n26381), .B2(
        data_in[5]), .ZN(n16038) );
  INV_X1 U11599 ( .A(n16039), .ZN(n20108) );
  AOI22_X1 U11600 ( .A1(\mem[749][6] ), .A2(n16033), .B1(n26381), .B2(
        data_in[6]), .ZN(n16039) );
  INV_X1 U11601 ( .A(n16040), .ZN(n20107) );
  AOI22_X1 U11602 ( .A1(\mem[749][7] ), .A2(n16033), .B1(n26381), .B2(
        data_in[7]), .ZN(n16040) );
  INV_X1 U11603 ( .A(n16041), .ZN(n20106) );
  AOI22_X1 U11604 ( .A1(\mem[750][0] ), .A2(n16042), .B1(n26380), .B2(
        data_in[0]), .ZN(n16041) );
  INV_X1 U11605 ( .A(n16043), .ZN(n20105) );
  AOI22_X1 U11606 ( .A1(\mem[750][1] ), .A2(n16042), .B1(n26380), .B2(
        data_in[1]), .ZN(n16043) );
  INV_X1 U11607 ( .A(n16044), .ZN(n20104) );
  AOI22_X1 U11608 ( .A1(\mem[750][2] ), .A2(n16042), .B1(n26380), .B2(
        data_in[2]), .ZN(n16044) );
  INV_X1 U11609 ( .A(n16045), .ZN(n20103) );
  AOI22_X1 U11610 ( .A1(\mem[750][3] ), .A2(n16042), .B1(n26380), .B2(
        data_in[3]), .ZN(n16045) );
  INV_X1 U11611 ( .A(n16046), .ZN(n20102) );
  AOI22_X1 U11612 ( .A1(\mem[750][4] ), .A2(n16042), .B1(n26380), .B2(
        data_in[4]), .ZN(n16046) );
  INV_X1 U11613 ( .A(n16047), .ZN(n20101) );
  AOI22_X1 U11614 ( .A1(\mem[750][5] ), .A2(n16042), .B1(n26380), .B2(
        data_in[5]), .ZN(n16047) );
  INV_X1 U11615 ( .A(n16048), .ZN(n20100) );
  AOI22_X1 U11616 ( .A1(\mem[750][6] ), .A2(n16042), .B1(n26380), .B2(
        data_in[6]), .ZN(n16048) );
  INV_X1 U11617 ( .A(n16049), .ZN(n20099) );
  AOI22_X1 U11618 ( .A1(\mem[750][7] ), .A2(n16042), .B1(n26380), .B2(
        data_in[7]), .ZN(n16049) );
  INV_X1 U11619 ( .A(n16050), .ZN(n20098) );
  AOI22_X1 U11620 ( .A1(\mem[751][0] ), .A2(n16051), .B1(n26379), .B2(
        data_in[0]), .ZN(n16050) );
  INV_X1 U11621 ( .A(n16052), .ZN(n20097) );
  AOI22_X1 U11622 ( .A1(\mem[751][1] ), .A2(n16051), .B1(n26379), .B2(
        data_in[1]), .ZN(n16052) );
  INV_X1 U11623 ( .A(n16053), .ZN(n20096) );
  AOI22_X1 U11624 ( .A1(\mem[751][2] ), .A2(n16051), .B1(n26379), .B2(
        data_in[2]), .ZN(n16053) );
  INV_X1 U11625 ( .A(n16054), .ZN(n20095) );
  AOI22_X1 U11626 ( .A1(\mem[751][3] ), .A2(n16051), .B1(n26379), .B2(
        data_in[3]), .ZN(n16054) );
  INV_X1 U11627 ( .A(n16055), .ZN(n20094) );
  AOI22_X1 U11628 ( .A1(\mem[751][4] ), .A2(n16051), .B1(n26379), .B2(
        data_in[4]), .ZN(n16055) );
  INV_X1 U11629 ( .A(n16056), .ZN(n20093) );
  AOI22_X1 U11630 ( .A1(\mem[751][5] ), .A2(n16051), .B1(n26379), .B2(
        data_in[5]), .ZN(n16056) );
  INV_X1 U11631 ( .A(n16057), .ZN(n20092) );
  AOI22_X1 U11632 ( .A1(\mem[751][6] ), .A2(n16051), .B1(n26379), .B2(
        data_in[6]), .ZN(n16057) );
  INV_X1 U11633 ( .A(n16058), .ZN(n20091) );
  AOI22_X1 U11634 ( .A1(\mem[751][7] ), .A2(n16051), .B1(n26379), .B2(
        data_in[7]), .ZN(n16058) );
  INV_X1 U11635 ( .A(n16059), .ZN(n20090) );
  AOI22_X1 U11636 ( .A1(\mem[752][0] ), .A2(n16060), .B1(n26378), .B2(
        data_in[0]), .ZN(n16059) );
  INV_X1 U11637 ( .A(n16061), .ZN(n20089) );
  AOI22_X1 U11638 ( .A1(\mem[752][1] ), .A2(n16060), .B1(n26378), .B2(
        data_in[1]), .ZN(n16061) );
  INV_X1 U11639 ( .A(n16062), .ZN(n20088) );
  AOI22_X1 U11640 ( .A1(\mem[752][2] ), .A2(n16060), .B1(n26378), .B2(
        data_in[2]), .ZN(n16062) );
  INV_X1 U11641 ( .A(n16063), .ZN(n20087) );
  AOI22_X1 U11642 ( .A1(\mem[752][3] ), .A2(n16060), .B1(n26378), .B2(
        data_in[3]), .ZN(n16063) );
  INV_X1 U11643 ( .A(n16064), .ZN(n20086) );
  AOI22_X1 U11644 ( .A1(\mem[752][4] ), .A2(n16060), .B1(n26378), .B2(
        data_in[4]), .ZN(n16064) );
  INV_X1 U11645 ( .A(n16065), .ZN(n20085) );
  AOI22_X1 U11646 ( .A1(\mem[752][5] ), .A2(n16060), .B1(n26378), .B2(
        data_in[5]), .ZN(n16065) );
  INV_X1 U11647 ( .A(n16066), .ZN(n20084) );
  AOI22_X1 U11648 ( .A1(\mem[752][6] ), .A2(n16060), .B1(n26378), .B2(
        data_in[6]), .ZN(n16066) );
  INV_X1 U11649 ( .A(n16067), .ZN(n20083) );
  AOI22_X1 U11650 ( .A1(\mem[752][7] ), .A2(n16060), .B1(n26378), .B2(
        data_in[7]), .ZN(n16067) );
  INV_X1 U11651 ( .A(n16068), .ZN(n20082) );
  AOI22_X1 U11652 ( .A1(\mem[753][0] ), .A2(n16069), .B1(n26377), .B2(
        data_in[0]), .ZN(n16068) );
  INV_X1 U11653 ( .A(n16070), .ZN(n20081) );
  AOI22_X1 U11654 ( .A1(\mem[753][1] ), .A2(n16069), .B1(n26377), .B2(
        data_in[1]), .ZN(n16070) );
  INV_X1 U11655 ( .A(n16071), .ZN(n20080) );
  AOI22_X1 U11656 ( .A1(\mem[753][2] ), .A2(n16069), .B1(n26377), .B2(
        data_in[2]), .ZN(n16071) );
  INV_X1 U11657 ( .A(n16072), .ZN(n20079) );
  AOI22_X1 U11658 ( .A1(\mem[753][3] ), .A2(n16069), .B1(n26377), .B2(
        data_in[3]), .ZN(n16072) );
  INV_X1 U11659 ( .A(n16073), .ZN(n20078) );
  AOI22_X1 U11660 ( .A1(\mem[753][4] ), .A2(n16069), .B1(n26377), .B2(
        data_in[4]), .ZN(n16073) );
  INV_X1 U11661 ( .A(n16074), .ZN(n20077) );
  AOI22_X1 U11662 ( .A1(\mem[753][5] ), .A2(n16069), .B1(n26377), .B2(
        data_in[5]), .ZN(n16074) );
  INV_X1 U11663 ( .A(n16075), .ZN(n20076) );
  AOI22_X1 U11664 ( .A1(\mem[753][6] ), .A2(n16069), .B1(n26377), .B2(
        data_in[6]), .ZN(n16075) );
  INV_X1 U11665 ( .A(n16076), .ZN(n20075) );
  AOI22_X1 U11666 ( .A1(\mem[753][7] ), .A2(n16069), .B1(n26377), .B2(
        data_in[7]), .ZN(n16076) );
  INV_X1 U11667 ( .A(n16077), .ZN(n20074) );
  AOI22_X1 U11668 ( .A1(\mem[754][0] ), .A2(n16078), .B1(n26376), .B2(
        data_in[0]), .ZN(n16077) );
  INV_X1 U11669 ( .A(n16079), .ZN(n20073) );
  AOI22_X1 U11670 ( .A1(\mem[754][1] ), .A2(n16078), .B1(n26376), .B2(
        data_in[1]), .ZN(n16079) );
  INV_X1 U11671 ( .A(n16080), .ZN(n20072) );
  AOI22_X1 U11672 ( .A1(\mem[754][2] ), .A2(n16078), .B1(n26376), .B2(
        data_in[2]), .ZN(n16080) );
  INV_X1 U11673 ( .A(n16081), .ZN(n20071) );
  AOI22_X1 U11674 ( .A1(\mem[754][3] ), .A2(n16078), .B1(n26376), .B2(
        data_in[3]), .ZN(n16081) );
  INV_X1 U11675 ( .A(n16082), .ZN(n20070) );
  AOI22_X1 U11676 ( .A1(\mem[754][4] ), .A2(n16078), .B1(n26376), .B2(
        data_in[4]), .ZN(n16082) );
  INV_X1 U11677 ( .A(n16083), .ZN(n20069) );
  AOI22_X1 U11678 ( .A1(\mem[754][5] ), .A2(n16078), .B1(n26376), .B2(
        data_in[5]), .ZN(n16083) );
  INV_X1 U11679 ( .A(n16084), .ZN(n20068) );
  AOI22_X1 U11680 ( .A1(\mem[754][6] ), .A2(n16078), .B1(n26376), .B2(
        data_in[6]), .ZN(n16084) );
  INV_X1 U11681 ( .A(n16085), .ZN(n20067) );
  AOI22_X1 U11682 ( .A1(\mem[754][7] ), .A2(n16078), .B1(n26376), .B2(
        data_in[7]), .ZN(n16085) );
  INV_X1 U11683 ( .A(n16086), .ZN(n20066) );
  AOI22_X1 U11684 ( .A1(\mem[755][0] ), .A2(n16087), .B1(n26375), .B2(
        data_in[0]), .ZN(n16086) );
  INV_X1 U11685 ( .A(n16088), .ZN(n20065) );
  AOI22_X1 U11686 ( .A1(\mem[755][1] ), .A2(n16087), .B1(n26375), .B2(
        data_in[1]), .ZN(n16088) );
  INV_X1 U11687 ( .A(n16089), .ZN(n20064) );
  AOI22_X1 U11688 ( .A1(\mem[755][2] ), .A2(n16087), .B1(n26375), .B2(
        data_in[2]), .ZN(n16089) );
  INV_X1 U11689 ( .A(n16090), .ZN(n20063) );
  AOI22_X1 U11690 ( .A1(\mem[755][3] ), .A2(n16087), .B1(n26375), .B2(
        data_in[3]), .ZN(n16090) );
  INV_X1 U11691 ( .A(n16091), .ZN(n20062) );
  AOI22_X1 U11692 ( .A1(\mem[755][4] ), .A2(n16087), .B1(n26375), .B2(
        data_in[4]), .ZN(n16091) );
  INV_X1 U11693 ( .A(n16092), .ZN(n20061) );
  AOI22_X1 U11694 ( .A1(\mem[755][5] ), .A2(n16087), .B1(n26375), .B2(
        data_in[5]), .ZN(n16092) );
  INV_X1 U11695 ( .A(n16093), .ZN(n20060) );
  AOI22_X1 U11696 ( .A1(\mem[755][6] ), .A2(n16087), .B1(n26375), .B2(
        data_in[6]), .ZN(n16093) );
  INV_X1 U11697 ( .A(n16094), .ZN(n20059) );
  AOI22_X1 U11698 ( .A1(\mem[755][7] ), .A2(n16087), .B1(n26375), .B2(
        data_in[7]), .ZN(n16094) );
  INV_X1 U11699 ( .A(n16095), .ZN(n20058) );
  AOI22_X1 U11700 ( .A1(\mem[756][0] ), .A2(n16096), .B1(n26374), .B2(
        data_in[0]), .ZN(n16095) );
  INV_X1 U11701 ( .A(n16097), .ZN(n20057) );
  AOI22_X1 U11702 ( .A1(\mem[756][1] ), .A2(n16096), .B1(n26374), .B2(
        data_in[1]), .ZN(n16097) );
  INV_X1 U11703 ( .A(n16098), .ZN(n20056) );
  AOI22_X1 U11704 ( .A1(\mem[756][2] ), .A2(n16096), .B1(n26374), .B2(
        data_in[2]), .ZN(n16098) );
  INV_X1 U11705 ( .A(n16099), .ZN(n20055) );
  AOI22_X1 U11706 ( .A1(\mem[756][3] ), .A2(n16096), .B1(n26374), .B2(
        data_in[3]), .ZN(n16099) );
  INV_X1 U11707 ( .A(n16100), .ZN(n20054) );
  AOI22_X1 U11708 ( .A1(\mem[756][4] ), .A2(n16096), .B1(n26374), .B2(
        data_in[4]), .ZN(n16100) );
  INV_X1 U11709 ( .A(n16101), .ZN(n20053) );
  AOI22_X1 U11710 ( .A1(\mem[756][5] ), .A2(n16096), .B1(n26374), .B2(
        data_in[5]), .ZN(n16101) );
  INV_X1 U11711 ( .A(n16102), .ZN(n20052) );
  AOI22_X1 U11712 ( .A1(\mem[756][6] ), .A2(n16096), .B1(n26374), .B2(
        data_in[6]), .ZN(n16102) );
  INV_X1 U11713 ( .A(n16103), .ZN(n20051) );
  AOI22_X1 U11714 ( .A1(\mem[756][7] ), .A2(n16096), .B1(n26374), .B2(
        data_in[7]), .ZN(n16103) );
  INV_X1 U11715 ( .A(n16104), .ZN(n20050) );
  AOI22_X1 U11716 ( .A1(\mem[757][0] ), .A2(n16105), .B1(n26373), .B2(
        data_in[0]), .ZN(n16104) );
  INV_X1 U11717 ( .A(n16106), .ZN(n20049) );
  AOI22_X1 U11718 ( .A1(\mem[757][1] ), .A2(n16105), .B1(n26373), .B2(
        data_in[1]), .ZN(n16106) );
  INV_X1 U11719 ( .A(n16107), .ZN(n20048) );
  AOI22_X1 U11720 ( .A1(\mem[757][2] ), .A2(n16105), .B1(n26373), .B2(
        data_in[2]), .ZN(n16107) );
  INV_X1 U11721 ( .A(n16108), .ZN(n20047) );
  AOI22_X1 U11722 ( .A1(\mem[757][3] ), .A2(n16105), .B1(n26373), .B2(
        data_in[3]), .ZN(n16108) );
  INV_X1 U11723 ( .A(n16109), .ZN(n20046) );
  AOI22_X1 U11724 ( .A1(\mem[757][4] ), .A2(n16105), .B1(n26373), .B2(
        data_in[4]), .ZN(n16109) );
  INV_X1 U11725 ( .A(n16110), .ZN(n20045) );
  AOI22_X1 U11726 ( .A1(\mem[757][5] ), .A2(n16105), .B1(n26373), .B2(
        data_in[5]), .ZN(n16110) );
  INV_X1 U11727 ( .A(n16111), .ZN(n20044) );
  AOI22_X1 U11728 ( .A1(\mem[757][6] ), .A2(n16105), .B1(n26373), .B2(
        data_in[6]), .ZN(n16111) );
  INV_X1 U11729 ( .A(n16112), .ZN(n20043) );
  AOI22_X1 U11730 ( .A1(\mem[757][7] ), .A2(n16105), .B1(n26373), .B2(
        data_in[7]), .ZN(n16112) );
  INV_X1 U11731 ( .A(n16113), .ZN(n20042) );
  AOI22_X1 U11732 ( .A1(\mem[758][0] ), .A2(n16114), .B1(n26372), .B2(
        data_in[0]), .ZN(n16113) );
  INV_X1 U11733 ( .A(n16115), .ZN(n20041) );
  AOI22_X1 U11734 ( .A1(\mem[758][1] ), .A2(n16114), .B1(n26372), .B2(
        data_in[1]), .ZN(n16115) );
  INV_X1 U11735 ( .A(n16116), .ZN(n20040) );
  AOI22_X1 U11736 ( .A1(\mem[758][2] ), .A2(n16114), .B1(n26372), .B2(
        data_in[2]), .ZN(n16116) );
  INV_X1 U11737 ( .A(n16117), .ZN(n20039) );
  AOI22_X1 U11738 ( .A1(\mem[758][3] ), .A2(n16114), .B1(n26372), .B2(
        data_in[3]), .ZN(n16117) );
  INV_X1 U11739 ( .A(n16118), .ZN(n20038) );
  AOI22_X1 U11740 ( .A1(\mem[758][4] ), .A2(n16114), .B1(n26372), .B2(
        data_in[4]), .ZN(n16118) );
  INV_X1 U11741 ( .A(n16119), .ZN(n20037) );
  AOI22_X1 U11742 ( .A1(\mem[758][5] ), .A2(n16114), .B1(n26372), .B2(
        data_in[5]), .ZN(n16119) );
  INV_X1 U11743 ( .A(n16120), .ZN(n20036) );
  AOI22_X1 U11744 ( .A1(\mem[758][6] ), .A2(n16114), .B1(n26372), .B2(
        data_in[6]), .ZN(n16120) );
  INV_X1 U11745 ( .A(n16121), .ZN(n20035) );
  AOI22_X1 U11746 ( .A1(\mem[758][7] ), .A2(n16114), .B1(n26372), .B2(
        data_in[7]), .ZN(n16121) );
  INV_X1 U11747 ( .A(n16122), .ZN(n20034) );
  AOI22_X1 U11748 ( .A1(\mem[759][0] ), .A2(n16123), .B1(n26371), .B2(
        data_in[0]), .ZN(n16122) );
  INV_X1 U11749 ( .A(n16124), .ZN(n20033) );
  AOI22_X1 U11750 ( .A1(\mem[759][1] ), .A2(n16123), .B1(n26371), .B2(
        data_in[1]), .ZN(n16124) );
  INV_X1 U11751 ( .A(n16125), .ZN(n20032) );
  AOI22_X1 U11752 ( .A1(\mem[759][2] ), .A2(n16123), .B1(n26371), .B2(
        data_in[2]), .ZN(n16125) );
  INV_X1 U11753 ( .A(n16126), .ZN(n20031) );
  AOI22_X1 U11754 ( .A1(\mem[759][3] ), .A2(n16123), .B1(n26371), .B2(
        data_in[3]), .ZN(n16126) );
  INV_X1 U11755 ( .A(n16127), .ZN(n20030) );
  AOI22_X1 U11756 ( .A1(\mem[759][4] ), .A2(n16123), .B1(n26371), .B2(
        data_in[4]), .ZN(n16127) );
  INV_X1 U11757 ( .A(n16128), .ZN(n20029) );
  AOI22_X1 U11758 ( .A1(\mem[759][5] ), .A2(n16123), .B1(n26371), .B2(
        data_in[5]), .ZN(n16128) );
  INV_X1 U11759 ( .A(n16129), .ZN(n20028) );
  AOI22_X1 U11760 ( .A1(\mem[759][6] ), .A2(n16123), .B1(n26371), .B2(
        data_in[6]), .ZN(n16129) );
  INV_X1 U11761 ( .A(n16130), .ZN(n20027) );
  AOI22_X1 U11762 ( .A1(\mem[759][7] ), .A2(n16123), .B1(n26371), .B2(
        data_in[7]), .ZN(n16130) );
  INV_X1 U11763 ( .A(n16131), .ZN(n20026) );
  AOI22_X1 U11764 ( .A1(\mem[760][0] ), .A2(n16132), .B1(n26370), .B2(
        data_in[0]), .ZN(n16131) );
  INV_X1 U11765 ( .A(n16133), .ZN(n20025) );
  AOI22_X1 U11766 ( .A1(\mem[760][1] ), .A2(n16132), .B1(n26370), .B2(
        data_in[1]), .ZN(n16133) );
  INV_X1 U11767 ( .A(n16134), .ZN(n20024) );
  AOI22_X1 U11768 ( .A1(\mem[760][2] ), .A2(n16132), .B1(n26370), .B2(
        data_in[2]), .ZN(n16134) );
  INV_X1 U11769 ( .A(n16135), .ZN(n20023) );
  AOI22_X1 U11770 ( .A1(\mem[760][3] ), .A2(n16132), .B1(n26370), .B2(
        data_in[3]), .ZN(n16135) );
  INV_X1 U11771 ( .A(n16136), .ZN(n20022) );
  AOI22_X1 U11772 ( .A1(\mem[760][4] ), .A2(n16132), .B1(n26370), .B2(
        data_in[4]), .ZN(n16136) );
  INV_X1 U11773 ( .A(n16137), .ZN(n20021) );
  AOI22_X1 U11774 ( .A1(\mem[760][5] ), .A2(n16132), .B1(n26370), .B2(
        data_in[5]), .ZN(n16137) );
  INV_X1 U11775 ( .A(n16138), .ZN(n20020) );
  AOI22_X1 U11776 ( .A1(\mem[760][6] ), .A2(n16132), .B1(n26370), .B2(
        data_in[6]), .ZN(n16138) );
  INV_X1 U11777 ( .A(n16139), .ZN(n20019) );
  AOI22_X1 U11778 ( .A1(\mem[760][7] ), .A2(n16132), .B1(n26370), .B2(
        data_in[7]), .ZN(n16139) );
  INV_X1 U11779 ( .A(n16140), .ZN(n20018) );
  AOI22_X1 U11780 ( .A1(\mem[761][0] ), .A2(n16141), .B1(n26369), .B2(
        data_in[0]), .ZN(n16140) );
  INV_X1 U11781 ( .A(n16142), .ZN(n20017) );
  AOI22_X1 U11782 ( .A1(\mem[761][1] ), .A2(n16141), .B1(n26369), .B2(
        data_in[1]), .ZN(n16142) );
  INV_X1 U11783 ( .A(n16143), .ZN(n20016) );
  AOI22_X1 U11784 ( .A1(\mem[761][2] ), .A2(n16141), .B1(n26369), .B2(
        data_in[2]), .ZN(n16143) );
  INV_X1 U11785 ( .A(n16144), .ZN(n20015) );
  AOI22_X1 U11786 ( .A1(\mem[761][3] ), .A2(n16141), .B1(n26369), .B2(
        data_in[3]), .ZN(n16144) );
  INV_X1 U11787 ( .A(n16145), .ZN(n20014) );
  AOI22_X1 U11788 ( .A1(\mem[761][4] ), .A2(n16141), .B1(n26369), .B2(
        data_in[4]), .ZN(n16145) );
  INV_X1 U11789 ( .A(n16146), .ZN(n20013) );
  AOI22_X1 U11790 ( .A1(\mem[761][5] ), .A2(n16141), .B1(n26369), .B2(
        data_in[5]), .ZN(n16146) );
  INV_X1 U11791 ( .A(n16147), .ZN(n20012) );
  AOI22_X1 U11792 ( .A1(\mem[761][6] ), .A2(n16141), .B1(n26369), .B2(
        data_in[6]), .ZN(n16147) );
  INV_X1 U11793 ( .A(n16148), .ZN(n20011) );
  AOI22_X1 U11794 ( .A1(\mem[761][7] ), .A2(n16141), .B1(n26369), .B2(
        data_in[7]), .ZN(n16148) );
  INV_X1 U11795 ( .A(n16149), .ZN(n20010) );
  AOI22_X1 U11796 ( .A1(\mem[762][0] ), .A2(n16150), .B1(n26368), .B2(
        data_in[0]), .ZN(n16149) );
  INV_X1 U11797 ( .A(n16151), .ZN(n20009) );
  AOI22_X1 U11798 ( .A1(\mem[762][1] ), .A2(n16150), .B1(n26368), .B2(
        data_in[1]), .ZN(n16151) );
  INV_X1 U11799 ( .A(n16152), .ZN(n20008) );
  AOI22_X1 U11800 ( .A1(\mem[762][2] ), .A2(n16150), .B1(n26368), .B2(
        data_in[2]), .ZN(n16152) );
  INV_X1 U11801 ( .A(n16153), .ZN(n20007) );
  AOI22_X1 U11802 ( .A1(\mem[762][3] ), .A2(n16150), .B1(n26368), .B2(
        data_in[3]), .ZN(n16153) );
  INV_X1 U11803 ( .A(n16154), .ZN(n20006) );
  AOI22_X1 U11804 ( .A1(\mem[762][4] ), .A2(n16150), .B1(n26368), .B2(
        data_in[4]), .ZN(n16154) );
  INV_X1 U11805 ( .A(n16155), .ZN(n20005) );
  AOI22_X1 U11806 ( .A1(\mem[762][5] ), .A2(n16150), .B1(n26368), .B2(
        data_in[5]), .ZN(n16155) );
  INV_X1 U11807 ( .A(n16156), .ZN(n20004) );
  AOI22_X1 U11808 ( .A1(\mem[762][6] ), .A2(n16150), .B1(n26368), .B2(
        data_in[6]), .ZN(n16156) );
  INV_X1 U11809 ( .A(n16157), .ZN(n20003) );
  AOI22_X1 U11810 ( .A1(\mem[762][7] ), .A2(n16150), .B1(n26368), .B2(
        data_in[7]), .ZN(n16157) );
  INV_X1 U11811 ( .A(n16158), .ZN(n20002) );
  AOI22_X1 U11812 ( .A1(\mem[763][0] ), .A2(n16159), .B1(n26367), .B2(
        data_in[0]), .ZN(n16158) );
  INV_X1 U11813 ( .A(n16160), .ZN(n20001) );
  AOI22_X1 U11814 ( .A1(\mem[763][1] ), .A2(n16159), .B1(n26367), .B2(
        data_in[1]), .ZN(n16160) );
  INV_X1 U11815 ( .A(n16161), .ZN(n20000) );
  AOI22_X1 U11816 ( .A1(\mem[763][2] ), .A2(n16159), .B1(n26367), .B2(
        data_in[2]), .ZN(n16161) );
  INV_X1 U11817 ( .A(n16162), .ZN(n19999) );
  AOI22_X1 U11818 ( .A1(\mem[763][3] ), .A2(n16159), .B1(n26367), .B2(
        data_in[3]), .ZN(n16162) );
  INV_X1 U11819 ( .A(n16163), .ZN(n19998) );
  AOI22_X1 U11820 ( .A1(\mem[763][4] ), .A2(n16159), .B1(n26367), .B2(
        data_in[4]), .ZN(n16163) );
  INV_X1 U11821 ( .A(n16164), .ZN(n19997) );
  AOI22_X1 U11822 ( .A1(\mem[763][5] ), .A2(n16159), .B1(n26367), .B2(
        data_in[5]), .ZN(n16164) );
  INV_X1 U11823 ( .A(n16165), .ZN(n19996) );
  AOI22_X1 U11824 ( .A1(\mem[763][6] ), .A2(n16159), .B1(n26367), .B2(
        data_in[6]), .ZN(n16165) );
  INV_X1 U11825 ( .A(n16166), .ZN(n19995) );
  AOI22_X1 U11826 ( .A1(\mem[763][7] ), .A2(n16159), .B1(n26367), .B2(
        data_in[7]), .ZN(n16166) );
  INV_X1 U11827 ( .A(n16167), .ZN(n19994) );
  AOI22_X1 U11828 ( .A1(\mem[764][0] ), .A2(n16168), .B1(n26366), .B2(
        data_in[0]), .ZN(n16167) );
  INV_X1 U11829 ( .A(n16169), .ZN(n19993) );
  AOI22_X1 U11830 ( .A1(\mem[764][1] ), .A2(n16168), .B1(n26366), .B2(
        data_in[1]), .ZN(n16169) );
  INV_X1 U11831 ( .A(n16170), .ZN(n19992) );
  AOI22_X1 U11832 ( .A1(\mem[764][2] ), .A2(n16168), .B1(n26366), .B2(
        data_in[2]), .ZN(n16170) );
  INV_X1 U11833 ( .A(n16171), .ZN(n19991) );
  AOI22_X1 U11834 ( .A1(\mem[764][3] ), .A2(n16168), .B1(n26366), .B2(
        data_in[3]), .ZN(n16171) );
  INV_X1 U11835 ( .A(n16172), .ZN(n19990) );
  AOI22_X1 U11836 ( .A1(\mem[764][4] ), .A2(n16168), .B1(n26366), .B2(
        data_in[4]), .ZN(n16172) );
  INV_X1 U11837 ( .A(n16173), .ZN(n19989) );
  AOI22_X1 U11838 ( .A1(\mem[764][5] ), .A2(n16168), .B1(n26366), .B2(
        data_in[5]), .ZN(n16173) );
  INV_X1 U11839 ( .A(n16174), .ZN(n19988) );
  AOI22_X1 U11840 ( .A1(\mem[764][6] ), .A2(n16168), .B1(n26366), .B2(
        data_in[6]), .ZN(n16174) );
  INV_X1 U11841 ( .A(n16175), .ZN(n19987) );
  AOI22_X1 U11842 ( .A1(\mem[764][7] ), .A2(n16168), .B1(n26366), .B2(
        data_in[7]), .ZN(n16175) );
  INV_X1 U11843 ( .A(n16176), .ZN(n19986) );
  AOI22_X1 U11844 ( .A1(\mem[765][0] ), .A2(n16177), .B1(n26365), .B2(
        data_in[0]), .ZN(n16176) );
  INV_X1 U11845 ( .A(n16178), .ZN(n19985) );
  AOI22_X1 U11846 ( .A1(\mem[765][1] ), .A2(n16177), .B1(n26365), .B2(
        data_in[1]), .ZN(n16178) );
  INV_X1 U11847 ( .A(n16179), .ZN(n19984) );
  AOI22_X1 U11848 ( .A1(\mem[765][2] ), .A2(n16177), .B1(n26365), .B2(
        data_in[2]), .ZN(n16179) );
  INV_X1 U11849 ( .A(n16180), .ZN(n19983) );
  AOI22_X1 U11850 ( .A1(\mem[765][3] ), .A2(n16177), .B1(n26365), .B2(
        data_in[3]), .ZN(n16180) );
  INV_X1 U11851 ( .A(n16181), .ZN(n19982) );
  AOI22_X1 U11852 ( .A1(\mem[765][4] ), .A2(n16177), .B1(n26365), .B2(
        data_in[4]), .ZN(n16181) );
  INV_X1 U11853 ( .A(n16182), .ZN(n19981) );
  AOI22_X1 U11854 ( .A1(\mem[765][5] ), .A2(n16177), .B1(n26365), .B2(
        data_in[5]), .ZN(n16182) );
  INV_X1 U11855 ( .A(n16183), .ZN(n19980) );
  AOI22_X1 U11856 ( .A1(\mem[765][6] ), .A2(n16177), .B1(n26365), .B2(
        data_in[6]), .ZN(n16183) );
  INV_X1 U11857 ( .A(n16184), .ZN(n19979) );
  AOI22_X1 U11858 ( .A1(\mem[765][7] ), .A2(n16177), .B1(n26365), .B2(
        data_in[7]), .ZN(n16184) );
  INV_X1 U11859 ( .A(n16185), .ZN(n19978) );
  AOI22_X1 U11860 ( .A1(\mem[766][0] ), .A2(n16186), .B1(n26364), .B2(
        data_in[0]), .ZN(n16185) );
  INV_X1 U11861 ( .A(n16187), .ZN(n19977) );
  AOI22_X1 U11862 ( .A1(\mem[766][1] ), .A2(n16186), .B1(n26364), .B2(
        data_in[1]), .ZN(n16187) );
  INV_X1 U11863 ( .A(n16188), .ZN(n19976) );
  AOI22_X1 U11864 ( .A1(\mem[766][2] ), .A2(n16186), .B1(n26364), .B2(
        data_in[2]), .ZN(n16188) );
  INV_X1 U11865 ( .A(n16189), .ZN(n19975) );
  AOI22_X1 U11866 ( .A1(\mem[766][3] ), .A2(n16186), .B1(n26364), .B2(
        data_in[3]), .ZN(n16189) );
  INV_X1 U11867 ( .A(n16190), .ZN(n19974) );
  AOI22_X1 U11868 ( .A1(\mem[766][4] ), .A2(n16186), .B1(n26364), .B2(
        data_in[4]), .ZN(n16190) );
  INV_X1 U11869 ( .A(n16191), .ZN(n19973) );
  AOI22_X1 U11870 ( .A1(\mem[766][5] ), .A2(n16186), .B1(n26364), .B2(
        data_in[5]), .ZN(n16191) );
  INV_X1 U11871 ( .A(n16192), .ZN(n19972) );
  AOI22_X1 U11872 ( .A1(\mem[766][6] ), .A2(n16186), .B1(n26364), .B2(
        data_in[6]), .ZN(n16192) );
  INV_X1 U11873 ( .A(n16193), .ZN(n19971) );
  AOI22_X1 U11874 ( .A1(\mem[766][7] ), .A2(n16186), .B1(n26364), .B2(
        data_in[7]), .ZN(n16193) );
  INV_X1 U11875 ( .A(n16194), .ZN(n19970) );
  AOI22_X1 U11876 ( .A1(\mem[767][0] ), .A2(n16195), .B1(n26363), .B2(
        data_in[0]), .ZN(n16194) );
  INV_X1 U11877 ( .A(n16196), .ZN(n19969) );
  AOI22_X1 U11878 ( .A1(\mem[767][1] ), .A2(n16195), .B1(n26363), .B2(
        data_in[1]), .ZN(n16196) );
  INV_X1 U11879 ( .A(n16197), .ZN(n19968) );
  AOI22_X1 U11880 ( .A1(\mem[767][2] ), .A2(n16195), .B1(n26363), .B2(
        data_in[2]), .ZN(n16197) );
  INV_X1 U11881 ( .A(n16198), .ZN(n19967) );
  AOI22_X1 U11882 ( .A1(\mem[767][3] ), .A2(n16195), .B1(n26363), .B2(
        data_in[3]), .ZN(n16198) );
  INV_X1 U11883 ( .A(n16199), .ZN(n19966) );
  AOI22_X1 U11884 ( .A1(\mem[767][4] ), .A2(n16195), .B1(n26363), .B2(
        data_in[4]), .ZN(n16199) );
  INV_X1 U11885 ( .A(n16200), .ZN(n19965) );
  AOI22_X1 U11886 ( .A1(\mem[767][5] ), .A2(n16195), .B1(n26363), .B2(
        data_in[5]), .ZN(n16200) );
  INV_X1 U11887 ( .A(n16201), .ZN(n19964) );
  AOI22_X1 U11888 ( .A1(\mem[767][6] ), .A2(n16195), .B1(n26363), .B2(
        data_in[6]), .ZN(n16201) );
  INV_X1 U11889 ( .A(n16202), .ZN(n19963) );
  AOI22_X1 U11890 ( .A1(\mem[767][7] ), .A2(n16195), .B1(n26363), .B2(
        data_in[7]), .ZN(n16202) );
  INV_X1 U11891 ( .A(n16276), .ZN(n19898) );
  AOI22_X1 U11892 ( .A1(\mem[776][0] ), .A2(n16277), .B1(n26354), .B2(
        data_in[0]), .ZN(n16276) );
  INV_X1 U11893 ( .A(n16278), .ZN(n19897) );
  AOI22_X1 U11894 ( .A1(\mem[776][1] ), .A2(n16277), .B1(n26354), .B2(
        data_in[1]), .ZN(n16278) );
  INV_X1 U11895 ( .A(n16279), .ZN(n19896) );
  AOI22_X1 U11896 ( .A1(\mem[776][2] ), .A2(n16277), .B1(n26354), .B2(
        data_in[2]), .ZN(n16279) );
  INV_X1 U11897 ( .A(n16280), .ZN(n19895) );
  AOI22_X1 U11898 ( .A1(\mem[776][3] ), .A2(n16277), .B1(n26354), .B2(
        data_in[3]), .ZN(n16280) );
  INV_X1 U11899 ( .A(n16281), .ZN(n19894) );
  AOI22_X1 U11900 ( .A1(\mem[776][4] ), .A2(n16277), .B1(n26354), .B2(
        data_in[4]), .ZN(n16281) );
  INV_X1 U11901 ( .A(n16282), .ZN(n19893) );
  AOI22_X1 U11902 ( .A1(\mem[776][5] ), .A2(n16277), .B1(n26354), .B2(
        data_in[5]), .ZN(n16282) );
  INV_X1 U11903 ( .A(n16283), .ZN(n19892) );
  AOI22_X1 U11904 ( .A1(\mem[776][6] ), .A2(n16277), .B1(n26354), .B2(
        data_in[6]), .ZN(n16283) );
  INV_X1 U11905 ( .A(n16284), .ZN(n19891) );
  AOI22_X1 U11906 ( .A1(\mem[776][7] ), .A2(n16277), .B1(n26354), .B2(
        data_in[7]), .ZN(n16284) );
  INV_X1 U11907 ( .A(n16285), .ZN(n19890) );
  AOI22_X1 U11908 ( .A1(\mem[777][0] ), .A2(n16286), .B1(n26353), .B2(
        data_in[0]), .ZN(n16285) );
  INV_X1 U11909 ( .A(n16287), .ZN(n19889) );
  AOI22_X1 U11910 ( .A1(\mem[777][1] ), .A2(n16286), .B1(n26353), .B2(
        data_in[1]), .ZN(n16287) );
  INV_X1 U11911 ( .A(n16288), .ZN(n19888) );
  AOI22_X1 U11912 ( .A1(\mem[777][2] ), .A2(n16286), .B1(n26353), .B2(
        data_in[2]), .ZN(n16288) );
  INV_X1 U11913 ( .A(n16289), .ZN(n19887) );
  AOI22_X1 U11914 ( .A1(\mem[777][3] ), .A2(n16286), .B1(n26353), .B2(
        data_in[3]), .ZN(n16289) );
  INV_X1 U11915 ( .A(n16290), .ZN(n19886) );
  AOI22_X1 U11916 ( .A1(\mem[777][4] ), .A2(n16286), .B1(n26353), .B2(
        data_in[4]), .ZN(n16290) );
  INV_X1 U11917 ( .A(n16291), .ZN(n19885) );
  AOI22_X1 U11918 ( .A1(\mem[777][5] ), .A2(n16286), .B1(n26353), .B2(
        data_in[5]), .ZN(n16291) );
  INV_X1 U11919 ( .A(n16292), .ZN(n19884) );
  AOI22_X1 U11920 ( .A1(\mem[777][6] ), .A2(n16286), .B1(n26353), .B2(
        data_in[6]), .ZN(n16292) );
  INV_X1 U11921 ( .A(n16293), .ZN(n19883) );
  AOI22_X1 U11922 ( .A1(\mem[777][7] ), .A2(n16286), .B1(n26353), .B2(
        data_in[7]), .ZN(n16293) );
  INV_X1 U11923 ( .A(n16294), .ZN(n19882) );
  AOI22_X1 U11924 ( .A1(\mem[778][0] ), .A2(n16295), .B1(n26352), .B2(
        data_in[0]), .ZN(n16294) );
  INV_X1 U11925 ( .A(n16296), .ZN(n19881) );
  AOI22_X1 U11926 ( .A1(\mem[778][1] ), .A2(n16295), .B1(n26352), .B2(
        data_in[1]), .ZN(n16296) );
  INV_X1 U11927 ( .A(n16297), .ZN(n19880) );
  AOI22_X1 U11928 ( .A1(\mem[778][2] ), .A2(n16295), .B1(n26352), .B2(
        data_in[2]), .ZN(n16297) );
  INV_X1 U11929 ( .A(n16298), .ZN(n19879) );
  AOI22_X1 U11930 ( .A1(\mem[778][3] ), .A2(n16295), .B1(n26352), .B2(
        data_in[3]), .ZN(n16298) );
  INV_X1 U11931 ( .A(n16299), .ZN(n19878) );
  AOI22_X1 U11932 ( .A1(\mem[778][4] ), .A2(n16295), .B1(n26352), .B2(
        data_in[4]), .ZN(n16299) );
  INV_X1 U11933 ( .A(n16300), .ZN(n19877) );
  AOI22_X1 U11934 ( .A1(\mem[778][5] ), .A2(n16295), .B1(n26352), .B2(
        data_in[5]), .ZN(n16300) );
  INV_X1 U11935 ( .A(n16301), .ZN(n19876) );
  AOI22_X1 U11936 ( .A1(\mem[778][6] ), .A2(n16295), .B1(n26352), .B2(
        data_in[6]), .ZN(n16301) );
  INV_X1 U11937 ( .A(n16302), .ZN(n19875) );
  AOI22_X1 U11938 ( .A1(\mem[778][7] ), .A2(n16295), .B1(n26352), .B2(
        data_in[7]), .ZN(n16302) );
  INV_X1 U11939 ( .A(n16303), .ZN(n19874) );
  AOI22_X1 U11940 ( .A1(\mem[779][0] ), .A2(n16304), .B1(n26351), .B2(
        data_in[0]), .ZN(n16303) );
  INV_X1 U11941 ( .A(n16305), .ZN(n19873) );
  AOI22_X1 U11942 ( .A1(\mem[779][1] ), .A2(n16304), .B1(n26351), .B2(
        data_in[1]), .ZN(n16305) );
  INV_X1 U11943 ( .A(n16306), .ZN(n19872) );
  AOI22_X1 U11944 ( .A1(\mem[779][2] ), .A2(n16304), .B1(n26351), .B2(
        data_in[2]), .ZN(n16306) );
  INV_X1 U11945 ( .A(n16307), .ZN(n19871) );
  AOI22_X1 U11946 ( .A1(\mem[779][3] ), .A2(n16304), .B1(n26351), .B2(
        data_in[3]), .ZN(n16307) );
  INV_X1 U11947 ( .A(n16308), .ZN(n19870) );
  AOI22_X1 U11948 ( .A1(\mem[779][4] ), .A2(n16304), .B1(n26351), .B2(
        data_in[4]), .ZN(n16308) );
  INV_X1 U11949 ( .A(n16309), .ZN(n19869) );
  AOI22_X1 U11950 ( .A1(\mem[779][5] ), .A2(n16304), .B1(n26351), .B2(
        data_in[5]), .ZN(n16309) );
  INV_X1 U11951 ( .A(n16310), .ZN(n19868) );
  AOI22_X1 U11952 ( .A1(\mem[779][6] ), .A2(n16304), .B1(n26351), .B2(
        data_in[6]), .ZN(n16310) );
  INV_X1 U11953 ( .A(n16311), .ZN(n19867) );
  AOI22_X1 U11954 ( .A1(\mem[779][7] ), .A2(n16304), .B1(n26351), .B2(
        data_in[7]), .ZN(n16311) );
  INV_X1 U11955 ( .A(n16312), .ZN(n19866) );
  AOI22_X1 U11956 ( .A1(\mem[780][0] ), .A2(n16313), .B1(n26350), .B2(
        data_in[0]), .ZN(n16312) );
  INV_X1 U11957 ( .A(n16314), .ZN(n19865) );
  AOI22_X1 U11958 ( .A1(\mem[780][1] ), .A2(n16313), .B1(n26350), .B2(
        data_in[1]), .ZN(n16314) );
  INV_X1 U11959 ( .A(n16315), .ZN(n19864) );
  AOI22_X1 U11960 ( .A1(\mem[780][2] ), .A2(n16313), .B1(n26350), .B2(
        data_in[2]), .ZN(n16315) );
  INV_X1 U11961 ( .A(n16316), .ZN(n19863) );
  AOI22_X1 U11962 ( .A1(\mem[780][3] ), .A2(n16313), .B1(n26350), .B2(
        data_in[3]), .ZN(n16316) );
  INV_X1 U11963 ( .A(n16317), .ZN(n19862) );
  AOI22_X1 U11964 ( .A1(\mem[780][4] ), .A2(n16313), .B1(n26350), .B2(
        data_in[4]), .ZN(n16317) );
  INV_X1 U11965 ( .A(n16318), .ZN(n19861) );
  AOI22_X1 U11966 ( .A1(\mem[780][5] ), .A2(n16313), .B1(n26350), .B2(
        data_in[5]), .ZN(n16318) );
  INV_X1 U11967 ( .A(n16319), .ZN(n19860) );
  AOI22_X1 U11968 ( .A1(\mem[780][6] ), .A2(n16313), .B1(n26350), .B2(
        data_in[6]), .ZN(n16319) );
  INV_X1 U11969 ( .A(n16320), .ZN(n19859) );
  AOI22_X1 U11970 ( .A1(\mem[780][7] ), .A2(n16313), .B1(n26350), .B2(
        data_in[7]), .ZN(n16320) );
  INV_X1 U11971 ( .A(n16321), .ZN(n19858) );
  AOI22_X1 U11972 ( .A1(\mem[781][0] ), .A2(n16322), .B1(n26349), .B2(
        data_in[0]), .ZN(n16321) );
  INV_X1 U11973 ( .A(n16323), .ZN(n19857) );
  AOI22_X1 U11974 ( .A1(\mem[781][1] ), .A2(n16322), .B1(n26349), .B2(
        data_in[1]), .ZN(n16323) );
  INV_X1 U11975 ( .A(n16324), .ZN(n19856) );
  AOI22_X1 U11976 ( .A1(\mem[781][2] ), .A2(n16322), .B1(n26349), .B2(
        data_in[2]), .ZN(n16324) );
  INV_X1 U11977 ( .A(n16325), .ZN(n19855) );
  AOI22_X1 U11978 ( .A1(\mem[781][3] ), .A2(n16322), .B1(n26349), .B2(
        data_in[3]), .ZN(n16325) );
  INV_X1 U11979 ( .A(n16326), .ZN(n19854) );
  AOI22_X1 U11980 ( .A1(\mem[781][4] ), .A2(n16322), .B1(n26349), .B2(
        data_in[4]), .ZN(n16326) );
  INV_X1 U11981 ( .A(n16327), .ZN(n19853) );
  AOI22_X1 U11982 ( .A1(\mem[781][5] ), .A2(n16322), .B1(n26349), .B2(
        data_in[5]), .ZN(n16327) );
  INV_X1 U11983 ( .A(n16328), .ZN(n19852) );
  AOI22_X1 U11984 ( .A1(\mem[781][6] ), .A2(n16322), .B1(n26349), .B2(
        data_in[6]), .ZN(n16328) );
  INV_X1 U11985 ( .A(n16329), .ZN(n19851) );
  AOI22_X1 U11986 ( .A1(\mem[781][7] ), .A2(n16322), .B1(n26349), .B2(
        data_in[7]), .ZN(n16329) );
  INV_X1 U11987 ( .A(n16330), .ZN(n19850) );
  AOI22_X1 U11988 ( .A1(\mem[782][0] ), .A2(n16331), .B1(n26348), .B2(
        data_in[0]), .ZN(n16330) );
  INV_X1 U11989 ( .A(n16332), .ZN(n19849) );
  AOI22_X1 U11990 ( .A1(\mem[782][1] ), .A2(n16331), .B1(n26348), .B2(
        data_in[1]), .ZN(n16332) );
  INV_X1 U11991 ( .A(n16333), .ZN(n19848) );
  AOI22_X1 U11992 ( .A1(\mem[782][2] ), .A2(n16331), .B1(n26348), .B2(
        data_in[2]), .ZN(n16333) );
  INV_X1 U11993 ( .A(n16334), .ZN(n19847) );
  AOI22_X1 U11994 ( .A1(\mem[782][3] ), .A2(n16331), .B1(n26348), .B2(
        data_in[3]), .ZN(n16334) );
  INV_X1 U11995 ( .A(n16335), .ZN(n19846) );
  AOI22_X1 U11996 ( .A1(\mem[782][4] ), .A2(n16331), .B1(n26348), .B2(
        data_in[4]), .ZN(n16335) );
  INV_X1 U11997 ( .A(n16336), .ZN(n19845) );
  AOI22_X1 U11998 ( .A1(\mem[782][5] ), .A2(n16331), .B1(n26348), .B2(
        data_in[5]), .ZN(n16336) );
  INV_X1 U11999 ( .A(n16337), .ZN(n19844) );
  AOI22_X1 U12000 ( .A1(\mem[782][6] ), .A2(n16331), .B1(n26348), .B2(
        data_in[6]), .ZN(n16337) );
  INV_X1 U12001 ( .A(n16338), .ZN(n19843) );
  AOI22_X1 U12002 ( .A1(\mem[782][7] ), .A2(n16331), .B1(n26348), .B2(
        data_in[7]), .ZN(n16338) );
  INV_X1 U12003 ( .A(n16339), .ZN(n19842) );
  AOI22_X1 U12004 ( .A1(\mem[783][0] ), .A2(n16340), .B1(n26347), .B2(
        data_in[0]), .ZN(n16339) );
  INV_X1 U12005 ( .A(n16341), .ZN(n19841) );
  AOI22_X1 U12006 ( .A1(\mem[783][1] ), .A2(n16340), .B1(n26347), .B2(
        data_in[1]), .ZN(n16341) );
  INV_X1 U12007 ( .A(n16342), .ZN(n19840) );
  AOI22_X1 U12008 ( .A1(\mem[783][2] ), .A2(n16340), .B1(n26347), .B2(
        data_in[2]), .ZN(n16342) );
  INV_X1 U12009 ( .A(n16343), .ZN(n19839) );
  AOI22_X1 U12010 ( .A1(\mem[783][3] ), .A2(n16340), .B1(n26347), .B2(
        data_in[3]), .ZN(n16343) );
  INV_X1 U12011 ( .A(n16344), .ZN(n19838) );
  AOI22_X1 U12012 ( .A1(\mem[783][4] ), .A2(n16340), .B1(n26347), .B2(
        data_in[4]), .ZN(n16344) );
  INV_X1 U12013 ( .A(n16345), .ZN(n19837) );
  AOI22_X1 U12014 ( .A1(\mem[783][5] ), .A2(n16340), .B1(n26347), .B2(
        data_in[5]), .ZN(n16345) );
  INV_X1 U12015 ( .A(n16346), .ZN(n19836) );
  AOI22_X1 U12016 ( .A1(\mem[783][6] ), .A2(n16340), .B1(n26347), .B2(
        data_in[6]), .ZN(n16346) );
  INV_X1 U12017 ( .A(n16347), .ZN(n19835) );
  AOI22_X1 U12018 ( .A1(\mem[783][7] ), .A2(n16340), .B1(n26347), .B2(
        data_in[7]), .ZN(n16347) );
  INV_X1 U12019 ( .A(n16348), .ZN(n19834) );
  AOI22_X1 U12020 ( .A1(\mem[784][0] ), .A2(n16349), .B1(n26346), .B2(
        data_in[0]), .ZN(n16348) );
  INV_X1 U12021 ( .A(n16350), .ZN(n19833) );
  AOI22_X1 U12022 ( .A1(\mem[784][1] ), .A2(n16349), .B1(n26346), .B2(
        data_in[1]), .ZN(n16350) );
  INV_X1 U12023 ( .A(n16351), .ZN(n19832) );
  AOI22_X1 U12024 ( .A1(\mem[784][2] ), .A2(n16349), .B1(n26346), .B2(
        data_in[2]), .ZN(n16351) );
  INV_X1 U12025 ( .A(n16352), .ZN(n19831) );
  AOI22_X1 U12026 ( .A1(\mem[784][3] ), .A2(n16349), .B1(n26346), .B2(
        data_in[3]), .ZN(n16352) );
  INV_X1 U12027 ( .A(n16353), .ZN(n19830) );
  AOI22_X1 U12028 ( .A1(\mem[784][4] ), .A2(n16349), .B1(n26346), .B2(
        data_in[4]), .ZN(n16353) );
  INV_X1 U12029 ( .A(n16354), .ZN(n19829) );
  AOI22_X1 U12030 ( .A1(\mem[784][5] ), .A2(n16349), .B1(n26346), .B2(
        data_in[5]), .ZN(n16354) );
  INV_X1 U12031 ( .A(n16355), .ZN(n19828) );
  AOI22_X1 U12032 ( .A1(\mem[784][6] ), .A2(n16349), .B1(n26346), .B2(
        data_in[6]), .ZN(n16355) );
  INV_X1 U12033 ( .A(n16356), .ZN(n19827) );
  AOI22_X1 U12034 ( .A1(\mem[784][7] ), .A2(n16349), .B1(n26346), .B2(
        data_in[7]), .ZN(n16356) );
  INV_X1 U12035 ( .A(n16357), .ZN(n19826) );
  AOI22_X1 U12036 ( .A1(\mem[785][0] ), .A2(n16358), .B1(n26345), .B2(
        data_in[0]), .ZN(n16357) );
  INV_X1 U12037 ( .A(n16359), .ZN(n19825) );
  AOI22_X1 U12038 ( .A1(\mem[785][1] ), .A2(n16358), .B1(n26345), .B2(
        data_in[1]), .ZN(n16359) );
  INV_X1 U12039 ( .A(n16360), .ZN(n19824) );
  AOI22_X1 U12040 ( .A1(\mem[785][2] ), .A2(n16358), .B1(n26345), .B2(
        data_in[2]), .ZN(n16360) );
  INV_X1 U12041 ( .A(n16361), .ZN(n19823) );
  AOI22_X1 U12042 ( .A1(\mem[785][3] ), .A2(n16358), .B1(n26345), .B2(
        data_in[3]), .ZN(n16361) );
  INV_X1 U12043 ( .A(n16362), .ZN(n19822) );
  AOI22_X1 U12044 ( .A1(\mem[785][4] ), .A2(n16358), .B1(n26345), .B2(
        data_in[4]), .ZN(n16362) );
  INV_X1 U12045 ( .A(n16363), .ZN(n19821) );
  AOI22_X1 U12046 ( .A1(\mem[785][5] ), .A2(n16358), .B1(n26345), .B2(
        data_in[5]), .ZN(n16363) );
  INV_X1 U12047 ( .A(n16364), .ZN(n19820) );
  AOI22_X1 U12048 ( .A1(\mem[785][6] ), .A2(n16358), .B1(n26345), .B2(
        data_in[6]), .ZN(n16364) );
  INV_X1 U12049 ( .A(n16365), .ZN(n19819) );
  AOI22_X1 U12050 ( .A1(\mem[785][7] ), .A2(n16358), .B1(n26345), .B2(
        data_in[7]), .ZN(n16365) );
  INV_X1 U12051 ( .A(n16366), .ZN(n19818) );
  AOI22_X1 U12052 ( .A1(\mem[786][0] ), .A2(n16367), .B1(n26344), .B2(
        data_in[0]), .ZN(n16366) );
  INV_X1 U12053 ( .A(n16368), .ZN(n19817) );
  AOI22_X1 U12054 ( .A1(\mem[786][1] ), .A2(n16367), .B1(n26344), .B2(
        data_in[1]), .ZN(n16368) );
  INV_X1 U12055 ( .A(n16369), .ZN(n19816) );
  AOI22_X1 U12056 ( .A1(\mem[786][2] ), .A2(n16367), .B1(n26344), .B2(
        data_in[2]), .ZN(n16369) );
  INV_X1 U12057 ( .A(n16370), .ZN(n19815) );
  AOI22_X1 U12058 ( .A1(\mem[786][3] ), .A2(n16367), .B1(n26344), .B2(
        data_in[3]), .ZN(n16370) );
  INV_X1 U12059 ( .A(n16371), .ZN(n19814) );
  AOI22_X1 U12060 ( .A1(\mem[786][4] ), .A2(n16367), .B1(n26344), .B2(
        data_in[4]), .ZN(n16371) );
  INV_X1 U12061 ( .A(n16372), .ZN(n19813) );
  AOI22_X1 U12062 ( .A1(\mem[786][5] ), .A2(n16367), .B1(n26344), .B2(
        data_in[5]), .ZN(n16372) );
  INV_X1 U12063 ( .A(n16373), .ZN(n19812) );
  AOI22_X1 U12064 ( .A1(\mem[786][6] ), .A2(n16367), .B1(n26344), .B2(
        data_in[6]), .ZN(n16373) );
  INV_X1 U12065 ( .A(n16374), .ZN(n19811) );
  AOI22_X1 U12066 ( .A1(\mem[786][7] ), .A2(n16367), .B1(n26344), .B2(
        data_in[7]), .ZN(n16374) );
  INV_X1 U12067 ( .A(n16375), .ZN(n19810) );
  AOI22_X1 U12068 ( .A1(\mem[787][0] ), .A2(n16376), .B1(n26343), .B2(
        data_in[0]), .ZN(n16375) );
  INV_X1 U12069 ( .A(n16377), .ZN(n19809) );
  AOI22_X1 U12070 ( .A1(\mem[787][1] ), .A2(n16376), .B1(n26343), .B2(
        data_in[1]), .ZN(n16377) );
  INV_X1 U12071 ( .A(n16378), .ZN(n19808) );
  AOI22_X1 U12072 ( .A1(\mem[787][2] ), .A2(n16376), .B1(n26343), .B2(
        data_in[2]), .ZN(n16378) );
  INV_X1 U12073 ( .A(n16379), .ZN(n19807) );
  AOI22_X1 U12074 ( .A1(\mem[787][3] ), .A2(n16376), .B1(n26343), .B2(
        data_in[3]), .ZN(n16379) );
  INV_X1 U12075 ( .A(n16380), .ZN(n19806) );
  AOI22_X1 U12076 ( .A1(\mem[787][4] ), .A2(n16376), .B1(n26343), .B2(
        data_in[4]), .ZN(n16380) );
  INV_X1 U12077 ( .A(n16381), .ZN(n19805) );
  AOI22_X1 U12078 ( .A1(\mem[787][5] ), .A2(n16376), .B1(n26343), .B2(
        data_in[5]), .ZN(n16381) );
  INV_X1 U12079 ( .A(n16382), .ZN(n19804) );
  AOI22_X1 U12080 ( .A1(\mem[787][6] ), .A2(n16376), .B1(n26343), .B2(
        data_in[6]), .ZN(n16382) );
  INV_X1 U12081 ( .A(n16383), .ZN(n19803) );
  AOI22_X1 U12082 ( .A1(\mem[787][7] ), .A2(n16376), .B1(n26343), .B2(
        data_in[7]), .ZN(n16383) );
  INV_X1 U12083 ( .A(n16384), .ZN(n19802) );
  AOI22_X1 U12084 ( .A1(\mem[788][0] ), .A2(n16385), .B1(n26342), .B2(
        data_in[0]), .ZN(n16384) );
  INV_X1 U12085 ( .A(n16386), .ZN(n19801) );
  AOI22_X1 U12086 ( .A1(\mem[788][1] ), .A2(n16385), .B1(n26342), .B2(
        data_in[1]), .ZN(n16386) );
  INV_X1 U12087 ( .A(n16387), .ZN(n19800) );
  AOI22_X1 U12088 ( .A1(\mem[788][2] ), .A2(n16385), .B1(n26342), .B2(
        data_in[2]), .ZN(n16387) );
  INV_X1 U12089 ( .A(n16388), .ZN(n19799) );
  AOI22_X1 U12090 ( .A1(\mem[788][3] ), .A2(n16385), .B1(n26342), .B2(
        data_in[3]), .ZN(n16388) );
  INV_X1 U12091 ( .A(n16389), .ZN(n19798) );
  AOI22_X1 U12092 ( .A1(\mem[788][4] ), .A2(n16385), .B1(n26342), .B2(
        data_in[4]), .ZN(n16389) );
  INV_X1 U12093 ( .A(n16390), .ZN(n19797) );
  AOI22_X1 U12094 ( .A1(\mem[788][5] ), .A2(n16385), .B1(n26342), .B2(
        data_in[5]), .ZN(n16390) );
  INV_X1 U12095 ( .A(n16391), .ZN(n19796) );
  AOI22_X1 U12096 ( .A1(\mem[788][6] ), .A2(n16385), .B1(n26342), .B2(
        data_in[6]), .ZN(n16391) );
  INV_X1 U12097 ( .A(n16392), .ZN(n19795) );
  AOI22_X1 U12098 ( .A1(\mem[788][7] ), .A2(n16385), .B1(n26342), .B2(
        data_in[7]), .ZN(n16392) );
  INV_X1 U12099 ( .A(n16393), .ZN(n19794) );
  AOI22_X1 U12100 ( .A1(\mem[789][0] ), .A2(n16394), .B1(n26341), .B2(
        data_in[0]), .ZN(n16393) );
  INV_X1 U12101 ( .A(n16395), .ZN(n19793) );
  AOI22_X1 U12102 ( .A1(\mem[789][1] ), .A2(n16394), .B1(n26341), .B2(
        data_in[1]), .ZN(n16395) );
  INV_X1 U12103 ( .A(n16396), .ZN(n19792) );
  AOI22_X1 U12104 ( .A1(\mem[789][2] ), .A2(n16394), .B1(n26341), .B2(
        data_in[2]), .ZN(n16396) );
  INV_X1 U12105 ( .A(n16397), .ZN(n19791) );
  AOI22_X1 U12106 ( .A1(\mem[789][3] ), .A2(n16394), .B1(n26341), .B2(
        data_in[3]), .ZN(n16397) );
  INV_X1 U12107 ( .A(n16398), .ZN(n19790) );
  AOI22_X1 U12108 ( .A1(\mem[789][4] ), .A2(n16394), .B1(n26341), .B2(
        data_in[4]), .ZN(n16398) );
  INV_X1 U12109 ( .A(n16399), .ZN(n19789) );
  AOI22_X1 U12110 ( .A1(\mem[789][5] ), .A2(n16394), .B1(n26341), .B2(
        data_in[5]), .ZN(n16399) );
  INV_X1 U12111 ( .A(n16400), .ZN(n19788) );
  AOI22_X1 U12112 ( .A1(\mem[789][6] ), .A2(n16394), .B1(n26341), .B2(
        data_in[6]), .ZN(n16400) );
  INV_X1 U12113 ( .A(n16401), .ZN(n19787) );
  AOI22_X1 U12114 ( .A1(\mem[789][7] ), .A2(n16394), .B1(n26341), .B2(
        data_in[7]), .ZN(n16401) );
  INV_X1 U12115 ( .A(n16402), .ZN(n19786) );
  AOI22_X1 U12116 ( .A1(\mem[790][0] ), .A2(n16403), .B1(n26340), .B2(
        data_in[0]), .ZN(n16402) );
  INV_X1 U12117 ( .A(n16404), .ZN(n19785) );
  AOI22_X1 U12118 ( .A1(\mem[790][1] ), .A2(n16403), .B1(n26340), .B2(
        data_in[1]), .ZN(n16404) );
  INV_X1 U12119 ( .A(n16405), .ZN(n19784) );
  AOI22_X1 U12120 ( .A1(\mem[790][2] ), .A2(n16403), .B1(n26340), .B2(
        data_in[2]), .ZN(n16405) );
  INV_X1 U12121 ( .A(n16406), .ZN(n19783) );
  AOI22_X1 U12122 ( .A1(\mem[790][3] ), .A2(n16403), .B1(n26340), .B2(
        data_in[3]), .ZN(n16406) );
  INV_X1 U12123 ( .A(n16407), .ZN(n19782) );
  AOI22_X1 U12124 ( .A1(\mem[790][4] ), .A2(n16403), .B1(n26340), .B2(
        data_in[4]), .ZN(n16407) );
  INV_X1 U12125 ( .A(n16408), .ZN(n19781) );
  AOI22_X1 U12126 ( .A1(\mem[790][5] ), .A2(n16403), .B1(n26340), .B2(
        data_in[5]), .ZN(n16408) );
  INV_X1 U12127 ( .A(n16409), .ZN(n19780) );
  AOI22_X1 U12128 ( .A1(\mem[790][6] ), .A2(n16403), .B1(n26340), .B2(
        data_in[6]), .ZN(n16409) );
  INV_X1 U12129 ( .A(n16410), .ZN(n19779) );
  AOI22_X1 U12130 ( .A1(\mem[790][7] ), .A2(n16403), .B1(n26340), .B2(
        data_in[7]), .ZN(n16410) );
  INV_X1 U12131 ( .A(n16411), .ZN(n19778) );
  AOI22_X1 U12132 ( .A1(\mem[791][0] ), .A2(n16412), .B1(n26339), .B2(
        data_in[0]), .ZN(n16411) );
  INV_X1 U12133 ( .A(n16413), .ZN(n19777) );
  AOI22_X1 U12134 ( .A1(\mem[791][1] ), .A2(n16412), .B1(n26339), .B2(
        data_in[1]), .ZN(n16413) );
  INV_X1 U12135 ( .A(n16414), .ZN(n19776) );
  AOI22_X1 U12136 ( .A1(\mem[791][2] ), .A2(n16412), .B1(n26339), .B2(
        data_in[2]), .ZN(n16414) );
  INV_X1 U12137 ( .A(n16415), .ZN(n19775) );
  AOI22_X1 U12138 ( .A1(\mem[791][3] ), .A2(n16412), .B1(n26339), .B2(
        data_in[3]), .ZN(n16415) );
  INV_X1 U12139 ( .A(n16416), .ZN(n19774) );
  AOI22_X1 U12140 ( .A1(\mem[791][4] ), .A2(n16412), .B1(n26339), .B2(
        data_in[4]), .ZN(n16416) );
  INV_X1 U12141 ( .A(n16417), .ZN(n19773) );
  AOI22_X1 U12142 ( .A1(\mem[791][5] ), .A2(n16412), .B1(n26339), .B2(
        data_in[5]), .ZN(n16417) );
  INV_X1 U12143 ( .A(n16418), .ZN(n19772) );
  AOI22_X1 U12144 ( .A1(\mem[791][6] ), .A2(n16412), .B1(n26339), .B2(
        data_in[6]), .ZN(n16418) );
  INV_X1 U12145 ( .A(n16419), .ZN(n19771) );
  AOI22_X1 U12146 ( .A1(\mem[791][7] ), .A2(n16412), .B1(n26339), .B2(
        data_in[7]), .ZN(n16419) );
  INV_X1 U12147 ( .A(n16420), .ZN(n19770) );
  AOI22_X1 U12148 ( .A1(\mem[792][0] ), .A2(n16421), .B1(n26338), .B2(
        data_in[0]), .ZN(n16420) );
  INV_X1 U12149 ( .A(n16422), .ZN(n19769) );
  AOI22_X1 U12150 ( .A1(\mem[792][1] ), .A2(n16421), .B1(n26338), .B2(
        data_in[1]), .ZN(n16422) );
  INV_X1 U12151 ( .A(n16423), .ZN(n19768) );
  AOI22_X1 U12152 ( .A1(\mem[792][2] ), .A2(n16421), .B1(n26338), .B2(
        data_in[2]), .ZN(n16423) );
  INV_X1 U12153 ( .A(n16424), .ZN(n19767) );
  AOI22_X1 U12154 ( .A1(\mem[792][3] ), .A2(n16421), .B1(n26338), .B2(
        data_in[3]), .ZN(n16424) );
  INV_X1 U12155 ( .A(n16425), .ZN(n19766) );
  AOI22_X1 U12156 ( .A1(\mem[792][4] ), .A2(n16421), .B1(n26338), .B2(
        data_in[4]), .ZN(n16425) );
  INV_X1 U12157 ( .A(n16426), .ZN(n19765) );
  AOI22_X1 U12158 ( .A1(\mem[792][5] ), .A2(n16421), .B1(n26338), .B2(
        data_in[5]), .ZN(n16426) );
  INV_X1 U12159 ( .A(n16427), .ZN(n19764) );
  AOI22_X1 U12160 ( .A1(\mem[792][6] ), .A2(n16421), .B1(n26338), .B2(
        data_in[6]), .ZN(n16427) );
  INV_X1 U12161 ( .A(n16428), .ZN(n19763) );
  AOI22_X1 U12162 ( .A1(\mem[792][7] ), .A2(n16421), .B1(n26338), .B2(
        data_in[7]), .ZN(n16428) );
  INV_X1 U12163 ( .A(n16429), .ZN(n19762) );
  AOI22_X1 U12164 ( .A1(\mem[793][0] ), .A2(n16430), .B1(n26337), .B2(
        data_in[0]), .ZN(n16429) );
  INV_X1 U12165 ( .A(n16431), .ZN(n19761) );
  AOI22_X1 U12166 ( .A1(\mem[793][1] ), .A2(n16430), .B1(n26337), .B2(
        data_in[1]), .ZN(n16431) );
  INV_X1 U12167 ( .A(n16432), .ZN(n19760) );
  AOI22_X1 U12168 ( .A1(\mem[793][2] ), .A2(n16430), .B1(n26337), .B2(
        data_in[2]), .ZN(n16432) );
  INV_X1 U12169 ( .A(n16433), .ZN(n19759) );
  AOI22_X1 U12170 ( .A1(\mem[793][3] ), .A2(n16430), .B1(n26337), .B2(
        data_in[3]), .ZN(n16433) );
  INV_X1 U12171 ( .A(n16434), .ZN(n19758) );
  AOI22_X1 U12172 ( .A1(\mem[793][4] ), .A2(n16430), .B1(n26337), .B2(
        data_in[4]), .ZN(n16434) );
  INV_X1 U12173 ( .A(n16435), .ZN(n19757) );
  AOI22_X1 U12174 ( .A1(\mem[793][5] ), .A2(n16430), .B1(n26337), .B2(
        data_in[5]), .ZN(n16435) );
  INV_X1 U12175 ( .A(n16436), .ZN(n19756) );
  AOI22_X1 U12176 ( .A1(\mem[793][6] ), .A2(n16430), .B1(n26337), .B2(
        data_in[6]), .ZN(n16436) );
  INV_X1 U12177 ( .A(n16437), .ZN(n19755) );
  AOI22_X1 U12178 ( .A1(\mem[793][7] ), .A2(n16430), .B1(n26337), .B2(
        data_in[7]), .ZN(n16437) );
  INV_X1 U12179 ( .A(n16438), .ZN(n19754) );
  AOI22_X1 U12180 ( .A1(\mem[794][0] ), .A2(n16439), .B1(n26336), .B2(
        data_in[0]), .ZN(n16438) );
  INV_X1 U12181 ( .A(n16440), .ZN(n19753) );
  AOI22_X1 U12182 ( .A1(\mem[794][1] ), .A2(n16439), .B1(n26336), .B2(
        data_in[1]), .ZN(n16440) );
  INV_X1 U12183 ( .A(n16441), .ZN(n19752) );
  AOI22_X1 U12184 ( .A1(\mem[794][2] ), .A2(n16439), .B1(n26336), .B2(
        data_in[2]), .ZN(n16441) );
  INV_X1 U12185 ( .A(n16442), .ZN(n19751) );
  AOI22_X1 U12186 ( .A1(\mem[794][3] ), .A2(n16439), .B1(n26336), .B2(
        data_in[3]), .ZN(n16442) );
  INV_X1 U12187 ( .A(n16443), .ZN(n19750) );
  AOI22_X1 U12188 ( .A1(\mem[794][4] ), .A2(n16439), .B1(n26336), .B2(
        data_in[4]), .ZN(n16443) );
  INV_X1 U12189 ( .A(n16444), .ZN(n19749) );
  AOI22_X1 U12190 ( .A1(\mem[794][5] ), .A2(n16439), .B1(n26336), .B2(
        data_in[5]), .ZN(n16444) );
  INV_X1 U12191 ( .A(n16445), .ZN(n19748) );
  AOI22_X1 U12192 ( .A1(\mem[794][6] ), .A2(n16439), .B1(n26336), .B2(
        data_in[6]), .ZN(n16445) );
  INV_X1 U12193 ( .A(n16446), .ZN(n19747) );
  AOI22_X1 U12194 ( .A1(\mem[794][7] ), .A2(n16439), .B1(n26336), .B2(
        data_in[7]), .ZN(n16446) );
  INV_X1 U12195 ( .A(n16447), .ZN(n19746) );
  AOI22_X1 U12196 ( .A1(\mem[795][0] ), .A2(n16448), .B1(n26335), .B2(
        data_in[0]), .ZN(n16447) );
  INV_X1 U12197 ( .A(n16449), .ZN(n19745) );
  AOI22_X1 U12198 ( .A1(\mem[795][1] ), .A2(n16448), .B1(n26335), .B2(
        data_in[1]), .ZN(n16449) );
  INV_X1 U12199 ( .A(n16450), .ZN(n19744) );
  AOI22_X1 U12200 ( .A1(\mem[795][2] ), .A2(n16448), .B1(n26335), .B2(
        data_in[2]), .ZN(n16450) );
  INV_X1 U12201 ( .A(n16451), .ZN(n19743) );
  AOI22_X1 U12202 ( .A1(\mem[795][3] ), .A2(n16448), .B1(n26335), .B2(
        data_in[3]), .ZN(n16451) );
  INV_X1 U12203 ( .A(n16452), .ZN(n19742) );
  AOI22_X1 U12204 ( .A1(\mem[795][4] ), .A2(n16448), .B1(n26335), .B2(
        data_in[4]), .ZN(n16452) );
  INV_X1 U12205 ( .A(n16453), .ZN(n19741) );
  AOI22_X1 U12206 ( .A1(\mem[795][5] ), .A2(n16448), .B1(n26335), .B2(
        data_in[5]), .ZN(n16453) );
  INV_X1 U12207 ( .A(n16454), .ZN(n19740) );
  AOI22_X1 U12208 ( .A1(\mem[795][6] ), .A2(n16448), .B1(n26335), .B2(
        data_in[6]), .ZN(n16454) );
  INV_X1 U12209 ( .A(n16455), .ZN(n19739) );
  AOI22_X1 U12210 ( .A1(\mem[795][7] ), .A2(n16448), .B1(n26335), .B2(
        data_in[7]), .ZN(n16455) );
  INV_X1 U12211 ( .A(n16456), .ZN(n19738) );
  AOI22_X1 U12212 ( .A1(\mem[796][0] ), .A2(n16457), .B1(n26334), .B2(
        data_in[0]), .ZN(n16456) );
  INV_X1 U12213 ( .A(n16458), .ZN(n19737) );
  AOI22_X1 U12214 ( .A1(\mem[796][1] ), .A2(n16457), .B1(n26334), .B2(
        data_in[1]), .ZN(n16458) );
  INV_X1 U12215 ( .A(n16459), .ZN(n19736) );
  AOI22_X1 U12216 ( .A1(\mem[796][2] ), .A2(n16457), .B1(n26334), .B2(
        data_in[2]), .ZN(n16459) );
  INV_X1 U12217 ( .A(n16460), .ZN(n19735) );
  AOI22_X1 U12218 ( .A1(\mem[796][3] ), .A2(n16457), .B1(n26334), .B2(
        data_in[3]), .ZN(n16460) );
  INV_X1 U12219 ( .A(n16461), .ZN(n19734) );
  AOI22_X1 U12220 ( .A1(\mem[796][4] ), .A2(n16457), .B1(n26334), .B2(
        data_in[4]), .ZN(n16461) );
  INV_X1 U12221 ( .A(n16462), .ZN(n19733) );
  AOI22_X1 U12222 ( .A1(\mem[796][5] ), .A2(n16457), .B1(n26334), .B2(
        data_in[5]), .ZN(n16462) );
  INV_X1 U12223 ( .A(n16463), .ZN(n19732) );
  AOI22_X1 U12224 ( .A1(\mem[796][6] ), .A2(n16457), .B1(n26334), .B2(
        data_in[6]), .ZN(n16463) );
  INV_X1 U12225 ( .A(n16464), .ZN(n19731) );
  AOI22_X1 U12226 ( .A1(\mem[796][7] ), .A2(n16457), .B1(n26334), .B2(
        data_in[7]), .ZN(n16464) );
  INV_X1 U12227 ( .A(n16465), .ZN(n19730) );
  AOI22_X1 U12228 ( .A1(\mem[797][0] ), .A2(n16466), .B1(n26333), .B2(
        data_in[0]), .ZN(n16465) );
  INV_X1 U12229 ( .A(n16467), .ZN(n19729) );
  AOI22_X1 U12230 ( .A1(\mem[797][1] ), .A2(n16466), .B1(n26333), .B2(
        data_in[1]), .ZN(n16467) );
  INV_X1 U12231 ( .A(n16468), .ZN(n19728) );
  AOI22_X1 U12232 ( .A1(\mem[797][2] ), .A2(n16466), .B1(n26333), .B2(
        data_in[2]), .ZN(n16468) );
  INV_X1 U12233 ( .A(n16469), .ZN(n19727) );
  AOI22_X1 U12234 ( .A1(\mem[797][3] ), .A2(n16466), .B1(n26333), .B2(
        data_in[3]), .ZN(n16469) );
  INV_X1 U12235 ( .A(n16470), .ZN(n19726) );
  AOI22_X1 U12236 ( .A1(\mem[797][4] ), .A2(n16466), .B1(n26333), .B2(
        data_in[4]), .ZN(n16470) );
  INV_X1 U12237 ( .A(n16471), .ZN(n19725) );
  AOI22_X1 U12238 ( .A1(\mem[797][5] ), .A2(n16466), .B1(n26333), .B2(
        data_in[5]), .ZN(n16471) );
  INV_X1 U12239 ( .A(n16472), .ZN(n19724) );
  AOI22_X1 U12240 ( .A1(\mem[797][6] ), .A2(n16466), .B1(n26333), .B2(
        data_in[6]), .ZN(n16472) );
  INV_X1 U12241 ( .A(n16473), .ZN(n19723) );
  AOI22_X1 U12242 ( .A1(\mem[797][7] ), .A2(n16466), .B1(n26333), .B2(
        data_in[7]), .ZN(n16473) );
  INV_X1 U12243 ( .A(n16474), .ZN(n19722) );
  AOI22_X1 U12244 ( .A1(\mem[798][0] ), .A2(n16475), .B1(n26332), .B2(
        data_in[0]), .ZN(n16474) );
  INV_X1 U12245 ( .A(n16476), .ZN(n19721) );
  AOI22_X1 U12246 ( .A1(\mem[798][1] ), .A2(n16475), .B1(n26332), .B2(
        data_in[1]), .ZN(n16476) );
  INV_X1 U12247 ( .A(n16477), .ZN(n19720) );
  AOI22_X1 U12248 ( .A1(\mem[798][2] ), .A2(n16475), .B1(n26332), .B2(
        data_in[2]), .ZN(n16477) );
  INV_X1 U12249 ( .A(n16478), .ZN(n19719) );
  AOI22_X1 U12250 ( .A1(\mem[798][3] ), .A2(n16475), .B1(n26332), .B2(
        data_in[3]), .ZN(n16478) );
  INV_X1 U12251 ( .A(n16479), .ZN(n19718) );
  AOI22_X1 U12252 ( .A1(\mem[798][4] ), .A2(n16475), .B1(n26332), .B2(
        data_in[4]), .ZN(n16479) );
  INV_X1 U12253 ( .A(n16480), .ZN(n19717) );
  AOI22_X1 U12254 ( .A1(\mem[798][5] ), .A2(n16475), .B1(n26332), .B2(
        data_in[5]), .ZN(n16480) );
  INV_X1 U12255 ( .A(n16481), .ZN(n19716) );
  AOI22_X1 U12256 ( .A1(\mem[798][6] ), .A2(n16475), .B1(n26332), .B2(
        data_in[6]), .ZN(n16481) );
  INV_X1 U12257 ( .A(n16482), .ZN(n19715) );
  AOI22_X1 U12258 ( .A1(\mem[798][7] ), .A2(n16475), .B1(n26332), .B2(
        data_in[7]), .ZN(n16482) );
  INV_X1 U12259 ( .A(n16483), .ZN(n19714) );
  AOI22_X1 U12260 ( .A1(\mem[799][0] ), .A2(n16484), .B1(n26331), .B2(
        data_in[0]), .ZN(n16483) );
  INV_X1 U12261 ( .A(n16485), .ZN(n19713) );
  AOI22_X1 U12262 ( .A1(\mem[799][1] ), .A2(n16484), .B1(n26331), .B2(
        data_in[1]), .ZN(n16485) );
  INV_X1 U12263 ( .A(n16486), .ZN(n19712) );
  AOI22_X1 U12264 ( .A1(\mem[799][2] ), .A2(n16484), .B1(n26331), .B2(
        data_in[2]), .ZN(n16486) );
  INV_X1 U12265 ( .A(n16487), .ZN(n19711) );
  AOI22_X1 U12266 ( .A1(\mem[799][3] ), .A2(n16484), .B1(n26331), .B2(
        data_in[3]), .ZN(n16487) );
  INV_X1 U12267 ( .A(n16488), .ZN(n19710) );
  AOI22_X1 U12268 ( .A1(\mem[799][4] ), .A2(n16484), .B1(n26331), .B2(
        data_in[4]), .ZN(n16488) );
  INV_X1 U12269 ( .A(n16489), .ZN(n19709) );
  AOI22_X1 U12270 ( .A1(\mem[799][5] ), .A2(n16484), .B1(n26331), .B2(
        data_in[5]), .ZN(n16489) );
  INV_X1 U12271 ( .A(n16490), .ZN(n19708) );
  AOI22_X1 U12272 ( .A1(\mem[799][6] ), .A2(n16484), .B1(n26331), .B2(
        data_in[6]), .ZN(n16490) );
  INV_X1 U12273 ( .A(n16491), .ZN(n19707) );
  AOI22_X1 U12274 ( .A1(\mem[799][7] ), .A2(n16484), .B1(n26331), .B2(
        data_in[7]), .ZN(n16491) );
  INV_X1 U12275 ( .A(n16566), .ZN(n19642) );
  AOI22_X1 U12276 ( .A1(\mem[808][0] ), .A2(n16567), .B1(n26322), .B2(
        data_in[0]), .ZN(n16566) );
  INV_X1 U12277 ( .A(n16568), .ZN(n19641) );
  AOI22_X1 U12278 ( .A1(\mem[808][1] ), .A2(n16567), .B1(n26322), .B2(
        data_in[1]), .ZN(n16568) );
  INV_X1 U12279 ( .A(n16569), .ZN(n19640) );
  AOI22_X1 U12280 ( .A1(\mem[808][2] ), .A2(n16567), .B1(n26322), .B2(
        data_in[2]), .ZN(n16569) );
  INV_X1 U12281 ( .A(n16570), .ZN(n19639) );
  AOI22_X1 U12282 ( .A1(\mem[808][3] ), .A2(n16567), .B1(n26322), .B2(
        data_in[3]), .ZN(n16570) );
  INV_X1 U12283 ( .A(n16571), .ZN(n19638) );
  AOI22_X1 U12284 ( .A1(\mem[808][4] ), .A2(n16567), .B1(n26322), .B2(
        data_in[4]), .ZN(n16571) );
  INV_X1 U12285 ( .A(n16572), .ZN(n19637) );
  AOI22_X1 U12286 ( .A1(\mem[808][5] ), .A2(n16567), .B1(n26322), .B2(
        data_in[5]), .ZN(n16572) );
  INV_X1 U12287 ( .A(n16573), .ZN(n19636) );
  AOI22_X1 U12288 ( .A1(\mem[808][6] ), .A2(n16567), .B1(n26322), .B2(
        data_in[6]), .ZN(n16573) );
  INV_X1 U12289 ( .A(n16574), .ZN(n19635) );
  AOI22_X1 U12290 ( .A1(\mem[808][7] ), .A2(n16567), .B1(n26322), .B2(
        data_in[7]), .ZN(n16574) );
  INV_X1 U12291 ( .A(n16575), .ZN(n19634) );
  AOI22_X1 U12292 ( .A1(\mem[809][0] ), .A2(n16576), .B1(n26321), .B2(
        data_in[0]), .ZN(n16575) );
  INV_X1 U12293 ( .A(n16577), .ZN(n19633) );
  AOI22_X1 U12294 ( .A1(\mem[809][1] ), .A2(n16576), .B1(n26321), .B2(
        data_in[1]), .ZN(n16577) );
  INV_X1 U12295 ( .A(n16578), .ZN(n19632) );
  AOI22_X1 U12296 ( .A1(\mem[809][2] ), .A2(n16576), .B1(n26321), .B2(
        data_in[2]), .ZN(n16578) );
  INV_X1 U12297 ( .A(n16579), .ZN(n19631) );
  AOI22_X1 U12298 ( .A1(\mem[809][3] ), .A2(n16576), .B1(n26321), .B2(
        data_in[3]), .ZN(n16579) );
  INV_X1 U12299 ( .A(n16580), .ZN(n19630) );
  AOI22_X1 U12300 ( .A1(\mem[809][4] ), .A2(n16576), .B1(n26321), .B2(
        data_in[4]), .ZN(n16580) );
  INV_X1 U12301 ( .A(n16581), .ZN(n19629) );
  AOI22_X1 U12302 ( .A1(\mem[809][5] ), .A2(n16576), .B1(n26321), .B2(
        data_in[5]), .ZN(n16581) );
  INV_X1 U12303 ( .A(n16582), .ZN(n19628) );
  AOI22_X1 U12304 ( .A1(\mem[809][6] ), .A2(n16576), .B1(n26321), .B2(
        data_in[6]), .ZN(n16582) );
  INV_X1 U12305 ( .A(n16583), .ZN(n19627) );
  AOI22_X1 U12306 ( .A1(\mem[809][7] ), .A2(n16576), .B1(n26321), .B2(
        data_in[7]), .ZN(n16583) );
  INV_X1 U12307 ( .A(n16584), .ZN(n19626) );
  AOI22_X1 U12308 ( .A1(\mem[810][0] ), .A2(n16585), .B1(n26320), .B2(
        data_in[0]), .ZN(n16584) );
  INV_X1 U12309 ( .A(n16586), .ZN(n19625) );
  AOI22_X1 U12310 ( .A1(\mem[810][1] ), .A2(n16585), .B1(n26320), .B2(
        data_in[1]), .ZN(n16586) );
  INV_X1 U12311 ( .A(n16587), .ZN(n19624) );
  AOI22_X1 U12312 ( .A1(\mem[810][2] ), .A2(n16585), .B1(n26320), .B2(
        data_in[2]), .ZN(n16587) );
  INV_X1 U12313 ( .A(n16588), .ZN(n19623) );
  AOI22_X1 U12314 ( .A1(\mem[810][3] ), .A2(n16585), .B1(n26320), .B2(
        data_in[3]), .ZN(n16588) );
  INV_X1 U12315 ( .A(n16589), .ZN(n19622) );
  AOI22_X1 U12316 ( .A1(\mem[810][4] ), .A2(n16585), .B1(n26320), .B2(
        data_in[4]), .ZN(n16589) );
  INV_X1 U12317 ( .A(n16590), .ZN(n19621) );
  AOI22_X1 U12318 ( .A1(\mem[810][5] ), .A2(n16585), .B1(n26320), .B2(
        data_in[5]), .ZN(n16590) );
  INV_X1 U12319 ( .A(n16591), .ZN(n19620) );
  AOI22_X1 U12320 ( .A1(\mem[810][6] ), .A2(n16585), .B1(n26320), .B2(
        data_in[6]), .ZN(n16591) );
  INV_X1 U12321 ( .A(n16592), .ZN(n19619) );
  AOI22_X1 U12322 ( .A1(\mem[810][7] ), .A2(n16585), .B1(n26320), .B2(
        data_in[7]), .ZN(n16592) );
  INV_X1 U12323 ( .A(n16593), .ZN(n19618) );
  AOI22_X1 U12324 ( .A1(\mem[811][0] ), .A2(n16594), .B1(n26319), .B2(
        data_in[0]), .ZN(n16593) );
  INV_X1 U12325 ( .A(n16595), .ZN(n19617) );
  AOI22_X1 U12326 ( .A1(\mem[811][1] ), .A2(n16594), .B1(n26319), .B2(
        data_in[1]), .ZN(n16595) );
  INV_X1 U12327 ( .A(n16596), .ZN(n19616) );
  AOI22_X1 U12328 ( .A1(\mem[811][2] ), .A2(n16594), .B1(n26319), .B2(
        data_in[2]), .ZN(n16596) );
  INV_X1 U12329 ( .A(n16597), .ZN(n19615) );
  AOI22_X1 U12330 ( .A1(\mem[811][3] ), .A2(n16594), .B1(n26319), .B2(
        data_in[3]), .ZN(n16597) );
  INV_X1 U12331 ( .A(n16598), .ZN(n19614) );
  AOI22_X1 U12332 ( .A1(\mem[811][4] ), .A2(n16594), .B1(n26319), .B2(
        data_in[4]), .ZN(n16598) );
  INV_X1 U12333 ( .A(n16599), .ZN(n19613) );
  AOI22_X1 U12334 ( .A1(\mem[811][5] ), .A2(n16594), .B1(n26319), .B2(
        data_in[5]), .ZN(n16599) );
  INV_X1 U12335 ( .A(n16600), .ZN(n19612) );
  AOI22_X1 U12336 ( .A1(\mem[811][6] ), .A2(n16594), .B1(n26319), .B2(
        data_in[6]), .ZN(n16600) );
  INV_X1 U12337 ( .A(n16601), .ZN(n19611) );
  AOI22_X1 U12338 ( .A1(\mem[811][7] ), .A2(n16594), .B1(n26319), .B2(
        data_in[7]), .ZN(n16601) );
  INV_X1 U12339 ( .A(n16602), .ZN(n19610) );
  AOI22_X1 U12340 ( .A1(\mem[812][0] ), .A2(n16603), .B1(n26318), .B2(
        data_in[0]), .ZN(n16602) );
  INV_X1 U12341 ( .A(n16604), .ZN(n19609) );
  AOI22_X1 U12342 ( .A1(\mem[812][1] ), .A2(n16603), .B1(n26318), .B2(
        data_in[1]), .ZN(n16604) );
  INV_X1 U12343 ( .A(n16605), .ZN(n19608) );
  AOI22_X1 U12344 ( .A1(\mem[812][2] ), .A2(n16603), .B1(n26318), .B2(
        data_in[2]), .ZN(n16605) );
  INV_X1 U12345 ( .A(n16606), .ZN(n19607) );
  AOI22_X1 U12346 ( .A1(\mem[812][3] ), .A2(n16603), .B1(n26318), .B2(
        data_in[3]), .ZN(n16606) );
  INV_X1 U12347 ( .A(n16607), .ZN(n19606) );
  AOI22_X1 U12348 ( .A1(\mem[812][4] ), .A2(n16603), .B1(n26318), .B2(
        data_in[4]), .ZN(n16607) );
  INV_X1 U12349 ( .A(n16608), .ZN(n19605) );
  AOI22_X1 U12350 ( .A1(\mem[812][5] ), .A2(n16603), .B1(n26318), .B2(
        data_in[5]), .ZN(n16608) );
  INV_X1 U12351 ( .A(n16609), .ZN(n19604) );
  AOI22_X1 U12352 ( .A1(\mem[812][6] ), .A2(n16603), .B1(n26318), .B2(
        data_in[6]), .ZN(n16609) );
  INV_X1 U12353 ( .A(n16610), .ZN(n19603) );
  AOI22_X1 U12354 ( .A1(\mem[812][7] ), .A2(n16603), .B1(n26318), .B2(
        data_in[7]), .ZN(n16610) );
  INV_X1 U12355 ( .A(n16611), .ZN(n19602) );
  AOI22_X1 U12356 ( .A1(\mem[813][0] ), .A2(n16612), .B1(n26317), .B2(
        data_in[0]), .ZN(n16611) );
  INV_X1 U12357 ( .A(n16613), .ZN(n19601) );
  AOI22_X1 U12358 ( .A1(\mem[813][1] ), .A2(n16612), .B1(n26317), .B2(
        data_in[1]), .ZN(n16613) );
  INV_X1 U12359 ( .A(n16614), .ZN(n19600) );
  AOI22_X1 U12360 ( .A1(\mem[813][2] ), .A2(n16612), .B1(n26317), .B2(
        data_in[2]), .ZN(n16614) );
  INV_X1 U12361 ( .A(n16615), .ZN(n19599) );
  AOI22_X1 U12362 ( .A1(\mem[813][3] ), .A2(n16612), .B1(n26317), .B2(
        data_in[3]), .ZN(n16615) );
  INV_X1 U12363 ( .A(n16616), .ZN(n19598) );
  AOI22_X1 U12364 ( .A1(\mem[813][4] ), .A2(n16612), .B1(n26317), .B2(
        data_in[4]), .ZN(n16616) );
  INV_X1 U12365 ( .A(n16617), .ZN(n19597) );
  AOI22_X1 U12366 ( .A1(\mem[813][5] ), .A2(n16612), .B1(n26317), .B2(
        data_in[5]), .ZN(n16617) );
  INV_X1 U12367 ( .A(n16618), .ZN(n19596) );
  AOI22_X1 U12368 ( .A1(\mem[813][6] ), .A2(n16612), .B1(n26317), .B2(
        data_in[6]), .ZN(n16618) );
  INV_X1 U12369 ( .A(n16619), .ZN(n19595) );
  AOI22_X1 U12370 ( .A1(\mem[813][7] ), .A2(n16612), .B1(n26317), .B2(
        data_in[7]), .ZN(n16619) );
  INV_X1 U12371 ( .A(n16620), .ZN(n19594) );
  AOI22_X1 U12372 ( .A1(\mem[814][0] ), .A2(n16621), .B1(n26316), .B2(
        data_in[0]), .ZN(n16620) );
  INV_X1 U12373 ( .A(n16622), .ZN(n19593) );
  AOI22_X1 U12374 ( .A1(\mem[814][1] ), .A2(n16621), .B1(n26316), .B2(
        data_in[1]), .ZN(n16622) );
  INV_X1 U12375 ( .A(n16623), .ZN(n19592) );
  AOI22_X1 U12376 ( .A1(\mem[814][2] ), .A2(n16621), .B1(n26316), .B2(
        data_in[2]), .ZN(n16623) );
  INV_X1 U12377 ( .A(n16624), .ZN(n19591) );
  AOI22_X1 U12378 ( .A1(\mem[814][3] ), .A2(n16621), .B1(n26316), .B2(
        data_in[3]), .ZN(n16624) );
  INV_X1 U12379 ( .A(n16625), .ZN(n19590) );
  AOI22_X1 U12380 ( .A1(\mem[814][4] ), .A2(n16621), .B1(n26316), .B2(
        data_in[4]), .ZN(n16625) );
  INV_X1 U12381 ( .A(n16626), .ZN(n19589) );
  AOI22_X1 U12382 ( .A1(\mem[814][5] ), .A2(n16621), .B1(n26316), .B2(
        data_in[5]), .ZN(n16626) );
  INV_X1 U12383 ( .A(n16627), .ZN(n19588) );
  AOI22_X1 U12384 ( .A1(\mem[814][6] ), .A2(n16621), .B1(n26316), .B2(
        data_in[6]), .ZN(n16627) );
  INV_X1 U12385 ( .A(n16628), .ZN(n19587) );
  AOI22_X1 U12386 ( .A1(\mem[814][7] ), .A2(n16621), .B1(n26316), .B2(
        data_in[7]), .ZN(n16628) );
  INV_X1 U12387 ( .A(n16629), .ZN(n19586) );
  AOI22_X1 U12388 ( .A1(\mem[815][0] ), .A2(n16630), .B1(n26315), .B2(
        data_in[0]), .ZN(n16629) );
  INV_X1 U12389 ( .A(n16631), .ZN(n19585) );
  AOI22_X1 U12390 ( .A1(\mem[815][1] ), .A2(n16630), .B1(n26315), .B2(
        data_in[1]), .ZN(n16631) );
  INV_X1 U12391 ( .A(n16632), .ZN(n19584) );
  AOI22_X1 U12392 ( .A1(\mem[815][2] ), .A2(n16630), .B1(n26315), .B2(
        data_in[2]), .ZN(n16632) );
  INV_X1 U12393 ( .A(n16633), .ZN(n19583) );
  AOI22_X1 U12394 ( .A1(\mem[815][3] ), .A2(n16630), .B1(n26315), .B2(
        data_in[3]), .ZN(n16633) );
  INV_X1 U12395 ( .A(n16634), .ZN(n19582) );
  AOI22_X1 U12396 ( .A1(\mem[815][4] ), .A2(n16630), .B1(n26315), .B2(
        data_in[4]), .ZN(n16634) );
  INV_X1 U12397 ( .A(n16635), .ZN(n19581) );
  AOI22_X1 U12398 ( .A1(\mem[815][5] ), .A2(n16630), .B1(n26315), .B2(
        data_in[5]), .ZN(n16635) );
  INV_X1 U12399 ( .A(n16636), .ZN(n19580) );
  AOI22_X1 U12400 ( .A1(\mem[815][6] ), .A2(n16630), .B1(n26315), .B2(
        data_in[6]), .ZN(n16636) );
  INV_X1 U12401 ( .A(n16637), .ZN(n19579) );
  AOI22_X1 U12402 ( .A1(\mem[815][7] ), .A2(n16630), .B1(n26315), .B2(
        data_in[7]), .ZN(n16637) );
  INV_X1 U12403 ( .A(n16638), .ZN(n19578) );
  AOI22_X1 U12404 ( .A1(\mem[816][0] ), .A2(n16639), .B1(n26314), .B2(
        data_in[0]), .ZN(n16638) );
  INV_X1 U12405 ( .A(n16640), .ZN(n19577) );
  AOI22_X1 U12406 ( .A1(\mem[816][1] ), .A2(n16639), .B1(n26314), .B2(
        data_in[1]), .ZN(n16640) );
  INV_X1 U12407 ( .A(n16641), .ZN(n19576) );
  AOI22_X1 U12408 ( .A1(\mem[816][2] ), .A2(n16639), .B1(n26314), .B2(
        data_in[2]), .ZN(n16641) );
  INV_X1 U12409 ( .A(n16642), .ZN(n19575) );
  AOI22_X1 U12410 ( .A1(\mem[816][3] ), .A2(n16639), .B1(n26314), .B2(
        data_in[3]), .ZN(n16642) );
  INV_X1 U12411 ( .A(n16643), .ZN(n19574) );
  AOI22_X1 U12412 ( .A1(\mem[816][4] ), .A2(n16639), .B1(n26314), .B2(
        data_in[4]), .ZN(n16643) );
  INV_X1 U12413 ( .A(n16644), .ZN(n19573) );
  AOI22_X1 U12414 ( .A1(\mem[816][5] ), .A2(n16639), .B1(n26314), .B2(
        data_in[5]), .ZN(n16644) );
  INV_X1 U12415 ( .A(n16645), .ZN(n19572) );
  AOI22_X1 U12416 ( .A1(\mem[816][6] ), .A2(n16639), .B1(n26314), .B2(
        data_in[6]), .ZN(n16645) );
  INV_X1 U12417 ( .A(n16646), .ZN(n19571) );
  AOI22_X1 U12418 ( .A1(\mem[816][7] ), .A2(n16639), .B1(n26314), .B2(
        data_in[7]), .ZN(n16646) );
  INV_X1 U12419 ( .A(n16647), .ZN(n19570) );
  AOI22_X1 U12420 ( .A1(\mem[817][0] ), .A2(n16648), .B1(n26313), .B2(
        data_in[0]), .ZN(n16647) );
  INV_X1 U12421 ( .A(n16649), .ZN(n19569) );
  AOI22_X1 U12422 ( .A1(\mem[817][1] ), .A2(n16648), .B1(n26313), .B2(
        data_in[1]), .ZN(n16649) );
  INV_X1 U12423 ( .A(n16650), .ZN(n19568) );
  AOI22_X1 U12424 ( .A1(\mem[817][2] ), .A2(n16648), .B1(n26313), .B2(
        data_in[2]), .ZN(n16650) );
  INV_X1 U12425 ( .A(n16651), .ZN(n19567) );
  AOI22_X1 U12426 ( .A1(\mem[817][3] ), .A2(n16648), .B1(n26313), .B2(
        data_in[3]), .ZN(n16651) );
  INV_X1 U12427 ( .A(n16652), .ZN(n19566) );
  AOI22_X1 U12428 ( .A1(\mem[817][4] ), .A2(n16648), .B1(n26313), .B2(
        data_in[4]), .ZN(n16652) );
  INV_X1 U12429 ( .A(n16653), .ZN(n19565) );
  AOI22_X1 U12430 ( .A1(\mem[817][5] ), .A2(n16648), .B1(n26313), .B2(
        data_in[5]), .ZN(n16653) );
  INV_X1 U12431 ( .A(n16654), .ZN(n19564) );
  AOI22_X1 U12432 ( .A1(\mem[817][6] ), .A2(n16648), .B1(n26313), .B2(
        data_in[6]), .ZN(n16654) );
  INV_X1 U12433 ( .A(n16655), .ZN(n19563) );
  AOI22_X1 U12434 ( .A1(\mem[817][7] ), .A2(n16648), .B1(n26313), .B2(
        data_in[7]), .ZN(n16655) );
  INV_X1 U12435 ( .A(n16656), .ZN(n19562) );
  AOI22_X1 U12436 ( .A1(\mem[818][0] ), .A2(n16657), .B1(n26312), .B2(
        data_in[0]), .ZN(n16656) );
  INV_X1 U12437 ( .A(n16658), .ZN(n19561) );
  AOI22_X1 U12438 ( .A1(\mem[818][1] ), .A2(n16657), .B1(n26312), .B2(
        data_in[1]), .ZN(n16658) );
  INV_X1 U12439 ( .A(n16659), .ZN(n19560) );
  AOI22_X1 U12440 ( .A1(\mem[818][2] ), .A2(n16657), .B1(n26312), .B2(
        data_in[2]), .ZN(n16659) );
  INV_X1 U12441 ( .A(n16660), .ZN(n19559) );
  AOI22_X1 U12442 ( .A1(\mem[818][3] ), .A2(n16657), .B1(n26312), .B2(
        data_in[3]), .ZN(n16660) );
  INV_X1 U12443 ( .A(n16661), .ZN(n19558) );
  AOI22_X1 U12444 ( .A1(\mem[818][4] ), .A2(n16657), .B1(n26312), .B2(
        data_in[4]), .ZN(n16661) );
  INV_X1 U12445 ( .A(n16662), .ZN(n19557) );
  AOI22_X1 U12446 ( .A1(\mem[818][5] ), .A2(n16657), .B1(n26312), .B2(
        data_in[5]), .ZN(n16662) );
  INV_X1 U12447 ( .A(n16663), .ZN(n19556) );
  AOI22_X1 U12448 ( .A1(\mem[818][6] ), .A2(n16657), .B1(n26312), .B2(
        data_in[6]), .ZN(n16663) );
  INV_X1 U12449 ( .A(n16664), .ZN(n19555) );
  AOI22_X1 U12450 ( .A1(\mem[818][7] ), .A2(n16657), .B1(n26312), .B2(
        data_in[7]), .ZN(n16664) );
  INV_X1 U12451 ( .A(n16665), .ZN(n19554) );
  AOI22_X1 U12452 ( .A1(\mem[819][0] ), .A2(n16666), .B1(n26311), .B2(
        data_in[0]), .ZN(n16665) );
  INV_X1 U12453 ( .A(n16667), .ZN(n19553) );
  AOI22_X1 U12454 ( .A1(\mem[819][1] ), .A2(n16666), .B1(n26311), .B2(
        data_in[1]), .ZN(n16667) );
  INV_X1 U12455 ( .A(n16668), .ZN(n19552) );
  AOI22_X1 U12456 ( .A1(\mem[819][2] ), .A2(n16666), .B1(n26311), .B2(
        data_in[2]), .ZN(n16668) );
  INV_X1 U12457 ( .A(n16669), .ZN(n19551) );
  AOI22_X1 U12458 ( .A1(\mem[819][3] ), .A2(n16666), .B1(n26311), .B2(
        data_in[3]), .ZN(n16669) );
  INV_X1 U12459 ( .A(n16670), .ZN(n19550) );
  AOI22_X1 U12460 ( .A1(\mem[819][4] ), .A2(n16666), .B1(n26311), .B2(
        data_in[4]), .ZN(n16670) );
  INV_X1 U12461 ( .A(n16671), .ZN(n19549) );
  AOI22_X1 U12462 ( .A1(\mem[819][5] ), .A2(n16666), .B1(n26311), .B2(
        data_in[5]), .ZN(n16671) );
  INV_X1 U12463 ( .A(n16672), .ZN(n19548) );
  AOI22_X1 U12464 ( .A1(\mem[819][6] ), .A2(n16666), .B1(n26311), .B2(
        data_in[6]), .ZN(n16672) );
  INV_X1 U12465 ( .A(n16673), .ZN(n19547) );
  AOI22_X1 U12466 ( .A1(\mem[819][7] ), .A2(n16666), .B1(n26311), .B2(
        data_in[7]), .ZN(n16673) );
  INV_X1 U12467 ( .A(n16674), .ZN(n19546) );
  AOI22_X1 U12468 ( .A1(\mem[820][0] ), .A2(n16675), .B1(n26310), .B2(
        data_in[0]), .ZN(n16674) );
  INV_X1 U12469 ( .A(n16676), .ZN(n19545) );
  AOI22_X1 U12470 ( .A1(\mem[820][1] ), .A2(n16675), .B1(n26310), .B2(
        data_in[1]), .ZN(n16676) );
  INV_X1 U12471 ( .A(n16677), .ZN(n19544) );
  AOI22_X1 U12472 ( .A1(\mem[820][2] ), .A2(n16675), .B1(n26310), .B2(
        data_in[2]), .ZN(n16677) );
  INV_X1 U12473 ( .A(n16678), .ZN(n19543) );
  AOI22_X1 U12474 ( .A1(\mem[820][3] ), .A2(n16675), .B1(n26310), .B2(
        data_in[3]), .ZN(n16678) );
  INV_X1 U12475 ( .A(n16679), .ZN(n19542) );
  AOI22_X1 U12476 ( .A1(\mem[820][4] ), .A2(n16675), .B1(n26310), .B2(
        data_in[4]), .ZN(n16679) );
  INV_X1 U12477 ( .A(n16680), .ZN(n19541) );
  AOI22_X1 U12478 ( .A1(\mem[820][5] ), .A2(n16675), .B1(n26310), .B2(
        data_in[5]), .ZN(n16680) );
  INV_X1 U12479 ( .A(n16681), .ZN(n19540) );
  AOI22_X1 U12480 ( .A1(\mem[820][6] ), .A2(n16675), .B1(n26310), .B2(
        data_in[6]), .ZN(n16681) );
  INV_X1 U12481 ( .A(n16682), .ZN(n19539) );
  AOI22_X1 U12482 ( .A1(\mem[820][7] ), .A2(n16675), .B1(n26310), .B2(
        data_in[7]), .ZN(n16682) );
  INV_X1 U12483 ( .A(n16683), .ZN(n19538) );
  AOI22_X1 U12484 ( .A1(\mem[821][0] ), .A2(n16684), .B1(n26309), .B2(
        data_in[0]), .ZN(n16683) );
  INV_X1 U12485 ( .A(n16685), .ZN(n19537) );
  AOI22_X1 U12486 ( .A1(\mem[821][1] ), .A2(n16684), .B1(n26309), .B2(
        data_in[1]), .ZN(n16685) );
  INV_X1 U12487 ( .A(n16686), .ZN(n19536) );
  AOI22_X1 U12488 ( .A1(\mem[821][2] ), .A2(n16684), .B1(n26309), .B2(
        data_in[2]), .ZN(n16686) );
  INV_X1 U12489 ( .A(n16687), .ZN(n19535) );
  AOI22_X1 U12490 ( .A1(\mem[821][3] ), .A2(n16684), .B1(n26309), .B2(
        data_in[3]), .ZN(n16687) );
  INV_X1 U12491 ( .A(n16688), .ZN(n19534) );
  AOI22_X1 U12492 ( .A1(\mem[821][4] ), .A2(n16684), .B1(n26309), .B2(
        data_in[4]), .ZN(n16688) );
  INV_X1 U12493 ( .A(n16689), .ZN(n19533) );
  AOI22_X1 U12494 ( .A1(\mem[821][5] ), .A2(n16684), .B1(n26309), .B2(
        data_in[5]), .ZN(n16689) );
  INV_X1 U12495 ( .A(n16690), .ZN(n19532) );
  AOI22_X1 U12496 ( .A1(\mem[821][6] ), .A2(n16684), .B1(n26309), .B2(
        data_in[6]), .ZN(n16690) );
  INV_X1 U12497 ( .A(n16691), .ZN(n19531) );
  AOI22_X1 U12498 ( .A1(\mem[821][7] ), .A2(n16684), .B1(n26309), .B2(
        data_in[7]), .ZN(n16691) );
  INV_X1 U12499 ( .A(n16692), .ZN(n19530) );
  AOI22_X1 U12500 ( .A1(\mem[822][0] ), .A2(n16693), .B1(n26308), .B2(
        data_in[0]), .ZN(n16692) );
  INV_X1 U12501 ( .A(n16694), .ZN(n19529) );
  AOI22_X1 U12502 ( .A1(\mem[822][1] ), .A2(n16693), .B1(n26308), .B2(
        data_in[1]), .ZN(n16694) );
  INV_X1 U12503 ( .A(n16695), .ZN(n19528) );
  AOI22_X1 U12504 ( .A1(\mem[822][2] ), .A2(n16693), .B1(n26308), .B2(
        data_in[2]), .ZN(n16695) );
  INV_X1 U12505 ( .A(n16696), .ZN(n19527) );
  AOI22_X1 U12506 ( .A1(\mem[822][3] ), .A2(n16693), .B1(n26308), .B2(
        data_in[3]), .ZN(n16696) );
  INV_X1 U12507 ( .A(n16697), .ZN(n19526) );
  AOI22_X1 U12508 ( .A1(\mem[822][4] ), .A2(n16693), .B1(n26308), .B2(
        data_in[4]), .ZN(n16697) );
  INV_X1 U12509 ( .A(n16698), .ZN(n19525) );
  AOI22_X1 U12510 ( .A1(\mem[822][5] ), .A2(n16693), .B1(n26308), .B2(
        data_in[5]), .ZN(n16698) );
  INV_X1 U12511 ( .A(n16699), .ZN(n19524) );
  AOI22_X1 U12512 ( .A1(\mem[822][6] ), .A2(n16693), .B1(n26308), .B2(
        data_in[6]), .ZN(n16699) );
  INV_X1 U12513 ( .A(n16700), .ZN(n19523) );
  AOI22_X1 U12514 ( .A1(\mem[822][7] ), .A2(n16693), .B1(n26308), .B2(
        data_in[7]), .ZN(n16700) );
  INV_X1 U12515 ( .A(n16701), .ZN(n19522) );
  AOI22_X1 U12516 ( .A1(\mem[823][0] ), .A2(n16702), .B1(n26307), .B2(
        data_in[0]), .ZN(n16701) );
  INV_X1 U12517 ( .A(n16703), .ZN(n19521) );
  AOI22_X1 U12518 ( .A1(\mem[823][1] ), .A2(n16702), .B1(n26307), .B2(
        data_in[1]), .ZN(n16703) );
  INV_X1 U12519 ( .A(n16704), .ZN(n19520) );
  AOI22_X1 U12520 ( .A1(\mem[823][2] ), .A2(n16702), .B1(n26307), .B2(
        data_in[2]), .ZN(n16704) );
  INV_X1 U12521 ( .A(n16705), .ZN(n19519) );
  AOI22_X1 U12522 ( .A1(\mem[823][3] ), .A2(n16702), .B1(n26307), .B2(
        data_in[3]), .ZN(n16705) );
  INV_X1 U12523 ( .A(n16706), .ZN(n19518) );
  AOI22_X1 U12524 ( .A1(\mem[823][4] ), .A2(n16702), .B1(n26307), .B2(
        data_in[4]), .ZN(n16706) );
  INV_X1 U12525 ( .A(n16707), .ZN(n19517) );
  AOI22_X1 U12526 ( .A1(\mem[823][5] ), .A2(n16702), .B1(n26307), .B2(
        data_in[5]), .ZN(n16707) );
  INV_X1 U12527 ( .A(n16708), .ZN(n19516) );
  AOI22_X1 U12528 ( .A1(\mem[823][6] ), .A2(n16702), .B1(n26307), .B2(
        data_in[6]), .ZN(n16708) );
  INV_X1 U12529 ( .A(n16709), .ZN(n19515) );
  AOI22_X1 U12530 ( .A1(\mem[823][7] ), .A2(n16702), .B1(n26307), .B2(
        data_in[7]), .ZN(n16709) );
  INV_X1 U12531 ( .A(n16710), .ZN(n19514) );
  AOI22_X1 U12532 ( .A1(\mem[824][0] ), .A2(n16711), .B1(n26306), .B2(
        data_in[0]), .ZN(n16710) );
  INV_X1 U12533 ( .A(n16712), .ZN(n19513) );
  AOI22_X1 U12534 ( .A1(\mem[824][1] ), .A2(n16711), .B1(n26306), .B2(
        data_in[1]), .ZN(n16712) );
  INV_X1 U12535 ( .A(n16713), .ZN(n19512) );
  AOI22_X1 U12536 ( .A1(\mem[824][2] ), .A2(n16711), .B1(n26306), .B2(
        data_in[2]), .ZN(n16713) );
  INV_X1 U12537 ( .A(n16714), .ZN(n19511) );
  AOI22_X1 U12538 ( .A1(\mem[824][3] ), .A2(n16711), .B1(n26306), .B2(
        data_in[3]), .ZN(n16714) );
  INV_X1 U12539 ( .A(n16715), .ZN(n19510) );
  AOI22_X1 U12540 ( .A1(\mem[824][4] ), .A2(n16711), .B1(n26306), .B2(
        data_in[4]), .ZN(n16715) );
  INV_X1 U12541 ( .A(n16716), .ZN(n19509) );
  AOI22_X1 U12542 ( .A1(\mem[824][5] ), .A2(n16711), .B1(n26306), .B2(
        data_in[5]), .ZN(n16716) );
  INV_X1 U12543 ( .A(n16717), .ZN(n19508) );
  AOI22_X1 U12544 ( .A1(\mem[824][6] ), .A2(n16711), .B1(n26306), .B2(
        data_in[6]), .ZN(n16717) );
  INV_X1 U12545 ( .A(n16718), .ZN(n19507) );
  AOI22_X1 U12546 ( .A1(\mem[824][7] ), .A2(n16711), .B1(n26306), .B2(
        data_in[7]), .ZN(n16718) );
  INV_X1 U12547 ( .A(n16719), .ZN(n19506) );
  AOI22_X1 U12548 ( .A1(\mem[825][0] ), .A2(n16720), .B1(n26305), .B2(
        data_in[0]), .ZN(n16719) );
  INV_X1 U12549 ( .A(n16721), .ZN(n19505) );
  AOI22_X1 U12550 ( .A1(\mem[825][1] ), .A2(n16720), .B1(n26305), .B2(
        data_in[1]), .ZN(n16721) );
  INV_X1 U12551 ( .A(n16722), .ZN(n19504) );
  AOI22_X1 U12552 ( .A1(\mem[825][2] ), .A2(n16720), .B1(n26305), .B2(
        data_in[2]), .ZN(n16722) );
  INV_X1 U12553 ( .A(n16723), .ZN(n19503) );
  AOI22_X1 U12554 ( .A1(\mem[825][3] ), .A2(n16720), .B1(n26305), .B2(
        data_in[3]), .ZN(n16723) );
  INV_X1 U12555 ( .A(n16724), .ZN(n19502) );
  AOI22_X1 U12556 ( .A1(\mem[825][4] ), .A2(n16720), .B1(n26305), .B2(
        data_in[4]), .ZN(n16724) );
  INV_X1 U12557 ( .A(n16725), .ZN(n19501) );
  AOI22_X1 U12558 ( .A1(\mem[825][5] ), .A2(n16720), .B1(n26305), .B2(
        data_in[5]), .ZN(n16725) );
  INV_X1 U12559 ( .A(n16726), .ZN(n19500) );
  AOI22_X1 U12560 ( .A1(\mem[825][6] ), .A2(n16720), .B1(n26305), .B2(
        data_in[6]), .ZN(n16726) );
  INV_X1 U12561 ( .A(n16727), .ZN(n19499) );
  AOI22_X1 U12562 ( .A1(\mem[825][7] ), .A2(n16720), .B1(n26305), .B2(
        data_in[7]), .ZN(n16727) );
  INV_X1 U12563 ( .A(n16728), .ZN(n19498) );
  AOI22_X1 U12564 ( .A1(\mem[826][0] ), .A2(n16729), .B1(n26304), .B2(
        data_in[0]), .ZN(n16728) );
  INV_X1 U12565 ( .A(n16730), .ZN(n19497) );
  AOI22_X1 U12566 ( .A1(\mem[826][1] ), .A2(n16729), .B1(n26304), .B2(
        data_in[1]), .ZN(n16730) );
  INV_X1 U12567 ( .A(n16731), .ZN(n19496) );
  AOI22_X1 U12568 ( .A1(\mem[826][2] ), .A2(n16729), .B1(n26304), .B2(
        data_in[2]), .ZN(n16731) );
  INV_X1 U12569 ( .A(n16732), .ZN(n19495) );
  AOI22_X1 U12570 ( .A1(\mem[826][3] ), .A2(n16729), .B1(n26304), .B2(
        data_in[3]), .ZN(n16732) );
  INV_X1 U12571 ( .A(n16733), .ZN(n19494) );
  AOI22_X1 U12572 ( .A1(\mem[826][4] ), .A2(n16729), .B1(n26304), .B2(
        data_in[4]), .ZN(n16733) );
  INV_X1 U12573 ( .A(n16734), .ZN(n19493) );
  AOI22_X1 U12574 ( .A1(\mem[826][5] ), .A2(n16729), .B1(n26304), .B2(
        data_in[5]), .ZN(n16734) );
  INV_X1 U12575 ( .A(n16735), .ZN(n19492) );
  AOI22_X1 U12576 ( .A1(\mem[826][6] ), .A2(n16729), .B1(n26304), .B2(
        data_in[6]), .ZN(n16735) );
  INV_X1 U12577 ( .A(n16736), .ZN(n19491) );
  AOI22_X1 U12578 ( .A1(\mem[826][7] ), .A2(n16729), .B1(n26304), .B2(
        data_in[7]), .ZN(n16736) );
  INV_X1 U12579 ( .A(n16737), .ZN(n19490) );
  AOI22_X1 U12580 ( .A1(\mem[827][0] ), .A2(n16738), .B1(n26303), .B2(
        data_in[0]), .ZN(n16737) );
  INV_X1 U12581 ( .A(n16739), .ZN(n19489) );
  AOI22_X1 U12582 ( .A1(\mem[827][1] ), .A2(n16738), .B1(n26303), .B2(
        data_in[1]), .ZN(n16739) );
  INV_X1 U12583 ( .A(n16740), .ZN(n19488) );
  AOI22_X1 U12584 ( .A1(\mem[827][2] ), .A2(n16738), .B1(n26303), .B2(
        data_in[2]), .ZN(n16740) );
  INV_X1 U12585 ( .A(n16741), .ZN(n19487) );
  AOI22_X1 U12586 ( .A1(\mem[827][3] ), .A2(n16738), .B1(n26303), .B2(
        data_in[3]), .ZN(n16741) );
  INV_X1 U12587 ( .A(n16742), .ZN(n19486) );
  AOI22_X1 U12588 ( .A1(\mem[827][4] ), .A2(n16738), .B1(n26303), .B2(
        data_in[4]), .ZN(n16742) );
  INV_X1 U12589 ( .A(n16743), .ZN(n19485) );
  AOI22_X1 U12590 ( .A1(\mem[827][5] ), .A2(n16738), .B1(n26303), .B2(
        data_in[5]), .ZN(n16743) );
  INV_X1 U12591 ( .A(n16744), .ZN(n19484) );
  AOI22_X1 U12592 ( .A1(\mem[827][6] ), .A2(n16738), .B1(n26303), .B2(
        data_in[6]), .ZN(n16744) );
  INV_X1 U12593 ( .A(n16745), .ZN(n19483) );
  AOI22_X1 U12594 ( .A1(\mem[827][7] ), .A2(n16738), .B1(n26303), .B2(
        data_in[7]), .ZN(n16745) );
  INV_X1 U12595 ( .A(n16746), .ZN(n19482) );
  AOI22_X1 U12596 ( .A1(\mem[828][0] ), .A2(n16747), .B1(n26302), .B2(
        data_in[0]), .ZN(n16746) );
  INV_X1 U12597 ( .A(n16748), .ZN(n19481) );
  AOI22_X1 U12598 ( .A1(\mem[828][1] ), .A2(n16747), .B1(n26302), .B2(
        data_in[1]), .ZN(n16748) );
  INV_X1 U12599 ( .A(n16749), .ZN(n19480) );
  AOI22_X1 U12600 ( .A1(\mem[828][2] ), .A2(n16747), .B1(n26302), .B2(
        data_in[2]), .ZN(n16749) );
  INV_X1 U12601 ( .A(n16750), .ZN(n19479) );
  AOI22_X1 U12602 ( .A1(\mem[828][3] ), .A2(n16747), .B1(n26302), .B2(
        data_in[3]), .ZN(n16750) );
  INV_X1 U12603 ( .A(n16751), .ZN(n19478) );
  AOI22_X1 U12604 ( .A1(\mem[828][4] ), .A2(n16747), .B1(n26302), .B2(
        data_in[4]), .ZN(n16751) );
  INV_X1 U12605 ( .A(n16752), .ZN(n19477) );
  AOI22_X1 U12606 ( .A1(\mem[828][5] ), .A2(n16747), .B1(n26302), .B2(
        data_in[5]), .ZN(n16752) );
  INV_X1 U12607 ( .A(n16753), .ZN(n19476) );
  AOI22_X1 U12608 ( .A1(\mem[828][6] ), .A2(n16747), .B1(n26302), .B2(
        data_in[6]), .ZN(n16753) );
  INV_X1 U12609 ( .A(n16754), .ZN(n19475) );
  AOI22_X1 U12610 ( .A1(\mem[828][7] ), .A2(n16747), .B1(n26302), .B2(
        data_in[7]), .ZN(n16754) );
  INV_X1 U12611 ( .A(n16755), .ZN(n19474) );
  AOI22_X1 U12612 ( .A1(\mem[829][0] ), .A2(n16756), .B1(n26301), .B2(
        data_in[0]), .ZN(n16755) );
  INV_X1 U12613 ( .A(n16757), .ZN(n19473) );
  AOI22_X1 U12614 ( .A1(\mem[829][1] ), .A2(n16756), .B1(n26301), .B2(
        data_in[1]), .ZN(n16757) );
  INV_X1 U12615 ( .A(n16758), .ZN(n19472) );
  AOI22_X1 U12616 ( .A1(\mem[829][2] ), .A2(n16756), .B1(n26301), .B2(
        data_in[2]), .ZN(n16758) );
  INV_X1 U12617 ( .A(n16759), .ZN(n19471) );
  AOI22_X1 U12618 ( .A1(\mem[829][3] ), .A2(n16756), .B1(n26301), .B2(
        data_in[3]), .ZN(n16759) );
  INV_X1 U12619 ( .A(n16760), .ZN(n19470) );
  AOI22_X1 U12620 ( .A1(\mem[829][4] ), .A2(n16756), .B1(n26301), .B2(
        data_in[4]), .ZN(n16760) );
  INV_X1 U12621 ( .A(n16761), .ZN(n19469) );
  AOI22_X1 U12622 ( .A1(\mem[829][5] ), .A2(n16756), .B1(n26301), .B2(
        data_in[5]), .ZN(n16761) );
  INV_X1 U12623 ( .A(n16762), .ZN(n19468) );
  AOI22_X1 U12624 ( .A1(\mem[829][6] ), .A2(n16756), .B1(n26301), .B2(
        data_in[6]), .ZN(n16762) );
  INV_X1 U12625 ( .A(n16763), .ZN(n19467) );
  AOI22_X1 U12626 ( .A1(\mem[829][7] ), .A2(n16756), .B1(n26301), .B2(
        data_in[7]), .ZN(n16763) );
  INV_X1 U12627 ( .A(n16764), .ZN(n19466) );
  AOI22_X1 U12628 ( .A1(\mem[830][0] ), .A2(n16765), .B1(n26300), .B2(
        data_in[0]), .ZN(n16764) );
  INV_X1 U12629 ( .A(n16766), .ZN(n19465) );
  AOI22_X1 U12630 ( .A1(\mem[830][1] ), .A2(n16765), .B1(n26300), .B2(
        data_in[1]), .ZN(n16766) );
  INV_X1 U12631 ( .A(n16767), .ZN(n19464) );
  AOI22_X1 U12632 ( .A1(\mem[830][2] ), .A2(n16765), .B1(n26300), .B2(
        data_in[2]), .ZN(n16767) );
  INV_X1 U12633 ( .A(n16768), .ZN(n19463) );
  AOI22_X1 U12634 ( .A1(\mem[830][3] ), .A2(n16765), .B1(n26300), .B2(
        data_in[3]), .ZN(n16768) );
  INV_X1 U12635 ( .A(n16769), .ZN(n19462) );
  AOI22_X1 U12636 ( .A1(\mem[830][4] ), .A2(n16765), .B1(n26300), .B2(
        data_in[4]), .ZN(n16769) );
  INV_X1 U12637 ( .A(n16770), .ZN(n19461) );
  AOI22_X1 U12638 ( .A1(\mem[830][5] ), .A2(n16765), .B1(n26300), .B2(
        data_in[5]), .ZN(n16770) );
  INV_X1 U12639 ( .A(n16771), .ZN(n19460) );
  AOI22_X1 U12640 ( .A1(\mem[830][6] ), .A2(n16765), .B1(n26300), .B2(
        data_in[6]), .ZN(n16771) );
  INV_X1 U12641 ( .A(n16772), .ZN(n19459) );
  AOI22_X1 U12642 ( .A1(\mem[830][7] ), .A2(n16765), .B1(n26300), .B2(
        data_in[7]), .ZN(n16772) );
  INV_X1 U12643 ( .A(n16773), .ZN(n19458) );
  AOI22_X1 U12644 ( .A1(\mem[831][0] ), .A2(n16774), .B1(n26299), .B2(
        data_in[0]), .ZN(n16773) );
  INV_X1 U12645 ( .A(n16775), .ZN(n19457) );
  AOI22_X1 U12646 ( .A1(\mem[831][1] ), .A2(n16774), .B1(n26299), .B2(
        data_in[1]), .ZN(n16775) );
  INV_X1 U12647 ( .A(n16776), .ZN(n19456) );
  AOI22_X1 U12648 ( .A1(\mem[831][2] ), .A2(n16774), .B1(n26299), .B2(
        data_in[2]), .ZN(n16776) );
  INV_X1 U12649 ( .A(n16777), .ZN(n19455) );
  AOI22_X1 U12650 ( .A1(\mem[831][3] ), .A2(n16774), .B1(n26299), .B2(
        data_in[3]), .ZN(n16777) );
  INV_X1 U12651 ( .A(n16778), .ZN(n19454) );
  AOI22_X1 U12652 ( .A1(\mem[831][4] ), .A2(n16774), .B1(n26299), .B2(
        data_in[4]), .ZN(n16778) );
  INV_X1 U12653 ( .A(n16779), .ZN(n19453) );
  AOI22_X1 U12654 ( .A1(\mem[831][5] ), .A2(n16774), .B1(n26299), .B2(
        data_in[5]), .ZN(n16779) );
  INV_X1 U12655 ( .A(n16780), .ZN(n19452) );
  AOI22_X1 U12656 ( .A1(\mem[831][6] ), .A2(n16774), .B1(n26299), .B2(
        data_in[6]), .ZN(n16780) );
  INV_X1 U12657 ( .A(n16781), .ZN(n19451) );
  AOI22_X1 U12658 ( .A1(\mem[831][7] ), .A2(n16774), .B1(n26299), .B2(
        data_in[7]), .ZN(n16781) );
  INV_X1 U12659 ( .A(n16855), .ZN(n19386) );
  AOI22_X1 U12660 ( .A1(\mem[840][0] ), .A2(n16856), .B1(n26290), .B2(
        data_in[0]), .ZN(n16855) );
  INV_X1 U12661 ( .A(n16857), .ZN(n19385) );
  AOI22_X1 U12662 ( .A1(\mem[840][1] ), .A2(n16856), .B1(n26290), .B2(
        data_in[1]), .ZN(n16857) );
  INV_X1 U12663 ( .A(n16858), .ZN(n19384) );
  AOI22_X1 U12664 ( .A1(\mem[840][2] ), .A2(n16856), .B1(n26290), .B2(
        data_in[2]), .ZN(n16858) );
  INV_X1 U12665 ( .A(n16859), .ZN(n19383) );
  AOI22_X1 U12666 ( .A1(\mem[840][3] ), .A2(n16856), .B1(n26290), .B2(
        data_in[3]), .ZN(n16859) );
  INV_X1 U12667 ( .A(n16860), .ZN(n19382) );
  AOI22_X1 U12668 ( .A1(\mem[840][4] ), .A2(n16856), .B1(n26290), .B2(
        data_in[4]), .ZN(n16860) );
  INV_X1 U12669 ( .A(n16861), .ZN(n19381) );
  AOI22_X1 U12670 ( .A1(\mem[840][5] ), .A2(n16856), .B1(n26290), .B2(
        data_in[5]), .ZN(n16861) );
  INV_X1 U12671 ( .A(n16862), .ZN(n19380) );
  AOI22_X1 U12672 ( .A1(\mem[840][6] ), .A2(n16856), .B1(n26290), .B2(
        data_in[6]), .ZN(n16862) );
  INV_X1 U12673 ( .A(n16863), .ZN(n19379) );
  AOI22_X1 U12674 ( .A1(\mem[840][7] ), .A2(n16856), .B1(n26290), .B2(
        data_in[7]), .ZN(n16863) );
  INV_X1 U12675 ( .A(n16864), .ZN(n19378) );
  AOI22_X1 U12676 ( .A1(\mem[841][0] ), .A2(n16865), .B1(n26289), .B2(
        data_in[0]), .ZN(n16864) );
  INV_X1 U12677 ( .A(n16866), .ZN(n19377) );
  AOI22_X1 U12678 ( .A1(\mem[841][1] ), .A2(n16865), .B1(n26289), .B2(
        data_in[1]), .ZN(n16866) );
  INV_X1 U12679 ( .A(n16867), .ZN(n19376) );
  AOI22_X1 U12680 ( .A1(\mem[841][2] ), .A2(n16865), .B1(n26289), .B2(
        data_in[2]), .ZN(n16867) );
  INV_X1 U12681 ( .A(n16868), .ZN(n19375) );
  AOI22_X1 U12682 ( .A1(\mem[841][3] ), .A2(n16865), .B1(n26289), .B2(
        data_in[3]), .ZN(n16868) );
  INV_X1 U12683 ( .A(n16869), .ZN(n19374) );
  AOI22_X1 U12684 ( .A1(\mem[841][4] ), .A2(n16865), .B1(n26289), .B2(
        data_in[4]), .ZN(n16869) );
  INV_X1 U12685 ( .A(n16870), .ZN(n19373) );
  AOI22_X1 U12686 ( .A1(\mem[841][5] ), .A2(n16865), .B1(n26289), .B2(
        data_in[5]), .ZN(n16870) );
  INV_X1 U12687 ( .A(n16871), .ZN(n19372) );
  AOI22_X1 U12688 ( .A1(\mem[841][6] ), .A2(n16865), .B1(n26289), .B2(
        data_in[6]), .ZN(n16871) );
  INV_X1 U12689 ( .A(n16872), .ZN(n19371) );
  AOI22_X1 U12690 ( .A1(\mem[841][7] ), .A2(n16865), .B1(n26289), .B2(
        data_in[7]), .ZN(n16872) );
  INV_X1 U12691 ( .A(n16873), .ZN(n19370) );
  AOI22_X1 U12692 ( .A1(\mem[842][0] ), .A2(n16874), .B1(n26288), .B2(
        data_in[0]), .ZN(n16873) );
  INV_X1 U12693 ( .A(n16875), .ZN(n19369) );
  AOI22_X1 U12694 ( .A1(\mem[842][1] ), .A2(n16874), .B1(n26288), .B2(
        data_in[1]), .ZN(n16875) );
  INV_X1 U12695 ( .A(n16876), .ZN(n19368) );
  AOI22_X1 U12696 ( .A1(\mem[842][2] ), .A2(n16874), .B1(n26288), .B2(
        data_in[2]), .ZN(n16876) );
  INV_X1 U12697 ( .A(n16877), .ZN(n19367) );
  AOI22_X1 U12698 ( .A1(\mem[842][3] ), .A2(n16874), .B1(n26288), .B2(
        data_in[3]), .ZN(n16877) );
  INV_X1 U12699 ( .A(n16878), .ZN(n19366) );
  AOI22_X1 U12700 ( .A1(\mem[842][4] ), .A2(n16874), .B1(n26288), .B2(
        data_in[4]), .ZN(n16878) );
  INV_X1 U12701 ( .A(n16879), .ZN(n19365) );
  AOI22_X1 U12702 ( .A1(\mem[842][5] ), .A2(n16874), .B1(n26288), .B2(
        data_in[5]), .ZN(n16879) );
  INV_X1 U12703 ( .A(n16880), .ZN(n19364) );
  AOI22_X1 U12704 ( .A1(\mem[842][6] ), .A2(n16874), .B1(n26288), .B2(
        data_in[6]), .ZN(n16880) );
  INV_X1 U12705 ( .A(n16881), .ZN(n19363) );
  AOI22_X1 U12706 ( .A1(\mem[842][7] ), .A2(n16874), .B1(n26288), .B2(
        data_in[7]), .ZN(n16881) );
  INV_X1 U12707 ( .A(n16882), .ZN(n19362) );
  AOI22_X1 U12708 ( .A1(\mem[843][0] ), .A2(n16883), .B1(n26287), .B2(
        data_in[0]), .ZN(n16882) );
  INV_X1 U12709 ( .A(n16884), .ZN(n19361) );
  AOI22_X1 U12710 ( .A1(\mem[843][1] ), .A2(n16883), .B1(n26287), .B2(
        data_in[1]), .ZN(n16884) );
  INV_X1 U12711 ( .A(n16885), .ZN(n19360) );
  AOI22_X1 U12712 ( .A1(\mem[843][2] ), .A2(n16883), .B1(n26287), .B2(
        data_in[2]), .ZN(n16885) );
  INV_X1 U12713 ( .A(n16886), .ZN(n19359) );
  AOI22_X1 U12714 ( .A1(\mem[843][3] ), .A2(n16883), .B1(n26287), .B2(
        data_in[3]), .ZN(n16886) );
  INV_X1 U12715 ( .A(n16887), .ZN(n19358) );
  AOI22_X1 U12716 ( .A1(\mem[843][4] ), .A2(n16883), .B1(n26287), .B2(
        data_in[4]), .ZN(n16887) );
  INV_X1 U12717 ( .A(n16888), .ZN(n19357) );
  AOI22_X1 U12718 ( .A1(\mem[843][5] ), .A2(n16883), .B1(n26287), .B2(
        data_in[5]), .ZN(n16888) );
  INV_X1 U12719 ( .A(n16889), .ZN(n19356) );
  AOI22_X1 U12720 ( .A1(\mem[843][6] ), .A2(n16883), .B1(n26287), .B2(
        data_in[6]), .ZN(n16889) );
  INV_X1 U12721 ( .A(n16890), .ZN(n19355) );
  AOI22_X1 U12722 ( .A1(\mem[843][7] ), .A2(n16883), .B1(n26287), .B2(
        data_in[7]), .ZN(n16890) );
  INV_X1 U12723 ( .A(n16891), .ZN(n19354) );
  AOI22_X1 U12724 ( .A1(\mem[844][0] ), .A2(n16892), .B1(n26286), .B2(
        data_in[0]), .ZN(n16891) );
  INV_X1 U12725 ( .A(n16893), .ZN(n19353) );
  AOI22_X1 U12726 ( .A1(\mem[844][1] ), .A2(n16892), .B1(n26286), .B2(
        data_in[1]), .ZN(n16893) );
  INV_X1 U12727 ( .A(n16894), .ZN(n19352) );
  AOI22_X1 U12728 ( .A1(\mem[844][2] ), .A2(n16892), .B1(n26286), .B2(
        data_in[2]), .ZN(n16894) );
  INV_X1 U12729 ( .A(n16895), .ZN(n19351) );
  AOI22_X1 U12730 ( .A1(\mem[844][3] ), .A2(n16892), .B1(n26286), .B2(
        data_in[3]), .ZN(n16895) );
  INV_X1 U12731 ( .A(n16896), .ZN(n19350) );
  AOI22_X1 U12732 ( .A1(\mem[844][4] ), .A2(n16892), .B1(n26286), .B2(
        data_in[4]), .ZN(n16896) );
  INV_X1 U12733 ( .A(n16897), .ZN(n19349) );
  AOI22_X1 U12734 ( .A1(\mem[844][5] ), .A2(n16892), .B1(n26286), .B2(
        data_in[5]), .ZN(n16897) );
  INV_X1 U12735 ( .A(n16898), .ZN(n19348) );
  AOI22_X1 U12736 ( .A1(\mem[844][6] ), .A2(n16892), .B1(n26286), .B2(
        data_in[6]), .ZN(n16898) );
  INV_X1 U12737 ( .A(n16899), .ZN(n19347) );
  AOI22_X1 U12738 ( .A1(\mem[844][7] ), .A2(n16892), .B1(n26286), .B2(
        data_in[7]), .ZN(n16899) );
  INV_X1 U12739 ( .A(n16900), .ZN(n19346) );
  AOI22_X1 U12740 ( .A1(\mem[845][0] ), .A2(n16901), .B1(n26285), .B2(
        data_in[0]), .ZN(n16900) );
  INV_X1 U12741 ( .A(n16902), .ZN(n19345) );
  AOI22_X1 U12742 ( .A1(\mem[845][1] ), .A2(n16901), .B1(n26285), .B2(
        data_in[1]), .ZN(n16902) );
  INV_X1 U12743 ( .A(n16903), .ZN(n19344) );
  AOI22_X1 U12744 ( .A1(\mem[845][2] ), .A2(n16901), .B1(n26285), .B2(
        data_in[2]), .ZN(n16903) );
  INV_X1 U12745 ( .A(n16904), .ZN(n19343) );
  AOI22_X1 U12746 ( .A1(\mem[845][3] ), .A2(n16901), .B1(n26285), .B2(
        data_in[3]), .ZN(n16904) );
  INV_X1 U12747 ( .A(n16905), .ZN(n19342) );
  AOI22_X1 U12748 ( .A1(\mem[845][4] ), .A2(n16901), .B1(n26285), .B2(
        data_in[4]), .ZN(n16905) );
  INV_X1 U12749 ( .A(n16906), .ZN(n19341) );
  AOI22_X1 U12750 ( .A1(\mem[845][5] ), .A2(n16901), .B1(n26285), .B2(
        data_in[5]), .ZN(n16906) );
  INV_X1 U12751 ( .A(n16907), .ZN(n19340) );
  AOI22_X1 U12752 ( .A1(\mem[845][6] ), .A2(n16901), .B1(n26285), .B2(
        data_in[6]), .ZN(n16907) );
  INV_X1 U12753 ( .A(n16908), .ZN(n19339) );
  AOI22_X1 U12754 ( .A1(\mem[845][7] ), .A2(n16901), .B1(n26285), .B2(
        data_in[7]), .ZN(n16908) );
  INV_X1 U12755 ( .A(n16909), .ZN(n19338) );
  AOI22_X1 U12756 ( .A1(\mem[846][0] ), .A2(n16910), .B1(n26284), .B2(
        data_in[0]), .ZN(n16909) );
  INV_X1 U12757 ( .A(n16911), .ZN(n19337) );
  AOI22_X1 U12758 ( .A1(\mem[846][1] ), .A2(n16910), .B1(n26284), .B2(
        data_in[1]), .ZN(n16911) );
  INV_X1 U12759 ( .A(n16912), .ZN(n19336) );
  AOI22_X1 U12760 ( .A1(\mem[846][2] ), .A2(n16910), .B1(n26284), .B2(
        data_in[2]), .ZN(n16912) );
  INV_X1 U12761 ( .A(n16913), .ZN(n19335) );
  AOI22_X1 U12762 ( .A1(\mem[846][3] ), .A2(n16910), .B1(n26284), .B2(
        data_in[3]), .ZN(n16913) );
  INV_X1 U12763 ( .A(n16914), .ZN(n19334) );
  AOI22_X1 U12764 ( .A1(\mem[846][4] ), .A2(n16910), .B1(n26284), .B2(
        data_in[4]), .ZN(n16914) );
  INV_X1 U12765 ( .A(n16915), .ZN(n19333) );
  AOI22_X1 U12766 ( .A1(\mem[846][5] ), .A2(n16910), .B1(n26284), .B2(
        data_in[5]), .ZN(n16915) );
  INV_X1 U12767 ( .A(n16916), .ZN(n19332) );
  AOI22_X1 U12768 ( .A1(\mem[846][6] ), .A2(n16910), .B1(n26284), .B2(
        data_in[6]), .ZN(n16916) );
  INV_X1 U12769 ( .A(n16917), .ZN(n19331) );
  AOI22_X1 U12770 ( .A1(\mem[846][7] ), .A2(n16910), .B1(n26284), .B2(
        data_in[7]), .ZN(n16917) );
  INV_X1 U12771 ( .A(n16918), .ZN(n19330) );
  AOI22_X1 U12772 ( .A1(\mem[847][0] ), .A2(n16919), .B1(n26283), .B2(
        data_in[0]), .ZN(n16918) );
  INV_X1 U12773 ( .A(n16920), .ZN(n19329) );
  AOI22_X1 U12774 ( .A1(\mem[847][1] ), .A2(n16919), .B1(n26283), .B2(
        data_in[1]), .ZN(n16920) );
  INV_X1 U12775 ( .A(n16921), .ZN(n19328) );
  AOI22_X1 U12776 ( .A1(\mem[847][2] ), .A2(n16919), .B1(n26283), .B2(
        data_in[2]), .ZN(n16921) );
  INV_X1 U12777 ( .A(n16922), .ZN(n19327) );
  AOI22_X1 U12778 ( .A1(\mem[847][3] ), .A2(n16919), .B1(n26283), .B2(
        data_in[3]), .ZN(n16922) );
  INV_X1 U12779 ( .A(n16923), .ZN(n19326) );
  AOI22_X1 U12780 ( .A1(\mem[847][4] ), .A2(n16919), .B1(n26283), .B2(
        data_in[4]), .ZN(n16923) );
  INV_X1 U12781 ( .A(n16924), .ZN(n19325) );
  AOI22_X1 U12782 ( .A1(\mem[847][5] ), .A2(n16919), .B1(n26283), .B2(
        data_in[5]), .ZN(n16924) );
  INV_X1 U12783 ( .A(n16925), .ZN(n19324) );
  AOI22_X1 U12784 ( .A1(\mem[847][6] ), .A2(n16919), .B1(n26283), .B2(
        data_in[6]), .ZN(n16925) );
  INV_X1 U12785 ( .A(n16926), .ZN(n19323) );
  AOI22_X1 U12786 ( .A1(\mem[847][7] ), .A2(n16919), .B1(n26283), .B2(
        data_in[7]), .ZN(n16926) );
  INV_X1 U12787 ( .A(n16927), .ZN(n19322) );
  AOI22_X1 U12788 ( .A1(\mem[848][0] ), .A2(n16928), .B1(n26282), .B2(
        data_in[0]), .ZN(n16927) );
  INV_X1 U12789 ( .A(n16929), .ZN(n19321) );
  AOI22_X1 U12790 ( .A1(\mem[848][1] ), .A2(n16928), .B1(n26282), .B2(
        data_in[1]), .ZN(n16929) );
  INV_X1 U12791 ( .A(n16930), .ZN(n19320) );
  AOI22_X1 U12792 ( .A1(\mem[848][2] ), .A2(n16928), .B1(n26282), .B2(
        data_in[2]), .ZN(n16930) );
  INV_X1 U12793 ( .A(n16931), .ZN(n19319) );
  AOI22_X1 U12794 ( .A1(\mem[848][3] ), .A2(n16928), .B1(n26282), .B2(
        data_in[3]), .ZN(n16931) );
  INV_X1 U12795 ( .A(n16932), .ZN(n19318) );
  AOI22_X1 U12796 ( .A1(\mem[848][4] ), .A2(n16928), .B1(n26282), .B2(
        data_in[4]), .ZN(n16932) );
  INV_X1 U12797 ( .A(n16933), .ZN(n19317) );
  AOI22_X1 U12798 ( .A1(\mem[848][5] ), .A2(n16928), .B1(n26282), .B2(
        data_in[5]), .ZN(n16933) );
  INV_X1 U12799 ( .A(n16934), .ZN(n19316) );
  AOI22_X1 U12800 ( .A1(\mem[848][6] ), .A2(n16928), .B1(n26282), .B2(
        data_in[6]), .ZN(n16934) );
  INV_X1 U12801 ( .A(n16935), .ZN(n19315) );
  AOI22_X1 U12802 ( .A1(\mem[848][7] ), .A2(n16928), .B1(n26282), .B2(
        data_in[7]), .ZN(n16935) );
  INV_X1 U12803 ( .A(n16936), .ZN(n19314) );
  AOI22_X1 U12804 ( .A1(\mem[849][0] ), .A2(n16937), .B1(n26281), .B2(
        data_in[0]), .ZN(n16936) );
  INV_X1 U12805 ( .A(n16938), .ZN(n19313) );
  AOI22_X1 U12806 ( .A1(\mem[849][1] ), .A2(n16937), .B1(n26281), .B2(
        data_in[1]), .ZN(n16938) );
  INV_X1 U12807 ( .A(n16939), .ZN(n19312) );
  AOI22_X1 U12808 ( .A1(\mem[849][2] ), .A2(n16937), .B1(n26281), .B2(
        data_in[2]), .ZN(n16939) );
  INV_X1 U12809 ( .A(n16940), .ZN(n19311) );
  AOI22_X1 U12810 ( .A1(\mem[849][3] ), .A2(n16937), .B1(n26281), .B2(
        data_in[3]), .ZN(n16940) );
  INV_X1 U12811 ( .A(n16941), .ZN(n19310) );
  AOI22_X1 U12812 ( .A1(\mem[849][4] ), .A2(n16937), .B1(n26281), .B2(
        data_in[4]), .ZN(n16941) );
  INV_X1 U12813 ( .A(n16942), .ZN(n19309) );
  AOI22_X1 U12814 ( .A1(\mem[849][5] ), .A2(n16937), .B1(n26281), .B2(
        data_in[5]), .ZN(n16942) );
  INV_X1 U12815 ( .A(n16943), .ZN(n19308) );
  AOI22_X1 U12816 ( .A1(\mem[849][6] ), .A2(n16937), .B1(n26281), .B2(
        data_in[6]), .ZN(n16943) );
  INV_X1 U12817 ( .A(n16944), .ZN(n19307) );
  AOI22_X1 U12818 ( .A1(\mem[849][7] ), .A2(n16937), .B1(n26281), .B2(
        data_in[7]), .ZN(n16944) );
  INV_X1 U12819 ( .A(n16945), .ZN(n19306) );
  AOI22_X1 U12820 ( .A1(\mem[850][0] ), .A2(n16946), .B1(n26280), .B2(
        data_in[0]), .ZN(n16945) );
  INV_X1 U12821 ( .A(n16947), .ZN(n19305) );
  AOI22_X1 U12822 ( .A1(\mem[850][1] ), .A2(n16946), .B1(n26280), .B2(
        data_in[1]), .ZN(n16947) );
  INV_X1 U12823 ( .A(n16948), .ZN(n19304) );
  AOI22_X1 U12824 ( .A1(\mem[850][2] ), .A2(n16946), .B1(n26280), .B2(
        data_in[2]), .ZN(n16948) );
  INV_X1 U12825 ( .A(n16949), .ZN(n19303) );
  AOI22_X1 U12826 ( .A1(\mem[850][3] ), .A2(n16946), .B1(n26280), .B2(
        data_in[3]), .ZN(n16949) );
  INV_X1 U12827 ( .A(n16950), .ZN(n19302) );
  AOI22_X1 U12828 ( .A1(\mem[850][4] ), .A2(n16946), .B1(n26280), .B2(
        data_in[4]), .ZN(n16950) );
  INV_X1 U12829 ( .A(n16951), .ZN(n19301) );
  AOI22_X1 U12830 ( .A1(\mem[850][5] ), .A2(n16946), .B1(n26280), .B2(
        data_in[5]), .ZN(n16951) );
  INV_X1 U12831 ( .A(n16952), .ZN(n19300) );
  AOI22_X1 U12832 ( .A1(\mem[850][6] ), .A2(n16946), .B1(n26280), .B2(
        data_in[6]), .ZN(n16952) );
  INV_X1 U12833 ( .A(n16953), .ZN(n19299) );
  AOI22_X1 U12834 ( .A1(\mem[850][7] ), .A2(n16946), .B1(n26280), .B2(
        data_in[7]), .ZN(n16953) );
  INV_X1 U12835 ( .A(n16954), .ZN(n19298) );
  AOI22_X1 U12836 ( .A1(\mem[851][0] ), .A2(n16955), .B1(n26279), .B2(
        data_in[0]), .ZN(n16954) );
  INV_X1 U12837 ( .A(n16956), .ZN(n19297) );
  AOI22_X1 U12838 ( .A1(\mem[851][1] ), .A2(n16955), .B1(n26279), .B2(
        data_in[1]), .ZN(n16956) );
  INV_X1 U12839 ( .A(n16957), .ZN(n19296) );
  AOI22_X1 U12840 ( .A1(\mem[851][2] ), .A2(n16955), .B1(n26279), .B2(
        data_in[2]), .ZN(n16957) );
  INV_X1 U12841 ( .A(n16958), .ZN(n19295) );
  AOI22_X1 U12842 ( .A1(\mem[851][3] ), .A2(n16955), .B1(n26279), .B2(
        data_in[3]), .ZN(n16958) );
  INV_X1 U12843 ( .A(n16959), .ZN(n19294) );
  AOI22_X1 U12844 ( .A1(\mem[851][4] ), .A2(n16955), .B1(n26279), .B2(
        data_in[4]), .ZN(n16959) );
  INV_X1 U12845 ( .A(n16960), .ZN(n19293) );
  AOI22_X1 U12846 ( .A1(\mem[851][5] ), .A2(n16955), .B1(n26279), .B2(
        data_in[5]), .ZN(n16960) );
  INV_X1 U12847 ( .A(n16961), .ZN(n19292) );
  AOI22_X1 U12848 ( .A1(\mem[851][6] ), .A2(n16955), .B1(n26279), .B2(
        data_in[6]), .ZN(n16961) );
  INV_X1 U12849 ( .A(n16962), .ZN(n19291) );
  AOI22_X1 U12850 ( .A1(\mem[851][7] ), .A2(n16955), .B1(n26279), .B2(
        data_in[7]), .ZN(n16962) );
  INV_X1 U12851 ( .A(n16963), .ZN(n19290) );
  AOI22_X1 U12852 ( .A1(\mem[852][0] ), .A2(n16964), .B1(n26278), .B2(
        data_in[0]), .ZN(n16963) );
  INV_X1 U12853 ( .A(n16965), .ZN(n19289) );
  AOI22_X1 U12854 ( .A1(\mem[852][1] ), .A2(n16964), .B1(n26278), .B2(
        data_in[1]), .ZN(n16965) );
  INV_X1 U12855 ( .A(n16966), .ZN(n19288) );
  AOI22_X1 U12856 ( .A1(\mem[852][2] ), .A2(n16964), .B1(n26278), .B2(
        data_in[2]), .ZN(n16966) );
  INV_X1 U12857 ( .A(n16967), .ZN(n19287) );
  AOI22_X1 U12858 ( .A1(\mem[852][3] ), .A2(n16964), .B1(n26278), .B2(
        data_in[3]), .ZN(n16967) );
  INV_X1 U12859 ( .A(n16968), .ZN(n19286) );
  AOI22_X1 U12860 ( .A1(\mem[852][4] ), .A2(n16964), .B1(n26278), .B2(
        data_in[4]), .ZN(n16968) );
  INV_X1 U12861 ( .A(n16969), .ZN(n19285) );
  AOI22_X1 U12862 ( .A1(\mem[852][5] ), .A2(n16964), .B1(n26278), .B2(
        data_in[5]), .ZN(n16969) );
  INV_X1 U12863 ( .A(n16970), .ZN(n19284) );
  AOI22_X1 U12864 ( .A1(\mem[852][6] ), .A2(n16964), .B1(n26278), .B2(
        data_in[6]), .ZN(n16970) );
  INV_X1 U12865 ( .A(n16971), .ZN(n19283) );
  AOI22_X1 U12866 ( .A1(\mem[852][7] ), .A2(n16964), .B1(n26278), .B2(
        data_in[7]), .ZN(n16971) );
  INV_X1 U12867 ( .A(n16972), .ZN(n19282) );
  AOI22_X1 U12868 ( .A1(\mem[853][0] ), .A2(n16973), .B1(n26277), .B2(
        data_in[0]), .ZN(n16972) );
  INV_X1 U12869 ( .A(n16974), .ZN(n19281) );
  AOI22_X1 U12870 ( .A1(\mem[853][1] ), .A2(n16973), .B1(n26277), .B2(
        data_in[1]), .ZN(n16974) );
  INV_X1 U12871 ( .A(n16975), .ZN(n19280) );
  AOI22_X1 U12872 ( .A1(\mem[853][2] ), .A2(n16973), .B1(n26277), .B2(
        data_in[2]), .ZN(n16975) );
  INV_X1 U12873 ( .A(n16976), .ZN(n19279) );
  AOI22_X1 U12874 ( .A1(\mem[853][3] ), .A2(n16973), .B1(n26277), .B2(
        data_in[3]), .ZN(n16976) );
  INV_X1 U12875 ( .A(n16977), .ZN(n19278) );
  AOI22_X1 U12876 ( .A1(\mem[853][4] ), .A2(n16973), .B1(n26277), .B2(
        data_in[4]), .ZN(n16977) );
  INV_X1 U12877 ( .A(n16978), .ZN(n19277) );
  AOI22_X1 U12878 ( .A1(\mem[853][5] ), .A2(n16973), .B1(n26277), .B2(
        data_in[5]), .ZN(n16978) );
  INV_X1 U12879 ( .A(n16979), .ZN(n19276) );
  AOI22_X1 U12880 ( .A1(\mem[853][6] ), .A2(n16973), .B1(n26277), .B2(
        data_in[6]), .ZN(n16979) );
  INV_X1 U12881 ( .A(n16980), .ZN(n19275) );
  AOI22_X1 U12882 ( .A1(\mem[853][7] ), .A2(n16973), .B1(n26277), .B2(
        data_in[7]), .ZN(n16980) );
  INV_X1 U12883 ( .A(n16981), .ZN(n19274) );
  AOI22_X1 U12884 ( .A1(\mem[854][0] ), .A2(n16982), .B1(n26276), .B2(
        data_in[0]), .ZN(n16981) );
  INV_X1 U12885 ( .A(n16983), .ZN(n19273) );
  AOI22_X1 U12886 ( .A1(\mem[854][1] ), .A2(n16982), .B1(n26276), .B2(
        data_in[1]), .ZN(n16983) );
  INV_X1 U12887 ( .A(n16984), .ZN(n19272) );
  AOI22_X1 U12888 ( .A1(\mem[854][2] ), .A2(n16982), .B1(n26276), .B2(
        data_in[2]), .ZN(n16984) );
  INV_X1 U12889 ( .A(n16985), .ZN(n19271) );
  AOI22_X1 U12890 ( .A1(\mem[854][3] ), .A2(n16982), .B1(n26276), .B2(
        data_in[3]), .ZN(n16985) );
  INV_X1 U12891 ( .A(n16986), .ZN(n19270) );
  AOI22_X1 U12892 ( .A1(\mem[854][4] ), .A2(n16982), .B1(n26276), .B2(
        data_in[4]), .ZN(n16986) );
  INV_X1 U12893 ( .A(n16987), .ZN(n19269) );
  AOI22_X1 U12894 ( .A1(\mem[854][5] ), .A2(n16982), .B1(n26276), .B2(
        data_in[5]), .ZN(n16987) );
  INV_X1 U12895 ( .A(n16988), .ZN(n19268) );
  AOI22_X1 U12896 ( .A1(\mem[854][6] ), .A2(n16982), .B1(n26276), .B2(
        data_in[6]), .ZN(n16988) );
  INV_X1 U12897 ( .A(n16989), .ZN(n19267) );
  AOI22_X1 U12898 ( .A1(\mem[854][7] ), .A2(n16982), .B1(n26276), .B2(
        data_in[7]), .ZN(n16989) );
  INV_X1 U12899 ( .A(n16990), .ZN(n19266) );
  AOI22_X1 U12900 ( .A1(\mem[855][0] ), .A2(n16991), .B1(n26275), .B2(
        data_in[0]), .ZN(n16990) );
  INV_X1 U12901 ( .A(n16992), .ZN(n19265) );
  AOI22_X1 U12902 ( .A1(\mem[855][1] ), .A2(n16991), .B1(n26275), .B2(
        data_in[1]), .ZN(n16992) );
  INV_X1 U12903 ( .A(n16993), .ZN(n19264) );
  AOI22_X1 U12904 ( .A1(\mem[855][2] ), .A2(n16991), .B1(n26275), .B2(
        data_in[2]), .ZN(n16993) );
  INV_X1 U12905 ( .A(n16994), .ZN(n19263) );
  AOI22_X1 U12906 ( .A1(\mem[855][3] ), .A2(n16991), .B1(n26275), .B2(
        data_in[3]), .ZN(n16994) );
  INV_X1 U12907 ( .A(n16995), .ZN(n19262) );
  AOI22_X1 U12908 ( .A1(\mem[855][4] ), .A2(n16991), .B1(n26275), .B2(
        data_in[4]), .ZN(n16995) );
  INV_X1 U12909 ( .A(n16996), .ZN(n19261) );
  AOI22_X1 U12910 ( .A1(\mem[855][5] ), .A2(n16991), .B1(n26275), .B2(
        data_in[5]), .ZN(n16996) );
  INV_X1 U12911 ( .A(n16997), .ZN(n19260) );
  AOI22_X1 U12912 ( .A1(\mem[855][6] ), .A2(n16991), .B1(n26275), .B2(
        data_in[6]), .ZN(n16997) );
  INV_X1 U12913 ( .A(n16998), .ZN(n19259) );
  AOI22_X1 U12914 ( .A1(\mem[855][7] ), .A2(n16991), .B1(n26275), .B2(
        data_in[7]), .ZN(n16998) );
  INV_X1 U12915 ( .A(n16999), .ZN(n19258) );
  AOI22_X1 U12916 ( .A1(\mem[856][0] ), .A2(n17000), .B1(n26274), .B2(
        data_in[0]), .ZN(n16999) );
  INV_X1 U12917 ( .A(n17001), .ZN(n19257) );
  AOI22_X1 U12918 ( .A1(\mem[856][1] ), .A2(n17000), .B1(n26274), .B2(
        data_in[1]), .ZN(n17001) );
  INV_X1 U12919 ( .A(n17002), .ZN(n19256) );
  AOI22_X1 U12920 ( .A1(\mem[856][2] ), .A2(n17000), .B1(n26274), .B2(
        data_in[2]), .ZN(n17002) );
  INV_X1 U12921 ( .A(n17003), .ZN(n19255) );
  AOI22_X1 U12922 ( .A1(\mem[856][3] ), .A2(n17000), .B1(n26274), .B2(
        data_in[3]), .ZN(n17003) );
  INV_X1 U12923 ( .A(n17004), .ZN(n19254) );
  AOI22_X1 U12924 ( .A1(\mem[856][4] ), .A2(n17000), .B1(n26274), .B2(
        data_in[4]), .ZN(n17004) );
  INV_X1 U12925 ( .A(n17005), .ZN(n19253) );
  AOI22_X1 U12926 ( .A1(\mem[856][5] ), .A2(n17000), .B1(n26274), .B2(
        data_in[5]), .ZN(n17005) );
  INV_X1 U12927 ( .A(n17006), .ZN(n19252) );
  AOI22_X1 U12928 ( .A1(\mem[856][6] ), .A2(n17000), .B1(n26274), .B2(
        data_in[6]), .ZN(n17006) );
  INV_X1 U12929 ( .A(n17007), .ZN(n19251) );
  AOI22_X1 U12930 ( .A1(\mem[856][7] ), .A2(n17000), .B1(n26274), .B2(
        data_in[7]), .ZN(n17007) );
  INV_X1 U12931 ( .A(n17008), .ZN(n19250) );
  AOI22_X1 U12932 ( .A1(\mem[857][0] ), .A2(n17009), .B1(n26273), .B2(
        data_in[0]), .ZN(n17008) );
  INV_X1 U12933 ( .A(n17010), .ZN(n19249) );
  AOI22_X1 U12934 ( .A1(\mem[857][1] ), .A2(n17009), .B1(n26273), .B2(
        data_in[1]), .ZN(n17010) );
  INV_X1 U12935 ( .A(n17011), .ZN(n19248) );
  AOI22_X1 U12936 ( .A1(\mem[857][2] ), .A2(n17009), .B1(n26273), .B2(
        data_in[2]), .ZN(n17011) );
  INV_X1 U12937 ( .A(n17012), .ZN(n19247) );
  AOI22_X1 U12938 ( .A1(\mem[857][3] ), .A2(n17009), .B1(n26273), .B2(
        data_in[3]), .ZN(n17012) );
  INV_X1 U12939 ( .A(n17013), .ZN(n19246) );
  AOI22_X1 U12940 ( .A1(\mem[857][4] ), .A2(n17009), .B1(n26273), .B2(
        data_in[4]), .ZN(n17013) );
  INV_X1 U12941 ( .A(n17014), .ZN(n19245) );
  AOI22_X1 U12942 ( .A1(\mem[857][5] ), .A2(n17009), .B1(n26273), .B2(
        data_in[5]), .ZN(n17014) );
  INV_X1 U12943 ( .A(n17015), .ZN(n19244) );
  AOI22_X1 U12944 ( .A1(\mem[857][6] ), .A2(n17009), .B1(n26273), .B2(
        data_in[6]), .ZN(n17015) );
  INV_X1 U12945 ( .A(n17016), .ZN(n19243) );
  AOI22_X1 U12946 ( .A1(\mem[857][7] ), .A2(n17009), .B1(n26273), .B2(
        data_in[7]), .ZN(n17016) );
  INV_X1 U12947 ( .A(n17017), .ZN(n19242) );
  AOI22_X1 U12948 ( .A1(\mem[858][0] ), .A2(n17018), .B1(n26272), .B2(
        data_in[0]), .ZN(n17017) );
  INV_X1 U12949 ( .A(n17019), .ZN(n19241) );
  AOI22_X1 U12950 ( .A1(\mem[858][1] ), .A2(n17018), .B1(n26272), .B2(
        data_in[1]), .ZN(n17019) );
  INV_X1 U12951 ( .A(n17020), .ZN(n19240) );
  AOI22_X1 U12952 ( .A1(\mem[858][2] ), .A2(n17018), .B1(n26272), .B2(
        data_in[2]), .ZN(n17020) );
  INV_X1 U12953 ( .A(n17021), .ZN(n19239) );
  AOI22_X1 U12954 ( .A1(\mem[858][3] ), .A2(n17018), .B1(n26272), .B2(
        data_in[3]), .ZN(n17021) );
  INV_X1 U12955 ( .A(n17022), .ZN(n19238) );
  AOI22_X1 U12956 ( .A1(\mem[858][4] ), .A2(n17018), .B1(n26272), .B2(
        data_in[4]), .ZN(n17022) );
  INV_X1 U12957 ( .A(n17023), .ZN(n19237) );
  AOI22_X1 U12958 ( .A1(\mem[858][5] ), .A2(n17018), .B1(n26272), .B2(
        data_in[5]), .ZN(n17023) );
  INV_X1 U12959 ( .A(n17024), .ZN(n19236) );
  AOI22_X1 U12960 ( .A1(\mem[858][6] ), .A2(n17018), .B1(n26272), .B2(
        data_in[6]), .ZN(n17024) );
  INV_X1 U12961 ( .A(n17025), .ZN(n19235) );
  AOI22_X1 U12962 ( .A1(\mem[858][7] ), .A2(n17018), .B1(n26272), .B2(
        data_in[7]), .ZN(n17025) );
  INV_X1 U12963 ( .A(n17026), .ZN(n19234) );
  AOI22_X1 U12964 ( .A1(\mem[859][0] ), .A2(n17027), .B1(n26271), .B2(
        data_in[0]), .ZN(n17026) );
  INV_X1 U12965 ( .A(n17028), .ZN(n19233) );
  AOI22_X1 U12966 ( .A1(\mem[859][1] ), .A2(n17027), .B1(n26271), .B2(
        data_in[1]), .ZN(n17028) );
  INV_X1 U12967 ( .A(n17029), .ZN(n19232) );
  AOI22_X1 U12968 ( .A1(\mem[859][2] ), .A2(n17027), .B1(n26271), .B2(
        data_in[2]), .ZN(n17029) );
  INV_X1 U12969 ( .A(n17030), .ZN(n19231) );
  AOI22_X1 U12970 ( .A1(\mem[859][3] ), .A2(n17027), .B1(n26271), .B2(
        data_in[3]), .ZN(n17030) );
  INV_X1 U12971 ( .A(n17031), .ZN(n19230) );
  AOI22_X1 U12972 ( .A1(\mem[859][4] ), .A2(n17027), .B1(n26271), .B2(
        data_in[4]), .ZN(n17031) );
  INV_X1 U12973 ( .A(n17032), .ZN(n19229) );
  AOI22_X1 U12974 ( .A1(\mem[859][5] ), .A2(n17027), .B1(n26271), .B2(
        data_in[5]), .ZN(n17032) );
  INV_X1 U12975 ( .A(n17033), .ZN(n19228) );
  AOI22_X1 U12976 ( .A1(\mem[859][6] ), .A2(n17027), .B1(n26271), .B2(
        data_in[6]), .ZN(n17033) );
  INV_X1 U12977 ( .A(n17034), .ZN(n19227) );
  AOI22_X1 U12978 ( .A1(\mem[859][7] ), .A2(n17027), .B1(n26271), .B2(
        data_in[7]), .ZN(n17034) );
  INV_X1 U12979 ( .A(n17035), .ZN(n19226) );
  AOI22_X1 U12980 ( .A1(\mem[860][0] ), .A2(n17036), .B1(n26270), .B2(
        data_in[0]), .ZN(n17035) );
  INV_X1 U12981 ( .A(n17037), .ZN(n19225) );
  AOI22_X1 U12982 ( .A1(\mem[860][1] ), .A2(n17036), .B1(n26270), .B2(
        data_in[1]), .ZN(n17037) );
  INV_X1 U12983 ( .A(n17038), .ZN(n19224) );
  AOI22_X1 U12984 ( .A1(\mem[860][2] ), .A2(n17036), .B1(n26270), .B2(
        data_in[2]), .ZN(n17038) );
  INV_X1 U12985 ( .A(n17039), .ZN(n19223) );
  AOI22_X1 U12986 ( .A1(\mem[860][3] ), .A2(n17036), .B1(n26270), .B2(
        data_in[3]), .ZN(n17039) );
  INV_X1 U12987 ( .A(n17040), .ZN(n19222) );
  AOI22_X1 U12988 ( .A1(\mem[860][4] ), .A2(n17036), .B1(n26270), .B2(
        data_in[4]), .ZN(n17040) );
  INV_X1 U12989 ( .A(n17041), .ZN(n19221) );
  AOI22_X1 U12990 ( .A1(\mem[860][5] ), .A2(n17036), .B1(n26270), .B2(
        data_in[5]), .ZN(n17041) );
  INV_X1 U12991 ( .A(n17042), .ZN(n19220) );
  AOI22_X1 U12992 ( .A1(\mem[860][6] ), .A2(n17036), .B1(n26270), .B2(
        data_in[6]), .ZN(n17042) );
  INV_X1 U12993 ( .A(n17043), .ZN(n19219) );
  AOI22_X1 U12994 ( .A1(\mem[860][7] ), .A2(n17036), .B1(n26270), .B2(
        data_in[7]), .ZN(n17043) );
  INV_X1 U12995 ( .A(n17044), .ZN(n19218) );
  AOI22_X1 U12996 ( .A1(\mem[861][0] ), .A2(n17045), .B1(n26269), .B2(
        data_in[0]), .ZN(n17044) );
  INV_X1 U12997 ( .A(n17046), .ZN(n19217) );
  AOI22_X1 U12998 ( .A1(\mem[861][1] ), .A2(n17045), .B1(n26269), .B2(
        data_in[1]), .ZN(n17046) );
  INV_X1 U12999 ( .A(n17047), .ZN(n19216) );
  AOI22_X1 U13000 ( .A1(\mem[861][2] ), .A2(n17045), .B1(n26269), .B2(
        data_in[2]), .ZN(n17047) );
  INV_X1 U13001 ( .A(n17048), .ZN(n19215) );
  AOI22_X1 U13002 ( .A1(\mem[861][3] ), .A2(n17045), .B1(n26269), .B2(
        data_in[3]), .ZN(n17048) );
  INV_X1 U13003 ( .A(n17049), .ZN(n19214) );
  AOI22_X1 U13004 ( .A1(\mem[861][4] ), .A2(n17045), .B1(n26269), .B2(
        data_in[4]), .ZN(n17049) );
  INV_X1 U13005 ( .A(n17050), .ZN(n19213) );
  AOI22_X1 U13006 ( .A1(\mem[861][5] ), .A2(n17045), .B1(n26269), .B2(
        data_in[5]), .ZN(n17050) );
  INV_X1 U13007 ( .A(n17051), .ZN(n19212) );
  AOI22_X1 U13008 ( .A1(\mem[861][6] ), .A2(n17045), .B1(n26269), .B2(
        data_in[6]), .ZN(n17051) );
  INV_X1 U13009 ( .A(n17052), .ZN(n19211) );
  AOI22_X1 U13010 ( .A1(\mem[861][7] ), .A2(n17045), .B1(n26269), .B2(
        data_in[7]), .ZN(n17052) );
  INV_X1 U13011 ( .A(n17053), .ZN(n19210) );
  AOI22_X1 U13012 ( .A1(\mem[862][0] ), .A2(n17054), .B1(n26268), .B2(
        data_in[0]), .ZN(n17053) );
  INV_X1 U13013 ( .A(n17055), .ZN(n19209) );
  AOI22_X1 U13014 ( .A1(\mem[862][1] ), .A2(n17054), .B1(n26268), .B2(
        data_in[1]), .ZN(n17055) );
  INV_X1 U13015 ( .A(n17056), .ZN(n19208) );
  AOI22_X1 U13016 ( .A1(\mem[862][2] ), .A2(n17054), .B1(n26268), .B2(
        data_in[2]), .ZN(n17056) );
  INV_X1 U13017 ( .A(n17057), .ZN(n19207) );
  AOI22_X1 U13018 ( .A1(\mem[862][3] ), .A2(n17054), .B1(n26268), .B2(
        data_in[3]), .ZN(n17057) );
  INV_X1 U13019 ( .A(n17058), .ZN(n19206) );
  AOI22_X1 U13020 ( .A1(\mem[862][4] ), .A2(n17054), .B1(n26268), .B2(
        data_in[4]), .ZN(n17058) );
  INV_X1 U13021 ( .A(n17059), .ZN(n19205) );
  AOI22_X1 U13022 ( .A1(\mem[862][5] ), .A2(n17054), .B1(n26268), .B2(
        data_in[5]), .ZN(n17059) );
  INV_X1 U13023 ( .A(n17060), .ZN(n19204) );
  AOI22_X1 U13024 ( .A1(\mem[862][6] ), .A2(n17054), .B1(n26268), .B2(
        data_in[6]), .ZN(n17060) );
  INV_X1 U13025 ( .A(n17061), .ZN(n19203) );
  AOI22_X1 U13026 ( .A1(\mem[862][7] ), .A2(n17054), .B1(n26268), .B2(
        data_in[7]), .ZN(n17061) );
  INV_X1 U13027 ( .A(n17062), .ZN(n19202) );
  AOI22_X1 U13028 ( .A1(\mem[863][0] ), .A2(n17063), .B1(n26267), .B2(
        data_in[0]), .ZN(n17062) );
  INV_X1 U13029 ( .A(n17064), .ZN(n19201) );
  AOI22_X1 U13030 ( .A1(\mem[863][1] ), .A2(n17063), .B1(n26267), .B2(
        data_in[1]), .ZN(n17064) );
  INV_X1 U13031 ( .A(n17065), .ZN(n19200) );
  AOI22_X1 U13032 ( .A1(\mem[863][2] ), .A2(n17063), .B1(n26267), .B2(
        data_in[2]), .ZN(n17065) );
  INV_X1 U13033 ( .A(n17066), .ZN(n19199) );
  AOI22_X1 U13034 ( .A1(\mem[863][3] ), .A2(n17063), .B1(n26267), .B2(
        data_in[3]), .ZN(n17066) );
  INV_X1 U13035 ( .A(n17067), .ZN(n19198) );
  AOI22_X1 U13036 ( .A1(\mem[863][4] ), .A2(n17063), .B1(n26267), .B2(
        data_in[4]), .ZN(n17067) );
  INV_X1 U13037 ( .A(n17068), .ZN(n19197) );
  AOI22_X1 U13038 ( .A1(\mem[863][5] ), .A2(n17063), .B1(n26267), .B2(
        data_in[5]), .ZN(n17068) );
  INV_X1 U13039 ( .A(n17069), .ZN(n19196) );
  AOI22_X1 U13040 ( .A1(\mem[863][6] ), .A2(n17063), .B1(n26267), .B2(
        data_in[6]), .ZN(n17069) );
  INV_X1 U13041 ( .A(n17070), .ZN(n19195) );
  AOI22_X1 U13042 ( .A1(\mem[863][7] ), .A2(n17063), .B1(n26267), .B2(
        data_in[7]), .ZN(n17070) );
  INV_X1 U13043 ( .A(n17144), .ZN(n19130) );
  AOI22_X1 U13044 ( .A1(\mem[872][0] ), .A2(n17145), .B1(n26258), .B2(
        data_in[0]), .ZN(n17144) );
  INV_X1 U13045 ( .A(n17146), .ZN(n19129) );
  AOI22_X1 U13046 ( .A1(\mem[872][1] ), .A2(n17145), .B1(n26258), .B2(
        data_in[1]), .ZN(n17146) );
  INV_X1 U13047 ( .A(n17147), .ZN(n19128) );
  AOI22_X1 U13048 ( .A1(\mem[872][2] ), .A2(n17145), .B1(n26258), .B2(
        data_in[2]), .ZN(n17147) );
  INV_X1 U13049 ( .A(n17148), .ZN(n19127) );
  AOI22_X1 U13050 ( .A1(\mem[872][3] ), .A2(n17145), .B1(n26258), .B2(
        data_in[3]), .ZN(n17148) );
  INV_X1 U13051 ( .A(n17149), .ZN(n19126) );
  AOI22_X1 U13052 ( .A1(\mem[872][4] ), .A2(n17145), .B1(n26258), .B2(
        data_in[4]), .ZN(n17149) );
  INV_X1 U13053 ( .A(n17150), .ZN(n19125) );
  AOI22_X1 U13054 ( .A1(\mem[872][5] ), .A2(n17145), .B1(n26258), .B2(
        data_in[5]), .ZN(n17150) );
  INV_X1 U13055 ( .A(n17151), .ZN(n19124) );
  AOI22_X1 U13056 ( .A1(\mem[872][6] ), .A2(n17145), .B1(n26258), .B2(
        data_in[6]), .ZN(n17151) );
  INV_X1 U13057 ( .A(n17152), .ZN(n19123) );
  AOI22_X1 U13058 ( .A1(\mem[872][7] ), .A2(n17145), .B1(n26258), .B2(
        data_in[7]), .ZN(n17152) );
  INV_X1 U13059 ( .A(n17153), .ZN(n19122) );
  AOI22_X1 U13060 ( .A1(\mem[873][0] ), .A2(n17154), .B1(n26257), .B2(
        data_in[0]), .ZN(n17153) );
  INV_X1 U13061 ( .A(n17155), .ZN(n19121) );
  AOI22_X1 U13062 ( .A1(\mem[873][1] ), .A2(n17154), .B1(n26257), .B2(
        data_in[1]), .ZN(n17155) );
  INV_X1 U13063 ( .A(n17156), .ZN(n19120) );
  AOI22_X1 U13064 ( .A1(\mem[873][2] ), .A2(n17154), .B1(n26257), .B2(
        data_in[2]), .ZN(n17156) );
  INV_X1 U13065 ( .A(n17157), .ZN(n19119) );
  AOI22_X1 U13066 ( .A1(\mem[873][3] ), .A2(n17154), .B1(n26257), .B2(
        data_in[3]), .ZN(n17157) );
  INV_X1 U13067 ( .A(n17158), .ZN(n19118) );
  AOI22_X1 U13068 ( .A1(\mem[873][4] ), .A2(n17154), .B1(n26257), .B2(
        data_in[4]), .ZN(n17158) );
  INV_X1 U13069 ( .A(n17159), .ZN(n19117) );
  AOI22_X1 U13070 ( .A1(\mem[873][5] ), .A2(n17154), .B1(n26257), .B2(
        data_in[5]), .ZN(n17159) );
  INV_X1 U13071 ( .A(n17160), .ZN(n19116) );
  AOI22_X1 U13072 ( .A1(\mem[873][6] ), .A2(n17154), .B1(n26257), .B2(
        data_in[6]), .ZN(n17160) );
  INV_X1 U13073 ( .A(n17161), .ZN(n19115) );
  AOI22_X1 U13074 ( .A1(\mem[873][7] ), .A2(n17154), .B1(n26257), .B2(
        data_in[7]), .ZN(n17161) );
  INV_X1 U13075 ( .A(n17162), .ZN(n19114) );
  AOI22_X1 U13076 ( .A1(\mem[874][0] ), .A2(n17163), .B1(n26256), .B2(
        data_in[0]), .ZN(n17162) );
  INV_X1 U13077 ( .A(n17164), .ZN(n19113) );
  AOI22_X1 U13078 ( .A1(\mem[874][1] ), .A2(n17163), .B1(n26256), .B2(
        data_in[1]), .ZN(n17164) );
  INV_X1 U13079 ( .A(n17165), .ZN(n19112) );
  AOI22_X1 U13080 ( .A1(\mem[874][2] ), .A2(n17163), .B1(n26256), .B2(
        data_in[2]), .ZN(n17165) );
  INV_X1 U13081 ( .A(n17166), .ZN(n19111) );
  AOI22_X1 U13082 ( .A1(\mem[874][3] ), .A2(n17163), .B1(n26256), .B2(
        data_in[3]), .ZN(n17166) );
  INV_X1 U13083 ( .A(n17167), .ZN(n19110) );
  AOI22_X1 U13084 ( .A1(\mem[874][4] ), .A2(n17163), .B1(n26256), .B2(
        data_in[4]), .ZN(n17167) );
  INV_X1 U13085 ( .A(n17168), .ZN(n19109) );
  AOI22_X1 U13086 ( .A1(\mem[874][5] ), .A2(n17163), .B1(n26256), .B2(
        data_in[5]), .ZN(n17168) );
  INV_X1 U13087 ( .A(n17169), .ZN(n19108) );
  AOI22_X1 U13088 ( .A1(\mem[874][6] ), .A2(n17163), .B1(n26256), .B2(
        data_in[6]), .ZN(n17169) );
  INV_X1 U13089 ( .A(n17170), .ZN(n19107) );
  AOI22_X1 U13090 ( .A1(\mem[874][7] ), .A2(n17163), .B1(n26256), .B2(
        data_in[7]), .ZN(n17170) );
  INV_X1 U13091 ( .A(n17171), .ZN(n19106) );
  AOI22_X1 U13092 ( .A1(\mem[875][0] ), .A2(n17172), .B1(n26255), .B2(
        data_in[0]), .ZN(n17171) );
  INV_X1 U13093 ( .A(n17173), .ZN(n19105) );
  AOI22_X1 U13094 ( .A1(\mem[875][1] ), .A2(n17172), .B1(n26255), .B2(
        data_in[1]), .ZN(n17173) );
  INV_X1 U13095 ( .A(n17174), .ZN(n19104) );
  AOI22_X1 U13096 ( .A1(\mem[875][2] ), .A2(n17172), .B1(n26255), .B2(
        data_in[2]), .ZN(n17174) );
  INV_X1 U13097 ( .A(n17175), .ZN(n19103) );
  AOI22_X1 U13098 ( .A1(\mem[875][3] ), .A2(n17172), .B1(n26255), .B2(
        data_in[3]), .ZN(n17175) );
  INV_X1 U13099 ( .A(n17176), .ZN(n19102) );
  AOI22_X1 U13100 ( .A1(\mem[875][4] ), .A2(n17172), .B1(n26255), .B2(
        data_in[4]), .ZN(n17176) );
  INV_X1 U13101 ( .A(n17177), .ZN(n19101) );
  AOI22_X1 U13102 ( .A1(\mem[875][5] ), .A2(n17172), .B1(n26255), .B2(
        data_in[5]), .ZN(n17177) );
  INV_X1 U13103 ( .A(n17178), .ZN(n19100) );
  AOI22_X1 U13104 ( .A1(\mem[875][6] ), .A2(n17172), .B1(n26255), .B2(
        data_in[6]), .ZN(n17178) );
  INV_X1 U13105 ( .A(n17179), .ZN(n19099) );
  AOI22_X1 U13106 ( .A1(\mem[875][7] ), .A2(n17172), .B1(n26255), .B2(
        data_in[7]), .ZN(n17179) );
  INV_X1 U13107 ( .A(n17180), .ZN(n19098) );
  AOI22_X1 U13108 ( .A1(\mem[876][0] ), .A2(n17181), .B1(n26254), .B2(
        data_in[0]), .ZN(n17180) );
  INV_X1 U13109 ( .A(n17182), .ZN(n19097) );
  AOI22_X1 U13110 ( .A1(\mem[876][1] ), .A2(n17181), .B1(n26254), .B2(
        data_in[1]), .ZN(n17182) );
  INV_X1 U13111 ( .A(n17183), .ZN(n19096) );
  AOI22_X1 U13112 ( .A1(\mem[876][2] ), .A2(n17181), .B1(n26254), .B2(
        data_in[2]), .ZN(n17183) );
  INV_X1 U13113 ( .A(n17184), .ZN(n19095) );
  AOI22_X1 U13114 ( .A1(\mem[876][3] ), .A2(n17181), .B1(n26254), .B2(
        data_in[3]), .ZN(n17184) );
  INV_X1 U13115 ( .A(n17185), .ZN(n19094) );
  AOI22_X1 U13116 ( .A1(\mem[876][4] ), .A2(n17181), .B1(n26254), .B2(
        data_in[4]), .ZN(n17185) );
  INV_X1 U13117 ( .A(n17186), .ZN(n19093) );
  AOI22_X1 U13118 ( .A1(\mem[876][5] ), .A2(n17181), .B1(n26254), .B2(
        data_in[5]), .ZN(n17186) );
  INV_X1 U13119 ( .A(n17187), .ZN(n19092) );
  AOI22_X1 U13120 ( .A1(\mem[876][6] ), .A2(n17181), .B1(n26254), .B2(
        data_in[6]), .ZN(n17187) );
  INV_X1 U13121 ( .A(n17188), .ZN(n19091) );
  AOI22_X1 U13122 ( .A1(\mem[876][7] ), .A2(n17181), .B1(n26254), .B2(
        data_in[7]), .ZN(n17188) );
  INV_X1 U13123 ( .A(n17189), .ZN(n19090) );
  AOI22_X1 U13124 ( .A1(\mem[877][0] ), .A2(n17190), .B1(n26253), .B2(
        data_in[0]), .ZN(n17189) );
  INV_X1 U13125 ( .A(n17191), .ZN(n19089) );
  AOI22_X1 U13126 ( .A1(\mem[877][1] ), .A2(n17190), .B1(n26253), .B2(
        data_in[1]), .ZN(n17191) );
  INV_X1 U13127 ( .A(n17192), .ZN(n19088) );
  AOI22_X1 U13128 ( .A1(\mem[877][2] ), .A2(n17190), .B1(n26253), .B2(
        data_in[2]), .ZN(n17192) );
  INV_X1 U13129 ( .A(n17193), .ZN(n19087) );
  AOI22_X1 U13130 ( .A1(\mem[877][3] ), .A2(n17190), .B1(n26253), .B2(
        data_in[3]), .ZN(n17193) );
  INV_X1 U13131 ( .A(n17194), .ZN(n19086) );
  AOI22_X1 U13132 ( .A1(\mem[877][4] ), .A2(n17190), .B1(n26253), .B2(
        data_in[4]), .ZN(n17194) );
  INV_X1 U13133 ( .A(n17195), .ZN(n19085) );
  AOI22_X1 U13134 ( .A1(\mem[877][5] ), .A2(n17190), .B1(n26253), .B2(
        data_in[5]), .ZN(n17195) );
  INV_X1 U13135 ( .A(n17196), .ZN(n19084) );
  AOI22_X1 U13136 ( .A1(\mem[877][6] ), .A2(n17190), .B1(n26253), .B2(
        data_in[6]), .ZN(n17196) );
  INV_X1 U13137 ( .A(n17197), .ZN(n19083) );
  AOI22_X1 U13138 ( .A1(\mem[877][7] ), .A2(n17190), .B1(n26253), .B2(
        data_in[7]), .ZN(n17197) );
  INV_X1 U13139 ( .A(n17198), .ZN(n19082) );
  AOI22_X1 U13140 ( .A1(\mem[878][0] ), .A2(n17199), .B1(n26252), .B2(
        data_in[0]), .ZN(n17198) );
  INV_X1 U13141 ( .A(n17200), .ZN(n19081) );
  AOI22_X1 U13142 ( .A1(\mem[878][1] ), .A2(n17199), .B1(n26252), .B2(
        data_in[1]), .ZN(n17200) );
  INV_X1 U13143 ( .A(n17201), .ZN(n19080) );
  AOI22_X1 U13144 ( .A1(\mem[878][2] ), .A2(n17199), .B1(n26252), .B2(
        data_in[2]), .ZN(n17201) );
  INV_X1 U13145 ( .A(n17202), .ZN(n19079) );
  AOI22_X1 U13146 ( .A1(\mem[878][3] ), .A2(n17199), .B1(n26252), .B2(
        data_in[3]), .ZN(n17202) );
  INV_X1 U13147 ( .A(n17203), .ZN(n19078) );
  AOI22_X1 U13148 ( .A1(\mem[878][4] ), .A2(n17199), .B1(n26252), .B2(
        data_in[4]), .ZN(n17203) );
  INV_X1 U13149 ( .A(n17204), .ZN(n19077) );
  AOI22_X1 U13150 ( .A1(\mem[878][5] ), .A2(n17199), .B1(n26252), .B2(
        data_in[5]), .ZN(n17204) );
  INV_X1 U13151 ( .A(n17205), .ZN(n19076) );
  AOI22_X1 U13152 ( .A1(\mem[878][6] ), .A2(n17199), .B1(n26252), .B2(
        data_in[6]), .ZN(n17205) );
  INV_X1 U13153 ( .A(n17206), .ZN(n19075) );
  AOI22_X1 U13154 ( .A1(\mem[878][7] ), .A2(n17199), .B1(n26252), .B2(
        data_in[7]), .ZN(n17206) );
  INV_X1 U13155 ( .A(n17207), .ZN(n19074) );
  AOI22_X1 U13156 ( .A1(\mem[879][0] ), .A2(n17208), .B1(n26251), .B2(
        data_in[0]), .ZN(n17207) );
  INV_X1 U13157 ( .A(n17209), .ZN(n19073) );
  AOI22_X1 U13158 ( .A1(\mem[879][1] ), .A2(n17208), .B1(n26251), .B2(
        data_in[1]), .ZN(n17209) );
  INV_X1 U13159 ( .A(n17210), .ZN(n19072) );
  AOI22_X1 U13160 ( .A1(\mem[879][2] ), .A2(n17208), .B1(n26251), .B2(
        data_in[2]), .ZN(n17210) );
  INV_X1 U13161 ( .A(n17211), .ZN(n19071) );
  AOI22_X1 U13162 ( .A1(\mem[879][3] ), .A2(n17208), .B1(n26251), .B2(
        data_in[3]), .ZN(n17211) );
  INV_X1 U13163 ( .A(n17212), .ZN(n19070) );
  AOI22_X1 U13164 ( .A1(\mem[879][4] ), .A2(n17208), .B1(n26251), .B2(
        data_in[4]), .ZN(n17212) );
  INV_X1 U13165 ( .A(n17213), .ZN(n19069) );
  AOI22_X1 U13166 ( .A1(\mem[879][5] ), .A2(n17208), .B1(n26251), .B2(
        data_in[5]), .ZN(n17213) );
  INV_X1 U13167 ( .A(n17214), .ZN(n19068) );
  AOI22_X1 U13168 ( .A1(\mem[879][6] ), .A2(n17208), .B1(n26251), .B2(
        data_in[6]), .ZN(n17214) );
  INV_X1 U13169 ( .A(n17215), .ZN(n19067) );
  AOI22_X1 U13170 ( .A1(\mem[879][7] ), .A2(n17208), .B1(n26251), .B2(
        data_in[7]), .ZN(n17215) );
  INV_X1 U13171 ( .A(n17216), .ZN(n19066) );
  AOI22_X1 U13172 ( .A1(\mem[880][0] ), .A2(n17217), .B1(n26250), .B2(
        data_in[0]), .ZN(n17216) );
  INV_X1 U13173 ( .A(n17218), .ZN(n19065) );
  AOI22_X1 U13174 ( .A1(\mem[880][1] ), .A2(n17217), .B1(n26250), .B2(
        data_in[1]), .ZN(n17218) );
  INV_X1 U13175 ( .A(n17219), .ZN(n19064) );
  AOI22_X1 U13176 ( .A1(\mem[880][2] ), .A2(n17217), .B1(n26250), .B2(
        data_in[2]), .ZN(n17219) );
  INV_X1 U13177 ( .A(n17220), .ZN(n19063) );
  AOI22_X1 U13178 ( .A1(\mem[880][3] ), .A2(n17217), .B1(n26250), .B2(
        data_in[3]), .ZN(n17220) );
  INV_X1 U13179 ( .A(n17221), .ZN(n19062) );
  AOI22_X1 U13180 ( .A1(\mem[880][4] ), .A2(n17217), .B1(n26250), .B2(
        data_in[4]), .ZN(n17221) );
  INV_X1 U13181 ( .A(n17222), .ZN(n19061) );
  AOI22_X1 U13182 ( .A1(\mem[880][5] ), .A2(n17217), .B1(n26250), .B2(
        data_in[5]), .ZN(n17222) );
  INV_X1 U13183 ( .A(n17223), .ZN(n19060) );
  AOI22_X1 U13184 ( .A1(\mem[880][6] ), .A2(n17217), .B1(n26250), .B2(
        data_in[6]), .ZN(n17223) );
  INV_X1 U13185 ( .A(n17224), .ZN(n19059) );
  AOI22_X1 U13186 ( .A1(\mem[880][7] ), .A2(n17217), .B1(n26250), .B2(
        data_in[7]), .ZN(n17224) );
  INV_X1 U13187 ( .A(n17225), .ZN(n19058) );
  AOI22_X1 U13188 ( .A1(\mem[881][0] ), .A2(n17226), .B1(n26249), .B2(
        data_in[0]), .ZN(n17225) );
  INV_X1 U13189 ( .A(n17227), .ZN(n19057) );
  AOI22_X1 U13190 ( .A1(\mem[881][1] ), .A2(n17226), .B1(n26249), .B2(
        data_in[1]), .ZN(n17227) );
  INV_X1 U13191 ( .A(n17228), .ZN(n19056) );
  AOI22_X1 U13192 ( .A1(\mem[881][2] ), .A2(n17226), .B1(n26249), .B2(
        data_in[2]), .ZN(n17228) );
  INV_X1 U13193 ( .A(n17229), .ZN(n19055) );
  AOI22_X1 U13194 ( .A1(\mem[881][3] ), .A2(n17226), .B1(n26249), .B2(
        data_in[3]), .ZN(n17229) );
  INV_X1 U13195 ( .A(n17230), .ZN(n19054) );
  AOI22_X1 U13196 ( .A1(\mem[881][4] ), .A2(n17226), .B1(n26249), .B2(
        data_in[4]), .ZN(n17230) );
  INV_X1 U13197 ( .A(n17231), .ZN(n19053) );
  AOI22_X1 U13198 ( .A1(\mem[881][5] ), .A2(n17226), .B1(n26249), .B2(
        data_in[5]), .ZN(n17231) );
  INV_X1 U13199 ( .A(n17232), .ZN(n19052) );
  AOI22_X1 U13200 ( .A1(\mem[881][6] ), .A2(n17226), .B1(n26249), .B2(
        data_in[6]), .ZN(n17232) );
  INV_X1 U13201 ( .A(n17233), .ZN(n19051) );
  AOI22_X1 U13202 ( .A1(\mem[881][7] ), .A2(n17226), .B1(n26249), .B2(
        data_in[7]), .ZN(n17233) );
  INV_X1 U13203 ( .A(n17234), .ZN(n19050) );
  AOI22_X1 U13204 ( .A1(\mem[882][0] ), .A2(n17235), .B1(n26248), .B2(
        data_in[0]), .ZN(n17234) );
  INV_X1 U13205 ( .A(n17236), .ZN(n19049) );
  AOI22_X1 U13206 ( .A1(\mem[882][1] ), .A2(n17235), .B1(n26248), .B2(
        data_in[1]), .ZN(n17236) );
  INV_X1 U13207 ( .A(n17237), .ZN(n19048) );
  AOI22_X1 U13208 ( .A1(\mem[882][2] ), .A2(n17235), .B1(n26248), .B2(
        data_in[2]), .ZN(n17237) );
  INV_X1 U13209 ( .A(n17238), .ZN(n19047) );
  AOI22_X1 U13210 ( .A1(\mem[882][3] ), .A2(n17235), .B1(n26248), .B2(
        data_in[3]), .ZN(n17238) );
  INV_X1 U13211 ( .A(n17239), .ZN(n19046) );
  AOI22_X1 U13212 ( .A1(\mem[882][4] ), .A2(n17235), .B1(n26248), .B2(
        data_in[4]), .ZN(n17239) );
  INV_X1 U13213 ( .A(n17240), .ZN(n19045) );
  AOI22_X1 U13214 ( .A1(\mem[882][5] ), .A2(n17235), .B1(n26248), .B2(
        data_in[5]), .ZN(n17240) );
  INV_X1 U13215 ( .A(n17241), .ZN(n19044) );
  AOI22_X1 U13216 ( .A1(\mem[882][6] ), .A2(n17235), .B1(n26248), .B2(
        data_in[6]), .ZN(n17241) );
  INV_X1 U13217 ( .A(n17242), .ZN(n19043) );
  AOI22_X1 U13218 ( .A1(\mem[882][7] ), .A2(n17235), .B1(n26248), .B2(
        data_in[7]), .ZN(n17242) );
  INV_X1 U13219 ( .A(n17243), .ZN(n19042) );
  AOI22_X1 U13220 ( .A1(\mem[883][0] ), .A2(n17244), .B1(n26247), .B2(
        data_in[0]), .ZN(n17243) );
  INV_X1 U13221 ( .A(n17245), .ZN(n19041) );
  AOI22_X1 U13222 ( .A1(\mem[883][1] ), .A2(n17244), .B1(n26247), .B2(
        data_in[1]), .ZN(n17245) );
  INV_X1 U13223 ( .A(n17246), .ZN(n19040) );
  AOI22_X1 U13224 ( .A1(\mem[883][2] ), .A2(n17244), .B1(n26247), .B2(
        data_in[2]), .ZN(n17246) );
  INV_X1 U13225 ( .A(n17247), .ZN(n19039) );
  AOI22_X1 U13226 ( .A1(\mem[883][3] ), .A2(n17244), .B1(n26247), .B2(
        data_in[3]), .ZN(n17247) );
  INV_X1 U13227 ( .A(n17248), .ZN(n19038) );
  AOI22_X1 U13228 ( .A1(\mem[883][4] ), .A2(n17244), .B1(n26247), .B2(
        data_in[4]), .ZN(n17248) );
  INV_X1 U13229 ( .A(n17249), .ZN(n19037) );
  AOI22_X1 U13230 ( .A1(\mem[883][5] ), .A2(n17244), .B1(n26247), .B2(
        data_in[5]), .ZN(n17249) );
  INV_X1 U13231 ( .A(n17250), .ZN(n19036) );
  AOI22_X1 U13232 ( .A1(\mem[883][6] ), .A2(n17244), .B1(n26247), .B2(
        data_in[6]), .ZN(n17250) );
  INV_X1 U13233 ( .A(n17251), .ZN(n19035) );
  AOI22_X1 U13234 ( .A1(\mem[883][7] ), .A2(n17244), .B1(n26247), .B2(
        data_in[7]), .ZN(n17251) );
  INV_X1 U13235 ( .A(n17252), .ZN(n19034) );
  AOI22_X1 U13236 ( .A1(\mem[884][0] ), .A2(n17253), .B1(n26246), .B2(
        data_in[0]), .ZN(n17252) );
  INV_X1 U13237 ( .A(n17254), .ZN(n19033) );
  AOI22_X1 U13238 ( .A1(\mem[884][1] ), .A2(n17253), .B1(n26246), .B2(
        data_in[1]), .ZN(n17254) );
  INV_X1 U13239 ( .A(n17255), .ZN(n19032) );
  AOI22_X1 U13240 ( .A1(\mem[884][2] ), .A2(n17253), .B1(n26246), .B2(
        data_in[2]), .ZN(n17255) );
  INV_X1 U13241 ( .A(n17256), .ZN(n19031) );
  AOI22_X1 U13242 ( .A1(\mem[884][3] ), .A2(n17253), .B1(n26246), .B2(
        data_in[3]), .ZN(n17256) );
  INV_X1 U13243 ( .A(n17257), .ZN(n19030) );
  AOI22_X1 U13244 ( .A1(\mem[884][4] ), .A2(n17253), .B1(n26246), .B2(
        data_in[4]), .ZN(n17257) );
  INV_X1 U13245 ( .A(n17258), .ZN(n19029) );
  AOI22_X1 U13246 ( .A1(\mem[884][5] ), .A2(n17253), .B1(n26246), .B2(
        data_in[5]), .ZN(n17258) );
  INV_X1 U13247 ( .A(n17259), .ZN(n19028) );
  AOI22_X1 U13248 ( .A1(\mem[884][6] ), .A2(n17253), .B1(n26246), .B2(
        data_in[6]), .ZN(n17259) );
  INV_X1 U13249 ( .A(n17260), .ZN(n19027) );
  AOI22_X1 U13250 ( .A1(\mem[884][7] ), .A2(n17253), .B1(n26246), .B2(
        data_in[7]), .ZN(n17260) );
  INV_X1 U13251 ( .A(n17261), .ZN(n19026) );
  AOI22_X1 U13252 ( .A1(\mem[885][0] ), .A2(n17262), .B1(n26245), .B2(
        data_in[0]), .ZN(n17261) );
  INV_X1 U13253 ( .A(n17263), .ZN(n19025) );
  AOI22_X1 U13254 ( .A1(\mem[885][1] ), .A2(n17262), .B1(n26245), .B2(
        data_in[1]), .ZN(n17263) );
  INV_X1 U13255 ( .A(n17264), .ZN(n19024) );
  AOI22_X1 U13256 ( .A1(\mem[885][2] ), .A2(n17262), .B1(n26245), .B2(
        data_in[2]), .ZN(n17264) );
  INV_X1 U13257 ( .A(n17265), .ZN(n19023) );
  AOI22_X1 U13258 ( .A1(\mem[885][3] ), .A2(n17262), .B1(n26245), .B2(
        data_in[3]), .ZN(n17265) );
  INV_X1 U13259 ( .A(n17266), .ZN(n19022) );
  AOI22_X1 U13260 ( .A1(\mem[885][4] ), .A2(n17262), .B1(n26245), .B2(
        data_in[4]), .ZN(n17266) );
  INV_X1 U13261 ( .A(n17267), .ZN(n19021) );
  AOI22_X1 U13262 ( .A1(\mem[885][5] ), .A2(n17262), .B1(n26245), .B2(
        data_in[5]), .ZN(n17267) );
  INV_X1 U13263 ( .A(n17268), .ZN(n19020) );
  AOI22_X1 U13264 ( .A1(\mem[885][6] ), .A2(n17262), .B1(n26245), .B2(
        data_in[6]), .ZN(n17268) );
  INV_X1 U13265 ( .A(n17269), .ZN(n19019) );
  AOI22_X1 U13266 ( .A1(\mem[885][7] ), .A2(n17262), .B1(n26245), .B2(
        data_in[7]), .ZN(n17269) );
  INV_X1 U13267 ( .A(n17270), .ZN(n19018) );
  AOI22_X1 U13268 ( .A1(\mem[886][0] ), .A2(n17271), .B1(n26244), .B2(
        data_in[0]), .ZN(n17270) );
  INV_X1 U13269 ( .A(n17272), .ZN(n19017) );
  AOI22_X1 U13270 ( .A1(\mem[886][1] ), .A2(n17271), .B1(n26244), .B2(
        data_in[1]), .ZN(n17272) );
  INV_X1 U13271 ( .A(n17273), .ZN(n19016) );
  AOI22_X1 U13272 ( .A1(\mem[886][2] ), .A2(n17271), .B1(n26244), .B2(
        data_in[2]), .ZN(n17273) );
  INV_X1 U13273 ( .A(n17274), .ZN(n19015) );
  AOI22_X1 U13274 ( .A1(\mem[886][3] ), .A2(n17271), .B1(n26244), .B2(
        data_in[3]), .ZN(n17274) );
  INV_X1 U13275 ( .A(n17275), .ZN(n19014) );
  AOI22_X1 U13276 ( .A1(\mem[886][4] ), .A2(n17271), .B1(n26244), .B2(
        data_in[4]), .ZN(n17275) );
  INV_X1 U13277 ( .A(n17276), .ZN(n19013) );
  AOI22_X1 U13278 ( .A1(\mem[886][5] ), .A2(n17271), .B1(n26244), .B2(
        data_in[5]), .ZN(n17276) );
  INV_X1 U13279 ( .A(n17277), .ZN(n19012) );
  AOI22_X1 U13280 ( .A1(\mem[886][6] ), .A2(n17271), .B1(n26244), .B2(
        data_in[6]), .ZN(n17277) );
  INV_X1 U13281 ( .A(n17278), .ZN(n19011) );
  AOI22_X1 U13282 ( .A1(\mem[886][7] ), .A2(n17271), .B1(n26244), .B2(
        data_in[7]), .ZN(n17278) );
  INV_X1 U13283 ( .A(n17279), .ZN(n19010) );
  AOI22_X1 U13284 ( .A1(\mem[887][0] ), .A2(n17280), .B1(n26243), .B2(
        data_in[0]), .ZN(n17279) );
  INV_X1 U13285 ( .A(n17281), .ZN(n19009) );
  AOI22_X1 U13286 ( .A1(\mem[887][1] ), .A2(n17280), .B1(n26243), .B2(
        data_in[1]), .ZN(n17281) );
  INV_X1 U13287 ( .A(n17282), .ZN(n19008) );
  AOI22_X1 U13288 ( .A1(\mem[887][2] ), .A2(n17280), .B1(n26243), .B2(
        data_in[2]), .ZN(n17282) );
  INV_X1 U13289 ( .A(n17283), .ZN(n19007) );
  AOI22_X1 U13290 ( .A1(\mem[887][3] ), .A2(n17280), .B1(n26243), .B2(
        data_in[3]), .ZN(n17283) );
  INV_X1 U13291 ( .A(n17284), .ZN(n19006) );
  AOI22_X1 U13292 ( .A1(\mem[887][4] ), .A2(n17280), .B1(n26243), .B2(
        data_in[4]), .ZN(n17284) );
  INV_X1 U13293 ( .A(n17285), .ZN(n19005) );
  AOI22_X1 U13294 ( .A1(\mem[887][5] ), .A2(n17280), .B1(n26243), .B2(
        data_in[5]), .ZN(n17285) );
  INV_X1 U13295 ( .A(n17286), .ZN(n19004) );
  AOI22_X1 U13296 ( .A1(\mem[887][6] ), .A2(n17280), .B1(n26243), .B2(
        data_in[6]), .ZN(n17286) );
  INV_X1 U13297 ( .A(n17287), .ZN(n19003) );
  AOI22_X1 U13298 ( .A1(\mem[887][7] ), .A2(n17280), .B1(n26243), .B2(
        data_in[7]), .ZN(n17287) );
  INV_X1 U13299 ( .A(n17288), .ZN(n19002) );
  AOI22_X1 U13300 ( .A1(\mem[888][0] ), .A2(n17289), .B1(n26242), .B2(
        data_in[0]), .ZN(n17288) );
  INV_X1 U13301 ( .A(n17290), .ZN(n19001) );
  AOI22_X1 U13302 ( .A1(\mem[888][1] ), .A2(n17289), .B1(n26242), .B2(
        data_in[1]), .ZN(n17290) );
  INV_X1 U13303 ( .A(n17291), .ZN(n19000) );
  AOI22_X1 U13304 ( .A1(\mem[888][2] ), .A2(n17289), .B1(n26242), .B2(
        data_in[2]), .ZN(n17291) );
  INV_X1 U13305 ( .A(n17292), .ZN(n18999) );
  AOI22_X1 U13306 ( .A1(\mem[888][3] ), .A2(n17289), .B1(n26242), .B2(
        data_in[3]), .ZN(n17292) );
  INV_X1 U13307 ( .A(n17293), .ZN(n18998) );
  AOI22_X1 U13308 ( .A1(\mem[888][4] ), .A2(n17289), .B1(n26242), .B2(
        data_in[4]), .ZN(n17293) );
  INV_X1 U13309 ( .A(n17294), .ZN(n18997) );
  AOI22_X1 U13310 ( .A1(\mem[888][5] ), .A2(n17289), .B1(n26242), .B2(
        data_in[5]), .ZN(n17294) );
  INV_X1 U13311 ( .A(n17295), .ZN(n18996) );
  AOI22_X1 U13312 ( .A1(\mem[888][6] ), .A2(n17289), .B1(n26242), .B2(
        data_in[6]), .ZN(n17295) );
  INV_X1 U13313 ( .A(n17296), .ZN(n18995) );
  AOI22_X1 U13314 ( .A1(\mem[888][7] ), .A2(n17289), .B1(n26242), .B2(
        data_in[7]), .ZN(n17296) );
  INV_X1 U13315 ( .A(n17297), .ZN(n18994) );
  AOI22_X1 U13316 ( .A1(\mem[889][0] ), .A2(n17298), .B1(n26241), .B2(
        data_in[0]), .ZN(n17297) );
  INV_X1 U13317 ( .A(n17299), .ZN(n18993) );
  AOI22_X1 U13318 ( .A1(\mem[889][1] ), .A2(n17298), .B1(n26241), .B2(
        data_in[1]), .ZN(n17299) );
  INV_X1 U13319 ( .A(n17300), .ZN(n18992) );
  AOI22_X1 U13320 ( .A1(\mem[889][2] ), .A2(n17298), .B1(n26241), .B2(
        data_in[2]), .ZN(n17300) );
  INV_X1 U13321 ( .A(n17301), .ZN(n18991) );
  AOI22_X1 U13322 ( .A1(\mem[889][3] ), .A2(n17298), .B1(n26241), .B2(
        data_in[3]), .ZN(n17301) );
  INV_X1 U13323 ( .A(n17302), .ZN(n18990) );
  AOI22_X1 U13324 ( .A1(\mem[889][4] ), .A2(n17298), .B1(n26241), .B2(
        data_in[4]), .ZN(n17302) );
  INV_X1 U13325 ( .A(n17303), .ZN(n18989) );
  AOI22_X1 U13326 ( .A1(\mem[889][5] ), .A2(n17298), .B1(n26241), .B2(
        data_in[5]), .ZN(n17303) );
  INV_X1 U13327 ( .A(n17304), .ZN(n18988) );
  AOI22_X1 U13328 ( .A1(\mem[889][6] ), .A2(n17298), .B1(n26241), .B2(
        data_in[6]), .ZN(n17304) );
  INV_X1 U13329 ( .A(n17305), .ZN(n18987) );
  AOI22_X1 U13330 ( .A1(\mem[889][7] ), .A2(n17298), .B1(n26241), .B2(
        data_in[7]), .ZN(n17305) );
  INV_X1 U13331 ( .A(n17306), .ZN(n18986) );
  AOI22_X1 U13332 ( .A1(\mem[890][0] ), .A2(n17307), .B1(n26240), .B2(
        data_in[0]), .ZN(n17306) );
  INV_X1 U13333 ( .A(n17308), .ZN(n18985) );
  AOI22_X1 U13334 ( .A1(\mem[890][1] ), .A2(n17307), .B1(n26240), .B2(
        data_in[1]), .ZN(n17308) );
  INV_X1 U13335 ( .A(n17309), .ZN(n18984) );
  AOI22_X1 U13336 ( .A1(\mem[890][2] ), .A2(n17307), .B1(n26240), .B2(
        data_in[2]), .ZN(n17309) );
  INV_X1 U13337 ( .A(n17310), .ZN(n18983) );
  AOI22_X1 U13338 ( .A1(\mem[890][3] ), .A2(n17307), .B1(n26240), .B2(
        data_in[3]), .ZN(n17310) );
  INV_X1 U13339 ( .A(n17311), .ZN(n18982) );
  AOI22_X1 U13340 ( .A1(\mem[890][4] ), .A2(n17307), .B1(n26240), .B2(
        data_in[4]), .ZN(n17311) );
  INV_X1 U13341 ( .A(n17312), .ZN(n18981) );
  AOI22_X1 U13342 ( .A1(\mem[890][5] ), .A2(n17307), .B1(n26240), .B2(
        data_in[5]), .ZN(n17312) );
  INV_X1 U13343 ( .A(n17313), .ZN(n18980) );
  AOI22_X1 U13344 ( .A1(\mem[890][6] ), .A2(n17307), .B1(n26240), .B2(
        data_in[6]), .ZN(n17313) );
  INV_X1 U13345 ( .A(n17314), .ZN(n18979) );
  AOI22_X1 U13346 ( .A1(\mem[890][7] ), .A2(n17307), .B1(n26240), .B2(
        data_in[7]), .ZN(n17314) );
  INV_X1 U13347 ( .A(n17315), .ZN(n18978) );
  AOI22_X1 U13348 ( .A1(\mem[891][0] ), .A2(n17316), .B1(n26239), .B2(
        data_in[0]), .ZN(n17315) );
  INV_X1 U13349 ( .A(n17317), .ZN(n18977) );
  AOI22_X1 U13350 ( .A1(\mem[891][1] ), .A2(n17316), .B1(n26239), .B2(
        data_in[1]), .ZN(n17317) );
  INV_X1 U13351 ( .A(n17318), .ZN(n18976) );
  AOI22_X1 U13352 ( .A1(\mem[891][2] ), .A2(n17316), .B1(n26239), .B2(
        data_in[2]), .ZN(n17318) );
  INV_X1 U13353 ( .A(n17319), .ZN(n18975) );
  AOI22_X1 U13354 ( .A1(\mem[891][3] ), .A2(n17316), .B1(n26239), .B2(
        data_in[3]), .ZN(n17319) );
  INV_X1 U13355 ( .A(n17320), .ZN(n18974) );
  AOI22_X1 U13356 ( .A1(\mem[891][4] ), .A2(n17316), .B1(n26239), .B2(
        data_in[4]), .ZN(n17320) );
  INV_X1 U13357 ( .A(n17321), .ZN(n18973) );
  AOI22_X1 U13358 ( .A1(\mem[891][5] ), .A2(n17316), .B1(n26239), .B2(
        data_in[5]), .ZN(n17321) );
  INV_X1 U13359 ( .A(n17322), .ZN(n18972) );
  AOI22_X1 U13360 ( .A1(\mem[891][6] ), .A2(n17316), .B1(n26239), .B2(
        data_in[6]), .ZN(n17322) );
  INV_X1 U13361 ( .A(n17323), .ZN(n18971) );
  AOI22_X1 U13362 ( .A1(\mem[891][7] ), .A2(n17316), .B1(n26239), .B2(
        data_in[7]), .ZN(n17323) );
  INV_X1 U13363 ( .A(n17324), .ZN(n18970) );
  AOI22_X1 U13364 ( .A1(\mem[892][0] ), .A2(n17325), .B1(n26238), .B2(
        data_in[0]), .ZN(n17324) );
  INV_X1 U13365 ( .A(n17326), .ZN(n18969) );
  AOI22_X1 U13366 ( .A1(\mem[892][1] ), .A2(n17325), .B1(n26238), .B2(
        data_in[1]), .ZN(n17326) );
  INV_X1 U13367 ( .A(n17327), .ZN(n18968) );
  AOI22_X1 U13368 ( .A1(\mem[892][2] ), .A2(n17325), .B1(n26238), .B2(
        data_in[2]), .ZN(n17327) );
  INV_X1 U13369 ( .A(n17328), .ZN(n18967) );
  AOI22_X1 U13370 ( .A1(\mem[892][3] ), .A2(n17325), .B1(n26238), .B2(
        data_in[3]), .ZN(n17328) );
  INV_X1 U13371 ( .A(n17329), .ZN(n18966) );
  AOI22_X1 U13372 ( .A1(\mem[892][4] ), .A2(n17325), .B1(n26238), .B2(
        data_in[4]), .ZN(n17329) );
  INV_X1 U13373 ( .A(n17330), .ZN(n18965) );
  AOI22_X1 U13374 ( .A1(\mem[892][5] ), .A2(n17325), .B1(n26238), .B2(
        data_in[5]), .ZN(n17330) );
  INV_X1 U13375 ( .A(n17331), .ZN(n18964) );
  AOI22_X1 U13376 ( .A1(\mem[892][6] ), .A2(n17325), .B1(n26238), .B2(
        data_in[6]), .ZN(n17331) );
  INV_X1 U13377 ( .A(n17332), .ZN(n18963) );
  AOI22_X1 U13378 ( .A1(\mem[892][7] ), .A2(n17325), .B1(n26238), .B2(
        data_in[7]), .ZN(n17332) );
  INV_X1 U13379 ( .A(n17333), .ZN(n18962) );
  AOI22_X1 U13380 ( .A1(\mem[893][0] ), .A2(n17334), .B1(n26237), .B2(
        data_in[0]), .ZN(n17333) );
  INV_X1 U13381 ( .A(n17335), .ZN(n18961) );
  AOI22_X1 U13382 ( .A1(\mem[893][1] ), .A2(n17334), .B1(n26237), .B2(
        data_in[1]), .ZN(n17335) );
  INV_X1 U13383 ( .A(n17336), .ZN(n18960) );
  AOI22_X1 U13384 ( .A1(\mem[893][2] ), .A2(n17334), .B1(n26237), .B2(
        data_in[2]), .ZN(n17336) );
  INV_X1 U13385 ( .A(n17337), .ZN(n18959) );
  AOI22_X1 U13386 ( .A1(\mem[893][3] ), .A2(n17334), .B1(n26237), .B2(
        data_in[3]), .ZN(n17337) );
  INV_X1 U13387 ( .A(n17338), .ZN(n18958) );
  AOI22_X1 U13388 ( .A1(\mem[893][4] ), .A2(n17334), .B1(n26237), .B2(
        data_in[4]), .ZN(n17338) );
  INV_X1 U13389 ( .A(n17339), .ZN(n18957) );
  AOI22_X1 U13390 ( .A1(\mem[893][5] ), .A2(n17334), .B1(n26237), .B2(
        data_in[5]), .ZN(n17339) );
  INV_X1 U13391 ( .A(n17340), .ZN(n18956) );
  AOI22_X1 U13392 ( .A1(\mem[893][6] ), .A2(n17334), .B1(n26237), .B2(
        data_in[6]), .ZN(n17340) );
  INV_X1 U13393 ( .A(n17341), .ZN(n18955) );
  AOI22_X1 U13394 ( .A1(\mem[893][7] ), .A2(n17334), .B1(n26237), .B2(
        data_in[7]), .ZN(n17341) );
  INV_X1 U13395 ( .A(n17342), .ZN(n18954) );
  AOI22_X1 U13396 ( .A1(\mem[894][0] ), .A2(n17343), .B1(n26236), .B2(
        data_in[0]), .ZN(n17342) );
  INV_X1 U13397 ( .A(n17344), .ZN(n18953) );
  AOI22_X1 U13398 ( .A1(\mem[894][1] ), .A2(n17343), .B1(n26236), .B2(
        data_in[1]), .ZN(n17344) );
  INV_X1 U13399 ( .A(n17345), .ZN(n18952) );
  AOI22_X1 U13400 ( .A1(\mem[894][2] ), .A2(n17343), .B1(n26236), .B2(
        data_in[2]), .ZN(n17345) );
  INV_X1 U13401 ( .A(n17346), .ZN(n18951) );
  AOI22_X1 U13402 ( .A1(\mem[894][3] ), .A2(n17343), .B1(n26236), .B2(
        data_in[3]), .ZN(n17346) );
  INV_X1 U13403 ( .A(n17347), .ZN(n18950) );
  AOI22_X1 U13404 ( .A1(\mem[894][4] ), .A2(n17343), .B1(n26236), .B2(
        data_in[4]), .ZN(n17347) );
  INV_X1 U13405 ( .A(n17348), .ZN(n18949) );
  AOI22_X1 U13406 ( .A1(\mem[894][5] ), .A2(n17343), .B1(n26236), .B2(
        data_in[5]), .ZN(n17348) );
  INV_X1 U13407 ( .A(n17349), .ZN(n18948) );
  AOI22_X1 U13408 ( .A1(\mem[894][6] ), .A2(n17343), .B1(n26236), .B2(
        data_in[6]), .ZN(n17349) );
  INV_X1 U13409 ( .A(n17350), .ZN(n18947) );
  AOI22_X1 U13410 ( .A1(\mem[894][7] ), .A2(n17343), .B1(n26236), .B2(
        data_in[7]), .ZN(n17350) );
  INV_X1 U13411 ( .A(n17351), .ZN(n18946) );
  AOI22_X1 U13412 ( .A1(\mem[895][0] ), .A2(n17352), .B1(n26235), .B2(
        data_in[0]), .ZN(n17351) );
  INV_X1 U13413 ( .A(n17353), .ZN(n18945) );
  AOI22_X1 U13414 ( .A1(\mem[895][1] ), .A2(n17352), .B1(n26235), .B2(
        data_in[1]), .ZN(n17353) );
  INV_X1 U13415 ( .A(n17354), .ZN(n18944) );
  AOI22_X1 U13416 ( .A1(\mem[895][2] ), .A2(n17352), .B1(n26235), .B2(
        data_in[2]), .ZN(n17354) );
  INV_X1 U13417 ( .A(n17355), .ZN(n18943) );
  AOI22_X1 U13418 ( .A1(\mem[895][3] ), .A2(n17352), .B1(n26235), .B2(
        data_in[3]), .ZN(n17355) );
  INV_X1 U13419 ( .A(n17356), .ZN(n18942) );
  AOI22_X1 U13420 ( .A1(\mem[895][4] ), .A2(n17352), .B1(n26235), .B2(
        data_in[4]), .ZN(n17356) );
  INV_X1 U13421 ( .A(n17357), .ZN(n18941) );
  AOI22_X1 U13422 ( .A1(\mem[895][5] ), .A2(n17352), .B1(n26235), .B2(
        data_in[5]), .ZN(n17357) );
  INV_X1 U13423 ( .A(n17358), .ZN(n18940) );
  AOI22_X1 U13424 ( .A1(\mem[895][6] ), .A2(n17352), .B1(n26235), .B2(
        data_in[6]), .ZN(n17358) );
  INV_X1 U13425 ( .A(n17359), .ZN(n18939) );
  AOI22_X1 U13426 ( .A1(\mem[895][7] ), .A2(n17352), .B1(n26235), .B2(
        data_in[7]), .ZN(n17359) );
  INV_X1 U13427 ( .A(n17433), .ZN(n18874) );
  AOI22_X1 U13428 ( .A1(\mem[904][0] ), .A2(n17434), .B1(n26226), .B2(
        data_in[0]), .ZN(n17433) );
  INV_X1 U13429 ( .A(n17435), .ZN(n18873) );
  AOI22_X1 U13430 ( .A1(\mem[904][1] ), .A2(n17434), .B1(n26226), .B2(
        data_in[1]), .ZN(n17435) );
  INV_X1 U13431 ( .A(n17436), .ZN(n18872) );
  AOI22_X1 U13432 ( .A1(\mem[904][2] ), .A2(n17434), .B1(n26226), .B2(
        data_in[2]), .ZN(n17436) );
  INV_X1 U13433 ( .A(n17437), .ZN(n18871) );
  AOI22_X1 U13434 ( .A1(\mem[904][3] ), .A2(n17434), .B1(n26226), .B2(
        data_in[3]), .ZN(n17437) );
  INV_X1 U13435 ( .A(n17438), .ZN(n18870) );
  AOI22_X1 U13436 ( .A1(\mem[904][4] ), .A2(n17434), .B1(n26226), .B2(
        data_in[4]), .ZN(n17438) );
  INV_X1 U13437 ( .A(n17439), .ZN(n18869) );
  AOI22_X1 U13438 ( .A1(\mem[904][5] ), .A2(n17434), .B1(n26226), .B2(
        data_in[5]), .ZN(n17439) );
  INV_X1 U13439 ( .A(n17440), .ZN(n18868) );
  AOI22_X1 U13440 ( .A1(\mem[904][6] ), .A2(n17434), .B1(n26226), .B2(
        data_in[6]), .ZN(n17440) );
  INV_X1 U13441 ( .A(n17441), .ZN(n18867) );
  AOI22_X1 U13442 ( .A1(\mem[904][7] ), .A2(n17434), .B1(n26226), .B2(
        data_in[7]), .ZN(n17441) );
  INV_X1 U13443 ( .A(n17442), .ZN(n18866) );
  AOI22_X1 U13444 ( .A1(\mem[905][0] ), .A2(n17443), .B1(n26225), .B2(
        data_in[0]), .ZN(n17442) );
  INV_X1 U13445 ( .A(n17444), .ZN(n18865) );
  AOI22_X1 U13446 ( .A1(\mem[905][1] ), .A2(n17443), .B1(n26225), .B2(
        data_in[1]), .ZN(n17444) );
  INV_X1 U13447 ( .A(n17445), .ZN(n18864) );
  AOI22_X1 U13448 ( .A1(\mem[905][2] ), .A2(n17443), .B1(n26225), .B2(
        data_in[2]), .ZN(n17445) );
  INV_X1 U13449 ( .A(n17446), .ZN(n18863) );
  AOI22_X1 U13450 ( .A1(\mem[905][3] ), .A2(n17443), .B1(n26225), .B2(
        data_in[3]), .ZN(n17446) );
  INV_X1 U13451 ( .A(n17447), .ZN(n18862) );
  AOI22_X1 U13452 ( .A1(\mem[905][4] ), .A2(n17443), .B1(n26225), .B2(
        data_in[4]), .ZN(n17447) );
  INV_X1 U13453 ( .A(n17448), .ZN(n18861) );
  AOI22_X1 U13454 ( .A1(\mem[905][5] ), .A2(n17443), .B1(n26225), .B2(
        data_in[5]), .ZN(n17448) );
  INV_X1 U13455 ( .A(n17449), .ZN(n18860) );
  AOI22_X1 U13456 ( .A1(\mem[905][6] ), .A2(n17443), .B1(n26225), .B2(
        data_in[6]), .ZN(n17449) );
  INV_X1 U13457 ( .A(n17450), .ZN(n18859) );
  AOI22_X1 U13458 ( .A1(\mem[905][7] ), .A2(n17443), .B1(n26225), .B2(
        data_in[7]), .ZN(n17450) );
  INV_X1 U13459 ( .A(n17451), .ZN(n18858) );
  AOI22_X1 U13460 ( .A1(\mem[906][0] ), .A2(n17452), .B1(n26224), .B2(
        data_in[0]), .ZN(n17451) );
  INV_X1 U13461 ( .A(n17453), .ZN(n18857) );
  AOI22_X1 U13462 ( .A1(\mem[906][1] ), .A2(n17452), .B1(n26224), .B2(
        data_in[1]), .ZN(n17453) );
  INV_X1 U13463 ( .A(n17454), .ZN(n18856) );
  AOI22_X1 U13464 ( .A1(\mem[906][2] ), .A2(n17452), .B1(n26224), .B2(
        data_in[2]), .ZN(n17454) );
  INV_X1 U13465 ( .A(n17455), .ZN(n18855) );
  AOI22_X1 U13466 ( .A1(\mem[906][3] ), .A2(n17452), .B1(n26224), .B2(
        data_in[3]), .ZN(n17455) );
  INV_X1 U13467 ( .A(n17456), .ZN(n18854) );
  AOI22_X1 U13468 ( .A1(\mem[906][4] ), .A2(n17452), .B1(n26224), .B2(
        data_in[4]), .ZN(n17456) );
  INV_X1 U13469 ( .A(n17457), .ZN(n18853) );
  AOI22_X1 U13470 ( .A1(\mem[906][5] ), .A2(n17452), .B1(n26224), .B2(
        data_in[5]), .ZN(n17457) );
  INV_X1 U13471 ( .A(n17458), .ZN(n18852) );
  AOI22_X1 U13472 ( .A1(\mem[906][6] ), .A2(n17452), .B1(n26224), .B2(
        data_in[6]), .ZN(n17458) );
  INV_X1 U13473 ( .A(n17459), .ZN(n18851) );
  AOI22_X1 U13474 ( .A1(\mem[906][7] ), .A2(n17452), .B1(n26224), .B2(
        data_in[7]), .ZN(n17459) );
  INV_X1 U13475 ( .A(n17460), .ZN(n18850) );
  AOI22_X1 U13476 ( .A1(\mem[907][0] ), .A2(n17461), .B1(n26223), .B2(
        data_in[0]), .ZN(n17460) );
  INV_X1 U13477 ( .A(n17462), .ZN(n18849) );
  AOI22_X1 U13478 ( .A1(\mem[907][1] ), .A2(n17461), .B1(n26223), .B2(
        data_in[1]), .ZN(n17462) );
  INV_X1 U13479 ( .A(n17463), .ZN(n18848) );
  AOI22_X1 U13480 ( .A1(\mem[907][2] ), .A2(n17461), .B1(n26223), .B2(
        data_in[2]), .ZN(n17463) );
  INV_X1 U13481 ( .A(n17464), .ZN(n18847) );
  AOI22_X1 U13482 ( .A1(\mem[907][3] ), .A2(n17461), .B1(n26223), .B2(
        data_in[3]), .ZN(n17464) );
  INV_X1 U13483 ( .A(n17465), .ZN(n18846) );
  AOI22_X1 U13484 ( .A1(\mem[907][4] ), .A2(n17461), .B1(n26223), .B2(
        data_in[4]), .ZN(n17465) );
  INV_X1 U13485 ( .A(n17466), .ZN(n18845) );
  AOI22_X1 U13486 ( .A1(\mem[907][5] ), .A2(n17461), .B1(n26223), .B2(
        data_in[5]), .ZN(n17466) );
  INV_X1 U13487 ( .A(n17467), .ZN(n18844) );
  AOI22_X1 U13488 ( .A1(\mem[907][6] ), .A2(n17461), .B1(n26223), .B2(
        data_in[6]), .ZN(n17467) );
  INV_X1 U13489 ( .A(n17468), .ZN(n18843) );
  AOI22_X1 U13490 ( .A1(\mem[907][7] ), .A2(n17461), .B1(n26223), .B2(
        data_in[7]), .ZN(n17468) );
  INV_X1 U13491 ( .A(n17469), .ZN(n18842) );
  AOI22_X1 U13492 ( .A1(\mem[908][0] ), .A2(n17470), .B1(n26222), .B2(
        data_in[0]), .ZN(n17469) );
  INV_X1 U13493 ( .A(n17471), .ZN(n18841) );
  AOI22_X1 U13494 ( .A1(\mem[908][1] ), .A2(n17470), .B1(n26222), .B2(
        data_in[1]), .ZN(n17471) );
  INV_X1 U13495 ( .A(n17472), .ZN(n18840) );
  AOI22_X1 U13496 ( .A1(\mem[908][2] ), .A2(n17470), .B1(n26222), .B2(
        data_in[2]), .ZN(n17472) );
  INV_X1 U13497 ( .A(n17473), .ZN(n18839) );
  AOI22_X1 U13498 ( .A1(\mem[908][3] ), .A2(n17470), .B1(n26222), .B2(
        data_in[3]), .ZN(n17473) );
  INV_X1 U13499 ( .A(n17474), .ZN(n18838) );
  AOI22_X1 U13500 ( .A1(\mem[908][4] ), .A2(n17470), .B1(n26222), .B2(
        data_in[4]), .ZN(n17474) );
  INV_X1 U13501 ( .A(n17475), .ZN(n18837) );
  AOI22_X1 U13502 ( .A1(\mem[908][5] ), .A2(n17470), .B1(n26222), .B2(
        data_in[5]), .ZN(n17475) );
  INV_X1 U13503 ( .A(n17476), .ZN(n18836) );
  AOI22_X1 U13504 ( .A1(\mem[908][6] ), .A2(n17470), .B1(n26222), .B2(
        data_in[6]), .ZN(n17476) );
  INV_X1 U13505 ( .A(n17477), .ZN(n18835) );
  AOI22_X1 U13506 ( .A1(\mem[908][7] ), .A2(n17470), .B1(n26222), .B2(
        data_in[7]), .ZN(n17477) );
  INV_X1 U13507 ( .A(n17478), .ZN(n18834) );
  AOI22_X1 U13508 ( .A1(\mem[909][0] ), .A2(n17479), .B1(n26221), .B2(
        data_in[0]), .ZN(n17478) );
  INV_X1 U13509 ( .A(n17480), .ZN(n18833) );
  AOI22_X1 U13510 ( .A1(\mem[909][1] ), .A2(n17479), .B1(n26221), .B2(
        data_in[1]), .ZN(n17480) );
  INV_X1 U13511 ( .A(n17481), .ZN(n18832) );
  AOI22_X1 U13512 ( .A1(\mem[909][2] ), .A2(n17479), .B1(n26221), .B2(
        data_in[2]), .ZN(n17481) );
  INV_X1 U13513 ( .A(n17482), .ZN(n18831) );
  AOI22_X1 U13514 ( .A1(\mem[909][3] ), .A2(n17479), .B1(n26221), .B2(
        data_in[3]), .ZN(n17482) );
  INV_X1 U13515 ( .A(n17483), .ZN(n18830) );
  AOI22_X1 U13516 ( .A1(\mem[909][4] ), .A2(n17479), .B1(n26221), .B2(
        data_in[4]), .ZN(n17483) );
  INV_X1 U13517 ( .A(n17484), .ZN(n18829) );
  AOI22_X1 U13518 ( .A1(\mem[909][5] ), .A2(n17479), .B1(n26221), .B2(
        data_in[5]), .ZN(n17484) );
  INV_X1 U13519 ( .A(n17485), .ZN(n18828) );
  AOI22_X1 U13520 ( .A1(\mem[909][6] ), .A2(n17479), .B1(n26221), .B2(
        data_in[6]), .ZN(n17485) );
  INV_X1 U13521 ( .A(n17486), .ZN(n18827) );
  AOI22_X1 U13522 ( .A1(\mem[909][7] ), .A2(n17479), .B1(n26221), .B2(
        data_in[7]), .ZN(n17486) );
  INV_X1 U13523 ( .A(n17487), .ZN(n18826) );
  AOI22_X1 U13524 ( .A1(\mem[910][0] ), .A2(n17488), .B1(n26220), .B2(
        data_in[0]), .ZN(n17487) );
  INV_X1 U13525 ( .A(n17489), .ZN(n18825) );
  AOI22_X1 U13526 ( .A1(\mem[910][1] ), .A2(n17488), .B1(n26220), .B2(
        data_in[1]), .ZN(n17489) );
  INV_X1 U13527 ( .A(n17490), .ZN(n18824) );
  AOI22_X1 U13528 ( .A1(\mem[910][2] ), .A2(n17488), .B1(n26220), .B2(
        data_in[2]), .ZN(n17490) );
  INV_X1 U13529 ( .A(n17491), .ZN(n18823) );
  AOI22_X1 U13530 ( .A1(\mem[910][3] ), .A2(n17488), .B1(n26220), .B2(
        data_in[3]), .ZN(n17491) );
  INV_X1 U13531 ( .A(n17492), .ZN(n18822) );
  AOI22_X1 U13532 ( .A1(\mem[910][4] ), .A2(n17488), .B1(n26220), .B2(
        data_in[4]), .ZN(n17492) );
  INV_X1 U13533 ( .A(n17493), .ZN(n18821) );
  AOI22_X1 U13534 ( .A1(\mem[910][5] ), .A2(n17488), .B1(n26220), .B2(
        data_in[5]), .ZN(n17493) );
  INV_X1 U13535 ( .A(n17494), .ZN(n18820) );
  AOI22_X1 U13536 ( .A1(\mem[910][6] ), .A2(n17488), .B1(n26220), .B2(
        data_in[6]), .ZN(n17494) );
  INV_X1 U13537 ( .A(n17495), .ZN(n18819) );
  AOI22_X1 U13538 ( .A1(\mem[910][7] ), .A2(n17488), .B1(n26220), .B2(
        data_in[7]), .ZN(n17495) );
  INV_X1 U13539 ( .A(n17496), .ZN(n18818) );
  AOI22_X1 U13540 ( .A1(\mem[911][0] ), .A2(n17497), .B1(n26219), .B2(
        data_in[0]), .ZN(n17496) );
  INV_X1 U13541 ( .A(n17498), .ZN(n18817) );
  AOI22_X1 U13542 ( .A1(\mem[911][1] ), .A2(n17497), .B1(n26219), .B2(
        data_in[1]), .ZN(n17498) );
  INV_X1 U13543 ( .A(n17499), .ZN(n18816) );
  AOI22_X1 U13544 ( .A1(\mem[911][2] ), .A2(n17497), .B1(n26219), .B2(
        data_in[2]), .ZN(n17499) );
  INV_X1 U13545 ( .A(n17500), .ZN(n18815) );
  AOI22_X1 U13546 ( .A1(\mem[911][3] ), .A2(n17497), .B1(n26219), .B2(
        data_in[3]), .ZN(n17500) );
  INV_X1 U13547 ( .A(n17501), .ZN(n18814) );
  AOI22_X1 U13548 ( .A1(\mem[911][4] ), .A2(n17497), .B1(n26219), .B2(
        data_in[4]), .ZN(n17501) );
  INV_X1 U13549 ( .A(n17502), .ZN(n18813) );
  AOI22_X1 U13550 ( .A1(\mem[911][5] ), .A2(n17497), .B1(n26219), .B2(
        data_in[5]), .ZN(n17502) );
  INV_X1 U13551 ( .A(n17503), .ZN(n18812) );
  AOI22_X1 U13552 ( .A1(\mem[911][6] ), .A2(n17497), .B1(n26219), .B2(
        data_in[6]), .ZN(n17503) );
  INV_X1 U13553 ( .A(n17504), .ZN(n18811) );
  AOI22_X1 U13554 ( .A1(\mem[911][7] ), .A2(n17497), .B1(n26219), .B2(
        data_in[7]), .ZN(n17504) );
  INV_X1 U13555 ( .A(n17505), .ZN(n18810) );
  AOI22_X1 U13556 ( .A1(\mem[912][0] ), .A2(n17506), .B1(n26218), .B2(
        data_in[0]), .ZN(n17505) );
  INV_X1 U13557 ( .A(n17507), .ZN(n18809) );
  AOI22_X1 U13558 ( .A1(\mem[912][1] ), .A2(n17506), .B1(n26218), .B2(
        data_in[1]), .ZN(n17507) );
  INV_X1 U13559 ( .A(n17508), .ZN(n18808) );
  AOI22_X1 U13560 ( .A1(\mem[912][2] ), .A2(n17506), .B1(n26218), .B2(
        data_in[2]), .ZN(n17508) );
  INV_X1 U13561 ( .A(n17509), .ZN(n18807) );
  AOI22_X1 U13562 ( .A1(\mem[912][3] ), .A2(n17506), .B1(n26218), .B2(
        data_in[3]), .ZN(n17509) );
  INV_X1 U13563 ( .A(n17510), .ZN(n18806) );
  AOI22_X1 U13564 ( .A1(\mem[912][4] ), .A2(n17506), .B1(n26218), .B2(
        data_in[4]), .ZN(n17510) );
  INV_X1 U13565 ( .A(n17511), .ZN(n18805) );
  AOI22_X1 U13566 ( .A1(\mem[912][5] ), .A2(n17506), .B1(n26218), .B2(
        data_in[5]), .ZN(n17511) );
  INV_X1 U13567 ( .A(n17512), .ZN(n18804) );
  AOI22_X1 U13568 ( .A1(\mem[912][6] ), .A2(n17506), .B1(n26218), .B2(
        data_in[6]), .ZN(n17512) );
  INV_X1 U13569 ( .A(n17513), .ZN(n18803) );
  AOI22_X1 U13570 ( .A1(\mem[912][7] ), .A2(n17506), .B1(n26218), .B2(
        data_in[7]), .ZN(n17513) );
  INV_X1 U13571 ( .A(n17514), .ZN(n18802) );
  AOI22_X1 U13572 ( .A1(\mem[913][0] ), .A2(n17515), .B1(n26217), .B2(
        data_in[0]), .ZN(n17514) );
  INV_X1 U13573 ( .A(n17516), .ZN(n18801) );
  AOI22_X1 U13574 ( .A1(\mem[913][1] ), .A2(n17515), .B1(n26217), .B2(
        data_in[1]), .ZN(n17516) );
  INV_X1 U13575 ( .A(n17517), .ZN(n18800) );
  AOI22_X1 U13576 ( .A1(\mem[913][2] ), .A2(n17515), .B1(n26217), .B2(
        data_in[2]), .ZN(n17517) );
  INV_X1 U13577 ( .A(n17518), .ZN(n18799) );
  AOI22_X1 U13578 ( .A1(\mem[913][3] ), .A2(n17515), .B1(n26217), .B2(
        data_in[3]), .ZN(n17518) );
  INV_X1 U13579 ( .A(n17519), .ZN(n18798) );
  AOI22_X1 U13580 ( .A1(\mem[913][4] ), .A2(n17515), .B1(n26217), .B2(
        data_in[4]), .ZN(n17519) );
  INV_X1 U13581 ( .A(n17520), .ZN(n18797) );
  AOI22_X1 U13582 ( .A1(\mem[913][5] ), .A2(n17515), .B1(n26217), .B2(
        data_in[5]), .ZN(n17520) );
  INV_X1 U13583 ( .A(n17521), .ZN(n18796) );
  AOI22_X1 U13584 ( .A1(\mem[913][6] ), .A2(n17515), .B1(n26217), .B2(
        data_in[6]), .ZN(n17521) );
  INV_X1 U13585 ( .A(n17522), .ZN(n18795) );
  AOI22_X1 U13586 ( .A1(\mem[913][7] ), .A2(n17515), .B1(n26217), .B2(
        data_in[7]), .ZN(n17522) );
  INV_X1 U13587 ( .A(n17523), .ZN(n18794) );
  AOI22_X1 U13588 ( .A1(\mem[914][0] ), .A2(n17524), .B1(n26216), .B2(
        data_in[0]), .ZN(n17523) );
  INV_X1 U13589 ( .A(n17525), .ZN(n18793) );
  AOI22_X1 U13590 ( .A1(\mem[914][1] ), .A2(n17524), .B1(n26216), .B2(
        data_in[1]), .ZN(n17525) );
  INV_X1 U13591 ( .A(n17526), .ZN(n18792) );
  AOI22_X1 U13592 ( .A1(\mem[914][2] ), .A2(n17524), .B1(n26216), .B2(
        data_in[2]), .ZN(n17526) );
  INV_X1 U13593 ( .A(n17527), .ZN(n18791) );
  AOI22_X1 U13594 ( .A1(\mem[914][3] ), .A2(n17524), .B1(n26216), .B2(
        data_in[3]), .ZN(n17527) );
  INV_X1 U13595 ( .A(n17528), .ZN(n18790) );
  AOI22_X1 U13596 ( .A1(\mem[914][4] ), .A2(n17524), .B1(n26216), .B2(
        data_in[4]), .ZN(n17528) );
  INV_X1 U13597 ( .A(n17529), .ZN(n18789) );
  AOI22_X1 U13598 ( .A1(\mem[914][5] ), .A2(n17524), .B1(n26216), .B2(
        data_in[5]), .ZN(n17529) );
  INV_X1 U13599 ( .A(n17530), .ZN(n18788) );
  AOI22_X1 U13600 ( .A1(\mem[914][6] ), .A2(n17524), .B1(n26216), .B2(
        data_in[6]), .ZN(n17530) );
  INV_X1 U13601 ( .A(n17531), .ZN(n18787) );
  AOI22_X1 U13602 ( .A1(\mem[914][7] ), .A2(n17524), .B1(n26216), .B2(
        data_in[7]), .ZN(n17531) );
  INV_X1 U13603 ( .A(n17532), .ZN(n18786) );
  AOI22_X1 U13604 ( .A1(\mem[915][0] ), .A2(n17533), .B1(n26215), .B2(
        data_in[0]), .ZN(n17532) );
  INV_X1 U13605 ( .A(n17534), .ZN(n18785) );
  AOI22_X1 U13606 ( .A1(\mem[915][1] ), .A2(n17533), .B1(n26215), .B2(
        data_in[1]), .ZN(n17534) );
  INV_X1 U13607 ( .A(n17535), .ZN(n18784) );
  AOI22_X1 U13608 ( .A1(\mem[915][2] ), .A2(n17533), .B1(n26215), .B2(
        data_in[2]), .ZN(n17535) );
  INV_X1 U13609 ( .A(n17536), .ZN(n18783) );
  AOI22_X1 U13610 ( .A1(\mem[915][3] ), .A2(n17533), .B1(n26215), .B2(
        data_in[3]), .ZN(n17536) );
  INV_X1 U13611 ( .A(n17537), .ZN(n18782) );
  AOI22_X1 U13612 ( .A1(\mem[915][4] ), .A2(n17533), .B1(n26215), .B2(
        data_in[4]), .ZN(n17537) );
  INV_X1 U13613 ( .A(n17538), .ZN(n18781) );
  AOI22_X1 U13614 ( .A1(\mem[915][5] ), .A2(n17533), .B1(n26215), .B2(
        data_in[5]), .ZN(n17538) );
  INV_X1 U13615 ( .A(n17539), .ZN(n18780) );
  AOI22_X1 U13616 ( .A1(\mem[915][6] ), .A2(n17533), .B1(n26215), .B2(
        data_in[6]), .ZN(n17539) );
  INV_X1 U13617 ( .A(n17540), .ZN(n18779) );
  AOI22_X1 U13618 ( .A1(\mem[915][7] ), .A2(n17533), .B1(n26215), .B2(
        data_in[7]), .ZN(n17540) );
  INV_X1 U13619 ( .A(n17541), .ZN(n18778) );
  AOI22_X1 U13620 ( .A1(\mem[916][0] ), .A2(n17542), .B1(n26214), .B2(
        data_in[0]), .ZN(n17541) );
  INV_X1 U13621 ( .A(n17543), .ZN(n18777) );
  AOI22_X1 U13622 ( .A1(\mem[916][1] ), .A2(n17542), .B1(n26214), .B2(
        data_in[1]), .ZN(n17543) );
  INV_X1 U13623 ( .A(n17544), .ZN(n18776) );
  AOI22_X1 U13624 ( .A1(\mem[916][2] ), .A2(n17542), .B1(n26214), .B2(
        data_in[2]), .ZN(n17544) );
  INV_X1 U13625 ( .A(n17545), .ZN(n18775) );
  AOI22_X1 U13626 ( .A1(\mem[916][3] ), .A2(n17542), .B1(n26214), .B2(
        data_in[3]), .ZN(n17545) );
  INV_X1 U13627 ( .A(n17546), .ZN(n18774) );
  AOI22_X1 U13628 ( .A1(\mem[916][4] ), .A2(n17542), .B1(n26214), .B2(
        data_in[4]), .ZN(n17546) );
  INV_X1 U13629 ( .A(n17547), .ZN(n18773) );
  AOI22_X1 U13630 ( .A1(\mem[916][5] ), .A2(n17542), .B1(n26214), .B2(
        data_in[5]), .ZN(n17547) );
  INV_X1 U13631 ( .A(n17548), .ZN(n18772) );
  AOI22_X1 U13632 ( .A1(\mem[916][6] ), .A2(n17542), .B1(n26214), .B2(
        data_in[6]), .ZN(n17548) );
  INV_X1 U13633 ( .A(n17549), .ZN(n18771) );
  AOI22_X1 U13634 ( .A1(\mem[916][7] ), .A2(n17542), .B1(n26214), .B2(
        data_in[7]), .ZN(n17549) );
  INV_X1 U13635 ( .A(n17550), .ZN(n18770) );
  AOI22_X1 U13636 ( .A1(\mem[917][0] ), .A2(n17551), .B1(n26213), .B2(
        data_in[0]), .ZN(n17550) );
  INV_X1 U13637 ( .A(n17552), .ZN(n18769) );
  AOI22_X1 U13638 ( .A1(\mem[917][1] ), .A2(n17551), .B1(n26213), .B2(
        data_in[1]), .ZN(n17552) );
  INV_X1 U13639 ( .A(n17553), .ZN(n18768) );
  AOI22_X1 U13640 ( .A1(\mem[917][2] ), .A2(n17551), .B1(n26213), .B2(
        data_in[2]), .ZN(n17553) );
  INV_X1 U13641 ( .A(n17554), .ZN(n18767) );
  AOI22_X1 U13642 ( .A1(\mem[917][3] ), .A2(n17551), .B1(n26213), .B2(
        data_in[3]), .ZN(n17554) );
  INV_X1 U13643 ( .A(n17555), .ZN(n18766) );
  AOI22_X1 U13644 ( .A1(\mem[917][4] ), .A2(n17551), .B1(n26213), .B2(
        data_in[4]), .ZN(n17555) );
  INV_X1 U13645 ( .A(n17556), .ZN(n18765) );
  AOI22_X1 U13646 ( .A1(\mem[917][5] ), .A2(n17551), .B1(n26213), .B2(
        data_in[5]), .ZN(n17556) );
  INV_X1 U13647 ( .A(n17557), .ZN(n18764) );
  AOI22_X1 U13648 ( .A1(\mem[917][6] ), .A2(n17551), .B1(n26213), .B2(
        data_in[6]), .ZN(n17557) );
  INV_X1 U13649 ( .A(n17558), .ZN(n18763) );
  AOI22_X1 U13650 ( .A1(\mem[917][7] ), .A2(n17551), .B1(n26213), .B2(
        data_in[7]), .ZN(n17558) );
  INV_X1 U13651 ( .A(n17559), .ZN(n18762) );
  AOI22_X1 U13652 ( .A1(\mem[918][0] ), .A2(n17560), .B1(n26212), .B2(
        data_in[0]), .ZN(n17559) );
  INV_X1 U13653 ( .A(n17561), .ZN(n18761) );
  AOI22_X1 U13654 ( .A1(\mem[918][1] ), .A2(n17560), .B1(n26212), .B2(
        data_in[1]), .ZN(n17561) );
  INV_X1 U13655 ( .A(n17562), .ZN(n18760) );
  AOI22_X1 U13656 ( .A1(\mem[918][2] ), .A2(n17560), .B1(n26212), .B2(
        data_in[2]), .ZN(n17562) );
  INV_X1 U13657 ( .A(n17563), .ZN(n18759) );
  AOI22_X1 U13658 ( .A1(\mem[918][3] ), .A2(n17560), .B1(n26212), .B2(
        data_in[3]), .ZN(n17563) );
  INV_X1 U13659 ( .A(n17564), .ZN(n18758) );
  AOI22_X1 U13660 ( .A1(\mem[918][4] ), .A2(n17560), .B1(n26212), .B2(
        data_in[4]), .ZN(n17564) );
  INV_X1 U13661 ( .A(n17565), .ZN(n18757) );
  AOI22_X1 U13662 ( .A1(\mem[918][5] ), .A2(n17560), .B1(n26212), .B2(
        data_in[5]), .ZN(n17565) );
  INV_X1 U13663 ( .A(n17566), .ZN(n18756) );
  AOI22_X1 U13664 ( .A1(\mem[918][6] ), .A2(n17560), .B1(n26212), .B2(
        data_in[6]), .ZN(n17566) );
  INV_X1 U13665 ( .A(n17567), .ZN(n18755) );
  AOI22_X1 U13666 ( .A1(\mem[918][7] ), .A2(n17560), .B1(n26212), .B2(
        data_in[7]), .ZN(n17567) );
  INV_X1 U13667 ( .A(n17568), .ZN(n18754) );
  AOI22_X1 U13668 ( .A1(\mem[919][0] ), .A2(n17569), .B1(n26211), .B2(
        data_in[0]), .ZN(n17568) );
  INV_X1 U13669 ( .A(n17570), .ZN(n18753) );
  AOI22_X1 U13670 ( .A1(\mem[919][1] ), .A2(n17569), .B1(n26211), .B2(
        data_in[1]), .ZN(n17570) );
  INV_X1 U13671 ( .A(n17571), .ZN(n18752) );
  AOI22_X1 U13672 ( .A1(\mem[919][2] ), .A2(n17569), .B1(n26211), .B2(
        data_in[2]), .ZN(n17571) );
  INV_X1 U13673 ( .A(n17572), .ZN(n18751) );
  AOI22_X1 U13674 ( .A1(\mem[919][3] ), .A2(n17569), .B1(n26211), .B2(
        data_in[3]), .ZN(n17572) );
  INV_X1 U13675 ( .A(n17573), .ZN(n18750) );
  AOI22_X1 U13676 ( .A1(\mem[919][4] ), .A2(n17569), .B1(n26211), .B2(
        data_in[4]), .ZN(n17573) );
  INV_X1 U13677 ( .A(n17574), .ZN(n18749) );
  AOI22_X1 U13678 ( .A1(\mem[919][5] ), .A2(n17569), .B1(n26211), .B2(
        data_in[5]), .ZN(n17574) );
  INV_X1 U13679 ( .A(n17575), .ZN(n18748) );
  AOI22_X1 U13680 ( .A1(\mem[919][6] ), .A2(n17569), .B1(n26211), .B2(
        data_in[6]), .ZN(n17575) );
  INV_X1 U13681 ( .A(n17576), .ZN(n18747) );
  AOI22_X1 U13682 ( .A1(\mem[919][7] ), .A2(n17569), .B1(n26211), .B2(
        data_in[7]), .ZN(n17576) );
  INV_X1 U13683 ( .A(n17577), .ZN(n18746) );
  AOI22_X1 U13684 ( .A1(\mem[920][0] ), .A2(n17578), .B1(n26210), .B2(
        data_in[0]), .ZN(n17577) );
  INV_X1 U13685 ( .A(n17579), .ZN(n18745) );
  AOI22_X1 U13686 ( .A1(\mem[920][1] ), .A2(n17578), .B1(n26210), .B2(
        data_in[1]), .ZN(n17579) );
  INV_X1 U13687 ( .A(n17580), .ZN(n18744) );
  AOI22_X1 U13688 ( .A1(\mem[920][2] ), .A2(n17578), .B1(n26210), .B2(
        data_in[2]), .ZN(n17580) );
  INV_X1 U13689 ( .A(n17581), .ZN(n18743) );
  AOI22_X1 U13690 ( .A1(\mem[920][3] ), .A2(n17578), .B1(n26210), .B2(
        data_in[3]), .ZN(n17581) );
  INV_X1 U13691 ( .A(n17582), .ZN(n18742) );
  AOI22_X1 U13692 ( .A1(\mem[920][4] ), .A2(n17578), .B1(n26210), .B2(
        data_in[4]), .ZN(n17582) );
  INV_X1 U13693 ( .A(n17583), .ZN(n18741) );
  AOI22_X1 U13694 ( .A1(\mem[920][5] ), .A2(n17578), .B1(n26210), .B2(
        data_in[5]), .ZN(n17583) );
  INV_X1 U13695 ( .A(n17584), .ZN(n18740) );
  AOI22_X1 U13696 ( .A1(\mem[920][6] ), .A2(n17578), .B1(n26210), .B2(
        data_in[6]), .ZN(n17584) );
  INV_X1 U13697 ( .A(n17585), .ZN(n18739) );
  AOI22_X1 U13698 ( .A1(\mem[920][7] ), .A2(n17578), .B1(n26210), .B2(
        data_in[7]), .ZN(n17585) );
  INV_X1 U13699 ( .A(n17586), .ZN(n18738) );
  AOI22_X1 U13700 ( .A1(\mem[921][0] ), .A2(n17587), .B1(n26209), .B2(
        data_in[0]), .ZN(n17586) );
  INV_X1 U13701 ( .A(n17588), .ZN(n18737) );
  AOI22_X1 U13702 ( .A1(\mem[921][1] ), .A2(n17587), .B1(n26209), .B2(
        data_in[1]), .ZN(n17588) );
  INV_X1 U13703 ( .A(n17589), .ZN(n18736) );
  AOI22_X1 U13704 ( .A1(\mem[921][2] ), .A2(n17587), .B1(n26209), .B2(
        data_in[2]), .ZN(n17589) );
  INV_X1 U13705 ( .A(n17590), .ZN(n18735) );
  AOI22_X1 U13706 ( .A1(\mem[921][3] ), .A2(n17587), .B1(n26209), .B2(
        data_in[3]), .ZN(n17590) );
  INV_X1 U13707 ( .A(n17591), .ZN(n18734) );
  AOI22_X1 U13708 ( .A1(\mem[921][4] ), .A2(n17587), .B1(n26209), .B2(
        data_in[4]), .ZN(n17591) );
  INV_X1 U13709 ( .A(n17592), .ZN(n18733) );
  AOI22_X1 U13710 ( .A1(\mem[921][5] ), .A2(n17587), .B1(n26209), .B2(
        data_in[5]), .ZN(n17592) );
  INV_X1 U13711 ( .A(n17593), .ZN(n18732) );
  AOI22_X1 U13712 ( .A1(\mem[921][6] ), .A2(n17587), .B1(n26209), .B2(
        data_in[6]), .ZN(n17593) );
  INV_X1 U13713 ( .A(n17594), .ZN(n18731) );
  AOI22_X1 U13714 ( .A1(\mem[921][7] ), .A2(n17587), .B1(n26209), .B2(
        data_in[7]), .ZN(n17594) );
  INV_X1 U13715 ( .A(n17595), .ZN(n18730) );
  AOI22_X1 U13716 ( .A1(\mem[922][0] ), .A2(n17596), .B1(n26208), .B2(
        data_in[0]), .ZN(n17595) );
  INV_X1 U13717 ( .A(n17597), .ZN(n18729) );
  AOI22_X1 U13718 ( .A1(\mem[922][1] ), .A2(n17596), .B1(n26208), .B2(
        data_in[1]), .ZN(n17597) );
  INV_X1 U13719 ( .A(n17598), .ZN(n18728) );
  AOI22_X1 U13720 ( .A1(\mem[922][2] ), .A2(n17596), .B1(n26208), .B2(
        data_in[2]), .ZN(n17598) );
  INV_X1 U13721 ( .A(n17599), .ZN(n18727) );
  AOI22_X1 U13722 ( .A1(\mem[922][3] ), .A2(n17596), .B1(n26208), .B2(
        data_in[3]), .ZN(n17599) );
  INV_X1 U13723 ( .A(n17600), .ZN(n18726) );
  AOI22_X1 U13724 ( .A1(\mem[922][4] ), .A2(n17596), .B1(n26208), .B2(
        data_in[4]), .ZN(n17600) );
  INV_X1 U13725 ( .A(n17601), .ZN(n18725) );
  AOI22_X1 U13726 ( .A1(\mem[922][5] ), .A2(n17596), .B1(n26208), .B2(
        data_in[5]), .ZN(n17601) );
  INV_X1 U13727 ( .A(n17602), .ZN(n18724) );
  AOI22_X1 U13728 ( .A1(\mem[922][6] ), .A2(n17596), .B1(n26208), .B2(
        data_in[6]), .ZN(n17602) );
  INV_X1 U13729 ( .A(n17603), .ZN(n18723) );
  AOI22_X1 U13730 ( .A1(\mem[922][7] ), .A2(n17596), .B1(n26208), .B2(
        data_in[7]), .ZN(n17603) );
  INV_X1 U13731 ( .A(n17604), .ZN(n18722) );
  AOI22_X1 U13732 ( .A1(\mem[923][0] ), .A2(n17605), .B1(n26207), .B2(
        data_in[0]), .ZN(n17604) );
  INV_X1 U13733 ( .A(n17606), .ZN(n18721) );
  AOI22_X1 U13734 ( .A1(\mem[923][1] ), .A2(n17605), .B1(n26207), .B2(
        data_in[1]), .ZN(n17606) );
  INV_X1 U13735 ( .A(n17607), .ZN(n18720) );
  AOI22_X1 U13736 ( .A1(\mem[923][2] ), .A2(n17605), .B1(n26207), .B2(
        data_in[2]), .ZN(n17607) );
  INV_X1 U13737 ( .A(n17608), .ZN(n18719) );
  AOI22_X1 U13738 ( .A1(\mem[923][3] ), .A2(n17605), .B1(n26207), .B2(
        data_in[3]), .ZN(n17608) );
  INV_X1 U13739 ( .A(n17609), .ZN(n18718) );
  AOI22_X1 U13740 ( .A1(\mem[923][4] ), .A2(n17605), .B1(n26207), .B2(
        data_in[4]), .ZN(n17609) );
  INV_X1 U13741 ( .A(n17610), .ZN(n18717) );
  AOI22_X1 U13742 ( .A1(\mem[923][5] ), .A2(n17605), .B1(n26207), .B2(
        data_in[5]), .ZN(n17610) );
  INV_X1 U13743 ( .A(n17611), .ZN(n18716) );
  AOI22_X1 U13744 ( .A1(\mem[923][6] ), .A2(n17605), .B1(n26207), .B2(
        data_in[6]), .ZN(n17611) );
  INV_X1 U13745 ( .A(n17612), .ZN(n18715) );
  AOI22_X1 U13746 ( .A1(\mem[923][7] ), .A2(n17605), .B1(n26207), .B2(
        data_in[7]), .ZN(n17612) );
  INV_X1 U13747 ( .A(n17613), .ZN(n18714) );
  AOI22_X1 U13748 ( .A1(\mem[924][0] ), .A2(n17614), .B1(n26206), .B2(
        data_in[0]), .ZN(n17613) );
  INV_X1 U13749 ( .A(n17615), .ZN(n18713) );
  AOI22_X1 U13750 ( .A1(\mem[924][1] ), .A2(n17614), .B1(n26206), .B2(
        data_in[1]), .ZN(n17615) );
  INV_X1 U13751 ( .A(n17616), .ZN(n18712) );
  AOI22_X1 U13752 ( .A1(\mem[924][2] ), .A2(n17614), .B1(n26206), .B2(
        data_in[2]), .ZN(n17616) );
  INV_X1 U13753 ( .A(n17617), .ZN(n18711) );
  AOI22_X1 U13754 ( .A1(\mem[924][3] ), .A2(n17614), .B1(n26206), .B2(
        data_in[3]), .ZN(n17617) );
  INV_X1 U13755 ( .A(n17618), .ZN(n18710) );
  AOI22_X1 U13756 ( .A1(\mem[924][4] ), .A2(n17614), .B1(n26206), .B2(
        data_in[4]), .ZN(n17618) );
  INV_X1 U13757 ( .A(n17619), .ZN(n18709) );
  AOI22_X1 U13758 ( .A1(\mem[924][5] ), .A2(n17614), .B1(n26206), .B2(
        data_in[5]), .ZN(n17619) );
  INV_X1 U13759 ( .A(n17620), .ZN(n18708) );
  AOI22_X1 U13760 ( .A1(\mem[924][6] ), .A2(n17614), .B1(n26206), .B2(
        data_in[6]), .ZN(n17620) );
  INV_X1 U13761 ( .A(n17621), .ZN(n18707) );
  AOI22_X1 U13762 ( .A1(\mem[924][7] ), .A2(n17614), .B1(n26206), .B2(
        data_in[7]), .ZN(n17621) );
  INV_X1 U13763 ( .A(n17622), .ZN(n18706) );
  AOI22_X1 U13764 ( .A1(\mem[925][0] ), .A2(n17623), .B1(n26205), .B2(
        data_in[0]), .ZN(n17622) );
  INV_X1 U13765 ( .A(n17624), .ZN(n18705) );
  AOI22_X1 U13766 ( .A1(\mem[925][1] ), .A2(n17623), .B1(n26205), .B2(
        data_in[1]), .ZN(n17624) );
  INV_X1 U13767 ( .A(n17625), .ZN(n18704) );
  AOI22_X1 U13768 ( .A1(\mem[925][2] ), .A2(n17623), .B1(n26205), .B2(
        data_in[2]), .ZN(n17625) );
  INV_X1 U13769 ( .A(n17626), .ZN(n18703) );
  AOI22_X1 U13770 ( .A1(\mem[925][3] ), .A2(n17623), .B1(n26205), .B2(
        data_in[3]), .ZN(n17626) );
  INV_X1 U13771 ( .A(n17627), .ZN(n18702) );
  AOI22_X1 U13772 ( .A1(\mem[925][4] ), .A2(n17623), .B1(n26205), .B2(
        data_in[4]), .ZN(n17627) );
  INV_X1 U13773 ( .A(n17628), .ZN(n18701) );
  AOI22_X1 U13774 ( .A1(\mem[925][5] ), .A2(n17623), .B1(n26205), .B2(
        data_in[5]), .ZN(n17628) );
  INV_X1 U13775 ( .A(n17629), .ZN(n18700) );
  AOI22_X1 U13776 ( .A1(\mem[925][6] ), .A2(n17623), .B1(n26205), .B2(
        data_in[6]), .ZN(n17629) );
  INV_X1 U13777 ( .A(n17630), .ZN(n18699) );
  AOI22_X1 U13778 ( .A1(\mem[925][7] ), .A2(n17623), .B1(n26205), .B2(
        data_in[7]), .ZN(n17630) );
  INV_X1 U13779 ( .A(n17631), .ZN(n18698) );
  AOI22_X1 U13780 ( .A1(\mem[926][0] ), .A2(n17632), .B1(n26204), .B2(
        data_in[0]), .ZN(n17631) );
  INV_X1 U13781 ( .A(n17633), .ZN(n18697) );
  AOI22_X1 U13782 ( .A1(\mem[926][1] ), .A2(n17632), .B1(n26204), .B2(
        data_in[1]), .ZN(n17633) );
  INV_X1 U13783 ( .A(n17634), .ZN(n18696) );
  AOI22_X1 U13784 ( .A1(\mem[926][2] ), .A2(n17632), .B1(n26204), .B2(
        data_in[2]), .ZN(n17634) );
  INV_X1 U13785 ( .A(n17635), .ZN(n18695) );
  AOI22_X1 U13786 ( .A1(\mem[926][3] ), .A2(n17632), .B1(n26204), .B2(
        data_in[3]), .ZN(n17635) );
  INV_X1 U13787 ( .A(n17636), .ZN(n18694) );
  AOI22_X1 U13788 ( .A1(\mem[926][4] ), .A2(n17632), .B1(n26204), .B2(
        data_in[4]), .ZN(n17636) );
  INV_X1 U13789 ( .A(n17637), .ZN(n18693) );
  AOI22_X1 U13790 ( .A1(\mem[926][5] ), .A2(n17632), .B1(n26204), .B2(
        data_in[5]), .ZN(n17637) );
  INV_X1 U13791 ( .A(n17638), .ZN(n18692) );
  AOI22_X1 U13792 ( .A1(\mem[926][6] ), .A2(n17632), .B1(n26204), .B2(
        data_in[6]), .ZN(n17638) );
  INV_X1 U13793 ( .A(n17639), .ZN(n18691) );
  AOI22_X1 U13794 ( .A1(\mem[926][7] ), .A2(n17632), .B1(n26204), .B2(
        data_in[7]), .ZN(n17639) );
  INV_X1 U13795 ( .A(n17640), .ZN(n18690) );
  AOI22_X1 U13796 ( .A1(\mem[927][0] ), .A2(n17641), .B1(n26203), .B2(
        data_in[0]), .ZN(n17640) );
  INV_X1 U13797 ( .A(n17642), .ZN(n18689) );
  AOI22_X1 U13798 ( .A1(\mem[927][1] ), .A2(n17641), .B1(n26203), .B2(
        data_in[1]), .ZN(n17642) );
  INV_X1 U13799 ( .A(n17643), .ZN(n18688) );
  AOI22_X1 U13800 ( .A1(\mem[927][2] ), .A2(n17641), .B1(n26203), .B2(
        data_in[2]), .ZN(n17643) );
  INV_X1 U13801 ( .A(n17644), .ZN(n18687) );
  AOI22_X1 U13802 ( .A1(\mem[927][3] ), .A2(n17641), .B1(n26203), .B2(
        data_in[3]), .ZN(n17644) );
  INV_X1 U13803 ( .A(n17645), .ZN(n18686) );
  AOI22_X1 U13804 ( .A1(\mem[927][4] ), .A2(n17641), .B1(n26203), .B2(
        data_in[4]), .ZN(n17645) );
  INV_X1 U13805 ( .A(n17646), .ZN(n18685) );
  AOI22_X1 U13806 ( .A1(\mem[927][5] ), .A2(n17641), .B1(n26203), .B2(
        data_in[5]), .ZN(n17646) );
  INV_X1 U13807 ( .A(n17647), .ZN(n18684) );
  AOI22_X1 U13808 ( .A1(\mem[927][6] ), .A2(n17641), .B1(n26203), .B2(
        data_in[6]), .ZN(n17647) );
  INV_X1 U13809 ( .A(n17648), .ZN(n18683) );
  AOI22_X1 U13810 ( .A1(\mem[927][7] ), .A2(n17641), .B1(n26203), .B2(
        data_in[7]), .ZN(n17648) );
  INV_X1 U13811 ( .A(n17722), .ZN(n18618) );
  AOI22_X1 U13812 ( .A1(\mem[936][0] ), .A2(n17723), .B1(n26194), .B2(
        data_in[0]), .ZN(n17722) );
  INV_X1 U13813 ( .A(n17724), .ZN(n18617) );
  AOI22_X1 U13814 ( .A1(\mem[936][1] ), .A2(n17723), .B1(n26194), .B2(
        data_in[1]), .ZN(n17724) );
  INV_X1 U13815 ( .A(n17725), .ZN(n18616) );
  AOI22_X1 U13816 ( .A1(\mem[936][2] ), .A2(n17723), .B1(n26194), .B2(
        data_in[2]), .ZN(n17725) );
  INV_X1 U13817 ( .A(n17726), .ZN(n18615) );
  AOI22_X1 U13818 ( .A1(\mem[936][3] ), .A2(n17723), .B1(n26194), .B2(
        data_in[3]), .ZN(n17726) );
  INV_X1 U13819 ( .A(n17727), .ZN(n18614) );
  AOI22_X1 U13820 ( .A1(\mem[936][4] ), .A2(n17723), .B1(n26194), .B2(
        data_in[4]), .ZN(n17727) );
  INV_X1 U13821 ( .A(n17728), .ZN(n18613) );
  AOI22_X1 U13822 ( .A1(\mem[936][5] ), .A2(n17723), .B1(n26194), .B2(
        data_in[5]), .ZN(n17728) );
  INV_X1 U13823 ( .A(n17729), .ZN(n18612) );
  AOI22_X1 U13824 ( .A1(\mem[936][6] ), .A2(n17723), .B1(n26194), .B2(
        data_in[6]), .ZN(n17729) );
  INV_X1 U13825 ( .A(n17730), .ZN(n18611) );
  AOI22_X1 U13826 ( .A1(\mem[936][7] ), .A2(n17723), .B1(n26194), .B2(
        data_in[7]), .ZN(n17730) );
  INV_X1 U13827 ( .A(n17731), .ZN(n18610) );
  AOI22_X1 U13828 ( .A1(\mem[937][0] ), .A2(n17732), .B1(n26193), .B2(
        data_in[0]), .ZN(n17731) );
  INV_X1 U13829 ( .A(n17733), .ZN(n18609) );
  AOI22_X1 U13830 ( .A1(\mem[937][1] ), .A2(n17732), .B1(n26193), .B2(
        data_in[1]), .ZN(n17733) );
  INV_X1 U13831 ( .A(n17734), .ZN(n18608) );
  AOI22_X1 U13832 ( .A1(\mem[937][2] ), .A2(n17732), .B1(n26193), .B2(
        data_in[2]), .ZN(n17734) );
  INV_X1 U13833 ( .A(n17735), .ZN(n18607) );
  AOI22_X1 U13834 ( .A1(\mem[937][3] ), .A2(n17732), .B1(n26193), .B2(
        data_in[3]), .ZN(n17735) );
  INV_X1 U13835 ( .A(n17736), .ZN(n18606) );
  AOI22_X1 U13836 ( .A1(\mem[937][4] ), .A2(n17732), .B1(n26193), .B2(
        data_in[4]), .ZN(n17736) );
  INV_X1 U13837 ( .A(n17737), .ZN(n18605) );
  AOI22_X1 U13838 ( .A1(\mem[937][5] ), .A2(n17732), .B1(n26193), .B2(
        data_in[5]), .ZN(n17737) );
  INV_X1 U13839 ( .A(n17738), .ZN(n18604) );
  AOI22_X1 U13840 ( .A1(\mem[937][6] ), .A2(n17732), .B1(n26193), .B2(
        data_in[6]), .ZN(n17738) );
  INV_X1 U13841 ( .A(n17739), .ZN(n18603) );
  AOI22_X1 U13842 ( .A1(\mem[937][7] ), .A2(n17732), .B1(n26193), .B2(
        data_in[7]), .ZN(n17739) );
  INV_X1 U13843 ( .A(n17740), .ZN(n18602) );
  AOI22_X1 U13844 ( .A1(\mem[938][0] ), .A2(n17741), .B1(n26192), .B2(
        data_in[0]), .ZN(n17740) );
  INV_X1 U13845 ( .A(n17742), .ZN(n18601) );
  AOI22_X1 U13846 ( .A1(\mem[938][1] ), .A2(n17741), .B1(n26192), .B2(
        data_in[1]), .ZN(n17742) );
  INV_X1 U13847 ( .A(n17743), .ZN(n18600) );
  AOI22_X1 U13848 ( .A1(\mem[938][2] ), .A2(n17741), .B1(n26192), .B2(
        data_in[2]), .ZN(n17743) );
  INV_X1 U13849 ( .A(n17744), .ZN(n18599) );
  AOI22_X1 U13850 ( .A1(\mem[938][3] ), .A2(n17741), .B1(n26192), .B2(
        data_in[3]), .ZN(n17744) );
  INV_X1 U13851 ( .A(n17745), .ZN(n18598) );
  AOI22_X1 U13852 ( .A1(\mem[938][4] ), .A2(n17741), .B1(n26192), .B2(
        data_in[4]), .ZN(n17745) );
  INV_X1 U13853 ( .A(n17746), .ZN(n18597) );
  AOI22_X1 U13854 ( .A1(\mem[938][5] ), .A2(n17741), .B1(n26192), .B2(
        data_in[5]), .ZN(n17746) );
  INV_X1 U13855 ( .A(n17747), .ZN(n18596) );
  AOI22_X1 U13856 ( .A1(\mem[938][6] ), .A2(n17741), .B1(n26192), .B2(
        data_in[6]), .ZN(n17747) );
  INV_X1 U13857 ( .A(n17748), .ZN(n18595) );
  AOI22_X1 U13858 ( .A1(\mem[938][7] ), .A2(n17741), .B1(n26192), .B2(
        data_in[7]), .ZN(n17748) );
  INV_X1 U13859 ( .A(n17749), .ZN(n18594) );
  AOI22_X1 U13860 ( .A1(\mem[939][0] ), .A2(n17750), .B1(n26191), .B2(
        data_in[0]), .ZN(n17749) );
  INV_X1 U13861 ( .A(n17751), .ZN(n18593) );
  AOI22_X1 U13862 ( .A1(\mem[939][1] ), .A2(n17750), .B1(n26191), .B2(
        data_in[1]), .ZN(n17751) );
  INV_X1 U13863 ( .A(n17752), .ZN(n18592) );
  AOI22_X1 U13864 ( .A1(\mem[939][2] ), .A2(n17750), .B1(n26191), .B2(
        data_in[2]), .ZN(n17752) );
  INV_X1 U13865 ( .A(n17753), .ZN(n18591) );
  AOI22_X1 U13866 ( .A1(\mem[939][3] ), .A2(n17750), .B1(n26191), .B2(
        data_in[3]), .ZN(n17753) );
  INV_X1 U13867 ( .A(n17754), .ZN(n18590) );
  AOI22_X1 U13868 ( .A1(\mem[939][4] ), .A2(n17750), .B1(n26191), .B2(
        data_in[4]), .ZN(n17754) );
  INV_X1 U13869 ( .A(n17755), .ZN(n18589) );
  AOI22_X1 U13870 ( .A1(\mem[939][5] ), .A2(n17750), .B1(n26191), .B2(
        data_in[5]), .ZN(n17755) );
  INV_X1 U13871 ( .A(n17756), .ZN(n18588) );
  AOI22_X1 U13872 ( .A1(\mem[939][6] ), .A2(n17750), .B1(n26191), .B2(
        data_in[6]), .ZN(n17756) );
  INV_X1 U13873 ( .A(n17757), .ZN(n18587) );
  AOI22_X1 U13874 ( .A1(\mem[939][7] ), .A2(n17750), .B1(n26191), .B2(
        data_in[7]), .ZN(n17757) );
  INV_X1 U13875 ( .A(n17758), .ZN(n18586) );
  AOI22_X1 U13876 ( .A1(\mem[940][0] ), .A2(n17759), .B1(n26190), .B2(
        data_in[0]), .ZN(n17758) );
  INV_X1 U13877 ( .A(n17760), .ZN(n18585) );
  AOI22_X1 U13878 ( .A1(\mem[940][1] ), .A2(n17759), .B1(n26190), .B2(
        data_in[1]), .ZN(n17760) );
  INV_X1 U13879 ( .A(n17761), .ZN(n18584) );
  AOI22_X1 U13880 ( .A1(\mem[940][2] ), .A2(n17759), .B1(n26190), .B2(
        data_in[2]), .ZN(n17761) );
  INV_X1 U13881 ( .A(n17762), .ZN(n18583) );
  AOI22_X1 U13882 ( .A1(\mem[940][3] ), .A2(n17759), .B1(n26190), .B2(
        data_in[3]), .ZN(n17762) );
  INV_X1 U13883 ( .A(n17763), .ZN(n18582) );
  AOI22_X1 U13884 ( .A1(\mem[940][4] ), .A2(n17759), .B1(n26190), .B2(
        data_in[4]), .ZN(n17763) );
  INV_X1 U13885 ( .A(n17764), .ZN(n18581) );
  AOI22_X1 U13886 ( .A1(\mem[940][5] ), .A2(n17759), .B1(n26190), .B2(
        data_in[5]), .ZN(n17764) );
  INV_X1 U13887 ( .A(n17765), .ZN(n18580) );
  AOI22_X1 U13888 ( .A1(\mem[940][6] ), .A2(n17759), .B1(n26190), .B2(
        data_in[6]), .ZN(n17765) );
  INV_X1 U13889 ( .A(n17766), .ZN(n18579) );
  AOI22_X1 U13890 ( .A1(\mem[940][7] ), .A2(n17759), .B1(n26190), .B2(
        data_in[7]), .ZN(n17766) );
  INV_X1 U13891 ( .A(n17767), .ZN(n18578) );
  AOI22_X1 U13892 ( .A1(\mem[941][0] ), .A2(n17768), .B1(n26189), .B2(
        data_in[0]), .ZN(n17767) );
  INV_X1 U13893 ( .A(n17769), .ZN(n18577) );
  AOI22_X1 U13894 ( .A1(\mem[941][1] ), .A2(n17768), .B1(n26189), .B2(
        data_in[1]), .ZN(n17769) );
  INV_X1 U13895 ( .A(n17770), .ZN(n18576) );
  AOI22_X1 U13896 ( .A1(\mem[941][2] ), .A2(n17768), .B1(n26189), .B2(
        data_in[2]), .ZN(n17770) );
  INV_X1 U13897 ( .A(n17771), .ZN(n18575) );
  AOI22_X1 U13898 ( .A1(\mem[941][3] ), .A2(n17768), .B1(n26189), .B2(
        data_in[3]), .ZN(n17771) );
  INV_X1 U13899 ( .A(n17772), .ZN(n18574) );
  AOI22_X1 U13900 ( .A1(\mem[941][4] ), .A2(n17768), .B1(n26189), .B2(
        data_in[4]), .ZN(n17772) );
  INV_X1 U13901 ( .A(n17773), .ZN(n18573) );
  AOI22_X1 U13902 ( .A1(\mem[941][5] ), .A2(n17768), .B1(n26189), .B2(
        data_in[5]), .ZN(n17773) );
  INV_X1 U13903 ( .A(n17774), .ZN(n18572) );
  AOI22_X1 U13904 ( .A1(\mem[941][6] ), .A2(n17768), .B1(n26189), .B2(
        data_in[6]), .ZN(n17774) );
  INV_X1 U13905 ( .A(n17775), .ZN(n18571) );
  AOI22_X1 U13906 ( .A1(\mem[941][7] ), .A2(n17768), .B1(n26189), .B2(
        data_in[7]), .ZN(n17775) );
  INV_X1 U13907 ( .A(n17776), .ZN(n18570) );
  AOI22_X1 U13908 ( .A1(\mem[942][0] ), .A2(n17777), .B1(n26188), .B2(
        data_in[0]), .ZN(n17776) );
  INV_X1 U13909 ( .A(n17778), .ZN(n18569) );
  AOI22_X1 U13910 ( .A1(\mem[942][1] ), .A2(n17777), .B1(n26188), .B2(
        data_in[1]), .ZN(n17778) );
  INV_X1 U13911 ( .A(n17779), .ZN(n18568) );
  AOI22_X1 U13912 ( .A1(\mem[942][2] ), .A2(n17777), .B1(n26188), .B2(
        data_in[2]), .ZN(n17779) );
  INV_X1 U13913 ( .A(n17780), .ZN(n18567) );
  AOI22_X1 U13914 ( .A1(\mem[942][3] ), .A2(n17777), .B1(n26188), .B2(
        data_in[3]), .ZN(n17780) );
  INV_X1 U13915 ( .A(n17781), .ZN(n18566) );
  AOI22_X1 U13916 ( .A1(\mem[942][4] ), .A2(n17777), .B1(n26188), .B2(
        data_in[4]), .ZN(n17781) );
  INV_X1 U13917 ( .A(n17782), .ZN(n18565) );
  AOI22_X1 U13918 ( .A1(\mem[942][5] ), .A2(n17777), .B1(n26188), .B2(
        data_in[5]), .ZN(n17782) );
  INV_X1 U13919 ( .A(n17783), .ZN(n18564) );
  AOI22_X1 U13920 ( .A1(\mem[942][6] ), .A2(n17777), .B1(n26188), .B2(
        data_in[6]), .ZN(n17783) );
  INV_X1 U13921 ( .A(n17784), .ZN(n18563) );
  AOI22_X1 U13922 ( .A1(\mem[942][7] ), .A2(n17777), .B1(n26188), .B2(
        data_in[7]), .ZN(n17784) );
  INV_X1 U13923 ( .A(n17785), .ZN(n18562) );
  AOI22_X1 U13924 ( .A1(\mem[943][0] ), .A2(n17786), .B1(n26187), .B2(
        data_in[0]), .ZN(n17785) );
  INV_X1 U13925 ( .A(n17787), .ZN(n18561) );
  AOI22_X1 U13926 ( .A1(\mem[943][1] ), .A2(n17786), .B1(n26187), .B2(
        data_in[1]), .ZN(n17787) );
  INV_X1 U13927 ( .A(n17788), .ZN(n18560) );
  AOI22_X1 U13928 ( .A1(\mem[943][2] ), .A2(n17786), .B1(n26187), .B2(
        data_in[2]), .ZN(n17788) );
  INV_X1 U13929 ( .A(n17789), .ZN(n18559) );
  AOI22_X1 U13930 ( .A1(\mem[943][3] ), .A2(n17786), .B1(n26187), .B2(
        data_in[3]), .ZN(n17789) );
  INV_X1 U13931 ( .A(n17790), .ZN(n18558) );
  AOI22_X1 U13932 ( .A1(\mem[943][4] ), .A2(n17786), .B1(n26187), .B2(
        data_in[4]), .ZN(n17790) );
  INV_X1 U13933 ( .A(n17791), .ZN(n18557) );
  AOI22_X1 U13934 ( .A1(\mem[943][5] ), .A2(n17786), .B1(n26187), .B2(
        data_in[5]), .ZN(n17791) );
  INV_X1 U13935 ( .A(n17792), .ZN(n18556) );
  AOI22_X1 U13936 ( .A1(\mem[943][6] ), .A2(n17786), .B1(n26187), .B2(
        data_in[6]), .ZN(n17792) );
  INV_X1 U13937 ( .A(n17793), .ZN(n18555) );
  AOI22_X1 U13938 ( .A1(\mem[943][7] ), .A2(n17786), .B1(n26187), .B2(
        data_in[7]), .ZN(n17793) );
  INV_X1 U13939 ( .A(n17794), .ZN(n18554) );
  AOI22_X1 U13940 ( .A1(\mem[944][0] ), .A2(n17795), .B1(n26186), .B2(
        data_in[0]), .ZN(n17794) );
  INV_X1 U13941 ( .A(n17796), .ZN(n18553) );
  AOI22_X1 U13942 ( .A1(\mem[944][1] ), .A2(n17795), .B1(n26186), .B2(
        data_in[1]), .ZN(n17796) );
  INV_X1 U13943 ( .A(n17797), .ZN(n18552) );
  AOI22_X1 U13944 ( .A1(\mem[944][2] ), .A2(n17795), .B1(n26186), .B2(
        data_in[2]), .ZN(n17797) );
  INV_X1 U13945 ( .A(n17798), .ZN(n18551) );
  AOI22_X1 U13946 ( .A1(\mem[944][3] ), .A2(n17795), .B1(n26186), .B2(
        data_in[3]), .ZN(n17798) );
  INV_X1 U13947 ( .A(n17799), .ZN(n18550) );
  AOI22_X1 U13948 ( .A1(\mem[944][4] ), .A2(n17795), .B1(n26186), .B2(
        data_in[4]), .ZN(n17799) );
  INV_X1 U13949 ( .A(n17800), .ZN(n18549) );
  AOI22_X1 U13950 ( .A1(\mem[944][5] ), .A2(n17795), .B1(n26186), .B2(
        data_in[5]), .ZN(n17800) );
  INV_X1 U13951 ( .A(n17801), .ZN(n18548) );
  AOI22_X1 U13952 ( .A1(\mem[944][6] ), .A2(n17795), .B1(n26186), .B2(
        data_in[6]), .ZN(n17801) );
  INV_X1 U13953 ( .A(n17802), .ZN(n18547) );
  AOI22_X1 U13954 ( .A1(\mem[944][7] ), .A2(n17795), .B1(n26186), .B2(
        data_in[7]), .ZN(n17802) );
  INV_X1 U13955 ( .A(n17803), .ZN(n18546) );
  AOI22_X1 U13956 ( .A1(\mem[945][0] ), .A2(n17804), .B1(n26185), .B2(
        data_in[0]), .ZN(n17803) );
  INV_X1 U13957 ( .A(n17805), .ZN(n18545) );
  AOI22_X1 U13958 ( .A1(\mem[945][1] ), .A2(n17804), .B1(n26185), .B2(
        data_in[1]), .ZN(n17805) );
  INV_X1 U13959 ( .A(n17806), .ZN(n18544) );
  AOI22_X1 U13960 ( .A1(\mem[945][2] ), .A2(n17804), .B1(n26185), .B2(
        data_in[2]), .ZN(n17806) );
  INV_X1 U13961 ( .A(n17807), .ZN(n18543) );
  AOI22_X1 U13962 ( .A1(\mem[945][3] ), .A2(n17804), .B1(n26185), .B2(
        data_in[3]), .ZN(n17807) );
  INV_X1 U13963 ( .A(n17808), .ZN(n18542) );
  AOI22_X1 U13964 ( .A1(\mem[945][4] ), .A2(n17804), .B1(n26185), .B2(
        data_in[4]), .ZN(n17808) );
  INV_X1 U13965 ( .A(n17809), .ZN(n18541) );
  AOI22_X1 U13966 ( .A1(\mem[945][5] ), .A2(n17804), .B1(n26185), .B2(
        data_in[5]), .ZN(n17809) );
  INV_X1 U13967 ( .A(n17810), .ZN(n18540) );
  AOI22_X1 U13968 ( .A1(\mem[945][6] ), .A2(n17804), .B1(n26185), .B2(
        data_in[6]), .ZN(n17810) );
  INV_X1 U13969 ( .A(n17811), .ZN(n18539) );
  AOI22_X1 U13970 ( .A1(\mem[945][7] ), .A2(n17804), .B1(n26185), .B2(
        data_in[7]), .ZN(n17811) );
  INV_X1 U13971 ( .A(n17812), .ZN(n18538) );
  AOI22_X1 U13972 ( .A1(\mem[946][0] ), .A2(n17813), .B1(n26184), .B2(
        data_in[0]), .ZN(n17812) );
  INV_X1 U13973 ( .A(n17814), .ZN(n18537) );
  AOI22_X1 U13974 ( .A1(\mem[946][1] ), .A2(n17813), .B1(n26184), .B2(
        data_in[1]), .ZN(n17814) );
  INV_X1 U13975 ( .A(n17815), .ZN(n18536) );
  AOI22_X1 U13976 ( .A1(\mem[946][2] ), .A2(n17813), .B1(n26184), .B2(
        data_in[2]), .ZN(n17815) );
  INV_X1 U13977 ( .A(n17816), .ZN(n18535) );
  AOI22_X1 U13978 ( .A1(\mem[946][3] ), .A2(n17813), .B1(n26184), .B2(
        data_in[3]), .ZN(n17816) );
  INV_X1 U13979 ( .A(n17817), .ZN(n18534) );
  AOI22_X1 U13980 ( .A1(\mem[946][4] ), .A2(n17813), .B1(n26184), .B2(
        data_in[4]), .ZN(n17817) );
  INV_X1 U13981 ( .A(n17818), .ZN(n18533) );
  AOI22_X1 U13982 ( .A1(\mem[946][5] ), .A2(n17813), .B1(n26184), .B2(
        data_in[5]), .ZN(n17818) );
  INV_X1 U13983 ( .A(n17819), .ZN(n18532) );
  AOI22_X1 U13984 ( .A1(\mem[946][6] ), .A2(n17813), .B1(n26184), .B2(
        data_in[6]), .ZN(n17819) );
  INV_X1 U13985 ( .A(n17820), .ZN(n18531) );
  AOI22_X1 U13986 ( .A1(\mem[946][7] ), .A2(n17813), .B1(n26184), .B2(
        data_in[7]), .ZN(n17820) );
  INV_X1 U13987 ( .A(n17821), .ZN(n18530) );
  AOI22_X1 U13988 ( .A1(\mem[947][0] ), .A2(n17822), .B1(n26183), .B2(
        data_in[0]), .ZN(n17821) );
  INV_X1 U13989 ( .A(n17823), .ZN(n18529) );
  AOI22_X1 U13990 ( .A1(\mem[947][1] ), .A2(n17822), .B1(n26183), .B2(
        data_in[1]), .ZN(n17823) );
  INV_X1 U13991 ( .A(n17824), .ZN(n9222) );
  AOI22_X1 U13992 ( .A1(\mem[947][2] ), .A2(n17822), .B1(n26183), .B2(
        data_in[2]), .ZN(n17824) );
  INV_X1 U13993 ( .A(n17825), .ZN(n9221) );
  AOI22_X1 U13994 ( .A1(\mem[947][3] ), .A2(n17822), .B1(n26183), .B2(
        data_in[3]), .ZN(n17825) );
  INV_X1 U13995 ( .A(n17826), .ZN(n9220) );
  AOI22_X1 U13996 ( .A1(\mem[947][4] ), .A2(n17822), .B1(n26183), .B2(
        data_in[4]), .ZN(n17826) );
  INV_X1 U13997 ( .A(n17827), .ZN(n9219) );
  AOI22_X1 U13998 ( .A1(\mem[947][5] ), .A2(n17822), .B1(n26183), .B2(
        data_in[5]), .ZN(n17827) );
  INV_X1 U13999 ( .A(n17828), .ZN(n9218) );
  AOI22_X1 U14000 ( .A1(\mem[947][6] ), .A2(n17822), .B1(n26183), .B2(
        data_in[6]), .ZN(n17828) );
  INV_X1 U14001 ( .A(n17829), .ZN(n9217) );
  AOI22_X1 U14002 ( .A1(\mem[947][7] ), .A2(n17822), .B1(n26183), .B2(
        data_in[7]), .ZN(n17829) );
  INV_X1 U14003 ( .A(n17830), .ZN(n9216) );
  AOI22_X1 U14004 ( .A1(\mem[948][0] ), .A2(n17831), .B1(n26182), .B2(
        data_in[0]), .ZN(n17830) );
  INV_X1 U14005 ( .A(n17832), .ZN(n9215) );
  AOI22_X1 U14006 ( .A1(\mem[948][1] ), .A2(n17831), .B1(n26182), .B2(
        data_in[1]), .ZN(n17832) );
  INV_X1 U14007 ( .A(n17833), .ZN(n9214) );
  AOI22_X1 U14008 ( .A1(\mem[948][2] ), .A2(n17831), .B1(n26182), .B2(
        data_in[2]), .ZN(n17833) );
  INV_X1 U14009 ( .A(n17834), .ZN(n9213) );
  AOI22_X1 U14010 ( .A1(\mem[948][3] ), .A2(n17831), .B1(n26182), .B2(
        data_in[3]), .ZN(n17834) );
  INV_X1 U14011 ( .A(n17835), .ZN(n9212) );
  AOI22_X1 U14012 ( .A1(\mem[948][4] ), .A2(n17831), .B1(n26182), .B2(
        data_in[4]), .ZN(n17835) );
  INV_X1 U14013 ( .A(n17836), .ZN(n9211) );
  AOI22_X1 U14014 ( .A1(\mem[948][5] ), .A2(n17831), .B1(n26182), .B2(
        data_in[5]), .ZN(n17836) );
  INV_X1 U14015 ( .A(n17837), .ZN(n9210) );
  AOI22_X1 U14016 ( .A1(\mem[948][6] ), .A2(n17831), .B1(n26182), .B2(
        data_in[6]), .ZN(n17837) );
  INV_X1 U14017 ( .A(n17838), .ZN(n9209) );
  AOI22_X1 U14018 ( .A1(\mem[948][7] ), .A2(n17831), .B1(n26182), .B2(
        data_in[7]), .ZN(n17838) );
  INV_X1 U14019 ( .A(n17839), .ZN(n9208) );
  AOI22_X1 U14020 ( .A1(\mem[949][0] ), .A2(n17840), .B1(n26181), .B2(
        data_in[0]), .ZN(n17839) );
  INV_X1 U14021 ( .A(n17841), .ZN(n9207) );
  AOI22_X1 U14022 ( .A1(\mem[949][1] ), .A2(n17840), .B1(n26181), .B2(
        data_in[1]), .ZN(n17841) );
  INV_X1 U14023 ( .A(n17842), .ZN(n9206) );
  AOI22_X1 U14024 ( .A1(\mem[949][2] ), .A2(n17840), .B1(n26181), .B2(
        data_in[2]), .ZN(n17842) );
  INV_X1 U14025 ( .A(n17843), .ZN(n9205) );
  AOI22_X1 U14026 ( .A1(\mem[949][3] ), .A2(n17840), .B1(n26181), .B2(
        data_in[3]), .ZN(n17843) );
  INV_X1 U14027 ( .A(n17844), .ZN(n9204) );
  AOI22_X1 U14028 ( .A1(\mem[949][4] ), .A2(n17840), .B1(n26181), .B2(
        data_in[4]), .ZN(n17844) );
  INV_X1 U14029 ( .A(n17845), .ZN(n9203) );
  AOI22_X1 U14030 ( .A1(\mem[949][5] ), .A2(n17840), .B1(n26181), .B2(
        data_in[5]), .ZN(n17845) );
  INV_X1 U14031 ( .A(n17846), .ZN(n9202) );
  AOI22_X1 U14032 ( .A1(\mem[949][6] ), .A2(n17840), .B1(n26181), .B2(
        data_in[6]), .ZN(n17846) );
  INV_X1 U14033 ( .A(n17847), .ZN(n9201) );
  AOI22_X1 U14034 ( .A1(\mem[949][7] ), .A2(n17840), .B1(n26181), .B2(
        data_in[7]), .ZN(n17847) );
  INV_X1 U14035 ( .A(n17848), .ZN(n9200) );
  AOI22_X1 U14036 ( .A1(\mem[950][0] ), .A2(n17849), .B1(n26180), .B2(
        data_in[0]), .ZN(n17848) );
  INV_X1 U14037 ( .A(n17850), .ZN(n9199) );
  AOI22_X1 U14038 ( .A1(\mem[950][1] ), .A2(n17849), .B1(n26180), .B2(
        data_in[1]), .ZN(n17850) );
  INV_X1 U14039 ( .A(n17851), .ZN(n9198) );
  AOI22_X1 U14040 ( .A1(\mem[950][2] ), .A2(n17849), .B1(n26180), .B2(
        data_in[2]), .ZN(n17851) );
  INV_X1 U14041 ( .A(n17852), .ZN(n9197) );
  AOI22_X1 U14042 ( .A1(\mem[950][3] ), .A2(n17849), .B1(n26180), .B2(
        data_in[3]), .ZN(n17852) );
  INV_X1 U14043 ( .A(n17853), .ZN(n9196) );
  AOI22_X1 U14044 ( .A1(\mem[950][4] ), .A2(n17849), .B1(n26180), .B2(
        data_in[4]), .ZN(n17853) );
  INV_X1 U14045 ( .A(n17854), .ZN(n9195) );
  AOI22_X1 U14046 ( .A1(\mem[950][5] ), .A2(n17849), .B1(n26180), .B2(
        data_in[5]), .ZN(n17854) );
  INV_X1 U14047 ( .A(n17855), .ZN(n9194) );
  AOI22_X1 U14048 ( .A1(\mem[950][6] ), .A2(n17849), .B1(n26180), .B2(
        data_in[6]), .ZN(n17855) );
  INV_X1 U14049 ( .A(n17856), .ZN(n9193) );
  AOI22_X1 U14050 ( .A1(\mem[950][7] ), .A2(n17849), .B1(n26180), .B2(
        data_in[7]), .ZN(n17856) );
  INV_X1 U14051 ( .A(n17857), .ZN(n9192) );
  AOI22_X1 U14052 ( .A1(\mem[951][0] ), .A2(n17858), .B1(n26179), .B2(
        data_in[0]), .ZN(n17857) );
  INV_X1 U14053 ( .A(n17859), .ZN(n9191) );
  AOI22_X1 U14054 ( .A1(\mem[951][1] ), .A2(n17858), .B1(n26179), .B2(
        data_in[1]), .ZN(n17859) );
  INV_X1 U14055 ( .A(n17860), .ZN(n9190) );
  AOI22_X1 U14056 ( .A1(\mem[951][2] ), .A2(n17858), .B1(n26179), .B2(
        data_in[2]), .ZN(n17860) );
  INV_X1 U14057 ( .A(n17861), .ZN(n9189) );
  AOI22_X1 U14058 ( .A1(\mem[951][3] ), .A2(n17858), .B1(n26179), .B2(
        data_in[3]), .ZN(n17861) );
  INV_X1 U14059 ( .A(n17862), .ZN(n9188) );
  AOI22_X1 U14060 ( .A1(\mem[951][4] ), .A2(n17858), .B1(n26179), .B2(
        data_in[4]), .ZN(n17862) );
  INV_X1 U14061 ( .A(n17863), .ZN(n9187) );
  AOI22_X1 U14062 ( .A1(\mem[951][5] ), .A2(n17858), .B1(n26179), .B2(
        data_in[5]), .ZN(n17863) );
  INV_X1 U14063 ( .A(n17864), .ZN(n9186) );
  AOI22_X1 U14064 ( .A1(\mem[951][6] ), .A2(n17858), .B1(n26179), .B2(
        data_in[6]), .ZN(n17864) );
  INV_X1 U14065 ( .A(n17865), .ZN(n9185) );
  AOI22_X1 U14066 ( .A1(\mem[951][7] ), .A2(n17858), .B1(n26179), .B2(
        data_in[7]), .ZN(n17865) );
  INV_X1 U14067 ( .A(n17866), .ZN(n9184) );
  AOI22_X1 U14068 ( .A1(\mem[952][0] ), .A2(n17867), .B1(n26178), .B2(
        data_in[0]), .ZN(n17866) );
  INV_X1 U14069 ( .A(n17868), .ZN(n9183) );
  AOI22_X1 U14070 ( .A1(\mem[952][1] ), .A2(n17867), .B1(n26178), .B2(
        data_in[1]), .ZN(n17868) );
  INV_X1 U14071 ( .A(n17869), .ZN(n9182) );
  AOI22_X1 U14072 ( .A1(\mem[952][2] ), .A2(n17867), .B1(n26178), .B2(
        data_in[2]), .ZN(n17869) );
  INV_X1 U14073 ( .A(n17870), .ZN(n9181) );
  AOI22_X1 U14074 ( .A1(\mem[952][3] ), .A2(n17867), .B1(n26178), .B2(
        data_in[3]), .ZN(n17870) );
  INV_X1 U14075 ( .A(n17871), .ZN(n9180) );
  AOI22_X1 U14076 ( .A1(\mem[952][4] ), .A2(n17867), .B1(n26178), .B2(
        data_in[4]), .ZN(n17871) );
  INV_X1 U14077 ( .A(n17872), .ZN(n9179) );
  AOI22_X1 U14078 ( .A1(\mem[952][5] ), .A2(n17867), .B1(n26178), .B2(
        data_in[5]), .ZN(n17872) );
  INV_X1 U14079 ( .A(n17873), .ZN(n9178) );
  AOI22_X1 U14080 ( .A1(\mem[952][6] ), .A2(n17867), .B1(n26178), .B2(
        data_in[6]), .ZN(n17873) );
  INV_X1 U14081 ( .A(n17874), .ZN(n9177) );
  AOI22_X1 U14082 ( .A1(\mem[952][7] ), .A2(n17867), .B1(n26178), .B2(
        data_in[7]), .ZN(n17874) );
  INV_X1 U14083 ( .A(n17875), .ZN(n9176) );
  AOI22_X1 U14084 ( .A1(\mem[953][0] ), .A2(n17876), .B1(n26177), .B2(
        data_in[0]), .ZN(n17875) );
  INV_X1 U14085 ( .A(n17877), .ZN(n9175) );
  AOI22_X1 U14086 ( .A1(\mem[953][1] ), .A2(n17876), .B1(n26177), .B2(
        data_in[1]), .ZN(n17877) );
  INV_X1 U14087 ( .A(n17878), .ZN(n9174) );
  AOI22_X1 U14088 ( .A1(\mem[953][2] ), .A2(n17876), .B1(n26177), .B2(
        data_in[2]), .ZN(n17878) );
  INV_X1 U14089 ( .A(n17879), .ZN(n9173) );
  AOI22_X1 U14090 ( .A1(\mem[953][3] ), .A2(n17876), .B1(n26177), .B2(
        data_in[3]), .ZN(n17879) );
  INV_X1 U14091 ( .A(n17880), .ZN(n9172) );
  AOI22_X1 U14092 ( .A1(\mem[953][4] ), .A2(n17876), .B1(n26177), .B2(
        data_in[4]), .ZN(n17880) );
  INV_X1 U14093 ( .A(n17881), .ZN(n9171) );
  AOI22_X1 U14094 ( .A1(\mem[953][5] ), .A2(n17876), .B1(n26177), .B2(
        data_in[5]), .ZN(n17881) );
  INV_X1 U14095 ( .A(n17882), .ZN(n9170) );
  AOI22_X1 U14096 ( .A1(\mem[953][6] ), .A2(n17876), .B1(n26177), .B2(
        data_in[6]), .ZN(n17882) );
  INV_X1 U14097 ( .A(n17883), .ZN(n9169) );
  AOI22_X1 U14098 ( .A1(\mem[953][7] ), .A2(n17876), .B1(n26177), .B2(
        data_in[7]), .ZN(n17883) );
  INV_X1 U14099 ( .A(n17884), .ZN(n9168) );
  AOI22_X1 U14100 ( .A1(\mem[954][0] ), .A2(n17885), .B1(n26176), .B2(
        data_in[0]), .ZN(n17884) );
  INV_X1 U14101 ( .A(n17886), .ZN(n9167) );
  AOI22_X1 U14102 ( .A1(\mem[954][1] ), .A2(n17885), .B1(n26176), .B2(
        data_in[1]), .ZN(n17886) );
  INV_X1 U14103 ( .A(n17887), .ZN(n9166) );
  AOI22_X1 U14104 ( .A1(\mem[954][2] ), .A2(n17885), .B1(n26176), .B2(
        data_in[2]), .ZN(n17887) );
  INV_X1 U14105 ( .A(n17888), .ZN(n9165) );
  AOI22_X1 U14106 ( .A1(\mem[954][3] ), .A2(n17885), .B1(n26176), .B2(
        data_in[3]), .ZN(n17888) );
  INV_X1 U14107 ( .A(n17889), .ZN(n9164) );
  AOI22_X1 U14108 ( .A1(\mem[954][4] ), .A2(n17885), .B1(n26176), .B2(
        data_in[4]), .ZN(n17889) );
  INV_X1 U14109 ( .A(n17890), .ZN(n9163) );
  AOI22_X1 U14110 ( .A1(\mem[954][5] ), .A2(n17885), .B1(n26176), .B2(
        data_in[5]), .ZN(n17890) );
  INV_X1 U14111 ( .A(n17891), .ZN(n9162) );
  AOI22_X1 U14112 ( .A1(\mem[954][6] ), .A2(n17885), .B1(n26176), .B2(
        data_in[6]), .ZN(n17891) );
  INV_X1 U14113 ( .A(n17892), .ZN(n9161) );
  AOI22_X1 U14114 ( .A1(\mem[954][7] ), .A2(n17885), .B1(n26176), .B2(
        data_in[7]), .ZN(n17892) );
  INV_X1 U14115 ( .A(n17893), .ZN(n9160) );
  AOI22_X1 U14116 ( .A1(\mem[955][0] ), .A2(n17894), .B1(n26175), .B2(
        data_in[0]), .ZN(n17893) );
  INV_X1 U14117 ( .A(n17895), .ZN(n9159) );
  AOI22_X1 U14118 ( .A1(\mem[955][1] ), .A2(n17894), .B1(n26175), .B2(
        data_in[1]), .ZN(n17895) );
  INV_X1 U14119 ( .A(n17896), .ZN(n9158) );
  AOI22_X1 U14120 ( .A1(\mem[955][2] ), .A2(n17894), .B1(n26175), .B2(
        data_in[2]), .ZN(n17896) );
  INV_X1 U14121 ( .A(n17897), .ZN(n9157) );
  AOI22_X1 U14122 ( .A1(\mem[955][3] ), .A2(n17894), .B1(n26175), .B2(
        data_in[3]), .ZN(n17897) );
  INV_X1 U14123 ( .A(n17898), .ZN(n9156) );
  AOI22_X1 U14124 ( .A1(\mem[955][4] ), .A2(n17894), .B1(n26175), .B2(
        data_in[4]), .ZN(n17898) );
  INV_X1 U14125 ( .A(n17899), .ZN(n9155) );
  AOI22_X1 U14126 ( .A1(\mem[955][5] ), .A2(n17894), .B1(n26175), .B2(
        data_in[5]), .ZN(n17899) );
  INV_X1 U14127 ( .A(n17900), .ZN(n9154) );
  AOI22_X1 U14128 ( .A1(\mem[955][6] ), .A2(n17894), .B1(n26175), .B2(
        data_in[6]), .ZN(n17900) );
  INV_X1 U14129 ( .A(n17901), .ZN(n9153) );
  AOI22_X1 U14130 ( .A1(\mem[955][7] ), .A2(n17894), .B1(n26175), .B2(
        data_in[7]), .ZN(n17901) );
  INV_X1 U14131 ( .A(n17902), .ZN(n9152) );
  AOI22_X1 U14132 ( .A1(\mem[956][0] ), .A2(n17903), .B1(n26174), .B2(
        data_in[0]), .ZN(n17902) );
  INV_X1 U14133 ( .A(n17904), .ZN(n9151) );
  AOI22_X1 U14134 ( .A1(\mem[956][1] ), .A2(n17903), .B1(n26174), .B2(
        data_in[1]), .ZN(n17904) );
  INV_X1 U14135 ( .A(n17905), .ZN(n9150) );
  AOI22_X1 U14136 ( .A1(\mem[956][2] ), .A2(n17903), .B1(n26174), .B2(
        data_in[2]), .ZN(n17905) );
  INV_X1 U14137 ( .A(n17906), .ZN(n9149) );
  AOI22_X1 U14138 ( .A1(\mem[956][3] ), .A2(n17903), .B1(n26174), .B2(
        data_in[3]), .ZN(n17906) );
  INV_X1 U14139 ( .A(n17907), .ZN(n9148) );
  AOI22_X1 U14140 ( .A1(\mem[956][4] ), .A2(n17903), .B1(n26174), .B2(
        data_in[4]), .ZN(n17907) );
  INV_X1 U14141 ( .A(n17908), .ZN(n9147) );
  AOI22_X1 U14142 ( .A1(\mem[956][5] ), .A2(n17903), .B1(n26174), .B2(
        data_in[5]), .ZN(n17908) );
  INV_X1 U14143 ( .A(n17909), .ZN(n9146) );
  AOI22_X1 U14144 ( .A1(\mem[956][6] ), .A2(n17903), .B1(n26174), .B2(
        data_in[6]), .ZN(n17909) );
  INV_X1 U14145 ( .A(n17910), .ZN(n9145) );
  AOI22_X1 U14146 ( .A1(\mem[956][7] ), .A2(n17903), .B1(n26174), .B2(
        data_in[7]), .ZN(n17910) );
  INV_X1 U14147 ( .A(n17911), .ZN(n9144) );
  AOI22_X1 U14148 ( .A1(\mem[957][0] ), .A2(n17912), .B1(n26173), .B2(
        data_in[0]), .ZN(n17911) );
  INV_X1 U14149 ( .A(n17913), .ZN(n9143) );
  AOI22_X1 U14150 ( .A1(\mem[957][1] ), .A2(n17912), .B1(n26173), .B2(
        data_in[1]), .ZN(n17913) );
  INV_X1 U14151 ( .A(n17914), .ZN(n9142) );
  AOI22_X1 U14152 ( .A1(\mem[957][2] ), .A2(n17912), .B1(n26173), .B2(
        data_in[2]), .ZN(n17914) );
  INV_X1 U14153 ( .A(n17915), .ZN(n9141) );
  AOI22_X1 U14154 ( .A1(\mem[957][3] ), .A2(n17912), .B1(n26173), .B2(
        data_in[3]), .ZN(n17915) );
  INV_X1 U14155 ( .A(n17916), .ZN(n9140) );
  AOI22_X1 U14156 ( .A1(\mem[957][4] ), .A2(n17912), .B1(n26173), .B2(
        data_in[4]), .ZN(n17916) );
  INV_X1 U14157 ( .A(n17917), .ZN(n9139) );
  AOI22_X1 U14158 ( .A1(\mem[957][5] ), .A2(n17912), .B1(n26173), .B2(
        data_in[5]), .ZN(n17917) );
  INV_X1 U14159 ( .A(n17918), .ZN(n9138) );
  AOI22_X1 U14160 ( .A1(\mem[957][6] ), .A2(n17912), .B1(n26173), .B2(
        data_in[6]), .ZN(n17918) );
  INV_X1 U14161 ( .A(n17919), .ZN(n9137) );
  AOI22_X1 U14162 ( .A1(\mem[957][7] ), .A2(n17912), .B1(n26173), .B2(
        data_in[7]), .ZN(n17919) );
  INV_X1 U14163 ( .A(n17920), .ZN(n9136) );
  AOI22_X1 U14164 ( .A1(\mem[958][0] ), .A2(n17921), .B1(n26172), .B2(
        data_in[0]), .ZN(n17920) );
  INV_X1 U14165 ( .A(n17922), .ZN(n9135) );
  AOI22_X1 U14166 ( .A1(\mem[958][1] ), .A2(n17921), .B1(n26172), .B2(
        data_in[1]), .ZN(n17922) );
  INV_X1 U14167 ( .A(n17923), .ZN(n9134) );
  AOI22_X1 U14168 ( .A1(\mem[958][2] ), .A2(n17921), .B1(n26172), .B2(
        data_in[2]), .ZN(n17923) );
  INV_X1 U14169 ( .A(n17924), .ZN(n9133) );
  AOI22_X1 U14170 ( .A1(\mem[958][3] ), .A2(n17921), .B1(n26172), .B2(
        data_in[3]), .ZN(n17924) );
  INV_X1 U14171 ( .A(n17925), .ZN(n9132) );
  AOI22_X1 U14172 ( .A1(\mem[958][4] ), .A2(n17921), .B1(n26172), .B2(
        data_in[4]), .ZN(n17925) );
  INV_X1 U14173 ( .A(n17926), .ZN(n9131) );
  AOI22_X1 U14174 ( .A1(\mem[958][5] ), .A2(n17921), .B1(n26172), .B2(
        data_in[5]), .ZN(n17926) );
  INV_X1 U14175 ( .A(n17927), .ZN(n9130) );
  AOI22_X1 U14176 ( .A1(\mem[958][6] ), .A2(n17921), .B1(n26172), .B2(
        data_in[6]), .ZN(n17927) );
  INV_X1 U14177 ( .A(n17928), .ZN(n9129) );
  AOI22_X1 U14178 ( .A1(\mem[958][7] ), .A2(n17921), .B1(n26172), .B2(
        data_in[7]), .ZN(n17928) );
  INV_X1 U14179 ( .A(n17929), .ZN(n9128) );
  AOI22_X1 U14180 ( .A1(\mem[959][0] ), .A2(n17930), .B1(n26171), .B2(
        data_in[0]), .ZN(n17929) );
  INV_X1 U14181 ( .A(n17931), .ZN(n9127) );
  AOI22_X1 U14182 ( .A1(\mem[959][1] ), .A2(n17930), .B1(n26171), .B2(
        data_in[1]), .ZN(n17931) );
  INV_X1 U14183 ( .A(n17932), .ZN(n9126) );
  AOI22_X1 U14184 ( .A1(\mem[959][2] ), .A2(n17930), .B1(n26171), .B2(
        data_in[2]), .ZN(n17932) );
  INV_X1 U14185 ( .A(n17933), .ZN(n9125) );
  AOI22_X1 U14186 ( .A1(\mem[959][3] ), .A2(n17930), .B1(n26171), .B2(
        data_in[3]), .ZN(n17933) );
  INV_X1 U14187 ( .A(n17934), .ZN(n9124) );
  AOI22_X1 U14188 ( .A1(\mem[959][4] ), .A2(n17930), .B1(n26171), .B2(
        data_in[4]), .ZN(n17934) );
  INV_X1 U14189 ( .A(n17935), .ZN(n9123) );
  AOI22_X1 U14190 ( .A1(\mem[959][5] ), .A2(n17930), .B1(n26171), .B2(
        data_in[5]), .ZN(n17935) );
  INV_X1 U14191 ( .A(n17936), .ZN(n9122) );
  AOI22_X1 U14192 ( .A1(\mem[959][6] ), .A2(n17930), .B1(n26171), .B2(
        data_in[6]), .ZN(n17936) );
  INV_X1 U14193 ( .A(n17937), .ZN(n9121) );
  AOI22_X1 U14194 ( .A1(\mem[959][7] ), .A2(n17930), .B1(n26171), .B2(
        data_in[7]), .ZN(n17937) );
  INV_X1 U14195 ( .A(n18011), .ZN(n9056) );
  AOI22_X1 U14196 ( .A1(\mem[968][0] ), .A2(n18012), .B1(n26162), .B2(
        data_in[0]), .ZN(n18011) );
  INV_X1 U14197 ( .A(n18013), .ZN(n9055) );
  AOI22_X1 U14198 ( .A1(\mem[968][1] ), .A2(n18012), .B1(n26162), .B2(
        data_in[1]), .ZN(n18013) );
  INV_X1 U14199 ( .A(n18014), .ZN(n9054) );
  AOI22_X1 U14200 ( .A1(\mem[968][2] ), .A2(n18012), .B1(n26162), .B2(
        data_in[2]), .ZN(n18014) );
  INV_X1 U14201 ( .A(n18015), .ZN(n9053) );
  AOI22_X1 U14202 ( .A1(\mem[968][3] ), .A2(n18012), .B1(n26162), .B2(
        data_in[3]), .ZN(n18015) );
  INV_X1 U14203 ( .A(n18016), .ZN(n9052) );
  AOI22_X1 U14204 ( .A1(\mem[968][4] ), .A2(n18012), .B1(n26162), .B2(
        data_in[4]), .ZN(n18016) );
  INV_X1 U14205 ( .A(n18017), .ZN(n9051) );
  AOI22_X1 U14206 ( .A1(\mem[968][5] ), .A2(n18012), .B1(n26162), .B2(
        data_in[5]), .ZN(n18017) );
  INV_X1 U14207 ( .A(n18018), .ZN(n9050) );
  AOI22_X1 U14208 ( .A1(\mem[968][6] ), .A2(n18012), .B1(n26162), .B2(
        data_in[6]), .ZN(n18018) );
  INV_X1 U14209 ( .A(n18019), .ZN(n9049) );
  AOI22_X1 U14210 ( .A1(\mem[968][7] ), .A2(n18012), .B1(n26162), .B2(
        data_in[7]), .ZN(n18019) );
  INV_X1 U14211 ( .A(n18020), .ZN(n9048) );
  AOI22_X1 U14212 ( .A1(\mem[969][0] ), .A2(n18021), .B1(n26161), .B2(
        data_in[0]), .ZN(n18020) );
  INV_X1 U14213 ( .A(n18022), .ZN(n9047) );
  AOI22_X1 U14214 ( .A1(\mem[969][1] ), .A2(n18021), .B1(n26161), .B2(
        data_in[1]), .ZN(n18022) );
  INV_X1 U14215 ( .A(n18023), .ZN(n9046) );
  AOI22_X1 U14216 ( .A1(\mem[969][2] ), .A2(n18021), .B1(n26161), .B2(
        data_in[2]), .ZN(n18023) );
  INV_X1 U14217 ( .A(n18024), .ZN(n9045) );
  AOI22_X1 U14218 ( .A1(\mem[969][3] ), .A2(n18021), .B1(n26161), .B2(
        data_in[3]), .ZN(n18024) );
  INV_X1 U14219 ( .A(n18025), .ZN(n9044) );
  AOI22_X1 U14220 ( .A1(\mem[969][4] ), .A2(n18021), .B1(n26161), .B2(
        data_in[4]), .ZN(n18025) );
  INV_X1 U14221 ( .A(n18026), .ZN(n9043) );
  AOI22_X1 U14222 ( .A1(\mem[969][5] ), .A2(n18021), .B1(n26161), .B2(
        data_in[5]), .ZN(n18026) );
  INV_X1 U14223 ( .A(n18027), .ZN(n9042) );
  AOI22_X1 U14224 ( .A1(\mem[969][6] ), .A2(n18021), .B1(n26161), .B2(
        data_in[6]), .ZN(n18027) );
  INV_X1 U14225 ( .A(n18028), .ZN(n9041) );
  AOI22_X1 U14226 ( .A1(\mem[969][7] ), .A2(n18021), .B1(n26161), .B2(
        data_in[7]), .ZN(n18028) );
  INV_X1 U14227 ( .A(n18029), .ZN(n9040) );
  AOI22_X1 U14228 ( .A1(\mem[970][0] ), .A2(n18030), .B1(n26160), .B2(
        data_in[0]), .ZN(n18029) );
  INV_X1 U14229 ( .A(n18031), .ZN(n9039) );
  AOI22_X1 U14230 ( .A1(\mem[970][1] ), .A2(n18030), .B1(n26160), .B2(
        data_in[1]), .ZN(n18031) );
  INV_X1 U14231 ( .A(n18032), .ZN(n9038) );
  AOI22_X1 U14232 ( .A1(\mem[970][2] ), .A2(n18030), .B1(n26160), .B2(
        data_in[2]), .ZN(n18032) );
  INV_X1 U14233 ( .A(n18033), .ZN(n9037) );
  AOI22_X1 U14234 ( .A1(\mem[970][3] ), .A2(n18030), .B1(n26160), .B2(
        data_in[3]), .ZN(n18033) );
  INV_X1 U14235 ( .A(n18034), .ZN(n9036) );
  AOI22_X1 U14236 ( .A1(\mem[970][4] ), .A2(n18030), .B1(n26160), .B2(
        data_in[4]), .ZN(n18034) );
  INV_X1 U14237 ( .A(n18035), .ZN(n9035) );
  AOI22_X1 U14238 ( .A1(\mem[970][5] ), .A2(n18030), .B1(n26160), .B2(
        data_in[5]), .ZN(n18035) );
  INV_X1 U14239 ( .A(n18036), .ZN(n9034) );
  AOI22_X1 U14240 ( .A1(\mem[970][6] ), .A2(n18030), .B1(n26160), .B2(
        data_in[6]), .ZN(n18036) );
  INV_X1 U14241 ( .A(n18037), .ZN(n9033) );
  AOI22_X1 U14242 ( .A1(\mem[970][7] ), .A2(n18030), .B1(n26160), .B2(
        data_in[7]), .ZN(n18037) );
  INV_X1 U14243 ( .A(n18038), .ZN(n9032) );
  AOI22_X1 U14244 ( .A1(\mem[971][0] ), .A2(n18039), .B1(n26159), .B2(
        data_in[0]), .ZN(n18038) );
  INV_X1 U14245 ( .A(n18040), .ZN(n9031) );
  AOI22_X1 U14246 ( .A1(\mem[971][1] ), .A2(n18039), .B1(n26159), .B2(
        data_in[1]), .ZN(n18040) );
  INV_X1 U14247 ( .A(n18041), .ZN(n9030) );
  AOI22_X1 U14248 ( .A1(\mem[971][2] ), .A2(n18039), .B1(n26159), .B2(
        data_in[2]), .ZN(n18041) );
  INV_X1 U14249 ( .A(n18042), .ZN(n9029) );
  AOI22_X1 U14250 ( .A1(\mem[971][3] ), .A2(n18039), .B1(n26159), .B2(
        data_in[3]), .ZN(n18042) );
  INV_X1 U14251 ( .A(n18043), .ZN(n9028) );
  AOI22_X1 U14252 ( .A1(\mem[971][4] ), .A2(n18039), .B1(n26159), .B2(
        data_in[4]), .ZN(n18043) );
  INV_X1 U14253 ( .A(n18044), .ZN(n9027) );
  AOI22_X1 U14254 ( .A1(\mem[971][5] ), .A2(n18039), .B1(n26159), .B2(
        data_in[5]), .ZN(n18044) );
  INV_X1 U14255 ( .A(n18045), .ZN(n9026) );
  AOI22_X1 U14256 ( .A1(\mem[971][6] ), .A2(n18039), .B1(n26159), .B2(
        data_in[6]), .ZN(n18045) );
  INV_X1 U14257 ( .A(n18046), .ZN(n9025) );
  AOI22_X1 U14258 ( .A1(\mem[971][7] ), .A2(n18039), .B1(n26159), .B2(
        data_in[7]), .ZN(n18046) );
  INV_X1 U14259 ( .A(n18047), .ZN(n9024) );
  AOI22_X1 U14260 ( .A1(\mem[972][0] ), .A2(n18048), .B1(n26158), .B2(
        data_in[0]), .ZN(n18047) );
  INV_X1 U14261 ( .A(n18049), .ZN(n9023) );
  AOI22_X1 U14262 ( .A1(\mem[972][1] ), .A2(n18048), .B1(n26158), .B2(
        data_in[1]), .ZN(n18049) );
  INV_X1 U14263 ( .A(n18050), .ZN(n9022) );
  AOI22_X1 U14264 ( .A1(\mem[972][2] ), .A2(n18048), .B1(n26158), .B2(
        data_in[2]), .ZN(n18050) );
  INV_X1 U14265 ( .A(n18051), .ZN(n9021) );
  AOI22_X1 U14266 ( .A1(\mem[972][3] ), .A2(n18048), .B1(n26158), .B2(
        data_in[3]), .ZN(n18051) );
  INV_X1 U14267 ( .A(n18052), .ZN(n9020) );
  AOI22_X1 U14268 ( .A1(\mem[972][4] ), .A2(n18048), .B1(n26158), .B2(
        data_in[4]), .ZN(n18052) );
  INV_X1 U14269 ( .A(n18053), .ZN(n9019) );
  AOI22_X1 U14270 ( .A1(\mem[972][5] ), .A2(n18048), .B1(n26158), .B2(
        data_in[5]), .ZN(n18053) );
  INV_X1 U14271 ( .A(n18054), .ZN(n9018) );
  AOI22_X1 U14272 ( .A1(\mem[972][6] ), .A2(n18048), .B1(n26158), .B2(
        data_in[6]), .ZN(n18054) );
  INV_X1 U14273 ( .A(n18055), .ZN(n9017) );
  AOI22_X1 U14274 ( .A1(\mem[972][7] ), .A2(n18048), .B1(n26158), .B2(
        data_in[7]), .ZN(n18055) );
  INV_X1 U14275 ( .A(n18056), .ZN(n9016) );
  AOI22_X1 U14276 ( .A1(\mem[973][0] ), .A2(n18057), .B1(n26157), .B2(
        data_in[0]), .ZN(n18056) );
  INV_X1 U14277 ( .A(n18058), .ZN(n9015) );
  AOI22_X1 U14278 ( .A1(\mem[973][1] ), .A2(n18057), .B1(n26157), .B2(
        data_in[1]), .ZN(n18058) );
  INV_X1 U14279 ( .A(n18059), .ZN(n9014) );
  AOI22_X1 U14280 ( .A1(\mem[973][2] ), .A2(n18057), .B1(n26157), .B2(
        data_in[2]), .ZN(n18059) );
  INV_X1 U14281 ( .A(n18060), .ZN(n9013) );
  AOI22_X1 U14282 ( .A1(\mem[973][3] ), .A2(n18057), .B1(n26157), .B2(
        data_in[3]), .ZN(n18060) );
  INV_X1 U14283 ( .A(n18061), .ZN(n9012) );
  AOI22_X1 U14284 ( .A1(\mem[973][4] ), .A2(n18057), .B1(n26157), .B2(
        data_in[4]), .ZN(n18061) );
  INV_X1 U14285 ( .A(n18062), .ZN(n9011) );
  AOI22_X1 U14286 ( .A1(\mem[973][5] ), .A2(n18057), .B1(n26157), .B2(
        data_in[5]), .ZN(n18062) );
  INV_X1 U14287 ( .A(n18063), .ZN(n9010) );
  AOI22_X1 U14288 ( .A1(\mem[973][6] ), .A2(n18057), .B1(n26157), .B2(
        data_in[6]), .ZN(n18063) );
  INV_X1 U14289 ( .A(n18064), .ZN(n9009) );
  AOI22_X1 U14290 ( .A1(\mem[973][7] ), .A2(n18057), .B1(n26157), .B2(
        data_in[7]), .ZN(n18064) );
  INV_X1 U14291 ( .A(n18065), .ZN(n9008) );
  AOI22_X1 U14292 ( .A1(\mem[974][0] ), .A2(n18066), .B1(n26156), .B2(
        data_in[0]), .ZN(n18065) );
  INV_X1 U14293 ( .A(n18067), .ZN(n9007) );
  AOI22_X1 U14294 ( .A1(\mem[974][1] ), .A2(n18066), .B1(n26156), .B2(
        data_in[1]), .ZN(n18067) );
  INV_X1 U14295 ( .A(n18068), .ZN(n9006) );
  AOI22_X1 U14296 ( .A1(\mem[974][2] ), .A2(n18066), .B1(n26156), .B2(
        data_in[2]), .ZN(n18068) );
  INV_X1 U14297 ( .A(n18069), .ZN(n9005) );
  AOI22_X1 U14298 ( .A1(\mem[974][3] ), .A2(n18066), .B1(n26156), .B2(
        data_in[3]), .ZN(n18069) );
  INV_X1 U14299 ( .A(n18070), .ZN(n9004) );
  AOI22_X1 U14300 ( .A1(\mem[974][4] ), .A2(n18066), .B1(n26156), .B2(
        data_in[4]), .ZN(n18070) );
  INV_X1 U14301 ( .A(n18071), .ZN(n9003) );
  AOI22_X1 U14302 ( .A1(\mem[974][5] ), .A2(n18066), .B1(n26156), .B2(
        data_in[5]), .ZN(n18071) );
  INV_X1 U14303 ( .A(n18072), .ZN(n9002) );
  AOI22_X1 U14304 ( .A1(\mem[974][6] ), .A2(n18066), .B1(n26156), .B2(
        data_in[6]), .ZN(n18072) );
  INV_X1 U14305 ( .A(n18073), .ZN(n9001) );
  AOI22_X1 U14306 ( .A1(\mem[974][7] ), .A2(n18066), .B1(n26156), .B2(
        data_in[7]), .ZN(n18073) );
  INV_X1 U14307 ( .A(n18074), .ZN(n9000) );
  AOI22_X1 U14308 ( .A1(\mem[975][0] ), .A2(n18075), .B1(n26155), .B2(
        data_in[0]), .ZN(n18074) );
  INV_X1 U14309 ( .A(n18076), .ZN(n8999) );
  AOI22_X1 U14310 ( .A1(\mem[975][1] ), .A2(n18075), .B1(n26155), .B2(
        data_in[1]), .ZN(n18076) );
  INV_X1 U14311 ( .A(n18077), .ZN(n8998) );
  AOI22_X1 U14312 ( .A1(\mem[975][2] ), .A2(n18075), .B1(n26155), .B2(
        data_in[2]), .ZN(n18077) );
  INV_X1 U14313 ( .A(n18078), .ZN(n8997) );
  AOI22_X1 U14314 ( .A1(\mem[975][3] ), .A2(n18075), .B1(n26155), .B2(
        data_in[3]), .ZN(n18078) );
  INV_X1 U14315 ( .A(n18079), .ZN(n8996) );
  AOI22_X1 U14316 ( .A1(\mem[975][4] ), .A2(n18075), .B1(n26155), .B2(
        data_in[4]), .ZN(n18079) );
  INV_X1 U14317 ( .A(n18080), .ZN(n8995) );
  AOI22_X1 U14318 ( .A1(\mem[975][5] ), .A2(n18075), .B1(n26155), .B2(
        data_in[5]), .ZN(n18080) );
  INV_X1 U14319 ( .A(n18081), .ZN(n8994) );
  AOI22_X1 U14320 ( .A1(\mem[975][6] ), .A2(n18075), .B1(n26155), .B2(
        data_in[6]), .ZN(n18081) );
  INV_X1 U14321 ( .A(n18082), .ZN(n8993) );
  AOI22_X1 U14322 ( .A1(\mem[975][7] ), .A2(n18075), .B1(n26155), .B2(
        data_in[7]), .ZN(n18082) );
  INV_X1 U14323 ( .A(n18083), .ZN(n8992) );
  AOI22_X1 U14324 ( .A1(\mem[976][0] ), .A2(n18084), .B1(n26154), .B2(
        data_in[0]), .ZN(n18083) );
  INV_X1 U14325 ( .A(n18085), .ZN(n8991) );
  AOI22_X1 U14326 ( .A1(\mem[976][1] ), .A2(n18084), .B1(n26154), .B2(
        data_in[1]), .ZN(n18085) );
  INV_X1 U14327 ( .A(n18086), .ZN(n8990) );
  AOI22_X1 U14328 ( .A1(\mem[976][2] ), .A2(n18084), .B1(n26154), .B2(
        data_in[2]), .ZN(n18086) );
  INV_X1 U14329 ( .A(n18087), .ZN(n8989) );
  AOI22_X1 U14330 ( .A1(\mem[976][3] ), .A2(n18084), .B1(n26154), .B2(
        data_in[3]), .ZN(n18087) );
  INV_X1 U14331 ( .A(n18088), .ZN(n8988) );
  AOI22_X1 U14332 ( .A1(\mem[976][4] ), .A2(n18084), .B1(n26154), .B2(
        data_in[4]), .ZN(n18088) );
  INV_X1 U14333 ( .A(n18089), .ZN(n8987) );
  AOI22_X1 U14334 ( .A1(\mem[976][5] ), .A2(n18084), .B1(n26154), .B2(
        data_in[5]), .ZN(n18089) );
  INV_X1 U14335 ( .A(n18090), .ZN(n8986) );
  AOI22_X1 U14336 ( .A1(\mem[976][6] ), .A2(n18084), .B1(n26154), .B2(
        data_in[6]), .ZN(n18090) );
  INV_X1 U14337 ( .A(n18091), .ZN(n8985) );
  AOI22_X1 U14338 ( .A1(\mem[976][7] ), .A2(n18084), .B1(n26154), .B2(
        data_in[7]), .ZN(n18091) );
  INV_X1 U14339 ( .A(n18092), .ZN(n8984) );
  AOI22_X1 U14340 ( .A1(\mem[977][0] ), .A2(n18093), .B1(n26153), .B2(
        data_in[0]), .ZN(n18092) );
  INV_X1 U14341 ( .A(n18094), .ZN(n8983) );
  AOI22_X1 U14342 ( .A1(\mem[977][1] ), .A2(n18093), .B1(n26153), .B2(
        data_in[1]), .ZN(n18094) );
  INV_X1 U14343 ( .A(n18095), .ZN(n8982) );
  AOI22_X1 U14344 ( .A1(\mem[977][2] ), .A2(n18093), .B1(n26153), .B2(
        data_in[2]), .ZN(n18095) );
  INV_X1 U14345 ( .A(n18096), .ZN(n8981) );
  AOI22_X1 U14346 ( .A1(\mem[977][3] ), .A2(n18093), .B1(n26153), .B2(
        data_in[3]), .ZN(n18096) );
  INV_X1 U14347 ( .A(n18097), .ZN(n8980) );
  AOI22_X1 U14348 ( .A1(\mem[977][4] ), .A2(n18093), .B1(n26153), .B2(
        data_in[4]), .ZN(n18097) );
  INV_X1 U14349 ( .A(n18098), .ZN(n8979) );
  AOI22_X1 U14350 ( .A1(\mem[977][5] ), .A2(n18093), .B1(n26153), .B2(
        data_in[5]), .ZN(n18098) );
  INV_X1 U14351 ( .A(n18099), .ZN(n8978) );
  AOI22_X1 U14352 ( .A1(\mem[977][6] ), .A2(n18093), .B1(n26153), .B2(
        data_in[6]), .ZN(n18099) );
  INV_X1 U14353 ( .A(n18100), .ZN(n8977) );
  AOI22_X1 U14354 ( .A1(\mem[977][7] ), .A2(n18093), .B1(n26153), .B2(
        data_in[7]), .ZN(n18100) );
  INV_X1 U14355 ( .A(n18101), .ZN(n8976) );
  AOI22_X1 U14356 ( .A1(\mem[978][0] ), .A2(n18102), .B1(n26152), .B2(
        data_in[0]), .ZN(n18101) );
  INV_X1 U14357 ( .A(n18103), .ZN(n8975) );
  AOI22_X1 U14358 ( .A1(\mem[978][1] ), .A2(n18102), .B1(n26152), .B2(
        data_in[1]), .ZN(n18103) );
  INV_X1 U14359 ( .A(n18104), .ZN(n8974) );
  AOI22_X1 U14360 ( .A1(\mem[978][2] ), .A2(n18102), .B1(n26152), .B2(
        data_in[2]), .ZN(n18104) );
  INV_X1 U14361 ( .A(n18105), .ZN(n8973) );
  AOI22_X1 U14362 ( .A1(\mem[978][3] ), .A2(n18102), .B1(n26152), .B2(
        data_in[3]), .ZN(n18105) );
  INV_X1 U14363 ( .A(n18106), .ZN(n8972) );
  AOI22_X1 U14364 ( .A1(\mem[978][4] ), .A2(n18102), .B1(n26152), .B2(
        data_in[4]), .ZN(n18106) );
  INV_X1 U14365 ( .A(n18107), .ZN(n8971) );
  AOI22_X1 U14366 ( .A1(\mem[978][5] ), .A2(n18102), .B1(n26152), .B2(
        data_in[5]), .ZN(n18107) );
  INV_X1 U14367 ( .A(n18108), .ZN(n8970) );
  AOI22_X1 U14368 ( .A1(\mem[978][6] ), .A2(n18102), .B1(n26152), .B2(
        data_in[6]), .ZN(n18108) );
  INV_X1 U14369 ( .A(n18109), .ZN(n8969) );
  AOI22_X1 U14370 ( .A1(\mem[978][7] ), .A2(n18102), .B1(n26152), .B2(
        data_in[7]), .ZN(n18109) );
  INV_X1 U14371 ( .A(n18110), .ZN(n8968) );
  AOI22_X1 U14372 ( .A1(\mem[979][0] ), .A2(n18111), .B1(n26151), .B2(
        data_in[0]), .ZN(n18110) );
  INV_X1 U14373 ( .A(n18112), .ZN(n8967) );
  AOI22_X1 U14374 ( .A1(\mem[979][1] ), .A2(n18111), .B1(n26151), .B2(
        data_in[1]), .ZN(n18112) );
  INV_X1 U14375 ( .A(n18113), .ZN(n8966) );
  AOI22_X1 U14376 ( .A1(\mem[979][2] ), .A2(n18111), .B1(n26151), .B2(
        data_in[2]), .ZN(n18113) );
  INV_X1 U14377 ( .A(n18114), .ZN(n8965) );
  AOI22_X1 U14378 ( .A1(\mem[979][3] ), .A2(n18111), .B1(n26151), .B2(
        data_in[3]), .ZN(n18114) );
  INV_X1 U14379 ( .A(n18115), .ZN(n8964) );
  AOI22_X1 U14380 ( .A1(\mem[979][4] ), .A2(n18111), .B1(n26151), .B2(
        data_in[4]), .ZN(n18115) );
  INV_X1 U14381 ( .A(n18116), .ZN(n8963) );
  AOI22_X1 U14382 ( .A1(\mem[979][5] ), .A2(n18111), .B1(n26151), .B2(
        data_in[5]), .ZN(n18116) );
  INV_X1 U14383 ( .A(n18117), .ZN(n8962) );
  AOI22_X1 U14384 ( .A1(\mem[979][6] ), .A2(n18111), .B1(n26151), .B2(
        data_in[6]), .ZN(n18117) );
  INV_X1 U14385 ( .A(n18118), .ZN(n8961) );
  AOI22_X1 U14386 ( .A1(\mem[979][7] ), .A2(n18111), .B1(n26151), .B2(
        data_in[7]), .ZN(n18118) );
  INV_X1 U14387 ( .A(n18119), .ZN(n8960) );
  AOI22_X1 U14388 ( .A1(\mem[980][0] ), .A2(n18120), .B1(n26150), .B2(
        data_in[0]), .ZN(n18119) );
  INV_X1 U14389 ( .A(n18121), .ZN(n8959) );
  AOI22_X1 U14390 ( .A1(\mem[980][1] ), .A2(n18120), .B1(n26150), .B2(
        data_in[1]), .ZN(n18121) );
  INV_X1 U14391 ( .A(n18122), .ZN(n8958) );
  AOI22_X1 U14392 ( .A1(\mem[980][2] ), .A2(n18120), .B1(n26150), .B2(
        data_in[2]), .ZN(n18122) );
  INV_X1 U14393 ( .A(n18123), .ZN(n8957) );
  AOI22_X1 U14394 ( .A1(\mem[980][3] ), .A2(n18120), .B1(n26150), .B2(
        data_in[3]), .ZN(n18123) );
  INV_X1 U14395 ( .A(n18124), .ZN(n8956) );
  AOI22_X1 U14396 ( .A1(\mem[980][4] ), .A2(n18120), .B1(n26150), .B2(
        data_in[4]), .ZN(n18124) );
  INV_X1 U14397 ( .A(n18125), .ZN(n8955) );
  AOI22_X1 U14398 ( .A1(\mem[980][5] ), .A2(n18120), .B1(n26150), .B2(
        data_in[5]), .ZN(n18125) );
  INV_X1 U14399 ( .A(n18126), .ZN(n8954) );
  AOI22_X1 U14400 ( .A1(\mem[980][6] ), .A2(n18120), .B1(n26150), .B2(
        data_in[6]), .ZN(n18126) );
  INV_X1 U14401 ( .A(n18127), .ZN(n8953) );
  AOI22_X1 U14402 ( .A1(\mem[980][7] ), .A2(n18120), .B1(n26150), .B2(
        data_in[7]), .ZN(n18127) );
  INV_X1 U14403 ( .A(n18128), .ZN(n8952) );
  AOI22_X1 U14404 ( .A1(\mem[981][0] ), .A2(n18129), .B1(n26149), .B2(
        data_in[0]), .ZN(n18128) );
  INV_X1 U14405 ( .A(n18130), .ZN(n8951) );
  AOI22_X1 U14406 ( .A1(\mem[981][1] ), .A2(n18129), .B1(n26149), .B2(
        data_in[1]), .ZN(n18130) );
  INV_X1 U14407 ( .A(n18131), .ZN(n8950) );
  AOI22_X1 U14408 ( .A1(\mem[981][2] ), .A2(n18129), .B1(n26149), .B2(
        data_in[2]), .ZN(n18131) );
  INV_X1 U14409 ( .A(n18132), .ZN(n8949) );
  AOI22_X1 U14410 ( .A1(\mem[981][3] ), .A2(n18129), .B1(n26149), .B2(
        data_in[3]), .ZN(n18132) );
  INV_X1 U14411 ( .A(n18133), .ZN(n8948) );
  AOI22_X1 U14412 ( .A1(\mem[981][4] ), .A2(n18129), .B1(n26149), .B2(
        data_in[4]), .ZN(n18133) );
  INV_X1 U14413 ( .A(n18134), .ZN(n8947) );
  AOI22_X1 U14414 ( .A1(\mem[981][5] ), .A2(n18129), .B1(n26149), .B2(
        data_in[5]), .ZN(n18134) );
  INV_X1 U14415 ( .A(n18135), .ZN(n8946) );
  AOI22_X1 U14416 ( .A1(\mem[981][6] ), .A2(n18129), .B1(n26149), .B2(
        data_in[6]), .ZN(n18135) );
  INV_X1 U14417 ( .A(n18136), .ZN(n8945) );
  AOI22_X1 U14418 ( .A1(\mem[981][7] ), .A2(n18129), .B1(n26149), .B2(
        data_in[7]), .ZN(n18136) );
  INV_X1 U14419 ( .A(n18137), .ZN(n8944) );
  AOI22_X1 U14420 ( .A1(\mem[982][0] ), .A2(n18138), .B1(n26148), .B2(
        data_in[0]), .ZN(n18137) );
  INV_X1 U14421 ( .A(n18139), .ZN(n8943) );
  AOI22_X1 U14422 ( .A1(\mem[982][1] ), .A2(n18138), .B1(n26148), .B2(
        data_in[1]), .ZN(n18139) );
  INV_X1 U14423 ( .A(n18140), .ZN(n8942) );
  AOI22_X1 U14424 ( .A1(\mem[982][2] ), .A2(n18138), .B1(n26148), .B2(
        data_in[2]), .ZN(n18140) );
  INV_X1 U14425 ( .A(n18141), .ZN(n8941) );
  AOI22_X1 U14426 ( .A1(\mem[982][3] ), .A2(n18138), .B1(n26148), .B2(
        data_in[3]), .ZN(n18141) );
  INV_X1 U14427 ( .A(n18142), .ZN(n8940) );
  AOI22_X1 U14428 ( .A1(\mem[982][4] ), .A2(n18138), .B1(n26148), .B2(
        data_in[4]), .ZN(n18142) );
  INV_X1 U14429 ( .A(n18143), .ZN(n8939) );
  AOI22_X1 U14430 ( .A1(\mem[982][5] ), .A2(n18138), .B1(n26148), .B2(
        data_in[5]), .ZN(n18143) );
  INV_X1 U14431 ( .A(n18144), .ZN(n8938) );
  AOI22_X1 U14432 ( .A1(\mem[982][6] ), .A2(n18138), .B1(n26148), .B2(
        data_in[6]), .ZN(n18144) );
  INV_X1 U14433 ( .A(n18145), .ZN(n8937) );
  AOI22_X1 U14434 ( .A1(\mem[982][7] ), .A2(n18138), .B1(n26148), .B2(
        data_in[7]), .ZN(n18145) );
  INV_X1 U14435 ( .A(n18146), .ZN(n8936) );
  AOI22_X1 U14436 ( .A1(\mem[983][0] ), .A2(n18147), .B1(n26147), .B2(
        data_in[0]), .ZN(n18146) );
  INV_X1 U14437 ( .A(n18148), .ZN(n8935) );
  AOI22_X1 U14438 ( .A1(\mem[983][1] ), .A2(n18147), .B1(n26147), .B2(
        data_in[1]), .ZN(n18148) );
  INV_X1 U14439 ( .A(n18149), .ZN(n8934) );
  AOI22_X1 U14440 ( .A1(\mem[983][2] ), .A2(n18147), .B1(n26147), .B2(
        data_in[2]), .ZN(n18149) );
  INV_X1 U14441 ( .A(n18150), .ZN(n8933) );
  AOI22_X1 U14442 ( .A1(\mem[983][3] ), .A2(n18147), .B1(n26147), .B2(
        data_in[3]), .ZN(n18150) );
  INV_X1 U14443 ( .A(n18151), .ZN(n8932) );
  AOI22_X1 U14444 ( .A1(\mem[983][4] ), .A2(n18147), .B1(n26147), .B2(
        data_in[4]), .ZN(n18151) );
  INV_X1 U14445 ( .A(n18152), .ZN(n8931) );
  AOI22_X1 U14446 ( .A1(\mem[983][5] ), .A2(n18147), .B1(n26147), .B2(
        data_in[5]), .ZN(n18152) );
  INV_X1 U14447 ( .A(n18153), .ZN(n8930) );
  AOI22_X1 U14448 ( .A1(\mem[983][6] ), .A2(n18147), .B1(n26147), .B2(
        data_in[6]), .ZN(n18153) );
  INV_X1 U14449 ( .A(n18154), .ZN(n8929) );
  AOI22_X1 U14450 ( .A1(\mem[983][7] ), .A2(n18147), .B1(n26147), .B2(
        data_in[7]), .ZN(n18154) );
  INV_X1 U14451 ( .A(n18155), .ZN(n8928) );
  AOI22_X1 U14452 ( .A1(\mem[984][0] ), .A2(n18156), .B1(n26146), .B2(
        data_in[0]), .ZN(n18155) );
  INV_X1 U14453 ( .A(n18157), .ZN(n8927) );
  AOI22_X1 U14454 ( .A1(\mem[984][1] ), .A2(n18156), .B1(n26146), .B2(
        data_in[1]), .ZN(n18157) );
  INV_X1 U14455 ( .A(n18158), .ZN(n8926) );
  AOI22_X1 U14456 ( .A1(\mem[984][2] ), .A2(n18156), .B1(n26146), .B2(
        data_in[2]), .ZN(n18158) );
  INV_X1 U14457 ( .A(n18159), .ZN(n8925) );
  AOI22_X1 U14458 ( .A1(\mem[984][3] ), .A2(n18156), .B1(n26146), .B2(
        data_in[3]), .ZN(n18159) );
  INV_X1 U14459 ( .A(n18160), .ZN(n8924) );
  AOI22_X1 U14460 ( .A1(\mem[984][4] ), .A2(n18156), .B1(n26146), .B2(
        data_in[4]), .ZN(n18160) );
  INV_X1 U14461 ( .A(n18161), .ZN(n8923) );
  AOI22_X1 U14462 ( .A1(\mem[984][5] ), .A2(n18156), .B1(n26146), .B2(
        data_in[5]), .ZN(n18161) );
  INV_X1 U14463 ( .A(n18162), .ZN(n8922) );
  AOI22_X1 U14464 ( .A1(\mem[984][6] ), .A2(n18156), .B1(n26146), .B2(
        data_in[6]), .ZN(n18162) );
  INV_X1 U14465 ( .A(n18163), .ZN(n8921) );
  AOI22_X1 U14466 ( .A1(\mem[984][7] ), .A2(n18156), .B1(n26146), .B2(
        data_in[7]), .ZN(n18163) );
  INV_X1 U14467 ( .A(n18164), .ZN(n8920) );
  AOI22_X1 U14468 ( .A1(\mem[985][0] ), .A2(n18165), .B1(n26145), .B2(
        data_in[0]), .ZN(n18164) );
  INV_X1 U14469 ( .A(n18166), .ZN(n8919) );
  AOI22_X1 U14470 ( .A1(\mem[985][1] ), .A2(n18165), .B1(n26145), .B2(
        data_in[1]), .ZN(n18166) );
  INV_X1 U14471 ( .A(n18167), .ZN(n8918) );
  AOI22_X1 U14472 ( .A1(\mem[985][2] ), .A2(n18165), .B1(n26145), .B2(
        data_in[2]), .ZN(n18167) );
  INV_X1 U14473 ( .A(n18168), .ZN(n8917) );
  AOI22_X1 U14474 ( .A1(\mem[985][3] ), .A2(n18165), .B1(n26145), .B2(
        data_in[3]), .ZN(n18168) );
  INV_X1 U14475 ( .A(n18169), .ZN(n8916) );
  AOI22_X1 U14476 ( .A1(\mem[985][4] ), .A2(n18165), .B1(n26145), .B2(
        data_in[4]), .ZN(n18169) );
  INV_X1 U14477 ( .A(n18170), .ZN(n8915) );
  AOI22_X1 U14478 ( .A1(\mem[985][5] ), .A2(n18165), .B1(n26145), .B2(
        data_in[5]), .ZN(n18170) );
  INV_X1 U14479 ( .A(n18171), .ZN(n8914) );
  AOI22_X1 U14480 ( .A1(\mem[985][6] ), .A2(n18165), .B1(n26145), .B2(
        data_in[6]), .ZN(n18171) );
  INV_X1 U14481 ( .A(n18172), .ZN(n8913) );
  AOI22_X1 U14482 ( .A1(\mem[985][7] ), .A2(n18165), .B1(n26145), .B2(
        data_in[7]), .ZN(n18172) );
  INV_X1 U14483 ( .A(n18173), .ZN(n8912) );
  AOI22_X1 U14484 ( .A1(\mem[986][0] ), .A2(n18174), .B1(n26144), .B2(
        data_in[0]), .ZN(n18173) );
  INV_X1 U14485 ( .A(n18175), .ZN(n8911) );
  AOI22_X1 U14486 ( .A1(\mem[986][1] ), .A2(n18174), .B1(n26144), .B2(
        data_in[1]), .ZN(n18175) );
  INV_X1 U14487 ( .A(n18176), .ZN(n8910) );
  AOI22_X1 U14488 ( .A1(\mem[986][2] ), .A2(n18174), .B1(n26144), .B2(
        data_in[2]), .ZN(n18176) );
  INV_X1 U14489 ( .A(n18177), .ZN(n8909) );
  AOI22_X1 U14490 ( .A1(\mem[986][3] ), .A2(n18174), .B1(n26144), .B2(
        data_in[3]), .ZN(n18177) );
  INV_X1 U14491 ( .A(n18178), .ZN(n8908) );
  AOI22_X1 U14492 ( .A1(\mem[986][4] ), .A2(n18174), .B1(n26144), .B2(
        data_in[4]), .ZN(n18178) );
  INV_X1 U14493 ( .A(n18179), .ZN(n8907) );
  AOI22_X1 U14494 ( .A1(\mem[986][5] ), .A2(n18174), .B1(n26144), .B2(
        data_in[5]), .ZN(n18179) );
  INV_X1 U14495 ( .A(n18180), .ZN(n8906) );
  AOI22_X1 U14496 ( .A1(\mem[986][6] ), .A2(n18174), .B1(n26144), .B2(
        data_in[6]), .ZN(n18180) );
  INV_X1 U14497 ( .A(n18181), .ZN(n8905) );
  AOI22_X1 U14498 ( .A1(\mem[986][7] ), .A2(n18174), .B1(n26144), .B2(
        data_in[7]), .ZN(n18181) );
  INV_X1 U14499 ( .A(n18182), .ZN(n8904) );
  AOI22_X1 U14500 ( .A1(\mem[987][0] ), .A2(n18183), .B1(n26143), .B2(
        data_in[0]), .ZN(n18182) );
  INV_X1 U14501 ( .A(n18184), .ZN(n8903) );
  AOI22_X1 U14502 ( .A1(\mem[987][1] ), .A2(n18183), .B1(n26143), .B2(
        data_in[1]), .ZN(n18184) );
  INV_X1 U14503 ( .A(n18185), .ZN(n8902) );
  AOI22_X1 U14504 ( .A1(\mem[987][2] ), .A2(n18183), .B1(n26143), .B2(
        data_in[2]), .ZN(n18185) );
  INV_X1 U14505 ( .A(n18186), .ZN(n8901) );
  AOI22_X1 U14506 ( .A1(\mem[987][3] ), .A2(n18183), .B1(n26143), .B2(
        data_in[3]), .ZN(n18186) );
  INV_X1 U14507 ( .A(n18187), .ZN(n8900) );
  AOI22_X1 U14508 ( .A1(\mem[987][4] ), .A2(n18183), .B1(n26143), .B2(
        data_in[4]), .ZN(n18187) );
  INV_X1 U14509 ( .A(n18188), .ZN(n8899) );
  AOI22_X1 U14510 ( .A1(\mem[987][5] ), .A2(n18183), .B1(n26143), .B2(
        data_in[5]), .ZN(n18188) );
  INV_X1 U14511 ( .A(n18189), .ZN(n8898) );
  AOI22_X1 U14512 ( .A1(\mem[987][6] ), .A2(n18183), .B1(n26143), .B2(
        data_in[6]), .ZN(n18189) );
  INV_X1 U14513 ( .A(n18190), .ZN(n8897) );
  AOI22_X1 U14514 ( .A1(\mem[987][7] ), .A2(n18183), .B1(n26143), .B2(
        data_in[7]), .ZN(n18190) );
  INV_X1 U14515 ( .A(n18191), .ZN(n8896) );
  AOI22_X1 U14516 ( .A1(\mem[988][0] ), .A2(n18192), .B1(n26142), .B2(
        data_in[0]), .ZN(n18191) );
  INV_X1 U14517 ( .A(n18193), .ZN(n8895) );
  AOI22_X1 U14518 ( .A1(\mem[988][1] ), .A2(n18192), .B1(n26142), .B2(
        data_in[1]), .ZN(n18193) );
  INV_X1 U14519 ( .A(n18194), .ZN(n8894) );
  AOI22_X1 U14520 ( .A1(\mem[988][2] ), .A2(n18192), .B1(n26142), .B2(
        data_in[2]), .ZN(n18194) );
  INV_X1 U14521 ( .A(n18195), .ZN(n8893) );
  AOI22_X1 U14522 ( .A1(\mem[988][3] ), .A2(n18192), .B1(n26142), .B2(
        data_in[3]), .ZN(n18195) );
  INV_X1 U14523 ( .A(n18196), .ZN(n8892) );
  AOI22_X1 U14524 ( .A1(\mem[988][4] ), .A2(n18192), .B1(n26142), .B2(
        data_in[4]), .ZN(n18196) );
  INV_X1 U14525 ( .A(n18197), .ZN(n8891) );
  AOI22_X1 U14526 ( .A1(\mem[988][5] ), .A2(n18192), .B1(n26142), .B2(
        data_in[5]), .ZN(n18197) );
  INV_X1 U14527 ( .A(n18198), .ZN(n8890) );
  AOI22_X1 U14528 ( .A1(\mem[988][6] ), .A2(n18192), .B1(n26142), .B2(
        data_in[6]), .ZN(n18198) );
  INV_X1 U14529 ( .A(n18199), .ZN(n8889) );
  AOI22_X1 U14530 ( .A1(\mem[988][7] ), .A2(n18192), .B1(n26142), .B2(
        data_in[7]), .ZN(n18199) );
  INV_X1 U14531 ( .A(n18200), .ZN(n8888) );
  AOI22_X1 U14532 ( .A1(\mem[989][0] ), .A2(n18201), .B1(n26141), .B2(
        data_in[0]), .ZN(n18200) );
  INV_X1 U14533 ( .A(n18202), .ZN(n8887) );
  AOI22_X1 U14534 ( .A1(\mem[989][1] ), .A2(n18201), .B1(n26141), .B2(
        data_in[1]), .ZN(n18202) );
  INV_X1 U14535 ( .A(n18203), .ZN(n8886) );
  AOI22_X1 U14536 ( .A1(\mem[989][2] ), .A2(n18201), .B1(n26141), .B2(
        data_in[2]), .ZN(n18203) );
  INV_X1 U14537 ( .A(n18204), .ZN(n8885) );
  AOI22_X1 U14538 ( .A1(\mem[989][3] ), .A2(n18201), .B1(n26141), .B2(
        data_in[3]), .ZN(n18204) );
  INV_X1 U14539 ( .A(n18205), .ZN(n8884) );
  AOI22_X1 U14540 ( .A1(\mem[989][4] ), .A2(n18201), .B1(n26141), .B2(
        data_in[4]), .ZN(n18205) );
  INV_X1 U14541 ( .A(n18206), .ZN(n8883) );
  AOI22_X1 U14542 ( .A1(\mem[989][5] ), .A2(n18201), .B1(n26141), .B2(
        data_in[5]), .ZN(n18206) );
  INV_X1 U14543 ( .A(n18207), .ZN(n8882) );
  AOI22_X1 U14544 ( .A1(\mem[989][6] ), .A2(n18201), .B1(n26141), .B2(
        data_in[6]), .ZN(n18207) );
  INV_X1 U14545 ( .A(n18208), .ZN(n8881) );
  AOI22_X1 U14546 ( .A1(\mem[989][7] ), .A2(n18201), .B1(n26141), .B2(
        data_in[7]), .ZN(n18208) );
  INV_X1 U14547 ( .A(n18209), .ZN(n8880) );
  AOI22_X1 U14548 ( .A1(\mem[990][0] ), .A2(n18210), .B1(n26140), .B2(
        data_in[0]), .ZN(n18209) );
  INV_X1 U14549 ( .A(n18211), .ZN(n8879) );
  AOI22_X1 U14550 ( .A1(\mem[990][1] ), .A2(n18210), .B1(n26140), .B2(
        data_in[1]), .ZN(n18211) );
  INV_X1 U14551 ( .A(n18212), .ZN(n8878) );
  AOI22_X1 U14552 ( .A1(\mem[990][2] ), .A2(n18210), .B1(n26140), .B2(
        data_in[2]), .ZN(n18212) );
  INV_X1 U14553 ( .A(n18213), .ZN(n8877) );
  AOI22_X1 U14554 ( .A1(\mem[990][3] ), .A2(n18210), .B1(n26140), .B2(
        data_in[3]), .ZN(n18213) );
  INV_X1 U14555 ( .A(n18214), .ZN(n8876) );
  AOI22_X1 U14556 ( .A1(\mem[990][4] ), .A2(n18210), .B1(n26140), .B2(
        data_in[4]), .ZN(n18214) );
  INV_X1 U14557 ( .A(n18215), .ZN(n8875) );
  AOI22_X1 U14558 ( .A1(\mem[990][5] ), .A2(n18210), .B1(n26140), .B2(
        data_in[5]), .ZN(n18215) );
  INV_X1 U14559 ( .A(n18216), .ZN(n8874) );
  AOI22_X1 U14560 ( .A1(\mem[990][6] ), .A2(n18210), .B1(n26140), .B2(
        data_in[6]), .ZN(n18216) );
  INV_X1 U14561 ( .A(n18217), .ZN(n8873) );
  AOI22_X1 U14562 ( .A1(\mem[990][7] ), .A2(n18210), .B1(n26140), .B2(
        data_in[7]), .ZN(n18217) );
  INV_X1 U14563 ( .A(n18218), .ZN(n8872) );
  AOI22_X1 U14564 ( .A1(\mem[991][0] ), .A2(n18219), .B1(n26139), .B2(
        data_in[0]), .ZN(n18218) );
  INV_X1 U14565 ( .A(n18220), .ZN(n8871) );
  AOI22_X1 U14566 ( .A1(\mem[991][1] ), .A2(n18219), .B1(n26139), .B2(
        data_in[1]), .ZN(n18220) );
  INV_X1 U14567 ( .A(n18221), .ZN(n8870) );
  AOI22_X1 U14568 ( .A1(\mem[991][2] ), .A2(n18219), .B1(n26139), .B2(
        data_in[2]), .ZN(n18221) );
  INV_X1 U14569 ( .A(n18222), .ZN(n8869) );
  AOI22_X1 U14570 ( .A1(\mem[991][3] ), .A2(n18219), .B1(n26139), .B2(
        data_in[3]), .ZN(n18222) );
  INV_X1 U14571 ( .A(n18223), .ZN(n8868) );
  AOI22_X1 U14572 ( .A1(\mem[991][4] ), .A2(n18219), .B1(n26139), .B2(
        data_in[4]), .ZN(n18223) );
  INV_X1 U14573 ( .A(n18224), .ZN(n8867) );
  AOI22_X1 U14574 ( .A1(\mem[991][5] ), .A2(n18219), .B1(n26139), .B2(
        data_in[5]), .ZN(n18224) );
  INV_X1 U14575 ( .A(n18225), .ZN(n8866) );
  AOI22_X1 U14576 ( .A1(\mem[991][6] ), .A2(n18219), .B1(n26139), .B2(
        data_in[6]), .ZN(n18225) );
  INV_X1 U14577 ( .A(n18226), .ZN(n8865) );
  AOI22_X1 U14578 ( .A1(\mem[991][7] ), .A2(n18219), .B1(n26139), .B2(
        data_in[7]), .ZN(n18226) );
  INV_X1 U14579 ( .A(n18309), .ZN(n8800) );
  AOI22_X1 U14580 ( .A1(\mem[1000][0] ), .A2(n18310), .B1(n26130), .B2(
        data_in[0]), .ZN(n18309) );
  INV_X1 U14581 ( .A(n18311), .ZN(n8799) );
  AOI22_X1 U14582 ( .A1(\mem[1000][1] ), .A2(n18310), .B1(n26130), .B2(
        data_in[1]), .ZN(n18311) );
  INV_X1 U14583 ( .A(n18312), .ZN(n8798) );
  AOI22_X1 U14584 ( .A1(\mem[1000][2] ), .A2(n18310), .B1(n26130), .B2(
        data_in[2]), .ZN(n18312) );
  INV_X1 U14585 ( .A(n18313), .ZN(n8797) );
  AOI22_X1 U14586 ( .A1(\mem[1000][3] ), .A2(n18310), .B1(n26130), .B2(
        data_in[3]), .ZN(n18313) );
  INV_X1 U14587 ( .A(n18314), .ZN(n8796) );
  AOI22_X1 U14588 ( .A1(\mem[1000][4] ), .A2(n18310), .B1(n26130), .B2(
        data_in[4]), .ZN(n18314) );
  INV_X1 U14589 ( .A(n18315), .ZN(n8795) );
  AOI22_X1 U14590 ( .A1(\mem[1000][5] ), .A2(n18310), .B1(n26130), .B2(
        data_in[5]), .ZN(n18315) );
  INV_X1 U14591 ( .A(n18316), .ZN(n8794) );
  AOI22_X1 U14592 ( .A1(\mem[1000][6] ), .A2(n18310), .B1(n26130), .B2(
        data_in[6]), .ZN(n18316) );
  INV_X1 U14593 ( .A(n18317), .ZN(n8793) );
  AOI22_X1 U14594 ( .A1(\mem[1000][7] ), .A2(n18310), .B1(n26130), .B2(
        data_in[7]), .ZN(n18317) );
  INV_X1 U14595 ( .A(n18319), .ZN(n8792) );
  AOI22_X1 U14596 ( .A1(\mem[1001][0] ), .A2(n18320), .B1(n26129), .B2(
        data_in[0]), .ZN(n18319) );
  INV_X1 U14597 ( .A(n18321), .ZN(n8791) );
  AOI22_X1 U14598 ( .A1(\mem[1001][1] ), .A2(n18320), .B1(n26129), .B2(
        data_in[1]), .ZN(n18321) );
  INV_X1 U14599 ( .A(n18322), .ZN(n8790) );
  AOI22_X1 U14600 ( .A1(\mem[1001][2] ), .A2(n18320), .B1(n26129), .B2(
        data_in[2]), .ZN(n18322) );
  INV_X1 U14601 ( .A(n18323), .ZN(n8789) );
  AOI22_X1 U14602 ( .A1(\mem[1001][3] ), .A2(n18320), .B1(n26129), .B2(
        data_in[3]), .ZN(n18323) );
  INV_X1 U14603 ( .A(n18324), .ZN(n8788) );
  AOI22_X1 U14604 ( .A1(\mem[1001][4] ), .A2(n18320), .B1(n26129), .B2(
        data_in[4]), .ZN(n18324) );
  INV_X1 U14605 ( .A(n18325), .ZN(n8787) );
  AOI22_X1 U14606 ( .A1(\mem[1001][5] ), .A2(n18320), .B1(n26129), .B2(
        data_in[5]), .ZN(n18325) );
  INV_X1 U14607 ( .A(n18326), .ZN(n8786) );
  AOI22_X1 U14608 ( .A1(\mem[1001][6] ), .A2(n18320), .B1(n26129), .B2(
        data_in[6]), .ZN(n18326) );
  INV_X1 U14609 ( .A(n18327), .ZN(n8785) );
  AOI22_X1 U14610 ( .A1(\mem[1001][7] ), .A2(n18320), .B1(n26129), .B2(
        data_in[7]), .ZN(n18327) );
  INV_X1 U14611 ( .A(n18328), .ZN(n8784) );
  AOI22_X1 U14612 ( .A1(\mem[1002][0] ), .A2(n18329), .B1(n26128), .B2(
        data_in[0]), .ZN(n18328) );
  INV_X1 U14613 ( .A(n18330), .ZN(n8783) );
  AOI22_X1 U14614 ( .A1(\mem[1002][1] ), .A2(n18329), .B1(n26128), .B2(
        data_in[1]), .ZN(n18330) );
  INV_X1 U14615 ( .A(n18331), .ZN(n8782) );
  AOI22_X1 U14616 ( .A1(\mem[1002][2] ), .A2(n18329), .B1(n26128), .B2(
        data_in[2]), .ZN(n18331) );
  INV_X1 U14617 ( .A(n18332), .ZN(n8781) );
  AOI22_X1 U14618 ( .A1(\mem[1002][3] ), .A2(n18329), .B1(n26128), .B2(
        data_in[3]), .ZN(n18332) );
  INV_X1 U14619 ( .A(n18333), .ZN(n8780) );
  AOI22_X1 U14620 ( .A1(\mem[1002][4] ), .A2(n18329), .B1(n26128), .B2(
        data_in[4]), .ZN(n18333) );
  INV_X1 U14621 ( .A(n18334), .ZN(n8779) );
  AOI22_X1 U14622 ( .A1(\mem[1002][5] ), .A2(n18329), .B1(n26128), .B2(
        data_in[5]), .ZN(n18334) );
  INV_X1 U14623 ( .A(n18335), .ZN(n8778) );
  AOI22_X1 U14624 ( .A1(\mem[1002][6] ), .A2(n18329), .B1(n26128), .B2(
        data_in[6]), .ZN(n18335) );
  INV_X1 U14625 ( .A(n18336), .ZN(n8777) );
  AOI22_X1 U14626 ( .A1(\mem[1002][7] ), .A2(n18329), .B1(n26128), .B2(
        data_in[7]), .ZN(n18336) );
  INV_X1 U14627 ( .A(n18337), .ZN(n8776) );
  AOI22_X1 U14628 ( .A1(\mem[1003][0] ), .A2(n18338), .B1(n26127), .B2(
        data_in[0]), .ZN(n18337) );
  INV_X1 U14629 ( .A(n18339), .ZN(n8775) );
  AOI22_X1 U14630 ( .A1(\mem[1003][1] ), .A2(n18338), .B1(n26127), .B2(
        data_in[1]), .ZN(n18339) );
  INV_X1 U14631 ( .A(n18340), .ZN(n8774) );
  AOI22_X1 U14632 ( .A1(\mem[1003][2] ), .A2(n18338), .B1(n26127), .B2(
        data_in[2]), .ZN(n18340) );
  INV_X1 U14633 ( .A(n18341), .ZN(n8773) );
  AOI22_X1 U14634 ( .A1(\mem[1003][3] ), .A2(n18338), .B1(n26127), .B2(
        data_in[3]), .ZN(n18341) );
  INV_X1 U14635 ( .A(n18342), .ZN(n8772) );
  AOI22_X1 U14636 ( .A1(\mem[1003][4] ), .A2(n18338), .B1(n26127), .B2(
        data_in[4]), .ZN(n18342) );
  INV_X1 U14637 ( .A(n18343), .ZN(n8771) );
  AOI22_X1 U14638 ( .A1(\mem[1003][5] ), .A2(n18338), .B1(n26127), .B2(
        data_in[5]), .ZN(n18343) );
  INV_X1 U14639 ( .A(n18344), .ZN(n8770) );
  AOI22_X1 U14640 ( .A1(\mem[1003][6] ), .A2(n18338), .B1(n26127), .B2(
        data_in[6]), .ZN(n18344) );
  INV_X1 U14641 ( .A(n18345), .ZN(n8769) );
  AOI22_X1 U14642 ( .A1(\mem[1003][7] ), .A2(n18338), .B1(n26127), .B2(
        data_in[7]), .ZN(n18345) );
  INV_X1 U14643 ( .A(n18346), .ZN(n8768) );
  AOI22_X1 U14644 ( .A1(\mem[1004][0] ), .A2(n18347), .B1(n26126), .B2(
        data_in[0]), .ZN(n18346) );
  INV_X1 U14645 ( .A(n18348), .ZN(n8767) );
  AOI22_X1 U14646 ( .A1(\mem[1004][1] ), .A2(n18347), .B1(n26126), .B2(
        data_in[1]), .ZN(n18348) );
  INV_X1 U14647 ( .A(n18349), .ZN(n8766) );
  AOI22_X1 U14648 ( .A1(\mem[1004][2] ), .A2(n18347), .B1(n26126), .B2(
        data_in[2]), .ZN(n18349) );
  INV_X1 U14649 ( .A(n18350), .ZN(n8765) );
  AOI22_X1 U14650 ( .A1(\mem[1004][3] ), .A2(n18347), .B1(n26126), .B2(
        data_in[3]), .ZN(n18350) );
  INV_X1 U14651 ( .A(n18351), .ZN(n8764) );
  AOI22_X1 U14652 ( .A1(\mem[1004][4] ), .A2(n18347), .B1(n26126), .B2(
        data_in[4]), .ZN(n18351) );
  INV_X1 U14653 ( .A(n18352), .ZN(n8763) );
  AOI22_X1 U14654 ( .A1(\mem[1004][5] ), .A2(n18347), .B1(n26126), .B2(
        data_in[5]), .ZN(n18352) );
  INV_X1 U14655 ( .A(n18353), .ZN(n8762) );
  AOI22_X1 U14656 ( .A1(\mem[1004][6] ), .A2(n18347), .B1(n26126), .B2(
        data_in[6]), .ZN(n18353) );
  INV_X1 U14657 ( .A(n18354), .ZN(n8761) );
  AOI22_X1 U14658 ( .A1(\mem[1004][7] ), .A2(n18347), .B1(n26126), .B2(
        data_in[7]), .ZN(n18354) );
  INV_X1 U14659 ( .A(n18355), .ZN(n8760) );
  AOI22_X1 U14660 ( .A1(\mem[1005][0] ), .A2(n18356), .B1(n26125), .B2(
        data_in[0]), .ZN(n18355) );
  INV_X1 U14661 ( .A(n18357), .ZN(n8759) );
  AOI22_X1 U14662 ( .A1(\mem[1005][1] ), .A2(n18356), .B1(n26125), .B2(
        data_in[1]), .ZN(n18357) );
  INV_X1 U14663 ( .A(n18358), .ZN(n8758) );
  AOI22_X1 U14664 ( .A1(\mem[1005][2] ), .A2(n18356), .B1(n26125), .B2(
        data_in[2]), .ZN(n18358) );
  INV_X1 U14665 ( .A(n18359), .ZN(n8757) );
  AOI22_X1 U14666 ( .A1(\mem[1005][3] ), .A2(n18356), .B1(n26125), .B2(
        data_in[3]), .ZN(n18359) );
  INV_X1 U14667 ( .A(n18360), .ZN(n8756) );
  AOI22_X1 U14668 ( .A1(\mem[1005][4] ), .A2(n18356), .B1(n26125), .B2(
        data_in[4]), .ZN(n18360) );
  INV_X1 U14669 ( .A(n18361), .ZN(n8755) );
  AOI22_X1 U14670 ( .A1(\mem[1005][5] ), .A2(n18356), .B1(n26125), .B2(
        data_in[5]), .ZN(n18361) );
  INV_X1 U14671 ( .A(n18362), .ZN(n8754) );
  AOI22_X1 U14672 ( .A1(\mem[1005][6] ), .A2(n18356), .B1(n26125), .B2(
        data_in[6]), .ZN(n18362) );
  INV_X1 U14673 ( .A(n18363), .ZN(n8753) );
  AOI22_X1 U14674 ( .A1(\mem[1005][7] ), .A2(n18356), .B1(n26125), .B2(
        data_in[7]), .ZN(n18363) );
  INV_X1 U14675 ( .A(n18364), .ZN(n8752) );
  AOI22_X1 U14676 ( .A1(\mem[1006][0] ), .A2(n18365), .B1(n26124), .B2(
        data_in[0]), .ZN(n18364) );
  INV_X1 U14677 ( .A(n18366), .ZN(n8751) );
  AOI22_X1 U14678 ( .A1(\mem[1006][1] ), .A2(n18365), .B1(n26124), .B2(
        data_in[1]), .ZN(n18366) );
  INV_X1 U14679 ( .A(n18367), .ZN(n8750) );
  AOI22_X1 U14680 ( .A1(\mem[1006][2] ), .A2(n18365), .B1(n26124), .B2(
        data_in[2]), .ZN(n18367) );
  INV_X1 U14681 ( .A(n18368), .ZN(n8749) );
  AOI22_X1 U14682 ( .A1(\mem[1006][3] ), .A2(n18365), .B1(n26124), .B2(
        data_in[3]), .ZN(n18368) );
  INV_X1 U14683 ( .A(n18369), .ZN(n8748) );
  AOI22_X1 U14684 ( .A1(\mem[1006][4] ), .A2(n18365), .B1(n26124), .B2(
        data_in[4]), .ZN(n18369) );
  INV_X1 U14685 ( .A(n18370), .ZN(n8747) );
  AOI22_X1 U14686 ( .A1(\mem[1006][5] ), .A2(n18365), .B1(n26124), .B2(
        data_in[5]), .ZN(n18370) );
  INV_X1 U14687 ( .A(n18371), .ZN(n8746) );
  AOI22_X1 U14688 ( .A1(\mem[1006][6] ), .A2(n18365), .B1(n26124), .B2(
        data_in[6]), .ZN(n18371) );
  INV_X1 U14689 ( .A(n18372), .ZN(n8745) );
  AOI22_X1 U14690 ( .A1(\mem[1006][7] ), .A2(n18365), .B1(n26124), .B2(
        data_in[7]), .ZN(n18372) );
  INV_X1 U14691 ( .A(n18373), .ZN(n8744) );
  AOI22_X1 U14692 ( .A1(\mem[1007][0] ), .A2(n18374), .B1(n26123), .B2(
        data_in[0]), .ZN(n18373) );
  INV_X1 U14693 ( .A(n18375), .ZN(n8743) );
  AOI22_X1 U14694 ( .A1(\mem[1007][1] ), .A2(n18374), .B1(n26123), .B2(
        data_in[1]), .ZN(n18375) );
  INV_X1 U14695 ( .A(n18376), .ZN(n8742) );
  AOI22_X1 U14696 ( .A1(\mem[1007][2] ), .A2(n18374), .B1(n26123), .B2(
        data_in[2]), .ZN(n18376) );
  INV_X1 U14697 ( .A(n18377), .ZN(n8741) );
  AOI22_X1 U14698 ( .A1(\mem[1007][3] ), .A2(n18374), .B1(n26123), .B2(
        data_in[3]), .ZN(n18377) );
  INV_X1 U14699 ( .A(n18378), .ZN(n8740) );
  AOI22_X1 U14700 ( .A1(\mem[1007][4] ), .A2(n18374), .B1(n26123), .B2(
        data_in[4]), .ZN(n18378) );
  INV_X1 U14701 ( .A(n18379), .ZN(n8739) );
  AOI22_X1 U14702 ( .A1(\mem[1007][5] ), .A2(n18374), .B1(n26123), .B2(
        data_in[5]), .ZN(n18379) );
  INV_X1 U14703 ( .A(n18380), .ZN(n8738) );
  AOI22_X1 U14704 ( .A1(\mem[1007][6] ), .A2(n18374), .B1(n26123), .B2(
        data_in[6]), .ZN(n18380) );
  INV_X1 U14705 ( .A(n18381), .ZN(n8737) );
  AOI22_X1 U14706 ( .A1(\mem[1007][7] ), .A2(n18374), .B1(n26123), .B2(
        data_in[7]), .ZN(n18381) );
  INV_X1 U14707 ( .A(n18382), .ZN(n8736) );
  AOI22_X1 U14708 ( .A1(\mem[1008][0] ), .A2(n18383), .B1(n26122), .B2(
        data_in[0]), .ZN(n18382) );
  INV_X1 U14709 ( .A(n18384), .ZN(n8735) );
  AOI22_X1 U14710 ( .A1(\mem[1008][1] ), .A2(n18383), .B1(n26122), .B2(
        data_in[1]), .ZN(n18384) );
  INV_X1 U14711 ( .A(n18385), .ZN(n8734) );
  AOI22_X1 U14712 ( .A1(\mem[1008][2] ), .A2(n18383), .B1(n26122), .B2(
        data_in[2]), .ZN(n18385) );
  INV_X1 U14713 ( .A(n18386), .ZN(n8733) );
  AOI22_X1 U14714 ( .A1(\mem[1008][3] ), .A2(n18383), .B1(n26122), .B2(
        data_in[3]), .ZN(n18386) );
  INV_X1 U14715 ( .A(n18387), .ZN(n8732) );
  AOI22_X1 U14716 ( .A1(\mem[1008][4] ), .A2(n18383), .B1(n26122), .B2(
        data_in[4]), .ZN(n18387) );
  INV_X1 U14717 ( .A(n18388), .ZN(n8731) );
  AOI22_X1 U14718 ( .A1(\mem[1008][5] ), .A2(n18383), .B1(n26122), .B2(
        data_in[5]), .ZN(n18388) );
  INV_X1 U14719 ( .A(n18389), .ZN(n8730) );
  AOI22_X1 U14720 ( .A1(\mem[1008][6] ), .A2(n18383), .B1(n26122), .B2(
        data_in[6]), .ZN(n18389) );
  INV_X1 U14721 ( .A(n18390), .ZN(n8729) );
  AOI22_X1 U14722 ( .A1(\mem[1008][7] ), .A2(n18383), .B1(n26122), .B2(
        data_in[7]), .ZN(n18390) );
  INV_X1 U14723 ( .A(n18392), .ZN(n8728) );
  AOI22_X1 U14724 ( .A1(\mem[1009][0] ), .A2(n18393), .B1(n26121), .B2(
        data_in[0]), .ZN(n18392) );
  INV_X1 U14725 ( .A(n18394), .ZN(n8727) );
  AOI22_X1 U14726 ( .A1(\mem[1009][1] ), .A2(n18393), .B1(n26121), .B2(
        data_in[1]), .ZN(n18394) );
  INV_X1 U14727 ( .A(n18395), .ZN(n8726) );
  AOI22_X1 U14728 ( .A1(\mem[1009][2] ), .A2(n18393), .B1(n26121), .B2(
        data_in[2]), .ZN(n18395) );
  INV_X1 U14729 ( .A(n18396), .ZN(n8725) );
  AOI22_X1 U14730 ( .A1(\mem[1009][3] ), .A2(n18393), .B1(n26121), .B2(
        data_in[3]), .ZN(n18396) );
  INV_X1 U14731 ( .A(n18397), .ZN(n8724) );
  AOI22_X1 U14732 ( .A1(\mem[1009][4] ), .A2(n18393), .B1(n26121), .B2(
        data_in[4]), .ZN(n18397) );
  INV_X1 U14733 ( .A(n18398), .ZN(n8723) );
  AOI22_X1 U14734 ( .A1(\mem[1009][5] ), .A2(n18393), .B1(n26121), .B2(
        data_in[5]), .ZN(n18398) );
  INV_X1 U14735 ( .A(n18399), .ZN(n8722) );
  AOI22_X1 U14736 ( .A1(\mem[1009][6] ), .A2(n18393), .B1(n26121), .B2(
        data_in[6]), .ZN(n18399) );
  INV_X1 U14737 ( .A(n18400), .ZN(n8721) );
  AOI22_X1 U14738 ( .A1(\mem[1009][7] ), .A2(n18393), .B1(n26121), .B2(
        data_in[7]), .ZN(n18400) );
  INV_X1 U14739 ( .A(n18401), .ZN(n8720) );
  AOI22_X1 U14740 ( .A1(\mem[1010][0] ), .A2(n18402), .B1(n26120), .B2(
        data_in[0]), .ZN(n18401) );
  INV_X1 U14741 ( .A(n18403), .ZN(n8719) );
  AOI22_X1 U14742 ( .A1(\mem[1010][1] ), .A2(n18402), .B1(n26120), .B2(
        data_in[1]), .ZN(n18403) );
  INV_X1 U14743 ( .A(n18404), .ZN(n8718) );
  AOI22_X1 U14744 ( .A1(\mem[1010][2] ), .A2(n18402), .B1(n26120), .B2(
        data_in[2]), .ZN(n18404) );
  INV_X1 U14745 ( .A(n18405), .ZN(n8717) );
  AOI22_X1 U14746 ( .A1(\mem[1010][3] ), .A2(n18402), .B1(n26120), .B2(
        data_in[3]), .ZN(n18405) );
  INV_X1 U14747 ( .A(n18406), .ZN(n8716) );
  AOI22_X1 U14748 ( .A1(\mem[1010][4] ), .A2(n18402), .B1(n26120), .B2(
        data_in[4]), .ZN(n18406) );
  INV_X1 U14749 ( .A(n18407), .ZN(n8715) );
  AOI22_X1 U14750 ( .A1(\mem[1010][5] ), .A2(n18402), .B1(n26120), .B2(
        data_in[5]), .ZN(n18407) );
  INV_X1 U14751 ( .A(n18408), .ZN(n8714) );
  AOI22_X1 U14752 ( .A1(\mem[1010][6] ), .A2(n18402), .B1(n26120), .B2(
        data_in[6]), .ZN(n18408) );
  INV_X1 U14753 ( .A(n18409), .ZN(n8713) );
  AOI22_X1 U14754 ( .A1(\mem[1010][7] ), .A2(n18402), .B1(n26120), .B2(
        data_in[7]), .ZN(n18409) );
  INV_X1 U14755 ( .A(n18410), .ZN(n8712) );
  AOI22_X1 U14756 ( .A1(\mem[1011][0] ), .A2(n18411), .B1(n26119), .B2(
        data_in[0]), .ZN(n18410) );
  INV_X1 U14757 ( .A(n18412), .ZN(n8711) );
  AOI22_X1 U14758 ( .A1(\mem[1011][1] ), .A2(n18411), .B1(n26119), .B2(
        data_in[1]), .ZN(n18412) );
  INV_X1 U14759 ( .A(n18413), .ZN(n8710) );
  AOI22_X1 U14760 ( .A1(\mem[1011][2] ), .A2(n18411), .B1(n26119), .B2(
        data_in[2]), .ZN(n18413) );
  INV_X1 U14761 ( .A(n18414), .ZN(n8709) );
  AOI22_X1 U14762 ( .A1(\mem[1011][3] ), .A2(n18411), .B1(n26119), .B2(
        data_in[3]), .ZN(n18414) );
  INV_X1 U14763 ( .A(n18415), .ZN(n8708) );
  AOI22_X1 U14764 ( .A1(\mem[1011][4] ), .A2(n18411), .B1(n26119), .B2(
        data_in[4]), .ZN(n18415) );
  INV_X1 U14765 ( .A(n18416), .ZN(n8707) );
  AOI22_X1 U14766 ( .A1(\mem[1011][5] ), .A2(n18411), .B1(n26119), .B2(
        data_in[5]), .ZN(n18416) );
  INV_X1 U14767 ( .A(n18417), .ZN(n8706) );
  AOI22_X1 U14768 ( .A1(\mem[1011][6] ), .A2(n18411), .B1(n26119), .B2(
        data_in[6]), .ZN(n18417) );
  INV_X1 U14769 ( .A(n18418), .ZN(n8705) );
  AOI22_X1 U14770 ( .A1(\mem[1011][7] ), .A2(n18411), .B1(n26119), .B2(
        data_in[7]), .ZN(n18418) );
  INV_X1 U14771 ( .A(n18419), .ZN(n8704) );
  AOI22_X1 U14772 ( .A1(\mem[1012][0] ), .A2(n18420), .B1(n26118), .B2(
        data_in[0]), .ZN(n18419) );
  INV_X1 U14773 ( .A(n18421), .ZN(n8703) );
  AOI22_X1 U14774 ( .A1(\mem[1012][1] ), .A2(n18420), .B1(n26118), .B2(
        data_in[1]), .ZN(n18421) );
  INV_X1 U14775 ( .A(n18422), .ZN(n8702) );
  AOI22_X1 U14776 ( .A1(\mem[1012][2] ), .A2(n18420), .B1(n26118), .B2(
        data_in[2]), .ZN(n18422) );
  INV_X1 U14777 ( .A(n18423), .ZN(n8701) );
  AOI22_X1 U14778 ( .A1(\mem[1012][3] ), .A2(n18420), .B1(n26118), .B2(
        data_in[3]), .ZN(n18423) );
  INV_X1 U14779 ( .A(n18424), .ZN(n8700) );
  AOI22_X1 U14780 ( .A1(\mem[1012][4] ), .A2(n18420), .B1(n26118), .B2(
        data_in[4]), .ZN(n18424) );
  INV_X1 U14781 ( .A(n18425), .ZN(n8699) );
  AOI22_X1 U14782 ( .A1(\mem[1012][5] ), .A2(n18420), .B1(n26118), .B2(
        data_in[5]), .ZN(n18425) );
  INV_X1 U14783 ( .A(n18426), .ZN(n8698) );
  AOI22_X1 U14784 ( .A1(\mem[1012][6] ), .A2(n18420), .B1(n26118), .B2(
        data_in[6]), .ZN(n18426) );
  INV_X1 U14785 ( .A(n18427), .ZN(n8697) );
  AOI22_X1 U14786 ( .A1(\mem[1012][7] ), .A2(n18420), .B1(n26118), .B2(
        data_in[7]), .ZN(n18427) );
  INV_X1 U14787 ( .A(n18428), .ZN(n8696) );
  AOI22_X1 U14788 ( .A1(\mem[1013][0] ), .A2(n18429), .B1(n26117), .B2(
        data_in[0]), .ZN(n18428) );
  INV_X1 U14789 ( .A(n18430), .ZN(n8695) );
  AOI22_X1 U14790 ( .A1(\mem[1013][1] ), .A2(n18429), .B1(n26117), .B2(
        data_in[1]), .ZN(n18430) );
  INV_X1 U14791 ( .A(n18431), .ZN(n8694) );
  AOI22_X1 U14792 ( .A1(\mem[1013][2] ), .A2(n18429), .B1(n26117), .B2(
        data_in[2]), .ZN(n18431) );
  INV_X1 U14793 ( .A(n18432), .ZN(n8693) );
  AOI22_X1 U14794 ( .A1(\mem[1013][3] ), .A2(n18429), .B1(n26117), .B2(
        data_in[3]), .ZN(n18432) );
  INV_X1 U14795 ( .A(n18433), .ZN(n8692) );
  AOI22_X1 U14796 ( .A1(\mem[1013][4] ), .A2(n18429), .B1(n26117), .B2(
        data_in[4]), .ZN(n18433) );
  INV_X1 U14797 ( .A(n18434), .ZN(n8691) );
  AOI22_X1 U14798 ( .A1(\mem[1013][5] ), .A2(n18429), .B1(n26117), .B2(
        data_in[5]), .ZN(n18434) );
  INV_X1 U14799 ( .A(n18435), .ZN(n8690) );
  AOI22_X1 U14800 ( .A1(\mem[1013][6] ), .A2(n18429), .B1(n26117), .B2(
        data_in[6]), .ZN(n18435) );
  INV_X1 U14801 ( .A(n18436), .ZN(n8689) );
  AOI22_X1 U14802 ( .A1(\mem[1013][7] ), .A2(n18429), .B1(n26117), .B2(
        data_in[7]), .ZN(n18436) );
  INV_X1 U14803 ( .A(n18437), .ZN(n8688) );
  AOI22_X1 U14804 ( .A1(\mem[1014][0] ), .A2(n18438), .B1(n26116), .B2(
        data_in[0]), .ZN(n18437) );
  INV_X1 U14805 ( .A(n18439), .ZN(n8687) );
  AOI22_X1 U14806 ( .A1(\mem[1014][1] ), .A2(n18438), .B1(n26116), .B2(
        data_in[1]), .ZN(n18439) );
  INV_X1 U14807 ( .A(n18440), .ZN(n8686) );
  AOI22_X1 U14808 ( .A1(\mem[1014][2] ), .A2(n18438), .B1(n26116), .B2(
        data_in[2]), .ZN(n18440) );
  INV_X1 U14809 ( .A(n18441), .ZN(n8685) );
  AOI22_X1 U14810 ( .A1(\mem[1014][3] ), .A2(n18438), .B1(n26116), .B2(
        data_in[3]), .ZN(n18441) );
  INV_X1 U14811 ( .A(n18442), .ZN(n8684) );
  AOI22_X1 U14812 ( .A1(\mem[1014][4] ), .A2(n18438), .B1(n26116), .B2(
        data_in[4]), .ZN(n18442) );
  INV_X1 U14813 ( .A(n18443), .ZN(n8683) );
  AOI22_X1 U14814 ( .A1(\mem[1014][5] ), .A2(n18438), .B1(n26116), .B2(
        data_in[5]), .ZN(n18443) );
  INV_X1 U14815 ( .A(n18444), .ZN(n8682) );
  AOI22_X1 U14816 ( .A1(\mem[1014][6] ), .A2(n18438), .B1(n26116), .B2(
        data_in[6]), .ZN(n18444) );
  INV_X1 U14817 ( .A(n18445), .ZN(n8681) );
  AOI22_X1 U14818 ( .A1(\mem[1014][7] ), .A2(n18438), .B1(n26116), .B2(
        data_in[7]), .ZN(n18445) );
  INV_X1 U14819 ( .A(n18446), .ZN(n8680) );
  AOI22_X1 U14820 ( .A1(\mem[1015][0] ), .A2(n18447), .B1(n26115), .B2(
        data_in[0]), .ZN(n18446) );
  INV_X1 U14821 ( .A(n18448), .ZN(n8679) );
  AOI22_X1 U14822 ( .A1(\mem[1015][1] ), .A2(n18447), .B1(n26115), .B2(
        data_in[1]), .ZN(n18448) );
  INV_X1 U14823 ( .A(n18449), .ZN(n8678) );
  AOI22_X1 U14824 ( .A1(\mem[1015][2] ), .A2(n18447), .B1(n26115), .B2(
        data_in[2]), .ZN(n18449) );
  INV_X1 U14825 ( .A(n18450), .ZN(n8677) );
  AOI22_X1 U14826 ( .A1(\mem[1015][3] ), .A2(n18447), .B1(n26115), .B2(
        data_in[3]), .ZN(n18450) );
  INV_X1 U14827 ( .A(n18451), .ZN(n8676) );
  AOI22_X1 U14828 ( .A1(\mem[1015][4] ), .A2(n18447), .B1(n26115), .B2(
        data_in[4]), .ZN(n18451) );
  INV_X1 U14829 ( .A(n18452), .ZN(n8675) );
  AOI22_X1 U14830 ( .A1(\mem[1015][5] ), .A2(n18447), .B1(n26115), .B2(
        data_in[5]), .ZN(n18452) );
  INV_X1 U14831 ( .A(n18453), .ZN(n8674) );
  AOI22_X1 U14832 ( .A1(\mem[1015][6] ), .A2(n18447), .B1(n26115), .B2(
        data_in[6]), .ZN(n18453) );
  INV_X1 U14833 ( .A(n18454), .ZN(n8673) );
  AOI22_X1 U14834 ( .A1(\mem[1015][7] ), .A2(n18447), .B1(n26115), .B2(
        data_in[7]), .ZN(n18454) );
  INV_X1 U14835 ( .A(n18455), .ZN(n8672) );
  AOI22_X1 U14836 ( .A1(\mem[1016][0] ), .A2(n18456), .B1(n26114), .B2(
        data_in[0]), .ZN(n18455) );
  INV_X1 U14837 ( .A(n18457), .ZN(n8671) );
  AOI22_X1 U14838 ( .A1(\mem[1016][1] ), .A2(n18456), .B1(n26114), .B2(
        data_in[1]), .ZN(n18457) );
  INV_X1 U14839 ( .A(n18458), .ZN(n8670) );
  AOI22_X1 U14840 ( .A1(\mem[1016][2] ), .A2(n18456), .B1(n26114), .B2(
        data_in[2]), .ZN(n18458) );
  INV_X1 U14841 ( .A(n18459), .ZN(n8669) );
  AOI22_X1 U14842 ( .A1(\mem[1016][3] ), .A2(n18456), .B1(n26114), .B2(
        data_in[3]), .ZN(n18459) );
  INV_X1 U14843 ( .A(n18460), .ZN(n8668) );
  AOI22_X1 U14844 ( .A1(\mem[1016][4] ), .A2(n18456), .B1(n26114), .B2(
        data_in[4]), .ZN(n18460) );
  INV_X1 U14845 ( .A(n18461), .ZN(n8667) );
  AOI22_X1 U14846 ( .A1(\mem[1016][5] ), .A2(n18456), .B1(n26114), .B2(
        data_in[5]), .ZN(n18461) );
  INV_X1 U14847 ( .A(n18462), .ZN(n8666) );
  AOI22_X1 U14848 ( .A1(\mem[1016][6] ), .A2(n18456), .B1(n26114), .B2(
        data_in[6]), .ZN(n18462) );
  INV_X1 U14849 ( .A(n18463), .ZN(n8665) );
  AOI22_X1 U14850 ( .A1(\mem[1016][7] ), .A2(n18456), .B1(n26114), .B2(
        data_in[7]), .ZN(n18463) );
  INV_X1 U14851 ( .A(n18465), .ZN(n8664) );
  AOI22_X1 U14852 ( .A1(\mem[1017][0] ), .A2(n18466), .B1(n26113), .B2(
        data_in[0]), .ZN(n18465) );
  INV_X1 U14853 ( .A(n18467), .ZN(n8663) );
  AOI22_X1 U14854 ( .A1(\mem[1017][1] ), .A2(n18466), .B1(n26113), .B2(
        data_in[1]), .ZN(n18467) );
  INV_X1 U14855 ( .A(n18468), .ZN(n8662) );
  AOI22_X1 U14856 ( .A1(\mem[1017][2] ), .A2(n18466), .B1(n26113), .B2(
        data_in[2]), .ZN(n18468) );
  INV_X1 U14857 ( .A(n18469), .ZN(n8661) );
  AOI22_X1 U14858 ( .A1(\mem[1017][3] ), .A2(n18466), .B1(n26113), .B2(
        data_in[3]), .ZN(n18469) );
  INV_X1 U14859 ( .A(n18470), .ZN(n8660) );
  AOI22_X1 U14860 ( .A1(\mem[1017][4] ), .A2(n18466), .B1(n26113), .B2(
        data_in[4]), .ZN(n18470) );
  INV_X1 U14861 ( .A(n18471), .ZN(n8659) );
  AOI22_X1 U14862 ( .A1(\mem[1017][5] ), .A2(n18466), .B1(n26113), .B2(
        data_in[5]), .ZN(n18471) );
  INV_X1 U14863 ( .A(n18472), .ZN(n8658) );
  AOI22_X1 U14864 ( .A1(\mem[1017][6] ), .A2(n18466), .B1(n26113), .B2(
        data_in[6]), .ZN(n18472) );
  INV_X1 U14865 ( .A(n18473), .ZN(n8657) );
  AOI22_X1 U14866 ( .A1(\mem[1017][7] ), .A2(n18466), .B1(n26113), .B2(
        data_in[7]), .ZN(n18473) );
  INV_X1 U14867 ( .A(n18474), .ZN(n8656) );
  AOI22_X1 U14868 ( .A1(\mem[1018][0] ), .A2(n18475), .B1(n26112), .B2(
        data_in[0]), .ZN(n18474) );
  INV_X1 U14869 ( .A(n18476), .ZN(n8655) );
  AOI22_X1 U14870 ( .A1(\mem[1018][1] ), .A2(n18475), .B1(n26112), .B2(
        data_in[1]), .ZN(n18476) );
  INV_X1 U14871 ( .A(n18477), .ZN(n8654) );
  AOI22_X1 U14872 ( .A1(\mem[1018][2] ), .A2(n18475), .B1(n26112), .B2(
        data_in[2]), .ZN(n18477) );
  INV_X1 U14873 ( .A(n18478), .ZN(n8653) );
  AOI22_X1 U14874 ( .A1(\mem[1018][3] ), .A2(n18475), .B1(n26112), .B2(
        data_in[3]), .ZN(n18478) );
  INV_X1 U14875 ( .A(n18479), .ZN(n8652) );
  AOI22_X1 U14876 ( .A1(\mem[1018][4] ), .A2(n18475), .B1(n26112), .B2(
        data_in[4]), .ZN(n18479) );
  INV_X1 U14877 ( .A(n18480), .ZN(n8651) );
  AOI22_X1 U14878 ( .A1(\mem[1018][5] ), .A2(n18475), .B1(n26112), .B2(
        data_in[5]), .ZN(n18480) );
  INV_X1 U14879 ( .A(n18481), .ZN(n8650) );
  AOI22_X1 U14880 ( .A1(\mem[1018][6] ), .A2(n18475), .B1(n26112), .B2(
        data_in[6]), .ZN(n18481) );
  INV_X1 U14881 ( .A(n18482), .ZN(n8649) );
  AOI22_X1 U14882 ( .A1(\mem[1018][7] ), .A2(n18475), .B1(n26112), .B2(
        data_in[7]), .ZN(n18482) );
  INV_X1 U14883 ( .A(n18483), .ZN(n8648) );
  AOI22_X1 U14884 ( .A1(\mem[1019][0] ), .A2(n18484), .B1(n26111), .B2(
        data_in[0]), .ZN(n18483) );
  INV_X1 U14885 ( .A(n18485), .ZN(n8647) );
  AOI22_X1 U14886 ( .A1(\mem[1019][1] ), .A2(n18484), .B1(n26111), .B2(
        data_in[1]), .ZN(n18485) );
  INV_X1 U14887 ( .A(n18486), .ZN(n8646) );
  AOI22_X1 U14888 ( .A1(\mem[1019][2] ), .A2(n18484), .B1(n26111), .B2(
        data_in[2]), .ZN(n18486) );
  INV_X1 U14889 ( .A(n18487), .ZN(n8645) );
  AOI22_X1 U14890 ( .A1(\mem[1019][3] ), .A2(n18484), .B1(n26111), .B2(
        data_in[3]), .ZN(n18487) );
  INV_X1 U14891 ( .A(n18488), .ZN(n8644) );
  AOI22_X1 U14892 ( .A1(\mem[1019][4] ), .A2(n18484), .B1(n26111), .B2(
        data_in[4]), .ZN(n18488) );
  INV_X1 U14893 ( .A(n18489), .ZN(n8643) );
  AOI22_X1 U14894 ( .A1(\mem[1019][5] ), .A2(n18484), .B1(n26111), .B2(
        data_in[5]), .ZN(n18489) );
  INV_X1 U14895 ( .A(n18490), .ZN(n8642) );
  AOI22_X1 U14896 ( .A1(\mem[1019][6] ), .A2(n18484), .B1(n26111), .B2(
        data_in[6]), .ZN(n18490) );
  INV_X1 U14897 ( .A(n18491), .ZN(n8641) );
  AOI22_X1 U14898 ( .A1(\mem[1019][7] ), .A2(n18484), .B1(n26111), .B2(
        data_in[7]), .ZN(n18491) );
  INV_X1 U14899 ( .A(n18492), .ZN(n8640) );
  AOI22_X1 U14900 ( .A1(\mem[1020][0] ), .A2(n18493), .B1(n26110), .B2(
        data_in[0]), .ZN(n18492) );
  INV_X1 U14901 ( .A(n18494), .ZN(n8639) );
  AOI22_X1 U14902 ( .A1(\mem[1020][1] ), .A2(n18493), .B1(n26110), .B2(
        data_in[1]), .ZN(n18494) );
  INV_X1 U14903 ( .A(n18495), .ZN(n8638) );
  AOI22_X1 U14904 ( .A1(\mem[1020][2] ), .A2(n18493), .B1(n26110), .B2(
        data_in[2]), .ZN(n18495) );
  INV_X1 U14905 ( .A(n18496), .ZN(n8637) );
  AOI22_X1 U14906 ( .A1(\mem[1020][3] ), .A2(n18493), .B1(n26110), .B2(
        data_in[3]), .ZN(n18496) );
  INV_X1 U14907 ( .A(n18497), .ZN(n8636) );
  AOI22_X1 U14908 ( .A1(\mem[1020][4] ), .A2(n18493), .B1(n26110), .B2(
        data_in[4]), .ZN(n18497) );
  INV_X1 U14909 ( .A(n18498), .ZN(n8635) );
  AOI22_X1 U14910 ( .A1(\mem[1020][5] ), .A2(n18493), .B1(n26110), .B2(
        data_in[5]), .ZN(n18498) );
  INV_X1 U14911 ( .A(n18499), .ZN(n8634) );
  AOI22_X1 U14912 ( .A1(\mem[1020][6] ), .A2(n18493), .B1(n26110), .B2(
        data_in[6]), .ZN(n18499) );
  INV_X1 U14913 ( .A(n18500), .ZN(n8633) );
  AOI22_X1 U14914 ( .A1(\mem[1020][7] ), .A2(n18493), .B1(n26110), .B2(
        data_in[7]), .ZN(n18500) );
  INV_X1 U14915 ( .A(n18501), .ZN(n8632) );
  AOI22_X1 U14916 ( .A1(\mem[1021][0] ), .A2(n18502), .B1(n26109), .B2(
        data_in[0]), .ZN(n18501) );
  INV_X1 U14917 ( .A(n18503), .ZN(n8631) );
  AOI22_X1 U14918 ( .A1(\mem[1021][1] ), .A2(n18502), .B1(n26109), .B2(
        data_in[1]), .ZN(n18503) );
  INV_X1 U14919 ( .A(n18504), .ZN(n8630) );
  AOI22_X1 U14920 ( .A1(\mem[1021][2] ), .A2(n18502), .B1(n26109), .B2(
        data_in[2]), .ZN(n18504) );
  INV_X1 U14921 ( .A(n18505), .ZN(n8629) );
  AOI22_X1 U14922 ( .A1(\mem[1021][3] ), .A2(n18502), .B1(n26109), .B2(
        data_in[3]), .ZN(n18505) );
  INV_X1 U14923 ( .A(n18506), .ZN(n8628) );
  AOI22_X1 U14924 ( .A1(\mem[1021][4] ), .A2(n18502), .B1(n26109), .B2(
        data_in[4]), .ZN(n18506) );
  INV_X1 U14925 ( .A(n18507), .ZN(n8627) );
  AOI22_X1 U14926 ( .A1(\mem[1021][5] ), .A2(n18502), .B1(n26109), .B2(
        data_in[5]), .ZN(n18507) );
  INV_X1 U14927 ( .A(n18508), .ZN(n8626) );
  AOI22_X1 U14928 ( .A1(\mem[1021][6] ), .A2(n18502), .B1(n26109), .B2(
        data_in[6]), .ZN(n18508) );
  INV_X1 U14929 ( .A(n18509), .ZN(n8625) );
  AOI22_X1 U14930 ( .A1(\mem[1021][7] ), .A2(n18502), .B1(n26109), .B2(
        data_in[7]), .ZN(n18509) );
  INV_X1 U14931 ( .A(n18510), .ZN(n8624) );
  AOI22_X1 U14932 ( .A1(\mem[1022][0] ), .A2(n18511), .B1(n26108), .B2(
        data_in[0]), .ZN(n18510) );
  INV_X1 U14933 ( .A(n18512), .ZN(n8623) );
  AOI22_X1 U14934 ( .A1(\mem[1022][1] ), .A2(n18511), .B1(n26108), .B2(
        data_in[1]), .ZN(n18512) );
  INV_X1 U14935 ( .A(n18513), .ZN(n8622) );
  AOI22_X1 U14936 ( .A1(\mem[1022][2] ), .A2(n18511), .B1(n26108), .B2(
        data_in[2]), .ZN(n18513) );
  INV_X1 U14937 ( .A(n18514), .ZN(n8621) );
  AOI22_X1 U14938 ( .A1(\mem[1022][3] ), .A2(n18511), .B1(n26108), .B2(
        data_in[3]), .ZN(n18514) );
  INV_X1 U14939 ( .A(n18515), .ZN(n8620) );
  AOI22_X1 U14940 ( .A1(\mem[1022][4] ), .A2(n18511), .B1(n26108), .B2(
        data_in[4]), .ZN(n18515) );
  INV_X1 U14941 ( .A(n18516), .ZN(n8619) );
  AOI22_X1 U14942 ( .A1(\mem[1022][5] ), .A2(n18511), .B1(n26108), .B2(
        data_in[5]), .ZN(n18516) );
  INV_X1 U14943 ( .A(n18517), .ZN(n8618) );
  AOI22_X1 U14944 ( .A1(\mem[1022][6] ), .A2(n18511), .B1(n26108), .B2(
        data_in[6]), .ZN(n18517) );
  INV_X1 U14945 ( .A(n18518), .ZN(n8617) );
  AOI22_X1 U14946 ( .A1(\mem[1022][7] ), .A2(n18511), .B1(n26108), .B2(
        data_in[7]), .ZN(n18518) );
  INV_X1 U14947 ( .A(n18519), .ZN(n8616) );
  AOI22_X1 U14948 ( .A1(\mem[1023][0] ), .A2(n18520), .B1(n26107), .B2(
        data_in[0]), .ZN(n18519) );
  INV_X1 U14949 ( .A(n18521), .ZN(n8615) );
  AOI22_X1 U14950 ( .A1(\mem[1023][1] ), .A2(n18520), .B1(n26107), .B2(
        data_in[1]), .ZN(n18521) );
  INV_X1 U14951 ( .A(n18522), .ZN(n8614) );
  AOI22_X1 U14952 ( .A1(\mem[1023][2] ), .A2(n18520), .B1(n26107), .B2(
        data_in[2]), .ZN(n18522) );
  INV_X1 U14953 ( .A(n18523), .ZN(n8613) );
  AOI22_X1 U14954 ( .A1(\mem[1023][3] ), .A2(n18520), .B1(n26107), .B2(
        data_in[3]), .ZN(n18523) );
  INV_X1 U14955 ( .A(n18524), .ZN(n8612) );
  AOI22_X1 U14956 ( .A1(\mem[1023][4] ), .A2(n18520), .B1(n26107), .B2(
        data_in[4]), .ZN(n18524) );
  INV_X1 U14957 ( .A(n18525), .ZN(n8611) );
  AOI22_X1 U14958 ( .A1(\mem[1023][5] ), .A2(n18520), .B1(n26107), .B2(
        data_in[5]), .ZN(n18525) );
  INV_X1 U14959 ( .A(n18526), .ZN(n8610) );
  AOI22_X1 U14960 ( .A1(\mem[1023][6] ), .A2(n18520), .B1(n26107), .B2(
        data_in[6]), .ZN(n18526) );
  INV_X1 U14961 ( .A(n18527), .ZN(n8609) );
  AOI22_X1 U14962 ( .A1(\mem[1023][7] ), .A2(n18520), .B1(n26107), .B2(
        data_in[7]), .ZN(n18527) );
  INV_X1 U14963 ( .A(n9547), .ZN(n25850) );
  AOI22_X1 U14964 ( .A1(\mem[32][0] ), .A2(n9548), .B1(n27098), .B2(data_in[0]), .ZN(n9547) );
  INV_X1 U14965 ( .A(n9549), .ZN(n25849) );
  AOI22_X1 U14966 ( .A1(\mem[32][1] ), .A2(n9548), .B1(n27098), .B2(data_in[1]), .ZN(n9549) );
  INV_X1 U14967 ( .A(n9550), .ZN(n25848) );
  AOI22_X1 U14968 ( .A1(\mem[32][2] ), .A2(n9548), .B1(n27098), .B2(data_in[2]), .ZN(n9550) );
  INV_X1 U14969 ( .A(n9551), .ZN(n25847) );
  AOI22_X1 U14970 ( .A1(\mem[32][3] ), .A2(n9548), .B1(n27098), .B2(data_in[3]), .ZN(n9551) );
  INV_X1 U14971 ( .A(n9552), .ZN(n25846) );
  AOI22_X1 U14972 ( .A1(\mem[32][4] ), .A2(n9548), .B1(n27098), .B2(data_in[4]), .ZN(n9552) );
  INV_X1 U14973 ( .A(n9553), .ZN(n25845) );
  AOI22_X1 U14974 ( .A1(\mem[32][5] ), .A2(n9548), .B1(n27098), .B2(data_in[5]), .ZN(n9553) );
  INV_X1 U14975 ( .A(n9554), .ZN(n25844) );
  AOI22_X1 U14976 ( .A1(\mem[32][6] ), .A2(n9548), .B1(n27098), .B2(data_in[6]), .ZN(n9554) );
  INV_X1 U14977 ( .A(n9555), .ZN(n25843) );
  AOI22_X1 U14978 ( .A1(\mem[32][7] ), .A2(n9548), .B1(n27098), .B2(data_in[7]), .ZN(n9555) );
  INV_X1 U14979 ( .A(n9557), .ZN(n25842) );
  AOI22_X1 U14980 ( .A1(\mem[33][0] ), .A2(n9558), .B1(n27097), .B2(data_in[0]), .ZN(n9557) );
  INV_X1 U14981 ( .A(n9559), .ZN(n25841) );
  AOI22_X1 U14982 ( .A1(\mem[33][1] ), .A2(n9558), .B1(n27097), .B2(data_in[1]), .ZN(n9559) );
  INV_X1 U14983 ( .A(n9560), .ZN(n25840) );
  AOI22_X1 U14984 ( .A1(\mem[33][2] ), .A2(n9558), .B1(n27097), .B2(data_in[2]), .ZN(n9560) );
  INV_X1 U14985 ( .A(n9561), .ZN(n25839) );
  AOI22_X1 U14986 ( .A1(\mem[33][3] ), .A2(n9558), .B1(n27097), .B2(data_in[3]), .ZN(n9561) );
  INV_X1 U14987 ( .A(n9562), .ZN(n25838) );
  AOI22_X1 U14988 ( .A1(\mem[33][4] ), .A2(n9558), .B1(n27097), .B2(data_in[4]), .ZN(n9562) );
  INV_X1 U14989 ( .A(n9563), .ZN(n25837) );
  AOI22_X1 U14990 ( .A1(\mem[33][5] ), .A2(n9558), .B1(n27097), .B2(data_in[5]), .ZN(n9563) );
  INV_X1 U14991 ( .A(n9564), .ZN(n25836) );
  AOI22_X1 U14992 ( .A1(\mem[33][6] ), .A2(n9558), .B1(n27097), .B2(data_in[6]), .ZN(n9564) );
  INV_X1 U14993 ( .A(n9565), .ZN(n25835) );
  AOI22_X1 U14994 ( .A1(\mem[33][7] ), .A2(n9558), .B1(n27097), .B2(data_in[7]), .ZN(n9565) );
  INV_X1 U14995 ( .A(n9566), .ZN(n25834) );
  AOI22_X1 U14996 ( .A1(\mem[34][0] ), .A2(n9567), .B1(n27096), .B2(data_in[0]), .ZN(n9566) );
  INV_X1 U14997 ( .A(n9568), .ZN(n25833) );
  AOI22_X1 U14998 ( .A1(\mem[34][1] ), .A2(n9567), .B1(n27096), .B2(data_in[1]), .ZN(n9568) );
  INV_X1 U14999 ( .A(n9569), .ZN(n25832) );
  AOI22_X1 U15000 ( .A1(\mem[34][2] ), .A2(n9567), .B1(n27096), .B2(data_in[2]), .ZN(n9569) );
  INV_X1 U15001 ( .A(n9570), .ZN(n25831) );
  AOI22_X1 U15002 ( .A1(\mem[34][3] ), .A2(n9567), .B1(n27096), .B2(data_in[3]), .ZN(n9570) );
  INV_X1 U15003 ( .A(n9571), .ZN(n25830) );
  AOI22_X1 U15004 ( .A1(\mem[34][4] ), .A2(n9567), .B1(n27096), .B2(data_in[4]), .ZN(n9571) );
  INV_X1 U15005 ( .A(n9572), .ZN(n25829) );
  AOI22_X1 U15006 ( .A1(\mem[34][5] ), .A2(n9567), .B1(n27096), .B2(data_in[5]), .ZN(n9572) );
  INV_X1 U15007 ( .A(n9573), .ZN(n25828) );
  AOI22_X1 U15008 ( .A1(\mem[34][6] ), .A2(n9567), .B1(n27096), .B2(data_in[6]), .ZN(n9573) );
  INV_X1 U15009 ( .A(n9574), .ZN(n25827) );
  AOI22_X1 U15010 ( .A1(\mem[34][7] ), .A2(n9567), .B1(n27096), .B2(data_in[7]), .ZN(n9574) );
  INV_X1 U15011 ( .A(n9575), .ZN(n25826) );
  AOI22_X1 U15012 ( .A1(\mem[35][0] ), .A2(n9576), .B1(n27095), .B2(data_in[0]), .ZN(n9575) );
  INV_X1 U15013 ( .A(n9577), .ZN(n25825) );
  AOI22_X1 U15014 ( .A1(\mem[35][1] ), .A2(n9576), .B1(n27095), .B2(data_in[1]), .ZN(n9577) );
  INV_X1 U15015 ( .A(n9578), .ZN(n25824) );
  AOI22_X1 U15016 ( .A1(\mem[35][2] ), .A2(n9576), .B1(n27095), .B2(data_in[2]), .ZN(n9578) );
  INV_X1 U15017 ( .A(n9579), .ZN(n25823) );
  AOI22_X1 U15018 ( .A1(\mem[35][3] ), .A2(n9576), .B1(n27095), .B2(data_in[3]), .ZN(n9579) );
  INV_X1 U15019 ( .A(n9580), .ZN(n25822) );
  AOI22_X1 U15020 ( .A1(\mem[35][4] ), .A2(n9576), .B1(n27095), .B2(data_in[4]), .ZN(n9580) );
  INV_X1 U15021 ( .A(n9581), .ZN(n25821) );
  AOI22_X1 U15022 ( .A1(\mem[35][5] ), .A2(n9576), .B1(n27095), .B2(data_in[5]), .ZN(n9581) );
  INV_X1 U15023 ( .A(n9582), .ZN(n25820) );
  AOI22_X1 U15024 ( .A1(\mem[35][6] ), .A2(n9576), .B1(n27095), .B2(data_in[6]), .ZN(n9582) );
  INV_X1 U15025 ( .A(n9583), .ZN(n25819) );
  AOI22_X1 U15026 ( .A1(\mem[35][7] ), .A2(n9576), .B1(n27095), .B2(data_in[7]), .ZN(n9583) );
  INV_X1 U15027 ( .A(n9584), .ZN(n25818) );
  AOI22_X1 U15028 ( .A1(\mem[36][0] ), .A2(n9585), .B1(n27094), .B2(data_in[0]), .ZN(n9584) );
  INV_X1 U15029 ( .A(n9586), .ZN(n25817) );
  AOI22_X1 U15030 ( .A1(\mem[36][1] ), .A2(n9585), .B1(n27094), .B2(data_in[1]), .ZN(n9586) );
  INV_X1 U15031 ( .A(n9587), .ZN(n25816) );
  AOI22_X1 U15032 ( .A1(\mem[36][2] ), .A2(n9585), .B1(n27094), .B2(data_in[2]), .ZN(n9587) );
  INV_X1 U15033 ( .A(n9588), .ZN(n25815) );
  AOI22_X1 U15034 ( .A1(\mem[36][3] ), .A2(n9585), .B1(n27094), .B2(data_in[3]), .ZN(n9588) );
  INV_X1 U15035 ( .A(n9589), .ZN(n25814) );
  AOI22_X1 U15036 ( .A1(\mem[36][4] ), .A2(n9585), .B1(n27094), .B2(data_in[4]), .ZN(n9589) );
  INV_X1 U15037 ( .A(n9590), .ZN(n25813) );
  AOI22_X1 U15038 ( .A1(\mem[36][5] ), .A2(n9585), .B1(n27094), .B2(data_in[5]), .ZN(n9590) );
  INV_X1 U15039 ( .A(n9591), .ZN(n25812) );
  AOI22_X1 U15040 ( .A1(\mem[36][6] ), .A2(n9585), .B1(n27094), .B2(data_in[6]), .ZN(n9591) );
  INV_X1 U15041 ( .A(n9592), .ZN(n25811) );
  AOI22_X1 U15042 ( .A1(\mem[36][7] ), .A2(n9585), .B1(n27094), .B2(data_in[7]), .ZN(n9592) );
  INV_X1 U15043 ( .A(n9593), .ZN(n25810) );
  AOI22_X1 U15044 ( .A1(\mem[37][0] ), .A2(n9594), .B1(n27093), .B2(data_in[0]), .ZN(n9593) );
  INV_X1 U15045 ( .A(n9595), .ZN(n25809) );
  AOI22_X1 U15046 ( .A1(\mem[37][1] ), .A2(n9594), .B1(n27093), .B2(data_in[1]), .ZN(n9595) );
  INV_X1 U15047 ( .A(n9596), .ZN(n25808) );
  AOI22_X1 U15048 ( .A1(\mem[37][2] ), .A2(n9594), .B1(n27093), .B2(data_in[2]), .ZN(n9596) );
  INV_X1 U15049 ( .A(n9597), .ZN(n25807) );
  AOI22_X1 U15050 ( .A1(\mem[37][3] ), .A2(n9594), .B1(n27093), .B2(data_in[3]), .ZN(n9597) );
  INV_X1 U15051 ( .A(n9598), .ZN(n25806) );
  AOI22_X1 U15052 ( .A1(\mem[37][4] ), .A2(n9594), .B1(n27093), .B2(data_in[4]), .ZN(n9598) );
  INV_X1 U15053 ( .A(n9599), .ZN(n25805) );
  AOI22_X1 U15054 ( .A1(\mem[37][5] ), .A2(n9594), .B1(n27093), .B2(data_in[5]), .ZN(n9599) );
  INV_X1 U15055 ( .A(n9600), .ZN(n25804) );
  AOI22_X1 U15056 ( .A1(\mem[37][6] ), .A2(n9594), .B1(n27093), .B2(data_in[6]), .ZN(n9600) );
  INV_X1 U15057 ( .A(n9601), .ZN(n25803) );
  AOI22_X1 U15058 ( .A1(\mem[37][7] ), .A2(n9594), .B1(n27093), .B2(data_in[7]), .ZN(n9601) );
  INV_X1 U15059 ( .A(n9602), .ZN(n25802) );
  AOI22_X1 U15060 ( .A1(\mem[38][0] ), .A2(n9603), .B1(n27092), .B2(data_in[0]), .ZN(n9602) );
  INV_X1 U15061 ( .A(n9604), .ZN(n25801) );
  AOI22_X1 U15062 ( .A1(\mem[38][1] ), .A2(n9603), .B1(n27092), .B2(data_in[1]), .ZN(n9604) );
  INV_X1 U15063 ( .A(n9605), .ZN(n25800) );
  AOI22_X1 U15064 ( .A1(\mem[38][2] ), .A2(n9603), .B1(n27092), .B2(data_in[2]), .ZN(n9605) );
  INV_X1 U15065 ( .A(n9606), .ZN(n25799) );
  AOI22_X1 U15066 ( .A1(\mem[38][3] ), .A2(n9603), .B1(n27092), .B2(data_in[3]), .ZN(n9606) );
  INV_X1 U15067 ( .A(n9607), .ZN(n25798) );
  AOI22_X1 U15068 ( .A1(\mem[38][4] ), .A2(n9603), .B1(n27092), .B2(data_in[4]), .ZN(n9607) );
  INV_X1 U15069 ( .A(n9608), .ZN(n25797) );
  AOI22_X1 U15070 ( .A1(\mem[38][5] ), .A2(n9603), .B1(n27092), .B2(data_in[5]), .ZN(n9608) );
  INV_X1 U15071 ( .A(n9609), .ZN(n25796) );
  AOI22_X1 U15072 ( .A1(\mem[38][6] ), .A2(n9603), .B1(n27092), .B2(data_in[6]), .ZN(n9609) );
  INV_X1 U15073 ( .A(n9610), .ZN(n25795) );
  AOI22_X1 U15074 ( .A1(\mem[38][7] ), .A2(n9603), .B1(n27092), .B2(data_in[7]), .ZN(n9610) );
  INV_X1 U15075 ( .A(n9611), .ZN(n25794) );
  AOI22_X1 U15076 ( .A1(\mem[39][0] ), .A2(n9612), .B1(n27091), .B2(data_in[0]), .ZN(n9611) );
  INV_X1 U15077 ( .A(n9613), .ZN(n25793) );
  AOI22_X1 U15078 ( .A1(\mem[39][1] ), .A2(n9612), .B1(n27091), .B2(data_in[1]), .ZN(n9613) );
  INV_X1 U15079 ( .A(n9614), .ZN(n25792) );
  AOI22_X1 U15080 ( .A1(\mem[39][2] ), .A2(n9612), .B1(n27091), .B2(data_in[2]), .ZN(n9614) );
  INV_X1 U15081 ( .A(n9615), .ZN(n25791) );
  AOI22_X1 U15082 ( .A1(\mem[39][3] ), .A2(n9612), .B1(n27091), .B2(data_in[3]), .ZN(n9615) );
  INV_X1 U15083 ( .A(n9616), .ZN(n25790) );
  AOI22_X1 U15084 ( .A1(\mem[39][4] ), .A2(n9612), .B1(n27091), .B2(data_in[4]), .ZN(n9616) );
  INV_X1 U15085 ( .A(n9617), .ZN(n25789) );
  AOI22_X1 U15086 ( .A1(\mem[39][5] ), .A2(n9612), .B1(n27091), .B2(data_in[5]), .ZN(n9617) );
  INV_X1 U15087 ( .A(n9618), .ZN(n25788) );
  AOI22_X1 U15088 ( .A1(\mem[39][6] ), .A2(n9612), .B1(n27091), .B2(data_in[6]), .ZN(n9618) );
  INV_X1 U15089 ( .A(n9619), .ZN(n25787) );
  AOI22_X1 U15090 ( .A1(\mem[39][7] ), .A2(n9612), .B1(n27091), .B2(data_in[7]), .ZN(n9619) );
  INV_X1 U15091 ( .A(n9837), .ZN(n25594) );
  AOI22_X1 U15092 ( .A1(\mem[64][0] ), .A2(n9838), .B1(n27066), .B2(data_in[0]), .ZN(n9837) );
  INV_X1 U15093 ( .A(n9839), .ZN(n25593) );
  AOI22_X1 U15094 ( .A1(\mem[64][1] ), .A2(n9838), .B1(n27066), .B2(data_in[1]), .ZN(n9839) );
  INV_X1 U15095 ( .A(n9840), .ZN(n25592) );
  AOI22_X1 U15096 ( .A1(\mem[64][2] ), .A2(n9838), .B1(n27066), .B2(data_in[2]), .ZN(n9840) );
  INV_X1 U15097 ( .A(n9841), .ZN(n25591) );
  AOI22_X1 U15098 ( .A1(\mem[64][3] ), .A2(n9838), .B1(n27066), .B2(data_in[3]), .ZN(n9841) );
  INV_X1 U15099 ( .A(n9842), .ZN(n25590) );
  AOI22_X1 U15100 ( .A1(\mem[64][4] ), .A2(n9838), .B1(n27066), .B2(data_in[4]), .ZN(n9842) );
  INV_X1 U15101 ( .A(n9843), .ZN(n25589) );
  AOI22_X1 U15102 ( .A1(\mem[64][5] ), .A2(n9838), .B1(n27066), .B2(data_in[5]), .ZN(n9843) );
  INV_X1 U15103 ( .A(n9844), .ZN(n25588) );
  AOI22_X1 U15104 ( .A1(\mem[64][6] ), .A2(n9838), .B1(n27066), .B2(data_in[6]), .ZN(n9844) );
  INV_X1 U15105 ( .A(n9845), .ZN(n25587) );
  AOI22_X1 U15106 ( .A1(\mem[64][7] ), .A2(n9838), .B1(n27066), .B2(data_in[7]), .ZN(n9845) );
  INV_X1 U15107 ( .A(n9847), .ZN(n25586) );
  AOI22_X1 U15108 ( .A1(\mem[65][0] ), .A2(n9848), .B1(n27065), .B2(data_in[0]), .ZN(n9847) );
  INV_X1 U15109 ( .A(n9849), .ZN(n25585) );
  AOI22_X1 U15110 ( .A1(\mem[65][1] ), .A2(n9848), .B1(n27065), .B2(data_in[1]), .ZN(n9849) );
  INV_X1 U15111 ( .A(n9850), .ZN(n25584) );
  AOI22_X1 U15112 ( .A1(\mem[65][2] ), .A2(n9848), .B1(n27065), .B2(data_in[2]), .ZN(n9850) );
  INV_X1 U15113 ( .A(n9851), .ZN(n25583) );
  AOI22_X1 U15114 ( .A1(\mem[65][3] ), .A2(n9848), .B1(n27065), .B2(data_in[3]), .ZN(n9851) );
  INV_X1 U15115 ( .A(n9852), .ZN(n25582) );
  AOI22_X1 U15116 ( .A1(\mem[65][4] ), .A2(n9848), .B1(n27065), .B2(data_in[4]), .ZN(n9852) );
  INV_X1 U15117 ( .A(n9853), .ZN(n25581) );
  AOI22_X1 U15118 ( .A1(\mem[65][5] ), .A2(n9848), .B1(n27065), .B2(data_in[5]), .ZN(n9853) );
  INV_X1 U15119 ( .A(n9854), .ZN(n25580) );
  AOI22_X1 U15120 ( .A1(\mem[65][6] ), .A2(n9848), .B1(n27065), .B2(data_in[6]), .ZN(n9854) );
  INV_X1 U15121 ( .A(n9855), .ZN(n25579) );
  AOI22_X1 U15122 ( .A1(\mem[65][7] ), .A2(n9848), .B1(n27065), .B2(data_in[7]), .ZN(n9855) );
  INV_X1 U15123 ( .A(n9856), .ZN(n25578) );
  AOI22_X1 U15124 ( .A1(\mem[66][0] ), .A2(n9857), .B1(n27064), .B2(data_in[0]), .ZN(n9856) );
  INV_X1 U15125 ( .A(n9858), .ZN(n25577) );
  AOI22_X1 U15126 ( .A1(\mem[66][1] ), .A2(n9857), .B1(n27064), .B2(data_in[1]), .ZN(n9858) );
  INV_X1 U15127 ( .A(n9859), .ZN(n25576) );
  AOI22_X1 U15128 ( .A1(\mem[66][2] ), .A2(n9857), .B1(n27064), .B2(data_in[2]), .ZN(n9859) );
  INV_X1 U15129 ( .A(n9860), .ZN(n25575) );
  AOI22_X1 U15130 ( .A1(\mem[66][3] ), .A2(n9857), .B1(n27064), .B2(data_in[3]), .ZN(n9860) );
  INV_X1 U15131 ( .A(n9861), .ZN(n25574) );
  AOI22_X1 U15132 ( .A1(\mem[66][4] ), .A2(n9857), .B1(n27064), .B2(data_in[4]), .ZN(n9861) );
  INV_X1 U15133 ( .A(n9862), .ZN(n25573) );
  AOI22_X1 U15134 ( .A1(\mem[66][5] ), .A2(n9857), .B1(n27064), .B2(data_in[5]), .ZN(n9862) );
  INV_X1 U15135 ( .A(n9863), .ZN(n25572) );
  AOI22_X1 U15136 ( .A1(\mem[66][6] ), .A2(n9857), .B1(n27064), .B2(data_in[6]), .ZN(n9863) );
  INV_X1 U15137 ( .A(n9864), .ZN(n25571) );
  AOI22_X1 U15138 ( .A1(\mem[66][7] ), .A2(n9857), .B1(n27064), .B2(data_in[7]), .ZN(n9864) );
  INV_X1 U15139 ( .A(n9865), .ZN(n25570) );
  AOI22_X1 U15140 ( .A1(\mem[67][0] ), .A2(n9866), .B1(n27063), .B2(data_in[0]), .ZN(n9865) );
  INV_X1 U15141 ( .A(n9867), .ZN(n25569) );
  AOI22_X1 U15142 ( .A1(\mem[67][1] ), .A2(n9866), .B1(n27063), .B2(data_in[1]), .ZN(n9867) );
  INV_X1 U15143 ( .A(n9868), .ZN(n25568) );
  AOI22_X1 U15144 ( .A1(\mem[67][2] ), .A2(n9866), .B1(n27063), .B2(data_in[2]), .ZN(n9868) );
  INV_X1 U15145 ( .A(n9869), .ZN(n25567) );
  AOI22_X1 U15146 ( .A1(\mem[67][3] ), .A2(n9866), .B1(n27063), .B2(data_in[3]), .ZN(n9869) );
  INV_X1 U15147 ( .A(n9870), .ZN(n25566) );
  AOI22_X1 U15148 ( .A1(\mem[67][4] ), .A2(n9866), .B1(n27063), .B2(data_in[4]), .ZN(n9870) );
  INV_X1 U15149 ( .A(n9871), .ZN(n25565) );
  AOI22_X1 U15150 ( .A1(\mem[67][5] ), .A2(n9866), .B1(n27063), .B2(data_in[5]), .ZN(n9871) );
  INV_X1 U15151 ( .A(n9872), .ZN(n25564) );
  AOI22_X1 U15152 ( .A1(\mem[67][6] ), .A2(n9866), .B1(n27063), .B2(data_in[6]), .ZN(n9872) );
  INV_X1 U15153 ( .A(n9873), .ZN(n25563) );
  AOI22_X1 U15154 ( .A1(\mem[67][7] ), .A2(n9866), .B1(n27063), .B2(data_in[7]), .ZN(n9873) );
  INV_X1 U15155 ( .A(n9874), .ZN(n25562) );
  AOI22_X1 U15156 ( .A1(\mem[68][0] ), .A2(n9875), .B1(n27062), .B2(data_in[0]), .ZN(n9874) );
  INV_X1 U15157 ( .A(n9876), .ZN(n25561) );
  AOI22_X1 U15158 ( .A1(\mem[68][1] ), .A2(n9875), .B1(n27062), .B2(data_in[1]), .ZN(n9876) );
  INV_X1 U15159 ( .A(n9877), .ZN(n25560) );
  AOI22_X1 U15160 ( .A1(\mem[68][2] ), .A2(n9875), .B1(n27062), .B2(data_in[2]), .ZN(n9877) );
  INV_X1 U15161 ( .A(n9878), .ZN(n25559) );
  AOI22_X1 U15162 ( .A1(\mem[68][3] ), .A2(n9875), .B1(n27062), .B2(data_in[3]), .ZN(n9878) );
  INV_X1 U15163 ( .A(n9879), .ZN(n25558) );
  AOI22_X1 U15164 ( .A1(\mem[68][4] ), .A2(n9875), .B1(n27062), .B2(data_in[4]), .ZN(n9879) );
  INV_X1 U15165 ( .A(n9880), .ZN(n25557) );
  AOI22_X1 U15166 ( .A1(\mem[68][5] ), .A2(n9875), .B1(n27062), .B2(data_in[5]), .ZN(n9880) );
  INV_X1 U15167 ( .A(n9881), .ZN(n25556) );
  AOI22_X1 U15168 ( .A1(\mem[68][6] ), .A2(n9875), .B1(n27062), .B2(data_in[6]), .ZN(n9881) );
  INV_X1 U15169 ( .A(n9882), .ZN(n25555) );
  AOI22_X1 U15170 ( .A1(\mem[68][7] ), .A2(n9875), .B1(n27062), .B2(data_in[7]), .ZN(n9882) );
  INV_X1 U15171 ( .A(n9883), .ZN(n25554) );
  AOI22_X1 U15172 ( .A1(\mem[69][0] ), .A2(n9884), .B1(n27061), .B2(data_in[0]), .ZN(n9883) );
  INV_X1 U15173 ( .A(n9885), .ZN(n25553) );
  AOI22_X1 U15174 ( .A1(\mem[69][1] ), .A2(n9884), .B1(n27061), .B2(data_in[1]), .ZN(n9885) );
  INV_X1 U15175 ( .A(n9886), .ZN(n25552) );
  AOI22_X1 U15176 ( .A1(\mem[69][2] ), .A2(n9884), .B1(n27061), .B2(data_in[2]), .ZN(n9886) );
  INV_X1 U15177 ( .A(n9887), .ZN(n25551) );
  AOI22_X1 U15178 ( .A1(\mem[69][3] ), .A2(n9884), .B1(n27061), .B2(data_in[3]), .ZN(n9887) );
  INV_X1 U15179 ( .A(n9888), .ZN(n25550) );
  AOI22_X1 U15180 ( .A1(\mem[69][4] ), .A2(n9884), .B1(n27061), .B2(data_in[4]), .ZN(n9888) );
  INV_X1 U15181 ( .A(n9889), .ZN(n25549) );
  AOI22_X1 U15182 ( .A1(\mem[69][5] ), .A2(n9884), .B1(n27061), .B2(data_in[5]), .ZN(n9889) );
  INV_X1 U15183 ( .A(n9890), .ZN(n25548) );
  AOI22_X1 U15184 ( .A1(\mem[69][6] ), .A2(n9884), .B1(n27061), .B2(data_in[6]), .ZN(n9890) );
  INV_X1 U15185 ( .A(n9891), .ZN(n25547) );
  AOI22_X1 U15186 ( .A1(\mem[69][7] ), .A2(n9884), .B1(n27061), .B2(data_in[7]), .ZN(n9891) );
  INV_X1 U15187 ( .A(n9892), .ZN(n25546) );
  AOI22_X1 U15188 ( .A1(\mem[70][0] ), .A2(n9893), .B1(n27060), .B2(data_in[0]), .ZN(n9892) );
  INV_X1 U15189 ( .A(n9894), .ZN(n25545) );
  AOI22_X1 U15190 ( .A1(\mem[70][1] ), .A2(n9893), .B1(n27060), .B2(data_in[1]), .ZN(n9894) );
  INV_X1 U15191 ( .A(n9895), .ZN(n25544) );
  AOI22_X1 U15192 ( .A1(\mem[70][2] ), .A2(n9893), .B1(n27060), .B2(data_in[2]), .ZN(n9895) );
  INV_X1 U15193 ( .A(n9896), .ZN(n25543) );
  AOI22_X1 U15194 ( .A1(\mem[70][3] ), .A2(n9893), .B1(n27060), .B2(data_in[3]), .ZN(n9896) );
  INV_X1 U15195 ( .A(n9897), .ZN(n25542) );
  AOI22_X1 U15196 ( .A1(\mem[70][4] ), .A2(n9893), .B1(n27060), .B2(data_in[4]), .ZN(n9897) );
  INV_X1 U15197 ( .A(n9898), .ZN(n25541) );
  AOI22_X1 U15198 ( .A1(\mem[70][5] ), .A2(n9893), .B1(n27060), .B2(data_in[5]), .ZN(n9898) );
  INV_X1 U15199 ( .A(n9899), .ZN(n25540) );
  AOI22_X1 U15200 ( .A1(\mem[70][6] ), .A2(n9893), .B1(n27060), .B2(data_in[6]), .ZN(n9899) );
  INV_X1 U15201 ( .A(n9900), .ZN(n25539) );
  AOI22_X1 U15202 ( .A1(\mem[70][7] ), .A2(n9893), .B1(n27060), .B2(data_in[7]), .ZN(n9900) );
  INV_X1 U15203 ( .A(n9901), .ZN(n25538) );
  AOI22_X1 U15204 ( .A1(\mem[71][0] ), .A2(n9902), .B1(n27059), .B2(data_in[0]), .ZN(n9901) );
  INV_X1 U15205 ( .A(n9903), .ZN(n25537) );
  AOI22_X1 U15206 ( .A1(\mem[71][1] ), .A2(n9902), .B1(n27059), .B2(data_in[1]), .ZN(n9903) );
  INV_X1 U15207 ( .A(n9904), .ZN(n25536) );
  AOI22_X1 U15208 ( .A1(\mem[71][2] ), .A2(n9902), .B1(n27059), .B2(data_in[2]), .ZN(n9904) );
  INV_X1 U15209 ( .A(n9905), .ZN(n25535) );
  AOI22_X1 U15210 ( .A1(\mem[71][3] ), .A2(n9902), .B1(n27059), .B2(data_in[3]), .ZN(n9905) );
  INV_X1 U15211 ( .A(n9906), .ZN(n25534) );
  AOI22_X1 U15212 ( .A1(\mem[71][4] ), .A2(n9902), .B1(n27059), .B2(data_in[4]), .ZN(n9906) );
  INV_X1 U15213 ( .A(n9907), .ZN(n25533) );
  AOI22_X1 U15214 ( .A1(\mem[71][5] ), .A2(n9902), .B1(n27059), .B2(data_in[5]), .ZN(n9907) );
  INV_X1 U15215 ( .A(n9908), .ZN(n25532) );
  AOI22_X1 U15216 ( .A1(\mem[71][6] ), .A2(n9902), .B1(n27059), .B2(data_in[6]), .ZN(n9908) );
  INV_X1 U15217 ( .A(n9909), .ZN(n25531) );
  AOI22_X1 U15218 ( .A1(\mem[71][7] ), .A2(n9902), .B1(n27059), .B2(data_in[7]), .ZN(n9909) );
  INV_X1 U15219 ( .A(n10127), .ZN(n25338) );
  AOI22_X1 U15220 ( .A1(\mem[96][0] ), .A2(n10128), .B1(n27034), .B2(
        data_in[0]), .ZN(n10127) );
  INV_X1 U15221 ( .A(n10129), .ZN(n25337) );
  AOI22_X1 U15222 ( .A1(\mem[96][1] ), .A2(n10128), .B1(n27034), .B2(
        data_in[1]), .ZN(n10129) );
  INV_X1 U15223 ( .A(n10130), .ZN(n25336) );
  AOI22_X1 U15224 ( .A1(\mem[96][2] ), .A2(n10128), .B1(n27034), .B2(
        data_in[2]), .ZN(n10130) );
  INV_X1 U15225 ( .A(n10131), .ZN(n25335) );
  AOI22_X1 U15226 ( .A1(\mem[96][3] ), .A2(n10128), .B1(n27034), .B2(
        data_in[3]), .ZN(n10131) );
  INV_X1 U15227 ( .A(n10132), .ZN(n25334) );
  AOI22_X1 U15228 ( .A1(\mem[96][4] ), .A2(n10128), .B1(n27034), .B2(
        data_in[4]), .ZN(n10132) );
  INV_X1 U15229 ( .A(n10133), .ZN(n25333) );
  AOI22_X1 U15230 ( .A1(\mem[96][5] ), .A2(n10128), .B1(n27034), .B2(
        data_in[5]), .ZN(n10133) );
  INV_X1 U15231 ( .A(n10134), .ZN(n25332) );
  AOI22_X1 U15232 ( .A1(\mem[96][6] ), .A2(n10128), .B1(n27034), .B2(
        data_in[6]), .ZN(n10134) );
  INV_X1 U15233 ( .A(n10135), .ZN(n25331) );
  AOI22_X1 U15234 ( .A1(\mem[96][7] ), .A2(n10128), .B1(n27034), .B2(
        data_in[7]), .ZN(n10135) );
  INV_X1 U15235 ( .A(n10137), .ZN(n25330) );
  AOI22_X1 U15236 ( .A1(\mem[97][0] ), .A2(n10138), .B1(n27033), .B2(
        data_in[0]), .ZN(n10137) );
  INV_X1 U15237 ( .A(n10139), .ZN(n25329) );
  AOI22_X1 U15238 ( .A1(\mem[97][1] ), .A2(n10138), .B1(n27033), .B2(
        data_in[1]), .ZN(n10139) );
  INV_X1 U15239 ( .A(n10140), .ZN(n25328) );
  AOI22_X1 U15240 ( .A1(\mem[97][2] ), .A2(n10138), .B1(n27033), .B2(
        data_in[2]), .ZN(n10140) );
  INV_X1 U15241 ( .A(n10141), .ZN(n25327) );
  AOI22_X1 U15242 ( .A1(\mem[97][3] ), .A2(n10138), .B1(n27033), .B2(
        data_in[3]), .ZN(n10141) );
  INV_X1 U15243 ( .A(n10142), .ZN(n25326) );
  AOI22_X1 U15244 ( .A1(\mem[97][4] ), .A2(n10138), .B1(n27033), .B2(
        data_in[4]), .ZN(n10142) );
  INV_X1 U15245 ( .A(n10143), .ZN(n25325) );
  AOI22_X1 U15246 ( .A1(\mem[97][5] ), .A2(n10138), .B1(n27033), .B2(
        data_in[5]), .ZN(n10143) );
  INV_X1 U15247 ( .A(n10144), .ZN(n25324) );
  AOI22_X1 U15248 ( .A1(\mem[97][6] ), .A2(n10138), .B1(n27033), .B2(
        data_in[6]), .ZN(n10144) );
  INV_X1 U15249 ( .A(n10145), .ZN(n25323) );
  AOI22_X1 U15250 ( .A1(\mem[97][7] ), .A2(n10138), .B1(n27033), .B2(
        data_in[7]), .ZN(n10145) );
  INV_X1 U15251 ( .A(n10146), .ZN(n25322) );
  AOI22_X1 U15252 ( .A1(\mem[98][0] ), .A2(n10147), .B1(n27032), .B2(
        data_in[0]), .ZN(n10146) );
  INV_X1 U15253 ( .A(n10148), .ZN(n25321) );
  AOI22_X1 U15254 ( .A1(\mem[98][1] ), .A2(n10147), .B1(n27032), .B2(
        data_in[1]), .ZN(n10148) );
  INV_X1 U15255 ( .A(n10149), .ZN(n25320) );
  AOI22_X1 U15256 ( .A1(\mem[98][2] ), .A2(n10147), .B1(n27032), .B2(
        data_in[2]), .ZN(n10149) );
  INV_X1 U15257 ( .A(n10150), .ZN(n25319) );
  AOI22_X1 U15258 ( .A1(\mem[98][3] ), .A2(n10147), .B1(n27032), .B2(
        data_in[3]), .ZN(n10150) );
  INV_X1 U15259 ( .A(n10151), .ZN(n25318) );
  AOI22_X1 U15260 ( .A1(\mem[98][4] ), .A2(n10147), .B1(n27032), .B2(
        data_in[4]), .ZN(n10151) );
  INV_X1 U15261 ( .A(n10152), .ZN(n25317) );
  AOI22_X1 U15262 ( .A1(\mem[98][5] ), .A2(n10147), .B1(n27032), .B2(
        data_in[5]), .ZN(n10152) );
  INV_X1 U15263 ( .A(n10153), .ZN(n25316) );
  AOI22_X1 U15264 ( .A1(\mem[98][6] ), .A2(n10147), .B1(n27032), .B2(
        data_in[6]), .ZN(n10153) );
  INV_X1 U15265 ( .A(n10154), .ZN(n25315) );
  AOI22_X1 U15266 ( .A1(\mem[98][7] ), .A2(n10147), .B1(n27032), .B2(
        data_in[7]), .ZN(n10154) );
  INV_X1 U15267 ( .A(n10155), .ZN(n25314) );
  AOI22_X1 U15268 ( .A1(\mem[99][0] ), .A2(n10156), .B1(n27031), .B2(
        data_in[0]), .ZN(n10155) );
  INV_X1 U15269 ( .A(n10157), .ZN(n25313) );
  AOI22_X1 U15270 ( .A1(\mem[99][1] ), .A2(n10156), .B1(n27031), .B2(
        data_in[1]), .ZN(n10157) );
  INV_X1 U15271 ( .A(n10158), .ZN(n25312) );
  AOI22_X1 U15272 ( .A1(\mem[99][2] ), .A2(n10156), .B1(n27031), .B2(
        data_in[2]), .ZN(n10158) );
  INV_X1 U15273 ( .A(n10159), .ZN(n25311) );
  AOI22_X1 U15274 ( .A1(\mem[99][3] ), .A2(n10156), .B1(n27031), .B2(
        data_in[3]), .ZN(n10159) );
  INV_X1 U15275 ( .A(n10160), .ZN(n25310) );
  AOI22_X1 U15276 ( .A1(\mem[99][4] ), .A2(n10156), .B1(n27031), .B2(
        data_in[4]), .ZN(n10160) );
  INV_X1 U15277 ( .A(n10161), .ZN(n25309) );
  AOI22_X1 U15278 ( .A1(\mem[99][5] ), .A2(n10156), .B1(n27031), .B2(
        data_in[5]), .ZN(n10161) );
  INV_X1 U15279 ( .A(n10162), .ZN(n25308) );
  AOI22_X1 U15280 ( .A1(\mem[99][6] ), .A2(n10156), .B1(n27031), .B2(
        data_in[6]), .ZN(n10162) );
  INV_X1 U15281 ( .A(n10163), .ZN(n25307) );
  AOI22_X1 U15282 ( .A1(\mem[99][7] ), .A2(n10156), .B1(n27031), .B2(
        data_in[7]), .ZN(n10163) );
  INV_X1 U15283 ( .A(n10164), .ZN(n25306) );
  AOI22_X1 U15284 ( .A1(\mem[100][0] ), .A2(n10165), .B1(n27030), .B2(
        data_in[0]), .ZN(n10164) );
  INV_X1 U15285 ( .A(n10166), .ZN(n25305) );
  AOI22_X1 U15286 ( .A1(\mem[100][1] ), .A2(n10165), .B1(n27030), .B2(
        data_in[1]), .ZN(n10166) );
  INV_X1 U15287 ( .A(n10167), .ZN(n25304) );
  AOI22_X1 U15288 ( .A1(\mem[100][2] ), .A2(n10165), .B1(n27030), .B2(
        data_in[2]), .ZN(n10167) );
  INV_X1 U15289 ( .A(n10168), .ZN(n25303) );
  AOI22_X1 U15290 ( .A1(\mem[100][3] ), .A2(n10165), .B1(n27030), .B2(
        data_in[3]), .ZN(n10168) );
  INV_X1 U15291 ( .A(n10169), .ZN(n25302) );
  AOI22_X1 U15292 ( .A1(\mem[100][4] ), .A2(n10165), .B1(n27030), .B2(
        data_in[4]), .ZN(n10169) );
  INV_X1 U15293 ( .A(n10170), .ZN(n25301) );
  AOI22_X1 U15294 ( .A1(\mem[100][5] ), .A2(n10165), .B1(n27030), .B2(
        data_in[5]), .ZN(n10170) );
  INV_X1 U15295 ( .A(n10171), .ZN(n25300) );
  AOI22_X1 U15296 ( .A1(\mem[100][6] ), .A2(n10165), .B1(n27030), .B2(
        data_in[6]), .ZN(n10171) );
  INV_X1 U15297 ( .A(n10172), .ZN(n25299) );
  AOI22_X1 U15298 ( .A1(\mem[100][7] ), .A2(n10165), .B1(n27030), .B2(
        data_in[7]), .ZN(n10172) );
  INV_X1 U15299 ( .A(n10173), .ZN(n25298) );
  AOI22_X1 U15300 ( .A1(\mem[101][0] ), .A2(n10174), .B1(n27029), .B2(
        data_in[0]), .ZN(n10173) );
  INV_X1 U15301 ( .A(n10175), .ZN(n25297) );
  AOI22_X1 U15302 ( .A1(\mem[101][1] ), .A2(n10174), .B1(n27029), .B2(
        data_in[1]), .ZN(n10175) );
  INV_X1 U15303 ( .A(n10176), .ZN(n25296) );
  AOI22_X1 U15304 ( .A1(\mem[101][2] ), .A2(n10174), .B1(n27029), .B2(
        data_in[2]), .ZN(n10176) );
  INV_X1 U15305 ( .A(n10177), .ZN(n25295) );
  AOI22_X1 U15306 ( .A1(\mem[101][3] ), .A2(n10174), .B1(n27029), .B2(
        data_in[3]), .ZN(n10177) );
  INV_X1 U15307 ( .A(n10178), .ZN(n25294) );
  AOI22_X1 U15308 ( .A1(\mem[101][4] ), .A2(n10174), .B1(n27029), .B2(
        data_in[4]), .ZN(n10178) );
  INV_X1 U15309 ( .A(n10179), .ZN(n25293) );
  AOI22_X1 U15310 ( .A1(\mem[101][5] ), .A2(n10174), .B1(n27029), .B2(
        data_in[5]), .ZN(n10179) );
  INV_X1 U15311 ( .A(n10180), .ZN(n25292) );
  AOI22_X1 U15312 ( .A1(\mem[101][6] ), .A2(n10174), .B1(n27029), .B2(
        data_in[6]), .ZN(n10180) );
  INV_X1 U15313 ( .A(n10181), .ZN(n25291) );
  AOI22_X1 U15314 ( .A1(\mem[101][7] ), .A2(n10174), .B1(n27029), .B2(
        data_in[7]), .ZN(n10181) );
  INV_X1 U15315 ( .A(n10182), .ZN(n25290) );
  AOI22_X1 U15316 ( .A1(\mem[102][0] ), .A2(n10183), .B1(n27028), .B2(
        data_in[0]), .ZN(n10182) );
  INV_X1 U15317 ( .A(n10184), .ZN(n25289) );
  AOI22_X1 U15318 ( .A1(\mem[102][1] ), .A2(n10183), .B1(n27028), .B2(
        data_in[1]), .ZN(n10184) );
  INV_X1 U15319 ( .A(n10185), .ZN(n25288) );
  AOI22_X1 U15320 ( .A1(\mem[102][2] ), .A2(n10183), .B1(n27028), .B2(
        data_in[2]), .ZN(n10185) );
  INV_X1 U15321 ( .A(n10186), .ZN(n25287) );
  AOI22_X1 U15322 ( .A1(\mem[102][3] ), .A2(n10183), .B1(n27028), .B2(
        data_in[3]), .ZN(n10186) );
  INV_X1 U15323 ( .A(n10187), .ZN(n25286) );
  AOI22_X1 U15324 ( .A1(\mem[102][4] ), .A2(n10183), .B1(n27028), .B2(
        data_in[4]), .ZN(n10187) );
  INV_X1 U15325 ( .A(n10188), .ZN(n25285) );
  AOI22_X1 U15326 ( .A1(\mem[102][5] ), .A2(n10183), .B1(n27028), .B2(
        data_in[5]), .ZN(n10188) );
  INV_X1 U15327 ( .A(n10189), .ZN(n25284) );
  AOI22_X1 U15328 ( .A1(\mem[102][6] ), .A2(n10183), .B1(n27028), .B2(
        data_in[6]), .ZN(n10189) );
  INV_X1 U15329 ( .A(n10190), .ZN(n25283) );
  AOI22_X1 U15330 ( .A1(\mem[102][7] ), .A2(n10183), .B1(n27028), .B2(
        data_in[7]), .ZN(n10190) );
  INV_X1 U15331 ( .A(n10191), .ZN(n25282) );
  AOI22_X1 U15332 ( .A1(\mem[103][0] ), .A2(n10192), .B1(n27027), .B2(
        data_in[0]), .ZN(n10191) );
  INV_X1 U15333 ( .A(n10193), .ZN(n25281) );
  AOI22_X1 U15334 ( .A1(\mem[103][1] ), .A2(n10192), .B1(n27027), .B2(
        data_in[1]), .ZN(n10193) );
  INV_X1 U15335 ( .A(n10194), .ZN(n25280) );
  AOI22_X1 U15336 ( .A1(\mem[103][2] ), .A2(n10192), .B1(n27027), .B2(
        data_in[2]), .ZN(n10194) );
  INV_X1 U15337 ( .A(n10195), .ZN(n25279) );
  AOI22_X1 U15338 ( .A1(\mem[103][3] ), .A2(n10192), .B1(n27027), .B2(
        data_in[3]), .ZN(n10195) );
  INV_X1 U15339 ( .A(n10196), .ZN(n25278) );
  AOI22_X1 U15340 ( .A1(\mem[103][4] ), .A2(n10192), .B1(n27027), .B2(
        data_in[4]), .ZN(n10196) );
  INV_X1 U15341 ( .A(n10197), .ZN(n25277) );
  AOI22_X1 U15342 ( .A1(\mem[103][5] ), .A2(n10192), .B1(n27027), .B2(
        data_in[5]), .ZN(n10197) );
  INV_X1 U15343 ( .A(n10198), .ZN(n25276) );
  AOI22_X1 U15344 ( .A1(\mem[103][6] ), .A2(n10192), .B1(n27027), .B2(
        data_in[6]), .ZN(n10198) );
  INV_X1 U15345 ( .A(n10199), .ZN(n25275) );
  AOI22_X1 U15346 ( .A1(\mem[103][7] ), .A2(n10192), .B1(n27027), .B2(
        data_in[7]), .ZN(n10199) );
  INV_X1 U15347 ( .A(n10417), .ZN(n25082) );
  AOI22_X1 U15348 ( .A1(\mem[128][0] ), .A2(n10418), .B1(n27002), .B2(
        data_in[0]), .ZN(n10417) );
  INV_X1 U15349 ( .A(n10419), .ZN(n25081) );
  AOI22_X1 U15350 ( .A1(\mem[128][1] ), .A2(n10418), .B1(n27002), .B2(
        data_in[1]), .ZN(n10419) );
  INV_X1 U15351 ( .A(n10420), .ZN(n25080) );
  AOI22_X1 U15352 ( .A1(\mem[128][2] ), .A2(n10418), .B1(n27002), .B2(
        data_in[2]), .ZN(n10420) );
  INV_X1 U15353 ( .A(n10421), .ZN(n25079) );
  AOI22_X1 U15354 ( .A1(\mem[128][3] ), .A2(n10418), .B1(n27002), .B2(
        data_in[3]), .ZN(n10421) );
  INV_X1 U15355 ( .A(n10422), .ZN(n25078) );
  AOI22_X1 U15356 ( .A1(\mem[128][4] ), .A2(n10418), .B1(n27002), .B2(
        data_in[4]), .ZN(n10422) );
  INV_X1 U15357 ( .A(n10423), .ZN(n25077) );
  AOI22_X1 U15358 ( .A1(\mem[128][5] ), .A2(n10418), .B1(n27002), .B2(
        data_in[5]), .ZN(n10423) );
  INV_X1 U15359 ( .A(n10424), .ZN(n25076) );
  AOI22_X1 U15360 ( .A1(\mem[128][6] ), .A2(n10418), .B1(n27002), .B2(
        data_in[6]), .ZN(n10424) );
  INV_X1 U15361 ( .A(n10425), .ZN(n25075) );
  AOI22_X1 U15362 ( .A1(\mem[128][7] ), .A2(n10418), .B1(n27002), .B2(
        data_in[7]), .ZN(n10425) );
  INV_X1 U15363 ( .A(n10427), .ZN(n25074) );
  AOI22_X1 U15364 ( .A1(\mem[129][0] ), .A2(n10428), .B1(n27001), .B2(
        data_in[0]), .ZN(n10427) );
  INV_X1 U15365 ( .A(n10429), .ZN(n25073) );
  AOI22_X1 U15366 ( .A1(\mem[129][1] ), .A2(n10428), .B1(n27001), .B2(
        data_in[1]), .ZN(n10429) );
  INV_X1 U15367 ( .A(n10430), .ZN(n25072) );
  AOI22_X1 U15368 ( .A1(\mem[129][2] ), .A2(n10428), .B1(n27001), .B2(
        data_in[2]), .ZN(n10430) );
  INV_X1 U15369 ( .A(n10431), .ZN(n25071) );
  AOI22_X1 U15370 ( .A1(\mem[129][3] ), .A2(n10428), .B1(n27001), .B2(
        data_in[3]), .ZN(n10431) );
  INV_X1 U15371 ( .A(n10432), .ZN(n25070) );
  AOI22_X1 U15372 ( .A1(\mem[129][4] ), .A2(n10428), .B1(n27001), .B2(
        data_in[4]), .ZN(n10432) );
  INV_X1 U15373 ( .A(n10433), .ZN(n25069) );
  AOI22_X1 U15374 ( .A1(\mem[129][5] ), .A2(n10428), .B1(n27001), .B2(
        data_in[5]), .ZN(n10433) );
  INV_X1 U15375 ( .A(n10434), .ZN(n25068) );
  AOI22_X1 U15376 ( .A1(\mem[129][6] ), .A2(n10428), .B1(n27001), .B2(
        data_in[6]), .ZN(n10434) );
  INV_X1 U15377 ( .A(n10435), .ZN(n25067) );
  AOI22_X1 U15378 ( .A1(\mem[129][7] ), .A2(n10428), .B1(n27001), .B2(
        data_in[7]), .ZN(n10435) );
  INV_X1 U15379 ( .A(n10436), .ZN(n25066) );
  AOI22_X1 U15380 ( .A1(\mem[130][0] ), .A2(n10437), .B1(n27000), .B2(
        data_in[0]), .ZN(n10436) );
  INV_X1 U15381 ( .A(n10438), .ZN(n25065) );
  AOI22_X1 U15382 ( .A1(\mem[130][1] ), .A2(n10437), .B1(n27000), .B2(
        data_in[1]), .ZN(n10438) );
  INV_X1 U15383 ( .A(n10439), .ZN(n25064) );
  AOI22_X1 U15384 ( .A1(\mem[130][2] ), .A2(n10437), .B1(n27000), .B2(
        data_in[2]), .ZN(n10439) );
  INV_X1 U15385 ( .A(n10440), .ZN(n25063) );
  AOI22_X1 U15386 ( .A1(\mem[130][3] ), .A2(n10437), .B1(n27000), .B2(
        data_in[3]), .ZN(n10440) );
  INV_X1 U15387 ( .A(n10441), .ZN(n25062) );
  AOI22_X1 U15388 ( .A1(\mem[130][4] ), .A2(n10437), .B1(n27000), .B2(
        data_in[4]), .ZN(n10441) );
  INV_X1 U15389 ( .A(n10442), .ZN(n25061) );
  AOI22_X1 U15390 ( .A1(\mem[130][5] ), .A2(n10437), .B1(n27000), .B2(
        data_in[5]), .ZN(n10442) );
  INV_X1 U15391 ( .A(n10443), .ZN(n25060) );
  AOI22_X1 U15392 ( .A1(\mem[130][6] ), .A2(n10437), .B1(n27000), .B2(
        data_in[6]), .ZN(n10443) );
  INV_X1 U15393 ( .A(n10444), .ZN(n25059) );
  AOI22_X1 U15394 ( .A1(\mem[130][7] ), .A2(n10437), .B1(n27000), .B2(
        data_in[7]), .ZN(n10444) );
  INV_X1 U15395 ( .A(n10445), .ZN(n25058) );
  AOI22_X1 U15396 ( .A1(\mem[131][0] ), .A2(n10446), .B1(n26999), .B2(
        data_in[0]), .ZN(n10445) );
  INV_X1 U15397 ( .A(n10447), .ZN(n25057) );
  AOI22_X1 U15398 ( .A1(\mem[131][1] ), .A2(n10446), .B1(n26999), .B2(
        data_in[1]), .ZN(n10447) );
  INV_X1 U15399 ( .A(n10448), .ZN(n25056) );
  AOI22_X1 U15400 ( .A1(\mem[131][2] ), .A2(n10446), .B1(n26999), .B2(
        data_in[2]), .ZN(n10448) );
  INV_X1 U15401 ( .A(n10449), .ZN(n25055) );
  AOI22_X1 U15402 ( .A1(\mem[131][3] ), .A2(n10446), .B1(n26999), .B2(
        data_in[3]), .ZN(n10449) );
  INV_X1 U15403 ( .A(n10450), .ZN(n25054) );
  AOI22_X1 U15404 ( .A1(\mem[131][4] ), .A2(n10446), .B1(n26999), .B2(
        data_in[4]), .ZN(n10450) );
  INV_X1 U15405 ( .A(n10451), .ZN(n25053) );
  AOI22_X1 U15406 ( .A1(\mem[131][5] ), .A2(n10446), .B1(n26999), .B2(
        data_in[5]), .ZN(n10451) );
  INV_X1 U15407 ( .A(n10452), .ZN(n25052) );
  AOI22_X1 U15408 ( .A1(\mem[131][6] ), .A2(n10446), .B1(n26999), .B2(
        data_in[6]), .ZN(n10452) );
  INV_X1 U15409 ( .A(n10453), .ZN(n25051) );
  AOI22_X1 U15410 ( .A1(\mem[131][7] ), .A2(n10446), .B1(n26999), .B2(
        data_in[7]), .ZN(n10453) );
  INV_X1 U15411 ( .A(n10454), .ZN(n25050) );
  AOI22_X1 U15412 ( .A1(\mem[132][0] ), .A2(n10455), .B1(n26998), .B2(
        data_in[0]), .ZN(n10454) );
  INV_X1 U15413 ( .A(n10456), .ZN(n25049) );
  AOI22_X1 U15414 ( .A1(\mem[132][1] ), .A2(n10455), .B1(n26998), .B2(
        data_in[1]), .ZN(n10456) );
  INV_X1 U15415 ( .A(n10457), .ZN(n25048) );
  AOI22_X1 U15416 ( .A1(\mem[132][2] ), .A2(n10455), .B1(n26998), .B2(
        data_in[2]), .ZN(n10457) );
  INV_X1 U15417 ( .A(n10458), .ZN(n25047) );
  AOI22_X1 U15418 ( .A1(\mem[132][3] ), .A2(n10455), .B1(n26998), .B2(
        data_in[3]), .ZN(n10458) );
  INV_X1 U15419 ( .A(n10459), .ZN(n25046) );
  AOI22_X1 U15420 ( .A1(\mem[132][4] ), .A2(n10455), .B1(n26998), .B2(
        data_in[4]), .ZN(n10459) );
  INV_X1 U15421 ( .A(n10460), .ZN(n25045) );
  AOI22_X1 U15422 ( .A1(\mem[132][5] ), .A2(n10455), .B1(n26998), .B2(
        data_in[5]), .ZN(n10460) );
  INV_X1 U15423 ( .A(n10461), .ZN(n25044) );
  AOI22_X1 U15424 ( .A1(\mem[132][6] ), .A2(n10455), .B1(n26998), .B2(
        data_in[6]), .ZN(n10461) );
  INV_X1 U15425 ( .A(n10462), .ZN(n25043) );
  AOI22_X1 U15426 ( .A1(\mem[132][7] ), .A2(n10455), .B1(n26998), .B2(
        data_in[7]), .ZN(n10462) );
  INV_X1 U15427 ( .A(n10463), .ZN(n25042) );
  AOI22_X1 U15428 ( .A1(\mem[133][0] ), .A2(n10464), .B1(n26997), .B2(
        data_in[0]), .ZN(n10463) );
  INV_X1 U15429 ( .A(n10465), .ZN(n25041) );
  AOI22_X1 U15430 ( .A1(\mem[133][1] ), .A2(n10464), .B1(n26997), .B2(
        data_in[1]), .ZN(n10465) );
  INV_X1 U15431 ( .A(n10466), .ZN(n25040) );
  AOI22_X1 U15432 ( .A1(\mem[133][2] ), .A2(n10464), .B1(n26997), .B2(
        data_in[2]), .ZN(n10466) );
  INV_X1 U15433 ( .A(n10467), .ZN(n25039) );
  AOI22_X1 U15434 ( .A1(\mem[133][3] ), .A2(n10464), .B1(n26997), .B2(
        data_in[3]), .ZN(n10467) );
  INV_X1 U15435 ( .A(n10468), .ZN(n25038) );
  AOI22_X1 U15436 ( .A1(\mem[133][4] ), .A2(n10464), .B1(n26997), .B2(
        data_in[4]), .ZN(n10468) );
  INV_X1 U15437 ( .A(n10469), .ZN(n25037) );
  AOI22_X1 U15438 ( .A1(\mem[133][5] ), .A2(n10464), .B1(n26997), .B2(
        data_in[5]), .ZN(n10469) );
  INV_X1 U15439 ( .A(n10470), .ZN(n25036) );
  AOI22_X1 U15440 ( .A1(\mem[133][6] ), .A2(n10464), .B1(n26997), .B2(
        data_in[6]), .ZN(n10470) );
  INV_X1 U15441 ( .A(n10471), .ZN(n25035) );
  AOI22_X1 U15442 ( .A1(\mem[133][7] ), .A2(n10464), .B1(n26997), .B2(
        data_in[7]), .ZN(n10471) );
  INV_X1 U15443 ( .A(n10472), .ZN(n25034) );
  AOI22_X1 U15444 ( .A1(\mem[134][0] ), .A2(n10473), .B1(n26996), .B2(
        data_in[0]), .ZN(n10472) );
  INV_X1 U15445 ( .A(n10474), .ZN(n25033) );
  AOI22_X1 U15446 ( .A1(\mem[134][1] ), .A2(n10473), .B1(n26996), .B2(
        data_in[1]), .ZN(n10474) );
  INV_X1 U15447 ( .A(n10475), .ZN(n25032) );
  AOI22_X1 U15448 ( .A1(\mem[134][2] ), .A2(n10473), .B1(n26996), .B2(
        data_in[2]), .ZN(n10475) );
  INV_X1 U15449 ( .A(n10476), .ZN(n25031) );
  AOI22_X1 U15450 ( .A1(\mem[134][3] ), .A2(n10473), .B1(n26996), .B2(
        data_in[3]), .ZN(n10476) );
  INV_X1 U15451 ( .A(n10477), .ZN(n25030) );
  AOI22_X1 U15452 ( .A1(\mem[134][4] ), .A2(n10473), .B1(n26996), .B2(
        data_in[4]), .ZN(n10477) );
  INV_X1 U15453 ( .A(n10478), .ZN(n25029) );
  AOI22_X1 U15454 ( .A1(\mem[134][5] ), .A2(n10473), .B1(n26996), .B2(
        data_in[5]), .ZN(n10478) );
  INV_X1 U15455 ( .A(n10479), .ZN(n25028) );
  AOI22_X1 U15456 ( .A1(\mem[134][6] ), .A2(n10473), .B1(n26996), .B2(
        data_in[6]), .ZN(n10479) );
  INV_X1 U15457 ( .A(n10480), .ZN(n25027) );
  AOI22_X1 U15458 ( .A1(\mem[134][7] ), .A2(n10473), .B1(n26996), .B2(
        data_in[7]), .ZN(n10480) );
  INV_X1 U15459 ( .A(n10481), .ZN(n25026) );
  AOI22_X1 U15460 ( .A1(\mem[135][0] ), .A2(n10482), .B1(n26995), .B2(
        data_in[0]), .ZN(n10481) );
  INV_X1 U15461 ( .A(n10483), .ZN(n25025) );
  AOI22_X1 U15462 ( .A1(\mem[135][1] ), .A2(n10482), .B1(n26995), .B2(
        data_in[1]), .ZN(n10483) );
  INV_X1 U15463 ( .A(n10484), .ZN(n25024) );
  AOI22_X1 U15464 ( .A1(\mem[135][2] ), .A2(n10482), .B1(n26995), .B2(
        data_in[2]), .ZN(n10484) );
  INV_X1 U15465 ( .A(n10485), .ZN(n25023) );
  AOI22_X1 U15466 ( .A1(\mem[135][3] ), .A2(n10482), .B1(n26995), .B2(
        data_in[3]), .ZN(n10485) );
  INV_X1 U15467 ( .A(n10486), .ZN(n25022) );
  AOI22_X1 U15468 ( .A1(\mem[135][4] ), .A2(n10482), .B1(n26995), .B2(
        data_in[4]), .ZN(n10486) );
  INV_X1 U15469 ( .A(n10487), .ZN(n25021) );
  AOI22_X1 U15470 ( .A1(\mem[135][5] ), .A2(n10482), .B1(n26995), .B2(
        data_in[5]), .ZN(n10487) );
  INV_X1 U15471 ( .A(n10488), .ZN(n25020) );
  AOI22_X1 U15472 ( .A1(\mem[135][6] ), .A2(n10482), .B1(n26995), .B2(
        data_in[6]), .ZN(n10488) );
  INV_X1 U15473 ( .A(n10489), .ZN(n25019) );
  AOI22_X1 U15474 ( .A1(\mem[135][7] ), .A2(n10482), .B1(n26995), .B2(
        data_in[7]), .ZN(n10489) );
  INV_X1 U15475 ( .A(n10707), .ZN(n24826) );
  AOI22_X1 U15476 ( .A1(\mem[160][0] ), .A2(n10708), .B1(n26970), .B2(
        data_in[0]), .ZN(n10707) );
  INV_X1 U15477 ( .A(n10709), .ZN(n24825) );
  AOI22_X1 U15478 ( .A1(\mem[160][1] ), .A2(n10708), .B1(n26970), .B2(
        data_in[1]), .ZN(n10709) );
  INV_X1 U15479 ( .A(n10710), .ZN(n24824) );
  AOI22_X1 U15480 ( .A1(\mem[160][2] ), .A2(n10708), .B1(n26970), .B2(
        data_in[2]), .ZN(n10710) );
  INV_X1 U15481 ( .A(n10711), .ZN(n24823) );
  AOI22_X1 U15482 ( .A1(\mem[160][3] ), .A2(n10708), .B1(n26970), .B2(
        data_in[3]), .ZN(n10711) );
  INV_X1 U15483 ( .A(n10712), .ZN(n24822) );
  AOI22_X1 U15484 ( .A1(\mem[160][4] ), .A2(n10708), .B1(n26970), .B2(
        data_in[4]), .ZN(n10712) );
  INV_X1 U15485 ( .A(n10713), .ZN(n24821) );
  AOI22_X1 U15486 ( .A1(\mem[160][5] ), .A2(n10708), .B1(n26970), .B2(
        data_in[5]), .ZN(n10713) );
  INV_X1 U15487 ( .A(n10714), .ZN(n24820) );
  AOI22_X1 U15488 ( .A1(\mem[160][6] ), .A2(n10708), .B1(n26970), .B2(
        data_in[6]), .ZN(n10714) );
  INV_X1 U15489 ( .A(n10715), .ZN(n24819) );
  AOI22_X1 U15490 ( .A1(\mem[160][7] ), .A2(n10708), .B1(n26970), .B2(
        data_in[7]), .ZN(n10715) );
  INV_X1 U15491 ( .A(n10717), .ZN(n24818) );
  AOI22_X1 U15492 ( .A1(\mem[161][0] ), .A2(n10718), .B1(n26969), .B2(
        data_in[0]), .ZN(n10717) );
  INV_X1 U15493 ( .A(n10719), .ZN(n24817) );
  AOI22_X1 U15494 ( .A1(\mem[161][1] ), .A2(n10718), .B1(n26969), .B2(
        data_in[1]), .ZN(n10719) );
  INV_X1 U15495 ( .A(n10720), .ZN(n24816) );
  AOI22_X1 U15496 ( .A1(\mem[161][2] ), .A2(n10718), .B1(n26969), .B2(
        data_in[2]), .ZN(n10720) );
  INV_X1 U15497 ( .A(n10721), .ZN(n24815) );
  AOI22_X1 U15498 ( .A1(\mem[161][3] ), .A2(n10718), .B1(n26969), .B2(
        data_in[3]), .ZN(n10721) );
  INV_X1 U15499 ( .A(n10722), .ZN(n24814) );
  AOI22_X1 U15500 ( .A1(\mem[161][4] ), .A2(n10718), .B1(n26969), .B2(
        data_in[4]), .ZN(n10722) );
  INV_X1 U15501 ( .A(n10723), .ZN(n24813) );
  AOI22_X1 U15502 ( .A1(\mem[161][5] ), .A2(n10718), .B1(n26969), .B2(
        data_in[5]), .ZN(n10723) );
  INV_X1 U15503 ( .A(n10724), .ZN(n24812) );
  AOI22_X1 U15504 ( .A1(\mem[161][6] ), .A2(n10718), .B1(n26969), .B2(
        data_in[6]), .ZN(n10724) );
  INV_X1 U15505 ( .A(n10725), .ZN(n24811) );
  AOI22_X1 U15506 ( .A1(\mem[161][7] ), .A2(n10718), .B1(n26969), .B2(
        data_in[7]), .ZN(n10725) );
  INV_X1 U15507 ( .A(n10726), .ZN(n24810) );
  AOI22_X1 U15508 ( .A1(\mem[162][0] ), .A2(n10727), .B1(n26968), .B2(
        data_in[0]), .ZN(n10726) );
  INV_X1 U15509 ( .A(n10728), .ZN(n24809) );
  AOI22_X1 U15510 ( .A1(\mem[162][1] ), .A2(n10727), .B1(n26968), .B2(
        data_in[1]), .ZN(n10728) );
  INV_X1 U15511 ( .A(n10729), .ZN(n24808) );
  AOI22_X1 U15512 ( .A1(\mem[162][2] ), .A2(n10727), .B1(n26968), .B2(
        data_in[2]), .ZN(n10729) );
  INV_X1 U15513 ( .A(n10730), .ZN(n24807) );
  AOI22_X1 U15514 ( .A1(\mem[162][3] ), .A2(n10727), .B1(n26968), .B2(
        data_in[3]), .ZN(n10730) );
  INV_X1 U15515 ( .A(n10731), .ZN(n24806) );
  AOI22_X1 U15516 ( .A1(\mem[162][4] ), .A2(n10727), .B1(n26968), .B2(
        data_in[4]), .ZN(n10731) );
  INV_X1 U15517 ( .A(n10732), .ZN(n24805) );
  AOI22_X1 U15518 ( .A1(\mem[162][5] ), .A2(n10727), .B1(n26968), .B2(
        data_in[5]), .ZN(n10732) );
  INV_X1 U15519 ( .A(n10733), .ZN(n24804) );
  AOI22_X1 U15520 ( .A1(\mem[162][6] ), .A2(n10727), .B1(n26968), .B2(
        data_in[6]), .ZN(n10733) );
  INV_X1 U15521 ( .A(n10734), .ZN(n24803) );
  AOI22_X1 U15522 ( .A1(\mem[162][7] ), .A2(n10727), .B1(n26968), .B2(
        data_in[7]), .ZN(n10734) );
  INV_X1 U15523 ( .A(n10735), .ZN(n24802) );
  AOI22_X1 U15524 ( .A1(\mem[163][0] ), .A2(n10736), .B1(n26967), .B2(
        data_in[0]), .ZN(n10735) );
  INV_X1 U15525 ( .A(n10737), .ZN(n24801) );
  AOI22_X1 U15526 ( .A1(\mem[163][1] ), .A2(n10736), .B1(n26967), .B2(
        data_in[1]), .ZN(n10737) );
  INV_X1 U15527 ( .A(n10738), .ZN(n24800) );
  AOI22_X1 U15528 ( .A1(\mem[163][2] ), .A2(n10736), .B1(n26967), .B2(
        data_in[2]), .ZN(n10738) );
  INV_X1 U15529 ( .A(n10739), .ZN(n24799) );
  AOI22_X1 U15530 ( .A1(\mem[163][3] ), .A2(n10736), .B1(n26967), .B2(
        data_in[3]), .ZN(n10739) );
  INV_X1 U15531 ( .A(n10740), .ZN(n24798) );
  AOI22_X1 U15532 ( .A1(\mem[163][4] ), .A2(n10736), .B1(n26967), .B2(
        data_in[4]), .ZN(n10740) );
  INV_X1 U15533 ( .A(n10741), .ZN(n24797) );
  AOI22_X1 U15534 ( .A1(\mem[163][5] ), .A2(n10736), .B1(n26967), .B2(
        data_in[5]), .ZN(n10741) );
  INV_X1 U15535 ( .A(n10742), .ZN(n24796) );
  AOI22_X1 U15536 ( .A1(\mem[163][6] ), .A2(n10736), .B1(n26967), .B2(
        data_in[6]), .ZN(n10742) );
  INV_X1 U15537 ( .A(n10743), .ZN(n24795) );
  AOI22_X1 U15538 ( .A1(\mem[163][7] ), .A2(n10736), .B1(n26967), .B2(
        data_in[7]), .ZN(n10743) );
  INV_X1 U15539 ( .A(n10744), .ZN(n24794) );
  AOI22_X1 U15540 ( .A1(\mem[164][0] ), .A2(n10745), .B1(n26966), .B2(
        data_in[0]), .ZN(n10744) );
  INV_X1 U15541 ( .A(n10746), .ZN(n24793) );
  AOI22_X1 U15542 ( .A1(\mem[164][1] ), .A2(n10745), .B1(n26966), .B2(
        data_in[1]), .ZN(n10746) );
  INV_X1 U15543 ( .A(n10747), .ZN(n24792) );
  AOI22_X1 U15544 ( .A1(\mem[164][2] ), .A2(n10745), .B1(n26966), .B2(
        data_in[2]), .ZN(n10747) );
  INV_X1 U15545 ( .A(n10748), .ZN(n24791) );
  AOI22_X1 U15546 ( .A1(\mem[164][3] ), .A2(n10745), .B1(n26966), .B2(
        data_in[3]), .ZN(n10748) );
  INV_X1 U15547 ( .A(n10749), .ZN(n24790) );
  AOI22_X1 U15548 ( .A1(\mem[164][4] ), .A2(n10745), .B1(n26966), .B2(
        data_in[4]), .ZN(n10749) );
  INV_X1 U15549 ( .A(n10750), .ZN(n24789) );
  AOI22_X1 U15550 ( .A1(\mem[164][5] ), .A2(n10745), .B1(n26966), .B2(
        data_in[5]), .ZN(n10750) );
  INV_X1 U15551 ( .A(n10751), .ZN(n24788) );
  AOI22_X1 U15552 ( .A1(\mem[164][6] ), .A2(n10745), .B1(n26966), .B2(
        data_in[6]), .ZN(n10751) );
  INV_X1 U15553 ( .A(n10752), .ZN(n24787) );
  AOI22_X1 U15554 ( .A1(\mem[164][7] ), .A2(n10745), .B1(n26966), .B2(
        data_in[7]), .ZN(n10752) );
  INV_X1 U15555 ( .A(n10753), .ZN(n24786) );
  AOI22_X1 U15556 ( .A1(\mem[165][0] ), .A2(n10754), .B1(n26965), .B2(
        data_in[0]), .ZN(n10753) );
  INV_X1 U15557 ( .A(n10755), .ZN(n24785) );
  AOI22_X1 U15558 ( .A1(\mem[165][1] ), .A2(n10754), .B1(n26965), .B2(
        data_in[1]), .ZN(n10755) );
  INV_X1 U15559 ( .A(n10756), .ZN(n24784) );
  AOI22_X1 U15560 ( .A1(\mem[165][2] ), .A2(n10754), .B1(n26965), .B2(
        data_in[2]), .ZN(n10756) );
  INV_X1 U15561 ( .A(n10757), .ZN(n24783) );
  AOI22_X1 U15562 ( .A1(\mem[165][3] ), .A2(n10754), .B1(n26965), .B2(
        data_in[3]), .ZN(n10757) );
  INV_X1 U15563 ( .A(n10758), .ZN(n24782) );
  AOI22_X1 U15564 ( .A1(\mem[165][4] ), .A2(n10754), .B1(n26965), .B2(
        data_in[4]), .ZN(n10758) );
  INV_X1 U15565 ( .A(n10759), .ZN(n24781) );
  AOI22_X1 U15566 ( .A1(\mem[165][5] ), .A2(n10754), .B1(n26965), .B2(
        data_in[5]), .ZN(n10759) );
  INV_X1 U15567 ( .A(n10760), .ZN(n24780) );
  AOI22_X1 U15568 ( .A1(\mem[165][6] ), .A2(n10754), .B1(n26965), .B2(
        data_in[6]), .ZN(n10760) );
  INV_X1 U15569 ( .A(n10761), .ZN(n24779) );
  AOI22_X1 U15570 ( .A1(\mem[165][7] ), .A2(n10754), .B1(n26965), .B2(
        data_in[7]), .ZN(n10761) );
  INV_X1 U15571 ( .A(n10762), .ZN(n24778) );
  AOI22_X1 U15572 ( .A1(\mem[166][0] ), .A2(n10763), .B1(n26964), .B2(
        data_in[0]), .ZN(n10762) );
  INV_X1 U15573 ( .A(n10764), .ZN(n24777) );
  AOI22_X1 U15574 ( .A1(\mem[166][1] ), .A2(n10763), .B1(n26964), .B2(
        data_in[1]), .ZN(n10764) );
  INV_X1 U15575 ( .A(n10765), .ZN(n24776) );
  AOI22_X1 U15576 ( .A1(\mem[166][2] ), .A2(n10763), .B1(n26964), .B2(
        data_in[2]), .ZN(n10765) );
  INV_X1 U15577 ( .A(n10766), .ZN(n24775) );
  AOI22_X1 U15578 ( .A1(\mem[166][3] ), .A2(n10763), .B1(n26964), .B2(
        data_in[3]), .ZN(n10766) );
  INV_X1 U15579 ( .A(n10767), .ZN(n24774) );
  AOI22_X1 U15580 ( .A1(\mem[166][4] ), .A2(n10763), .B1(n26964), .B2(
        data_in[4]), .ZN(n10767) );
  INV_X1 U15581 ( .A(n10768), .ZN(n24773) );
  AOI22_X1 U15582 ( .A1(\mem[166][5] ), .A2(n10763), .B1(n26964), .B2(
        data_in[5]), .ZN(n10768) );
  INV_X1 U15583 ( .A(n10769), .ZN(n24772) );
  AOI22_X1 U15584 ( .A1(\mem[166][6] ), .A2(n10763), .B1(n26964), .B2(
        data_in[6]), .ZN(n10769) );
  INV_X1 U15585 ( .A(n10770), .ZN(n24771) );
  AOI22_X1 U15586 ( .A1(\mem[166][7] ), .A2(n10763), .B1(n26964), .B2(
        data_in[7]), .ZN(n10770) );
  INV_X1 U15587 ( .A(n10771), .ZN(n24770) );
  AOI22_X1 U15588 ( .A1(\mem[167][0] ), .A2(n10772), .B1(n26963), .B2(
        data_in[0]), .ZN(n10771) );
  INV_X1 U15589 ( .A(n10773), .ZN(n24769) );
  AOI22_X1 U15590 ( .A1(\mem[167][1] ), .A2(n10772), .B1(n26963), .B2(
        data_in[1]), .ZN(n10773) );
  INV_X1 U15591 ( .A(n10774), .ZN(n24768) );
  AOI22_X1 U15592 ( .A1(\mem[167][2] ), .A2(n10772), .B1(n26963), .B2(
        data_in[2]), .ZN(n10774) );
  INV_X1 U15593 ( .A(n10775), .ZN(n24767) );
  AOI22_X1 U15594 ( .A1(\mem[167][3] ), .A2(n10772), .B1(n26963), .B2(
        data_in[3]), .ZN(n10775) );
  INV_X1 U15595 ( .A(n10776), .ZN(n24766) );
  AOI22_X1 U15596 ( .A1(\mem[167][4] ), .A2(n10772), .B1(n26963), .B2(
        data_in[4]), .ZN(n10776) );
  INV_X1 U15597 ( .A(n10777), .ZN(n24765) );
  AOI22_X1 U15598 ( .A1(\mem[167][5] ), .A2(n10772), .B1(n26963), .B2(
        data_in[5]), .ZN(n10777) );
  INV_X1 U15599 ( .A(n10778), .ZN(n24764) );
  AOI22_X1 U15600 ( .A1(\mem[167][6] ), .A2(n10772), .B1(n26963), .B2(
        data_in[6]), .ZN(n10778) );
  INV_X1 U15601 ( .A(n10779), .ZN(n24763) );
  AOI22_X1 U15602 ( .A1(\mem[167][7] ), .A2(n10772), .B1(n26963), .B2(
        data_in[7]), .ZN(n10779) );
  INV_X1 U15603 ( .A(n10997), .ZN(n24570) );
  AOI22_X1 U15604 ( .A1(\mem[192][0] ), .A2(n10998), .B1(n26938), .B2(
        data_in[0]), .ZN(n10997) );
  INV_X1 U15605 ( .A(n10999), .ZN(n24569) );
  AOI22_X1 U15606 ( .A1(\mem[192][1] ), .A2(n10998), .B1(n26938), .B2(
        data_in[1]), .ZN(n10999) );
  INV_X1 U15607 ( .A(n11000), .ZN(n24568) );
  AOI22_X1 U15608 ( .A1(\mem[192][2] ), .A2(n10998), .B1(n26938), .B2(
        data_in[2]), .ZN(n11000) );
  INV_X1 U15609 ( .A(n11001), .ZN(n24567) );
  AOI22_X1 U15610 ( .A1(\mem[192][3] ), .A2(n10998), .B1(n26938), .B2(
        data_in[3]), .ZN(n11001) );
  INV_X1 U15611 ( .A(n11002), .ZN(n24566) );
  AOI22_X1 U15612 ( .A1(\mem[192][4] ), .A2(n10998), .B1(n26938), .B2(
        data_in[4]), .ZN(n11002) );
  INV_X1 U15613 ( .A(n11003), .ZN(n24565) );
  AOI22_X1 U15614 ( .A1(\mem[192][5] ), .A2(n10998), .B1(n26938), .B2(
        data_in[5]), .ZN(n11003) );
  INV_X1 U15615 ( .A(n11004), .ZN(n24564) );
  AOI22_X1 U15616 ( .A1(\mem[192][6] ), .A2(n10998), .B1(n26938), .B2(
        data_in[6]), .ZN(n11004) );
  INV_X1 U15617 ( .A(n11005), .ZN(n24563) );
  AOI22_X1 U15618 ( .A1(\mem[192][7] ), .A2(n10998), .B1(n26938), .B2(
        data_in[7]), .ZN(n11005) );
  INV_X1 U15619 ( .A(n11007), .ZN(n24562) );
  AOI22_X1 U15620 ( .A1(\mem[193][0] ), .A2(n11008), .B1(n26937), .B2(
        data_in[0]), .ZN(n11007) );
  INV_X1 U15621 ( .A(n11009), .ZN(n24561) );
  AOI22_X1 U15622 ( .A1(\mem[193][1] ), .A2(n11008), .B1(n26937), .B2(
        data_in[1]), .ZN(n11009) );
  INV_X1 U15623 ( .A(n11010), .ZN(n24560) );
  AOI22_X1 U15624 ( .A1(\mem[193][2] ), .A2(n11008), .B1(n26937), .B2(
        data_in[2]), .ZN(n11010) );
  INV_X1 U15625 ( .A(n11011), .ZN(n24559) );
  AOI22_X1 U15626 ( .A1(\mem[193][3] ), .A2(n11008), .B1(n26937), .B2(
        data_in[3]), .ZN(n11011) );
  INV_X1 U15627 ( .A(n11012), .ZN(n24558) );
  AOI22_X1 U15628 ( .A1(\mem[193][4] ), .A2(n11008), .B1(n26937), .B2(
        data_in[4]), .ZN(n11012) );
  INV_X1 U15629 ( .A(n11013), .ZN(n24557) );
  AOI22_X1 U15630 ( .A1(\mem[193][5] ), .A2(n11008), .B1(n26937), .B2(
        data_in[5]), .ZN(n11013) );
  INV_X1 U15631 ( .A(n11014), .ZN(n24556) );
  AOI22_X1 U15632 ( .A1(\mem[193][6] ), .A2(n11008), .B1(n26937), .B2(
        data_in[6]), .ZN(n11014) );
  INV_X1 U15633 ( .A(n11015), .ZN(n24555) );
  AOI22_X1 U15634 ( .A1(\mem[193][7] ), .A2(n11008), .B1(n26937), .B2(
        data_in[7]), .ZN(n11015) );
  INV_X1 U15635 ( .A(n11016), .ZN(n24554) );
  AOI22_X1 U15636 ( .A1(\mem[194][0] ), .A2(n11017), .B1(n26936), .B2(
        data_in[0]), .ZN(n11016) );
  INV_X1 U15637 ( .A(n11018), .ZN(n24553) );
  AOI22_X1 U15638 ( .A1(\mem[194][1] ), .A2(n11017), .B1(n26936), .B2(
        data_in[1]), .ZN(n11018) );
  INV_X1 U15639 ( .A(n11019), .ZN(n24552) );
  AOI22_X1 U15640 ( .A1(\mem[194][2] ), .A2(n11017), .B1(n26936), .B2(
        data_in[2]), .ZN(n11019) );
  INV_X1 U15641 ( .A(n11020), .ZN(n24551) );
  AOI22_X1 U15642 ( .A1(\mem[194][3] ), .A2(n11017), .B1(n26936), .B2(
        data_in[3]), .ZN(n11020) );
  INV_X1 U15643 ( .A(n11021), .ZN(n24550) );
  AOI22_X1 U15644 ( .A1(\mem[194][4] ), .A2(n11017), .B1(n26936), .B2(
        data_in[4]), .ZN(n11021) );
  INV_X1 U15645 ( .A(n11022), .ZN(n24549) );
  AOI22_X1 U15646 ( .A1(\mem[194][5] ), .A2(n11017), .B1(n26936), .B2(
        data_in[5]), .ZN(n11022) );
  INV_X1 U15647 ( .A(n11023), .ZN(n24548) );
  AOI22_X1 U15648 ( .A1(\mem[194][6] ), .A2(n11017), .B1(n26936), .B2(
        data_in[6]), .ZN(n11023) );
  INV_X1 U15649 ( .A(n11024), .ZN(n24547) );
  AOI22_X1 U15650 ( .A1(\mem[194][7] ), .A2(n11017), .B1(n26936), .B2(
        data_in[7]), .ZN(n11024) );
  INV_X1 U15651 ( .A(n11025), .ZN(n24546) );
  AOI22_X1 U15652 ( .A1(\mem[195][0] ), .A2(n11026), .B1(n26935), .B2(
        data_in[0]), .ZN(n11025) );
  INV_X1 U15653 ( .A(n11027), .ZN(n24545) );
  AOI22_X1 U15654 ( .A1(\mem[195][1] ), .A2(n11026), .B1(n26935), .B2(
        data_in[1]), .ZN(n11027) );
  INV_X1 U15655 ( .A(n11028), .ZN(n24544) );
  AOI22_X1 U15656 ( .A1(\mem[195][2] ), .A2(n11026), .B1(n26935), .B2(
        data_in[2]), .ZN(n11028) );
  INV_X1 U15657 ( .A(n11029), .ZN(n24543) );
  AOI22_X1 U15658 ( .A1(\mem[195][3] ), .A2(n11026), .B1(n26935), .B2(
        data_in[3]), .ZN(n11029) );
  INV_X1 U15659 ( .A(n11030), .ZN(n24542) );
  AOI22_X1 U15660 ( .A1(\mem[195][4] ), .A2(n11026), .B1(n26935), .B2(
        data_in[4]), .ZN(n11030) );
  INV_X1 U15661 ( .A(n11031), .ZN(n24541) );
  AOI22_X1 U15662 ( .A1(\mem[195][5] ), .A2(n11026), .B1(n26935), .B2(
        data_in[5]), .ZN(n11031) );
  INV_X1 U15663 ( .A(n11032), .ZN(n24540) );
  AOI22_X1 U15664 ( .A1(\mem[195][6] ), .A2(n11026), .B1(n26935), .B2(
        data_in[6]), .ZN(n11032) );
  INV_X1 U15665 ( .A(n11033), .ZN(n24539) );
  AOI22_X1 U15666 ( .A1(\mem[195][7] ), .A2(n11026), .B1(n26935), .B2(
        data_in[7]), .ZN(n11033) );
  INV_X1 U15667 ( .A(n11034), .ZN(n24538) );
  AOI22_X1 U15668 ( .A1(\mem[196][0] ), .A2(n11035), .B1(n26934), .B2(
        data_in[0]), .ZN(n11034) );
  INV_X1 U15669 ( .A(n11036), .ZN(n24537) );
  AOI22_X1 U15670 ( .A1(\mem[196][1] ), .A2(n11035), .B1(n26934), .B2(
        data_in[1]), .ZN(n11036) );
  INV_X1 U15671 ( .A(n11037), .ZN(n24536) );
  AOI22_X1 U15672 ( .A1(\mem[196][2] ), .A2(n11035), .B1(n26934), .B2(
        data_in[2]), .ZN(n11037) );
  INV_X1 U15673 ( .A(n11038), .ZN(n24535) );
  AOI22_X1 U15674 ( .A1(\mem[196][3] ), .A2(n11035), .B1(n26934), .B2(
        data_in[3]), .ZN(n11038) );
  INV_X1 U15675 ( .A(n11039), .ZN(n24534) );
  AOI22_X1 U15676 ( .A1(\mem[196][4] ), .A2(n11035), .B1(n26934), .B2(
        data_in[4]), .ZN(n11039) );
  INV_X1 U15677 ( .A(n11040), .ZN(n24533) );
  AOI22_X1 U15678 ( .A1(\mem[196][5] ), .A2(n11035), .B1(n26934), .B2(
        data_in[5]), .ZN(n11040) );
  INV_X1 U15679 ( .A(n11041), .ZN(n24532) );
  AOI22_X1 U15680 ( .A1(\mem[196][6] ), .A2(n11035), .B1(n26934), .B2(
        data_in[6]), .ZN(n11041) );
  INV_X1 U15681 ( .A(n11042), .ZN(n24531) );
  AOI22_X1 U15682 ( .A1(\mem[196][7] ), .A2(n11035), .B1(n26934), .B2(
        data_in[7]), .ZN(n11042) );
  INV_X1 U15683 ( .A(n11043), .ZN(n24530) );
  AOI22_X1 U15684 ( .A1(\mem[197][0] ), .A2(n11044), .B1(n26933), .B2(
        data_in[0]), .ZN(n11043) );
  INV_X1 U15685 ( .A(n11045), .ZN(n24529) );
  AOI22_X1 U15686 ( .A1(\mem[197][1] ), .A2(n11044), .B1(n26933), .B2(
        data_in[1]), .ZN(n11045) );
  INV_X1 U15687 ( .A(n11046), .ZN(n24528) );
  AOI22_X1 U15688 ( .A1(\mem[197][2] ), .A2(n11044), .B1(n26933), .B2(
        data_in[2]), .ZN(n11046) );
  INV_X1 U15689 ( .A(n11047), .ZN(n24527) );
  AOI22_X1 U15690 ( .A1(\mem[197][3] ), .A2(n11044), .B1(n26933), .B2(
        data_in[3]), .ZN(n11047) );
  INV_X1 U15691 ( .A(n11048), .ZN(n24526) );
  AOI22_X1 U15692 ( .A1(\mem[197][4] ), .A2(n11044), .B1(n26933), .B2(
        data_in[4]), .ZN(n11048) );
  INV_X1 U15693 ( .A(n11049), .ZN(n24525) );
  AOI22_X1 U15694 ( .A1(\mem[197][5] ), .A2(n11044), .B1(n26933), .B2(
        data_in[5]), .ZN(n11049) );
  INV_X1 U15695 ( .A(n11050), .ZN(n24524) );
  AOI22_X1 U15696 ( .A1(\mem[197][6] ), .A2(n11044), .B1(n26933), .B2(
        data_in[6]), .ZN(n11050) );
  INV_X1 U15697 ( .A(n11051), .ZN(n24523) );
  AOI22_X1 U15698 ( .A1(\mem[197][7] ), .A2(n11044), .B1(n26933), .B2(
        data_in[7]), .ZN(n11051) );
  INV_X1 U15699 ( .A(n11052), .ZN(n24522) );
  AOI22_X1 U15700 ( .A1(\mem[198][0] ), .A2(n11053), .B1(n26932), .B2(
        data_in[0]), .ZN(n11052) );
  INV_X1 U15701 ( .A(n11054), .ZN(n24521) );
  AOI22_X1 U15702 ( .A1(\mem[198][1] ), .A2(n11053), .B1(n26932), .B2(
        data_in[1]), .ZN(n11054) );
  INV_X1 U15703 ( .A(n11055), .ZN(n24520) );
  AOI22_X1 U15704 ( .A1(\mem[198][2] ), .A2(n11053), .B1(n26932), .B2(
        data_in[2]), .ZN(n11055) );
  INV_X1 U15705 ( .A(n11056), .ZN(n24519) );
  AOI22_X1 U15706 ( .A1(\mem[198][3] ), .A2(n11053), .B1(n26932), .B2(
        data_in[3]), .ZN(n11056) );
  INV_X1 U15707 ( .A(n11057), .ZN(n24518) );
  AOI22_X1 U15708 ( .A1(\mem[198][4] ), .A2(n11053), .B1(n26932), .B2(
        data_in[4]), .ZN(n11057) );
  INV_X1 U15709 ( .A(n11058), .ZN(n24517) );
  AOI22_X1 U15710 ( .A1(\mem[198][5] ), .A2(n11053), .B1(n26932), .B2(
        data_in[5]), .ZN(n11058) );
  INV_X1 U15711 ( .A(n11059), .ZN(n24516) );
  AOI22_X1 U15712 ( .A1(\mem[198][6] ), .A2(n11053), .B1(n26932), .B2(
        data_in[6]), .ZN(n11059) );
  INV_X1 U15713 ( .A(n11060), .ZN(n24515) );
  AOI22_X1 U15714 ( .A1(\mem[198][7] ), .A2(n11053), .B1(n26932), .B2(
        data_in[7]), .ZN(n11060) );
  INV_X1 U15715 ( .A(n11061), .ZN(n24514) );
  AOI22_X1 U15716 ( .A1(\mem[199][0] ), .A2(n11062), .B1(n26931), .B2(
        data_in[0]), .ZN(n11061) );
  INV_X1 U15717 ( .A(n11063), .ZN(n24513) );
  AOI22_X1 U15718 ( .A1(\mem[199][1] ), .A2(n11062), .B1(n26931), .B2(
        data_in[1]), .ZN(n11063) );
  INV_X1 U15719 ( .A(n11064), .ZN(n24512) );
  AOI22_X1 U15720 ( .A1(\mem[199][2] ), .A2(n11062), .B1(n26931), .B2(
        data_in[2]), .ZN(n11064) );
  INV_X1 U15721 ( .A(n11065), .ZN(n24511) );
  AOI22_X1 U15722 ( .A1(\mem[199][3] ), .A2(n11062), .B1(n26931), .B2(
        data_in[3]), .ZN(n11065) );
  INV_X1 U15723 ( .A(n11066), .ZN(n24510) );
  AOI22_X1 U15724 ( .A1(\mem[199][4] ), .A2(n11062), .B1(n26931), .B2(
        data_in[4]), .ZN(n11066) );
  INV_X1 U15725 ( .A(n11067), .ZN(n24509) );
  AOI22_X1 U15726 ( .A1(\mem[199][5] ), .A2(n11062), .B1(n26931), .B2(
        data_in[5]), .ZN(n11067) );
  INV_X1 U15727 ( .A(n11068), .ZN(n24508) );
  AOI22_X1 U15728 ( .A1(\mem[199][6] ), .A2(n11062), .B1(n26931), .B2(
        data_in[6]), .ZN(n11068) );
  INV_X1 U15729 ( .A(n11069), .ZN(n24507) );
  AOI22_X1 U15730 ( .A1(\mem[199][7] ), .A2(n11062), .B1(n26931), .B2(
        data_in[7]), .ZN(n11069) );
  INV_X1 U15731 ( .A(n11287), .ZN(n24314) );
  AOI22_X1 U15732 ( .A1(\mem[224][0] ), .A2(n11288), .B1(n26906), .B2(
        data_in[0]), .ZN(n11287) );
  INV_X1 U15733 ( .A(n11289), .ZN(n24313) );
  AOI22_X1 U15734 ( .A1(\mem[224][1] ), .A2(n11288), .B1(n26906), .B2(
        data_in[1]), .ZN(n11289) );
  INV_X1 U15735 ( .A(n11290), .ZN(n24312) );
  AOI22_X1 U15736 ( .A1(\mem[224][2] ), .A2(n11288), .B1(n26906), .B2(
        data_in[2]), .ZN(n11290) );
  INV_X1 U15737 ( .A(n11291), .ZN(n24311) );
  AOI22_X1 U15738 ( .A1(\mem[224][3] ), .A2(n11288), .B1(n26906), .B2(
        data_in[3]), .ZN(n11291) );
  INV_X1 U15739 ( .A(n11292), .ZN(n24310) );
  AOI22_X1 U15740 ( .A1(\mem[224][4] ), .A2(n11288), .B1(n26906), .B2(
        data_in[4]), .ZN(n11292) );
  INV_X1 U15741 ( .A(n11293), .ZN(n24309) );
  AOI22_X1 U15742 ( .A1(\mem[224][5] ), .A2(n11288), .B1(n26906), .B2(
        data_in[5]), .ZN(n11293) );
  INV_X1 U15743 ( .A(n11294), .ZN(n24308) );
  AOI22_X1 U15744 ( .A1(\mem[224][6] ), .A2(n11288), .B1(n26906), .B2(
        data_in[6]), .ZN(n11294) );
  INV_X1 U15745 ( .A(n11295), .ZN(n24307) );
  AOI22_X1 U15746 ( .A1(\mem[224][7] ), .A2(n11288), .B1(n26906), .B2(
        data_in[7]), .ZN(n11295) );
  INV_X1 U15747 ( .A(n11297), .ZN(n24306) );
  AOI22_X1 U15748 ( .A1(\mem[225][0] ), .A2(n11298), .B1(n26905), .B2(
        data_in[0]), .ZN(n11297) );
  INV_X1 U15749 ( .A(n11299), .ZN(n24305) );
  AOI22_X1 U15750 ( .A1(\mem[225][1] ), .A2(n11298), .B1(n26905), .B2(
        data_in[1]), .ZN(n11299) );
  INV_X1 U15751 ( .A(n11300), .ZN(n24304) );
  AOI22_X1 U15752 ( .A1(\mem[225][2] ), .A2(n11298), .B1(n26905), .B2(
        data_in[2]), .ZN(n11300) );
  INV_X1 U15753 ( .A(n11301), .ZN(n24303) );
  AOI22_X1 U15754 ( .A1(\mem[225][3] ), .A2(n11298), .B1(n26905), .B2(
        data_in[3]), .ZN(n11301) );
  INV_X1 U15755 ( .A(n11302), .ZN(n24302) );
  AOI22_X1 U15756 ( .A1(\mem[225][4] ), .A2(n11298), .B1(n26905), .B2(
        data_in[4]), .ZN(n11302) );
  INV_X1 U15757 ( .A(n11303), .ZN(n24301) );
  AOI22_X1 U15758 ( .A1(\mem[225][5] ), .A2(n11298), .B1(n26905), .B2(
        data_in[5]), .ZN(n11303) );
  INV_X1 U15759 ( .A(n11304), .ZN(n24300) );
  AOI22_X1 U15760 ( .A1(\mem[225][6] ), .A2(n11298), .B1(n26905), .B2(
        data_in[6]), .ZN(n11304) );
  INV_X1 U15761 ( .A(n11305), .ZN(n24299) );
  AOI22_X1 U15762 ( .A1(\mem[225][7] ), .A2(n11298), .B1(n26905), .B2(
        data_in[7]), .ZN(n11305) );
  INV_X1 U15763 ( .A(n11306), .ZN(n24298) );
  AOI22_X1 U15764 ( .A1(\mem[226][0] ), .A2(n11307), .B1(n26904), .B2(
        data_in[0]), .ZN(n11306) );
  INV_X1 U15765 ( .A(n11308), .ZN(n24297) );
  AOI22_X1 U15766 ( .A1(\mem[226][1] ), .A2(n11307), .B1(n26904), .B2(
        data_in[1]), .ZN(n11308) );
  INV_X1 U15767 ( .A(n11309), .ZN(n24296) );
  AOI22_X1 U15768 ( .A1(\mem[226][2] ), .A2(n11307), .B1(n26904), .B2(
        data_in[2]), .ZN(n11309) );
  INV_X1 U15769 ( .A(n11310), .ZN(n24295) );
  AOI22_X1 U15770 ( .A1(\mem[226][3] ), .A2(n11307), .B1(n26904), .B2(
        data_in[3]), .ZN(n11310) );
  INV_X1 U15771 ( .A(n11311), .ZN(n24294) );
  AOI22_X1 U15772 ( .A1(\mem[226][4] ), .A2(n11307), .B1(n26904), .B2(
        data_in[4]), .ZN(n11311) );
  INV_X1 U15773 ( .A(n11312), .ZN(n24293) );
  AOI22_X1 U15774 ( .A1(\mem[226][5] ), .A2(n11307), .B1(n26904), .B2(
        data_in[5]), .ZN(n11312) );
  INV_X1 U15775 ( .A(n11313), .ZN(n24292) );
  AOI22_X1 U15776 ( .A1(\mem[226][6] ), .A2(n11307), .B1(n26904), .B2(
        data_in[6]), .ZN(n11313) );
  INV_X1 U15777 ( .A(n11314), .ZN(n24291) );
  AOI22_X1 U15778 ( .A1(\mem[226][7] ), .A2(n11307), .B1(n26904), .B2(
        data_in[7]), .ZN(n11314) );
  INV_X1 U15779 ( .A(n11315), .ZN(n24290) );
  AOI22_X1 U15780 ( .A1(\mem[227][0] ), .A2(n11316), .B1(n26903), .B2(
        data_in[0]), .ZN(n11315) );
  INV_X1 U15781 ( .A(n11317), .ZN(n24289) );
  AOI22_X1 U15782 ( .A1(\mem[227][1] ), .A2(n11316), .B1(n26903), .B2(
        data_in[1]), .ZN(n11317) );
  INV_X1 U15783 ( .A(n11318), .ZN(n24288) );
  AOI22_X1 U15784 ( .A1(\mem[227][2] ), .A2(n11316), .B1(n26903), .B2(
        data_in[2]), .ZN(n11318) );
  INV_X1 U15785 ( .A(n11319), .ZN(n24287) );
  AOI22_X1 U15786 ( .A1(\mem[227][3] ), .A2(n11316), .B1(n26903), .B2(
        data_in[3]), .ZN(n11319) );
  INV_X1 U15787 ( .A(n11320), .ZN(n24286) );
  AOI22_X1 U15788 ( .A1(\mem[227][4] ), .A2(n11316), .B1(n26903), .B2(
        data_in[4]), .ZN(n11320) );
  INV_X1 U15789 ( .A(n11321), .ZN(n24285) );
  AOI22_X1 U15790 ( .A1(\mem[227][5] ), .A2(n11316), .B1(n26903), .B2(
        data_in[5]), .ZN(n11321) );
  INV_X1 U15791 ( .A(n11322), .ZN(n24284) );
  AOI22_X1 U15792 ( .A1(\mem[227][6] ), .A2(n11316), .B1(n26903), .B2(
        data_in[6]), .ZN(n11322) );
  INV_X1 U15793 ( .A(n11323), .ZN(n24283) );
  AOI22_X1 U15794 ( .A1(\mem[227][7] ), .A2(n11316), .B1(n26903), .B2(
        data_in[7]), .ZN(n11323) );
  INV_X1 U15795 ( .A(n11324), .ZN(n24282) );
  AOI22_X1 U15796 ( .A1(\mem[228][0] ), .A2(n11325), .B1(n26902), .B2(
        data_in[0]), .ZN(n11324) );
  INV_X1 U15797 ( .A(n11326), .ZN(n24281) );
  AOI22_X1 U15798 ( .A1(\mem[228][1] ), .A2(n11325), .B1(n26902), .B2(
        data_in[1]), .ZN(n11326) );
  INV_X1 U15799 ( .A(n11327), .ZN(n24280) );
  AOI22_X1 U15800 ( .A1(\mem[228][2] ), .A2(n11325), .B1(n26902), .B2(
        data_in[2]), .ZN(n11327) );
  INV_X1 U15801 ( .A(n11328), .ZN(n24279) );
  AOI22_X1 U15802 ( .A1(\mem[228][3] ), .A2(n11325), .B1(n26902), .B2(
        data_in[3]), .ZN(n11328) );
  INV_X1 U15803 ( .A(n11329), .ZN(n24278) );
  AOI22_X1 U15804 ( .A1(\mem[228][4] ), .A2(n11325), .B1(n26902), .B2(
        data_in[4]), .ZN(n11329) );
  INV_X1 U15805 ( .A(n11330), .ZN(n24277) );
  AOI22_X1 U15806 ( .A1(\mem[228][5] ), .A2(n11325), .B1(n26902), .B2(
        data_in[5]), .ZN(n11330) );
  INV_X1 U15807 ( .A(n11331), .ZN(n24276) );
  AOI22_X1 U15808 ( .A1(\mem[228][6] ), .A2(n11325), .B1(n26902), .B2(
        data_in[6]), .ZN(n11331) );
  INV_X1 U15809 ( .A(n11332), .ZN(n24275) );
  AOI22_X1 U15810 ( .A1(\mem[228][7] ), .A2(n11325), .B1(n26902), .B2(
        data_in[7]), .ZN(n11332) );
  INV_X1 U15811 ( .A(n11333), .ZN(n24274) );
  AOI22_X1 U15812 ( .A1(\mem[229][0] ), .A2(n11334), .B1(n26901), .B2(
        data_in[0]), .ZN(n11333) );
  INV_X1 U15813 ( .A(n11335), .ZN(n24273) );
  AOI22_X1 U15814 ( .A1(\mem[229][1] ), .A2(n11334), .B1(n26901), .B2(
        data_in[1]), .ZN(n11335) );
  INV_X1 U15815 ( .A(n11336), .ZN(n24272) );
  AOI22_X1 U15816 ( .A1(\mem[229][2] ), .A2(n11334), .B1(n26901), .B2(
        data_in[2]), .ZN(n11336) );
  INV_X1 U15817 ( .A(n11337), .ZN(n24271) );
  AOI22_X1 U15818 ( .A1(\mem[229][3] ), .A2(n11334), .B1(n26901), .B2(
        data_in[3]), .ZN(n11337) );
  INV_X1 U15819 ( .A(n11338), .ZN(n24270) );
  AOI22_X1 U15820 ( .A1(\mem[229][4] ), .A2(n11334), .B1(n26901), .B2(
        data_in[4]), .ZN(n11338) );
  INV_X1 U15821 ( .A(n11339), .ZN(n24269) );
  AOI22_X1 U15822 ( .A1(\mem[229][5] ), .A2(n11334), .B1(n26901), .B2(
        data_in[5]), .ZN(n11339) );
  INV_X1 U15823 ( .A(n11340), .ZN(n24268) );
  AOI22_X1 U15824 ( .A1(\mem[229][6] ), .A2(n11334), .B1(n26901), .B2(
        data_in[6]), .ZN(n11340) );
  INV_X1 U15825 ( .A(n11341), .ZN(n24267) );
  AOI22_X1 U15826 ( .A1(\mem[229][7] ), .A2(n11334), .B1(n26901), .B2(
        data_in[7]), .ZN(n11341) );
  INV_X1 U15827 ( .A(n11342), .ZN(n24266) );
  AOI22_X1 U15828 ( .A1(\mem[230][0] ), .A2(n11343), .B1(n26900), .B2(
        data_in[0]), .ZN(n11342) );
  INV_X1 U15829 ( .A(n11344), .ZN(n24265) );
  AOI22_X1 U15830 ( .A1(\mem[230][1] ), .A2(n11343), .B1(n26900), .B2(
        data_in[1]), .ZN(n11344) );
  INV_X1 U15831 ( .A(n11345), .ZN(n24264) );
  AOI22_X1 U15832 ( .A1(\mem[230][2] ), .A2(n11343), .B1(n26900), .B2(
        data_in[2]), .ZN(n11345) );
  INV_X1 U15833 ( .A(n11346), .ZN(n24263) );
  AOI22_X1 U15834 ( .A1(\mem[230][3] ), .A2(n11343), .B1(n26900), .B2(
        data_in[3]), .ZN(n11346) );
  INV_X1 U15835 ( .A(n11347), .ZN(n24262) );
  AOI22_X1 U15836 ( .A1(\mem[230][4] ), .A2(n11343), .B1(n26900), .B2(
        data_in[4]), .ZN(n11347) );
  INV_X1 U15837 ( .A(n11348), .ZN(n24261) );
  AOI22_X1 U15838 ( .A1(\mem[230][5] ), .A2(n11343), .B1(n26900), .B2(
        data_in[5]), .ZN(n11348) );
  INV_X1 U15839 ( .A(n11349), .ZN(n24260) );
  AOI22_X1 U15840 ( .A1(\mem[230][6] ), .A2(n11343), .B1(n26900), .B2(
        data_in[6]), .ZN(n11349) );
  INV_X1 U15841 ( .A(n11350), .ZN(n24259) );
  AOI22_X1 U15842 ( .A1(\mem[230][7] ), .A2(n11343), .B1(n26900), .B2(
        data_in[7]), .ZN(n11350) );
  INV_X1 U15843 ( .A(n11351), .ZN(n24258) );
  AOI22_X1 U15844 ( .A1(\mem[231][0] ), .A2(n11352), .B1(n26899), .B2(
        data_in[0]), .ZN(n11351) );
  INV_X1 U15845 ( .A(n11353), .ZN(n24257) );
  AOI22_X1 U15846 ( .A1(\mem[231][1] ), .A2(n11352), .B1(n26899), .B2(
        data_in[1]), .ZN(n11353) );
  INV_X1 U15847 ( .A(n11354), .ZN(n24256) );
  AOI22_X1 U15848 ( .A1(\mem[231][2] ), .A2(n11352), .B1(n26899), .B2(
        data_in[2]), .ZN(n11354) );
  INV_X1 U15849 ( .A(n11355), .ZN(n24255) );
  AOI22_X1 U15850 ( .A1(\mem[231][3] ), .A2(n11352), .B1(n26899), .B2(
        data_in[3]), .ZN(n11355) );
  INV_X1 U15851 ( .A(n11356), .ZN(n24254) );
  AOI22_X1 U15852 ( .A1(\mem[231][4] ), .A2(n11352), .B1(n26899), .B2(
        data_in[4]), .ZN(n11356) );
  INV_X1 U15853 ( .A(n11357), .ZN(n24253) );
  AOI22_X1 U15854 ( .A1(\mem[231][5] ), .A2(n11352), .B1(n26899), .B2(
        data_in[5]), .ZN(n11357) );
  INV_X1 U15855 ( .A(n11358), .ZN(n24252) );
  AOI22_X1 U15856 ( .A1(\mem[231][6] ), .A2(n11352), .B1(n26899), .B2(
        data_in[6]), .ZN(n11358) );
  INV_X1 U15857 ( .A(n11359), .ZN(n24251) );
  AOI22_X1 U15858 ( .A1(\mem[231][7] ), .A2(n11352), .B1(n26899), .B2(
        data_in[7]), .ZN(n11359) );
  INV_X1 U15859 ( .A(n11577), .ZN(n24058) );
  AOI22_X1 U15860 ( .A1(\mem[256][0] ), .A2(n11578), .B1(n26874), .B2(
        data_in[0]), .ZN(n11577) );
  INV_X1 U15861 ( .A(n11579), .ZN(n24057) );
  AOI22_X1 U15862 ( .A1(\mem[256][1] ), .A2(n11578), .B1(n26874), .B2(
        data_in[1]), .ZN(n11579) );
  INV_X1 U15863 ( .A(n11580), .ZN(n24056) );
  AOI22_X1 U15864 ( .A1(\mem[256][2] ), .A2(n11578), .B1(n26874), .B2(
        data_in[2]), .ZN(n11580) );
  INV_X1 U15865 ( .A(n11581), .ZN(n24055) );
  AOI22_X1 U15866 ( .A1(\mem[256][3] ), .A2(n11578), .B1(n26874), .B2(
        data_in[3]), .ZN(n11581) );
  INV_X1 U15867 ( .A(n11582), .ZN(n24054) );
  AOI22_X1 U15868 ( .A1(\mem[256][4] ), .A2(n11578), .B1(n26874), .B2(
        data_in[4]), .ZN(n11582) );
  INV_X1 U15869 ( .A(n11583), .ZN(n24053) );
  AOI22_X1 U15870 ( .A1(\mem[256][5] ), .A2(n11578), .B1(n26874), .B2(
        data_in[5]), .ZN(n11583) );
  INV_X1 U15871 ( .A(n11584), .ZN(n24052) );
  AOI22_X1 U15872 ( .A1(\mem[256][6] ), .A2(n11578), .B1(n26874), .B2(
        data_in[6]), .ZN(n11584) );
  INV_X1 U15873 ( .A(n11585), .ZN(n24051) );
  AOI22_X1 U15874 ( .A1(\mem[256][7] ), .A2(n11578), .B1(n26874), .B2(
        data_in[7]), .ZN(n11585) );
  INV_X1 U15875 ( .A(n11587), .ZN(n24050) );
  AOI22_X1 U15876 ( .A1(\mem[257][0] ), .A2(n11588), .B1(n26873), .B2(
        data_in[0]), .ZN(n11587) );
  INV_X1 U15877 ( .A(n11589), .ZN(n24049) );
  AOI22_X1 U15878 ( .A1(\mem[257][1] ), .A2(n11588), .B1(n26873), .B2(
        data_in[1]), .ZN(n11589) );
  INV_X1 U15879 ( .A(n11590), .ZN(n24048) );
  AOI22_X1 U15880 ( .A1(\mem[257][2] ), .A2(n11588), .B1(n26873), .B2(
        data_in[2]), .ZN(n11590) );
  INV_X1 U15881 ( .A(n11591), .ZN(n24047) );
  AOI22_X1 U15882 ( .A1(\mem[257][3] ), .A2(n11588), .B1(n26873), .B2(
        data_in[3]), .ZN(n11591) );
  INV_X1 U15883 ( .A(n11592), .ZN(n24046) );
  AOI22_X1 U15884 ( .A1(\mem[257][4] ), .A2(n11588), .B1(n26873), .B2(
        data_in[4]), .ZN(n11592) );
  INV_X1 U15885 ( .A(n11593), .ZN(n24045) );
  AOI22_X1 U15886 ( .A1(\mem[257][5] ), .A2(n11588), .B1(n26873), .B2(
        data_in[5]), .ZN(n11593) );
  INV_X1 U15887 ( .A(n11594), .ZN(n24044) );
  AOI22_X1 U15888 ( .A1(\mem[257][6] ), .A2(n11588), .B1(n26873), .B2(
        data_in[6]), .ZN(n11594) );
  INV_X1 U15889 ( .A(n11595), .ZN(n24043) );
  AOI22_X1 U15890 ( .A1(\mem[257][7] ), .A2(n11588), .B1(n26873), .B2(
        data_in[7]), .ZN(n11595) );
  INV_X1 U15891 ( .A(n11596), .ZN(n24042) );
  AOI22_X1 U15892 ( .A1(\mem[258][0] ), .A2(n11597), .B1(n26872), .B2(
        data_in[0]), .ZN(n11596) );
  INV_X1 U15893 ( .A(n11598), .ZN(n24041) );
  AOI22_X1 U15894 ( .A1(\mem[258][1] ), .A2(n11597), .B1(n26872), .B2(
        data_in[1]), .ZN(n11598) );
  INV_X1 U15895 ( .A(n11599), .ZN(n24040) );
  AOI22_X1 U15896 ( .A1(\mem[258][2] ), .A2(n11597), .B1(n26872), .B2(
        data_in[2]), .ZN(n11599) );
  INV_X1 U15897 ( .A(n11600), .ZN(n24039) );
  AOI22_X1 U15898 ( .A1(\mem[258][3] ), .A2(n11597), .B1(n26872), .B2(
        data_in[3]), .ZN(n11600) );
  INV_X1 U15899 ( .A(n11601), .ZN(n24038) );
  AOI22_X1 U15900 ( .A1(\mem[258][4] ), .A2(n11597), .B1(n26872), .B2(
        data_in[4]), .ZN(n11601) );
  INV_X1 U15901 ( .A(n11602), .ZN(n24037) );
  AOI22_X1 U15902 ( .A1(\mem[258][5] ), .A2(n11597), .B1(n26872), .B2(
        data_in[5]), .ZN(n11602) );
  INV_X1 U15903 ( .A(n11603), .ZN(n24036) );
  AOI22_X1 U15904 ( .A1(\mem[258][6] ), .A2(n11597), .B1(n26872), .B2(
        data_in[6]), .ZN(n11603) );
  INV_X1 U15905 ( .A(n11604), .ZN(n24035) );
  AOI22_X1 U15906 ( .A1(\mem[258][7] ), .A2(n11597), .B1(n26872), .B2(
        data_in[7]), .ZN(n11604) );
  INV_X1 U15907 ( .A(n11605), .ZN(n24034) );
  AOI22_X1 U15908 ( .A1(\mem[259][0] ), .A2(n11606), .B1(n26871), .B2(
        data_in[0]), .ZN(n11605) );
  INV_X1 U15909 ( .A(n11607), .ZN(n24033) );
  AOI22_X1 U15910 ( .A1(\mem[259][1] ), .A2(n11606), .B1(n26871), .B2(
        data_in[1]), .ZN(n11607) );
  INV_X1 U15911 ( .A(n11608), .ZN(n24032) );
  AOI22_X1 U15912 ( .A1(\mem[259][2] ), .A2(n11606), .B1(n26871), .B2(
        data_in[2]), .ZN(n11608) );
  INV_X1 U15913 ( .A(n11609), .ZN(n24031) );
  AOI22_X1 U15914 ( .A1(\mem[259][3] ), .A2(n11606), .B1(n26871), .B2(
        data_in[3]), .ZN(n11609) );
  INV_X1 U15915 ( .A(n11610), .ZN(n24030) );
  AOI22_X1 U15916 ( .A1(\mem[259][4] ), .A2(n11606), .B1(n26871), .B2(
        data_in[4]), .ZN(n11610) );
  INV_X1 U15917 ( .A(n11611), .ZN(n24029) );
  AOI22_X1 U15918 ( .A1(\mem[259][5] ), .A2(n11606), .B1(n26871), .B2(
        data_in[5]), .ZN(n11611) );
  INV_X1 U15919 ( .A(n11612), .ZN(n24028) );
  AOI22_X1 U15920 ( .A1(\mem[259][6] ), .A2(n11606), .B1(n26871), .B2(
        data_in[6]), .ZN(n11612) );
  INV_X1 U15921 ( .A(n11613), .ZN(n24027) );
  AOI22_X1 U15922 ( .A1(\mem[259][7] ), .A2(n11606), .B1(n26871), .B2(
        data_in[7]), .ZN(n11613) );
  INV_X1 U15923 ( .A(n11614), .ZN(n24026) );
  AOI22_X1 U15924 ( .A1(\mem[260][0] ), .A2(n11615), .B1(n26870), .B2(
        data_in[0]), .ZN(n11614) );
  INV_X1 U15925 ( .A(n11616), .ZN(n24025) );
  AOI22_X1 U15926 ( .A1(\mem[260][1] ), .A2(n11615), .B1(n26870), .B2(
        data_in[1]), .ZN(n11616) );
  INV_X1 U15927 ( .A(n11617), .ZN(n24024) );
  AOI22_X1 U15928 ( .A1(\mem[260][2] ), .A2(n11615), .B1(n26870), .B2(
        data_in[2]), .ZN(n11617) );
  INV_X1 U15929 ( .A(n11618), .ZN(n24023) );
  AOI22_X1 U15930 ( .A1(\mem[260][3] ), .A2(n11615), .B1(n26870), .B2(
        data_in[3]), .ZN(n11618) );
  INV_X1 U15931 ( .A(n11619), .ZN(n24022) );
  AOI22_X1 U15932 ( .A1(\mem[260][4] ), .A2(n11615), .B1(n26870), .B2(
        data_in[4]), .ZN(n11619) );
  INV_X1 U15933 ( .A(n11620), .ZN(n24021) );
  AOI22_X1 U15934 ( .A1(\mem[260][5] ), .A2(n11615), .B1(n26870), .B2(
        data_in[5]), .ZN(n11620) );
  INV_X1 U15935 ( .A(n11621), .ZN(n24020) );
  AOI22_X1 U15936 ( .A1(\mem[260][6] ), .A2(n11615), .B1(n26870), .B2(
        data_in[6]), .ZN(n11621) );
  INV_X1 U15937 ( .A(n11622), .ZN(n24019) );
  AOI22_X1 U15938 ( .A1(\mem[260][7] ), .A2(n11615), .B1(n26870), .B2(
        data_in[7]), .ZN(n11622) );
  INV_X1 U15939 ( .A(n11623), .ZN(n24018) );
  AOI22_X1 U15940 ( .A1(\mem[261][0] ), .A2(n11624), .B1(n26869), .B2(
        data_in[0]), .ZN(n11623) );
  INV_X1 U15941 ( .A(n11625), .ZN(n24017) );
  AOI22_X1 U15942 ( .A1(\mem[261][1] ), .A2(n11624), .B1(n26869), .B2(
        data_in[1]), .ZN(n11625) );
  INV_X1 U15943 ( .A(n11626), .ZN(n24016) );
  AOI22_X1 U15944 ( .A1(\mem[261][2] ), .A2(n11624), .B1(n26869), .B2(
        data_in[2]), .ZN(n11626) );
  INV_X1 U15945 ( .A(n11627), .ZN(n24015) );
  AOI22_X1 U15946 ( .A1(\mem[261][3] ), .A2(n11624), .B1(n26869), .B2(
        data_in[3]), .ZN(n11627) );
  INV_X1 U15947 ( .A(n11628), .ZN(n24014) );
  AOI22_X1 U15948 ( .A1(\mem[261][4] ), .A2(n11624), .B1(n26869), .B2(
        data_in[4]), .ZN(n11628) );
  INV_X1 U15949 ( .A(n11629), .ZN(n24013) );
  AOI22_X1 U15950 ( .A1(\mem[261][5] ), .A2(n11624), .B1(n26869), .B2(
        data_in[5]), .ZN(n11629) );
  INV_X1 U15951 ( .A(n11630), .ZN(n24012) );
  AOI22_X1 U15952 ( .A1(\mem[261][6] ), .A2(n11624), .B1(n26869), .B2(
        data_in[6]), .ZN(n11630) );
  INV_X1 U15953 ( .A(n11631), .ZN(n24011) );
  AOI22_X1 U15954 ( .A1(\mem[261][7] ), .A2(n11624), .B1(n26869), .B2(
        data_in[7]), .ZN(n11631) );
  INV_X1 U15955 ( .A(n11632), .ZN(n24010) );
  AOI22_X1 U15956 ( .A1(\mem[262][0] ), .A2(n11633), .B1(n26868), .B2(
        data_in[0]), .ZN(n11632) );
  INV_X1 U15957 ( .A(n11634), .ZN(n24009) );
  AOI22_X1 U15958 ( .A1(\mem[262][1] ), .A2(n11633), .B1(n26868), .B2(
        data_in[1]), .ZN(n11634) );
  INV_X1 U15959 ( .A(n11635), .ZN(n24008) );
  AOI22_X1 U15960 ( .A1(\mem[262][2] ), .A2(n11633), .B1(n26868), .B2(
        data_in[2]), .ZN(n11635) );
  INV_X1 U15961 ( .A(n11636), .ZN(n24007) );
  AOI22_X1 U15962 ( .A1(\mem[262][3] ), .A2(n11633), .B1(n26868), .B2(
        data_in[3]), .ZN(n11636) );
  INV_X1 U15963 ( .A(n11637), .ZN(n24006) );
  AOI22_X1 U15964 ( .A1(\mem[262][4] ), .A2(n11633), .B1(n26868), .B2(
        data_in[4]), .ZN(n11637) );
  INV_X1 U15965 ( .A(n11638), .ZN(n24005) );
  AOI22_X1 U15966 ( .A1(\mem[262][5] ), .A2(n11633), .B1(n26868), .B2(
        data_in[5]), .ZN(n11638) );
  INV_X1 U15967 ( .A(n11639), .ZN(n24004) );
  AOI22_X1 U15968 ( .A1(\mem[262][6] ), .A2(n11633), .B1(n26868), .B2(
        data_in[6]), .ZN(n11639) );
  INV_X1 U15969 ( .A(n11640), .ZN(n24003) );
  AOI22_X1 U15970 ( .A1(\mem[262][7] ), .A2(n11633), .B1(n26868), .B2(
        data_in[7]), .ZN(n11640) );
  INV_X1 U15971 ( .A(n11641), .ZN(n24002) );
  AOI22_X1 U15972 ( .A1(\mem[263][0] ), .A2(n11642), .B1(n26867), .B2(
        data_in[0]), .ZN(n11641) );
  INV_X1 U15973 ( .A(n11643), .ZN(n24001) );
  AOI22_X1 U15974 ( .A1(\mem[263][1] ), .A2(n11642), .B1(n26867), .B2(
        data_in[1]), .ZN(n11643) );
  INV_X1 U15975 ( .A(n11644), .ZN(n24000) );
  AOI22_X1 U15976 ( .A1(\mem[263][2] ), .A2(n11642), .B1(n26867), .B2(
        data_in[2]), .ZN(n11644) );
  INV_X1 U15977 ( .A(n11645), .ZN(n23999) );
  AOI22_X1 U15978 ( .A1(\mem[263][3] ), .A2(n11642), .B1(n26867), .B2(
        data_in[3]), .ZN(n11645) );
  INV_X1 U15979 ( .A(n11646), .ZN(n23998) );
  AOI22_X1 U15980 ( .A1(\mem[263][4] ), .A2(n11642), .B1(n26867), .B2(
        data_in[4]), .ZN(n11646) );
  INV_X1 U15981 ( .A(n11647), .ZN(n23997) );
  AOI22_X1 U15982 ( .A1(\mem[263][5] ), .A2(n11642), .B1(n26867), .B2(
        data_in[5]), .ZN(n11647) );
  INV_X1 U15983 ( .A(n11648), .ZN(n23996) );
  AOI22_X1 U15984 ( .A1(\mem[263][6] ), .A2(n11642), .B1(n26867), .B2(
        data_in[6]), .ZN(n11648) );
  INV_X1 U15985 ( .A(n11649), .ZN(n23995) );
  AOI22_X1 U15986 ( .A1(\mem[263][7] ), .A2(n11642), .B1(n26867), .B2(
        data_in[7]), .ZN(n11649) );
  INV_X1 U15987 ( .A(n11867), .ZN(n23802) );
  AOI22_X1 U15988 ( .A1(\mem[288][0] ), .A2(n11868), .B1(n26842), .B2(
        data_in[0]), .ZN(n11867) );
  INV_X1 U15989 ( .A(n11869), .ZN(n23801) );
  AOI22_X1 U15990 ( .A1(\mem[288][1] ), .A2(n11868), .B1(n26842), .B2(
        data_in[1]), .ZN(n11869) );
  INV_X1 U15991 ( .A(n11870), .ZN(n23800) );
  AOI22_X1 U15992 ( .A1(\mem[288][2] ), .A2(n11868), .B1(n26842), .B2(
        data_in[2]), .ZN(n11870) );
  INV_X1 U15993 ( .A(n11871), .ZN(n23799) );
  AOI22_X1 U15994 ( .A1(\mem[288][3] ), .A2(n11868), .B1(n26842), .B2(
        data_in[3]), .ZN(n11871) );
  INV_X1 U15995 ( .A(n11872), .ZN(n23798) );
  AOI22_X1 U15996 ( .A1(\mem[288][4] ), .A2(n11868), .B1(n26842), .B2(
        data_in[4]), .ZN(n11872) );
  INV_X1 U15997 ( .A(n11873), .ZN(n23797) );
  AOI22_X1 U15998 ( .A1(\mem[288][5] ), .A2(n11868), .B1(n26842), .B2(
        data_in[5]), .ZN(n11873) );
  INV_X1 U15999 ( .A(n11874), .ZN(n23796) );
  AOI22_X1 U16000 ( .A1(\mem[288][6] ), .A2(n11868), .B1(n26842), .B2(
        data_in[6]), .ZN(n11874) );
  INV_X1 U16001 ( .A(n11875), .ZN(n23795) );
  AOI22_X1 U16002 ( .A1(\mem[288][7] ), .A2(n11868), .B1(n26842), .B2(
        data_in[7]), .ZN(n11875) );
  INV_X1 U16003 ( .A(n11877), .ZN(n23794) );
  AOI22_X1 U16004 ( .A1(\mem[289][0] ), .A2(n11878), .B1(n26841), .B2(
        data_in[0]), .ZN(n11877) );
  INV_X1 U16005 ( .A(n11879), .ZN(n23793) );
  AOI22_X1 U16006 ( .A1(\mem[289][1] ), .A2(n11878), .B1(n26841), .B2(
        data_in[1]), .ZN(n11879) );
  INV_X1 U16007 ( .A(n11880), .ZN(n23792) );
  AOI22_X1 U16008 ( .A1(\mem[289][2] ), .A2(n11878), .B1(n26841), .B2(
        data_in[2]), .ZN(n11880) );
  INV_X1 U16009 ( .A(n11881), .ZN(n23791) );
  AOI22_X1 U16010 ( .A1(\mem[289][3] ), .A2(n11878), .B1(n26841), .B2(
        data_in[3]), .ZN(n11881) );
  INV_X1 U16011 ( .A(n11882), .ZN(n23790) );
  AOI22_X1 U16012 ( .A1(\mem[289][4] ), .A2(n11878), .B1(n26841), .B2(
        data_in[4]), .ZN(n11882) );
  INV_X1 U16013 ( .A(n11883), .ZN(n23789) );
  AOI22_X1 U16014 ( .A1(\mem[289][5] ), .A2(n11878), .B1(n26841), .B2(
        data_in[5]), .ZN(n11883) );
  INV_X1 U16015 ( .A(n11884), .ZN(n23788) );
  AOI22_X1 U16016 ( .A1(\mem[289][6] ), .A2(n11878), .B1(n26841), .B2(
        data_in[6]), .ZN(n11884) );
  INV_X1 U16017 ( .A(n11885), .ZN(n23787) );
  AOI22_X1 U16018 ( .A1(\mem[289][7] ), .A2(n11878), .B1(n26841), .B2(
        data_in[7]), .ZN(n11885) );
  INV_X1 U16019 ( .A(n11886), .ZN(n23786) );
  AOI22_X1 U16020 ( .A1(\mem[290][0] ), .A2(n11887), .B1(n26840), .B2(
        data_in[0]), .ZN(n11886) );
  INV_X1 U16021 ( .A(n11888), .ZN(n23785) );
  AOI22_X1 U16022 ( .A1(\mem[290][1] ), .A2(n11887), .B1(n26840), .B2(
        data_in[1]), .ZN(n11888) );
  INV_X1 U16023 ( .A(n11889), .ZN(n23784) );
  AOI22_X1 U16024 ( .A1(\mem[290][2] ), .A2(n11887), .B1(n26840), .B2(
        data_in[2]), .ZN(n11889) );
  INV_X1 U16025 ( .A(n11890), .ZN(n23783) );
  AOI22_X1 U16026 ( .A1(\mem[290][3] ), .A2(n11887), .B1(n26840), .B2(
        data_in[3]), .ZN(n11890) );
  INV_X1 U16027 ( .A(n11891), .ZN(n23782) );
  AOI22_X1 U16028 ( .A1(\mem[290][4] ), .A2(n11887), .B1(n26840), .B2(
        data_in[4]), .ZN(n11891) );
  INV_X1 U16029 ( .A(n11892), .ZN(n23781) );
  AOI22_X1 U16030 ( .A1(\mem[290][5] ), .A2(n11887), .B1(n26840), .B2(
        data_in[5]), .ZN(n11892) );
  INV_X1 U16031 ( .A(n11893), .ZN(n23780) );
  AOI22_X1 U16032 ( .A1(\mem[290][6] ), .A2(n11887), .B1(n26840), .B2(
        data_in[6]), .ZN(n11893) );
  INV_X1 U16033 ( .A(n11894), .ZN(n23779) );
  AOI22_X1 U16034 ( .A1(\mem[290][7] ), .A2(n11887), .B1(n26840), .B2(
        data_in[7]), .ZN(n11894) );
  INV_X1 U16035 ( .A(n11895), .ZN(n23778) );
  AOI22_X1 U16036 ( .A1(\mem[291][0] ), .A2(n11896), .B1(n26839), .B2(
        data_in[0]), .ZN(n11895) );
  INV_X1 U16037 ( .A(n11897), .ZN(n23777) );
  AOI22_X1 U16038 ( .A1(\mem[291][1] ), .A2(n11896), .B1(n26839), .B2(
        data_in[1]), .ZN(n11897) );
  INV_X1 U16039 ( .A(n11898), .ZN(n23776) );
  AOI22_X1 U16040 ( .A1(\mem[291][2] ), .A2(n11896), .B1(n26839), .B2(
        data_in[2]), .ZN(n11898) );
  INV_X1 U16041 ( .A(n11899), .ZN(n23775) );
  AOI22_X1 U16042 ( .A1(\mem[291][3] ), .A2(n11896), .B1(n26839), .B2(
        data_in[3]), .ZN(n11899) );
  INV_X1 U16043 ( .A(n11900), .ZN(n23774) );
  AOI22_X1 U16044 ( .A1(\mem[291][4] ), .A2(n11896), .B1(n26839), .B2(
        data_in[4]), .ZN(n11900) );
  INV_X1 U16045 ( .A(n11901), .ZN(n23773) );
  AOI22_X1 U16046 ( .A1(\mem[291][5] ), .A2(n11896), .B1(n26839), .B2(
        data_in[5]), .ZN(n11901) );
  INV_X1 U16047 ( .A(n11902), .ZN(n23772) );
  AOI22_X1 U16048 ( .A1(\mem[291][6] ), .A2(n11896), .B1(n26839), .B2(
        data_in[6]), .ZN(n11902) );
  INV_X1 U16049 ( .A(n11903), .ZN(n23771) );
  AOI22_X1 U16050 ( .A1(\mem[291][7] ), .A2(n11896), .B1(n26839), .B2(
        data_in[7]), .ZN(n11903) );
  INV_X1 U16051 ( .A(n11904), .ZN(n23770) );
  AOI22_X1 U16052 ( .A1(\mem[292][0] ), .A2(n11905), .B1(n26838), .B2(
        data_in[0]), .ZN(n11904) );
  INV_X1 U16053 ( .A(n11906), .ZN(n23769) );
  AOI22_X1 U16054 ( .A1(\mem[292][1] ), .A2(n11905), .B1(n26838), .B2(
        data_in[1]), .ZN(n11906) );
  INV_X1 U16055 ( .A(n11907), .ZN(n23768) );
  AOI22_X1 U16056 ( .A1(\mem[292][2] ), .A2(n11905), .B1(n26838), .B2(
        data_in[2]), .ZN(n11907) );
  INV_X1 U16057 ( .A(n11908), .ZN(n23767) );
  AOI22_X1 U16058 ( .A1(\mem[292][3] ), .A2(n11905), .B1(n26838), .B2(
        data_in[3]), .ZN(n11908) );
  INV_X1 U16059 ( .A(n11909), .ZN(n23766) );
  AOI22_X1 U16060 ( .A1(\mem[292][4] ), .A2(n11905), .B1(n26838), .B2(
        data_in[4]), .ZN(n11909) );
  INV_X1 U16061 ( .A(n11910), .ZN(n23765) );
  AOI22_X1 U16062 ( .A1(\mem[292][5] ), .A2(n11905), .B1(n26838), .B2(
        data_in[5]), .ZN(n11910) );
  INV_X1 U16063 ( .A(n11911), .ZN(n23764) );
  AOI22_X1 U16064 ( .A1(\mem[292][6] ), .A2(n11905), .B1(n26838), .B2(
        data_in[6]), .ZN(n11911) );
  INV_X1 U16065 ( .A(n11912), .ZN(n23763) );
  AOI22_X1 U16066 ( .A1(\mem[292][7] ), .A2(n11905), .B1(n26838), .B2(
        data_in[7]), .ZN(n11912) );
  INV_X1 U16067 ( .A(n11913), .ZN(n23762) );
  AOI22_X1 U16068 ( .A1(\mem[293][0] ), .A2(n11914), .B1(n26837), .B2(
        data_in[0]), .ZN(n11913) );
  INV_X1 U16069 ( .A(n11915), .ZN(n23761) );
  AOI22_X1 U16070 ( .A1(\mem[293][1] ), .A2(n11914), .B1(n26837), .B2(
        data_in[1]), .ZN(n11915) );
  INV_X1 U16071 ( .A(n11916), .ZN(n23760) );
  AOI22_X1 U16072 ( .A1(\mem[293][2] ), .A2(n11914), .B1(n26837), .B2(
        data_in[2]), .ZN(n11916) );
  INV_X1 U16073 ( .A(n11917), .ZN(n23759) );
  AOI22_X1 U16074 ( .A1(\mem[293][3] ), .A2(n11914), .B1(n26837), .B2(
        data_in[3]), .ZN(n11917) );
  INV_X1 U16075 ( .A(n11918), .ZN(n23758) );
  AOI22_X1 U16076 ( .A1(\mem[293][4] ), .A2(n11914), .B1(n26837), .B2(
        data_in[4]), .ZN(n11918) );
  INV_X1 U16077 ( .A(n11919), .ZN(n23757) );
  AOI22_X1 U16078 ( .A1(\mem[293][5] ), .A2(n11914), .B1(n26837), .B2(
        data_in[5]), .ZN(n11919) );
  INV_X1 U16079 ( .A(n11920), .ZN(n23756) );
  AOI22_X1 U16080 ( .A1(\mem[293][6] ), .A2(n11914), .B1(n26837), .B2(
        data_in[6]), .ZN(n11920) );
  INV_X1 U16081 ( .A(n11921), .ZN(n23755) );
  AOI22_X1 U16082 ( .A1(\mem[293][7] ), .A2(n11914), .B1(n26837), .B2(
        data_in[7]), .ZN(n11921) );
  INV_X1 U16083 ( .A(n11922), .ZN(n23754) );
  AOI22_X1 U16084 ( .A1(\mem[294][0] ), .A2(n11923), .B1(n26836), .B2(
        data_in[0]), .ZN(n11922) );
  INV_X1 U16085 ( .A(n11924), .ZN(n23753) );
  AOI22_X1 U16086 ( .A1(\mem[294][1] ), .A2(n11923), .B1(n26836), .B2(
        data_in[1]), .ZN(n11924) );
  INV_X1 U16087 ( .A(n11925), .ZN(n23752) );
  AOI22_X1 U16088 ( .A1(\mem[294][2] ), .A2(n11923), .B1(n26836), .B2(
        data_in[2]), .ZN(n11925) );
  INV_X1 U16089 ( .A(n11926), .ZN(n23751) );
  AOI22_X1 U16090 ( .A1(\mem[294][3] ), .A2(n11923), .B1(n26836), .B2(
        data_in[3]), .ZN(n11926) );
  INV_X1 U16091 ( .A(n11927), .ZN(n23750) );
  AOI22_X1 U16092 ( .A1(\mem[294][4] ), .A2(n11923), .B1(n26836), .B2(
        data_in[4]), .ZN(n11927) );
  INV_X1 U16093 ( .A(n11928), .ZN(n23749) );
  AOI22_X1 U16094 ( .A1(\mem[294][5] ), .A2(n11923), .B1(n26836), .B2(
        data_in[5]), .ZN(n11928) );
  INV_X1 U16095 ( .A(n11929), .ZN(n23748) );
  AOI22_X1 U16096 ( .A1(\mem[294][6] ), .A2(n11923), .B1(n26836), .B2(
        data_in[6]), .ZN(n11929) );
  INV_X1 U16097 ( .A(n11930), .ZN(n23747) );
  AOI22_X1 U16098 ( .A1(\mem[294][7] ), .A2(n11923), .B1(n26836), .B2(
        data_in[7]), .ZN(n11930) );
  INV_X1 U16099 ( .A(n11931), .ZN(n23746) );
  AOI22_X1 U16100 ( .A1(\mem[295][0] ), .A2(n11932), .B1(n26835), .B2(
        data_in[0]), .ZN(n11931) );
  INV_X1 U16101 ( .A(n11933), .ZN(n23745) );
  AOI22_X1 U16102 ( .A1(\mem[295][1] ), .A2(n11932), .B1(n26835), .B2(
        data_in[1]), .ZN(n11933) );
  INV_X1 U16103 ( .A(n11934), .ZN(n23744) );
  AOI22_X1 U16104 ( .A1(\mem[295][2] ), .A2(n11932), .B1(n26835), .B2(
        data_in[2]), .ZN(n11934) );
  INV_X1 U16105 ( .A(n11935), .ZN(n23743) );
  AOI22_X1 U16106 ( .A1(\mem[295][3] ), .A2(n11932), .B1(n26835), .B2(
        data_in[3]), .ZN(n11935) );
  INV_X1 U16107 ( .A(n11936), .ZN(n23742) );
  AOI22_X1 U16108 ( .A1(\mem[295][4] ), .A2(n11932), .B1(n26835), .B2(
        data_in[4]), .ZN(n11936) );
  INV_X1 U16109 ( .A(n11937), .ZN(n23741) );
  AOI22_X1 U16110 ( .A1(\mem[295][5] ), .A2(n11932), .B1(n26835), .B2(
        data_in[5]), .ZN(n11937) );
  INV_X1 U16111 ( .A(n11938), .ZN(n23740) );
  AOI22_X1 U16112 ( .A1(\mem[295][6] ), .A2(n11932), .B1(n26835), .B2(
        data_in[6]), .ZN(n11938) );
  INV_X1 U16113 ( .A(n11939), .ZN(n23739) );
  AOI22_X1 U16114 ( .A1(\mem[295][7] ), .A2(n11932), .B1(n26835), .B2(
        data_in[7]), .ZN(n11939) );
  INV_X1 U16115 ( .A(n12156), .ZN(n23546) );
  AOI22_X1 U16116 ( .A1(\mem[320][0] ), .A2(n12157), .B1(n26810), .B2(
        data_in[0]), .ZN(n12156) );
  INV_X1 U16117 ( .A(n12158), .ZN(n23545) );
  AOI22_X1 U16118 ( .A1(\mem[320][1] ), .A2(n12157), .B1(n26810), .B2(
        data_in[1]), .ZN(n12158) );
  INV_X1 U16119 ( .A(n12159), .ZN(n23544) );
  AOI22_X1 U16120 ( .A1(\mem[320][2] ), .A2(n12157), .B1(n26810), .B2(
        data_in[2]), .ZN(n12159) );
  INV_X1 U16121 ( .A(n12160), .ZN(n23543) );
  AOI22_X1 U16122 ( .A1(\mem[320][3] ), .A2(n12157), .B1(n26810), .B2(
        data_in[3]), .ZN(n12160) );
  INV_X1 U16123 ( .A(n12161), .ZN(n23542) );
  AOI22_X1 U16124 ( .A1(\mem[320][4] ), .A2(n12157), .B1(n26810), .B2(
        data_in[4]), .ZN(n12161) );
  INV_X1 U16125 ( .A(n12162), .ZN(n23541) );
  AOI22_X1 U16126 ( .A1(\mem[320][5] ), .A2(n12157), .B1(n26810), .B2(
        data_in[5]), .ZN(n12162) );
  INV_X1 U16127 ( .A(n12163), .ZN(n23540) );
  AOI22_X1 U16128 ( .A1(\mem[320][6] ), .A2(n12157), .B1(n26810), .B2(
        data_in[6]), .ZN(n12163) );
  INV_X1 U16129 ( .A(n12164), .ZN(n23539) );
  AOI22_X1 U16130 ( .A1(\mem[320][7] ), .A2(n12157), .B1(n26810), .B2(
        data_in[7]), .ZN(n12164) );
  INV_X1 U16131 ( .A(n12166), .ZN(n23538) );
  AOI22_X1 U16132 ( .A1(\mem[321][0] ), .A2(n12167), .B1(n26809), .B2(
        data_in[0]), .ZN(n12166) );
  INV_X1 U16133 ( .A(n12168), .ZN(n23537) );
  AOI22_X1 U16134 ( .A1(\mem[321][1] ), .A2(n12167), .B1(n26809), .B2(
        data_in[1]), .ZN(n12168) );
  INV_X1 U16135 ( .A(n12169), .ZN(n23536) );
  AOI22_X1 U16136 ( .A1(\mem[321][2] ), .A2(n12167), .B1(n26809), .B2(
        data_in[2]), .ZN(n12169) );
  INV_X1 U16137 ( .A(n12170), .ZN(n23535) );
  AOI22_X1 U16138 ( .A1(\mem[321][3] ), .A2(n12167), .B1(n26809), .B2(
        data_in[3]), .ZN(n12170) );
  INV_X1 U16139 ( .A(n12171), .ZN(n23534) );
  AOI22_X1 U16140 ( .A1(\mem[321][4] ), .A2(n12167), .B1(n26809), .B2(
        data_in[4]), .ZN(n12171) );
  INV_X1 U16141 ( .A(n12172), .ZN(n23533) );
  AOI22_X1 U16142 ( .A1(\mem[321][5] ), .A2(n12167), .B1(n26809), .B2(
        data_in[5]), .ZN(n12172) );
  INV_X1 U16143 ( .A(n12173), .ZN(n23532) );
  AOI22_X1 U16144 ( .A1(\mem[321][6] ), .A2(n12167), .B1(n26809), .B2(
        data_in[6]), .ZN(n12173) );
  INV_X1 U16145 ( .A(n12174), .ZN(n23531) );
  AOI22_X1 U16146 ( .A1(\mem[321][7] ), .A2(n12167), .B1(n26809), .B2(
        data_in[7]), .ZN(n12174) );
  INV_X1 U16147 ( .A(n12175), .ZN(n23530) );
  AOI22_X1 U16148 ( .A1(\mem[322][0] ), .A2(n12176), .B1(n26808), .B2(
        data_in[0]), .ZN(n12175) );
  INV_X1 U16149 ( .A(n12177), .ZN(n23529) );
  AOI22_X1 U16150 ( .A1(\mem[322][1] ), .A2(n12176), .B1(n26808), .B2(
        data_in[1]), .ZN(n12177) );
  INV_X1 U16151 ( .A(n12178), .ZN(n23528) );
  AOI22_X1 U16152 ( .A1(\mem[322][2] ), .A2(n12176), .B1(n26808), .B2(
        data_in[2]), .ZN(n12178) );
  INV_X1 U16153 ( .A(n12179), .ZN(n23527) );
  AOI22_X1 U16154 ( .A1(\mem[322][3] ), .A2(n12176), .B1(n26808), .B2(
        data_in[3]), .ZN(n12179) );
  INV_X1 U16155 ( .A(n12180), .ZN(n23526) );
  AOI22_X1 U16156 ( .A1(\mem[322][4] ), .A2(n12176), .B1(n26808), .B2(
        data_in[4]), .ZN(n12180) );
  INV_X1 U16157 ( .A(n12181), .ZN(n23525) );
  AOI22_X1 U16158 ( .A1(\mem[322][5] ), .A2(n12176), .B1(n26808), .B2(
        data_in[5]), .ZN(n12181) );
  INV_X1 U16159 ( .A(n12182), .ZN(n23524) );
  AOI22_X1 U16160 ( .A1(\mem[322][6] ), .A2(n12176), .B1(n26808), .B2(
        data_in[6]), .ZN(n12182) );
  INV_X1 U16161 ( .A(n12183), .ZN(n23523) );
  AOI22_X1 U16162 ( .A1(\mem[322][7] ), .A2(n12176), .B1(n26808), .B2(
        data_in[7]), .ZN(n12183) );
  INV_X1 U16163 ( .A(n12184), .ZN(n23522) );
  AOI22_X1 U16164 ( .A1(\mem[323][0] ), .A2(n12185), .B1(n26807), .B2(
        data_in[0]), .ZN(n12184) );
  INV_X1 U16165 ( .A(n12186), .ZN(n23521) );
  AOI22_X1 U16166 ( .A1(\mem[323][1] ), .A2(n12185), .B1(n26807), .B2(
        data_in[1]), .ZN(n12186) );
  INV_X1 U16167 ( .A(n12187), .ZN(n23520) );
  AOI22_X1 U16168 ( .A1(\mem[323][2] ), .A2(n12185), .B1(n26807), .B2(
        data_in[2]), .ZN(n12187) );
  INV_X1 U16169 ( .A(n12188), .ZN(n23519) );
  AOI22_X1 U16170 ( .A1(\mem[323][3] ), .A2(n12185), .B1(n26807), .B2(
        data_in[3]), .ZN(n12188) );
  INV_X1 U16171 ( .A(n12189), .ZN(n23518) );
  AOI22_X1 U16172 ( .A1(\mem[323][4] ), .A2(n12185), .B1(n26807), .B2(
        data_in[4]), .ZN(n12189) );
  INV_X1 U16173 ( .A(n12190), .ZN(n23517) );
  AOI22_X1 U16174 ( .A1(\mem[323][5] ), .A2(n12185), .B1(n26807), .B2(
        data_in[5]), .ZN(n12190) );
  INV_X1 U16175 ( .A(n12191), .ZN(n23516) );
  AOI22_X1 U16176 ( .A1(\mem[323][6] ), .A2(n12185), .B1(n26807), .B2(
        data_in[6]), .ZN(n12191) );
  INV_X1 U16177 ( .A(n12192), .ZN(n23515) );
  AOI22_X1 U16178 ( .A1(\mem[323][7] ), .A2(n12185), .B1(n26807), .B2(
        data_in[7]), .ZN(n12192) );
  INV_X1 U16179 ( .A(n12193), .ZN(n23514) );
  AOI22_X1 U16180 ( .A1(\mem[324][0] ), .A2(n12194), .B1(n26806), .B2(
        data_in[0]), .ZN(n12193) );
  INV_X1 U16181 ( .A(n12195), .ZN(n23513) );
  AOI22_X1 U16182 ( .A1(\mem[324][1] ), .A2(n12194), .B1(n26806), .B2(
        data_in[1]), .ZN(n12195) );
  INV_X1 U16183 ( .A(n12196), .ZN(n23512) );
  AOI22_X1 U16184 ( .A1(\mem[324][2] ), .A2(n12194), .B1(n26806), .B2(
        data_in[2]), .ZN(n12196) );
  INV_X1 U16185 ( .A(n12197), .ZN(n23511) );
  AOI22_X1 U16186 ( .A1(\mem[324][3] ), .A2(n12194), .B1(n26806), .B2(
        data_in[3]), .ZN(n12197) );
  INV_X1 U16187 ( .A(n12198), .ZN(n23510) );
  AOI22_X1 U16188 ( .A1(\mem[324][4] ), .A2(n12194), .B1(n26806), .B2(
        data_in[4]), .ZN(n12198) );
  INV_X1 U16189 ( .A(n12199), .ZN(n23509) );
  AOI22_X1 U16190 ( .A1(\mem[324][5] ), .A2(n12194), .B1(n26806), .B2(
        data_in[5]), .ZN(n12199) );
  INV_X1 U16191 ( .A(n12200), .ZN(n23508) );
  AOI22_X1 U16192 ( .A1(\mem[324][6] ), .A2(n12194), .B1(n26806), .B2(
        data_in[6]), .ZN(n12200) );
  INV_X1 U16193 ( .A(n12201), .ZN(n23507) );
  AOI22_X1 U16194 ( .A1(\mem[324][7] ), .A2(n12194), .B1(n26806), .B2(
        data_in[7]), .ZN(n12201) );
  INV_X1 U16195 ( .A(n12202), .ZN(n23506) );
  AOI22_X1 U16196 ( .A1(\mem[325][0] ), .A2(n12203), .B1(n26805), .B2(
        data_in[0]), .ZN(n12202) );
  INV_X1 U16197 ( .A(n12204), .ZN(n23505) );
  AOI22_X1 U16198 ( .A1(\mem[325][1] ), .A2(n12203), .B1(n26805), .B2(
        data_in[1]), .ZN(n12204) );
  INV_X1 U16199 ( .A(n12205), .ZN(n23504) );
  AOI22_X1 U16200 ( .A1(\mem[325][2] ), .A2(n12203), .B1(n26805), .B2(
        data_in[2]), .ZN(n12205) );
  INV_X1 U16201 ( .A(n12206), .ZN(n23503) );
  AOI22_X1 U16202 ( .A1(\mem[325][3] ), .A2(n12203), .B1(n26805), .B2(
        data_in[3]), .ZN(n12206) );
  INV_X1 U16203 ( .A(n12207), .ZN(n23502) );
  AOI22_X1 U16204 ( .A1(\mem[325][4] ), .A2(n12203), .B1(n26805), .B2(
        data_in[4]), .ZN(n12207) );
  INV_X1 U16205 ( .A(n12208), .ZN(n23501) );
  AOI22_X1 U16206 ( .A1(\mem[325][5] ), .A2(n12203), .B1(n26805), .B2(
        data_in[5]), .ZN(n12208) );
  INV_X1 U16207 ( .A(n12209), .ZN(n23500) );
  AOI22_X1 U16208 ( .A1(\mem[325][6] ), .A2(n12203), .B1(n26805), .B2(
        data_in[6]), .ZN(n12209) );
  INV_X1 U16209 ( .A(n12210), .ZN(n23499) );
  AOI22_X1 U16210 ( .A1(\mem[325][7] ), .A2(n12203), .B1(n26805), .B2(
        data_in[7]), .ZN(n12210) );
  INV_X1 U16211 ( .A(n12211), .ZN(n23498) );
  AOI22_X1 U16212 ( .A1(\mem[326][0] ), .A2(n12212), .B1(n26804), .B2(
        data_in[0]), .ZN(n12211) );
  INV_X1 U16213 ( .A(n12213), .ZN(n23497) );
  AOI22_X1 U16214 ( .A1(\mem[326][1] ), .A2(n12212), .B1(n26804), .B2(
        data_in[1]), .ZN(n12213) );
  INV_X1 U16215 ( .A(n12214), .ZN(n23496) );
  AOI22_X1 U16216 ( .A1(\mem[326][2] ), .A2(n12212), .B1(n26804), .B2(
        data_in[2]), .ZN(n12214) );
  INV_X1 U16217 ( .A(n12215), .ZN(n23495) );
  AOI22_X1 U16218 ( .A1(\mem[326][3] ), .A2(n12212), .B1(n26804), .B2(
        data_in[3]), .ZN(n12215) );
  INV_X1 U16219 ( .A(n12216), .ZN(n23494) );
  AOI22_X1 U16220 ( .A1(\mem[326][4] ), .A2(n12212), .B1(n26804), .B2(
        data_in[4]), .ZN(n12216) );
  INV_X1 U16221 ( .A(n12217), .ZN(n23493) );
  AOI22_X1 U16222 ( .A1(\mem[326][5] ), .A2(n12212), .B1(n26804), .B2(
        data_in[5]), .ZN(n12217) );
  INV_X1 U16223 ( .A(n12218), .ZN(n23492) );
  AOI22_X1 U16224 ( .A1(\mem[326][6] ), .A2(n12212), .B1(n26804), .B2(
        data_in[6]), .ZN(n12218) );
  INV_X1 U16225 ( .A(n12219), .ZN(n23491) );
  AOI22_X1 U16226 ( .A1(\mem[326][7] ), .A2(n12212), .B1(n26804), .B2(
        data_in[7]), .ZN(n12219) );
  INV_X1 U16227 ( .A(n12220), .ZN(n23490) );
  AOI22_X1 U16228 ( .A1(\mem[327][0] ), .A2(n12221), .B1(n26803), .B2(
        data_in[0]), .ZN(n12220) );
  INV_X1 U16229 ( .A(n12222), .ZN(n23489) );
  AOI22_X1 U16230 ( .A1(\mem[327][1] ), .A2(n12221), .B1(n26803), .B2(
        data_in[1]), .ZN(n12222) );
  INV_X1 U16231 ( .A(n12223), .ZN(n23488) );
  AOI22_X1 U16232 ( .A1(\mem[327][2] ), .A2(n12221), .B1(n26803), .B2(
        data_in[2]), .ZN(n12223) );
  INV_X1 U16233 ( .A(n12224), .ZN(n23487) );
  AOI22_X1 U16234 ( .A1(\mem[327][3] ), .A2(n12221), .B1(n26803), .B2(
        data_in[3]), .ZN(n12224) );
  INV_X1 U16235 ( .A(n12225), .ZN(n23486) );
  AOI22_X1 U16236 ( .A1(\mem[327][4] ), .A2(n12221), .B1(n26803), .B2(
        data_in[4]), .ZN(n12225) );
  INV_X1 U16237 ( .A(n12226), .ZN(n23485) );
  AOI22_X1 U16238 ( .A1(\mem[327][5] ), .A2(n12221), .B1(n26803), .B2(
        data_in[5]), .ZN(n12226) );
  INV_X1 U16239 ( .A(n12227), .ZN(n23484) );
  AOI22_X1 U16240 ( .A1(\mem[327][6] ), .A2(n12221), .B1(n26803), .B2(
        data_in[6]), .ZN(n12227) );
  INV_X1 U16241 ( .A(n12228), .ZN(n23483) );
  AOI22_X1 U16242 ( .A1(\mem[327][7] ), .A2(n12221), .B1(n26803), .B2(
        data_in[7]), .ZN(n12228) );
  INV_X1 U16243 ( .A(n12445), .ZN(n23290) );
  AOI22_X1 U16244 ( .A1(\mem[352][0] ), .A2(n12446), .B1(n26778), .B2(
        data_in[0]), .ZN(n12445) );
  INV_X1 U16245 ( .A(n12447), .ZN(n23289) );
  AOI22_X1 U16246 ( .A1(\mem[352][1] ), .A2(n12446), .B1(n26778), .B2(
        data_in[1]), .ZN(n12447) );
  INV_X1 U16247 ( .A(n12448), .ZN(n23288) );
  AOI22_X1 U16248 ( .A1(\mem[352][2] ), .A2(n12446), .B1(n26778), .B2(
        data_in[2]), .ZN(n12448) );
  INV_X1 U16249 ( .A(n12449), .ZN(n23287) );
  AOI22_X1 U16250 ( .A1(\mem[352][3] ), .A2(n12446), .B1(n26778), .B2(
        data_in[3]), .ZN(n12449) );
  INV_X1 U16251 ( .A(n12450), .ZN(n23286) );
  AOI22_X1 U16252 ( .A1(\mem[352][4] ), .A2(n12446), .B1(n26778), .B2(
        data_in[4]), .ZN(n12450) );
  INV_X1 U16253 ( .A(n12451), .ZN(n23285) );
  AOI22_X1 U16254 ( .A1(\mem[352][5] ), .A2(n12446), .B1(n26778), .B2(
        data_in[5]), .ZN(n12451) );
  INV_X1 U16255 ( .A(n12452), .ZN(n23284) );
  AOI22_X1 U16256 ( .A1(\mem[352][6] ), .A2(n12446), .B1(n26778), .B2(
        data_in[6]), .ZN(n12452) );
  INV_X1 U16257 ( .A(n12453), .ZN(n23283) );
  AOI22_X1 U16258 ( .A1(\mem[352][7] ), .A2(n12446), .B1(n26778), .B2(
        data_in[7]), .ZN(n12453) );
  INV_X1 U16259 ( .A(n12455), .ZN(n23282) );
  AOI22_X1 U16260 ( .A1(\mem[353][0] ), .A2(n12456), .B1(n26777), .B2(
        data_in[0]), .ZN(n12455) );
  INV_X1 U16261 ( .A(n12457), .ZN(n23281) );
  AOI22_X1 U16262 ( .A1(\mem[353][1] ), .A2(n12456), .B1(n26777), .B2(
        data_in[1]), .ZN(n12457) );
  INV_X1 U16263 ( .A(n12458), .ZN(n23280) );
  AOI22_X1 U16264 ( .A1(\mem[353][2] ), .A2(n12456), .B1(n26777), .B2(
        data_in[2]), .ZN(n12458) );
  INV_X1 U16265 ( .A(n12459), .ZN(n23279) );
  AOI22_X1 U16266 ( .A1(\mem[353][3] ), .A2(n12456), .B1(n26777), .B2(
        data_in[3]), .ZN(n12459) );
  INV_X1 U16267 ( .A(n12460), .ZN(n23278) );
  AOI22_X1 U16268 ( .A1(\mem[353][4] ), .A2(n12456), .B1(n26777), .B2(
        data_in[4]), .ZN(n12460) );
  INV_X1 U16269 ( .A(n12461), .ZN(n23277) );
  AOI22_X1 U16270 ( .A1(\mem[353][5] ), .A2(n12456), .B1(n26777), .B2(
        data_in[5]), .ZN(n12461) );
  INV_X1 U16271 ( .A(n12462), .ZN(n23276) );
  AOI22_X1 U16272 ( .A1(\mem[353][6] ), .A2(n12456), .B1(n26777), .B2(
        data_in[6]), .ZN(n12462) );
  INV_X1 U16273 ( .A(n12463), .ZN(n23275) );
  AOI22_X1 U16274 ( .A1(\mem[353][7] ), .A2(n12456), .B1(n26777), .B2(
        data_in[7]), .ZN(n12463) );
  INV_X1 U16275 ( .A(n12464), .ZN(n23274) );
  AOI22_X1 U16276 ( .A1(\mem[354][0] ), .A2(n12465), .B1(n26776), .B2(
        data_in[0]), .ZN(n12464) );
  INV_X1 U16277 ( .A(n12466), .ZN(n23273) );
  AOI22_X1 U16278 ( .A1(\mem[354][1] ), .A2(n12465), .B1(n26776), .B2(
        data_in[1]), .ZN(n12466) );
  INV_X1 U16279 ( .A(n12467), .ZN(n23272) );
  AOI22_X1 U16280 ( .A1(\mem[354][2] ), .A2(n12465), .B1(n26776), .B2(
        data_in[2]), .ZN(n12467) );
  INV_X1 U16281 ( .A(n12468), .ZN(n23271) );
  AOI22_X1 U16282 ( .A1(\mem[354][3] ), .A2(n12465), .B1(n26776), .B2(
        data_in[3]), .ZN(n12468) );
  INV_X1 U16283 ( .A(n12469), .ZN(n23270) );
  AOI22_X1 U16284 ( .A1(\mem[354][4] ), .A2(n12465), .B1(n26776), .B2(
        data_in[4]), .ZN(n12469) );
  INV_X1 U16285 ( .A(n12470), .ZN(n23269) );
  AOI22_X1 U16286 ( .A1(\mem[354][5] ), .A2(n12465), .B1(n26776), .B2(
        data_in[5]), .ZN(n12470) );
  INV_X1 U16287 ( .A(n12471), .ZN(n23268) );
  AOI22_X1 U16288 ( .A1(\mem[354][6] ), .A2(n12465), .B1(n26776), .B2(
        data_in[6]), .ZN(n12471) );
  INV_X1 U16289 ( .A(n12472), .ZN(n23267) );
  AOI22_X1 U16290 ( .A1(\mem[354][7] ), .A2(n12465), .B1(n26776), .B2(
        data_in[7]), .ZN(n12472) );
  INV_X1 U16291 ( .A(n12473), .ZN(n23266) );
  AOI22_X1 U16292 ( .A1(\mem[355][0] ), .A2(n12474), .B1(n26775), .B2(
        data_in[0]), .ZN(n12473) );
  INV_X1 U16293 ( .A(n12475), .ZN(n23265) );
  AOI22_X1 U16294 ( .A1(\mem[355][1] ), .A2(n12474), .B1(n26775), .B2(
        data_in[1]), .ZN(n12475) );
  INV_X1 U16295 ( .A(n12476), .ZN(n23264) );
  AOI22_X1 U16296 ( .A1(\mem[355][2] ), .A2(n12474), .B1(n26775), .B2(
        data_in[2]), .ZN(n12476) );
  INV_X1 U16297 ( .A(n12477), .ZN(n23263) );
  AOI22_X1 U16298 ( .A1(\mem[355][3] ), .A2(n12474), .B1(n26775), .B2(
        data_in[3]), .ZN(n12477) );
  INV_X1 U16299 ( .A(n12478), .ZN(n23262) );
  AOI22_X1 U16300 ( .A1(\mem[355][4] ), .A2(n12474), .B1(n26775), .B2(
        data_in[4]), .ZN(n12478) );
  INV_X1 U16301 ( .A(n12479), .ZN(n23261) );
  AOI22_X1 U16302 ( .A1(\mem[355][5] ), .A2(n12474), .B1(n26775), .B2(
        data_in[5]), .ZN(n12479) );
  INV_X1 U16303 ( .A(n12480), .ZN(n23260) );
  AOI22_X1 U16304 ( .A1(\mem[355][6] ), .A2(n12474), .B1(n26775), .B2(
        data_in[6]), .ZN(n12480) );
  INV_X1 U16305 ( .A(n12481), .ZN(n23259) );
  AOI22_X1 U16306 ( .A1(\mem[355][7] ), .A2(n12474), .B1(n26775), .B2(
        data_in[7]), .ZN(n12481) );
  INV_X1 U16307 ( .A(n12482), .ZN(n23258) );
  AOI22_X1 U16308 ( .A1(\mem[356][0] ), .A2(n12483), .B1(n26774), .B2(
        data_in[0]), .ZN(n12482) );
  INV_X1 U16309 ( .A(n12484), .ZN(n23257) );
  AOI22_X1 U16310 ( .A1(\mem[356][1] ), .A2(n12483), .B1(n26774), .B2(
        data_in[1]), .ZN(n12484) );
  INV_X1 U16311 ( .A(n12485), .ZN(n23256) );
  AOI22_X1 U16312 ( .A1(\mem[356][2] ), .A2(n12483), .B1(n26774), .B2(
        data_in[2]), .ZN(n12485) );
  INV_X1 U16313 ( .A(n12486), .ZN(n23255) );
  AOI22_X1 U16314 ( .A1(\mem[356][3] ), .A2(n12483), .B1(n26774), .B2(
        data_in[3]), .ZN(n12486) );
  INV_X1 U16315 ( .A(n12487), .ZN(n23254) );
  AOI22_X1 U16316 ( .A1(\mem[356][4] ), .A2(n12483), .B1(n26774), .B2(
        data_in[4]), .ZN(n12487) );
  INV_X1 U16317 ( .A(n12488), .ZN(n23253) );
  AOI22_X1 U16318 ( .A1(\mem[356][5] ), .A2(n12483), .B1(n26774), .B2(
        data_in[5]), .ZN(n12488) );
  INV_X1 U16319 ( .A(n12489), .ZN(n23252) );
  AOI22_X1 U16320 ( .A1(\mem[356][6] ), .A2(n12483), .B1(n26774), .B2(
        data_in[6]), .ZN(n12489) );
  INV_X1 U16321 ( .A(n12490), .ZN(n23251) );
  AOI22_X1 U16322 ( .A1(\mem[356][7] ), .A2(n12483), .B1(n26774), .B2(
        data_in[7]), .ZN(n12490) );
  INV_X1 U16323 ( .A(n12491), .ZN(n23250) );
  AOI22_X1 U16324 ( .A1(\mem[357][0] ), .A2(n12492), .B1(n26773), .B2(
        data_in[0]), .ZN(n12491) );
  INV_X1 U16325 ( .A(n12493), .ZN(n23249) );
  AOI22_X1 U16326 ( .A1(\mem[357][1] ), .A2(n12492), .B1(n26773), .B2(
        data_in[1]), .ZN(n12493) );
  INV_X1 U16327 ( .A(n12494), .ZN(n23248) );
  AOI22_X1 U16328 ( .A1(\mem[357][2] ), .A2(n12492), .B1(n26773), .B2(
        data_in[2]), .ZN(n12494) );
  INV_X1 U16329 ( .A(n12495), .ZN(n23247) );
  AOI22_X1 U16330 ( .A1(\mem[357][3] ), .A2(n12492), .B1(n26773), .B2(
        data_in[3]), .ZN(n12495) );
  INV_X1 U16331 ( .A(n12496), .ZN(n23246) );
  AOI22_X1 U16332 ( .A1(\mem[357][4] ), .A2(n12492), .B1(n26773), .B2(
        data_in[4]), .ZN(n12496) );
  INV_X1 U16333 ( .A(n12497), .ZN(n23245) );
  AOI22_X1 U16334 ( .A1(\mem[357][5] ), .A2(n12492), .B1(n26773), .B2(
        data_in[5]), .ZN(n12497) );
  INV_X1 U16335 ( .A(n12498), .ZN(n23244) );
  AOI22_X1 U16336 ( .A1(\mem[357][6] ), .A2(n12492), .B1(n26773), .B2(
        data_in[6]), .ZN(n12498) );
  INV_X1 U16337 ( .A(n12499), .ZN(n23243) );
  AOI22_X1 U16338 ( .A1(\mem[357][7] ), .A2(n12492), .B1(n26773), .B2(
        data_in[7]), .ZN(n12499) );
  INV_X1 U16339 ( .A(n12500), .ZN(n23242) );
  AOI22_X1 U16340 ( .A1(\mem[358][0] ), .A2(n12501), .B1(n26772), .B2(
        data_in[0]), .ZN(n12500) );
  INV_X1 U16341 ( .A(n12502), .ZN(n23241) );
  AOI22_X1 U16342 ( .A1(\mem[358][1] ), .A2(n12501), .B1(n26772), .B2(
        data_in[1]), .ZN(n12502) );
  INV_X1 U16343 ( .A(n12503), .ZN(n23240) );
  AOI22_X1 U16344 ( .A1(\mem[358][2] ), .A2(n12501), .B1(n26772), .B2(
        data_in[2]), .ZN(n12503) );
  INV_X1 U16345 ( .A(n12504), .ZN(n23239) );
  AOI22_X1 U16346 ( .A1(\mem[358][3] ), .A2(n12501), .B1(n26772), .B2(
        data_in[3]), .ZN(n12504) );
  INV_X1 U16347 ( .A(n12505), .ZN(n23238) );
  AOI22_X1 U16348 ( .A1(\mem[358][4] ), .A2(n12501), .B1(n26772), .B2(
        data_in[4]), .ZN(n12505) );
  INV_X1 U16349 ( .A(n12506), .ZN(n23237) );
  AOI22_X1 U16350 ( .A1(\mem[358][5] ), .A2(n12501), .B1(n26772), .B2(
        data_in[5]), .ZN(n12506) );
  INV_X1 U16351 ( .A(n12507), .ZN(n23236) );
  AOI22_X1 U16352 ( .A1(\mem[358][6] ), .A2(n12501), .B1(n26772), .B2(
        data_in[6]), .ZN(n12507) );
  INV_X1 U16353 ( .A(n12508), .ZN(n23235) );
  AOI22_X1 U16354 ( .A1(\mem[358][7] ), .A2(n12501), .B1(n26772), .B2(
        data_in[7]), .ZN(n12508) );
  INV_X1 U16355 ( .A(n12509), .ZN(n23234) );
  AOI22_X1 U16356 ( .A1(\mem[359][0] ), .A2(n12510), .B1(n26771), .B2(
        data_in[0]), .ZN(n12509) );
  INV_X1 U16357 ( .A(n12511), .ZN(n23233) );
  AOI22_X1 U16358 ( .A1(\mem[359][1] ), .A2(n12510), .B1(n26771), .B2(
        data_in[1]), .ZN(n12511) );
  INV_X1 U16359 ( .A(n12512), .ZN(n23232) );
  AOI22_X1 U16360 ( .A1(\mem[359][2] ), .A2(n12510), .B1(n26771), .B2(
        data_in[2]), .ZN(n12512) );
  INV_X1 U16361 ( .A(n12513), .ZN(n23231) );
  AOI22_X1 U16362 ( .A1(\mem[359][3] ), .A2(n12510), .B1(n26771), .B2(
        data_in[3]), .ZN(n12513) );
  INV_X1 U16363 ( .A(n12514), .ZN(n23230) );
  AOI22_X1 U16364 ( .A1(\mem[359][4] ), .A2(n12510), .B1(n26771), .B2(
        data_in[4]), .ZN(n12514) );
  INV_X1 U16365 ( .A(n12515), .ZN(n23229) );
  AOI22_X1 U16366 ( .A1(\mem[359][5] ), .A2(n12510), .B1(n26771), .B2(
        data_in[5]), .ZN(n12515) );
  INV_X1 U16367 ( .A(n12516), .ZN(n23228) );
  AOI22_X1 U16368 ( .A1(\mem[359][6] ), .A2(n12510), .B1(n26771), .B2(
        data_in[6]), .ZN(n12516) );
  INV_X1 U16369 ( .A(n12517), .ZN(n23227) );
  AOI22_X1 U16370 ( .A1(\mem[359][7] ), .A2(n12510), .B1(n26771), .B2(
        data_in[7]), .ZN(n12517) );
  INV_X1 U16371 ( .A(n12734), .ZN(n23034) );
  AOI22_X1 U16372 ( .A1(\mem[384][0] ), .A2(n12735), .B1(n26746), .B2(
        data_in[0]), .ZN(n12734) );
  INV_X1 U16373 ( .A(n12736), .ZN(n23033) );
  AOI22_X1 U16374 ( .A1(\mem[384][1] ), .A2(n12735), .B1(n26746), .B2(
        data_in[1]), .ZN(n12736) );
  INV_X1 U16375 ( .A(n12737), .ZN(n23032) );
  AOI22_X1 U16376 ( .A1(\mem[384][2] ), .A2(n12735), .B1(n26746), .B2(
        data_in[2]), .ZN(n12737) );
  INV_X1 U16377 ( .A(n12738), .ZN(n23031) );
  AOI22_X1 U16378 ( .A1(\mem[384][3] ), .A2(n12735), .B1(n26746), .B2(
        data_in[3]), .ZN(n12738) );
  INV_X1 U16379 ( .A(n12739), .ZN(n23030) );
  AOI22_X1 U16380 ( .A1(\mem[384][4] ), .A2(n12735), .B1(n26746), .B2(
        data_in[4]), .ZN(n12739) );
  INV_X1 U16381 ( .A(n12740), .ZN(n23029) );
  AOI22_X1 U16382 ( .A1(\mem[384][5] ), .A2(n12735), .B1(n26746), .B2(
        data_in[5]), .ZN(n12740) );
  INV_X1 U16383 ( .A(n12741), .ZN(n23028) );
  AOI22_X1 U16384 ( .A1(\mem[384][6] ), .A2(n12735), .B1(n26746), .B2(
        data_in[6]), .ZN(n12741) );
  INV_X1 U16385 ( .A(n12742), .ZN(n23027) );
  AOI22_X1 U16386 ( .A1(\mem[384][7] ), .A2(n12735), .B1(n26746), .B2(
        data_in[7]), .ZN(n12742) );
  INV_X1 U16387 ( .A(n12744), .ZN(n23026) );
  AOI22_X1 U16388 ( .A1(\mem[385][0] ), .A2(n12745), .B1(n26745), .B2(
        data_in[0]), .ZN(n12744) );
  INV_X1 U16389 ( .A(n12746), .ZN(n23025) );
  AOI22_X1 U16390 ( .A1(\mem[385][1] ), .A2(n12745), .B1(n26745), .B2(
        data_in[1]), .ZN(n12746) );
  INV_X1 U16391 ( .A(n12747), .ZN(n23024) );
  AOI22_X1 U16392 ( .A1(\mem[385][2] ), .A2(n12745), .B1(n26745), .B2(
        data_in[2]), .ZN(n12747) );
  INV_X1 U16393 ( .A(n12748), .ZN(n23023) );
  AOI22_X1 U16394 ( .A1(\mem[385][3] ), .A2(n12745), .B1(n26745), .B2(
        data_in[3]), .ZN(n12748) );
  INV_X1 U16395 ( .A(n12749), .ZN(n23022) );
  AOI22_X1 U16396 ( .A1(\mem[385][4] ), .A2(n12745), .B1(n26745), .B2(
        data_in[4]), .ZN(n12749) );
  INV_X1 U16397 ( .A(n12750), .ZN(n23021) );
  AOI22_X1 U16398 ( .A1(\mem[385][5] ), .A2(n12745), .B1(n26745), .B2(
        data_in[5]), .ZN(n12750) );
  INV_X1 U16399 ( .A(n12751), .ZN(n23020) );
  AOI22_X1 U16400 ( .A1(\mem[385][6] ), .A2(n12745), .B1(n26745), .B2(
        data_in[6]), .ZN(n12751) );
  INV_X1 U16401 ( .A(n12752), .ZN(n23019) );
  AOI22_X1 U16402 ( .A1(\mem[385][7] ), .A2(n12745), .B1(n26745), .B2(
        data_in[7]), .ZN(n12752) );
  INV_X1 U16403 ( .A(n12753), .ZN(n23018) );
  AOI22_X1 U16404 ( .A1(\mem[386][0] ), .A2(n12754), .B1(n26744), .B2(
        data_in[0]), .ZN(n12753) );
  INV_X1 U16405 ( .A(n12755), .ZN(n23017) );
  AOI22_X1 U16406 ( .A1(\mem[386][1] ), .A2(n12754), .B1(n26744), .B2(
        data_in[1]), .ZN(n12755) );
  INV_X1 U16407 ( .A(n12756), .ZN(n23016) );
  AOI22_X1 U16408 ( .A1(\mem[386][2] ), .A2(n12754), .B1(n26744), .B2(
        data_in[2]), .ZN(n12756) );
  INV_X1 U16409 ( .A(n12757), .ZN(n23015) );
  AOI22_X1 U16410 ( .A1(\mem[386][3] ), .A2(n12754), .B1(n26744), .B2(
        data_in[3]), .ZN(n12757) );
  INV_X1 U16411 ( .A(n12758), .ZN(n23014) );
  AOI22_X1 U16412 ( .A1(\mem[386][4] ), .A2(n12754), .B1(n26744), .B2(
        data_in[4]), .ZN(n12758) );
  INV_X1 U16413 ( .A(n12759), .ZN(n23013) );
  AOI22_X1 U16414 ( .A1(\mem[386][5] ), .A2(n12754), .B1(n26744), .B2(
        data_in[5]), .ZN(n12759) );
  INV_X1 U16415 ( .A(n12760), .ZN(n23012) );
  AOI22_X1 U16416 ( .A1(\mem[386][6] ), .A2(n12754), .B1(n26744), .B2(
        data_in[6]), .ZN(n12760) );
  INV_X1 U16417 ( .A(n12761), .ZN(n23011) );
  AOI22_X1 U16418 ( .A1(\mem[386][7] ), .A2(n12754), .B1(n26744), .B2(
        data_in[7]), .ZN(n12761) );
  INV_X1 U16419 ( .A(n12762), .ZN(n23010) );
  AOI22_X1 U16420 ( .A1(\mem[387][0] ), .A2(n12763), .B1(n26743), .B2(
        data_in[0]), .ZN(n12762) );
  INV_X1 U16421 ( .A(n12764), .ZN(n23009) );
  AOI22_X1 U16422 ( .A1(\mem[387][1] ), .A2(n12763), .B1(n26743), .B2(
        data_in[1]), .ZN(n12764) );
  INV_X1 U16423 ( .A(n12765), .ZN(n23008) );
  AOI22_X1 U16424 ( .A1(\mem[387][2] ), .A2(n12763), .B1(n26743), .B2(
        data_in[2]), .ZN(n12765) );
  INV_X1 U16425 ( .A(n12766), .ZN(n23007) );
  AOI22_X1 U16426 ( .A1(\mem[387][3] ), .A2(n12763), .B1(n26743), .B2(
        data_in[3]), .ZN(n12766) );
  INV_X1 U16427 ( .A(n12767), .ZN(n23006) );
  AOI22_X1 U16428 ( .A1(\mem[387][4] ), .A2(n12763), .B1(n26743), .B2(
        data_in[4]), .ZN(n12767) );
  INV_X1 U16429 ( .A(n12768), .ZN(n23005) );
  AOI22_X1 U16430 ( .A1(\mem[387][5] ), .A2(n12763), .B1(n26743), .B2(
        data_in[5]), .ZN(n12768) );
  INV_X1 U16431 ( .A(n12769), .ZN(n23004) );
  AOI22_X1 U16432 ( .A1(\mem[387][6] ), .A2(n12763), .B1(n26743), .B2(
        data_in[6]), .ZN(n12769) );
  INV_X1 U16433 ( .A(n12770), .ZN(n23003) );
  AOI22_X1 U16434 ( .A1(\mem[387][7] ), .A2(n12763), .B1(n26743), .B2(
        data_in[7]), .ZN(n12770) );
  INV_X1 U16435 ( .A(n12771), .ZN(n23002) );
  AOI22_X1 U16436 ( .A1(\mem[388][0] ), .A2(n12772), .B1(n26742), .B2(
        data_in[0]), .ZN(n12771) );
  INV_X1 U16437 ( .A(n12773), .ZN(n23001) );
  AOI22_X1 U16438 ( .A1(\mem[388][1] ), .A2(n12772), .B1(n26742), .B2(
        data_in[1]), .ZN(n12773) );
  INV_X1 U16439 ( .A(n12774), .ZN(n23000) );
  AOI22_X1 U16440 ( .A1(\mem[388][2] ), .A2(n12772), .B1(n26742), .B2(
        data_in[2]), .ZN(n12774) );
  INV_X1 U16441 ( .A(n12775), .ZN(n22999) );
  AOI22_X1 U16442 ( .A1(\mem[388][3] ), .A2(n12772), .B1(n26742), .B2(
        data_in[3]), .ZN(n12775) );
  INV_X1 U16443 ( .A(n12776), .ZN(n22998) );
  AOI22_X1 U16444 ( .A1(\mem[388][4] ), .A2(n12772), .B1(n26742), .B2(
        data_in[4]), .ZN(n12776) );
  INV_X1 U16445 ( .A(n12777), .ZN(n22997) );
  AOI22_X1 U16446 ( .A1(\mem[388][5] ), .A2(n12772), .B1(n26742), .B2(
        data_in[5]), .ZN(n12777) );
  INV_X1 U16447 ( .A(n12778), .ZN(n22996) );
  AOI22_X1 U16448 ( .A1(\mem[388][6] ), .A2(n12772), .B1(n26742), .B2(
        data_in[6]), .ZN(n12778) );
  INV_X1 U16449 ( .A(n12779), .ZN(n22995) );
  AOI22_X1 U16450 ( .A1(\mem[388][7] ), .A2(n12772), .B1(n26742), .B2(
        data_in[7]), .ZN(n12779) );
  INV_X1 U16451 ( .A(n12780), .ZN(n22994) );
  AOI22_X1 U16452 ( .A1(\mem[389][0] ), .A2(n12781), .B1(n26741), .B2(
        data_in[0]), .ZN(n12780) );
  INV_X1 U16453 ( .A(n12782), .ZN(n22993) );
  AOI22_X1 U16454 ( .A1(\mem[389][1] ), .A2(n12781), .B1(n26741), .B2(
        data_in[1]), .ZN(n12782) );
  INV_X1 U16455 ( .A(n12783), .ZN(n22992) );
  AOI22_X1 U16456 ( .A1(\mem[389][2] ), .A2(n12781), .B1(n26741), .B2(
        data_in[2]), .ZN(n12783) );
  INV_X1 U16457 ( .A(n12784), .ZN(n22991) );
  AOI22_X1 U16458 ( .A1(\mem[389][3] ), .A2(n12781), .B1(n26741), .B2(
        data_in[3]), .ZN(n12784) );
  INV_X1 U16459 ( .A(n12785), .ZN(n22990) );
  AOI22_X1 U16460 ( .A1(\mem[389][4] ), .A2(n12781), .B1(n26741), .B2(
        data_in[4]), .ZN(n12785) );
  INV_X1 U16461 ( .A(n12786), .ZN(n22989) );
  AOI22_X1 U16462 ( .A1(\mem[389][5] ), .A2(n12781), .B1(n26741), .B2(
        data_in[5]), .ZN(n12786) );
  INV_X1 U16463 ( .A(n12787), .ZN(n22988) );
  AOI22_X1 U16464 ( .A1(\mem[389][6] ), .A2(n12781), .B1(n26741), .B2(
        data_in[6]), .ZN(n12787) );
  INV_X1 U16465 ( .A(n12788), .ZN(n22987) );
  AOI22_X1 U16466 ( .A1(\mem[389][7] ), .A2(n12781), .B1(n26741), .B2(
        data_in[7]), .ZN(n12788) );
  INV_X1 U16467 ( .A(n12789), .ZN(n22986) );
  AOI22_X1 U16468 ( .A1(\mem[390][0] ), .A2(n12790), .B1(n26740), .B2(
        data_in[0]), .ZN(n12789) );
  INV_X1 U16469 ( .A(n12791), .ZN(n22985) );
  AOI22_X1 U16470 ( .A1(\mem[390][1] ), .A2(n12790), .B1(n26740), .B2(
        data_in[1]), .ZN(n12791) );
  INV_X1 U16471 ( .A(n12792), .ZN(n22984) );
  AOI22_X1 U16472 ( .A1(\mem[390][2] ), .A2(n12790), .B1(n26740), .B2(
        data_in[2]), .ZN(n12792) );
  INV_X1 U16473 ( .A(n12793), .ZN(n22983) );
  AOI22_X1 U16474 ( .A1(\mem[390][3] ), .A2(n12790), .B1(n26740), .B2(
        data_in[3]), .ZN(n12793) );
  INV_X1 U16475 ( .A(n12794), .ZN(n22982) );
  AOI22_X1 U16476 ( .A1(\mem[390][4] ), .A2(n12790), .B1(n26740), .B2(
        data_in[4]), .ZN(n12794) );
  INV_X1 U16477 ( .A(n12795), .ZN(n22981) );
  AOI22_X1 U16478 ( .A1(\mem[390][5] ), .A2(n12790), .B1(n26740), .B2(
        data_in[5]), .ZN(n12795) );
  INV_X1 U16479 ( .A(n12796), .ZN(n22980) );
  AOI22_X1 U16480 ( .A1(\mem[390][6] ), .A2(n12790), .B1(n26740), .B2(
        data_in[6]), .ZN(n12796) );
  INV_X1 U16481 ( .A(n12797), .ZN(n22979) );
  AOI22_X1 U16482 ( .A1(\mem[390][7] ), .A2(n12790), .B1(n26740), .B2(
        data_in[7]), .ZN(n12797) );
  INV_X1 U16483 ( .A(n12798), .ZN(n22978) );
  AOI22_X1 U16484 ( .A1(\mem[391][0] ), .A2(n12799), .B1(n26739), .B2(
        data_in[0]), .ZN(n12798) );
  INV_X1 U16485 ( .A(n12800), .ZN(n22977) );
  AOI22_X1 U16486 ( .A1(\mem[391][1] ), .A2(n12799), .B1(n26739), .B2(
        data_in[1]), .ZN(n12800) );
  INV_X1 U16487 ( .A(n12801), .ZN(n22976) );
  AOI22_X1 U16488 ( .A1(\mem[391][2] ), .A2(n12799), .B1(n26739), .B2(
        data_in[2]), .ZN(n12801) );
  INV_X1 U16489 ( .A(n12802), .ZN(n22975) );
  AOI22_X1 U16490 ( .A1(\mem[391][3] ), .A2(n12799), .B1(n26739), .B2(
        data_in[3]), .ZN(n12802) );
  INV_X1 U16491 ( .A(n12803), .ZN(n22974) );
  AOI22_X1 U16492 ( .A1(\mem[391][4] ), .A2(n12799), .B1(n26739), .B2(
        data_in[4]), .ZN(n12803) );
  INV_X1 U16493 ( .A(n12804), .ZN(n22973) );
  AOI22_X1 U16494 ( .A1(\mem[391][5] ), .A2(n12799), .B1(n26739), .B2(
        data_in[5]), .ZN(n12804) );
  INV_X1 U16495 ( .A(n12805), .ZN(n22972) );
  AOI22_X1 U16496 ( .A1(\mem[391][6] ), .A2(n12799), .B1(n26739), .B2(
        data_in[6]), .ZN(n12805) );
  INV_X1 U16497 ( .A(n12806), .ZN(n22971) );
  AOI22_X1 U16498 ( .A1(\mem[391][7] ), .A2(n12799), .B1(n26739), .B2(
        data_in[7]), .ZN(n12806) );
  INV_X1 U16499 ( .A(n13023), .ZN(n22778) );
  AOI22_X1 U16500 ( .A1(\mem[416][0] ), .A2(n13024), .B1(n26714), .B2(
        data_in[0]), .ZN(n13023) );
  INV_X1 U16501 ( .A(n13025), .ZN(n22777) );
  AOI22_X1 U16502 ( .A1(\mem[416][1] ), .A2(n13024), .B1(n26714), .B2(
        data_in[1]), .ZN(n13025) );
  INV_X1 U16503 ( .A(n13026), .ZN(n22776) );
  AOI22_X1 U16504 ( .A1(\mem[416][2] ), .A2(n13024), .B1(n26714), .B2(
        data_in[2]), .ZN(n13026) );
  INV_X1 U16505 ( .A(n13027), .ZN(n22775) );
  AOI22_X1 U16506 ( .A1(\mem[416][3] ), .A2(n13024), .B1(n26714), .B2(
        data_in[3]), .ZN(n13027) );
  INV_X1 U16507 ( .A(n13028), .ZN(n22774) );
  AOI22_X1 U16508 ( .A1(\mem[416][4] ), .A2(n13024), .B1(n26714), .B2(
        data_in[4]), .ZN(n13028) );
  INV_X1 U16509 ( .A(n13029), .ZN(n22773) );
  AOI22_X1 U16510 ( .A1(\mem[416][5] ), .A2(n13024), .B1(n26714), .B2(
        data_in[5]), .ZN(n13029) );
  INV_X1 U16511 ( .A(n13030), .ZN(n22772) );
  AOI22_X1 U16512 ( .A1(\mem[416][6] ), .A2(n13024), .B1(n26714), .B2(
        data_in[6]), .ZN(n13030) );
  INV_X1 U16513 ( .A(n13031), .ZN(n22771) );
  AOI22_X1 U16514 ( .A1(\mem[416][7] ), .A2(n13024), .B1(n26714), .B2(
        data_in[7]), .ZN(n13031) );
  INV_X1 U16515 ( .A(n13033), .ZN(n22770) );
  AOI22_X1 U16516 ( .A1(\mem[417][0] ), .A2(n13034), .B1(n26713), .B2(
        data_in[0]), .ZN(n13033) );
  INV_X1 U16517 ( .A(n13035), .ZN(n22769) );
  AOI22_X1 U16518 ( .A1(\mem[417][1] ), .A2(n13034), .B1(n26713), .B2(
        data_in[1]), .ZN(n13035) );
  INV_X1 U16519 ( .A(n13036), .ZN(n22768) );
  AOI22_X1 U16520 ( .A1(\mem[417][2] ), .A2(n13034), .B1(n26713), .B2(
        data_in[2]), .ZN(n13036) );
  INV_X1 U16521 ( .A(n13037), .ZN(n22767) );
  AOI22_X1 U16522 ( .A1(\mem[417][3] ), .A2(n13034), .B1(n26713), .B2(
        data_in[3]), .ZN(n13037) );
  INV_X1 U16523 ( .A(n13038), .ZN(n22766) );
  AOI22_X1 U16524 ( .A1(\mem[417][4] ), .A2(n13034), .B1(n26713), .B2(
        data_in[4]), .ZN(n13038) );
  INV_X1 U16525 ( .A(n13039), .ZN(n22765) );
  AOI22_X1 U16526 ( .A1(\mem[417][5] ), .A2(n13034), .B1(n26713), .B2(
        data_in[5]), .ZN(n13039) );
  INV_X1 U16527 ( .A(n13040), .ZN(n22764) );
  AOI22_X1 U16528 ( .A1(\mem[417][6] ), .A2(n13034), .B1(n26713), .B2(
        data_in[6]), .ZN(n13040) );
  INV_X1 U16529 ( .A(n13041), .ZN(n22763) );
  AOI22_X1 U16530 ( .A1(\mem[417][7] ), .A2(n13034), .B1(n26713), .B2(
        data_in[7]), .ZN(n13041) );
  INV_X1 U16531 ( .A(n13042), .ZN(n22762) );
  AOI22_X1 U16532 ( .A1(\mem[418][0] ), .A2(n13043), .B1(n26712), .B2(
        data_in[0]), .ZN(n13042) );
  INV_X1 U16533 ( .A(n13044), .ZN(n22761) );
  AOI22_X1 U16534 ( .A1(\mem[418][1] ), .A2(n13043), .B1(n26712), .B2(
        data_in[1]), .ZN(n13044) );
  INV_X1 U16535 ( .A(n13045), .ZN(n22760) );
  AOI22_X1 U16536 ( .A1(\mem[418][2] ), .A2(n13043), .B1(n26712), .B2(
        data_in[2]), .ZN(n13045) );
  INV_X1 U16537 ( .A(n13046), .ZN(n22759) );
  AOI22_X1 U16538 ( .A1(\mem[418][3] ), .A2(n13043), .B1(n26712), .B2(
        data_in[3]), .ZN(n13046) );
  INV_X1 U16539 ( .A(n13047), .ZN(n22758) );
  AOI22_X1 U16540 ( .A1(\mem[418][4] ), .A2(n13043), .B1(n26712), .B2(
        data_in[4]), .ZN(n13047) );
  INV_X1 U16541 ( .A(n13048), .ZN(n22757) );
  AOI22_X1 U16542 ( .A1(\mem[418][5] ), .A2(n13043), .B1(n26712), .B2(
        data_in[5]), .ZN(n13048) );
  INV_X1 U16543 ( .A(n13049), .ZN(n22756) );
  AOI22_X1 U16544 ( .A1(\mem[418][6] ), .A2(n13043), .B1(n26712), .B2(
        data_in[6]), .ZN(n13049) );
  INV_X1 U16545 ( .A(n13050), .ZN(n22755) );
  AOI22_X1 U16546 ( .A1(\mem[418][7] ), .A2(n13043), .B1(n26712), .B2(
        data_in[7]), .ZN(n13050) );
  INV_X1 U16547 ( .A(n13051), .ZN(n22754) );
  AOI22_X1 U16548 ( .A1(\mem[419][0] ), .A2(n13052), .B1(n26711), .B2(
        data_in[0]), .ZN(n13051) );
  INV_X1 U16549 ( .A(n13053), .ZN(n22753) );
  AOI22_X1 U16550 ( .A1(\mem[419][1] ), .A2(n13052), .B1(n26711), .B2(
        data_in[1]), .ZN(n13053) );
  INV_X1 U16551 ( .A(n13054), .ZN(n22752) );
  AOI22_X1 U16552 ( .A1(\mem[419][2] ), .A2(n13052), .B1(n26711), .B2(
        data_in[2]), .ZN(n13054) );
  INV_X1 U16553 ( .A(n13055), .ZN(n22751) );
  AOI22_X1 U16554 ( .A1(\mem[419][3] ), .A2(n13052), .B1(n26711), .B2(
        data_in[3]), .ZN(n13055) );
  INV_X1 U16555 ( .A(n13056), .ZN(n22750) );
  AOI22_X1 U16556 ( .A1(\mem[419][4] ), .A2(n13052), .B1(n26711), .B2(
        data_in[4]), .ZN(n13056) );
  INV_X1 U16557 ( .A(n13057), .ZN(n22749) );
  AOI22_X1 U16558 ( .A1(\mem[419][5] ), .A2(n13052), .B1(n26711), .B2(
        data_in[5]), .ZN(n13057) );
  INV_X1 U16559 ( .A(n13058), .ZN(n22748) );
  AOI22_X1 U16560 ( .A1(\mem[419][6] ), .A2(n13052), .B1(n26711), .B2(
        data_in[6]), .ZN(n13058) );
  INV_X1 U16561 ( .A(n13059), .ZN(n22747) );
  AOI22_X1 U16562 ( .A1(\mem[419][7] ), .A2(n13052), .B1(n26711), .B2(
        data_in[7]), .ZN(n13059) );
  INV_X1 U16563 ( .A(n13060), .ZN(n22746) );
  AOI22_X1 U16564 ( .A1(\mem[420][0] ), .A2(n13061), .B1(n26710), .B2(
        data_in[0]), .ZN(n13060) );
  INV_X1 U16565 ( .A(n13062), .ZN(n22745) );
  AOI22_X1 U16566 ( .A1(\mem[420][1] ), .A2(n13061), .B1(n26710), .B2(
        data_in[1]), .ZN(n13062) );
  INV_X1 U16567 ( .A(n13063), .ZN(n22744) );
  AOI22_X1 U16568 ( .A1(\mem[420][2] ), .A2(n13061), .B1(n26710), .B2(
        data_in[2]), .ZN(n13063) );
  INV_X1 U16569 ( .A(n13064), .ZN(n22743) );
  AOI22_X1 U16570 ( .A1(\mem[420][3] ), .A2(n13061), .B1(n26710), .B2(
        data_in[3]), .ZN(n13064) );
  INV_X1 U16571 ( .A(n13065), .ZN(n22742) );
  AOI22_X1 U16572 ( .A1(\mem[420][4] ), .A2(n13061), .B1(n26710), .B2(
        data_in[4]), .ZN(n13065) );
  INV_X1 U16573 ( .A(n13066), .ZN(n22741) );
  AOI22_X1 U16574 ( .A1(\mem[420][5] ), .A2(n13061), .B1(n26710), .B2(
        data_in[5]), .ZN(n13066) );
  INV_X1 U16575 ( .A(n13067), .ZN(n22740) );
  AOI22_X1 U16576 ( .A1(\mem[420][6] ), .A2(n13061), .B1(n26710), .B2(
        data_in[6]), .ZN(n13067) );
  INV_X1 U16577 ( .A(n13068), .ZN(n22739) );
  AOI22_X1 U16578 ( .A1(\mem[420][7] ), .A2(n13061), .B1(n26710), .B2(
        data_in[7]), .ZN(n13068) );
  INV_X1 U16579 ( .A(n13069), .ZN(n22738) );
  AOI22_X1 U16580 ( .A1(\mem[421][0] ), .A2(n13070), .B1(n26709), .B2(
        data_in[0]), .ZN(n13069) );
  INV_X1 U16581 ( .A(n13071), .ZN(n22737) );
  AOI22_X1 U16582 ( .A1(\mem[421][1] ), .A2(n13070), .B1(n26709), .B2(
        data_in[1]), .ZN(n13071) );
  INV_X1 U16583 ( .A(n13072), .ZN(n22736) );
  AOI22_X1 U16584 ( .A1(\mem[421][2] ), .A2(n13070), .B1(n26709), .B2(
        data_in[2]), .ZN(n13072) );
  INV_X1 U16585 ( .A(n13073), .ZN(n22735) );
  AOI22_X1 U16586 ( .A1(\mem[421][3] ), .A2(n13070), .B1(n26709), .B2(
        data_in[3]), .ZN(n13073) );
  INV_X1 U16587 ( .A(n13074), .ZN(n22734) );
  AOI22_X1 U16588 ( .A1(\mem[421][4] ), .A2(n13070), .B1(n26709), .B2(
        data_in[4]), .ZN(n13074) );
  INV_X1 U16589 ( .A(n13075), .ZN(n22733) );
  AOI22_X1 U16590 ( .A1(\mem[421][5] ), .A2(n13070), .B1(n26709), .B2(
        data_in[5]), .ZN(n13075) );
  INV_X1 U16591 ( .A(n13076), .ZN(n22732) );
  AOI22_X1 U16592 ( .A1(\mem[421][6] ), .A2(n13070), .B1(n26709), .B2(
        data_in[6]), .ZN(n13076) );
  INV_X1 U16593 ( .A(n13077), .ZN(n22731) );
  AOI22_X1 U16594 ( .A1(\mem[421][7] ), .A2(n13070), .B1(n26709), .B2(
        data_in[7]), .ZN(n13077) );
  INV_X1 U16595 ( .A(n13078), .ZN(n22730) );
  AOI22_X1 U16596 ( .A1(\mem[422][0] ), .A2(n13079), .B1(n26708), .B2(
        data_in[0]), .ZN(n13078) );
  INV_X1 U16597 ( .A(n13080), .ZN(n22729) );
  AOI22_X1 U16598 ( .A1(\mem[422][1] ), .A2(n13079), .B1(n26708), .B2(
        data_in[1]), .ZN(n13080) );
  INV_X1 U16599 ( .A(n13081), .ZN(n22728) );
  AOI22_X1 U16600 ( .A1(\mem[422][2] ), .A2(n13079), .B1(n26708), .B2(
        data_in[2]), .ZN(n13081) );
  INV_X1 U16601 ( .A(n13082), .ZN(n22727) );
  AOI22_X1 U16602 ( .A1(\mem[422][3] ), .A2(n13079), .B1(n26708), .B2(
        data_in[3]), .ZN(n13082) );
  INV_X1 U16603 ( .A(n13083), .ZN(n22726) );
  AOI22_X1 U16604 ( .A1(\mem[422][4] ), .A2(n13079), .B1(n26708), .B2(
        data_in[4]), .ZN(n13083) );
  INV_X1 U16605 ( .A(n13084), .ZN(n22725) );
  AOI22_X1 U16606 ( .A1(\mem[422][5] ), .A2(n13079), .B1(n26708), .B2(
        data_in[5]), .ZN(n13084) );
  INV_X1 U16607 ( .A(n13085), .ZN(n22724) );
  AOI22_X1 U16608 ( .A1(\mem[422][6] ), .A2(n13079), .B1(n26708), .B2(
        data_in[6]), .ZN(n13085) );
  INV_X1 U16609 ( .A(n13086), .ZN(n22723) );
  AOI22_X1 U16610 ( .A1(\mem[422][7] ), .A2(n13079), .B1(n26708), .B2(
        data_in[7]), .ZN(n13086) );
  INV_X1 U16611 ( .A(n13087), .ZN(n22722) );
  AOI22_X1 U16612 ( .A1(\mem[423][0] ), .A2(n13088), .B1(n26707), .B2(
        data_in[0]), .ZN(n13087) );
  INV_X1 U16613 ( .A(n13089), .ZN(n22721) );
  AOI22_X1 U16614 ( .A1(\mem[423][1] ), .A2(n13088), .B1(n26707), .B2(
        data_in[1]), .ZN(n13089) );
  INV_X1 U16615 ( .A(n13090), .ZN(n22720) );
  AOI22_X1 U16616 ( .A1(\mem[423][2] ), .A2(n13088), .B1(n26707), .B2(
        data_in[2]), .ZN(n13090) );
  INV_X1 U16617 ( .A(n13091), .ZN(n22719) );
  AOI22_X1 U16618 ( .A1(\mem[423][3] ), .A2(n13088), .B1(n26707), .B2(
        data_in[3]), .ZN(n13091) );
  INV_X1 U16619 ( .A(n13092), .ZN(n22718) );
  AOI22_X1 U16620 ( .A1(\mem[423][4] ), .A2(n13088), .B1(n26707), .B2(
        data_in[4]), .ZN(n13092) );
  INV_X1 U16621 ( .A(n13093), .ZN(n22717) );
  AOI22_X1 U16622 ( .A1(\mem[423][5] ), .A2(n13088), .B1(n26707), .B2(
        data_in[5]), .ZN(n13093) );
  INV_X1 U16623 ( .A(n13094), .ZN(n22716) );
  AOI22_X1 U16624 ( .A1(\mem[423][6] ), .A2(n13088), .B1(n26707), .B2(
        data_in[6]), .ZN(n13094) );
  INV_X1 U16625 ( .A(n13095), .ZN(n22715) );
  AOI22_X1 U16626 ( .A1(\mem[423][7] ), .A2(n13088), .B1(n26707), .B2(
        data_in[7]), .ZN(n13095) );
  INV_X1 U16627 ( .A(n13312), .ZN(n22522) );
  AOI22_X1 U16628 ( .A1(\mem[448][0] ), .A2(n13313), .B1(n26682), .B2(
        data_in[0]), .ZN(n13312) );
  INV_X1 U16629 ( .A(n13314), .ZN(n22521) );
  AOI22_X1 U16630 ( .A1(\mem[448][1] ), .A2(n13313), .B1(n26682), .B2(
        data_in[1]), .ZN(n13314) );
  INV_X1 U16631 ( .A(n13315), .ZN(n22520) );
  AOI22_X1 U16632 ( .A1(\mem[448][2] ), .A2(n13313), .B1(n26682), .B2(
        data_in[2]), .ZN(n13315) );
  INV_X1 U16633 ( .A(n13316), .ZN(n22519) );
  AOI22_X1 U16634 ( .A1(\mem[448][3] ), .A2(n13313), .B1(n26682), .B2(
        data_in[3]), .ZN(n13316) );
  INV_X1 U16635 ( .A(n13317), .ZN(n22518) );
  AOI22_X1 U16636 ( .A1(\mem[448][4] ), .A2(n13313), .B1(n26682), .B2(
        data_in[4]), .ZN(n13317) );
  INV_X1 U16637 ( .A(n13318), .ZN(n22517) );
  AOI22_X1 U16638 ( .A1(\mem[448][5] ), .A2(n13313), .B1(n26682), .B2(
        data_in[5]), .ZN(n13318) );
  INV_X1 U16639 ( .A(n13319), .ZN(n22516) );
  AOI22_X1 U16640 ( .A1(\mem[448][6] ), .A2(n13313), .B1(n26682), .B2(
        data_in[6]), .ZN(n13319) );
  INV_X1 U16641 ( .A(n13320), .ZN(n22515) );
  AOI22_X1 U16642 ( .A1(\mem[448][7] ), .A2(n13313), .B1(n26682), .B2(
        data_in[7]), .ZN(n13320) );
  INV_X1 U16643 ( .A(n13322), .ZN(n22514) );
  AOI22_X1 U16644 ( .A1(\mem[449][0] ), .A2(n13323), .B1(n26681), .B2(
        data_in[0]), .ZN(n13322) );
  INV_X1 U16645 ( .A(n13324), .ZN(n22513) );
  AOI22_X1 U16646 ( .A1(\mem[449][1] ), .A2(n13323), .B1(n26681), .B2(
        data_in[1]), .ZN(n13324) );
  INV_X1 U16647 ( .A(n13325), .ZN(n22512) );
  AOI22_X1 U16648 ( .A1(\mem[449][2] ), .A2(n13323), .B1(n26681), .B2(
        data_in[2]), .ZN(n13325) );
  INV_X1 U16649 ( .A(n13326), .ZN(n22511) );
  AOI22_X1 U16650 ( .A1(\mem[449][3] ), .A2(n13323), .B1(n26681), .B2(
        data_in[3]), .ZN(n13326) );
  INV_X1 U16651 ( .A(n13327), .ZN(n22510) );
  AOI22_X1 U16652 ( .A1(\mem[449][4] ), .A2(n13323), .B1(n26681), .B2(
        data_in[4]), .ZN(n13327) );
  INV_X1 U16653 ( .A(n13328), .ZN(n22509) );
  AOI22_X1 U16654 ( .A1(\mem[449][5] ), .A2(n13323), .B1(n26681), .B2(
        data_in[5]), .ZN(n13328) );
  INV_X1 U16655 ( .A(n13329), .ZN(n22508) );
  AOI22_X1 U16656 ( .A1(\mem[449][6] ), .A2(n13323), .B1(n26681), .B2(
        data_in[6]), .ZN(n13329) );
  INV_X1 U16657 ( .A(n13330), .ZN(n22507) );
  AOI22_X1 U16658 ( .A1(\mem[449][7] ), .A2(n13323), .B1(n26681), .B2(
        data_in[7]), .ZN(n13330) );
  INV_X1 U16659 ( .A(n13331), .ZN(n22506) );
  AOI22_X1 U16660 ( .A1(\mem[450][0] ), .A2(n13332), .B1(n26680), .B2(
        data_in[0]), .ZN(n13331) );
  INV_X1 U16661 ( .A(n13333), .ZN(n22505) );
  AOI22_X1 U16662 ( .A1(\mem[450][1] ), .A2(n13332), .B1(n26680), .B2(
        data_in[1]), .ZN(n13333) );
  INV_X1 U16663 ( .A(n13334), .ZN(n22504) );
  AOI22_X1 U16664 ( .A1(\mem[450][2] ), .A2(n13332), .B1(n26680), .B2(
        data_in[2]), .ZN(n13334) );
  INV_X1 U16665 ( .A(n13335), .ZN(n22503) );
  AOI22_X1 U16666 ( .A1(\mem[450][3] ), .A2(n13332), .B1(n26680), .B2(
        data_in[3]), .ZN(n13335) );
  INV_X1 U16667 ( .A(n13336), .ZN(n22502) );
  AOI22_X1 U16668 ( .A1(\mem[450][4] ), .A2(n13332), .B1(n26680), .B2(
        data_in[4]), .ZN(n13336) );
  INV_X1 U16669 ( .A(n13337), .ZN(n22501) );
  AOI22_X1 U16670 ( .A1(\mem[450][5] ), .A2(n13332), .B1(n26680), .B2(
        data_in[5]), .ZN(n13337) );
  INV_X1 U16671 ( .A(n13338), .ZN(n22500) );
  AOI22_X1 U16672 ( .A1(\mem[450][6] ), .A2(n13332), .B1(n26680), .B2(
        data_in[6]), .ZN(n13338) );
  INV_X1 U16673 ( .A(n13339), .ZN(n22499) );
  AOI22_X1 U16674 ( .A1(\mem[450][7] ), .A2(n13332), .B1(n26680), .B2(
        data_in[7]), .ZN(n13339) );
  INV_X1 U16675 ( .A(n13340), .ZN(n22498) );
  AOI22_X1 U16676 ( .A1(\mem[451][0] ), .A2(n13341), .B1(n26679), .B2(
        data_in[0]), .ZN(n13340) );
  INV_X1 U16677 ( .A(n13342), .ZN(n22497) );
  AOI22_X1 U16678 ( .A1(\mem[451][1] ), .A2(n13341), .B1(n26679), .B2(
        data_in[1]), .ZN(n13342) );
  INV_X1 U16679 ( .A(n13343), .ZN(n22496) );
  AOI22_X1 U16680 ( .A1(\mem[451][2] ), .A2(n13341), .B1(n26679), .B2(
        data_in[2]), .ZN(n13343) );
  INV_X1 U16681 ( .A(n13344), .ZN(n22495) );
  AOI22_X1 U16682 ( .A1(\mem[451][3] ), .A2(n13341), .B1(n26679), .B2(
        data_in[3]), .ZN(n13344) );
  INV_X1 U16683 ( .A(n13345), .ZN(n22494) );
  AOI22_X1 U16684 ( .A1(\mem[451][4] ), .A2(n13341), .B1(n26679), .B2(
        data_in[4]), .ZN(n13345) );
  INV_X1 U16685 ( .A(n13346), .ZN(n22493) );
  AOI22_X1 U16686 ( .A1(\mem[451][5] ), .A2(n13341), .B1(n26679), .B2(
        data_in[5]), .ZN(n13346) );
  INV_X1 U16687 ( .A(n13347), .ZN(n22492) );
  AOI22_X1 U16688 ( .A1(\mem[451][6] ), .A2(n13341), .B1(n26679), .B2(
        data_in[6]), .ZN(n13347) );
  INV_X1 U16689 ( .A(n13348), .ZN(n22491) );
  AOI22_X1 U16690 ( .A1(\mem[451][7] ), .A2(n13341), .B1(n26679), .B2(
        data_in[7]), .ZN(n13348) );
  INV_X1 U16691 ( .A(n13349), .ZN(n22490) );
  AOI22_X1 U16692 ( .A1(\mem[452][0] ), .A2(n13350), .B1(n26678), .B2(
        data_in[0]), .ZN(n13349) );
  INV_X1 U16693 ( .A(n13351), .ZN(n22489) );
  AOI22_X1 U16694 ( .A1(\mem[452][1] ), .A2(n13350), .B1(n26678), .B2(
        data_in[1]), .ZN(n13351) );
  INV_X1 U16695 ( .A(n13352), .ZN(n22488) );
  AOI22_X1 U16696 ( .A1(\mem[452][2] ), .A2(n13350), .B1(n26678), .B2(
        data_in[2]), .ZN(n13352) );
  INV_X1 U16697 ( .A(n13353), .ZN(n22487) );
  AOI22_X1 U16698 ( .A1(\mem[452][3] ), .A2(n13350), .B1(n26678), .B2(
        data_in[3]), .ZN(n13353) );
  INV_X1 U16699 ( .A(n13354), .ZN(n22486) );
  AOI22_X1 U16700 ( .A1(\mem[452][4] ), .A2(n13350), .B1(n26678), .B2(
        data_in[4]), .ZN(n13354) );
  INV_X1 U16701 ( .A(n13355), .ZN(n22485) );
  AOI22_X1 U16702 ( .A1(\mem[452][5] ), .A2(n13350), .B1(n26678), .B2(
        data_in[5]), .ZN(n13355) );
  INV_X1 U16703 ( .A(n13356), .ZN(n22484) );
  AOI22_X1 U16704 ( .A1(\mem[452][6] ), .A2(n13350), .B1(n26678), .B2(
        data_in[6]), .ZN(n13356) );
  INV_X1 U16705 ( .A(n13357), .ZN(n22483) );
  AOI22_X1 U16706 ( .A1(\mem[452][7] ), .A2(n13350), .B1(n26678), .B2(
        data_in[7]), .ZN(n13357) );
  INV_X1 U16707 ( .A(n13358), .ZN(n22482) );
  AOI22_X1 U16708 ( .A1(\mem[453][0] ), .A2(n13359), .B1(n26677), .B2(
        data_in[0]), .ZN(n13358) );
  INV_X1 U16709 ( .A(n13360), .ZN(n22481) );
  AOI22_X1 U16710 ( .A1(\mem[453][1] ), .A2(n13359), .B1(n26677), .B2(
        data_in[1]), .ZN(n13360) );
  INV_X1 U16711 ( .A(n13361), .ZN(n22480) );
  AOI22_X1 U16712 ( .A1(\mem[453][2] ), .A2(n13359), .B1(n26677), .B2(
        data_in[2]), .ZN(n13361) );
  INV_X1 U16713 ( .A(n13362), .ZN(n22479) );
  AOI22_X1 U16714 ( .A1(\mem[453][3] ), .A2(n13359), .B1(n26677), .B2(
        data_in[3]), .ZN(n13362) );
  INV_X1 U16715 ( .A(n13363), .ZN(n22478) );
  AOI22_X1 U16716 ( .A1(\mem[453][4] ), .A2(n13359), .B1(n26677), .B2(
        data_in[4]), .ZN(n13363) );
  INV_X1 U16717 ( .A(n13364), .ZN(n22477) );
  AOI22_X1 U16718 ( .A1(\mem[453][5] ), .A2(n13359), .B1(n26677), .B2(
        data_in[5]), .ZN(n13364) );
  INV_X1 U16719 ( .A(n13365), .ZN(n22476) );
  AOI22_X1 U16720 ( .A1(\mem[453][6] ), .A2(n13359), .B1(n26677), .B2(
        data_in[6]), .ZN(n13365) );
  INV_X1 U16721 ( .A(n13366), .ZN(n22475) );
  AOI22_X1 U16722 ( .A1(\mem[453][7] ), .A2(n13359), .B1(n26677), .B2(
        data_in[7]), .ZN(n13366) );
  INV_X1 U16723 ( .A(n13367), .ZN(n22474) );
  AOI22_X1 U16724 ( .A1(\mem[454][0] ), .A2(n13368), .B1(n26676), .B2(
        data_in[0]), .ZN(n13367) );
  INV_X1 U16725 ( .A(n13369), .ZN(n22473) );
  AOI22_X1 U16726 ( .A1(\mem[454][1] ), .A2(n13368), .B1(n26676), .B2(
        data_in[1]), .ZN(n13369) );
  INV_X1 U16727 ( .A(n13370), .ZN(n22472) );
  AOI22_X1 U16728 ( .A1(\mem[454][2] ), .A2(n13368), .B1(n26676), .B2(
        data_in[2]), .ZN(n13370) );
  INV_X1 U16729 ( .A(n13371), .ZN(n22471) );
  AOI22_X1 U16730 ( .A1(\mem[454][3] ), .A2(n13368), .B1(n26676), .B2(
        data_in[3]), .ZN(n13371) );
  INV_X1 U16731 ( .A(n13372), .ZN(n22470) );
  AOI22_X1 U16732 ( .A1(\mem[454][4] ), .A2(n13368), .B1(n26676), .B2(
        data_in[4]), .ZN(n13372) );
  INV_X1 U16733 ( .A(n13373), .ZN(n22469) );
  AOI22_X1 U16734 ( .A1(\mem[454][5] ), .A2(n13368), .B1(n26676), .B2(
        data_in[5]), .ZN(n13373) );
  INV_X1 U16735 ( .A(n13374), .ZN(n22468) );
  AOI22_X1 U16736 ( .A1(\mem[454][6] ), .A2(n13368), .B1(n26676), .B2(
        data_in[6]), .ZN(n13374) );
  INV_X1 U16737 ( .A(n13375), .ZN(n22467) );
  AOI22_X1 U16738 ( .A1(\mem[454][7] ), .A2(n13368), .B1(n26676), .B2(
        data_in[7]), .ZN(n13375) );
  INV_X1 U16739 ( .A(n13376), .ZN(n22466) );
  AOI22_X1 U16740 ( .A1(\mem[455][0] ), .A2(n13377), .B1(n26675), .B2(
        data_in[0]), .ZN(n13376) );
  INV_X1 U16741 ( .A(n13378), .ZN(n22465) );
  AOI22_X1 U16742 ( .A1(\mem[455][1] ), .A2(n13377), .B1(n26675), .B2(
        data_in[1]), .ZN(n13378) );
  INV_X1 U16743 ( .A(n13379), .ZN(n22464) );
  AOI22_X1 U16744 ( .A1(\mem[455][2] ), .A2(n13377), .B1(n26675), .B2(
        data_in[2]), .ZN(n13379) );
  INV_X1 U16745 ( .A(n13380), .ZN(n22463) );
  AOI22_X1 U16746 ( .A1(\mem[455][3] ), .A2(n13377), .B1(n26675), .B2(
        data_in[3]), .ZN(n13380) );
  INV_X1 U16747 ( .A(n13381), .ZN(n22462) );
  AOI22_X1 U16748 ( .A1(\mem[455][4] ), .A2(n13377), .B1(n26675), .B2(
        data_in[4]), .ZN(n13381) );
  INV_X1 U16749 ( .A(n13382), .ZN(n22461) );
  AOI22_X1 U16750 ( .A1(\mem[455][5] ), .A2(n13377), .B1(n26675), .B2(
        data_in[5]), .ZN(n13382) );
  INV_X1 U16751 ( .A(n13383), .ZN(n22460) );
  AOI22_X1 U16752 ( .A1(\mem[455][6] ), .A2(n13377), .B1(n26675), .B2(
        data_in[6]), .ZN(n13383) );
  INV_X1 U16753 ( .A(n13384), .ZN(n22459) );
  AOI22_X1 U16754 ( .A1(\mem[455][7] ), .A2(n13377), .B1(n26675), .B2(
        data_in[7]), .ZN(n13384) );
  INV_X1 U16755 ( .A(n13601), .ZN(n22266) );
  AOI22_X1 U16756 ( .A1(\mem[480][0] ), .A2(n13602), .B1(n26650), .B2(
        data_in[0]), .ZN(n13601) );
  INV_X1 U16757 ( .A(n13603), .ZN(n22265) );
  AOI22_X1 U16758 ( .A1(\mem[480][1] ), .A2(n13602), .B1(n26650), .B2(
        data_in[1]), .ZN(n13603) );
  INV_X1 U16759 ( .A(n13604), .ZN(n22264) );
  AOI22_X1 U16760 ( .A1(\mem[480][2] ), .A2(n13602), .B1(n26650), .B2(
        data_in[2]), .ZN(n13604) );
  INV_X1 U16761 ( .A(n13605), .ZN(n22263) );
  AOI22_X1 U16762 ( .A1(\mem[480][3] ), .A2(n13602), .B1(n26650), .B2(
        data_in[3]), .ZN(n13605) );
  INV_X1 U16763 ( .A(n13606), .ZN(n22262) );
  AOI22_X1 U16764 ( .A1(\mem[480][4] ), .A2(n13602), .B1(n26650), .B2(
        data_in[4]), .ZN(n13606) );
  INV_X1 U16765 ( .A(n13607), .ZN(n22261) );
  AOI22_X1 U16766 ( .A1(\mem[480][5] ), .A2(n13602), .B1(n26650), .B2(
        data_in[5]), .ZN(n13607) );
  INV_X1 U16767 ( .A(n13608), .ZN(n22260) );
  AOI22_X1 U16768 ( .A1(\mem[480][6] ), .A2(n13602), .B1(n26650), .B2(
        data_in[6]), .ZN(n13608) );
  INV_X1 U16769 ( .A(n13609), .ZN(n22259) );
  AOI22_X1 U16770 ( .A1(\mem[480][7] ), .A2(n13602), .B1(n26650), .B2(
        data_in[7]), .ZN(n13609) );
  INV_X1 U16771 ( .A(n13611), .ZN(n22258) );
  AOI22_X1 U16772 ( .A1(\mem[481][0] ), .A2(n13612), .B1(n26649), .B2(
        data_in[0]), .ZN(n13611) );
  INV_X1 U16773 ( .A(n13613), .ZN(n22257) );
  AOI22_X1 U16774 ( .A1(\mem[481][1] ), .A2(n13612), .B1(n26649), .B2(
        data_in[1]), .ZN(n13613) );
  INV_X1 U16775 ( .A(n13614), .ZN(n22256) );
  AOI22_X1 U16776 ( .A1(\mem[481][2] ), .A2(n13612), .B1(n26649), .B2(
        data_in[2]), .ZN(n13614) );
  INV_X1 U16777 ( .A(n13615), .ZN(n22255) );
  AOI22_X1 U16778 ( .A1(\mem[481][3] ), .A2(n13612), .B1(n26649), .B2(
        data_in[3]), .ZN(n13615) );
  INV_X1 U16779 ( .A(n13616), .ZN(n22254) );
  AOI22_X1 U16780 ( .A1(\mem[481][4] ), .A2(n13612), .B1(n26649), .B2(
        data_in[4]), .ZN(n13616) );
  INV_X1 U16781 ( .A(n13617), .ZN(n22253) );
  AOI22_X1 U16782 ( .A1(\mem[481][5] ), .A2(n13612), .B1(n26649), .B2(
        data_in[5]), .ZN(n13617) );
  INV_X1 U16783 ( .A(n13618), .ZN(n22252) );
  AOI22_X1 U16784 ( .A1(\mem[481][6] ), .A2(n13612), .B1(n26649), .B2(
        data_in[6]), .ZN(n13618) );
  INV_X1 U16785 ( .A(n13619), .ZN(n22251) );
  AOI22_X1 U16786 ( .A1(\mem[481][7] ), .A2(n13612), .B1(n26649), .B2(
        data_in[7]), .ZN(n13619) );
  INV_X1 U16787 ( .A(n13620), .ZN(n22250) );
  AOI22_X1 U16788 ( .A1(\mem[482][0] ), .A2(n13621), .B1(n26648), .B2(
        data_in[0]), .ZN(n13620) );
  INV_X1 U16789 ( .A(n13622), .ZN(n22249) );
  AOI22_X1 U16790 ( .A1(\mem[482][1] ), .A2(n13621), .B1(n26648), .B2(
        data_in[1]), .ZN(n13622) );
  INV_X1 U16791 ( .A(n13623), .ZN(n22248) );
  AOI22_X1 U16792 ( .A1(\mem[482][2] ), .A2(n13621), .B1(n26648), .B2(
        data_in[2]), .ZN(n13623) );
  INV_X1 U16793 ( .A(n13624), .ZN(n22247) );
  AOI22_X1 U16794 ( .A1(\mem[482][3] ), .A2(n13621), .B1(n26648), .B2(
        data_in[3]), .ZN(n13624) );
  INV_X1 U16795 ( .A(n13625), .ZN(n22246) );
  AOI22_X1 U16796 ( .A1(\mem[482][4] ), .A2(n13621), .B1(n26648), .B2(
        data_in[4]), .ZN(n13625) );
  INV_X1 U16797 ( .A(n13626), .ZN(n22245) );
  AOI22_X1 U16798 ( .A1(\mem[482][5] ), .A2(n13621), .B1(n26648), .B2(
        data_in[5]), .ZN(n13626) );
  INV_X1 U16799 ( .A(n13627), .ZN(n22244) );
  AOI22_X1 U16800 ( .A1(\mem[482][6] ), .A2(n13621), .B1(n26648), .B2(
        data_in[6]), .ZN(n13627) );
  INV_X1 U16801 ( .A(n13628), .ZN(n22243) );
  AOI22_X1 U16802 ( .A1(\mem[482][7] ), .A2(n13621), .B1(n26648), .B2(
        data_in[7]), .ZN(n13628) );
  INV_X1 U16803 ( .A(n13629), .ZN(n22242) );
  AOI22_X1 U16804 ( .A1(\mem[483][0] ), .A2(n13630), .B1(n26647), .B2(
        data_in[0]), .ZN(n13629) );
  INV_X1 U16805 ( .A(n13631), .ZN(n22241) );
  AOI22_X1 U16806 ( .A1(\mem[483][1] ), .A2(n13630), .B1(n26647), .B2(
        data_in[1]), .ZN(n13631) );
  INV_X1 U16807 ( .A(n13632), .ZN(n22240) );
  AOI22_X1 U16808 ( .A1(\mem[483][2] ), .A2(n13630), .B1(n26647), .B2(
        data_in[2]), .ZN(n13632) );
  INV_X1 U16809 ( .A(n13633), .ZN(n22239) );
  AOI22_X1 U16810 ( .A1(\mem[483][3] ), .A2(n13630), .B1(n26647), .B2(
        data_in[3]), .ZN(n13633) );
  INV_X1 U16811 ( .A(n13634), .ZN(n22238) );
  AOI22_X1 U16812 ( .A1(\mem[483][4] ), .A2(n13630), .B1(n26647), .B2(
        data_in[4]), .ZN(n13634) );
  INV_X1 U16813 ( .A(n13635), .ZN(n22237) );
  AOI22_X1 U16814 ( .A1(\mem[483][5] ), .A2(n13630), .B1(n26647), .B2(
        data_in[5]), .ZN(n13635) );
  INV_X1 U16815 ( .A(n13636), .ZN(n22236) );
  AOI22_X1 U16816 ( .A1(\mem[483][6] ), .A2(n13630), .B1(n26647), .B2(
        data_in[6]), .ZN(n13636) );
  INV_X1 U16817 ( .A(n13637), .ZN(n22235) );
  AOI22_X1 U16818 ( .A1(\mem[483][7] ), .A2(n13630), .B1(n26647), .B2(
        data_in[7]), .ZN(n13637) );
  INV_X1 U16819 ( .A(n13638), .ZN(n22234) );
  AOI22_X1 U16820 ( .A1(\mem[484][0] ), .A2(n13639), .B1(n26646), .B2(
        data_in[0]), .ZN(n13638) );
  INV_X1 U16821 ( .A(n13640), .ZN(n22233) );
  AOI22_X1 U16822 ( .A1(\mem[484][1] ), .A2(n13639), .B1(n26646), .B2(
        data_in[1]), .ZN(n13640) );
  INV_X1 U16823 ( .A(n13641), .ZN(n22232) );
  AOI22_X1 U16824 ( .A1(\mem[484][2] ), .A2(n13639), .B1(n26646), .B2(
        data_in[2]), .ZN(n13641) );
  INV_X1 U16825 ( .A(n13642), .ZN(n22231) );
  AOI22_X1 U16826 ( .A1(\mem[484][3] ), .A2(n13639), .B1(n26646), .B2(
        data_in[3]), .ZN(n13642) );
  INV_X1 U16827 ( .A(n13643), .ZN(n22230) );
  AOI22_X1 U16828 ( .A1(\mem[484][4] ), .A2(n13639), .B1(n26646), .B2(
        data_in[4]), .ZN(n13643) );
  INV_X1 U16829 ( .A(n13644), .ZN(n22229) );
  AOI22_X1 U16830 ( .A1(\mem[484][5] ), .A2(n13639), .B1(n26646), .B2(
        data_in[5]), .ZN(n13644) );
  INV_X1 U16831 ( .A(n13645), .ZN(n22228) );
  AOI22_X1 U16832 ( .A1(\mem[484][6] ), .A2(n13639), .B1(n26646), .B2(
        data_in[6]), .ZN(n13645) );
  INV_X1 U16833 ( .A(n13646), .ZN(n22227) );
  AOI22_X1 U16834 ( .A1(\mem[484][7] ), .A2(n13639), .B1(n26646), .B2(
        data_in[7]), .ZN(n13646) );
  INV_X1 U16835 ( .A(n13647), .ZN(n22226) );
  AOI22_X1 U16836 ( .A1(\mem[485][0] ), .A2(n13648), .B1(n26645), .B2(
        data_in[0]), .ZN(n13647) );
  INV_X1 U16837 ( .A(n13649), .ZN(n22225) );
  AOI22_X1 U16838 ( .A1(\mem[485][1] ), .A2(n13648), .B1(n26645), .B2(
        data_in[1]), .ZN(n13649) );
  INV_X1 U16839 ( .A(n13650), .ZN(n22224) );
  AOI22_X1 U16840 ( .A1(\mem[485][2] ), .A2(n13648), .B1(n26645), .B2(
        data_in[2]), .ZN(n13650) );
  INV_X1 U16841 ( .A(n13651), .ZN(n22223) );
  AOI22_X1 U16842 ( .A1(\mem[485][3] ), .A2(n13648), .B1(n26645), .B2(
        data_in[3]), .ZN(n13651) );
  INV_X1 U16843 ( .A(n13652), .ZN(n22222) );
  AOI22_X1 U16844 ( .A1(\mem[485][4] ), .A2(n13648), .B1(n26645), .B2(
        data_in[4]), .ZN(n13652) );
  INV_X1 U16845 ( .A(n13653), .ZN(n22221) );
  AOI22_X1 U16846 ( .A1(\mem[485][5] ), .A2(n13648), .B1(n26645), .B2(
        data_in[5]), .ZN(n13653) );
  INV_X1 U16847 ( .A(n13654), .ZN(n22220) );
  AOI22_X1 U16848 ( .A1(\mem[485][6] ), .A2(n13648), .B1(n26645), .B2(
        data_in[6]), .ZN(n13654) );
  INV_X1 U16849 ( .A(n13655), .ZN(n22219) );
  AOI22_X1 U16850 ( .A1(\mem[485][7] ), .A2(n13648), .B1(n26645), .B2(
        data_in[7]), .ZN(n13655) );
  INV_X1 U16851 ( .A(n13656), .ZN(n22218) );
  AOI22_X1 U16852 ( .A1(\mem[486][0] ), .A2(n13657), .B1(n26644), .B2(
        data_in[0]), .ZN(n13656) );
  INV_X1 U16853 ( .A(n13658), .ZN(n22217) );
  AOI22_X1 U16854 ( .A1(\mem[486][1] ), .A2(n13657), .B1(n26644), .B2(
        data_in[1]), .ZN(n13658) );
  INV_X1 U16855 ( .A(n13659), .ZN(n22216) );
  AOI22_X1 U16856 ( .A1(\mem[486][2] ), .A2(n13657), .B1(n26644), .B2(
        data_in[2]), .ZN(n13659) );
  INV_X1 U16857 ( .A(n13660), .ZN(n22215) );
  AOI22_X1 U16858 ( .A1(\mem[486][3] ), .A2(n13657), .B1(n26644), .B2(
        data_in[3]), .ZN(n13660) );
  INV_X1 U16859 ( .A(n13661), .ZN(n22214) );
  AOI22_X1 U16860 ( .A1(\mem[486][4] ), .A2(n13657), .B1(n26644), .B2(
        data_in[4]), .ZN(n13661) );
  INV_X1 U16861 ( .A(n13662), .ZN(n22213) );
  AOI22_X1 U16862 ( .A1(\mem[486][5] ), .A2(n13657), .B1(n26644), .B2(
        data_in[5]), .ZN(n13662) );
  INV_X1 U16863 ( .A(n13663), .ZN(n22212) );
  AOI22_X1 U16864 ( .A1(\mem[486][6] ), .A2(n13657), .B1(n26644), .B2(
        data_in[6]), .ZN(n13663) );
  INV_X1 U16865 ( .A(n13664), .ZN(n22211) );
  AOI22_X1 U16866 ( .A1(\mem[486][7] ), .A2(n13657), .B1(n26644), .B2(
        data_in[7]), .ZN(n13664) );
  INV_X1 U16867 ( .A(n13665), .ZN(n22210) );
  AOI22_X1 U16868 ( .A1(\mem[487][0] ), .A2(n13666), .B1(n26643), .B2(
        data_in[0]), .ZN(n13665) );
  INV_X1 U16869 ( .A(n13667), .ZN(n22209) );
  AOI22_X1 U16870 ( .A1(\mem[487][1] ), .A2(n13666), .B1(n26643), .B2(
        data_in[1]), .ZN(n13667) );
  INV_X1 U16871 ( .A(n13668), .ZN(n22208) );
  AOI22_X1 U16872 ( .A1(\mem[487][2] ), .A2(n13666), .B1(n26643), .B2(
        data_in[2]), .ZN(n13668) );
  INV_X1 U16873 ( .A(n13669), .ZN(n22207) );
  AOI22_X1 U16874 ( .A1(\mem[487][3] ), .A2(n13666), .B1(n26643), .B2(
        data_in[3]), .ZN(n13669) );
  INV_X1 U16875 ( .A(n13670), .ZN(n22206) );
  AOI22_X1 U16876 ( .A1(\mem[487][4] ), .A2(n13666), .B1(n26643), .B2(
        data_in[4]), .ZN(n13670) );
  INV_X1 U16877 ( .A(n13671), .ZN(n22205) );
  AOI22_X1 U16878 ( .A1(\mem[487][5] ), .A2(n13666), .B1(n26643), .B2(
        data_in[5]), .ZN(n13671) );
  INV_X1 U16879 ( .A(n13672), .ZN(n22204) );
  AOI22_X1 U16880 ( .A1(\mem[487][6] ), .A2(n13666), .B1(n26643), .B2(
        data_in[6]), .ZN(n13672) );
  INV_X1 U16881 ( .A(n13673), .ZN(n22203) );
  AOI22_X1 U16882 ( .A1(\mem[487][7] ), .A2(n13666), .B1(n26643), .B2(
        data_in[7]), .ZN(n13673) );
  INV_X1 U16883 ( .A(n13890), .ZN(n22010) );
  AOI22_X1 U16884 ( .A1(\mem[512][0] ), .A2(n13891), .B1(n26618), .B2(
        data_in[0]), .ZN(n13890) );
  INV_X1 U16885 ( .A(n13892), .ZN(n22009) );
  AOI22_X1 U16886 ( .A1(\mem[512][1] ), .A2(n13891), .B1(n26618), .B2(
        data_in[1]), .ZN(n13892) );
  INV_X1 U16887 ( .A(n13893), .ZN(n22008) );
  AOI22_X1 U16888 ( .A1(\mem[512][2] ), .A2(n13891), .B1(n26618), .B2(
        data_in[2]), .ZN(n13893) );
  INV_X1 U16889 ( .A(n13894), .ZN(n22007) );
  AOI22_X1 U16890 ( .A1(\mem[512][3] ), .A2(n13891), .B1(n26618), .B2(
        data_in[3]), .ZN(n13894) );
  INV_X1 U16891 ( .A(n13895), .ZN(n22006) );
  AOI22_X1 U16892 ( .A1(\mem[512][4] ), .A2(n13891), .B1(n26618), .B2(
        data_in[4]), .ZN(n13895) );
  INV_X1 U16893 ( .A(n13896), .ZN(n22005) );
  AOI22_X1 U16894 ( .A1(\mem[512][5] ), .A2(n13891), .B1(n26618), .B2(
        data_in[5]), .ZN(n13896) );
  INV_X1 U16895 ( .A(n13897), .ZN(n22004) );
  AOI22_X1 U16896 ( .A1(\mem[512][6] ), .A2(n13891), .B1(n26618), .B2(
        data_in[6]), .ZN(n13897) );
  INV_X1 U16897 ( .A(n13898), .ZN(n22003) );
  AOI22_X1 U16898 ( .A1(\mem[512][7] ), .A2(n13891), .B1(n26618), .B2(
        data_in[7]), .ZN(n13898) );
  INV_X1 U16899 ( .A(n13900), .ZN(n22002) );
  AOI22_X1 U16900 ( .A1(\mem[513][0] ), .A2(n13901), .B1(n26617), .B2(
        data_in[0]), .ZN(n13900) );
  INV_X1 U16901 ( .A(n13902), .ZN(n22001) );
  AOI22_X1 U16902 ( .A1(\mem[513][1] ), .A2(n13901), .B1(n26617), .B2(
        data_in[1]), .ZN(n13902) );
  INV_X1 U16903 ( .A(n13903), .ZN(n22000) );
  AOI22_X1 U16904 ( .A1(\mem[513][2] ), .A2(n13901), .B1(n26617), .B2(
        data_in[2]), .ZN(n13903) );
  INV_X1 U16905 ( .A(n13904), .ZN(n21999) );
  AOI22_X1 U16906 ( .A1(\mem[513][3] ), .A2(n13901), .B1(n26617), .B2(
        data_in[3]), .ZN(n13904) );
  INV_X1 U16907 ( .A(n13905), .ZN(n21998) );
  AOI22_X1 U16908 ( .A1(\mem[513][4] ), .A2(n13901), .B1(n26617), .B2(
        data_in[4]), .ZN(n13905) );
  INV_X1 U16909 ( .A(n13906), .ZN(n21997) );
  AOI22_X1 U16910 ( .A1(\mem[513][5] ), .A2(n13901), .B1(n26617), .B2(
        data_in[5]), .ZN(n13906) );
  INV_X1 U16911 ( .A(n13907), .ZN(n21996) );
  AOI22_X1 U16912 ( .A1(\mem[513][6] ), .A2(n13901), .B1(n26617), .B2(
        data_in[6]), .ZN(n13907) );
  INV_X1 U16913 ( .A(n13908), .ZN(n21995) );
  AOI22_X1 U16914 ( .A1(\mem[513][7] ), .A2(n13901), .B1(n26617), .B2(
        data_in[7]), .ZN(n13908) );
  INV_X1 U16915 ( .A(n13909), .ZN(n21994) );
  AOI22_X1 U16916 ( .A1(\mem[514][0] ), .A2(n13910), .B1(n26616), .B2(
        data_in[0]), .ZN(n13909) );
  INV_X1 U16917 ( .A(n13911), .ZN(n21993) );
  AOI22_X1 U16918 ( .A1(\mem[514][1] ), .A2(n13910), .B1(n26616), .B2(
        data_in[1]), .ZN(n13911) );
  INV_X1 U16919 ( .A(n13912), .ZN(n21992) );
  AOI22_X1 U16920 ( .A1(\mem[514][2] ), .A2(n13910), .B1(n26616), .B2(
        data_in[2]), .ZN(n13912) );
  INV_X1 U16921 ( .A(n13913), .ZN(n21991) );
  AOI22_X1 U16922 ( .A1(\mem[514][3] ), .A2(n13910), .B1(n26616), .B2(
        data_in[3]), .ZN(n13913) );
  INV_X1 U16923 ( .A(n13914), .ZN(n21990) );
  AOI22_X1 U16924 ( .A1(\mem[514][4] ), .A2(n13910), .B1(n26616), .B2(
        data_in[4]), .ZN(n13914) );
  INV_X1 U16925 ( .A(n13915), .ZN(n21989) );
  AOI22_X1 U16926 ( .A1(\mem[514][5] ), .A2(n13910), .B1(n26616), .B2(
        data_in[5]), .ZN(n13915) );
  INV_X1 U16927 ( .A(n13916), .ZN(n21988) );
  AOI22_X1 U16928 ( .A1(\mem[514][6] ), .A2(n13910), .B1(n26616), .B2(
        data_in[6]), .ZN(n13916) );
  INV_X1 U16929 ( .A(n13917), .ZN(n21987) );
  AOI22_X1 U16930 ( .A1(\mem[514][7] ), .A2(n13910), .B1(n26616), .B2(
        data_in[7]), .ZN(n13917) );
  INV_X1 U16931 ( .A(n13918), .ZN(n21986) );
  AOI22_X1 U16932 ( .A1(\mem[515][0] ), .A2(n13919), .B1(n26615), .B2(
        data_in[0]), .ZN(n13918) );
  INV_X1 U16933 ( .A(n13920), .ZN(n21985) );
  AOI22_X1 U16934 ( .A1(\mem[515][1] ), .A2(n13919), .B1(n26615), .B2(
        data_in[1]), .ZN(n13920) );
  INV_X1 U16935 ( .A(n13921), .ZN(n21984) );
  AOI22_X1 U16936 ( .A1(\mem[515][2] ), .A2(n13919), .B1(n26615), .B2(
        data_in[2]), .ZN(n13921) );
  INV_X1 U16937 ( .A(n13922), .ZN(n21983) );
  AOI22_X1 U16938 ( .A1(\mem[515][3] ), .A2(n13919), .B1(n26615), .B2(
        data_in[3]), .ZN(n13922) );
  INV_X1 U16939 ( .A(n13923), .ZN(n21982) );
  AOI22_X1 U16940 ( .A1(\mem[515][4] ), .A2(n13919), .B1(n26615), .B2(
        data_in[4]), .ZN(n13923) );
  INV_X1 U16941 ( .A(n13924), .ZN(n21981) );
  AOI22_X1 U16942 ( .A1(\mem[515][5] ), .A2(n13919), .B1(n26615), .B2(
        data_in[5]), .ZN(n13924) );
  INV_X1 U16943 ( .A(n13925), .ZN(n21980) );
  AOI22_X1 U16944 ( .A1(\mem[515][6] ), .A2(n13919), .B1(n26615), .B2(
        data_in[6]), .ZN(n13925) );
  INV_X1 U16945 ( .A(n13926), .ZN(n21979) );
  AOI22_X1 U16946 ( .A1(\mem[515][7] ), .A2(n13919), .B1(n26615), .B2(
        data_in[7]), .ZN(n13926) );
  INV_X1 U16947 ( .A(n13927), .ZN(n21978) );
  AOI22_X1 U16948 ( .A1(\mem[516][0] ), .A2(n13928), .B1(n26614), .B2(
        data_in[0]), .ZN(n13927) );
  INV_X1 U16949 ( .A(n13929), .ZN(n21977) );
  AOI22_X1 U16950 ( .A1(\mem[516][1] ), .A2(n13928), .B1(n26614), .B2(
        data_in[1]), .ZN(n13929) );
  INV_X1 U16951 ( .A(n13930), .ZN(n21976) );
  AOI22_X1 U16952 ( .A1(\mem[516][2] ), .A2(n13928), .B1(n26614), .B2(
        data_in[2]), .ZN(n13930) );
  INV_X1 U16953 ( .A(n13931), .ZN(n21975) );
  AOI22_X1 U16954 ( .A1(\mem[516][3] ), .A2(n13928), .B1(n26614), .B2(
        data_in[3]), .ZN(n13931) );
  INV_X1 U16955 ( .A(n13932), .ZN(n21974) );
  AOI22_X1 U16956 ( .A1(\mem[516][4] ), .A2(n13928), .B1(n26614), .B2(
        data_in[4]), .ZN(n13932) );
  INV_X1 U16957 ( .A(n13933), .ZN(n21973) );
  AOI22_X1 U16958 ( .A1(\mem[516][5] ), .A2(n13928), .B1(n26614), .B2(
        data_in[5]), .ZN(n13933) );
  INV_X1 U16959 ( .A(n13934), .ZN(n21972) );
  AOI22_X1 U16960 ( .A1(\mem[516][6] ), .A2(n13928), .B1(n26614), .B2(
        data_in[6]), .ZN(n13934) );
  INV_X1 U16961 ( .A(n13935), .ZN(n21971) );
  AOI22_X1 U16962 ( .A1(\mem[516][7] ), .A2(n13928), .B1(n26614), .B2(
        data_in[7]), .ZN(n13935) );
  INV_X1 U16963 ( .A(n13936), .ZN(n21970) );
  AOI22_X1 U16964 ( .A1(\mem[517][0] ), .A2(n13937), .B1(n26613), .B2(
        data_in[0]), .ZN(n13936) );
  INV_X1 U16965 ( .A(n13938), .ZN(n21969) );
  AOI22_X1 U16966 ( .A1(\mem[517][1] ), .A2(n13937), .B1(n26613), .B2(
        data_in[1]), .ZN(n13938) );
  INV_X1 U16967 ( .A(n13939), .ZN(n21968) );
  AOI22_X1 U16968 ( .A1(\mem[517][2] ), .A2(n13937), .B1(n26613), .B2(
        data_in[2]), .ZN(n13939) );
  INV_X1 U16969 ( .A(n13940), .ZN(n21967) );
  AOI22_X1 U16970 ( .A1(\mem[517][3] ), .A2(n13937), .B1(n26613), .B2(
        data_in[3]), .ZN(n13940) );
  INV_X1 U16971 ( .A(n13941), .ZN(n21966) );
  AOI22_X1 U16972 ( .A1(\mem[517][4] ), .A2(n13937), .B1(n26613), .B2(
        data_in[4]), .ZN(n13941) );
  INV_X1 U16973 ( .A(n13942), .ZN(n21965) );
  AOI22_X1 U16974 ( .A1(\mem[517][5] ), .A2(n13937), .B1(n26613), .B2(
        data_in[5]), .ZN(n13942) );
  INV_X1 U16975 ( .A(n13943), .ZN(n21964) );
  AOI22_X1 U16976 ( .A1(\mem[517][6] ), .A2(n13937), .B1(n26613), .B2(
        data_in[6]), .ZN(n13943) );
  INV_X1 U16977 ( .A(n13944), .ZN(n21963) );
  AOI22_X1 U16978 ( .A1(\mem[517][7] ), .A2(n13937), .B1(n26613), .B2(
        data_in[7]), .ZN(n13944) );
  INV_X1 U16979 ( .A(n13945), .ZN(n21962) );
  AOI22_X1 U16980 ( .A1(\mem[518][0] ), .A2(n13946), .B1(n26612), .B2(
        data_in[0]), .ZN(n13945) );
  INV_X1 U16981 ( .A(n13947), .ZN(n21961) );
  AOI22_X1 U16982 ( .A1(\mem[518][1] ), .A2(n13946), .B1(n26612), .B2(
        data_in[1]), .ZN(n13947) );
  INV_X1 U16983 ( .A(n13948), .ZN(n21960) );
  AOI22_X1 U16984 ( .A1(\mem[518][2] ), .A2(n13946), .B1(n26612), .B2(
        data_in[2]), .ZN(n13948) );
  INV_X1 U16985 ( .A(n13949), .ZN(n21959) );
  AOI22_X1 U16986 ( .A1(\mem[518][3] ), .A2(n13946), .B1(n26612), .B2(
        data_in[3]), .ZN(n13949) );
  INV_X1 U16987 ( .A(n13950), .ZN(n21958) );
  AOI22_X1 U16988 ( .A1(\mem[518][4] ), .A2(n13946), .B1(n26612), .B2(
        data_in[4]), .ZN(n13950) );
  INV_X1 U16989 ( .A(n13951), .ZN(n21957) );
  AOI22_X1 U16990 ( .A1(\mem[518][5] ), .A2(n13946), .B1(n26612), .B2(
        data_in[5]), .ZN(n13951) );
  INV_X1 U16991 ( .A(n13952), .ZN(n21956) );
  AOI22_X1 U16992 ( .A1(\mem[518][6] ), .A2(n13946), .B1(n26612), .B2(
        data_in[6]), .ZN(n13952) );
  INV_X1 U16993 ( .A(n13953), .ZN(n21955) );
  AOI22_X1 U16994 ( .A1(\mem[518][7] ), .A2(n13946), .B1(n26612), .B2(
        data_in[7]), .ZN(n13953) );
  INV_X1 U16995 ( .A(n13954), .ZN(n21954) );
  AOI22_X1 U16996 ( .A1(\mem[519][0] ), .A2(n13955), .B1(n26611), .B2(
        data_in[0]), .ZN(n13954) );
  INV_X1 U16997 ( .A(n13956), .ZN(n21953) );
  AOI22_X1 U16998 ( .A1(\mem[519][1] ), .A2(n13955), .B1(n26611), .B2(
        data_in[1]), .ZN(n13956) );
  INV_X1 U16999 ( .A(n13957), .ZN(n21952) );
  AOI22_X1 U17000 ( .A1(\mem[519][2] ), .A2(n13955), .B1(n26611), .B2(
        data_in[2]), .ZN(n13957) );
  INV_X1 U17001 ( .A(n13958), .ZN(n21951) );
  AOI22_X1 U17002 ( .A1(\mem[519][3] ), .A2(n13955), .B1(n26611), .B2(
        data_in[3]), .ZN(n13958) );
  INV_X1 U17003 ( .A(n13959), .ZN(n21950) );
  AOI22_X1 U17004 ( .A1(\mem[519][4] ), .A2(n13955), .B1(n26611), .B2(
        data_in[4]), .ZN(n13959) );
  INV_X1 U17005 ( .A(n13960), .ZN(n21949) );
  AOI22_X1 U17006 ( .A1(\mem[519][5] ), .A2(n13955), .B1(n26611), .B2(
        data_in[5]), .ZN(n13960) );
  INV_X1 U17007 ( .A(n13961), .ZN(n21948) );
  AOI22_X1 U17008 ( .A1(\mem[519][6] ), .A2(n13955), .B1(n26611), .B2(
        data_in[6]), .ZN(n13961) );
  INV_X1 U17009 ( .A(n13962), .ZN(n21947) );
  AOI22_X1 U17010 ( .A1(\mem[519][7] ), .A2(n13955), .B1(n26611), .B2(
        data_in[7]), .ZN(n13962) );
  INV_X1 U17011 ( .A(n14180), .ZN(n21754) );
  AOI22_X1 U17012 ( .A1(\mem[544][0] ), .A2(n14181), .B1(n26586), .B2(
        data_in[0]), .ZN(n14180) );
  INV_X1 U17013 ( .A(n14182), .ZN(n21753) );
  AOI22_X1 U17014 ( .A1(\mem[544][1] ), .A2(n14181), .B1(n26586), .B2(
        data_in[1]), .ZN(n14182) );
  INV_X1 U17015 ( .A(n14183), .ZN(n21752) );
  AOI22_X1 U17016 ( .A1(\mem[544][2] ), .A2(n14181), .B1(n26586), .B2(
        data_in[2]), .ZN(n14183) );
  INV_X1 U17017 ( .A(n14184), .ZN(n21751) );
  AOI22_X1 U17018 ( .A1(\mem[544][3] ), .A2(n14181), .B1(n26586), .B2(
        data_in[3]), .ZN(n14184) );
  INV_X1 U17019 ( .A(n14185), .ZN(n21750) );
  AOI22_X1 U17020 ( .A1(\mem[544][4] ), .A2(n14181), .B1(n26586), .B2(
        data_in[4]), .ZN(n14185) );
  INV_X1 U17021 ( .A(n14186), .ZN(n21749) );
  AOI22_X1 U17022 ( .A1(\mem[544][5] ), .A2(n14181), .B1(n26586), .B2(
        data_in[5]), .ZN(n14186) );
  INV_X1 U17023 ( .A(n14187), .ZN(n21748) );
  AOI22_X1 U17024 ( .A1(\mem[544][6] ), .A2(n14181), .B1(n26586), .B2(
        data_in[6]), .ZN(n14187) );
  INV_X1 U17025 ( .A(n14188), .ZN(n21747) );
  AOI22_X1 U17026 ( .A1(\mem[544][7] ), .A2(n14181), .B1(n26586), .B2(
        data_in[7]), .ZN(n14188) );
  INV_X1 U17027 ( .A(n14190), .ZN(n21746) );
  AOI22_X1 U17028 ( .A1(\mem[545][0] ), .A2(n14191), .B1(n26585), .B2(
        data_in[0]), .ZN(n14190) );
  INV_X1 U17029 ( .A(n14192), .ZN(n21745) );
  AOI22_X1 U17030 ( .A1(\mem[545][1] ), .A2(n14191), .B1(n26585), .B2(
        data_in[1]), .ZN(n14192) );
  INV_X1 U17031 ( .A(n14193), .ZN(n21744) );
  AOI22_X1 U17032 ( .A1(\mem[545][2] ), .A2(n14191), .B1(n26585), .B2(
        data_in[2]), .ZN(n14193) );
  INV_X1 U17033 ( .A(n14194), .ZN(n21743) );
  AOI22_X1 U17034 ( .A1(\mem[545][3] ), .A2(n14191), .B1(n26585), .B2(
        data_in[3]), .ZN(n14194) );
  INV_X1 U17035 ( .A(n14195), .ZN(n21742) );
  AOI22_X1 U17036 ( .A1(\mem[545][4] ), .A2(n14191), .B1(n26585), .B2(
        data_in[4]), .ZN(n14195) );
  INV_X1 U17037 ( .A(n14196), .ZN(n21741) );
  AOI22_X1 U17038 ( .A1(\mem[545][5] ), .A2(n14191), .B1(n26585), .B2(
        data_in[5]), .ZN(n14196) );
  INV_X1 U17039 ( .A(n14197), .ZN(n21740) );
  AOI22_X1 U17040 ( .A1(\mem[545][6] ), .A2(n14191), .B1(n26585), .B2(
        data_in[6]), .ZN(n14197) );
  INV_X1 U17041 ( .A(n14198), .ZN(n21739) );
  AOI22_X1 U17042 ( .A1(\mem[545][7] ), .A2(n14191), .B1(n26585), .B2(
        data_in[7]), .ZN(n14198) );
  INV_X1 U17043 ( .A(n14199), .ZN(n21738) );
  AOI22_X1 U17044 ( .A1(\mem[546][0] ), .A2(n14200), .B1(n26584), .B2(
        data_in[0]), .ZN(n14199) );
  INV_X1 U17045 ( .A(n14201), .ZN(n21737) );
  AOI22_X1 U17046 ( .A1(\mem[546][1] ), .A2(n14200), .B1(n26584), .B2(
        data_in[1]), .ZN(n14201) );
  INV_X1 U17047 ( .A(n14202), .ZN(n21736) );
  AOI22_X1 U17048 ( .A1(\mem[546][2] ), .A2(n14200), .B1(n26584), .B2(
        data_in[2]), .ZN(n14202) );
  INV_X1 U17049 ( .A(n14203), .ZN(n21735) );
  AOI22_X1 U17050 ( .A1(\mem[546][3] ), .A2(n14200), .B1(n26584), .B2(
        data_in[3]), .ZN(n14203) );
  INV_X1 U17051 ( .A(n14204), .ZN(n21734) );
  AOI22_X1 U17052 ( .A1(\mem[546][4] ), .A2(n14200), .B1(n26584), .B2(
        data_in[4]), .ZN(n14204) );
  INV_X1 U17053 ( .A(n14205), .ZN(n21733) );
  AOI22_X1 U17054 ( .A1(\mem[546][5] ), .A2(n14200), .B1(n26584), .B2(
        data_in[5]), .ZN(n14205) );
  INV_X1 U17055 ( .A(n14206), .ZN(n21732) );
  AOI22_X1 U17056 ( .A1(\mem[546][6] ), .A2(n14200), .B1(n26584), .B2(
        data_in[6]), .ZN(n14206) );
  INV_X1 U17057 ( .A(n14207), .ZN(n21731) );
  AOI22_X1 U17058 ( .A1(\mem[546][7] ), .A2(n14200), .B1(n26584), .B2(
        data_in[7]), .ZN(n14207) );
  INV_X1 U17059 ( .A(n14208), .ZN(n21730) );
  AOI22_X1 U17060 ( .A1(\mem[547][0] ), .A2(n14209), .B1(n26583), .B2(
        data_in[0]), .ZN(n14208) );
  INV_X1 U17061 ( .A(n14210), .ZN(n21729) );
  AOI22_X1 U17062 ( .A1(\mem[547][1] ), .A2(n14209), .B1(n26583), .B2(
        data_in[1]), .ZN(n14210) );
  INV_X1 U17063 ( .A(n14211), .ZN(n21728) );
  AOI22_X1 U17064 ( .A1(\mem[547][2] ), .A2(n14209), .B1(n26583), .B2(
        data_in[2]), .ZN(n14211) );
  INV_X1 U17065 ( .A(n14212), .ZN(n21727) );
  AOI22_X1 U17066 ( .A1(\mem[547][3] ), .A2(n14209), .B1(n26583), .B2(
        data_in[3]), .ZN(n14212) );
  INV_X1 U17067 ( .A(n14213), .ZN(n21726) );
  AOI22_X1 U17068 ( .A1(\mem[547][4] ), .A2(n14209), .B1(n26583), .B2(
        data_in[4]), .ZN(n14213) );
  INV_X1 U17069 ( .A(n14214), .ZN(n21725) );
  AOI22_X1 U17070 ( .A1(\mem[547][5] ), .A2(n14209), .B1(n26583), .B2(
        data_in[5]), .ZN(n14214) );
  INV_X1 U17071 ( .A(n14215), .ZN(n21724) );
  AOI22_X1 U17072 ( .A1(\mem[547][6] ), .A2(n14209), .B1(n26583), .B2(
        data_in[6]), .ZN(n14215) );
  INV_X1 U17073 ( .A(n14216), .ZN(n21723) );
  AOI22_X1 U17074 ( .A1(\mem[547][7] ), .A2(n14209), .B1(n26583), .B2(
        data_in[7]), .ZN(n14216) );
  INV_X1 U17075 ( .A(n14217), .ZN(n21722) );
  AOI22_X1 U17076 ( .A1(\mem[548][0] ), .A2(n14218), .B1(n26582), .B2(
        data_in[0]), .ZN(n14217) );
  INV_X1 U17077 ( .A(n14219), .ZN(n21721) );
  AOI22_X1 U17078 ( .A1(\mem[548][1] ), .A2(n14218), .B1(n26582), .B2(
        data_in[1]), .ZN(n14219) );
  INV_X1 U17079 ( .A(n14220), .ZN(n21720) );
  AOI22_X1 U17080 ( .A1(\mem[548][2] ), .A2(n14218), .B1(n26582), .B2(
        data_in[2]), .ZN(n14220) );
  INV_X1 U17081 ( .A(n14221), .ZN(n21719) );
  AOI22_X1 U17082 ( .A1(\mem[548][3] ), .A2(n14218), .B1(n26582), .B2(
        data_in[3]), .ZN(n14221) );
  INV_X1 U17083 ( .A(n14222), .ZN(n21718) );
  AOI22_X1 U17084 ( .A1(\mem[548][4] ), .A2(n14218), .B1(n26582), .B2(
        data_in[4]), .ZN(n14222) );
  INV_X1 U17085 ( .A(n14223), .ZN(n21717) );
  AOI22_X1 U17086 ( .A1(\mem[548][5] ), .A2(n14218), .B1(n26582), .B2(
        data_in[5]), .ZN(n14223) );
  INV_X1 U17087 ( .A(n14224), .ZN(n21716) );
  AOI22_X1 U17088 ( .A1(\mem[548][6] ), .A2(n14218), .B1(n26582), .B2(
        data_in[6]), .ZN(n14224) );
  INV_X1 U17089 ( .A(n14225), .ZN(n21715) );
  AOI22_X1 U17090 ( .A1(\mem[548][7] ), .A2(n14218), .B1(n26582), .B2(
        data_in[7]), .ZN(n14225) );
  INV_X1 U17091 ( .A(n14226), .ZN(n21714) );
  AOI22_X1 U17092 ( .A1(\mem[549][0] ), .A2(n14227), .B1(n26581), .B2(
        data_in[0]), .ZN(n14226) );
  INV_X1 U17093 ( .A(n14228), .ZN(n21713) );
  AOI22_X1 U17094 ( .A1(\mem[549][1] ), .A2(n14227), .B1(n26581), .B2(
        data_in[1]), .ZN(n14228) );
  INV_X1 U17095 ( .A(n14229), .ZN(n21712) );
  AOI22_X1 U17096 ( .A1(\mem[549][2] ), .A2(n14227), .B1(n26581), .B2(
        data_in[2]), .ZN(n14229) );
  INV_X1 U17097 ( .A(n14230), .ZN(n21711) );
  AOI22_X1 U17098 ( .A1(\mem[549][3] ), .A2(n14227), .B1(n26581), .B2(
        data_in[3]), .ZN(n14230) );
  INV_X1 U17099 ( .A(n14231), .ZN(n21710) );
  AOI22_X1 U17100 ( .A1(\mem[549][4] ), .A2(n14227), .B1(n26581), .B2(
        data_in[4]), .ZN(n14231) );
  INV_X1 U17101 ( .A(n14232), .ZN(n21709) );
  AOI22_X1 U17102 ( .A1(\mem[549][5] ), .A2(n14227), .B1(n26581), .B2(
        data_in[5]), .ZN(n14232) );
  INV_X1 U17103 ( .A(n14233), .ZN(n21708) );
  AOI22_X1 U17104 ( .A1(\mem[549][6] ), .A2(n14227), .B1(n26581), .B2(
        data_in[6]), .ZN(n14233) );
  INV_X1 U17105 ( .A(n14234), .ZN(n21707) );
  AOI22_X1 U17106 ( .A1(\mem[549][7] ), .A2(n14227), .B1(n26581), .B2(
        data_in[7]), .ZN(n14234) );
  INV_X1 U17107 ( .A(n14235), .ZN(n21706) );
  AOI22_X1 U17108 ( .A1(\mem[550][0] ), .A2(n14236), .B1(n26580), .B2(
        data_in[0]), .ZN(n14235) );
  INV_X1 U17109 ( .A(n14237), .ZN(n21705) );
  AOI22_X1 U17110 ( .A1(\mem[550][1] ), .A2(n14236), .B1(n26580), .B2(
        data_in[1]), .ZN(n14237) );
  INV_X1 U17111 ( .A(n14238), .ZN(n21704) );
  AOI22_X1 U17112 ( .A1(\mem[550][2] ), .A2(n14236), .B1(n26580), .B2(
        data_in[2]), .ZN(n14238) );
  INV_X1 U17113 ( .A(n14239), .ZN(n21703) );
  AOI22_X1 U17114 ( .A1(\mem[550][3] ), .A2(n14236), .B1(n26580), .B2(
        data_in[3]), .ZN(n14239) );
  INV_X1 U17115 ( .A(n14240), .ZN(n21702) );
  AOI22_X1 U17116 ( .A1(\mem[550][4] ), .A2(n14236), .B1(n26580), .B2(
        data_in[4]), .ZN(n14240) );
  INV_X1 U17117 ( .A(n14241), .ZN(n21701) );
  AOI22_X1 U17118 ( .A1(\mem[550][5] ), .A2(n14236), .B1(n26580), .B2(
        data_in[5]), .ZN(n14241) );
  INV_X1 U17119 ( .A(n14242), .ZN(n21700) );
  AOI22_X1 U17120 ( .A1(\mem[550][6] ), .A2(n14236), .B1(n26580), .B2(
        data_in[6]), .ZN(n14242) );
  INV_X1 U17121 ( .A(n14243), .ZN(n21699) );
  AOI22_X1 U17122 ( .A1(\mem[550][7] ), .A2(n14236), .B1(n26580), .B2(
        data_in[7]), .ZN(n14243) );
  INV_X1 U17123 ( .A(n14244), .ZN(n21698) );
  AOI22_X1 U17124 ( .A1(\mem[551][0] ), .A2(n14245), .B1(n26579), .B2(
        data_in[0]), .ZN(n14244) );
  INV_X1 U17125 ( .A(n14246), .ZN(n21697) );
  AOI22_X1 U17126 ( .A1(\mem[551][1] ), .A2(n14245), .B1(n26579), .B2(
        data_in[1]), .ZN(n14246) );
  INV_X1 U17127 ( .A(n14247), .ZN(n21696) );
  AOI22_X1 U17128 ( .A1(\mem[551][2] ), .A2(n14245), .B1(n26579), .B2(
        data_in[2]), .ZN(n14247) );
  INV_X1 U17129 ( .A(n14248), .ZN(n21695) );
  AOI22_X1 U17130 ( .A1(\mem[551][3] ), .A2(n14245), .B1(n26579), .B2(
        data_in[3]), .ZN(n14248) );
  INV_X1 U17131 ( .A(n14249), .ZN(n21694) );
  AOI22_X1 U17132 ( .A1(\mem[551][4] ), .A2(n14245), .B1(n26579), .B2(
        data_in[4]), .ZN(n14249) );
  INV_X1 U17133 ( .A(n14250), .ZN(n21693) );
  AOI22_X1 U17134 ( .A1(\mem[551][5] ), .A2(n14245), .B1(n26579), .B2(
        data_in[5]), .ZN(n14250) );
  INV_X1 U17135 ( .A(n14251), .ZN(n21692) );
  AOI22_X1 U17136 ( .A1(\mem[551][6] ), .A2(n14245), .B1(n26579), .B2(
        data_in[6]), .ZN(n14251) );
  INV_X1 U17137 ( .A(n14252), .ZN(n21691) );
  AOI22_X1 U17138 ( .A1(\mem[551][7] ), .A2(n14245), .B1(n26579), .B2(
        data_in[7]), .ZN(n14252) );
  INV_X1 U17139 ( .A(n14469), .ZN(n21498) );
  AOI22_X1 U17140 ( .A1(\mem[576][0] ), .A2(n14470), .B1(n26554), .B2(
        data_in[0]), .ZN(n14469) );
  INV_X1 U17141 ( .A(n14471), .ZN(n21497) );
  AOI22_X1 U17142 ( .A1(\mem[576][1] ), .A2(n14470), .B1(n26554), .B2(
        data_in[1]), .ZN(n14471) );
  INV_X1 U17143 ( .A(n14472), .ZN(n21496) );
  AOI22_X1 U17144 ( .A1(\mem[576][2] ), .A2(n14470), .B1(n26554), .B2(
        data_in[2]), .ZN(n14472) );
  INV_X1 U17145 ( .A(n14473), .ZN(n21495) );
  AOI22_X1 U17146 ( .A1(\mem[576][3] ), .A2(n14470), .B1(n26554), .B2(
        data_in[3]), .ZN(n14473) );
  INV_X1 U17147 ( .A(n14474), .ZN(n21494) );
  AOI22_X1 U17148 ( .A1(\mem[576][4] ), .A2(n14470), .B1(n26554), .B2(
        data_in[4]), .ZN(n14474) );
  INV_X1 U17149 ( .A(n14475), .ZN(n21493) );
  AOI22_X1 U17150 ( .A1(\mem[576][5] ), .A2(n14470), .B1(n26554), .B2(
        data_in[5]), .ZN(n14475) );
  INV_X1 U17151 ( .A(n14476), .ZN(n21492) );
  AOI22_X1 U17152 ( .A1(\mem[576][6] ), .A2(n14470), .B1(n26554), .B2(
        data_in[6]), .ZN(n14476) );
  INV_X1 U17153 ( .A(n14477), .ZN(n21491) );
  AOI22_X1 U17154 ( .A1(\mem[576][7] ), .A2(n14470), .B1(n26554), .B2(
        data_in[7]), .ZN(n14477) );
  INV_X1 U17155 ( .A(n14479), .ZN(n21490) );
  AOI22_X1 U17156 ( .A1(\mem[577][0] ), .A2(n14480), .B1(n26553), .B2(
        data_in[0]), .ZN(n14479) );
  INV_X1 U17157 ( .A(n14481), .ZN(n21489) );
  AOI22_X1 U17158 ( .A1(\mem[577][1] ), .A2(n14480), .B1(n26553), .B2(
        data_in[1]), .ZN(n14481) );
  INV_X1 U17159 ( .A(n14482), .ZN(n21488) );
  AOI22_X1 U17160 ( .A1(\mem[577][2] ), .A2(n14480), .B1(n26553), .B2(
        data_in[2]), .ZN(n14482) );
  INV_X1 U17161 ( .A(n14483), .ZN(n21487) );
  AOI22_X1 U17162 ( .A1(\mem[577][3] ), .A2(n14480), .B1(n26553), .B2(
        data_in[3]), .ZN(n14483) );
  INV_X1 U17163 ( .A(n14484), .ZN(n21486) );
  AOI22_X1 U17164 ( .A1(\mem[577][4] ), .A2(n14480), .B1(n26553), .B2(
        data_in[4]), .ZN(n14484) );
  INV_X1 U17165 ( .A(n14485), .ZN(n21485) );
  AOI22_X1 U17166 ( .A1(\mem[577][5] ), .A2(n14480), .B1(n26553), .B2(
        data_in[5]), .ZN(n14485) );
  INV_X1 U17167 ( .A(n14486), .ZN(n21484) );
  AOI22_X1 U17168 ( .A1(\mem[577][6] ), .A2(n14480), .B1(n26553), .B2(
        data_in[6]), .ZN(n14486) );
  INV_X1 U17169 ( .A(n14487), .ZN(n21483) );
  AOI22_X1 U17170 ( .A1(\mem[577][7] ), .A2(n14480), .B1(n26553), .B2(
        data_in[7]), .ZN(n14487) );
  INV_X1 U17171 ( .A(n14488), .ZN(n21482) );
  AOI22_X1 U17172 ( .A1(\mem[578][0] ), .A2(n14489), .B1(n26552), .B2(
        data_in[0]), .ZN(n14488) );
  INV_X1 U17173 ( .A(n14490), .ZN(n21481) );
  AOI22_X1 U17174 ( .A1(\mem[578][1] ), .A2(n14489), .B1(n26552), .B2(
        data_in[1]), .ZN(n14490) );
  INV_X1 U17175 ( .A(n14491), .ZN(n21480) );
  AOI22_X1 U17176 ( .A1(\mem[578][2] ), .A2(n14489), .B1(n26552), .B2(
        data_in[2]), .ZN(n14491) );
  INV_X1 U17177 ( .A(n14492), .ZN(n21479) );
  AOI22_X1 U17178 ( .A1(\mem[578][3] ), .A2(n14489), .B1(n26552), .B2(
        data_in[3]), .ZN(n14492) );
  INV_X1 U17179 ( .A(n14493), .ZN(n21478) );
  AOI22_X1 U17180 ( .A1(\mem[578][4] ), .A2(n14489), .B1(n26552), .B2(
        data_in[4]), .ZN(n14493) );
  INV_X1 U17181 ( .A(n14494), .ZN(n21477) );
  AOI22_X1 U17182 ( .A1(\mem[578][5] ), .A2(n14489), .B1(n26552), .B2(
        data_in[5]), .ZN(n14494) );
  INV_X1 U17183 ( .A(n14495), .ZN(n21476) );
  AOI22_X1 U17184 ( .A1(\mem[578][6] ), .A2(n14489), .B1(n26552), .B2(
        data_in[6]), .ZN(n14495) );
  INV_X1 U17185 ( .A(n14496), .ZN(n21475) );
  AOI22_X1 U17186 ( .A1(\mem[578][7] ), .A2(n14489), .B1(n26552), .B2(
        data_in[7]), .ZN(n14496) );
  INV_X1 U17187 ( .A(n14497), .ZN(n21474) );
  AOI22_X1 U17188 ( .A1(\mem[579][0] ), .A2(n14498), .B1(n26551), .B2(
        data_in[0]), .ZN(n14497) );
  INV_X1 U17189 ( .A(n14499), .ZN(n21473) );
  AOI22_X1 U17190 ( .A1(\mem[579][1] ), .A2(n14498), .B1(n26551), .B2(
        data_in[1]), .ZN(n14499) );
  INV_X1 U17191 ( .A(n14500), .ZN(n21472) );
  AOI22_X1 U17192 ( .A1(\mem[579][2] ), .A2(n14498), .B1(n26551), .B2(
        data_in[2]), .ZN(n14500) );
  INV_X1 U17193 ( .A(n14501), .ZN(n21471) );
  AOI22_X1 U17194 ( .A1(\mem[579][3] ), .A2(n14498), .B1(n26551), .B2(
        data_in[3]), .ZN(n14501) );
  INV_X1 U17195 ( .A(n14502), .ZN(n21470) );
  AOI22_X1 U17196 ( .A1(\mem[579][4] ), .A2(n14498), .B1(n26551), .B2(
        data_in[4]), .ZN(n14502) );
  INV_X1 U17197 ( .A(n14503), .ZN(n21469) );
  AOI22_X1 U17198 ( .A1(\mem[579][5] ), .A2(n14498), .B1(n26551), .B2(
        data_in[5]), .ZN(n14503) );
  INV_X1 U17199 ( .A(n14504), .ZN(n21468) );
  AOI22_X1 U17200 ( .A1(\mem[579][6] ), .A2(n14498), .B1(n26551), .B2(
        data_in[6]), .ZN(n14504) );
  INV_X1 U17201 ( .A(n14505), .ZN(n21467) );
  AOI22_X1 U17202 ( .A1(\mem[579][7] ), .A2(n14498), .B1(n26551), .B2(
        data_in[7]), .ZN(n14505) );
  INV_X1 U17203 ( .A(n14506), .ZN(n21466) );
  AOI22_X1 U17204 ( .A1(\mem[580][0] ), .A2(n14507), .B1(n26550), .B2(
        data_in[0]), .ZN(n14506) );
  INV_X1 U17205 ( .A(n14508), .ZN(n21465) );
  AOI22_X1 U17206 ( .A1(\mem[580][1] ), .A2(n14507), .B1(n26550), .B2(
        data_in[1]), .ZN(n14508) );
  INV_X1 U17207 ( .A(n14509), .ZN(n21464) );
  AOI22_X1 U17208 ( .A1(\mem[580][2] ), .A2(n14507), .B1(n26550), .B2(
        data_in[2]), .ZN(n14509) );
  INV_X1 U17209 ( .A(n14510), .ZN(n21463) );
  AOI22_X1 U17210 ( .A1(\mem[580][3] ), .A2(n14507), .B1(n26550), .B2(
        data_in[3]), .ZN(n14510) );
  INV_X1 U17211 ( .A(n14511), .ZN(n21462) );
  AOI22_X1 U17212 ( .A1(\mem[580][4] ), .A2(n14507), .B1(n26550), .B2(
        data_in[4]), .ZN(n14511) );
  INV_X1 U17213 ( .A(n14512), .ZN(n21461) );
  AOI22_X1 U17214 ( .A1(\mem[580][5] ), .A2(n14507), .B1(n26550), .B2(
        data_in[5]), .ZN(n14512) );
  INV_X1 U17215 ( .A(n14513), .ZN(n21460) );
  AOI22_X1 U17216 ( .A1(\mem[580][6] ), .A2(n14507), .B1(n26550), .B2(
        data_in[6]), .ZN(n14513) );
  INV_X1 U17217 ( .A(n14514), .ZN(n21459) );
  AOI22_X1 U17218 ( .A1(\mem[580][7] ), .A2(n14507), .B1(n26550), .B2(
        data_in[7]), .ZN(n14514) );
  INV_X1 U17219 ( .A(n14515), .ZN(n21458) );
  AOI22_X1 U17220 ( .A1(\mem[581][0] ), .A2(n14516), .B1(n26549), .B2(
        data_in[0]), .ZN(n14515) );
  INV_X1 U17221 ( .A(n14517), .ZN(n21457) );
  AOI22_X1 U17222 ( .A1(\mem[581][1] ), .A2(n14516), .B1(n26549), .B2(
        data_in[1]), .ZN(n14517) );
  INV_X1 U17223 ( .A(n14518), .ZN(n21456) );
  AOI22_X1 U17224 ( .A1(\mem[581][2] ), .A2(n14516), .B1(n26549), .B2(
        data_in[2]), .ZN(n14518) );
  INV_X1 U17225 ( .A(n14519), .ZN(n21455) );
  AOI22_X1 U17226 ( .A1(\mem[581][3] ), .A2(n14516), .B1(n26549), .B2(
        data_in[3]), .ZN(n14519) );
  INV_X1 U17227 ( .A(n14520), .ZN(n21454) );
  AOI22_X1 U17228 ( .A1(\mem[581][4] ), .A2(n14516), .B1(n26549), .B2(
        data_in[4]), .ZN(n14520) );
  INV_X1 U17229 ( .A(n14521), .ZN(n21453) );
  AOI22_X1 U17230 ( .A1(\mem[581][5] ), .A2(n14516), .B1(n26549), .B2(
        data_in[5]), .ZN(n14521) );
  INV_X1 U17231 ( .A(n14522), .ZN(n21452) );
  AOI22_X1 U17232 ( .A1(\mem[581][6] ), .A2(n14516), .B1(n26549), .B2(
        data_in[6]), .ZN(n14522) );
  INV_X1 U17233 ( .A(n14523), .ZN(n21451) );
  AOI22_X1 U17234 ( .A1(\mem[581][7] ), .A2(n14516), .B1(n26549), .B2(
        data_in[7]), .ZN(n14523) );
  INV_X1 U17235 ( .A(n14524), .ZN(n21450) );
  AOI22_X1 U17236 ( .A1(\mem[582][0] ), .A2(n14525), .B1(n26548), .B2(
        data_in[0]), .ZN(n14524) );
  INV_X1 U17237 ( .A(n14526), .ZN(n21449) );
  AOI22_X1 U17238 ( .A1(\mem[582][1] ), .A2(n14525), .B1(n26548), .B2(
        data_in[1]), .ZN(n14526) );
  INV_X1 U17239 ( .A(n14527), .ZN(n21448) );
  AOI22_X1 U17240 ( .A1(\mem[582][2] ), .A2(n14525), .B1(n26548), .B2(
        data_in[2]), .ZN(n14527) );
  INV_X1 U17241 ( .A(n14528), .ZN(n21447) );
  AOI22_X1 U17242 ( .A1(\mem[582][3] ), .A2(n14525), .B1(n26548), .B2(
        data_in[3]), .ZN(n14528) );
  INV_X1 U17243 ( .A(n14529), .ZN(n21446) );
  AOI22_X1 U17244 ( .A1(\mem[582][4] ), .A2(n14525), .B1(n26548), .B2(
        data_in[4]), .ZN(n14529) );
  INV_X1 U17245 ( .A(n14530), .ZN(n21445) );
  AOI22_X1 U17246 ( .A1(\mem[582][5] ), .A2(n14525), .B1(n26548), .B2(
        data_in[5]), .ZN(n14530) );
  INV_X1 U17247 ( .A(n14531), .ZN(n21444) );
  AOI22_X1 U17248 ( .A1(\mem[582][6] ), .A2(n14525), .B1(n26548), .B2(
        data_in[6]), .ZN(n14531) );
  INV_X1 U17249 ( .A(n14532), .ZN(n21443) );
  AOI22_X1 U17250 ( .A1(\mem[582][7] ), .A2(n14525), .B1(n26548), .B2(
        data_in[7]), .ZN(n14532) );
  INV_X1 U17251 ( .A(n14533), .ZN(n21442) );
  AOI22_X1 U17252 ( .A1(\mem[583][0] ), .A2(n14534), .B1(n26547), .B2(
        data_in[0]), .ZN(n14533) );
  INV_X1 U17253 ( .A(n14535), .ZN(n21441) );
  AOI22_X1 U17254 ( .A1(\mem[583][1] ), .A2(n14534), .B1(n26547), .B2(
        data_in[1]), .ZN(n14535) );
  INV_X1 U17255 ( .A(n14536), .ZN(n21440) );
  AOI22_X1 U17256 ( .A1(\mem[583][2] ), .A2(n14534), .B1(n26547), .B2(
        data_in[2]), .ZN(n14536) );
  INV_X1 U17257 ( .A(n14537), .ZN(n21439) );
  AOI22_X1 U17258 ( .A1(\mem[583][3] ), .A2(n14534), .B1(n26547), .B2(
        data_in[3]), .ZN(n14537) );
  INV_X1 U17259 ( .A(n14538), .ZN(n21438) );
  AOI22_X1 U17260 ( .A1(\mem[583][4] ), .A2(n14534), .B1(n26547), .B2(
        data_in[4]), .ZN(n14538) );
  INV_X1 U17261 ( .A(n14539), .ZN(n21437) );
  AOI22_X1 U17262 ( .A1(\mem[583][5] ), .A2(n14534), .B1(n26547), .B2(
        data_in[5]), .ZN(n14539) );
  INV_X1 U17263 ( .A(n14540), .ZN(n21436) );
  AOI22_X1 U17264 ( .A1(\mem[583][6] ), .A2(n14534), .B1(n26547), .B2(
        data_in[6]), .ZN(n14540) );
  INV_X1 U17265 ( .A(n14541), .ZN(n21435) );
  AOI22_X1 U17266 ( .A1(\mem[583][7] ), .A2(n14534), .B1(n26547), .B2(
        data_in[7]), .ZN(n14541) );
  INV_X1 U17267 ( .A(n14758), .ZN(n21242) );
  AOI22_X1 U17268 ( .A1(\mem[608][0] ), .A2(n14759), .B1(n26522), .B2(
        data_in[0]), .ZN(n14758) );
  INV_X1 U17269 ( .A(n14760), .ZN(n21241) );
  AOI22_X1 U17270 ( .A1(\mem[608][1] ), .A2(n14759), .B1(n26522), .B2(
        data_in[1]), .ZN(n14760) );
  INV_X1 U17271 ( .A(n14761), .ZN(n21240) );
  AOI22_X1 U17272 ( .A1(\mem[608][2] ), .A2(n14759), .B1(n26522), .B2(
        data_in[2]), .ZN(n14761) );
  INV_X1 U17273 ( .A(n14762), .ZN(n21239) );
  AOI22_X1 U17274 ( .A1(\mem[608][3] ), .A2(n14759), .B1(n26522), .B2(
        data_in[3]), .ZN(n14762) );
  INV_X1 U17275 ( .A(n14763), .ZN(n21238) );
  AOI22_X1 U17276 ( .A1(\mem[608][4] ), .A2(n14759), .B1(n26522), .B2(
        data_in[4]), .ZN(n14763) );
  INV_X1 U17277 ( .A(n14764), .ZN(n21237) );
  AOI22_X1 U17278 ( .A1(\mem[608][5] ), .A2(n14759), .B1(n26522), .B2(
        data_in[5]), .ZN(n14764) );
  INV_X1 U17279 ( .A(n14765), .ZN(n21236) );
  AOI22_X1 U17280 ( .A1(\mem[608][6] ), .A2(n14759), .B1(n26522), .B2(
        data_in[6]), .ZN(n14765) );
  INV_X1 U17281 ( .A(n14766), .ZN(n21235) );
  AOI22_X1 U17282 ( .A1(\mem[608][7] ), .A2(n14759), .B1(n26522), .B2(
        data_in[7]), .ZN(n14766) );
  INV_X1 U17283 ( .A(n14768), .ZN(n21234) );
  AOI22_X1 U17284 ( .A1(\mem[609][0] ), .A2(n14769), .B1(n26521), .B2(
        data_in[0]), .ZN(n14768) );
  INV_X1 U17285 ( .A(n14770), .ZN(n21233) );
  AOI22_X1 U17286 ( .A1(\mem[609][1] ), .A2(n14769), .B1(n26521), .B2(
        data_in[1]), .ZN(n14770) );
  INV_X1 U17287 ( .A(n14771), .ZN(n21232) );
  AOI22_X1 U17288 ( .A1(\mem[609][2] ), .A2(n14769), .B1(n26521), .B2(
        data_in[2]), .ZN(n14771) );
  INV_X1 U17289 ( .A(n14772), .ZN(n21231) );
  AOI22_X1 U17290 ( .A1(\mem[609][3] ), .A2(n14769), .B1(n26521), .B2(
        data_in[3]), .ZN(n14772) );
  INV_X1 U17291 ( .A(n14773), .ZN(n21230) );
  AOI22_X1 U17292 ( .A1(\mem[609][4] ), .A2(n14769), .B1(n26521), .B2(
        data_in[4]), .ZN(n14773) );
  INV_X1 U17293 ( .A(n14774), .ZN(n21229) );
  AOI22_X1 U17294 ( .A1(\mem[609][5] ), .A2(n14769), .B1(n26521), .B2(
        data_in[5]), .ZN(n14774) );
  INV_X1 U17295 ( .A(n14775), .ZN(n21228) );
  AOI22_X1 U17296 ( .A1(\mem[609][6] ), .A2(n14769), .B1(n26521), .B2(
        data_in[6]), .ZN(n14775) );
  INV_X1 U17297 ( .A(n14776), .ZN(n21227) );
  AOI22_X1 U17298 ( .A1(\mem[609][7] ), .A2(n14769), .B1(n26521), .B2(
        data_in[7]), .ZN(n14776) );
  INV_X1 U17299 ( .A(n14777), .ZN(n21226) );
  AOI22_X1 U17300 ( .A1(\mem[610][0] ), .A2(n14778), .B1(n26520), .B2(
        data_in[0]), .ZN(n14777) );
  INV_X1 U17301 ( .A(n14779), .ZN(n21225) );
  AOI22_X1 U17302 ( .A1(\mem[610][1] ), .A2(n14778), .B1(n26520), .B2(
        data_in[1]), .ZN(n14779) );
  INV_X1 U17303 ( .A(n14780), .ZN(n21224) );
  AOI22_X1 U17304 ( .A1(\mem[610][2] ), .A2(n14778), .B1(n26520), .B2(
        data_in[2]), .ZN(n14780) );
  INV_X1 U17305 ( .A(n14781), .ZN(n21223) );
  AOI22_X1 U17306 ( .A1(\mem[610][3] ), .A2(n14778), .B1(n26520), .B2(
        data_in[3]), .ZN(n14781) );
  INV_X1 U17307 ( .A(n14782), .ZN(n21222) );
  AOI22_X1 U17308 ( .A1(\mem[610][4] ), .A2(n14778), .B1(n26520), .B2(
        data_in[4]), .ZN(n14782) );
  INV_X1 U17309 ( .A(n14783), .ZN(n21221) );
  AOI22_X1 U17310 ( .A1(\mem[610][5] ), .A2(n14778), .B1(n26520), .B2(
        data_in[5]), .ZN(n14783) );
  INV_X1 U17311 ( .A(n14784), .ZN(n21220) );
  AOI22_X1 U17312 ( .A1(\mem[610][6] ), .A2(n14778), .B1(n26520), .B2(
        data_in[6]), .ZN(n14784) );
  INV_X1 U17313 ( .A(n14785), .ZN(n21219) );
  AOI22_X1 U17314 ( .A1(\mem[610][7] ), .A2(n14778), .B1(n26520), .B2(
        data_in[7]), .ZN(n14785) );
  INV_X1 U17315 ( .A(n14786), .ZN(n21218) );
  AOI22_X1 U17316 ( .A1(\mem[611][0] ), .A2(n14787), .B1(n26519), .B2(
        data_in[0]), .ZN(n14786) );
  INV_X1 U17317 ( .A(n14788), .ZN(n21217) );
  AOI22_X1 U17318 ( .A1(\mem[611][1] ), .A2(n14787), .B1(n26519), .B2(
        data_in[1]), .ZN(n14788) );
  INV_X1 U17319 ( .A(n14789), .ZN(n21216) );
  AOI22_X1 U17320 ( .A1(\mem[611][2] ), .A2(n14787), .B1(n26519), .B2(
        data_in[2]), .ZN(n14789) );
  INV_X1 U17321 ( .A(n14790), .ZN(n21215) );
  AOI22_X1 U17322 ( .A1(\mem[611][3] ), .A2(n14787), .B1(n26519), .B2(
        data_in[3]), .ZN(n14790) );
  INV_X1 U17323 ( .A(n14791), .ZN(n21214) );
  AOI22_X1 U17324 ( .A1(\mem[611][4] ), .A2(n14787), .B1(n26519), .B2(
        data_in[4]), .ZN(n14791) );
  INV_X1 U17325 ( .A(n14792), .ZN(n21213) );
  AOI22_X1 U17326 ( .A1(\mem[611][5] ), .A2(n14787), .B1(n26519), .B2(
        data_in[5]), .ZN(n14792) );
  INV_X1 U17327 ( .A(n14793), .ZN(n21212) );
  AOI22_X1 U17328 ( .A1(\mem[611][6] ), .A2(n14787), .B1(n26519), .B2(
        data_in[6]), .ZN(n14793) );
  INV_X1 U17329 ( .A(n14794), .ZN(n21211) );
  AOI22_X1 U17330 ( .A1(\mem[611][7] ), .A2(n14787), .B1(n26519), .B2(
        data_in[7]), .ZN(n14794) );
  INV_X1 U17331 ( .A(n14795), .ZN(n21210) );
  AOI22_X1 U17332 ( .A1(\mem[612][0] ), .A2(n14796), .B1(n26518), .B2(
        data_in[0]), .ZN(n14795) );
  INV_X1 U17333 ( .A(n14797), .ZN(n21209) );
  AOI22_X1 U17334 ( .A1(\mem[612][1] ), .A2(n14796), .B1(n26518), .B2(
        data_in[1]), .ZN(n14797) );
  INV_X1 U17335 ( .A(n14798), .ZN(n21208) );
  AOI22_X1 U17336 ( .A1(\mem[612][2] ), .A2(n14796), .B1(n26518), .B2(
        data_in[2]), .ZN(n14798) );
  INV_X1 U17337 ( .A(n14799), .ZN(n21207) );
  AOI22_X1 U17338 ( .A1(\mem[612][3] ), .A2(n14796), .B1(n26518), .B2(
        data_in[3]), .ZN(n14799) );
  INV_X1 U17339 ( .A(n14800), .ZN(n21206) );
  AOI22_X1 U17340 ( .A1(\mem[612][4] ), .A2(n14796), .B1(n26518), .B2(
        data_in[4]), .ZN(n14800) );
  INV_X1 U17341 ( .A(n14801), .ZN(n21205) );
  AOI22_X1 U17342 ( .A1(\mem[612][5] ), .A2(n14796), .B1(n26518), .B2(
        data_in[5]), .ZN(n14801) );
  INV_X1 U17343 ( .A(n14802), .ZN(n21204) );
  AOI22_X1 U17344 ( .A1(\mem[612][6] ), .A2(n14796), .B1(n26518), .B2(
        data_in[6]), .ZN(n14802) );
  INV_X1 U17345 ( .A(n14803), .ZN(n21203) );
  AOI22_X1 U17346 ( .A1(\mem[612][7] ), .A2(n14796), .B1(n26518), .B2(
        data_in[7]), .ZN(n14803) );
  INV_X1 U17347 ( .A(n14804), .ZN(n21202) );
  AOI22_X1 U17348 ( .A1(\mem[613][0] ), .A2(n14805), .B1(n26517), .B2(
        data_in[0]), .ZN(n14804) );
  INV_X1 U17349 ( .A(n14806), .ZN(n21201) );
  AOI22_X1 U17350 ( .A1(\mem[613][1] ), .A2(n14805), .B1(n26517), .B2(
        data_in[1]), .ZN(n14806) );
  INV_X1 U17351 ( .A(n14807), .ZN(n21200) );
  AOI22_X1 U17352 ( .A1(\mem[613][2] ), .A2(n14805), .B1(n26517), .B2(
        data_in[2]), .ZN(n14807) );
  INV_X1 U17353 ( .A(n14808), .ZN(n21199) );
  AOI22_X1 U17354 ( .A1(\mem[613][3] ), .A2(n14805), .B1(n26517), .B2(
        data_in[3]), .ZN(n14808) );
  INV_X1 U17355 ( .A(n14809), .ZN(n21198) );
  AOI22_X1 U17356 ( .A1(\mem[613][4] ), .A2(n14805), .B1(n26517), .B2(
        data_in[4]), .ZN(n14809) );
  INV_X1 U17357 ( .A(n14810), .ZN(n21197) );
  AOI22_X1 U17358 ( .A1(\mem[613][5] ), .A2(n14805), .B1(n26517), .B2(
        data_in[5]), .ZN(n14810) );
  INV_X1 U17359 ( .A(n14811), .ZN(n21196) );
  AOI22_X1 U17360 ( .A1(\mem[613][6] ), .A2(n14805), .B1(n26517), .B2(
        data_in[6]), .ZN(n14811) );
  INV_X1 U17361 ( .A(n14812), .ZN(n21195) );
  AOI22_X1 U17362 ( .A1(\mem[613][7] ), .A2(n14805), .B1(n26517), .B2(
        data_in[7]), .ZN(n14812) );
  INV_X1 U17363 ( .A(n14813), .ZN(n21194) );
  AOI22_X1 U17364 ( .A1(\mem[614][0] ), .A2(n14814), .B1(n26516), .B2(
        data_in[0]), .ZN(n14813) );
  INV_X1 U17365 ( .A(n14815), .ZN(n21193) );
  AOI22_X1 U17366 ( .A1(\mem[614][1] ), .A2(n14814), .B1(n26516), .B2(
        data_in[1]), .ZN(n14815) );
  INV_X1 U17367 ( .A(n14816), .ZN(n21192) );
  AOI22_X1 U17368 ( .A1(\mem[614][2] ), .A2(n14814), .B1(n26516), .B2(
        data_in[2]), .ZN(n14816) );
  INV_X1 U17369 ( .A(n14817), .ZN(n21191) );
  AOI22_X1 U17370 ( .A1(\mem[614][3] ), .A2(n14814), .B1(n26516), .B2(
        data_in[3]), .ZN(n14817) );
  INV_X1 U17371 ( .A(n14818), .ZN(n21190) );
  AOI22_X1 U17372 ( .A1(\mem[614][4] ), .A2(n14814), .B1(n26516), .B2(
        data_in[4]), .ZN(n14818) );
  INV_X1 U17373 ( .A(n14819), .ZN(n21189) );
  AOI22_X1 U17374 ( .A1(\mem[614][5] ), .A2(n14814), .B1(n26516), .B2(
        data_in[5]), .ZN(n14819) );
  INV_X1 U17375 ( .A(n14820), .ZN(n21188) );
  AOI22_X1 U17376 ( .A1(\mem[614][6] ), .A2(n14814), .B1(n26516), .B2(
        data_in[6]), .ZN(n14820) );
  INV_X1 U17377 ( .A(n14821), .ZN(n21187) );
  AOI22_X1 U17378 ( .A1(\mem[614][7] ), .A2(n14814), .B1(n26516), .B2(
        data_in[7]), .ZN(n14821) );
  INV_X1 U17379 ( .A(n14822), .ZN(n21186) );
  AOI22_X1 U17380 ( .A1(\mem[615][0] ), .A2(n14823), .B1(n26515), .B2(
        data_in[0]), .ZN(n14822) );
  INV_X1 U17381 ( .A(n14824), .ZN(n21185) );
  AOI22_X1 U17382 ( .A1(\mem[615][1] ), .A2(n14823), .B1(n26515), .B2(
        data_in[1]), .ZN(n14824) );
  INV_X1 U17383 ( .A(n14825), .ZN(n21184) );
  AOI22_X1 U17384 ( .A1(\mem[615][2] ), .A2(n14823), .B1(n26515), .B2(
        data_in[2]), .ZN(n14825) );
  INV_X1 U17385 ( .A(n14826), .ZN(n21183) );
  AOI22_X1 U17386 ( .A1(\mem[615][3] ), .A2(n14823), .B1(n26515), .B2(
        data_in[3]), .ZN(n14826) );
  INV_X1 U17387 ( .A(n14827), .ZN(n21182) );
  AOI22_X1 U17388 ( .A1(\mem[615][4] ), .A2(n14823), .B1(n26515), .B2(
        data_in[4]), .ZN(n14827) );
  INV_X1 U17389 ( .A(n14828), .ZN(n21181) );
  AOI22_X1 U17390 ( .A1(\mem[615][5] ), .A2(n14823), .B1(n26515), .B2(
        data_in[5]), .ZN(n14828) );
  INV_X1 U17391 ( .A(n14829), .ZN(n21180) );
  AOI22_X1 U17392 ( .A1(\mem[615][6] ), .A2(n14823), .B1(n26515), .B2(
        data_in[6]), .ZN(n14829) );
  INV_X1 U17393 ( .A(n14830), .ZN(n21179) );
  AOI22_X1 U17394 ( .A1(\mem[615][7] ), .A2(n14823), .B1(n26515), .B2(
        data_in[7]), .ZN(n14830) );
  INV_X1 U17395 ( .A(n15047), .ZN(n20986) );
  AOI22_X1 U17396 ( .A1(\mem[640][0] ), .A2(n15048), .B1(n26490), .B2(
        data_in[0]), .ZN(n15047) );
  INV_X1 U17397 ( .A(n15049), .ZN(n20985) );
  AOI22_X1 U17398 ( .A1(\mem[640][1] ), .A2(n15048), .B1(n26490), .B2(
        data_in[1]), .ZN(n15049) );
  INV_X1 U17399 ( .A(n15050), .ZN(n20984) );
  AOI22_X1 U17400 ( .A1(\mem[640][2] ), .A2(n15048), .B1(n26490), .B2(
        data_in[2]), .ZN(n15050) );
  INV_X1 U17401 ( .A(n15051), .ZN(n20983) );
  AOI22_X1 U17402 ( .A1(\mem[640][3] ), .A2(n15048), .B1(n26490), .B2(
        data_in[3]), .ZN(n15051) );
  INV_X1 U17403 ( .A(n15052), .ZN(n20982) );
  AOI22_X1 U17404 ( .A1(\mem[640][4] ), .A2(n15048), .B1(n26490), .B2(
        data_in[4]), .ZN(n15052) );
  INV_X1 U17405 ( .A(n15053), .ZN(n20981) );
  AOI22_X1 U17406 ( .A1(\mem[640][5] ), .A2(n15048), .B1(n26490), .B2(
        data_in[5]), .ZN(n15053) );
  INV_X1 U17407 ( .A(n15054), .ZN(n20980) );
  AOI22_X1 U17408 ( .A1(\mem[640][6] ), .A2(n15048), .B1(n26490), .B2(
        data_in[6]), .ZN(n15054) );
  INV_X1 U17409 ( .A(n15055), .ZN(n20979) );
  AOI22_X1 U17410 ( .A1(\mem[640][7] ), .A2(n15048), .B1(n26490), .B2(
        data_in[7]), .ZN(n15055) );
  INV_X1 U17411 ( .A(n15057), .ZN(n20978) );
  AOI22_X1 U17412 ( .A1(\mem[641][0] ), .A2(n15058), .B1(n26489), .B2(
        data_in[0]), .ZN(n15057) );
  INV_X1 U17413 ( .A(n15059), .ZN(n20977) );
  AOI22_X1 U17414 ( .A1(\mem[641][1] ), .A2(n15058), .B1(n26489), .B2(
        data_in[1]), .ZN(n15059) );
  INV_X1 U17415 ( .A(n15060), .ZN(n20976) );
  AOI22_X1 U17416 ( .A1(\mem[641][2] ), .A2(n15058), .B1(n26489), .B2(
        data_in[2]), .ZN(n15060) );
  INV_X1 U17417 ( .A(n15061), .ZN(n20975) );
  AOI22_X1 U17418 ( .A1(\mem[641][3] ), .A2(n15058), .B1(n26489), .B2(
        data_in[3]), .ZN(n15061) );
  INV_X1 U17419 ( .A(n15062), .ZN(n20974) );
  AOI22_X1 U17420 ( .A1(\mem[641][4] ), .A2(n15058), .B1(n26489), .B2(
        data_in[4]), .ZN(n15062) );
  INV_X1 U17421 ( .A(n15063), .ZN(n20973) );
  AOI22_X1 U17422 ( .A1(\mem[641][5] ), .A2(n15058), .B1(n26489), .B2(
        data_in[5]), .ZN(n15063) );
  INV_X1 U17423 ( .A(n15064), .ZN(n20972) );
  AOI22_X1 U17424 ( .A1(\mem[641][6] ), .A2(n15058), .B1(n26489), .B2(
        data_in[6]), .ZN(n15064) );
  INV_X1 U17425 ( .A(n15065), .ZN(n20971) );
  AOI22_X1 U17426 ( .A1(\mem[641][7] ), .A2(n15058), .B1(n26489), .B2(
        data_in[7]), .ZN(n15065) );
  INV_X1 U17427 ( .A(n15066), .ZN(n20970) );
  AOI22_X1 U17428 ( .A1(\mem[642][0] ), .A2(n15067), .B1(n26488), .B2(
        data_in[0]), .ZN(n15066) );
  INV_X1 U17429 ( .A(n15068), .ZN(n20969) );
  AOI22_X1 U17430 ( .A1(\mem[642][1] ), .A2(n15067), .B1(n26488), .B2(
        data_in[1]), .ZN(n15068) );
  INV_X1 U17431 ( .A(n15069), .ZN(n20968) );
  AOI22_X1 U17432 ( .A1(\mem[642][2] ), .A2(n15067), .B1(n26488), .B2(
        data_in[2]), .ZN(n15069) );
  INV_X1 U17433 ( .A(n15070), .ZN(n20967) );
  AOI22_X1 U17434 ( .A1(\mem[642][3] ), .A2(n15067), .B1(n26488), .B2(
        data_in[3]), .ZN(n15070) );
  INV_X1 U17435 ( .A(n15071), .ZN(n20966) );
  AOI22_X1 U17436 ( .A1(\mem[642][4] ), .A2(n15067), .B1(n26488), .B2(
        data_in[4]), .ZN(n15071) );
  INV_X1 U17437 ( .A(n15072), .ZN(n20965) );
  AOI22_X1 U17438 ( .A1(\mem[642][5] ), .A2(n15067), .B1(n26488), .B2(
        data_in[5]), .ZN(n15072) );
  INV_X1 U17439 ( .A(n15073), .ZN(n20964) );
  AOI22_X1 U17440 ( .A1(\mem[642][6] ), .A2(n15067), .B1(n26488), .B2(
        data_in[6]), .ZN(n15073) );
  INV_X1 U17441 ( .A(n15074), .ZN(n20963) );
  AOI22_X1 U17442 ( .A1(\mem[642][7] ), .A2(n15067), .B1(n26488), .B2(
        data_in[7]), .ZN(n15074) );
  INV_X1 U17443 ( .A(n15075), .ZN(n20962) );
  AOI22_X1 U17444 ( .A1(\mem[643][0] ), .A2(n15076), .B1(n26487), .B2(
        data_in[0]), .ZN(n15075) );
  INV_X1 U17445 ( .A(n15077), .ZN(n20961) );
  AOI22_X1 U17446 ( .A1(\mem[643][1] ), .A2(n15076), .B1(n26487), .B2(
        data_in[1]), .ZN(n15077) );
  INV_X1 U17447 ( .A(n15078), .ZN(n20960) );
  AOI22_X1 U17448 ( .A1(\mem[643][2] ), .A2(n15076), .B1(n26487), .B2(
        data_in[2]), .ZN(n15078) );
  INV_X1 U17449 ( .A(n15079), .ZN(n20959) );
  AOI22_X1 U17450 ( .A1(\mem[643][3] ), .A2(n15076), .B1(n26487), .B2(
        data_in[3]), .ZN(n15079) );
  INV_X1 U17451 ( .A(n15080), .ZN(n20958) );
  AOI22_X1 U17452 ( .A1(\mem[643][4] ), .A2(n15076), .B1(n26487), .B2(
        data_in[4]), .ZN(n15080) );
  INV_X1 U17453 ( .A(n15081), .ZN(n20957) );
  AOI22_X1 U17454 ( .A1(\mem[643][5] ), .A2(n15076), .B1(n26487), .B2(
        data_in[5]), .ZN(n15081) );
  INV_X1 U17455 ( .A(n15082), .ZN(n20956) );
  AOI22_X1 U17456 ( .A1(\mem[643][6] ), .A2(n15076), .B1(n26487), .B2(
        data_in[6]), .ZN(n15082) );
  INV_X1 U17457 ( .A(n15083), .ZN(n20955) );
  AOI22_X1 U17458 ( .A1(\mem[643][7] ), .A2(n15076), .B1(n26487), .B2(
        data_in[7]), .ZN(n15083) );
  INV_X1 U17459 ( .A(n15084), .ZN(n20954) );
  AOI22_X1 U17460 ( .A1(\mem[644][0] ), .A2(n15085), .B1(n26486), .B2(
        data_in[0]), .ZN(n15084) );
  INV_X1 U17461 ( .A(n15086), .ZN(n20953) );
  AOI22_X1 U17462 ( .A1(\mem[644][1] ), .A2(n15085), .B1(n26486), .B2(
        data_in[1]), .ZN(n15086) );
  INV_X1 U17463 ( .A(n15087), .ZN(n20952) );
  AOI22_X1 U17464 ( .A1(\mem[644][2] ), .A2(n15085), .B1(n26486), .B2(
        data_in[2]), .ZN(n15087) );
  INV_X1 U17465 ( .A(n15088), .ZN(n20951) );
  AOI22_X1 U17466 ( .A1(\mem[644][3] ), .A2(n15085), .B1(n26486), .B2(
        data_in[3]), .ZN(n15088) );
  INV_X1 U17467 ( .A(n15089), .ZN(n20950) );
  AOI22_X1 U17468 ( .A1(\mem[644][4] ), .A2(n15085), .B1(n26486), .B2(
        data_in[4]), .ZN(n15089) );
  INV_X1 U17469 ( .A(n15090), .ZN(n20949) );
  AOI22_X1 U17470 ( .A1(\mem[644][5] ), .A2(n15085), .B1(n26486), .B2(
        data_in[5]), .ZN(n15090) );
  INV_X1 U17471 ( .A(n15091), .ZN(n20948) );
  AOI22_X1 U17472 ( .A1(\mem[644][6] ), .A2(n15085), .B1(n26486), .B2(
        data_in[6]), .ZN(n15091) );
  INV_X1 U17473 ( .A(n15092), .ZN(n20947) );
  AOI22_X1 U17474 ( .A1(\mem[644][7] ), .A2(n15085), .B1(n26486), .B2(
        data_in[7]), .ZN(n15092) );
  INV_X1 U17475 ( .A(n15093), .ZN(n20946) );
  AOI22_X1 U17476 ( .A1(\mem[645][0] ), .A2(n15094), .B1(n26485), .B2(
        data_in[0]), .ZN(n15093) );
  INV_X1 U17477 ( .A(n15095), .ZN(n20945) );
  AOI22_X1 U17478 ( .A1(\mem[645][1] ), .A2(n15094), .B1(n26485), .B2(
        data_in[1]), .ZN(n15095) );
  INV_X1 U17479 ( .A(n15096), .ZN(n20944) );
  AOI22_X1 U17480 ( .A1(\mem[645][2] ), .A2(n15094), .B1(n26485), .B2(
        data_in[2]), .ZN(n15096) );
  INV_X1 U17481 ( .A(n15097), .ZN(n20943) );
  AOI22_X1 U17482 ( .A1(\mem[645][3] ), .A2(n15094), .B1(n26485), .B2(
        data_in[3]), .ZN(n15097) );
  INV_X1 U17483 ( .A(n15098), .ZN(n20942) );
  AOI22_X1 U17484 ( .A1(\mem[645][4] ), .A2(n15094), .B1(n26485), .B2(
        data_in[4]), .ZN(n15098) );
  INV_X1 U17485 ( .A(n15099), .ZN(n20941) );
  AOI22_X1 U17486 ( .A1(\mem[645][5] ), .A2(n15094), .B1(n26485), .B2(
        data_in[5]), .ZN(n15099) );
  INV_X1 U17487 ( .A(n15100), .ZN(n20940) );
  AOI22_X1 U17488 ( .A1(\mem[645][6] ), .A2(n15094), .B1(n26485), .B2(
        data_in[6]), .ZN(n15100) );
  INV_X1 U17489 ( .A(n15101), .ZN(n20939) );
  AOI22_X1 U17490 ( .A1(\mem[645][7] ), .A2(n15094), .B1(n26485), .B2(
        data_in[7]), .ZN(n15101) );
  INV_X1 U17491 ( .A(n15102), .ZN(n20938) );
  AOI22_X1 U17492 ( .A1(\mem[646][0] ), .A2(n15103), .B1(n26484), .B2(
        data_in[0]), .ZN(n15102) );
  INV_X1 U17493 ( .A(n15104), .ZN(n20937) );
  AOI22_X1 U17494 ( .A1(\mem[646][1] ), .A2(n15103), .B1(n26484), .B2(
        data_in[1]), .ZN(n15104) );
  INV_X1 U17495 ( .A(n15105), .ZN(n20936) );
  AOI22_X1 U17496 ( .A1(\mem[646][2] ), .A2(n15103), .B1(n26484), .B2(
        data_in[2]), .ZN(n15105) );
  INV_X1 U17497 ( .A(n15106), .ZN(n20935) );
  AOI22_X1 U17498 ( .A1(\mem[646][3] ), .A2(n15103), .B1(n26484), .B2(
        data_in[3]), .ZN(n15106) );
  INV_X1 U17499 ( .A(n15107), .ZN(n20934) );
  AOI22_X1 U17500 ( .A1(\mem[646][4] ), .A2(n15103), .B1(n26484), .B2(
        data_in[4]), .ZN(n15107) );
  INV_X1 U17501 ( .A(n15108), .ZN(n20933) );
  AOI22_X1 U17502 ( .A1(\mem[646][5] ), .A2(n15103), .B1(n26484), .B2(
        data_in[5]), .ZN(n15108) );
  INV_X1 U17503 ( .A(n15109), .ZN(n20932) );
  AOI22_X1 U17504 ( .A1(\mem[646][6] ), .A2(n15103), .B1(n26484), .B2(
        data_in[6]), .ZN(n15109) );
  INV_X1 U17505 ( .A(n15110), .ZN(n20931) );
  AOI22_X1 U17506 ( .A1(\mem[646][7] ), .A2(n15103), .B1(n26484), .B2(
        data_in[7]), .ZN(n15110) );
  INV_X1 U17507 ( .A(n15111), .ZN(n20930) );
  AOI22_X1 U17508 ( .A1(\mem[647][0] ), .A2(n15112), .B1(n26483), .B2(
        data_in[0]), .ZN(n15111) );
  INV_X1 U17509 ( .A(n15113), .ZN(n20929) );
  AOI22_X1 U17510 ( .A1(\mem[647][1] ), .A2(n15112), .B1(n26483), .B2(
        data_in[1]), .ZN(n15113) );
  INV_X1 U17511 ( .A(n15114), .ZN(n20928) );
  AOI22_X1 U17512 ( .A1(\mem[647][2] ), .A2(n15112), .B1(n26483), .B2(
        data_in[2]), .ZN(n15114) );
  INV_X1 U17513 ( .A(n15115), .ZN(n20927) );
  AOI22_X1 U17514 ( .A1(\mem[647][3] ), .A2(n15112), .B1(n26483), .B2(
        data_in[3]), .ZN(n15115) );
  INV_X1 U17515 ( .A(n15116), .ZN(n20926) );
  AOI22_X1 U17516 ( .A1(\mem[647][4] ), .A2(n15112), .B1(n26483), .B2(
        data_in[4]), .ZN(n15116) );
  INV_X1 U17517 ( .A(n15117), .ZN(n20925) );
  AOI22_X1 U17518 ( .A1(\mem[647][5] ), .A2(n15112), .B1(n26483), .B2(
        data_in[5]), .ZN(n15117) );
  INV_X1 U17519 ( .A(n15118), .ZN(n20924) );
  AOI22_X1 U17520 ( .A1(\mem[647][6] ), .A2(n15112), .B1(n26483), .B2(
        data_in[6]), .ZN(n15118) );
  INV_X1 U17521 ( .A(n15119), .ZN(n20923) );
  AOI22_X1 U17522 ( .A1(\mem[647][7] ), .A2(n15112), .B1(n26483), .B2(
        data_in[7]), .ZN(n15119) );
  INV_X1 U17523 ( .A(n15336), .ZN(n20730) );
  AOI22_X1 U17524 ( .A1(\mem[672][0] ), .A2(n15337), .B1(n26458), .B2(
        data_in[0]), .ZN(n15336) );
  INV_X1 U17525 ( .A(n15338), .ZN(n20729) );
  AOI22_X1 U17526 ( .A1(\mem[672][1] ), .A2(n15337), .B1(n26458), .B2(
        data_in[1]), .ZN(n15338) );
  INV_X1 U17527 ( .A(n15339), .ZN(n20728) );
  AOI22_X1 U17528 ( .A1(\mem[672][2] ), .A2(n15337), .B1(n26458), .B2(
        data_in[2]), .ZN(n15339) );
  INV_X1 U17529 ( .A(n15340), .ZN(n20727) );
  AOI22_X1 U17530 ( .A1(\mem[672][3] ), .A2(n15337), .B1(n26458), .B2(
        data_in[3]), .ZN(n15340) );
  INV_X1 U17531 ( .A(n15341), .ZN(n20726) );
  AOI22_X1 U17532 ( .A1(\mem[672][4] ), .A2(n15337), .B1(n26458), .B2(
        data_in[4]), .ZN(n15341) );
  INV_X1 U17533 ( .A(n15342), .ZN(n20725) );
  AOI22_X1 U17534 ( .A1(\mem[672][5] ), .A2(n15337), .B1(n26458), .B2(
        data_in[5]), .ZN(n15342) );
  INV_X1 U17535 ( .A(n15343), .ZN(n20724) );
  AOI22_X1 U17536 ( .A1(\mem[672][6] ), .A2(n15337), .B1(n26458), .B2(
        data_in[6]), .ZN(n15343) );
  INV_X1 U17537 ( .A(n15344), .ZN(n20723) );
  AOI22_X1 U17538 ( .A1(\mem[672][7] ), .A2(n15337), .B1(n26458), .B2(
        data_in[7]), .ZN(n15344) );
  INV_X1 U17539 ( .A(n15346), .ZN(n20722) );
  AOI22_X1 U17540 ( .A1(\mem[673][0] ), .A2(n15347), .B1(n26457), .B2(
        data_in[0]), .ZN(n15346) );
  INV_X1 U17541 ( .A(n15348), .ZN(n20721) );
  AOI22_X1 U17542 ( .A1(\mem[673][1] ), .A2(n15347), .B1(n26457), .B2(
        data_in[1]), .ZN(n15348) );
  INV_X1 U17543 ( .A(n15349), .ZN(n20720) );
  AOI22_X1 U17544 ( .A1(\mem[673][2] ), .A2(n15347), .B1(n26457), .B2(
        data_in[2]), .ZN(n15349) );
  INV_X1 U17545 ( .A(n15350), .ZN(n20719) );
  AOI22_X1 U17546 ( .A1(\mem[673][3] ), .A2(n15347), .B1(n26457), .B2(
        data_in[3]), .ZN(n15350) );
  INV_X1 U17547 ( .A(n15351), .ZN(n20718) );
  AOI22_X1 U17548 ( .A1(\mem[673][4] ), .A2(n15347), .B1(n26457), .B2(
        data_in[4]), .ZN(n15351) );
  INV_X1 U17549 ( .A(n15352), .ZN(n20717) );
  AOI22_X1 U17550 ( .A1(\mem[673][5] ), .A2(n15347), .B1(n26457), .B2(
        data_in[5]), .ZN(n15352) );
  INV_X1 U17551 ( .A(n15353), .ZN(n20716) );
  AOI22_X1 U17552 ( .A1(\mem[673][6] ), .A2(n15347), .B1(n26457), .B2(
        data_in[6]), .ZN(n15353) );
  INV_X1 U17553 ( .A(n15354), .ZN(n20715) );
  AOI22_X1 U17554 ( .A1(\mem[673][7] ), .A2(n15347), .B1(n26457), .B2(
        data_in[7]), .ZN(n15354) );
  INV_X1 U17555 ( .A(n15355), .ZN(n20714) );
  AOI22_X1 U17556 ( .A1(\mem[674][0] ), .A2(n15356), .B1(n26456), .B2(
        data_in[0]), .ZN(n15355) );
  INV_X1 U17557 ( .A(n15357), .ZN(n20713) );
  AOI22_X1 U17558 ( .A1(\mem[674][1] ), .A2(n15356), .B1(n26456), .B2(
        data_in[1]), .ZN(n15357) );
  INV_X1 U17559 ( .A(n15358), .ZN(n20712) );
  AOI22_X1 U17560 ( .A1(\mem[674][2] ), .A2(n15356), .B1(n26456), .B2(
        data_in[2]), .ZN(n15358) );
  INV_X1 U17561 ( .A(n15359), .ZN(n20711) );
  AOI22_X1 U17562 ( .A1(\mem[674][3] ), .A2(n15356), .B1(n26456), .B2(
        data_in[3]), .ZN(n15359) );
  INV_X1 U17563 ( .A(n15360), .ZN(n20710) );
  AOI22_X1 U17564 ( .A1(\mem[674][4] ), .A2(n15356), .B1(n26456), .B2(
        data_in[4]), .ZN(n15360) );
  INV_X1 U17565 ( .A(n15361), .ZN(n20709) );
  AOI22_X1 U17566 ( .A1(\mem[674][5] ), .A2(n15356), .B1(n26456), .B2(
        data_in[5]), .ZN(n15361) );
  INV_X1 U17567 ( .A(n15362), .ZN(n20708) );
  AOI22_X1 U17568 ( .A1(\mem[674][6] ), .A2(n15356), .B1(n26456), .B2(
        data_in[6]), .ZN(n15362) );
  INV_X1 U17569 ( .A(n15363), .ZN(n20707) );
  AOI22_X1 U17570 ( .A1(\mem[674][7] ), .A2(n15356), .B1(n26456), .B2(
        data_in[7]), .ZN(n15363) );
  INV_X1 U17571 ( .A(n15364), .ZN(n20706) );
  AOI22_X1 U17572 ( .A1(\mem[675][0] ), .A2(n15365), .B1(n26455), .B2(
        data_in[0]), .ZN(n15364) );
  INV_X1 U17573 ( .A(n15366), .ZN(n20705) );
  AOI22_X1 U17574 ( .A1(\mem[675][1] ), .A2(n15365), .B1(n26455), .B2(
        data_in[1]), .ZN(n15366) );
  INV_X1 U17575 ( .A(n15367), .ZN(n20704) );
  AOI22_X1 U17576 ( .A1(\mem[675][2] ), .A2(n15365), .B1(n26455), .B2(
        data_in[2]), .ZN(n15367) );
  INV_X1 U17577 ( .A(n15368), .ZN(n20703) );
  AOI22_X1 U17578 ( .A1(\mem[675][3] ), .A2(n15365), .B1(n26455), .B2(
        data_in[3]), .ZN(n15368) );
  INV_X1 U17579 ( .A(n15369), .ZN(n20702) );
  AOI22_X1 U17580 ( .A1(\mem[675][4] ), .A2(n15365), .B1(n26455), .B2(
        data_in[4]), .ZN(n15369) );
  INV_X1 U17581 ( .A(n15370), .ZN(n20701) );
  AOI22_X1 U17582 ( .A1(\mem[675][5] ), .A2(n15365), .B1(n26455), .B2(
        data_in[5]), .ZN(n15370) );
  INV_X1 U17583 ( .A(n15371), .ZN(n20700) );
  AOI22_X1 U17584 ( .A1(\mem[675][6] ), .A2(n15365), .B1(n26455), .B2(
        data_in[6]), .ZN(n15371) );
  INV_X1 U17585 ( .A(n15372), .ZN(n20699) );
  AOI22_X1 U17586 ( .A1(\mem[675][7] ), .A2(n15365), .B1(n26455), .B2(
        data_in[7]), .ZN(n15372) );
  INV_X1 U17587 ( .A(n15373), .ZN(n20698) );
  AOI22_X1 U17588 ( .A1(\mem[676][0] ), .A2(n15374), .B1(n26454), .B2(
        data_in[0]), .ZN(n15373) );
  INV_X1 U17589 ( .A(n15375), .ZN(n20697) );
  AOI22_X1 U17590 ( .A1(\mem[676][1] ), .A2(n15374), .B1(n26454), .B2(
        data_in[1]), .ZN(n15375) );
  INV_X1 U17591 ( .A(n15376), .ZN(n20696) );
  AOI22_X1 U17592 ( .A1(\mem[676][2] ), .A2(n15374), .B1(n26454), .B2(
        data_in[2]), .ZN(n15376) );
  INV_X1 U17593 ( .A(n15377), .ZN(n20695) );
  AOI22_X1 U17594 ( .A1(\mem[676][3] ), .A2(n15374), .B1(n26454), .B2(
        data_in[3]), .ZN(n15377) );
  INV_X1 U17595 ( .A(n15378), .ZN(n20694) );
  AOI22_X1 U17596 ( .A1(\mem[676][4] ), .A2(n15374), .B1(n26454), .B2(
        data_in[4]), .ZN(n15378) );
  INV_X1 U17597 ( .A(n15379), .ZN(n20693) );
  AOI22_X1 U17598 ( .A1(\mem[676][5] ), .A2(n15374), .B1(n26454), .B2(
        data_in[5]), .ZN(n15379) );
  INV_X1 U17599 ( .A(n15380), .ZN(n20692) );
  AOI22_X1 U17600 ( .A1(\mem[676][6] ), .A2(n15374), .B1(n26454), .B2(
        data_in[6]), .ZN(n15380) );
  INV_X1 U17601 ( .A(n15381), .ZN(n20691) );
  AOI22_X1 U17602 ( .A1(\mem[676][7] ), .A2(n15374), .B1(n26454), .B2(
        data_in[7]), .ZN(n15381) );
  INV_X1 U17603 ( .A(n15382), .ZN(n20690) );
  AOI22_X1 U17604 ( .A1(\mem[677][0] ), .A2(n15383), .B1(n26453), .B2(
        data_in[0]), .ZN(n15382) );
  INV_X1 U17605 ( .A(n15384), .ZN(n20689) );
  AOI22_X1 U17606 ( .A1(\mem[677][1] ), .A2(n15383), .B1(n26453), .B2(
        data_in[1]), .ZN(n15384) );
  INV_X1 U17607 ( .A(n15385), .ZN(n20688) );
  AOI22_X1 U17608 ( .A1(\mem[677][2] ), .A2(n15383), .B1(n26453), .B2(
        data_in[2]), .ZN(n15385) );
  INV_X1 U17609 ( .A(n15386), .ZN(n20687) );
  AOI22_X1 U17610 ( .A1(\mem[677][3] ), .A2(n15383), .B1(n26453), .B2(
        data_in[3]), .ZN(n15386) );
  INV_X1 U17611 ( .A(n15387), .ZN(n20686) );
  AOI22_X1 U17612 ( .A1(\mem[677][4] ), .A2(n15383), .B1(n26453), .B2(
        data_in[4]), .ZN(n15387) );
  INV_X1 U17613 ( .A(n15388), .ZN(n20685) );
  AOI22_X1 U17614 ( .A1(\mem[677][5] ), .A2(n15383), .B1(n26453), .B2(
        data_in[5]), .ZN(n15388) );
  INV_X1 U17615 ( .A(n15389), .ZN(n20684) );
  AOI22_X1 U17616 ( .A1(\mem[677][6] ), .A2(n15383), .B1(n26453), .B2(
        data_in[6]), .ZN(n15389) );
  INV_X1 U17617 ( .A(n15390), .ZN(n20683) );
  AOI22_X1 U17618 ( .A1(\mem[677][7] ), .A2(n15383), .B1(n26453), .B2(
        data_in[7]), .ZN(n15390) );
  INV_X1 U17619 ( .A(n15391), .ZN(n20682) );
  AOI22_X1 U17620 ( .A1(\mem[678][0] ), .A2(n15392), .B1(n26452), .B2(
        data_in[0]), .ZN(n15391) );
  INV_X1 U17621 ( .A(n15393), .ZN(n20681) );
  AOI22_X1 U17622 ( .A1(\mem[678][1] ), .A2(n15392), .B1(n26452), .B2(
        data_in[1]), .ZN(n15393) );
  INV_X1 U17623 ( .A(n15394), .ZN(n20680) );
  AOI22_X1 U17624 ( .A1(\mem[678][2] ), .A2(n15392), .B1(n26452), .B2(
        data_in[2]), .ZN(n15394) );
  INV_X1 U17625 ( .A(n15395), .ZN(n20679) );
  AOI22_X1 U17626 ( .A1(\mem[678][3] ), .A2(n15392), .B1(n26452), .B2(
        data_in[3]), .ZN(n15395) );
  INV_X1 U17627 ( .A(n15396), .ZN(n20678) );
  AOI22_X1 U17628 ( .A1(\mem[678][4] ), .A2(n15392), .B1(n26452), .B2(
        data_in[4]), .ZN(n15396) );
  INV_X1 U17629 ( .A(n15397), .ZN(n20677) );
  AOI22_X1 U17630 ( .A1(\mem[678][5] ), .A2(n15392), .B1(n26452), .B2(
        data_in[5]), .ZN(n15397) );
  INV_X1 U17631 ( .A(n15398), .ZN(n20676) );
  AOI22_X1 U17632 ( .A1(\mem[678][6] ), .A2(n15392), .B1(n26452), .B2(
        data_in[6]), .ZN(n15398) );
  INV_X1 U17633 ( .A(n15399), .ZN(n20675) );
  AOI22_X1 U17634 ( .A1(\mem[678][7] ), .A2(n15392), .B1(n26452), .B2(
        data_in[7]), .ZN(n15399) );
  INV_X1 U17635 ( .A(n15400), .ZN(n20674) );
  AOI22_X1 U17636 ( .A1(\mem[679][0] ), .A2(n15401), .B1(n26451), .B2(
        data_in[0]), .ZN(n15400) );
  INV_X1 U17637 ( .A(n15402), .ZN(n20673) );
  AOI22_X1 U17638 ( .A1(\mem[679][1] ), .A2(n15401), .B1(n26451), .B2(
        data_in[1]), .ZN(n15402) );
  INV_X1 U17639 ( .A(n15403), .ZN(n20672) );
  AOI22_X1 U17640 ( .A1(\mem[679][2] ), .A2(n15401), .B1(n26451), .B2(
        data_in[2]), .ZN(n15403) );
  INV_X1 U17641 ( .A(n15404), .ZN(n20671) );
  AOI22_X1 U17642 ( .A1(\mem[679][3] ), .A2(n15401), .B1(n26451), .B2(
        data_in[3]), .ZN(n15404) );
  INV_X1 U17643 ( .A(n15405), .ZN(n20670) );
  AOI22_X1 U17644 ( .A1(\mem[679][4] ), .A2(n15401), .B1(n26451), .B2(
        data_in[4]), .ZN(n15405) );
  INV_X1 U17645 ( .A(n15406), .ZN(n20669) );
  AOI22_X1 U17646 ( .A1(\mem[679][5] ), .A2(n15401), .B1(n26451), .B2(
        data_in[5]), .ZN(n15406) );
  INV_X1 U17647 ( .A(n15407), .ZN(n20668) );
  AOI22_X1 U17648 ( .A1(\mem[679][6] ), .A2(n15401), .B1(n26451), .B2(
        data_in[6]), .ZN(n15407) );
  INV_X1 U17649 ( .A(n15408), .ZN(n20667) );
  AOI22_X1 U17650 ( .A1(\mem[679][7] ), .A2(n15401), .B1(n26451), .B2(
        data_in[7]), .ZN(n15408) );
  INV_X1 U17651 ( .A(n15625), .ZN(n20474) );
  AOI22_X1 U17652 ( .A1(\mem[704][0] ), .A2(n15626), .B1(n26426), .B2(
        data_in[0]), .ZN(n15625) );
  INV_X1 U17653 ( .A(n15627), .ZN(n20473) );
  AOI22_X1 U17654 ( .A1(\mem[704][1] ), .A2(n15626), .B1(n26426), .B2(
        data_in[1]), .ZN(n15627) );
  INV_X1 U17655 ( .A(n15628), .ZN(n20472) );
  AOI22_X1 U17656 ( .A1(\mem[704][2] ), .A2(n15626), .B1(n26426), .B2(
        data_in[2]), .ZN(n15628) );
  INV_X1 U17657 ( .A(n15629), .ZN(n20471) );
  AOI22_X1 U17658 ( .A1(\mem[704][3] ), .A2(n15626), .B1(n26426), .B2(
        data_in[3]), .ZN(n15629) );
  INV_X1 U17659 ( .A(n15630), .ZN(n20470) );
  AOI22_X1 U17660 ( .A1(\mem[704][4] ), .A2(n15626), .B1(n26426), .B2(
        data_in[4]), .ZN(n15630) );
  INV_X1 U17661 ( .A(n15631), .ZN(n20469) );
  AOI22_X1 U17662 ( .A1(\mem[704][5] ), .A2(n15626), .B1(n26426), .B2(
        data_in[5]), .ZN(n15631) );
  INV_X1 U17663 ( .A(n15632), .ZN(n20468) );
  AOI22_X1 U17664 ( .A1(\mem[704][6] ), .A2(n15626), .B1(n26426), .B2(
        data_in[6]), .ZN(n15632) );
  INV_X1 U17665 ( .A(n15633), .ZN(n20467) );
  AOI22_X1 U17666 ( .A1(\mem[704][7] ), .A2(n15626), .B1(n26426), .B2(
        data_in[7]), .ZN(n15633) );
  INV_X1 U17667 ( .A(n15635), .ZN(n20466) );
  AOI22_X1 U17668 ( .A1(\mem[705][0] ), .A2(n15636), .B1(n26425), .B2(
        data_in[0]), .ZN(n15635) );
  INV_X1 U17669 ( .A(n15637), .ZN(n20465) );
  AOI22_X1 U17670 ( .A1(\mem[705][1] ), .A2(n15636), .B1(n26425), .B2(
        data_in[1]), .ZN(n15637) );
  INV_X1 U17671 ( .A(n15638), .ZN(n20464) );
  AOI22_X1 U17672 ( .A1(\mem[705][2] ), .A2(n15636), .B1(n26425), .B2(
        data_in[2]), .ZN(n15638) );
  INV_X1 U17673 ( .A(n15639), .ZN(n20463) );
  AOI22_X1 U17674 ( .A1(\mem[705][3] ), .A2(n15636), .B1(n26425), .B2(
        data_in[3]), .ZN(n15639) );
  INV_X1 U17675 ( .A(n15640), .ZN(n20462) );
  AOI22_X1 U17676 ( .A1(\mem[705][4] ), .A2(n15636), .B1(n26425), .B2(
        data_in[4]), .ZN(n15640) );
  INV_X1 U17677 ( .A(n15641), .ZN(n20461) );
  AOI22_X1 U17678 ( .A1(\mem[705][5] ), .A2(n15636), .B1(n26425), .B2(
        data_in[5]), .ZN(n15641) );
  INV_X1 U17679 ( .A(n15642), .ZN(n20460) );
  AOI22_X1 U17680 ( .A1(\mem[705][6] ), .A2(n15636), .B1(n26425), .B2(
        data_in[6]), .ZN(n15642) );
  INV_X1 U17681 ( .A(n15643), .ZN(n20459) );
  AOI22_X1 U17682 ( .A1(\mem[705][7] ), .A2(n15636), .B1(n26425), .B2(
        data_in[7]), .ZN(n15643) );
  INV_X1 U17683 ( .A(n15644), .ZN(n20458) );
  AOI22_X1 U17684 ( .A1(\mem[706][0] ), .A2(n15645), .B1(n26424), .B2(
        data_in[0]), .ZN(n15644) );
  INV_X1 U17685 ( .A(n15646), .ZN(n20457) );
  AOI22_X1 U17686 ( .A1(\mem[706][1] ), .A2(n15645), .B1(n26424), .B2(
        data_in[1]), .ZN(n15646) );
  INV_X1 U17687 ( .A(n15647), .ZN(n20456) );
  AOI22_X1 U17688 ( .A1(\mem[706][2] ), .A2(n15645), .B1(n26424), .B2(
        data_in[2]), .ZN(n15647) );
  INV_X1 U17689 ( .A(n15648), .ZN(n20455) );
  AOI22_X1 U17690 ( .A1(\mem[706][3] ), .A2(n15645), .B1(n26424), .B2(
        data_in[3]), .ZN(n15648) );
  INV_X1 U17691 ( .A(n15649), .ZN(n20454) );
  AOI22_X1 U17692 ( .A1(\mem[706][4] ), .A2(n15645), .B1(n26424), .B2(
        data_in[4]), .ZN(n15649) );
  INV_X1 U17693 ( .A(n15650), .ZN(n20453) );
  AOI22_X1 U17694 ( .A1(\mem[706][5] ), .A2(n15645), .B1(n26424), .B2(
        data_in[5]), .ZN(n15650) );
  INV_X1 U17695 ( .A(n15651), .ZN(n20452) );
  AOI22_X1 U17696 ( .A1(\mem[706][6] ), .A2(n15645), .B1(n26424), .B2(
        data_in[6]), .ZN(n15651) );
  INV_X1 U17697 ( .A(n15652), .ZN(n20451) );
  AOI22_X1 U17698 ( .A1(\mem[706][7] ), .A2(n15645), .B1(n26424), .B2(
        data_in[7]), .ZN(n15652) );
  INV_X1 U17699 ( .A(n15653), .ZN(n20450) );
  AOI22_X1 U17700 ( .A1(\mem[707][0] ), .A2(n15654), .B1(n26423), .B2(
        data_in[0]), .ZN(n15653) );
  INV_X1 U17701 ( .A(n15655), .ZN(n20449) );
  AOI22_X1 U17702 ( .A1(\mem[707][1] ), .A2(n15654), .B1(n26423), .B2(
        data_in[1]), .ZN(n15655) );
  INV_X1 U17703 ( .A(n15656), .ZN(n20448) );
  AOI22_X1 U17704 ( .A1(\mem[707][2] ), .A2(n15654), .B1(n26423), .B2(
        data_in[2]), .ZN(n15656) );
  INV_X1 U17705 ( .A(n15657), .ZN(n20447) );
  AOI22_X1 U17706 ( .A1(\mem[707][3] ), .A2(n15654), .B1(n26423), .B2(
        data_in[3]), .ZN(n15657) );
  INV_X1 U17707 ( .A(n15658), .ZN(n20446) );
  AOI22_X1 U17708 ( .A1(\mem[707][4] ), .A2(n15654), .B1(n26423), .B2(
        data_in[4]), .ZN(n15658) );
  INV_X1 U17709 ( .A(n15659), .ZN(n20445) );
  AOI22_X1 U17710 ( .A1(\mem[707][5] ), .A2(n15654), .B1(n26423), .B2(
        data_in[5]), .ZN(n15659) );
  INV_X1 U17711 ( .A(n15660), .ZN(n20444) );
  AOI22_X1 U17712 ( .A1(\mem[707][6] ), .A2(n15654), .B1(n26423), .B2(
        data_in[6]), .ZN(n15660) );
  INV_X1 U17713 ( .A(n15661), .ZN(n20443) );
  AOI22_X1 U17714 ( .A1(\mem[707][7] ), .A2(n15654), .B1(n26423), .B2(
        data_in[7]), .ZN(n15661) );
  INV_X1 U17715 ( .A(n15662), .ZN(n20442) );
  AOI22_X1 U17716 ( .A1(\mem[708][0] ), .A2(n15663), .B1(n26422), .B2(
        data_in[0]), .ZN(n15662) );
  INV_X1 U17717 ( .A(n15664), .ZN(n20441) );
  AOI22_X1 U17718 ( .A1(\mem[708][1] ), .A2(n15663), .B1(n26422), .B2(
        data_in[1]), .ZN(n15664) );
  INV_X1 U17719 ( .A(n15665), .ZN(n20440) );
  AOI22_X1 U17720 ( .A1(\mem[708][2] ), .A2(n15663), .B1(n26422), .B2(
        data_in[2]), .ZN(n15665) );
  INV_X1 U17721 ( .A(n15666), .ZN(n20439) );
  AOI22_X1 U17722 ( .A1(\mem[708][3] ), .A2(n15663), .B1(n26422), .B2(
        data_in[3]), .ZN(n15666) );
  INV_X1 U17723 ( .A(n15667), .ZN(n20438) );
  AOI22_X1 U17724 ( .A1(\mem[708][4] ), .A2(n15663), .B1(n26422), .B2(
        data_in[4]), .ZN(n15667) );
  INV_X1 U17725 ( .A(n15668), .ZN(n20437) );
  AOI22_X1 U17726 ( .A1(\mem[708][5] ), .A2(n15663), .B1(n26422), .B2(
        data_in[5]), .ZN(n15668) );
  INV_X1 U17727 ( .A(n15669), .ZN(n20436) );
  AOI22_X1 U17728 ( .A1(\mem[708][6] ), .A2(n15663), .B1(n26422), .B2(
        data_in[6]), .ZN(n15669) );
  INV_X1 U17729 ( .A(n15670), .ZN(n20435) );
  AOI22_X1 U17730 ( .A1(\mem[708][7] ), .A2(n15663), .B1(n26422), .B2(
        data_in[7]), .ZN(n15670) );
  INV_X1 U17731 ( .A(n15671), .ZN(n20434) );
  AOI22_X1 U17732 ( .A1(\mem[709][0] ), .A2(n15672), .B1(n26421), .B2(
        data_in[0]), .ZN(n15671) );
  INV_X1 U17733 ( .A(n15673), .ZN(n20433) );
  AOI22_X1 U17734 ( .A1(\mem[709][1] ), .A2(n15672), .B1(n26421), .B2(
        data_in[1]), .ZN(n15673) );
  INV_X1 U17735 ( .A(n15674), .ZN(n20432) );
  AOI22_X1 U17736 ( .A1(\mem[709][2] ), .A2(n15672), .B1(n26421), .B2(
        data_in[2]), .ZN(n15674) );
  INV_X1 U17737 ( .A(n15675), .ZN(n20431) );
  AOI22_X1 U17738 ( .A1(\mem[709][3] ), .A2(n15672), .B1(n26421), .B2(
        data_in[3]), .ZN(n15675) );
  INV_X1 U17739 ( .A(n15676), .ZN(n20430) );
  AOI22_X1 U17740 ( .A1(\mem[709][4] ), .A2(n15672), .B1(n26421), .B2(
        data_in[4]), .ZN(n15676) );
  INV_X1 U17741 ( .A(n15677), .ZN(n20429) );
  AOI22_X1 U17742 ( .A1(\mem[709][5] ), .A2(n15672), .B1(n26421), .B2(
        data_in[5]), .ZN(n15677) );
  INV_X1 U17743 ( .A(n15678), .ZN(n20428) );
  AOI22_X1 U17744 ( .A1(\mem[709][6] ), .A2(n15672), .B1(n26421), .B2(
        data_in[6]), .ZN(n15678) );
  INV_X1 U17745 ( .A(n15679), .ZN(n20427) );
  AOI22_X1 U17746 ( .A1(\mem[709][7] ), .A2(n15672), .B1(n26421), .B2(
        data_in[7]), .ZN(n15679) );
  INV_X1 U17747 ( .A(n15680), .ZN(n20426) );
  AOI22_X1 U17748 ( .A1(\mem[710][0] ), .A2(n15681), .B1(n26420), .B2(
        data_in[0]), .ZN(n15680) );
  INV_X1 U17749 ( .A(n15682), .ZN(n20425) );
  AOI22_X1 U17750 ( .A1(\mem[710][1] ), .A2(n15681), .B1(n26420), .B2(
        data_in[1]), .ZN(n15682) );
  INV_X1 U17751 ( .A(n15683), .ZN(n20424) );
  AOI22_X1 U17752 ( .A1(\mem[710][2] ), .A2(n15681), .B1(n26420), .B2(
        data_in[2]), .ZN(n15683) );
  INV_X1 U17753 ( .A(n15684), .ZN(n20423) );
  AOI22_X1 U17754 ( .A1(\mem[710][3] ), .A2(n15681), .B1(n26420), .B2(
        data_in[3]), .ZN(n15684) );
  INV_X1 U17755 ( .A(n15685), .ZN(n20422) );
  AOI22_X1 U17756 ( .A1(\mem[710][4] ), .A2(n15681), .B1(n26420), .B2(
        data_in[4]), .ZN(n15685) );
  INV_X1 U17757 ( .A(n15686), .ZN(n20421) );
  AOI22_X1 U17758 ( .A1(\mem[710][5] ), .A2(n15681), .B1(n26420), .B2(
        data_in[5]), .ZN(n15686) );
  INV_X1 U17759 ( .A(n15687), .ZN(n20420) );
  AOI22_X1 U17760 ( .A1(\mem[710][6] ), .A2(n15681), .B1(n26420), .B2(
        data_in[6]), .ZN(n15687) );
  INV_X1 U17761 ( .A(n15688), .ZN(n20419) );
  AOI22_X1 U17762 ( .A1(\mem[710][7] ), .A2(n15681), .B1(n26420), .B2(
        data_in[7]), .ZN(n15688) );
  INV_X1 U17763 ( .A(n15689), .ZN(n20418) );
  AOI22_X1 U17764 ( .A1(\mem[711][0] ), .A2(n15690), .B1(n26419), .B2(
        data_in[0]), .ZN(n15689) );
  INV_X1 U17765 ( .A(n15691), .ZN(n20417) );
  AOI22_X1 U17766 ( .A1(\mem[711][1] ), .A2(n15690), .B1(n26419), .B2(
        data_in[1]), .ZN(n15691) );
  INV_X1 U17767 ( .A(n15692), .ZN(n20416) );
  AOI22_X1 U17768 ( .A1(\mem[711][2] ), .A2(n15690), .B1(n26419), .B2(
        data_in[2]), .ZN(n15692) );
  INV_X1 U17769 ( .A(n15693), .ZN(n20415) );
  AOI22_X1 U17770 ( .A1(\mem[711][3] ), .A2(n15690), .B1(n26419), .B2(
        data_in[3]), .ZN(n15693) );
  INV_X1 U17771 ( .A(n15694), .ZN(n20414) );
  AOI22_X1 U17772 ( .A1(\mem[711][4] ), .A2(n15690), .B1(n26419), .B2(
        data_in[4]), .ZN(n15694) );
  INV_X1 U17773 ( .A(n15695), .ZN(n20413) );
  AOI22_X1 U17774 ( .A1(\mem[711][5] ), .A2(n15690), .B1(n26419), .B2(
        data_in[5]), .ZN(n15695) );
  INV_X1 U17775 ( .A(n15696), .ZN(n20412) );
  AOI22_X1 U17776 ( .A1(\mem[711][6] ), .A2(n15690), .B1(n26419), .B2(
        data_in[6]), .ZN(n15696) );
  INV_X1 U17777 ( .A(n15697), .ZN(n20411) );
  AOI22_X1 U17778 ( .A1(\mem[711][7] ), .A2(n15690), .B1(n26419), .B2(
        data_in[7]), .ZN(n15697) );
  INV_X1 U17779 ( .A(n15914), .ZN(n20218) );
  AOI22_X1 U17780 ( .A1(\mem[736][0] ), .A2(n15915), .B1(n26394), .B2(
        data_in[0]), .ZN(n15914) );
  INV_X1 U17781 ( .A(n15916), .ZN(n20217) );
  AOI22_X1 U17782 ( .A1(\mem[736][1] ), .A2(n15915), .B1(n26394), .B2(
        data_in[1]), .ZN(n15916) );
  INV_X1 U17783 ( .A(n15917), .ZN(n20216) );
  AOI22_X1 U17784 ( .A1(\mem[736][2] ), .A2(n15915), .B1(n26394), .B2(
        data_in[2]), .ZN(n15917) );
  INV_X1 U17785 ( .A(n15918), .ZN(n20215) );
  AOI22_X1 U17786 ( .A1(\mem[736][3] ), .A2(n15915), .B1(n26394), .B2(
        data_in[3]), .ZN(n15918) );
  INV_X1 U17787 ( .A(n15919), .ZN(n20214) );
  AOI22_X1 U17788 ( .A1(\mem[736][4] ), .A2(n15915), .B1(n26394), .B2(
        data_in[4]), .ZN(n15919) );
  INV_X1 U17789 ( .A(n15920), .ZN(n20213) );
  AOI22_X1 U17790 ( .A1(\mem[736][5] ), .A2(n15915), .B1(n26394), .B2(
        data_in[5]), .ZN(n15920) );
  INV_X1 U17791 ( .A(n15921), .ZN(n20212) );
  AOI22_X1 U17792 ( .A1(\mem[736][6] ), .A2(n15915), .B1(n26394), .B2(
        data_in[6]), .ZN(n15921) );
  INV_X1 U17793 ( .A(n15922), .ZN(n20211) );
  AOI22_X1 U17794 ( .A1(\mem[736][7] ), .A2(n15915), .B1(n26394), .B2(
        data_in[7]), .ZN(n15922) );
  INV_X1 U17795 ( .A(n15924), .ZN(n20210) );
  AOI22_X1 U17796 ( .A1(\mem[737][0] ), .A2(n15925), .B1(n26393), .B2(
        data_in[0]), .ZN(n15924) );
  INV_X1 U17797 ( .A(n15926), .ZN(n20209) );
  AOI22_X1 U17798 ( .A1(\mem[737][1] ), .A2(n15925), .B1(n26393), .B2(
        data_in[1]), .ZN(n15926) );
  INV_X1 U17799 ( .A(n15927), .ZN(n20208) );
  AOI22_X1 U17800 ( .A1(\mem[737][2] ), .A2(n15925), .B1(n26393), .B2(
        data_in[2]), .ZN(n15927) );
  INV_X1 U17801 ( .A(n15928), .ZN(n20207) );
  AOI22_X1 U17802 ( .A1(\mem[737][3] ), .A2(n15925), .B1(n26393), .B2(
        data_in[3]), .ZN(n15928) );
  INV_X1 U17803 ( .A(n15929), .ZN(n20206) );
  AOI22_X1 U17804 ( .A1(\mem[737][4] ), .A2(n15925), .B1(n26393), .B2(
        data_in[4]), .ZN(n15929) );
  INV_X1 U17805 ( .A(n15930), .ZN(n20205) );
  AOI22_X1 U17806 ( .A1(\mem[737][5] ), .A2(n15925), .B1(n26393), .B2(
        data_in[5]), .ZN(n15930) );
  INV_X1 U17807 ( .A(n15931), .ZN(n20204) );
  AOI22_X1 U17808 ( .A1(\mem[737][6] ), .A2(n15925), .B1(n26393), .B2(
        data_in[6]), .ZN(n15931) );
  INV_X1 U17809 ( .A(n15932), .ZN(n20203) );
  AOI22_X1 U17810 ( .A1(\mem[737][7] ), .A2(n15925), .B1(n26393), .B2(
        data_in[7]), .ZN(n15932) );
  INV_X1 U17811 ( .A(n15933), .ZN(n20202) );
  AOI22_X1 U17812 ( .A1(\mem[738][0] ), .A2(n15934), .B1(n26392), .B2(
        data_in[0]), .ZN(n15933) );
  INV_X1 U17813 ( .A(n15935), .ZN(n20201) );
  AOI22_X1 U17814 ( .A1(\mem[738][1] ), .A2(n15934), .B1(n26392), .B2(
        data_in[1]), .ZN(n15935) );
  INV_X1 U17815 ( .A(n15936), .ZN(n20200) );
  AOI22_X1 U17816 ( .A1(\mem[738][2] ), .A2(n15934), .B1(n26392), .B2(
        data_in[2]), .ZN(n15936) );
  INV_X1 U17817 ( .A(n15937), .ZN(n20199) );
  AOI22_X1 U17818 ( .A1(\mem[738][3] ), .A2(n15934), .B1(n26392), .B2(
        data_in[3]), .ZN(n15937) );
  INV_X1 U17819 ( .A(n15938), .ZN(n20198) );
  AOI22_X1 U17820 ( .A1(\mem[738][4] ), .A2(n15934), .B1(n26392), .B2(
        data_in[4]), .ZN(n15938) );
  INV_X1 U17821 ( .A(n15939), .ZN(n20197) );
  AOI22_X1 U17822 ( .A1(\mem[738][5] ), .A2(n15934), .B1(n26392), .B2(
        data_in[5]), .ZN(n15939) );
  INV_X1 U17823 ( .A(n15940), .ZN(n20196) );
  AOI22_X1 U17824 ( .A1(\mem[738][6] ), .A2(n15934), .B1(n26392), .B2(
        data_in[6]), .ZN(n15940) );
  INV_X1 U17825 ( .A(n15941), .ZN(n20195) );
  AOI22_X1 U17826 ( .A1(\mem[738][7] ), .A2(n15934), .B1(n26392), .B2(
        data_in[7]), .ZN(n15941) );
  INV_X1 U17827 ( .A(n15942), .ZN(n20194) );
  AOI22_X1 U17828 ( .A1(\mem[739][0] ), .A2(n15943), .B1(n26391), .B2(
        data_in[0]), .ZN(n15942) );
  INV_X1 U17829 ( .A(n15944), .ZN(n20193) );
  AOI22_X1 U17830 ( .A1(\mem[739][1] ), .A2(n15943), .B1(n26391), .B2(
        data_in[1]), .ZN(n15944) );
  INV_X1 U17831 ( .A(n15945), .ZN(n20192) );
  AOI22_X1 U17832 ( .A1(\mem[739][2] ), .A2(n15943), .B1(n26391), .B2(
        data_in[2]), .ZN(n15945) );
  INV_X1 U17833 ( .A(n15946), .ZN(n20191) );
  AOI22_X1 U17834 ( .A1(\mem[739][3] ), .A2(n15943), .B1(n26391), .B2(
        data_in[3]), .ZN(n15946) );
  INV_X1 U17835 ( .A(n15947), .ZN(n20190) );
  AOI22_X1 U17836 ( .A1(\mem[739][4] ), .A2(n15943), .B1(n26391), .B2(
        data_in[4]), .ZN(n15947) );
  INV_X1 U17837 ( .A(n15948), .ZN(n20189) );
  AOI22_X1 U17838 ( .A1(\mem[739][5] ), .A2(n15943), .B1(n26391), .B2(
        data_in[5]), .ZN(n15948) );
  INV_X1 U17839 ( .A(n15949), .ZN(n20188) );
  AOI22_X1 U17840 ( .A1(\mem[739][6] ), .A2(n15943), .B1(n26391), .B2(
        data_in[6]), .ZN(n15949) );
  INV_X1 U17841 ( .A(n15950), .ZN(n20187) );
  AOI22_X1 U17842 ( .A1(\mem[739][7] ), .A2(n15943), .B1(n26391), .B2(
        data_in[7]), .ZN(n15950) );
  INV_X1 U17843 ( .A(n15951), .ZN(n20186) );
  AOI22_X1 U17844 ( .A1(\mem[740][0] ), .A2(n15952), .B1(n26390), .B2(
        data_in[0]), .ZN(n15951) );
  INV_X1 U17845 ( .A(n15953), .ZN(n20185) );
  AOI22_X1 U17846 ( .A1(\mem[740][1] ), .A2(n15952), .B1(n26390), .B2(
        data_in[1]), .ZN(n15953) );
  INV_X1 U17847 ( .A(n15954), .ZN(n20184) );
  AOI22_X1 U17848 ( .A1(\mem[740][2] ), .A2(n15952), .B1(n26390), .B2(
        data_in[2]), .ZN(n15954) );
  INV_X1 U17849 ( .A(n15955), .ZN(n20183) );
  AOI22_X1 U17850 ( .A1(\mem[740][3] ), .A2(n15952), .B1(n26390), .B2(
        data_in[3]), .ZN(n15955) );
  INV_X1 U17851 ( .A(n15956), .ZN(n20182) );
  AOI22_X1 U17852 ( .A1(\mem[740][4] ), .A2(n15952), .B1(n26390), .B2(
        data_in[4]), .ZN(n15956) );
  INV_X1 U17853 ( .A(n15957), .ZN(n20181) );
  AOI22_X1 U17854 ( .A1(\mem[740][5] ), .A2(n15952), .B1(n26390), .B2(
        data_in[5]), .ZN(n15957) );
  INV_X1 U17855 ( .A(n15958), .ZN(n20180) );
  AOI22_X1 U17856 ( .A1(\mem[740][6] ), .A2(n15952), .B1(n26390), .B2(
        data_in[6]), .ZN(n15958) );
  INV_X1 U17857 ( .A(n15959), .ZN(n20179) );
  AOI22_X1 U17858 ( .A1(\mem[740][7] ), .A2(n15952), .B1(n26390), .B2(
        data_in[7]), .ZN(n15959) );
  INV_X1 U17859 ( .A(n15960), .ZN(n20178) );
  AOI22_X1 U17860 ( .A1(\mem[741][0] ), .A2(n15961), .B1(n26389), .B2(
        data_in[0]), .ZN(n15960) );
  INV_X1 U17861 ( .A(n15962), .ZN(n20177) );
  AOI22_X1 U17862 ( .A1(\mem[741][1] ), .A2(n15961), .B1(n26389), .B2(
        data_in[1]), .ZN(n15962) );
  INV_X1 U17863 ( .A(n15963), .ZN(n20176) );
  AOI22_X1 U17864 ( .A1(\mem[741][2] ), .A2(n15961), .B1(n26389), .B2(
        data_in[2]), .ZN(n15963) );
  INV_X1 U17865 ( .A(n15964), .ZN(n20175) );
  AOI22_X1 U17866 ( .A1(\mem[741][3] ), .A2(n15961), .B1(n26389), .B2(
        data_in[3]), .ZN(n15964) );
  INV_X1 U17867 ( .A(n15965), .ZN(n20174) );
  AOI22_X1 U17868 ( .A1(\mem[741][4] ), .A2(n15961), .B1(n26389), .B2(
        data_in[4]), .ZN(n15965) );
  INV_X1 U17869 ( .A(n15966), .ZN(n20173) );
  AOI22_X1 U17870 ( .A1(\mem[741][5] ), .A2(n15961), .B1(n26389), .B2(
        data_in[5]), .ZN(n15966) );
  INV_X1 U17871 ( .A(n15967), .ZN(n20172) );
  AOI22_X1 U17872 ( .A1(\mem[741][6] ), .A2(n15961), .B1(n26389), .B2(
        data_in[6]), .ZN(n15967) );
  INV_X1 U17873 ( .A(n15968), .ZN(n20171) );
  AOI22_X1 U17874 ( .A1(\mem[741][7] ), .A2(n15961), .B1(n26389), .B2(
        data_in[7]), .ZN(n15968) );
  INV_X1 U17875 ( .A(n15969), .ZN(n20170) );
  AOI22_X1 U17876 ( .A1(\mem[742][0] ), .A2(n15970), .B1(n26388), .B2(
        data_in[0]), .ZN(n15969) );
  INV_X1 U17877 ( .A(n15971), .ZN(n20169) );
  AOI22_X1 U17878 ( .A1(\mem[742][1] ), .A2(n15970), .B1(n26388), .B2(
        data_in[1]), .ZN(n15971) );
  INV_X1 U17879 ( .A(n15972), .ZN(n20168) );
  AOI22_X1 U17880 ( .A1(\mem[742][2] ), .A2(n15970), .B1(n26388), .B2(
        data_in[2]), .ZN(n15972) );
  INV_X1 U17881 ( .A(n15973), .ZN(n20167) );
  AOI22_X1 U17882 ( .A1(\mem[742][3] ), .A2(n15970), .B1(n26388), .B2(
        data_in[3]), .ZN(n15973) );
  INV_X1 U17883 ( .A(n15974), .ZN(n20166) );
  AOI22_X1 U17884 ( .A1(\mem[742][4] ), .A2(n15970), .B1(n26388), .B2(
        data_in[4]), .ZN(n15974) );
  INV_X1 U17885 ( .A(n15975), .ZN(n20165) );
  AOI22_X1 U17886 ( .A1(\mem[742][5] ), .A2(n15970), .B1(n26388), .B2(
        data_in[5]), .ZN(n15975) );
  INV_X1 U17887 ( .A(n15976), .ZN(n20164) );
  AOI22_X1 U17888 ( .A1(\mem[742][6] ), .A2(n15970), .B1(n26388), .B2(
        data_in[6]), .ZN(n15976) );
  INV_X1 U17889 ( .A(n15977), .ZN(n20163) );
  AOI22_X1 U17890 ( .A1(\mem[742][7] ), .A2(n15970), .B1(n26388), .B2(
        data_in[7]), .ZN(n15977) );
  INV_X1 U17891 ( .A(n15978), .ZN(n20162) );
  AOI22_X1 U17892 ( .A1(\mem[743][0] ), .A2(n15979), .B1(n26387), .B2(
        data_in[0]), .ZN(n15978) );
  INV_X1 U17893 ( .A(n15980), .ZN(n20161) );
  AOI22_X1 U17894 ( .A1(\mem[743][1] ), .A2(n15979), .B1(n26387), .B2(
        data_in[1]), .ZN(n15980) );
  INV_X1 U17895 ( .A(n15981), .ZN(n20160) );
  AOI22_X1 U17896 ( .A1(\mem[743][2] ), .A2(n15979), .B1(n26387), .B2(
        data_in[2]), .ZN(n15981) );
  INV_X1 U17897 ( .A(n15982), .ZN(n20159) );
  AOI22_X1 U17898 ( .A1(\mem[743][3] ), .A2(n15979), .B1(n26387), .B2(
        data_in[3]), .ZN(n15982) );
  INV_X1 U17899 ( .A(n15983), .ZN(n20158) );
  AOI22_X1 U17900 ( .A1(\mem[743][4] ), .A2(n15979), .B1(n26387), .B2(
        data_in[4]), .ZN(n15983) );
  INV_X1 U17901 ( .A(n15984), .ZN(n20157) );
  AOI22_X1 U17902 ( .A1(\mem[743][5] ), .A2(n15979), .B1(n26387), .B2(
        data_in[5]), .ZN(n15984) );
  INV_X1 U17903 ( .A(n15985), .ZN(n20156) );
  AOI22_X1 U17904 ( .A1(\mem[743][6] ), .A2(n15979), .B1(n26387), .B2(
        data_in[6]), .ZN(n15985) );
  INV_X1 U17905 ( .A(n15986), .ZN(n20155) );
  AOI22_X1 U17906 ( .A1(\mem[743][7] ), .A2(n15979), .B1(n26387), .B2(
        data_in[7]), .ZN(n15986) );
  INV_X1 U17907 ( .A(n16203), .ZN(n19962) );
  AOI22_X1 U17908 ( .A1(\mem[768][0] ), .A2(n16204), .B1(n26362), .B2(
        data_in[0]), .ZN(n16203) );
  INV_X1 U17909 ( .A(n16205), .ZN(n19961) );
  AOI22_X1 U17910 ( .A1(\mem[768][1] ), .A2(n16204), .B1(n26362), .B2(
        data_in[1]), .ZN(n16205) );
  INV_X1 U17911 ( .A(n16206), .ZN(n19960) );
  AOI22_X1 U17912 ( .A1(\mem[768][2] ), .A2(n16204), .B1(n26362), .B2(
        data_in[2]), .ZN(n16206) );
  INV_X1 U17913 ( .A(n16207), .ZN(n19959) );
  AOI22_X1 U17914 ( .A1(\mem[768][3] ), .A2(n16204), .B1(n26362), .B2(
        data_in[3]), .ZN(n16207) );
  INV_X1 U17915 ( .A(n16208), .ZN(n19958) );
  AOI22_X1 U17916 ( .A1(\mem[768][4] ), .A2(n16204), .B1(n26362), .B2(
        data_in[4]), .ZN(n16208) );
  INV_X1 U17917 ( .A(n16209), .ZN(n19957) );
  AOI22_X1 U17918 ( .A1(\mem[768][5] ), .A2(n16204), .B1(n26362), .B2(
        data_in[5]), .ZN(n16209) );
  INV_X1 U17919 ( .A(n16210), .ZN(n19956) );
  AOI22_X1 U17920 ( .A1(\mem[768][6] ), .A2(n16204), .B1(n26362), .B2(
        data_in[6]), .ZN(n16210) );
  INV_X1 U17921 ( .A(n16211), .ZN(n19955) );
  AOI22_X1 U17922 ( .A1(\mem[768][7] ), .A2(n16204), .B1(n26362), .B2(
        data_in[7]), .ZN(n16211) );
  INV_X1 U17923 ( .A(n16213), .ZN(n19954) );
  AOI22_X1 U17924 ( .A1(\mem[769][0] ), .A2(n16214), .B1(n26361), .B2(
        data_in[0]), .ZN(n16213) );
  INV_X1 U17925 ( .A(n16215), .ZN(n19953) );
  AOI22_X1 U17926 ( .A1(\mem[769][1] ), .A2(n16214), .B1(n26361), .B2(
        data_in[1]), .ZN(n16215) );
  INV_X1 U17927 ( .A(n16216), .ZN(n19952) );
  AOI22_X1 U17928 ( .A1(\mem[769][2] ), .A2(n16214), .B1(n26361), .B2(
        data_in[2]), .ZN(n16216) );
  INV_X1 U17929 ( .A(n16217), .ZN(n19951) );
  AOI22_X1 U17930 ( .A1(\mem[769][3] ), .A2(n16214), .B1(n26361), .B2(
        data_in[3]), .ZN(n16217) );
  INV_X1 U17931 ( .A(n16218), .ZN(n19950) );
  AOI22_X1 U17932 ( .A1(\mem[769][4] ), .A2(n16214), .B1(n26361), .B2(
        data_in[4]), .ZN(n16218) );
  INV_X1 U17933 ( .A(n16219), .ZN(n19949) );
  AOI22_X1 U17934 ( .A1(\mem[769][5] ), .A2(n16214), .B1(n26361), .B2(
        data_in[5]), .ZN(n16219) );
  INV_X1 U17935 ( .A(n16220), .ZN(n19948) );
  AOI22_X1 U17936 ( .A1(\mem[769][6] ), .A2(n16214), .B1(n26361), .B2(
        data_in[6]), .ZN(n16220) );
  INV_X1 U17937 ( .A(n16221), .ZN(n19947) );
  AOI22_X1 U17938 ( .A1(\mem[769][7] ), .A2(n16214), .B1(n26361), .B2(
        data_in[7]), .ZN(n16221) );
  INV_X1 U17939 ( .A(n16222), .ZN(n19946) );
  AOI22_X1 U17940 ( .A1(\mem[770][0] ), .A2(n16223), .B1(n26360), .B2(
        data_in[0]), .ZN(n16222) );
  INV_X1 U17941 ( .A(n16224), .ZN(n19945) );
  AOI22_X1 U17942 ( .A1(\mem[770][1] ), .A2(n16223), .B1(n26360), .B2(
        data_in[1]), .ZN(n16224) );
  INV_X1 U17943 ( .A(n16225), .ZN(n19944) );
  AOI22_X1 U17944 ( .A1(\mem[770][2] ), .A2(n16223), .B1(n26360), .B2(
        data_in[2]), .ZN(n16225) );
  INV_X1 U17945 ( .A(n16226), .ZN(n19943) );
  AOI22_X1 U17946 ( .A1(\mem[770][3] ), .A2(n16223), .B1(n26360), .B2(
        data_in[3]), .ZN(n16226) );
  INV_X1 U17947 ( .A(n16227), .ZN(n19942) );
  AOI22_X1 U17948 ( .A1(\mem[770][4] ), .A2(n16223), .B1(n26360), .B2(
        data_in[4]), .ZN(n16227) );
  INV_X1 U17949 ( .A(n16228), .ZN(n19941) );
  AOI22_X1 U17950 ( .A1(\mem[770][5] ), .A2(n16223), .B1(n26360), .B2(
        data_in[5]), .ZN(n16228) );
  INV_X1 U17951 ( .A(n16229), .ZN(n19940) );
  AOI22_X1 U17952 ( .A1(\mem[770][6] ), .A2(n16223), .B1(n26360), .B2(
        data_in[6]), .ZN(n16229) );
  INV_X1 U17953 ( .A(n16230), .ZN(n19939) );
  AOI22_X1 U17954 ( .A1(\mem[770][7] ), .A2(n16223), .B1(n26360), .B2(
        data_in[7]), .ZN(n16230) );
  INV_X1 U17955 ( .A(n16231), .ZN(n19938) );
  AOI22_X1 U17956 ( .A1(\mem[771][0] ), .A2(n16232), .B1(n26359), .B2(
        data_in[0]), .ZN(n16231) );
  INV_X1 U17957 ( .A(n16233), .ZN(n19937) );
  AOI22_X1 U17958 ( .A1(\mem[771][1] ), .A2(n16232), .B1(n26359), .B2(
        data_in[1]), .ZN(n16233) );
  INV_X1 U17959 ( .A(n16234), .ZN(n19936) );
  AOI22_X1 U17960 ( .A1(\mem[771][2] ), .A2(n16232), .B1(n26359), .B2(
        data_in[2]), .ZN(n16234) );
  INV_X1 U17961 ( .A(n16235), .ZN(n19935) );
  AOI22_X1 U17962 ( .A1(\mem[771][3] ), .A2(n16232), .B1(n26359), .B2(
        data_in[3]), .ZN(n16235) );
  INV_X1 U17963 ( .A(n16236), .ZN(n19934) );
  AOI22_X1 U17964 ( .A1(\mem[771][4] ), .A2(n16232), .B1(n26359), .B2(
        data_in[4]), .ZN(n16236) );
  INV_X1 U17965 ( .A(n16237), .ZN(n19933) );
  AOI22_X1 U17966 ( .A1(\mem[771][5] ), .A2(n16232), .B1(n26359), .B2(
        data_in[5]), .ZN(n16237) );
  INV_X1 U17967 ( .A(n16238), .ZN(n19932) );
  AOI22_X1 U17968 ( .A1(\mem[771][6] ), .A2(n16232), .B1(n26359), .B2(
        data_in[6]), .ZN(n16238) );
  INV_X1 U17969 ( .A(n16239), .ZN(n19931) );
  AOI22_X1 U17970 ( .A1(\mem[771][7] ), .A2(n16232), .B1(n26359), .B2(
        data_in[7]), .ZN(n16239) );
  INV_X1 U17971 ( .A(n16240), .ZN(n19930) );
  AOI22_X1 U17972 ( .A1(\mem[772][0] ), .A2(n16241), .B1(n26358), .B2(
        data_in[0]), .ZN(n16240) );
  INV_X1 U17973 ( .A(n16242), .ZN(n19929) );
  AOI22_X1 U17974 ( .A1(\mem[772][1] ), .A2(n16241), .B1(n26358), .B2(
        data_in[1]), .ZN(n16242) );
  INV_X1 U17975 ( .A(n16243), .ZN(n19928) );
  AOI22_X1 U17976 ( .A1(\mem[772][2] ), .A2(n16241), .B1(n26358), .B2(
        data_in[2]), .ZN(n16243) );
  INV_X1 U17977 ( .A(n16244), .ZN(n19927) );
  AOI22_X1 U17978 ( .A1(\mem[772][3] ), .A2(n16241), .B1(n26358), .B2(
        data_in[3]), .ZN(n16244) );
  INV_X1 U17979 ( .A(n16245), .ZN(n19926) );
  AOI22_X1 U17980 ( .A1(\mem[772][4] ), .A2(n16241), .B1(n26358), .B2(
        data_in[4]), .ZN(n16245) );
  INV_X1 U17981 ( .A(n16246), .ZN(n19925) );
  AOI22_X1 U17982 ( .A1(\mem[772][5] ), .A2(n16241), .B1(n26358), .B2(
        data_in[5]), .ZN(n16246) );
  INV_X1 U17983 ( .A(n16247), .ZN(n19924) );
  AOI22_X1 U17984 ( .A1(\mem[772][6] ), .A2(n16241), .B1(n26358), .B2(
        data_in[6]), .ZN(n16247) );
  INV_X1 U17985 ( .A(n16248), .ZN(n19923) );
  AOI22_X1 U17986 ( .A1(\mem[772][7] ), .A2(n16241), .B1(n26358), .B2(
        data_in[7]), .ZN(n16248) );
  INV_X1 U17987 ( .A(n16249), .ZN(n19922) );
  AOI22_X1 U17988 ( .A1(\mem[773][0] ), .A2(n16250), .B1(n26357), .B2(
        data_in[0]), .ZN(n16249) );
  INV_X1 U17989 ( .A(n16251), .ZN(n19921) );
  AOI22_X1 U17990 ( .A1(\mem[773][1] ), .A2(n16250), .B1(n26357), .B2(
        data_in[1]), .ZN(n16251) );
  INV_X1 U17991 ( .A(n16252), .ZN(n19920) );
  AOI22_X1 U17992 ( .A1(\mem[773][2] ), .A2(n16250), .B1(n26357), .B2(
        data_in[2]), .ZN(n16252) );
  INV_X1 U17993 ( .A(n16253), .ZN(n19919) );
  AOI22_X1 U17994 ( .A1(\mem[773][3] ), .A2(n16250), .B1(n26357), .B2(
        data_in[3]), .ZN(n16253) );
  INV_X1 U17995 ( .A(n16254), .ZN(n19918) );
  AOI22_X1 U17996 ( .A1(\mem[773][4] ), .A2(n16250), .B1(n26357), .B2(
        data_in[4]), .ZN(n16254) );
  INV_X1 U17997 ( .A(n16255), .ZN(n19917) );
  AOI22_X1 U17998 ( .A1(\mem[773][5] ), .A2(n16250), .B1(n26357), .B2(
        data_in[5]), .ZN(n16255) );
  INV_X1 U17999 ( .A(n16256), .ZN(n19916) );
  AOI22_X1 U18000 ( .A1(\mem[773][6] ), .A2(n16250), .B1(n26357), .B2(
        data_in[6]), .ZN(n16256) );
  INV_X1 U18001 ( .A(n16257), .ZN(n19915) );
  AOI22_X1 U18002 ( .A1(\mem[773][7] ), .A2(n16250), .B1(n26357), .B2(
        data_in[7]), .ZN(n16257) );
  INV_X1 U18003 ( .A(n16258), .ZN(n19914) );
  AOI22_X1 U18004 ( .A1(\mem[774][0] ), .A2(n16259), .B1(n26356), .B2(
        data_in[0]), .ZN(n16258) );
  INV_X1 U18005 ( .A(n16260), .ZN(n19913) );
  AOI22_X1 U18006 ( .A1(\mem[774][1] ), .A2(n16259), .B1(n26356), .B2(
        data_in[1]), .ZN(n16260) );
  INV_X1 U18007 ( .A(n16261), .ZN(n19912) );
  AOI22_X1 U18008 ( .A1(\mem[774][2] ), .A2(n16259), .B1(n26356), .B2(
        data_in[2]), .ZN(n16261) );
  INV_X1 U18009 ( .A(n16262), .ZN(n19911) );
  AOI22_X1 U18010 ( .A1(\mem[774][3] ), .A2(n16259), .B1(n26356), .B2(
        data_in[3]), .ZN(n16262) );
  INV_X1 U18011 ( .A(n16263), .ZN(n19910) );
  AOI22_X1 U18012 ( .A1(\mem[774][4] ), .A2(n16259), .B1(n26356), .B2(
        data_in[4]), .ZN(n16263) );
  INV_X1 U18013 ( .A(n16264), .ZN(n19909) );
  AOI22_X1 U18014 ( .A1(\mem[774][5] ), .A2(n16259), .B1(n26356), .B2(
        data_in[5]), .ZN(n16264) );
  INV_X1 U18015 ( .A(n16265), .ZN(n19908) );
  AOI22_X1 U18016 ( .A1(\mem[774][6] ), .A2(n16259), .B1(n26356), .B2(
        data_in[6]), .ZN(n16265) );
  INV_X1 U18017 ( .A(n16266), .ZN(n19907) );
  AOI22_X1 U18018 ( .A1(\mem[774][7] ), .A2(n16259), .B1(n26356), .B2(
        data_in[7]), .ZN(n16266) );
  INV_X1 U18019 ( .A(n16267), .ZN(n19906) );
  AOI22_X1 U18020 ( .A1(\mem[775][0] ), .A2(n16268), .B1(n26355), .B2(
        data_in[0]), .ZN(n16267) );
  INV_X1 U18021 ( .A(n16269), .ZN(n19905) );
  AOI22_X1 U18022 ( .A1(\mem[775][1] ), .A2(n16268), .B1(n26355), .B2(
        data_in[1]), .ZN(n16269) );
  INV_X1 U18023 ( .A(n16270), .ZN(n19904) );
  AOI22_X1 U18024 ( .A1(\mem[775][2] ), .A2(n16268), .B1(n26355), .B2(
        data_in[2]), .ZN(n16270) );
  INV_X1 U18025 ( .A(n16271), .ZN(n19903) );
  AOI22_X1 U18026 ( .A1(\mem[775][3] ), .A2(n16268), .B1(n26355), .B2(
        data_in[3]), .ZN(n16271) );
  INV_X1 U18027 ( .A(n16272), .ZN(n19902) );
  AOI22_X1 U18028 ( .A1(\mem[775][4] ), .A2(n16268), .B1(n26355), .B2(
        data_in[4]), .ZN(n16272) );
  INV_X1 U18029 ( .A(n16273), .ZN(n19901) );
  AOI22_X1 U18030 ( .A1(\mem[775][5] ), .A2(n16268), .B1(n26355), .B2(
        data_in[5]), .ZN(n16273) );
  INV_X1 U18031 ( .A(n16274), .ZN(n19900) );
  AOI22_X1 U18032 ( .A1(\mem[775][6] ), .A2(n16268), .B1(n26355), .B2(
        data_in[6]), .ZN(n16274) );
  INV_X1 U18033 ( .A(n16275), .ZN(n19899) );
  AOI22_X1 U18034 ( .A1(\mem[775][7] ), .A2(n16268), .B1(n26355), .B2(
        data_in[7]), .ZN(n16275) );
  INV_X1 U18035 ( .A(n16493), .ZN(n19706) );
  AOI22_X1 U18036 ( .A1(\mem[800][0] ), .A2(n16494), .B1(n26330), .B2(
        data_in[0]), .ZN(n16493) );
  INV_X1 U18037 ( .A(n16495), .ZN(n19705) );
  AOI22_X1 U18038 ( .A1(\mem[800][1] ), .A2(n16494), .B1(n26330), .B2(
        data_in[1]), .ZN(n16495) );
  INV_X1 U18039 ( .A(n16496), .ZN(n19704) );
  AOI22_X1 U18040 ( .A1(\mem[800][2] ), .A2(n16494), .B1(n26330), .B2(
        data_in[2]), .ZN(n16496) );
  INV_X1 U18041 ( .A(n16497), .ZN(n19703) );
  AOI22_X1 U18042 ( .A1(\mem[800][3] ), .A2(n16494), .B1(n26330), .B2(
        data_in[3]), .ZN(n16497) );
  INV_X1 U18043 ( .A(n16498), .ZN(n19702) );
  AOI22_X1 U18044 ( .A1(\mem[800][4] ), .A2(n16494), .B1(n26330), .B2(
        data_in[4]), .ZN(n16498) );
  INV_X1 U18045 ( .A(n16499), .ZN(n19701) );
  AOI22_X1 U18046 ( .A1(\mem[800][5] ), .A2(n16494), .B1(n26330), .B2(
        data_in[5]), .ZN(n16499) );
  INV_X1 U18047 ( .A(n16500), .ZN(n19700) );
  AOI22_X1 U18048 ( .A1(\mem[800][6] ), .A2(n16494), .B1(n26330), .B2(
        data_in[6]), .ZN(n16500) );
  INV_X1 U18049 ( .A(n16501), .ZN(n19699) );
  AOI22_X1 U18050 ( .A1(\mem[800][7] ), .A2(n16494), .B1(n26330), .B2(
        data_in[7]), .ZN(n16501) );
  INV_X1 U18051 ( .A(n16503), .ZN(n19698) );
  AOI22_X1 U18052 ( .A1(\mem[801][0] ), .A2(n16504), .B1(n26329), .B2(
        data_in[0]), .ZN(n16503) );
  INV_X1 U18053 ( .A(n16505), .ZN(n19697) );
  AOI22_X1 U18054 ( .A1(\mem[801][1] ), .A2(n16504), .B1(n26329), .B2(
        data_in[1]), .ZN(n16505) );
  INV_X1 U18055 ( .A(n16506), .ZN(n19696) );
  AOI22_X1 U18056 ( .A1(\mem[801][2] ), .A2(n16504), .B1(n26329), .B2(
        data_in[2]), .ZN(n16506) );
  INV_X1 U18057 ( .A(n16507), .ZN(n19695) );
  AOI22_X1 U18058 ( .A1(\mem[801][3] ), .A2(n16504), .B1(n26329), .B2(
        data_in[3]), .ZN(n16507) );
  INV_X1 U18059 ( .A(n16508), .ZN(n19694) );
  AOI22_X1 U18060 ( .A1(\mem[801][4] ), .A2(n16504), .B1(n26329), .B2(
        data_in[4]), .ZN(n16508) );
  INV_X1 U18061 ( .A(n16509), .ZN(n19693) );
  AOI22_X1 U18062 ( .A1(\mem[801][5] ), .A2(n16504), .B1(n26329), .B2(
        data_in[5]), .ZN(n16509) );
  INV_X1 U18063 ( .A(n16510), .ZN(n19692) );
  AOI22_X1 U18064 ( .A1(\mem[801][6] ), .A2(n16504), .B1(n26329), .B2(
        data_in[6]), .ZN(n16510) );
  INV_X1 U18065 ( .A(n16511), .ZN(n19691) );
  AOI22_X1 U18066 ( .A1(\mem[801][7] ), .A2(n16504), .B1(n26329), .B2(
        data_in[7]), .ZN(n16511) );
  INV_X1 U18067 ( .A(n16512), .ZN(n19690) );
  AOI22_X1 U18068 ( .A1(\mem[802][0] ), .A2(n16513), .B1(n26328), .B2(
        data_in[0]), .ZN(n16512) );
  INV_X1 U18069 ( .A(n16514), .ZN(n19689) );
  AOI22_X1 U18070 ( .A1(\mem[802][1] ), .A2(n16513), .B1(n26328), .B2(
        data_in[1]), .ZN(n16514) );
  INV_X1 U18071 ( .A(n16515), .ZN(n19688) );
  AOI22_X1 U18072 ( .A1(\mem[802][2] ), .A2(n16513), .B1(n26328), .B2(
        data_in[2]), .ZN(n16515) );
  INV_X1 U18073 ( .A(n16516), .ZN(n19687) );
  AOI22_X1 U18074 ( .A1(\mem[802][3] ), .A2(n16513), .B1(n26328), .B2(
        data_in[3]), .ZN(n16516) );
  INV_X1 U18075 ( .A(n16517), .ZN(n19686) );
  AOI22_X1 U18076 ( .A1(\mem[802][4] ), .A2(n16513), .B1(n26328), .B2(
        data_in[4]), .ZN(n16517) );
  INV_X1 U18077 ( .A(n16518), .ZN(n19685) );
  AOI22_X1 U18078 ( .A1(\mem[802][5] ), .A2(n16513), .B1(n26328), .B2(
        data_in[5]), .ZN(n16518) );
  INV_X1 U18079 ( .A(n16519), .ZN(n19684) );
  AOI22_X1 U18080 ( .A1(\mem[802][6] ), .A2(n16513), .B1(n26328), .B2(
        data_in[6]), .ZN(n16519) );
  INV_X1 U18081 ( .A(n16520), .ZN(n19683) );
  AOI22_X1 U18082 ( .A1(\mem[802][7] ), .A2(n16513), .B1(n26328), .B2(
        data_in[7]), .ZN(n16520) );
  INV_X1 U18083 ( .A(n16521), .ZN(n19682) );
  AOI22_X1 U18084 ( .A1(\mem[803][0] ), .A2(n16522), .B1(n26327), .B2(
        data_in[0]), .ZN(n16521) );
  INV_X1 U18085 ( .A(n16523), .ZN(n19681) );
  AOI22_X1 U18086 ( .A1(\mem[803][1] ), .A2(n16522), .B1(n26327), .B2(
        data_in[1]), .ZN(n16523) );
  INV_X1 U18087 ( .A(n16524), .ZN(n19680) );
  AOI22_X1 U18088 ( .A1(\mem[803][2] ), .A2(n16522), .B1(n26327), .B2(
        data_in[2]), .ZN(n16524) );
  INV_X1 U18089 ( .A(n16525), .ZN(n19679) );
  AOI22_X1 U18090 ( .A1(\mem[803][3] ), .A2(n16522), .B1(n26327), .B2(
        data_in[3]), .ZN(n16525) );
  INV_X1 U18091 ( .A(n16526), .ZN(n19678) );
  AOI22_X1 U18092 ( .A1(\mem[803][4] ), .A2(n16522), .B1(n26327), .B2(
        data_in[4]), .ZN(n16526) );
  INV_X1 U18093 ( .A(n16527), .ZN(n19677) );
  AOI22_X1 U18094 ( .A1(\mem[803][5] ), .A2(n16522), .B1(n26327), .B2(
        data_in[5]), .ZN(n16527) );
  INV_X1 U18095 ( .A(n16528), .ZN(n19676) );
  AOI22_X1 U18096 ( .A1(\mem[803][6] ), .A2(n16522), .B1(n26327), .B2(
        data_in[6]), .ZN(n16528) );
  INV_X1 U18097 ( .A(n16529), .ZN(n19675) );
  AOI22_X1 U18098 ( .A1(\mem[803][7] ), .A2(n16522), .B1(n26327), .B2(
        data_in[7]), .ZN(n16529) );
  INV_X1 U18099 ( .A(n16530), .ZN(n19674) );
  AOI22_X1 U18100 ( .A1(\mem[804][0] ), .A2(n16531), .B1(n26326), .B2(
        data_in[0]), .ZN(n16530) );
  INV_X1 U18101 ( .A(n16532), .ZN(n19673) );
  AOI22_X1 U18102 ( .A1(\mem[804][1] ), .A2(n16531), .B1(n26326), .B2(
        data_in[1]), .ZN(n16532) );
  INV_X1 U18103 ( .A(n16533), .ZN(n19672) );
  AOI22_X1 U18104 ( .A1(\mem[804][2] ), .A2(n16531), .B1(n26326), .B2(
        data_in[2]), .ZN(n16533) );
  INV_X1 U18105 ( .A(n16534), .ZN(n19671) );
  AOI22_X1 U18106 ( .A1(\mem[804][3] ), .A2(n16531), .B1(n26326), .B2(
        data_in[3]), .ZN(n16534) );
  INV_X1 U18107 ( .A(n16535), .ZN(n19670) );
  AOI22_X1 U18108 ( .A1(\mem[804][4] ), .A2(n16531), .B1(n26326), .B2(
        data_in[4]), .ZN(n16535) );
  INV_X1 U18109 ( .A(n16536), .ZN(n19669) );
  AOI22_X1 U18110 ( .A1(\mem[804][5] ), .A2(n16531), .B1(n26326), .B2(
        data_in[5]), .ZN(n16536) );
  INV_X1 U18111 ( .A(n16537), .ZN(n19668) );
  AOI22_X1 U18112 ( .A1(\mem[804][6] ), .A2(n16531), .B1(n26326), .B2(
        data_in[6]), .ZN(n16537) );
  INV_X1 U18113 ( .A(n16538), .ZN(n19667) );
  AOI22_X1 U18114 ( .A1(\mem[804][7] ), .A2(n16531), .B1(n26326), .B2(
        data_in[7]), .ZN(n16538) );
  INV_X1 U18115 ( .A(n16539), .ZN(n19666) );
  AOI22_X1 U18116 ( .A1(\mem[805][0] ), .A2(n16540), .B1(n26325), .B2(
        data_in[0]), .ZN(n16539) );
  INV_X1 U18117 ( .A(n16541), .ZN(n19665) );
  AOI22_X1 U18118 ( .A1(\mem[805][1] ), .A2(n16540), .B1(n26325), .B2(
        data_in[1]), .ZN(n16541) );
  INV_X1 U18119 ( .A(n16542), .ZN(n19664) );
  AOI22_X1 U18120 ( .A1(\mem[805][2] ), .A2(n16540), .B1(n26325), .B2(
        data_in[2]), .ZN(n16542) );
  INV_X1 U18121 ( .A(n16543), .ZN(n19663) );
  AOI22_X1 U18122 ( .A1(\mem[805][3] ), .A2(n16540), .B1(n26325), .B2(
        data_in[3]), .ZN(n16543) );
  INV_X1 U18123 ( .A(n16544), .ZN(n19662) );
  AOI22_X1 U18124 ( .A1(\mem[805][4] ), .A2(n16540), .B1(n26325), .B2(
        data_in[4]), .ZN(n16544) );
  INV_X1 U18125 ( .A(n16545), .ZN(n19661) );
  AOI22_X1 U18126 ( .A1(\mem[805][5] ), .A2(n16540), .B1(n26325), .B2(
        data_in[5]), .ZN(n16545) );
  INV_X1 U18127 ( .A(n16546), .ZN(n19660) );
  AOI22_X1 U18128 ( .A1(\mem[805][6] ), .A2(n16540), .B1(n26325), .B2(
        data_in[6]), .ZN(n16546) );
  INV_X1 U18129 ( .A(n16547), .ZN(n19659) );
  AOI22_X1 U18130 ( .A1(\mem[805][7] ), .A2(n16540), .B1(n26325), .B2(
        data_in[7]), .ZN(n16547) );
  INV_X1 U18131 ( .A(n16548), .ZN(n19658) );
  AOI22_X1 U18132 ( .A1(\mem[806][0] ), .A2(n16549), .B1(n26324), .B2(
        data_in[0]), .ZN(n16548) );
  INV_X1 U18133 ( .A(n16550), .ZN(n19657) );
  AOI22_X1 U18134 ( .A1(\mem[806][1] ), .A2(n16549), .B1(n26324), .B2(
        data_in[1]), .ZN(n16550) );
  INV_X1 U18135 ( .A(n16551), .ZN(n19656) );
  AOI22_X1 U18136 ( .A1(\mem[806][2] ), .A2(n16549), .B1(n26324), .B2(
        data_in[2]), .ZN(n16551) );
  INV_X1 U18137 ( .A(n16552), .ZN(n19655) );
  AOI22_X1 U18138 ( .A1(\mem[806][3] ), .A2(n16549), .B1(n26324), .B2(
        data_in[3]), .ZN(n16552) );
  INV_X1 U18139 ( .A(n16553), .ZN(n19654) );
  AOI22_X1 U18140 ( .A1(\mem[806][4] ), .A2(n16549), .B1(n26324), .B2(
        data_in[4]), .ZN(n16553) );
  INV_X1 U18141 ( .A(n16554), .ZN(n19653) );
  AOI22_X1 U18142 ( .A1(\mem[806][5] ), .A2(n16549), .B1(n26324), .B2(
        data_in[5]), .ZN(n16554) );
  INV_X1 U18143 ( .A(n16555), .ZN(n19652) );
  AOI22_X1 U18144 ( .A1(\mem[806][6] ), .A2(n16549), .B1(n26324), .B2(
        data_in[6]), .ZN(n16555) );
  INV_X1 U18145 ( .A(n16556), .ZN(n19651) );
  AOI22_X1 U18146 ( .A1(\mem[806][7] ), .A2(n16549), .B1(n26324), .B2(
        data_in[7]), .ZN(n16556) );
  INV_X1 U18147 ( .A(n16557), .ZN(n19650) );
  AOI22_X1 U18148 ( .A1(\mem[807][0] ), .A2(n16558), .B1(n26323), .B2(
        data_in[0]), .ZN(n16557) );
  INV_X1 U18149 ( .A(n16559), .ZN(n19649) );
  AOI22_X1 U18150 ( .A1(\mem[807][1] ), .A2(n16558), .B1(n26323), .B2(
        data_in[1]), .ZN(n16559) );
  INV_X1 U18151 ( .A(n16560), .ZN(n19648) );
  AOI22_X1 U18152 ( .A1(\mem[807][2] ), .A2(n16558), .B1(n26323), .B2(
        data_in[2]), .ZN(n16560) );
  INV_X1 U18153 ( .A(n16561), .ZN(n19647) );
  AOI22_X1 U18154 ( .A1(\mem[807][3] ), .A2(n16558), .B1(n26323), .B2(
        data_in[3]), .ZN(n16561) );
  INV_X1 U18155 ( .A(n16562), .ZN(n19646) );
  AOI22_X1 U18156 ( .A1(\mem[807][4] ), .A2(n16558), .B1(n26323), .B2(
        data_in[4]), .ZN(n16562) );
  INV_X1 U18157 ( .A(n16563), .ZN(n19645) );
  AOI22_X1 U18158 ( .A1(\mem[807][5] ), .A2(n16558), .B1(n26323), .B2(
        data_in[5]), .ZN(n16563) );
  INV_X1 U18159 ( .A(n16564), .ZN(n19644) );
  AOI22_X1 U18160 ( .A1(\mem[807][6] ), .A2(n16558), .B1(n26323), .B2(
        data_in[6]), .ZN(n16564) );
  INV_X1 U18161 ( .A(n16565), .ZN(n19643) );
  AOI22_X1 U18162 ( .A1(\mem[807][7] ), .A2(n16558), .B1(n26323), .B2(
        data_in[7]), .ZN(n16565) );
  INV_X1 U18163 ( .A(n16782), .ZN(n19450) );
  AOI22_X1 U18164 ( .A1(\mem[832][0] ), .A2(n16783), .B1(n26298), .B2(
        data_in[0]), .ZN(n16782) );
  INV_X1 U18165 ( .A(n16784), .ZN(n19449) );
  AOI22_X1 U18166 ( .A1(\mem[832][1] ), .A2(n16783), .B1(n26298), .B2(
        data_in[1]), .ZN(n16784) );
  INV_X1 U18167 ( .A(n16785), .ZN(n19448) );
  AOI22_X1 U18168 ( .A1(\mem[832][2] ), .A2(n16783), .B1(n26298), .B2(
        data_in[2]), .ZN(n16785) );
  INV_X1 U18169 ( .A(n16786), .ZN(n19447) );
  AOI22_X1 U18170 ( .A1(\mem[832][3] ), .A2(n16783), .B1(n26298), .B2(
        data_in[3]), .ZN(n16786) );
  INV_X1 U18171 ( .A(n16787), .ZN(n19446) );
  AOI22_X1 U18172 ( .A1(\mem[832][4] ), .A2(n16783), .B1(n26298), .B2(
        data_in[4]), .ZN(n16787) );
  INV_X1 U18173 ( .A(n16788), .ZN(n19445) );
  AOI22_X1 U18174 ( .A1(\mem[832][5] ), .A2(n16783), .B1(n26298), .B2(
        data_in[5]), .ZN(n16788) );
  INV_X1 U18175 ( .A(n16789), .ZN(n19444) );
  AOI22_X1 U18176 ( .A1(\mem[832][6] ), .A2(n16783), .B1(n26298), .B2(
        data_in[6]), .ZN(n16789) );
  INV_X1 U18177 ( .A(n16790), .ZN(n19443) );
  AOI22_X1 U18178 ( .A1(\mem[832][7] ), .A2(n16783), .B1(n26298), .B2(
        data_in[7]), .ZN(n16790) );
  INV_X1 U18179 ( .A(n16792), .ZN(n19442) );
  AOI22_X1 U18180 ( .A1(\mem[833][0] ), .A2(n16793), .B1(n26297), .B2(
        data_in[0]), .ZN(n16792) );
  INV_X1 U18181 ( .A(n16794), .ZN(n19441) );
  AOI22_X1 U18182 ( .A1(\mem[833][1] ), .A2(n16793), .B1(n26297), .B2(
        data_in[1]), .ZN(n16794) );
  INV_X1 U18183 ( .A(n16795), .ZN(n19440) );
  AOI22_X1 U18184 ( .A1(\mem[833][2] ), .A2(n16793), .B1(n26297), .B2(
        data_in[2]), .ZN(n16795) );
  INV_X1 U18185 ( .A(n16796), .ZN(n19439) );
  AOI22_X1 U18186 ( .A1(\mem[833][3] ), .A2(n16793), .B1(n26297), .B2(
        data_in[3]), .ZN(n16796) );
  INV_X1 U18187 ( .A(n16797), .ZN(n19438) );
  AOI22_X1 U18188 ( .A1(\mem[833][4] ), .A2(n16793), .B1(n26297), .B2(
        data_in[4]), .ZN(n16797) );
  INV_X1 U18189 ( .A(n16798), .ZN(n19437) );
  AOI22_X1 U18190 ( .A1(\mem[833][5] ), .A2(n16793), .B1(n26297), .B2(
        data_in[5]), .ZN(n16798) );
  INV_X1 U18191 ( .A(n16799), .ZN(n19436) );
  AOI22_X1 U18192 ( .A1(\mem[833][6] ), .A2(n16793), .B1(n26297), .B2(
        data_in[6]), .ZN(n16799) );
  INV_X1 U18193 ( .A(n16800), .ZN(n19435) );
  AOI22_X1 U18194 ( .A1(\mem[833][7] ), .A2(n16793), .B1(n26297), .B2(
        data_in[7]), .ZN(n16800) );
  INV_X1 U18195 ( .A(n16801), .ZN(n19434) );
  AOI22_X1 U18196 ( .A1(\mem[834][0] ), .A2(n16802), .B1(n26296), .B2(
        data_in[0]), .ZN(n16801) );
  INV_X1 U18197 ( .A(n16803), .ZN(n19433) );
  AOI22_X1 U18198 ( .A1(\mem[834][1] ), .A2(n16802), .B1(n26296), .B2(
        data_in[1]), .ZN(n16803) );
  INV_X1 U18199 ( .A(n16804), .ZN(n19432) );
  AOI22_X1 U18200 ( .A1(\mem[834][2] ), .A2(n16802), .B1(n26296), .B2(
        data_in[2]), .ZN(n16804) );
  INV_X1 U18201 ( .A(n16805), .ZN(n19431) );
  AOI22_X1 U18202 ( .A1(\mem[834][3] ), .A2(n16802), .B1(n26296), .B2(
        data_in[3]), .ZN(n16805) );
  INV_X1 U18203 ( .A(n16806), .ZN(n19430) );
  AOI22_X1 U18204 ( .A1(\mem[834][4] ), .A2(n16802), .B1(n26296), .B2(
        data_in[4]), .ZN(n16806) );
  INV_X1 U18205 ( .A(n16807), .ZN(n19429) );
  AOI22_X1 U18206 ( .A1(\mem[834][5] ), .A2(n16802), .B1(n26296), .B2(
        data_in[5]), .ZN(n16807) );
  INV_X1 U18207 ( .A(n16808), .ZN(n19428) );
  AOI22_X1 U18208 ( .A1(\mem[834][6] ), .A2(n16802), .B1(n26296), .B2(
        data_in[6]), .ZN(n16808) );
  INV_X1 U18209 ( .A(n16809), .ZN(n19427) );
  AOI22_X1 U18210 ( .A1(\mem[834][7] ), .A2(n16802), .B1(n26296), .B2(
        data_in[7]), .ZN(n16809) );
  INV_X1 U18211 ( .A(n16810), .ZN(n19426) );
  AOI22_X1 U18212 ( .A1(\mem[835][0] ), .A2(n16811), .B1(n26295), .B2(
        data_in[0]), .ZN(n16810) );
  INV_X1 U18213 ( .A(n16812), .ZN(n19425) );
  AOI22_X1 U18214 ( .A1(\mem[835][1] ), .A2(n16811), .B1(n26295), .B2(
        data_in[1]), .ZN(n16812) );
  INV_X1 U18215 ( .A(n16813), .ZN(n19424) );
  AOI22_X1 U18216 ( .A1(\mem[835][2] ), .A2(n16811), .B1(n26295), .B2(
        data_in[2]), .ZN(n16813) );
  INV_X1 U18217 ( .A(n16814), .ZN(n19423) );
  AOI22_X1 U18218 ( .A1(\mem[835][3] ), .A2(n16811), .B1(n26295), .B2(
        data_in[3]), .ZN(n16814) );
  INV_X1 U18219 ( .A(n16815), .ZN(n19422) );
  AOI22_X1 U18220 ( .A1(\mem[835][4] ), .A2(n16811), .B1(n26295), .B2(
        data_in[4]), .ZN(n16815) );
  INV_X1 U18221 ( .A(n16816), .ZN(n19421) );
  AOI22_X1 U18222 ( .A1(\mem[835][5] ), .A2(n16811), .B1(n26295), .B2(
        data_in[5]), .ZN(n16816) );
  INV_X1 U18223 ( .A(n16817), .ZN(n19420) );
  AOI22_X1 U18224 ( .A1(\mem[835][6] ), .A2(n16811), .B1(n26295), .B2(
        data_in[6]), .ZN(n16817) );
  INV_X1 U18225 ( .A(n16818), .ZN(n19419) );
  AOI22_X1 U18226 ( .A1(\mem[835][7] ), .A2(n16811), .B1(n26295), .B2(
        data_in[7]), .ZN(n16818) );
  INV_X1 U18227 ( .A(n16819), .ZN(n19418) );
  AOI22_X1 U18228 ( .A1(\mem[836][0] ), .A2(n16820), .B1(n26294), .B2(
        data_in[0]), .ZN(n16819) );
  INV_X1 U18229 ( .A(n16821), .ZN(n19417) );
  AOI22_X1 U18230 ( .A1(\mem[836][1] ), .A2(n16820), .B1(n26294), .B2(
        data_in[1]), .ZN(n16821) );
  INV_X1 U18231 ( .A(n16822), .ZN(n19416) );
  AOI22_X1 U18232 ( .A1(\mem[836][2] ), .A2(n16820), .B1(n26294), .B2(
        data_in[2]), .ZN(n16822) );
  INV_X1 U18233 ( .A(n16823), .ZN(n19415) );
  AOI22_X1 U18234 ( .A1(\mem[836][3] ), .A2(n16820), .B1(n26294), .B2(
        data_in[3]), .ZN(n16823) );
  INV_X1 U18235 ( .A(n16824), .ZN(n19414) );
  AOI22_X1 U18236 ( .A1(\mem[836][4] ), .A2(n16820), .B1(n26294), .B2(
        data_in[4]), .ZN(n16824) );
  INV_X1 U18237 ( .A(n16825), .ZN(n19413) );
  AOI22_X1 U18238 ( .A1(\mem[836][5] ), .A2(n16820), .B1(n26294), .B2(
        data_in[5]), .ZN(n16825) );
  INV_X1 U18239 ( .A(n16826), .ZN(n19412) );
  AOI22_X1 U18240 ( .A1(\mem[836][6] ), .A2(n16820), .B1(n26294), .B2(
        data_in[6]), .ZN(n16826) );
  INV_X1 U18241 ( .A(n16827), .ZN(n19411) );
  AOI22_X1 U18242 ( .A1(\mem[836][7] ), .A2(n16820), .B1(n26294), .B2(
        data_in[7]), .ZN(n16827) );
  INV_X1 U18243 ( .A(n16828), .ZN(n19410) );
  AOI22_X1 U18244 ( .A1(\mem[837][0] ), .A2(n16829), .B1(n26293), .B2(
        data_in[0]), .ZN(n16828) );
  INV_X1 U18245 ( .A(n16830), .ZN(n19409) );
  AOI22_X1 U18246 ( .A1(\mem[837][1] ), .A2(n16829), .B1(n26293), .B2(
        data_in[1]), .ZN(n16830) );
  INV_X1 U18247 ( .A(n16831), .ZN(n19408) );
  AOI22_X1 U18248 ( .A1(\mem[837][2] ), .A2(n16829), .B1(n26293), .B2(
        data_in[2]), .ZN(n16831) );
  INV_X1 U18249 ( .A(n16832), .ZN(n19407) );
  AOI22_X1 U18250 ( .A1(\mem[837][3] ), .A2(n16829), .B1(n26293), .B2(
        data_in[3]), .ZN(n16832) );
  INV_X1 U18251 ( .A(n16833), .ZN(n19406) );
  AOI22_X1 U18252 ( .A1(\mem[837][4] ), .A2(n16829), .B1(n26293), .B2(
        data_in[4]), .ZN(n16833) );
  INV_X1 U18253 ( .A(n16834), .ZN(n19405) );
  AOI22_X1 U18254 ( .A1(\mem[837][5] ), .A2(n16829), .B1(n26293), .B2(
        data_in[5]), .ZN(n16834) );
  INV_X1 U18255 ( .A(n16835), .ZN(n19404) );
  AOI22_X1 U18256 ( .A1(\mem[837][6] ), .A2(n16829), .B1(n26293), .B2(
        data_in[6]), .ZN(n16835) );
  INV_X1 U18257 ( .A(n16836), .ZN(n19403) );
  AOI22_X1 U18258 ( .A1(\mem[837][7] ), .A2(n16829), .B1(n26293), .B2(
        data_in[7]), .ZN(n16836) );
  INV_X1 U18259 ( .A(n16837), .ZN(n19402) );
  AOI22_X1 U18260 ( .A1(\mem[838][0] ), .A2(n16838), .B1(n26292), .B2(
        data_in[0]), .ZN(n16837) );
  INV_X1 U18261 ( .A(n16839), .ZN(n19401) );
  AOI22_X1 U18262 ( .A1(\mem[838][1] ), .A2(n16838), .B1(n26292), .B2(
        data_in[1]), .ZN(n16839) );
  INV_X1 U18263 ( .A(n16840), .ZN(n19400) );
  AOI22_X1 U18264 ( .A1(\mem[838][2] ), .A2(n16838), .B1(n26292), .B2(
        data_in[2]), .ZN(n16840) );
  INV_X1 U18265 ( .A(n16841), .ZN(n19399) );
  AOI22_X1 U18266 ( .A1(\mem[838][3] ), .A2(n16838), .B1(n26292), .B2(
        data_in[3]), .ZN(n16841) );
  INV_X1 U18267 ( .A(n16842), .ZN(n19398) );
  AOI22_X1 U18268 ( .A1(\mem[838][4] ), .A2(n16838), .B1(n26292), .B2(
        data_in[4]), .ZN(n16842) );
  INV_X1 U18269 ( .A(n16843), .ZN(n19397) );
  AOI22_X1 U18270 ( .A1(\mem[838][5] ), .A2(n16838), .B1(n26292), .B2(
        data_in[5]), .ZN(n16843) );
  INV_X1 U18271 ( .A(n16844), .ZN(n19396) );
  AOI22_X1 U18272 ( .A1(\mem[838][6] ), .A2(n16838), .B1(n26292), .B2(
        data_in[6]), .ZN(n16844) );
  INV_X1 U18273 ( .A(n16845), .ZN(n19395) );
  AOI22_X1 U18274 ( .A1(\mem[838][7] ), .A2(n16838), .B1(n26292), .B2(
        data_in[7]), .ZN(n16845) );
  INV_X1 U18275 ( .A(n16846), .ZN(n19394) );
  AOI22_X1 U18276 ( .A1(\mem[839][0] ), .A2(n16847), .B1(n26291), .B2(
        data_in[0]), .ZN(n16846) );
  INV_X1 U18277 ( .A(n16848), .ZN(n19393) );
  AOI22_X1 U18278 ( .A1(\mem[839][1] ), .A2(n16847), .B1(n26291), .B2(
        data_in[1]), .ZN(n16848) );
  INV_X1 U18279 ( .A(n16849), .ZN(n19392) );
  AOI22_X1 U18280 ( .A1(\mem[839][2] ), .A2(n16847), .B1(n26291), .B2(
        data_in[2]), .ZN(n16849) );
  INV_X1 U18281 ( .A(n16850), .ZN(n19391) );
  AOI22_X1 U18282 ( .A1(\mem[839][3] ), .A2(n16847), .B1(n26291), .B2(
        data_in[3]), .ZN(n16850) );
  INV_X1 U18283 ( .A(n16851), .ZN(n19390) );
  AOI22_X1 U18284 ( .A1(\mem[839][4] ), .A2(n16847), .B1(n26291), .B2(
        data_in[4]), .ZN(n16851) );
  INV_X1 U18285 ( .A(n16852), .ZN(n19389) );
  AOI22_X1 U18286 ( .A1(\mem[839][5] ), .A2(n16847), .B1(n26291), .B2(
        data_in[5]), .ZN(n16852) );
  INV_X1 U18287 ( .A(n16853), .ZN(n19388) );
  AOI22_X1 U18288 ( .A1(\mem[839][6] ), .A2(n16847), .B1(n26291), .B2(
        data_in[6]), .ZN(n16853) );
  INV_X1 U18289 ( .A(n16854), .ZN(n19387) );
  AOI22_X1 U18290 ( .A1(\mem[839][7] ), .A2(n16847), .B1(n26291), .B2(
        data_in[7]), .ZN(n16854) );
  INV_X1 U18291 ( .A(n17071), .ZN(n19194) );
  AOI22_X1 U18292 ( .A1(\mem[864][0] ), .A2(n17072), .B1(n26266), .B2(
        data_in[0]), .ZN(n17071) );
  INV_X1 U18293 ( .A(n17073), .ZN(n19193) );
  AOI22_X1 U18294 ( .A1(\mem[864][1] ), .A2(n17072), .B1(n26266), .B2(
        data_in[1]), .ZN(n17073) );
  INV_X1 U18295 ( .A(n17074), .ZN(n19192) );
  AOI22_X1 U18296 ( .A1(\mem[864][2] ), .A2(n17072), .B1(n26266), .B2(
        data_in[2]), .ZN(n17074) );
  INV_X1 U18297 ( .A(n17075), .ZN(n19191) );
  AOI22_X1 U18298 ( .A1(\mem[864][3] ), .A2(n17072), .B1(n26266), .B2(
        data_in[3]), .ZN(n17075) );
  INV_X1 U18299 ( .A(n17076), .ZN(n19190) );
  AOI22_X1 U18300 ( .A1(\mem[864][4] ), .A2(n17072), .B1(n26266), .B2(
        data_in[4]), .ZN(n17076) );
  INV_X1 U18301 ( .A(n17077), .ZN(n19189) );
  AOI22_X1 U18302 ( .A1(\mem[864][5] ), .A2(n17072), .B1(n26266), .B2(
        data_in[5]), .ZN(n17077) );
  INV_X1 U18303 ( .A(n17078), .ZN(n19188) );
  AOI22_X1 U18304 ( .A1(\mem[864][6] ), .A2(n17072), .B1(n26266), .B2(
        data_in[6]), .ZN(n17078) );
  INV_X1 U18305 ( .A(n17079), .ZN(n19187) );
  AOI22_X1 U18306 ( .A1(\mem[864][7] ), .A2(n17072), .B1(n26266), .B2(
        data_in[7]), .ZN(n17079) );
  INV_X1 U18307 ( .A(n17081), .ZN(n19186) );
  AOI22_X1 U18308 ( .A1(\mem[865][0] ), .A2(n17082), .B1(n26265), .B2(
        data_in[0]), .ZN(n17081) );
  INV_X1 U18309 ( .A(n17083), .ZN(n19185) );
  AOI22_X1 U18310 ( .A1(\mem[865][1] ), .A2(n17082), .B1(n26265), .B2(
        data_in[1]), .ZN(n17083) );
  INV_X1 U18311 ( .A(n17084), .ZN(n19184) );
  AOI22_X1 U18312 ( .A1(\mem[865][2] ), .A2(n17082), .B1(n26265), .B2(
        data_in[2]), .ZN(n17084) );
  INV_X1 U18313 ( .A(n17085), .ZN(n19183) );
  AOI22_X1 U18314 ( .A1(\mem[865][3] ), .A2(n17082), .B1(n26265), .B2(
        data_in[3]), .ZN(n17085) );
  INV_X1 U18315 ( .A(n17086), .ZN(n19182) );
  AOI22_X1 U18316 ( .A1(\mem[865][4] ), .A2(n17082), .B1(n26265), .B2(
        data_in[4]), .ZN(n17086) );
  INV_X1 U18317 ( .A(n17087), .ZN(n19181) );
  AOI22_X1 U18318 ( .A1(\mem[865][5] ), .A2(n17082), .B1(n26265), .B2(
        data_in[5]), .ZN(n17087) );
  INV_X1 U18319 ( .A(n17088), .ZN(n19180) );
  AOI22_X1 U18320 ( .A1(\mem[865][6] ), .A2(n17082), .B1(n26265), .B2(
        data_in[6]), .ZN(n17088) );
  INV_X1 U18321 ( .A(n17089), .ZN(n19179) );
  AOI22_X1 U18322 ( .A1(\mem[865][7] ), .A2(n17082), .B1(n26265), .B2(
        data_in[7]), .ZN(n17089) );
  INV_X1 U18323 ( .A(n17090), .ZN(n19178) );
  AOI22_X1 U18324 ( .A1(\mem[866][0] ), .A2(n17091), .B1(n26264), .B2(
        data_in[0]), .ZN(n17090) );
  INV_X1 U18325 ( .A(n17092), .ZN(n19177) );
  AOI22_X1 U18326 ( .A1(\mem[866][1] ), .A2(n17091), .B1(n26264), .B2(
        data_in[1]), .ZN(n17092) );
  INV_X1 U18327 ( .A(n17093), .ZN(n19176) );
  AOI22_X1 U18328 ( .A1(\mem[866][2] ), .A2(n17091), .B1(n26264), .B2(
        data_in[2]), .ZN(n17093) );
  INV_X1 U18329 ( .A(n17094), .ZN(n19175) );
  AOI22_X1 U18330 ( .A1(\mem[866][3] ), .A2(n17091), .B1(n26264), .B2(
        data_in[3]), .ZN(n17094) );
  INV_X1 U18331 ( .A(n17095), .ZN(n19174) );
  AOI22_X1 U18332 ( .A1(\mem[866][4] ), .A2(n17091), .B1(n26264), .B2(
        data_in[4]), .ZN(n17095) );
  INV_X1 U18333 ( .A(n17096), .ZN(n19173) );
  AOI22_X1 U18334 ( .A1(\mem[866][5] ), .A2(n17091), .B1(n26264), .B2(
        data_in[5]), .ZN(n17096) );
  INV_X1 U18335 ( .A(n17097), .ZN(n19172) );
  AOI22_X1 U18336 ( .A1(\mem[866][6] ), .A2(n17091), .B1(n26264), .B2(
        data_in[6]), .ZN(n17097) );
  INV_X1 U18337 ( .A(n17098), .ZN(n19171) );
  AOI22_X1 U18338 ( .A1(\mem[866][7] ), .A2(n17091), .B1(n26264), .B2(
        data_in[7]), .ZN(n17098) );
  INV_X1 U18339 ( .A(n17099), .ZN(n19170) );
  AOI22_X1 U18340 ( .A1(\mem[867][0] ), .A2(n17100), .B1(n26263), .B2(
        data_in[0]), .ZN(n17099) );
  INV_X1 U18341 ( .A(n17101), .ZN(n19169) );
  AOI22_X1 U18342 ( .A1(\mem[867][1] ), .A2(n17100), .B1(n26263), .B2(
        data_in[1]), .ZN(n17101) );
  INV_X1 U18343 ( .A(n17102), .ZN(n19168) );
  AOI22_X1 U18344 ( .A1(\mem[867][2] ), .A2(n17100), .B1(n26263), .B2(
        data_in[2]), .ZN(n17102) );
  INV_X1 U18345 ( .A(n17103), .ZN(n19167) );
  AOI22_X1 U18346 ( .A1(\mem[867][3] ), .A2(n17100), .B1(n26263), .B2(
        data_in[3]), .ZN(n17103) );
  INV_X1 U18347 ( .A(n17104), .ZN(n19166) );
  AOI22_X1 U18348 ( .A1(\mem[867][4] ), .A2(n17100), .B1(n26263), .B2(
        data_in[4]), .ZN(n17104) );
  INV_X1 U18349 ( .A(n17105), .ZN(n19165) );
  AOI22_X1 U18350 ( .A1(\mem[867][5] ), .A2(n17100), .B1(n26263), .B2(
        data_in[5]), .ZN(n17105) );
  INV_X1 U18351 ( .A(n17106), .ZN(n19164) );
  AOI22_X1 U18352 ( .A1(\mem[867][6] ), .A2(n17100), .B1(n26263), .B2(
        data_in[6]), .ZN(n17106) );
  INV_X1 U18353 ( .A(n17107), .ZN(n19163) );
  AOI22_X1 U18354 ( .A1(\mem[867][7] ), .A2(n17100), .B1(n26263), .B2(
        data_in[7]), .ZN(n17107) );
  INV_X1 U18355 ( .A(n17108), .ZN(n19162) );
  AOI22_X1 U18356 ( .A1(\mem[868][0] ), .A2(n17109), .B1(n26262), .B2(
        data_in[0]), .ZN(n17108) );
  INV_X1 U18357 ( .A(n17110), .ZN(n19161) );
  AOI22_X1 U18358 ( .A1(\mem[868][1] ), .A2(n17109), .B1(n26262), .B2(
        data_in[1]), .ZN(n17110) );
  INV_X1 U18359 ( .A(n17111), .ZN(n19160) );
  AOI22_X1 U18360 ( .A1(\mem[868][2] ), .A2(n17109), .B1(n26262), .B2(
        data_in[2]), .ZN(n17111) );
  INV_X1 U18361 ( .A(n17112), .ZN(n19159) );
  AOI22_X1 U18362 ( .A1(\mem[868][3] ), .A2(n17109), .B1(n26262), .B2(
        data_in[3]), .ZN(n17112) );
  INV_X1 U18363 ( .A(n17113), .ZN(n19158) );
  AOI22_X1 U18364 ( .A1(\mem[868][4] ), .A2(n17109), .B1(n26262), .B2(
        data_in[4]), .ZN(n17113) );
  INV_X1 U18365 ( .A(n17114), .ZN(n19157) );
  AOI22_X1 U18366 ( .A1(\mem[868][5] ), .A2(n17109), .B1(n26262), .B2(
        data_in[5]), .ZN(n17114) );
  INV_X1 U18367 ( .A(n17115), .ZN(n19156) );
  AOI22_X1 U18368 ( .A1(\mem[868][6] ), .A2(n17109), .B1(n26262), .B2(
        data_in[6]), .ZN(n17115) );
  INV_X1 U18369 ( .A(n17116), .ZN(n19155) );
  AOI22_X1 U18370 ( .A1(\mem[868][7] ), .A2(n17109), .B1(n26262), .B2(
        data_in[7]), .ZN(n17116) );
  INV_X1 U18371 ( .A(n17117), .ZN(n19154) );
  AOI22_X1 U18372 ( .A1(\mem[869][0] ), .A2(n17118), .B1(n26261), .B2(
        data_in[0]), .ZN(n17117) );
  INV_X1 U18373 ( .A(n17119), .ZN(n19153) );
  AOI22_X1 U18374 ( .A1(\mem[869][1] ), .A2(n17118), .B1(n26261), .B2(
        data_in[1]), .ZN(n17119) );
  INV_X1 U18375 ( .A(n17120), .ZN(n19152) );
  AOI22_X1 U18376 ( .A1(\mem[869][2] ), .A2(n17118), .B1(n26261), .B2(
        data_in[2]), .ZN(n17120) );
  INV_X1 U18377 ( .A(n17121), .ZN(n19151) );
  AOI22_X1 U18378 ( .A1(\mem[869][3] ), .A2(n17118), .B1(n26261), .B2(
        data_in[3]), .ZN(n17121) );
  INV_X1 U18379 ( .A(n17122), .ZN(n19150) );
  AOI22_X1 U18380 ( .A1(\mem[869][4] ), .A2(n17118), .B1(n26261), .B2(
        data_in[4]), .ZN(n17122) );
  INV_X1 U18381 ( .A(n17123), .ZN(n19149) );
  AOI22_X1 U18382 ( .A1(\mem[869][5] ), .A2(n17118), .B1(n26261), .B2(
        data_in[5]), .ZN(n17123) );
  INV_X1 U18383 ( .A(n17124), .ZN(n19148) );
  AOI22_X1 U18384 ( .A1(\mem[869][6] ), .A2(n17118), .B1(n26261), .B2(
        data_in[6]), .ZN(n17124) );
  INV_X1 U18385 ( .A(n17125), .ZN(n19147) );
  AOI22_X1 U18386 ( .A1(\mem[869][7] ), .A2(n17118), .B1(n26261), .B2(
        data_in[7]), .ZN(n17125) );
  INV_X1 U18387 ( .A(n17126), .ZN(n19146) );
  AOI22_X1 U18388 ( .A1(\mem[870][0] ), .A2(n17127), .B1(n26260), .B2(
        data_in[0]), .ZN(n17126) );
  INV_X1 U18389 ( .A(n17128), .ZN(n19145) );
  AOI22_X1 U18390 ( .A1(\mem[870][1] ), .A2(n17127), .B1(n26260), .B2(
        data_in[1]), .ZN(n17128) );
  INV_X1 U18391 ( .A(n17129), .ZN(n19144) );
  AOI22_X1 U18392 ( .A1(\mem[870][2] ), .A2(n17127), .B1(n26260), .B2(
        data_in[2]), .ZN(n17129) );
  INV_X1 U18393 ( .A(n17130), .ZN(n19143) );
  AOI22_X1 U18394 ( .A1(\mem[870][3] ), .A2(n17127), .B1(n26260), .B2(
        data_in[3]), .ZN(n17130) );
  INV_X1 U18395 ( .A(n17131), .ZN(n19142) );
  AOI22_X1 U18396 ( .A1(\mem[870][4] ), .A2(n17127), .B1(n26260), .B2(
        data_in[4]), .ZN(n17131) );
  INV_X1 U18397 ( .A(n17132), .ZN(n19141) );
  AOI22_X1 U18398 ( .A1(\mem[870][5] ), .A2(n17127), .B1(n26260), .B2(
        data_in[5]), .ZN(n17132) );
  INV_X1 U18399 ( .A(n17133), .ZN(n19140) );
  AOI22_X1 U18400 ( .A1(\mem[870][6] ), .A2(n17127), .B1(n26260), .B2(
        data_in[6]), .ZN(n17133) );
  INV_X1 U18401 ( .A(n17134), .ZN(n19139) );
  AOI22_X1 U18402 ( .A1(\mem[870][7] ), .A2(n17127), .B1(n26260), .B2(
        data_in[7]), .ZN(n17134) );
  INV_X1 U18403 ( .A(n17135), .ZN(n19138) );
  AOI22_X1 U18404 ( .A1(\mem[871][0] ), .A2(n17136), .B1(n26259), .B2(
        data_in[0]), .ZN(n17135) );
  INV_X1 U18405 ( .A(n17137), .ZN(n19137) );
  AOI22_X1 U18406 ( .A1(\mem[871][1] ), .A2(n17136), .B1(n26259), .B2(
        data_in[1]), .ZN(n17137) );
  INV_X1 U18407 ( .A(n17138), .ZN(n19136) );
  AOI22_X1 U18408 ( .A1(\mem[871][2] ), .A2(n17136), .B1(n26259), .B2(
        data_in[2]), .ZN(n17138) );
  INV_X1 U18409 ( .A(n17139), .ZN(n19135) );
  AOI22_X1 U18410 ( .A1(\mem[871][3] ), .A2(n17136), .B1(n26259), .B2(
        data_in[3]), .ZN(n17139) );
  INV_X1 U18411 ( .A(n17140), .ZN(n19134) );
  AOI22_X1 U18412 ( .A1(\mem[871][4] ), .A2(n17136), .B1(n26259), .B2(
        data_in[4]), .ZN(n17140) );
  INV_X1 U18413 ( .A(n17141), .ZN(n19133) );
  AOI22_X1 U18414 ( .A1(\mem[871][5] ), .A2(n17136), .B1(n26259), .B2(
        data_in[5]), .ZN(n17141) );
  INV_X1 U18415 ( .A(n17142), .ZN(n19132) );
  AOI22_X1 U18416 ( .A1(\mem[871][6] ), .A2(n17136), .B1(n26259), .B2(
        data_in[6]), .ZN(n17142) );
  INV_X1 U18417 ( .A(n17143), .ZN(n19131) );
  AOI22_X1 U18418 ( .A1(\mem[871][7] ), .A2(n17136), .B1(n26259), .B2(
        data_in[7]), .ZN(n17143) );
  INV_X1 U18419 ( .A(n17360), .ZN(n18938) );
  AOI22_X1 U18420 ( .A1(\mem[896][0] ), .A2(n17361), .B1(n26234), .B2(
        data_in[0]), .ZN(n17360) );
  INV_X1 U18421 ( .A(n17362), .ZN(n18937) );
  AOI22_X1 U18422 ( .A1(\mem[896][1] ), .A2(n17361), .B1(n26234), .B2(
        data_in[1]), .ZN(n17362) );
  INV_X1 U18423 ( .A(n17363), .ZN(n18936) );
  AOI22_X1 U18424 ( .A1(\mem[896][2] ), .A2(n17361), .B1(n26234), .B2(
        data_in[2]), .ZN(n17363) );
  INV_X1 U18425 ( .A(n17364), .ZN(n18935) );
  AOI22_X1 U18426 ( .A1(\mem[896][3] ), .A2(n17361), .B1(n26234), .B2(
        data_in[3]), .ZN(n17364) );
  INV_X1 U18427 ( .A(n17365), .ZN(n18934) );
  AOI22_X1 U18428 ( .A1(\mem[896][4] ), .A2(n17361), .B1(n26234), .B2(
        data_in[4]), .ZN(n17365) );
  INV_X1 U18429 ( .A(n17366), .ZN(n18933) );
  AOI22_X1 U18430 ( .A1(\mem[896][5] ), .A2(n17361), .B1(n26234), .B2(
        data_in[5]), .ZN(n17366) );
  INV_X1 U18431 ( .A(n17367), .ZN(n18932) );
  AOI22_X1 U18432 ( .A1(\mem[896][6] ), .A2(n17361), .B1(n26234), .B2(
        data_in[6]), .ZN(n17367) );
  INV_X1 U18433 ( .A(n17368), .ZN(n18931) );
  AOI22_X1 U18434 ( .A1(\mem[896][7] ), .A2(n17361), .B1(n26234), .B2(
        data_in[7]), .ZN(n17368) );
  INV_X1 U18435 ( .A(n17370), .ZN(n18930) );
  AOI22_X1 U18436 ( .A1(\mem[897][0] ), .A2(n17371), .B1(n26233), .B2(
        data_in[0]), .ZN(n17370) );
  INV_X1 U18437 ( .A(n17372), .ZN(n18929) );
  AOI22_X1 U18438 ( .A1(\mem[897][1] ), .A2(n17371), .B1(n26233), .B2(
        data_in[1]), .ZN(n17372) );
  INV_X1 U18439 ( .A(n17373), .ZN(n18928) );
  AOI22_X1 U18440 ( .A1(\mem[897][2] ), .A2(n17371), .B1(n26233), .B2(
        data_in[2]), .ZN(n17373) );
  INV_X1 U18441 ( .A(n17374), .ZN(n18927) );
  AOI22_X1 U18442 ( .A1(\mem[897][3] ), .A2(n17371), .B1(n26233), .B2(
        data_in[3]), .ZN(n17374) );
  INV_X1 U18443 ( .A(n17375), .ZN(n18926) );
  AOI22_X1 U18444 ( .A1(\mem[897][4] ), .A2(n17371), .B1(n26233), .B2(
        data_in[4]), .ZN(n17375) );
  INV_X1 U18445 ( .A(n17376), .ZN(n18925) );
  AOI22_X1 U18446 ( .A1(\mem[897][5] ), .A2(n17371), .B1(n26233), .B2(
        data_in[5]), .ZN(n17376) );
  INV_X1 U18447 ( .A(n17377), .ZN(n18924) );
  AOI22_X1 U18448 ( .A1(\mem[897][6] ), .A2(n17371), .B1(n26233), .B2(
        data_in[6]), .ZN(n17377) );
  INV_X1 U18449 ( .A(n17378), .ZN(n18923) );
  AOI22_X1 U18450 ( .A1(\mem[897][7] ), .A2(n17371), .B1(n26233), .B2(
        data_in[7]), .ZN(n17378) );
  INV_X1 U18451 ( .A(n17379), .ZN(n18922) );
  AOI22_X1 U18452 ( .A1(\mem[898][0] ), .A2(n17380), .B1(n26232), .B2(
        data_in[0]), .ZN(n17379) );
  INV_X1 U18453 ( .A(n17381), .ZN(n18921) );
  AOI22_X1 U18454 ( .A1(\mem[898][1] ), .A2(n17380), .B1(n26232), .B2(
        data_in[1]), .ZN(n17381) );
  INV_X1 U18455 ( .A(n17382), .ZN(n18920) );
  AOI22_X1 U18456 ( .A1(\mem[898][2] ), .A2(n17380), .B1(n26232), .B2(
        data_in[2]), .ZN(n17382) );
  INV_X1 U18457 ( .A(n17383), .ZN(n18919) );
  AOI22_X1 U18458 ( .A1(\mem[898][3] ), .A2(n17380), .B1(n26232), .B2(
        data_in[3]), .ZN(n17383) );
  INV_X1 U18459 ( .A(n17384), .ZN(n18918) );
  AOI22_X1 U18460 ( .A1(\mem[898][4] ), .A2(n17380), .B1(n26232), .B2(
        data_in[4]), .ZN(n17384) );
  INV_X1 U18461 ( .A(n17385), .ZN(n18917) );
  AOI22_X1 U18462 ( .A1(\mem[898][5] ), .A2(n17380), .B1(n26232), .B2(
        data_in[5]), .ZN(n17385) );
  INV_X1 U18463 ( .A(n17386), .ZN(n18916) );
  AOI22_X1 U18464 ( .A1(\mem[898][6] ), .A2(n17380), .B1(n26232), .B2(
        data_in[6]), .ZN(n17386) );
  INV_X1 U18465 ( .A(n17387), .ZN(n18915) );
  AOI22_X1 U18466 ( .A1(\mem[898][7] ), .A2(n17380), .B1(n26232), .B2(
        data_in[7]), .ZN(n17387) );
  INV_X1 U18467 ( .A(n17388), .ZN(n18914) );
  AOI22_X1 U18468 ( .A1(\mem[899][0] ), .A2(n17389), .B1(n26231), .B2(
        data_in[0]), .ZN(n17388) );
  INV_X1 U18469 ( .A(n17390), .ZN(n18913) );
  AOI22_X1 U18470 ( .A1(\mem[899][1] ), .A2(n17389), .B1(n26231), .B2(
        data_in[1]), .ZN(n17390) );
  INV_X1 U18471 ( .A(n17391), .ZN(n18912) );
  AOI22_X1 U18472 ( .A1(\mem[899][2] ), .A2(n17389), .B1(n26231), .B2(
        data_in[2]), .ZN(n17391) );
  INV_X1 U18473 ( .A(n17392), .ZN(n18911) );
  AOI22_X1 U18474 ( .A1(\mem[899][3] ), .A2(n17389), .B1(n26231), .B2(
        data_in[3]), .ZN(n17392) );
  INV_X1 U18475 ( .A(n17393), .ZN(n18910) );
  AOI22_X1 U18476 ( .A1(\mem[899][4] ), .A2(n17389), .B1(n26231), .B2(
        data_in[4]), .ZN(n17393) );
  INV_X1 U18477 ( .A(n17394), .ZN(n18909) );
  AOI22_X1 U18478 ( .A1(\mem[899][5] ), .A2(n17389), .B1(n26231), .B2(
        data_in[5]), .ZN(n17394) );
  INV_X1 U18479 ( .A(n17395), .ZN(n18908) );
  AOI22_X1 U18480 ( .A1(\mem[899][6] ), .A2(n17389), .B1(n26231), .B2(
        data_in[6]), .ZN(n17395) );
  INV_X1 U18481 ( .A(n17396), .ZN(n18907) );
  AOI22_X1 U18482 ( .A1(\mem[899][7] ), .A2(n17389), .B1(n26231), .B2(
        data_in[7]), .ZN(n17396) );
  INV_X1 U18483 ( .A(n17397), .ZN(n18906) );
  AOI22_X1 U18484 ( .A1(\mem[900][0] ), .A2(n17398), .B1(n26230), .B2(
        data_in[0]), .ZN(n17397) );
  INV_X1 U18485 ( .A(n17399), .ZN(n18905) );
  AOI22_X1 U18486 ( .A1(\mem[900][1] ), .A2(n17398), .B1(n26230), .B2(
        data_in[1]), .ZN(n17399) );
  INV_X1 U18487 ( .A(n17400), .ZN(n18904) );
  AOI22_X1 U18488 ( .A1(\mem[900][2] ), .A2(n17398), .B1(n26230), .B2(
        data_in[2]), .ZN(n17400) );
  INV_X1 U18489 ( .A(n17401), .ZN(n18903) );
  AOI22_X1 U18490 ( .A1(\mem[900][3] ), .A2(n17398), .B1(n26230), .B2(
        data_in[3]), .ZN(n17401) );
  INV_X1 U18491 ( .A(n17402), .ZN(n18902) );
  AOI22_X1 U18492 ( .A1(\mem[900][4] ), .A2(n17398), .B1(n26230), .B2(
        data_in[4]), .ZN(n17402) );
  INV_X1 U18493 ( .A(n17403), .ZN(n18901) );
  AOI22_X1 U18494 ( .A1(\mem[900][5] ), .A2(n17398), .B1(n26230), .B2(
        data_in[5]), .ZN(n17403) );
  INV_X1 U18495 ( .A(n17404), .ZN(n18900) );
  AOI22_X1 U18496 ( .A1(\mem[900][6] ), .A2(n17398), .B1(n26230), .B2(
        data_in[6]), .ZN(n17404) );
  INV_X1 U18497 ( .A(n17405), .ZN(n18899) );
  AOI22_X1 U18498 ( .A1(\mem[900][7] ), .A2(n17398), .B1(n26230), .B2(
        data_in[7]), .ZN(n17405) );
  INV_X1 U18499 ( .A(n17406), .ZN(n18898) );
  AOI22_X1 U18500 ( .A1(\mem[901][0] ), .A2(n17407), .B1(n26229), .B2(
        data_in[0]), .ZN(n17406) );
  INV_X1 U18501 ( .A(n17408), .ZN(n18897) );
  AOI22_X1 U18502 ( .A1(\mem[901][1] ), .A2(n17407), .B1(n26229), .B2(
        data_in[1]), .ZN(n17408) );
  INV_X1 U18503 ( .A(n17409), .ZN(n18896) );
  AOI22_X1 U18504 ( .A1(\mem[901][2] ), .A2(n17407), .B1(n26229), .B2(
        data_in[2]), .ZN(n17409) );
  INV_X1 U18505 ( .A(n17410), .ZN(n18895) );
  AOI22_X1 U18506 ( .A1(\mem[901][3] ), .A2(n17407), .B1(n26229), .B2(
        data_in[3]), .ZN(n17410) );
  INV_X1 U18507 ( .A(n17411), .ZN(n18894) );
  AOI22_X1 U18508 ( .A1(\mem[901][4] ), .A2(n17407), .B1(n26229), .B2(
        data_in[4]), .ZN(n17411) );
  INV_X1 U18509 ( .A(n17412), .ZN(n18893) );
  AOI22_X1 U18510 ( .A1(\mem[901][5] ), .A2(n17407), .B1(n26229), .B2(
        data_in[5]), .ZN(n17412) );
  INV_X1 U18511 ( .A(n17413), .ZN(n18892) );
  AOI22_X1 U18512 ( .A1(\mem[901][6] ), .A2(n17407), .B1(n26229), .B2(
        data_in[6]), .ZN(n17413) );
  INV_X1 U18513 ( .A(n17414), .ZN(n18891) );
  AOI22_X1 U18514 ( .A1(\mem[901][7] ), .A2(n17407), .B1(n26229), .B2(
        data_in[7]), .ZN(n17414) );
  INV_X1 U18515 ( .A(n17415), .ZN(n18890) );
  AOI22_X1 U18516 ( .A1(\mem[902][0] ), .A2(n17416), .B1(n26228), .B2(
        data_in[0]), .ZN(n17415) );
  INV_X1 U18517 ( .A(n17417), .ZN(n18889) );
  AOI22_X1 U18518 ( .A1(\mem[902][1] ), .A2(n17416), .B1(n26228), .B2(
        data_in[1]), .ZN(n17417) );
  INV_X1 U18519 ( .A(n17418), .ZN(n18888) );
  AOI22_X1 U18520 ( .A1(\mem[902][2] ), .A2(n17416), .B1(n26228), .B2(
        data_in[2]), .ZN(n17418) );
  INV_X1 U18521 ( .A(n17419), .ZN(n18887) );
  AOI22_X1 U18522 ( .A1(\mem[902][3] ), .A2(n17416), .B1(n26228), .B2(
        data_in[3]), .ZN(n17419) );
  INV_X1 U18523 ( .A(n17420), .ZN(n18886) );
  AOI22_X1 U18524 ( .A1(\mem[902][4] ), .A2(n17416), .B1(n26228), .B2(
        data_in[4]), .ZN(n17420) );
  INV_X1 U18525 ( .A(n17421), .ZN(n18885) );
  AOI22_X1 U18526 ( .A1(\mem[902][5] ), .A2(n17416), .B1(n26228), .B2(
        data_in[5]), .ZN(n17421) );
  INV_X1 U18527 ( .A(n17422), .ZN(n18884) );
  AOI22_X1 U18528 ( .A1(\mem[902][6] ), .A2(n17416), .B1(n26228), .B2(
        data_in[6]), .ZN(n17422) );
  INV_X1 U18529 ( .A(n17423), .ZN(n18883) );
  AOI22_X1 U18530 ( .A1(\mem[902][7] ), .A2(n17416), .B1(n26228), .B2(
        data_in[7]), .ZN(n17423) );
  INV_X1 U18531 ( .A(n17424), .ZN(n18882) );
  AOI22_X1 U18532 ( .A1(\mem[903][0] ), .A2(n17425), .B1(n26227), .B2(
        data_in[0]), .ZN(n17424) );
  INV_X1 U18533 ( .A(n17426), .ZN(n18881) );
  AOI22_X1 U18534 ( .A1(\mem[903][1] ), .A2(n17425), .B1(n26227), .B2(
        data_in[1]), .ZN(n17426) );
  INV_X1 U18535 ( .A(n17427), .ZN(n18880) );
  AOI22_X1 U18536 ( .A1(\mem[903][2] ), .A2(n17425), .B1(n26227), .B2(
        data_in[2]), .ZN(n17427) );
  INV_X1 U18537 ( .A(n17428), .ZN(n18879) );
  AOI22_X1 U18538 ( .A1(\mem[903][3] ), .A2(n17425), .B1(n26227), .B2(
        data_in[3]), .ZN(n17428) );
  INV_X1 U18539 ( .A(n17429), .ZN(n18878) );
  AOI22_X1 U18540 ( .A1(\mem[903][4] ), .A2(n17425), .B1(n26227), .B2(
        data_in[4]), .ZN(n17429) );
  INV_X1 U18541 ( .A(n17430), .ZN(n18877) );
  AOI22_X1 U18542 ( .A1(\mem[903][5] ), .A2(n17425), .B1(n26227), .B2(
        data_in[5]), .ZN(n17430) );
  INV_X1 U18543 ( .A(n17431), .ZN(n18876) );
  AOI22_X1 U18544 ( .A1(\mem[903][6] ), .A2(n17425), .B1(n26227), .B2(
        data_in[6]), .ZN(n17431) );
  INV_X1 U18545 ( .A(n17432), .ZN(n18875) );
  AOI22_X1 U18546 ( .A1(\mem[903][7] ), .A2(n17425), .B1(n26227), .B2(
        data_in[7]), .ZN(n17432) );
  INV_X1 U18547 ( .A(n17649), .ZN(n18682) );
  AOI22_X1 U18548 ( .A1(\mem[928][0] ), .A2(n17650), .B1(n26202), .B2(
        data_in[0]), .ZN(n17649) );
  INV_X1 U18549 ( .A(n17651), .ZN(n18681) );
  AOI22_X1 U18550 ( .A1(\mem[928][1] ), .A2(n17650), .B1(n26202), .B2(
        data_in[1]), .ZN(n17651) );
  INV_X1 U18551 ( .A(n17652), .ZN(n18680) );
  AOI22_X1 U18552 ( .A1(\mem[928][2] ), .A2(n17650), .B1(n26202), .B2(
        data_in[2]), .ZN(n17652) );
  INV_X1 U18553 ( .A(n17653), .ZN(n18679) );
  AOI22_X1 U18554 ( .A1(\mem[928][3] ), .A2(n17650), .B1(n26202), .B2(
        data_in[3]), .ZN(n17653) );
  INV_X1 U18555 ( .A(n17654), .ZN(n18678) );
  AOI22_X1 U18556 ( .A1(\mem[928][4] ), .A2(n17650), .B1(n26202), .B2(
        data_in[4]), .ZN(n17654) );
  INV_X1 U18557 ( .A(n17655), .ZN(n18677) );
  AOI22_X1 U18558 ( .A1(\mem[928][5] ), .A2(n17650), .B1(n26202), .B2(
        data_in[5]), .ZN(n17655) );
  INV_X1 U18559 ( .A(n17656), .ZN(n18676) );
  AOI22_X1 U18560 ( .A1(\mem[928][6] ), .A2(n17650), .B1(n26202), .B2(
        data_in[6]), .ZN(n17656) );
  INV_X1 U18561 ( .A(n17657), .ZN(n18675) );
  AOI22_X1 U18562 ( .A1(\mem[928][7] ), .A2(n17650), .B1(n26202), .B2(
        data_in[7]), .ZN(n17657) );
  INV_X1 U18563 ( .A(n17659), .ZN(n18674) );
  AOI22_X1 U18564 ( .A1(\mem[929][0] ), .A2(n17660), .B1(n26201), .B2(
        data_in[0]), .ZN(n17659) );
  INV_X1 U18565 ( .A(n17661), .ZN(n18673) );
  AOI22_X1 U18566 ( .A1(\mem[929][1] ), .A2(n17660), .B1(n26201), .B2(
        data_in[1]), .ZN(n17661) );
  INV_X1 U18567 ( .A(n17662), .ZN(n18672) );
  AOI22_X1 U18568 ( .A1(\mem[929][2] ), .A2(n17660), .B1(n26201), .B2(
        data_in[2]), .ZN(n17662) );
  INV_X1 U18569 ( .A(n17663), .ZN(n18671) );
  AOI22_X1 U18570 ( .A1(\mem[929][3] ), .A2(n17660), .B1(n26201), .B2(
        data_in[3]), .ZN(n17663) );
  INV_X1 U18571 ( .A(n17664), .ZN(n18670) );
  AOI22_X1 U18572 ( .A1(\mem[929][4] ), .A2(n17660), .B1(n26201), .B2(
        data_in[4]), .ZN(n17664) );
  INV_X1 U18573 ( .A(n17665), .ZN(n18669) );
  AOI22_X1 U18574 ( .A1(\mem[929][5] ), .A2(n17660), .B1(n26201), .B2(
        data_in[5]), .ZN(n17665) );
  INV_X1 U18575 ( .A(n17666), .ZN(n18668) );
  AOI22_X1 U18576 ( .A1(\mem[929][6] ), .A2(n17660), .B1(n26201), .B2(
        data_in[6]), .ZN(n17666) );
  INV_X1 U18577 ( .A(n17667), .ZN(n18667) );
  AOI22_X1 U18578 ( .A1(\mem[929][7] ), .A2(n17660), .B1(n26201), .B2(
        data_in[7]), .ZN(n17667) );
  INV_X1 U18579 ( .A(n17668), .ZN(n18666) );
  AOI22_X1 U18580 ( .A1(\mem[930][0] ), .A2(n17669), .B1(n26200), .B2(
        data_in[0]), .ZN(n17668) );
  INV_X1 U18581 ( .A(n17670), .ZN(n18665) );
  AOI22_X1 U18582 ( .A1(\mem[930][1] ), .A2(n17669), .B1(n26200), .B2(
        data_in[1]), .ZN(n17670) );
  INV_X1 U18583 ( .A(n17671), .ZN(n18664) );
  AOI22_X1 U18584 ( .A1(\mem[930][2] ), .A2(n17669), .B1(n26200), .B2(
        data_in[2]), .ZN(n17671) );
  INV_X1 U18585 ( .A(n17672), .ZN(n18663) );
  AOI22_X1 U18586 ( .A1(\mem[930][3] ), .A2(n17669), .B1(n26200), .B2(
        data_in[3]), .ZN(n17672) );
  INV_X1 U18587 ( .A(n17673), .ZN(n18662) );
  AOI22_X1 U18588 ( .A1(\mem[930][4] ), .A2(n17669), .B1(n26200), .B2(
        data_in[4]), .ZN(n17673) );
  INV_X1 U18589 ( .A(n17674), .ZN(n18661) );
  AOI22_X1 U18590 ( .A1(\mem[930][5] ), .A2(n17669), .B1(n26200), .B2(
        data_in[5]), .ZN(n17674) );
  INV_X1 U18591 ( .A(n17675), .ZN(n18660) );
  AOI22_X1 U18592 ( .A1(\mem[930][6] ), .A2(n17669), .B1(n26200), .B2(
        data_in[6]), .ZN(n17675) );
  INV_X1 U18593 ( .A(n17676), .ZN(n18659) );
  AOI22_X1 U18594 ( .A1(\mem[930][7] ), .A2(n17669), .B1(n26200), .B2(
        data_in[7]), .ZN(n17676) );
  INV_X1 U18595 ( .A(n17677), .ZN(n18658) );
  AOI22_X1 U18596 ( .A1(\mem[931][0] ), .A2(n17678), .B1(n26199), .B2(
        data_in[0]), .ZN(n17677) );
  INV_X1 U18597 ( .A(n17679), .ZN(n18657) );
  AOI22_X1 U18598 ( .A1(\mem[931][1] ), .A2(n17678), .B1(n26199), .B2(
        data_in[1]), .ZN(n17679) );
  INV_X1 U18599 ( .A(n17680), .ZN(n18656) );
  AOI22_X1 U18600 ( .A1(\mem[931][2] ), .A2(n17678), .B1(n26199), .B2(
        data_in[2]), .ZN(n17680) );
  INV_X1 U18601 ( .A(n17681), .ZN(n18655) );
  AOI22_X1 U18602 ( .A1(\mem[931][3] ), .A2(n17678), .B1(n26199), .B2(
        data_in[3]), .ZN(n17681) );
  INV_X1 U18603 ( .A(n17682), .ZN(n18654) );
  AOI22_X1 U18604 ( .A1(\mem[931][4] ), .A2(n17678), .B1(n26199), .B2(
        data_in[4]), .ZN(n17682) );
  INV_X1 U18605 ( .A(n17683), .ZN(n18653) );
  AOI22_X1 U18606 ( .A1(\mem[931][5] ), .A2(n17678), .B1(n26199), .B2(
        data_in[5]), .ZN(n17683) );
  INV_X1 U18607 ( .A(n17684), .ZN(n18652) );
  AOI22_X1 U18608 ( .A1(\mem[931][6] ), .A2(n17678), .B1(n26199), .B2(
        data_in[6]), .ZN(n17684) );
  INV_X1 U18609 ( .A(n17685), .ZN(n18651) );
  AOI22_X1 U18610 ( .A1(\mem[931][7] ), .A2(n17678), .B1(n26199), .B2(
        data_in[7]), .ZN(n17685) );
  INV_X1 U18611 ( .A(n17686), .ZN(n18650) );
  AOI22_X1 U18612 ( .A1(\mem[932][0] ), .A2(n17687), .B1(n26198), .B2(
        data_in[0]), .ZN(n17686) );
  INV_X1 U18613 ( .A(n17688), .ZN(n18649) );
  AOI22_X1 U18614 ( .A1(\mem[932][1] ), .A2(n17687), .B1(n26198), .B2(
        data_in[1]), .ZN(n17688) );
  INV_X1 U18615 ( .A(n17689), .ZN(n18648) );
  AOI22_X1 U18616 ( .A1(\mem[932][2] ), .A2(n17687), .B1(n26198), .B2(
        data_in[2]), .ZN(n17689) );
  INV_X1 U18617 ( .A(n17690), .ZN(n18647) );
  AOI22_X1 U18618 ( .A1(\mem[932][3] ), .A2(n17687), .B1(n26198), .B2(
        data_in[3]), .ZN(n17690) );
  INV_X1 U18619 ( .A(n17691), .ZN(n18646) );
  AOI22_X1 U18620 ( .A1(\mem[932][4] ), .A2(n17687), .B1(n26198), .B2(
        data_in[4]), .ZN(n17691) );
  INV_X1 U18621 ( .A(n17692), .ZN(n18645) );
  AOI22_X1 U18622 ( .A1(\mem[932][5] ), .A2(n17687), .B1(n26198), .B2(
        data_in[5]), .ZN(n17692) );
  INV_X1 U18623 ( .A(n17693), .ZN(n18644) );
  AOI22_X1 U18624 ( .A1(\mem[932][6] ), .A2(n17687), .B1(n26198), .B2(
        data_in[6]), .ZN(n17693) );
  INV_X1 U18625 ( .A(n17694), .ZN(n18643) );
  AOI22_X1 U18626 ( .A1(\mem[932][7] ), .A2(n17687), .B1(n26198), .B2(
        data_in[7]), .ZN(n17694) );
  INV_X1 U18627 ( .A(n17695), .ZN(n18642) );
  AOI22_X1 U18628 ( .A1(\mem[933][0] ), .A2(n17696), .B1(n26197), .B2(
        data_in[0]), .ZN(n17695) );
  INV_X1 U18629 ( .A(n17697), .ZN(n18641) );
  AOI22_X1 U18630 ( .A1(\mem[933][1] ), .A2(n17696), .B1(n26197), .B2(
        data_in[1]), .ZN(n17697) );
  INV_X1 U18631 ( .A(n17698), .ZN(n18640) );
  AOI22_X1 U18632 ( .A1(\mem[933][2] ), .A2(n17696), .B1(n26197), .B2(
        data_in[2]), .ZN(n17698) );
  INV_X1 U18633 ( .A(n17699), .ZN(n18639) );
  AOI22_X1 U18634 ( .A1(\mem[933][3] ), .A2(n17696), .B1(n26197), .B2(
        data_in[3]), .ZN(n17699) );
  INV_X1 U18635 ( .A(n17700), .ZN(n18638) );
  AOI22_X1 U18636 ( .A1(\mem[933][4] ), .A2(n17696), .B1(n26197), .B2(
        data_in[4]), .ZN(n17700) );
  INV_X1 U18637 ( .A(n17701), .ZN(n18637) );
  AOI22_X1 U18638 ( .A1(\mem[933][5] ), .A2(n17696), .B1(n26197), .B2(
        data_in[5]), .ZN(n17701) );
  INV_X1 U18639 ( .A(n17702), .ZN(n18636) );
  AOI22_X1 U18640 ( .A1(\mem[933][6] ), .A2(n17696), .B1(n26197), .B2(
        data_in[6]), .ZN(n17702) );
  INV_X1 U18641 ( .A(n17703), .ZN(n18635) );
  AOI22_X1 U18642 ( .A1(\mem[933][7] ), .A2(n17696), .B1(n26197), .B2(
        data_in[7]), .ZN(n17703) );
  INV_X1 U18643 ( .A(n17704), .ZN(n18634) );
  AOI22_X1 U18644 ( .A1(\mem[934][0] ), .A2(n17705), .B1(n26196), .B2(
        data_in[0]), .ZN(n17704) );
  INV_X1 U18645 ( .A(n17706), .ZN(n18633) );
  AOI22_X1 U18646 ( .A1(\mem[934][1] ), .A2(n17705), .B1(n26196), .B2(
        data_in[1]), .ZN(n17706) );
  INV_X1 U18647 ( .A(n17707), .ZN(n18632) );
  AOI22_X1 U18648 ( .A1(\mem[934][2] ), .A2(n17705), .B1(n26196), .B2(
        data_in[2]), .ZN(n17707) );
  INV_X1 U18649 ( .A(n17708), .ZN(n18631) );
  AOI22_X1 U18650 ( .A1(\mem[934][3] ), .A2(n17705), .B1(n26196), .B2(
        data_in[3]), .ZN(n17708) );
  INV_X1 U18651 ( .A(n17709), .ZN(n18630) );
  AOI22_X1 U18652 ( .A1(\mem[934][4] ), .A2(n17705), .B1(n26196), .B2(
        data_in[4]), .ZN(n17709) );
  INV_X1 U18653 ( .A(n17710), .ZN(n18629) );
  AOI22_X1 U18654 ( .A1(\mem[934][5] ), .A2(n17705), .B1(n26196), .B2(
        data_in[5]), .ZN(n17710) );
  INV_X1 U18655 ( .A(n17711), .ZN(n18628) );
  AOI22_X1 U18656 ( .A1(\mem[934][6] ), .A2(n17705), .B1(n26196), .B2(
        data_in[6]), .ZN(n17711) );
  INV_X1 U18657 ( .A(n17712), .ZN(n18627) );
  AOI22_X1 U18658 ( .A1(\mem[934][7] ), .A2(n17705), .B1(n26196), .B2(
        data_in[7]), .ZN(n17712) );
  INV_X1 U18659 ( .A(n17713), .ZN(n18626) );
  AOI22_X1 U18660 ( .A1(\mem[935][0] ), .A2(n17714), .B1(n26195), .B2(
        data_in[0]), .ZN(n17713) );
  INV_X1 U18661 ( .A(n17715), .ZN(n18625) );
  AOI22_X1 U18662 ( .A1(\mem[935][1] ), .A2(n17714), .B1(n26195), .B2(
        data_in[1]), .ZN(n17715) );
  INV_X1 U18663 ( .A(n17716), .ZN(n18624) );
  AOI22_X1 U18664 ( .A1(\mem[935][2] ), .A2(n17714), .B1(n26195), .B2(
        data_in[2]), .ZN(n17716) );
  INV_X1 U18665 ( .A(n17717), .ZN(n18623) );
  AOI22_X1 U18666 ( .A1(\mem[935][3] ), .A2(n17714), .B1(n26195), .B2(
        data_in[3]), .ZN(n17717) );
  INV_X1 U18667 ( .A(n17718), .ZN(n18622) );
  AOI22_X1 U18668 ( .A1(\mem[935][4] ), .A2(n17714), .B1(n26195), .B2(
        data_in[4]), .ZN(n17718) );
  INV_X1 U18669 ( .A(n17719), .ZN(n18621) );
  AOI22_X1 U18670 ( .A1(\mem[935][5] ), .A2(n17714), .B1(n26195), .B2(
        data_in[5]), .ZN(n17719) );
  INV_X1 U18671 ( .A(n17720), .ZN(n18620) );
  AOI22_X1 U18672 ( .A1(\mem[935][6] ), .A2(n17714), .B1(n26195), .B2(
        data_in[6]), .ZN(n17720) );
  INV_X1 U18673 ( .A(n17721), .ZN(n18619) );
  AOI22_X1 U18674 ( .A1(\mem[935][7] ), .A2(n17714), .B1(n26195), .B2(
        data_in[7]), .ZN(n17721) );
  INV_X1 U18675 ( .A(n17938), .ZN(n9120) );
  AOI22_X1 U18676 ( .A1(\mem[960][0] ), .A2(n17939), .B1(n26170), .B2(
        data_in[0]), .ZN(n17938) );
  INV_X1 U18677 ( .A(n17940), .ZN(n9119) );
  AOI22_X1 U18678 ( .A1(\mem[960][1] ), .A2(n17939), .B1(n26170), .B2(
        data_in[1]), .ZN(n17940) );
  INV_X1 U18679 ( .A(n17941), .ZN(n9118) );
  AOI22_X1 U18680 ( .A1(\mem[960][2] ), .A2(n17939), .B1(n26170), .B2(
        data_in[2]), .ZN(n17941) );
  INV_X1 U18681 ( .A(n17942), .ZN(n9117) );
  AOI22_X1 U18682 ( .A1(\mem[960][3] ), .A2(n17939), .B1(n26170), .B2(
        data_in[3]), .ZN(n17942) );
  INV_X1 U18683 ( .A(n17943), .ZN(n9116) );
  AOI22_X1 U18684 ( .A1(\mem[960][4] ), .A2(n17939), .B1(n26170), .B2(
        data_in[4]), .ZN(n17943) );
  INV_X1 U18685 ( .A(n17944), .ZN(n9115) );
  AOI22_X1 U18686 ( .A1(\mem[960][5] ), .A2(n17939), .B1(n26170), .B2(
        data_in[5]), .ZN(n17944) );
  INV_X1 U18687 ( .A(n17945), .ZN(n9114) );
  AOI22_X1 U18688 ( .A1(\mem[960][6] ), .A2(n17939), .B1(n26170), .B2(
        data_in[6]), .ZN(n17945) );
  INV_X1 U18689 ( .A(n17946), .ZN(n9113) );
  AOI22_X1 U18690 ( .A1(\mem[960][7] ), .A2(n17939), .B1(n26170), .B2(
        data_in[7]), .ZN(n17946) );
  INV_X1 U18691 ( .A(n17948), .ZN(n9112) );
  AOI22_X1 U18692 ( .A1(\mem[961][0] ), .A2(n17949), .B1(n26169), .B2(
        data_in[0]), .ZN(n17948) );
  INV_X1 U18693 ( .A(n17950), .ZN(n9111) );
  AOI22_X1 U18694 ( .A1(\mem[961][1] ), .A2(n17949), .B1(n26169), .B2(
        data_in[1]), .ZN(n17950) );
  INV_X1 U18695 ( .A(n17951), .ZN(n9110) );
  AOI22_X1 U18696 ( .A1(\mem[961][2] ), .A2(n17949), .B1(n26169), .B2(
        data_in[2]), .ZN(n17951) );
  INV_X1 U18697 ( .A(n17952), .ZN(n9109) );
  AOI22_X1 U18698 ( .A1(\mem[961][3] ), .A2(n17949), .B1(n26169), .B2(
        data_in[3]), .ZN(n17952) );
  INV_X1 U18699 ( .A(n17953), .ZN(n9108) );
  AOI22_X1 U18700 ( .A1(\mem[961][4] ), .A2(n17949), .B1(n26169), .B2(
        data_in[4]), .ZN(n17953) );
  INV_X1 U18701 ( .A(n17954), .ZN(n9107) );
  AOI22_X1 U18702 ( .A1(\mem[961][5] ), .A2(n17949), .B1(n26169), .B2(
        data_in[5]), .ZN(n17954) );
  INV_X1 U18703 ( .A(n17955), .ZN(n9106) );
  AOI22_X1 U18704 ( .A1(\mem[961][6] ), .A2(n17949), .B1(n26169), .B2(
        data_in[6]), .ZN(n17955) );
  INV_X1 U18705 ( .A(n17956), .ZN(n9105) );
  AOI22_X1 U18706 ( .A1(\mem[961][7] ), .A2(n17949), .B1(n26169), .B2(
        data_in[7]), .ZN(n17956) );
  INV_X1 U18707 ( .A(n17957), .ZN(n9104) );
  AOI22_X1 U18708 ( .A1(\mem[962][0] ), .A2(n17958), .B1(n26168), .B2(
        data_in[0]), .ZN(n17957) );
  INV_X1 U18709 ( .A(n17959), .ZN(n9103) );
  AOI22_X1 U18710 ( .A1(\mem[962][1] ), .A2(n17958), .B1(n26168), .B2(
        data_in[1]), .ZN(n17959) );
  INV_X1 U18711 ( .A(n17960), .ZN(n9102) );
  AOI22_X1 U18712 ( .A1(\mem[962][2] ), .A2(n17958), .B1(n26168), .B2(
        data_in[2]), .ZN(n17960) );
  INV_X1 U18713 ( .A(n17961), .ZN(n9101) );
  AOI22_X1 U18714 ( .A1(\mem[962][3] ), .A2(n17958), .B1(n26168), .B2(
        data_in[3]), .ZN(n17961) );
  INV_X1 U18715 ( .A(n17962), .ZN(n9100) );
  AOI22_X1 U18716 ( .A1(\mem[962][4] ), .A2(n17958), .B1(n26168), .B2(
        data_in[4]), .ZN(n17962) );
  INV_X1 U18717 ( .A(n17963), .ZN(n9099) );
  AOI22_X1 U18718 ( .A1(\mem[962][5] ), .A2(n17958), .B1(n26168), .B2(
        data_in[5]), .ZN(n17963) );
  INV_X1 U18719 ( .A(n17964), .ZN(n9098) );
  AOI22_X1 U18720 ( .A1(\mem[962][6] ), .A2(n17958), .B1(n26168), .B2(
        data_in[6]), .ZN(n17964) );
  INV_X1 U18721 ( .A(n17965), .ZN(n9097) );
  AOI22_X1 U18722 ( .A1(\mem[962][7] ), .A2(n17958), .B1(n26168), .B2(
        data_in[7]), .ZN(n17965) );
  INV_X1 U18723 ( .A(n17966), .ZN(n9096) );
  AOI22_X1 U18724 ( .A1(\mem[963][0] ), .A2(n17967), .B1(n26167), .B2(
        data_in[0]), .ZN(n17966) );
  INV_X1 U18725 ( .A(n17968), .ZN(n9095) );
  AOI22_X1 U18726 ( .A1(\mem[963][1] ), .A2(n17967), .B1(n26167), .B2(
        data_in[1]), .ZN(n17968) );
  INV_X1 U18727 ( .A(n17969), .ZN(n9094) );
  AOI22_X1 U18728 ( .A1(\mem[963][2] ), .A2(n17967), .B1(n26167), .B2(
        data_in[2]), .ZN(n17969) );
  INV_X1 U18729 ( .A(n17970), .ZN(n9093) );
  AOI22_X1 U18730 ( .A1(\mem[963][3] ), .A2(n17967), .B1(n26167), .B2(
        data_in[3]), .ZN(n17970) );
  INV_X1 U18731 ( .A(n17971), .ZN(n9092) );
  AOI22_X1 U18732 ( .A1(\mem[963][4] ), .A2(n17967), .B1(n26167), .B2(
        data_in[4]), .ZN(n17971) );
  INV_X1 U18733 ( .A(n17972), .ZN(n9091) );
  AOI22_X1 U18734 ( .A1(\mem[963][5] ), .A2(n17967), .B1(n26167), .B2(
        data_in[5]), .ZN(n17972) );
  INV_X1 U18735 ( .A(n17973), .ZN(n9090) );
  AOI22_X1 U18736 ( .A1(\mem[963][6] ), .A2(n17967), .B1(n26167), .B2(
        data_in[6]), .ZN(n17973) );
  INV_X1 U18737 ( .A(n17974), .ZN(n9089) );
  AOI22_X1 U18738 ( .A1(\mem[963][7] ), .A2(n17967), .B1(n26167), .B2(
        data_in[7]), .ZN(n17974) );
  INV_X1 U18739 ( .A(n17975), .ZN(n9088) );
  AOI22_X1 U18740 ( .A1(\mem[964][0] ), .A2(n17976), .B1(n26166), .B2(
        data_in[0]), .ZN(n17975) );
  INV_X1 U18741 ( .A(n17977), .ZN(n9087) );
  AOI22_X1 U18742 ( .A1(\mem[964][1] ), .A2(n17976), .B1(n26166), .B2(
        data_in[1]), .ZN(n17977) );
  INV_X1 U18743 ( .A(n17978), .ZN(n9086) );
  AOI22_X1 U18744 ( .A1(\mem[964][2] ), .A2(n17976), .B1(n26166), .B2(
        data_in[2]), .ZN(n17978) );
  INV_X1 U18745 ( .A(n17979), .ZN(n9085) );
  AOI22_X1 U18746 ( .A1(\mem[964][3] ), .A2(n17976), .B1(n26166), .B2(
        data_in[3]), .ZN(n17979) );
  INV_X1 U18747 ( .A(n17980), .ZN(n9084) );
  AOI22_X1 U18748 ( .A1(\mem[964][4] ), .A2(n17976), .B1(n26166), .B2(
        data_in[4]), .ZN(n17980) );
  INV_X1 U18749 ( .A(n17981), .ZN(n9083) );
  AOI22_X1 U18750 ( .A1(\mem[964][5] ), .A2(n17976), .B1(n26166), .B2(
        data_in[5]), .ZN(n17981) );
  INV_X1 U18751 ( .A(n17982), .ZN(n9082) );
  AOI22_X1 U18752 ( .A1(\mem[964][6] ), .A2(n17976), .B1(n26166), .B2(
        data_in[6]), .ZN(n17982) );
  INV_X1 U18753 ( .A(n17983), .ZN(n9081) );
  AOI22_X1 U18754 ( .A1(\mem[964][7] ), .A2(n17976), .B1(n26166), .B2(
        data_in[7]), .ZN(n17983) );
  INV_X1 U18755 ( .A(n17984), .ZN(n9080) );
  AOI22_X1 U18756 ( .A1(\mem[965][0] ), .A2(n17985), .B1(n26165), .B2(
        data_in[0]), .ZN(n17984) );
  INV_X1 U18757 ( .A(n17986), .ZN(n9079) );
  AOI22_X1 U18758 ( .A1(\mem[965][1] ), .A2(n17985), .B1(n26165), .B2(
        data_in[1]), .ZN(n17986) );
  INV_X1 U18759 ( .A(n17987), .ZN(n9078) );
  AOI22_X1 U18760 ( .A1(\mem[965][2] ), .A2(n17985), .B1(n26165), .B2(
        data_in[2]), .ZN(n17987) );
  INV_X1 U18761 ( .A(n17988), .ZN(n9077) );
  AOI22_X1 U18762 ( .A1(\mem[965][3] ), .A2(n17985), .B1(n26165), .B2(
        data_in[3]), .ZN(n17988) );
  INV_X1 U18763 ( .A(n17989), .ZN(n9076) );
  AOI22_X1 U18764 ( .A1(\mem[965][4] ), .A2(n17985), .B1(n26165), .B2(
        data_in[4]), .ZN(n17989) );
  INV_X1 U18765 ( .A(n17990), .ZN(n9075) );
  AOI22_X1 U18766 ( .A1(\mem[965][5] ), .A2(n17985), .B1(n26165), .B2(
        data_in[5]), .ZN(n17990) );
  INV_X1 U18767 ( .A(n17991), .ZN(n9074) );
  AOI22_X1 U18768 ( .A1(\mem[965][6] ), .A2(n17985), .B1(n26165), .B2(
        data_in[6]), .ZN(n17991) );
  INV_X1 U18769 ( .A(n17992), .ZN(n9073) );
  AOI22_X1 U18770 ( .A1(\mem[965][7] ), .A2(n17985), .B1(n26165), .B2(
        data_in[7]), .ZN(n17992) );
  INV_X1 U18771 ( .A(n17993), .ZN(n9072) );
  AOI22_X1 U18772 ( .A1(\mem[966][0] ), .A2(n17994), .B1(n26164), .B2(
        data_in[0]), .ZN(n17993) );
  INV_X1 U18773 ( .A(n17995), .ZN(n9071) );
  AOI22_X1 U18774 ( .A1(\mem[966][1] ), .A2(n17994), .B1(n26164), .B2(
        data_in[1]), .ZN(n17995) );
  INV_X1 U18775 ( .A(n17996), .ZN(n9070) );
  AOI22_X1 U18776 ( .A1(\mem[966][2] ), .A2(n17994), .B1(n26164), .B2(
        data_in[2]), .ZN(n17996) );
  INV_X1 U18777 ( .A(n17997), .ZN(n9069) );
  AOI22_X1 U18778 ( .A1(\mem[966][3] ), .A2(n17994), .B1(n26164), .B2(
        data_in[3]), .ZN(n17997) );
  INV_X1 U18779 ( .A(n17998), .ZN(n9068) );
  AOI22_X1 U18780 ( .A1(\mem[966][4] ), .A2(n17994), .B1(n26164), .B2(
        data_in[4]), .ZN(n17998) );
  INV_X1 U18781 ( .A(n17999), .ZN(n9067) );
  AOI22_X1 U18782 ( .A1(\mem[966][5] ), .A2(n17994), .B1(n26164), .B2(
        data_in[5]), .ZN(n17999) );
  INV_X1 U18783 ( .A(n18000), .ZN(n9066) );
  AOI22_X1 U18784 ( .A1(\mem[966][6] ), .A2(n17994), .B1(n26164), .B2(
        data_in[6]), .ZN(n18000) );
  INV_X1 U18785 ( .A(n18001), .ZN(n9065) );
  AOI22_X1 U18786 ( .A1(\mem[966][7] ), .A2(n17994), .B1(n26164), .B2(
        data_in[7]), .ZN(n18001) );
  INV_X1 U18787 ( .A(n18002), .ZN(n9064) );
  AOI22_X1 U18788 ( .A1(\mem[967][0] ), .A2(n18003), .B1(n26163), .B2(
        data_in[0]), .ZN(n18002) );
  INV_X1 U18789 ( .A(n18004), .ZN(n9063) );
  AOI22_X1 U18790 ( .A1(\mem[967][1] ), .A2(n18003), .B1(n26163), .B2(
        data_in[1]), .ZN(n18004) );
  INV_X1 U18791 ( .A(n18005), .ZN(n9062) );
  AOI22_X1 U18792 ( .A1(\mem[967][2] ), .A2(n18003), .B1(n26163), .B2(
        data_in[2]), .ZN(n18005) );
  INV_X1 U18793 ( .A(n18006), .ZN(n9061) );
  AOI22_X1 U18794 ( .A1(\mem[967][3] ), .A2(n18003), .B1(n26163), .B2(
        data_in[3]), .ZN(n18006) );
  INV_X1 U18795 ( .A(n18007), .ZN(n9060) );
  AOI22_X1 U18796 ( .A1(\mem[967][4] ), .A2(n18003), .B1(n26163), .B2(
        data_in[4]), .ZN(n18007) );
  INV_X1 U18797 ( .A(n18008), .ZN(n9059) );
  AOI22_X1 U18798 ( .A1(\mem[967][5] ), .A2(n18003), .B1(n26163), .B2(
        data_in[5]), .ZN(n18008) );
  INV_X1 U18799 ( .A(n18009), .ZN(n9058) );
  AOI22_X1 U18800 ( .A1(\mem[967][6] ), .A2(n18003), .B1(n26163), .B2(
        data_in[6]), .ZN(n18009) );
  INV_X1 U18801 ( .A(n18010), .ZN(n9057) );
  AOI22_X1 U18802 ( .A1(\mem[967][7] ), .A2(n18003), .B1(n26163), .B2(
        data_in[7]), .ZN(n18010) );
  INV_X1 U18803 ( .A(n18227), .ZN(n8864) );
  AOI22_X1 U18804 ( .A1(\mem[992][0] ), .A2(n18228), .B1(n26138), .B2(
        data_in[0]), .ZN(n18227) );
  INV_X1 U18805 ( .A(n18229), .ZN(n8863) );
  AOI22_X1 U18806 ( .A1(\mem[992][1] ), .A2(n18228), .B1(n26138), .B2(
        data_in[1]), .ZN(n18229) );
  INV_X1 U18807 ( .A(n18230), .ZN(n8862) );
  AOI22_X1 U18808 ( .A1(\mem[992][2] ), .A2(n18228), .B1(n26138), .B2(
        data_in[2]), .ZN(n18230) );
  INV_X1 U18809 ( .A(n18231), .ZN(n8861) );
  AOI22_X1 U18810 ( .A1(\mem[992][3] ), .A2(n18228), .B1(n26138), .B2(
        data_in[3]), .ZN(n18231) );
  INV_X1 U18811 ( .A(n18232), .ZN(n8860) );
  AOI22_X1 U18812 ( .A1(\mem[992][4] ), .A2(n18228), .B1(n26138), .B2(
        data_in[4]), .ZN(n18232) );
  INV_X1 U18813 ( .A(n18233), .ZN(n8859) );
  AOI22_X1 U18814 ( .A1(\mem[992][5] ), .A2(n18228), .B1(n26138), .B2(
        data_in[5]), .ZN(n18233) );
  INV_X1 U18815 ( .A(n18234), .ZN(n8858) );
  AOI22_X1 U18816 ( .A1(\mem[992][6] ), .A2(n18228), .B1(n26138), .B2(
        data_in[6]), .ZN(n18234) );
  INV_X1 U18817 ( .A(n18235), .ZN(n8857) );
  AOI22_X1 U18818 ( .A1(\mem[992][7] ), .A2(n18228), .B1(n26138), .B2(
        data_in[7]), .ZN(n18235) );
  INV_X1 U18819 ( .A(n18239), .ZN(n8856) );
  AOI22_X1 U18820 ( .A1(\mem[993][0] ), .A2(n18240), .B1(n26137), .B2(
        data_in[0]), .ZN(n18239) );
  INV_X1 U18821 ( .A(n18241), .ZN(n8855) );
  AOI22_X1 U18822 ( .A1(\mem[993][1] ), .A2(n18240), .B1(n26137), .B2(
        data_in[1]), .ZN(n18241) );
  INV_X1 U18823 ( .A(n18242), .ZN(n8854) );
  AOI22_X1 U18824 ( .A1(\mem[993][2] ), .A2(n18240), .B1(n26137), .B2(
        data_in[2]), .ZN(n18242) );
  INV_X1 U18825 ( .A(n18243), .ZN(n8853) );
  AOI22_X1 U18826 ( .A1(\mem[993][3] ), .A2(n18240), .B1(n26137), .B2(
        data_in[3]), .ZN(n18243) );
  INV_X1 U18827 ( .A(n18244), .ZN(n8852) );
  AOI22_X1 U18828 ( .A1(\mem[993][4] ), .A2(n18240), .B1(n26137), .B2(
        data_in[4]), .ZN(n18244) );
  INV_X1 U18829 ( .A(n18245), .ZN(n8851) );
  AOI22_X1 U18830 ( .A1(\mem[993][5] ), .A2(n18240), .B1(n26137), .B2(
        data_in[5]), .ZN(n18245) );
  INV_X1 U18831 ( .A(n18246), .ZN(n8850) );
  AOI22_X1 U18832 ( .A1(\mem[993][6] ), .A2(n18240), .B1(n26137), .B2(
        data_in[6]), .ZN(n18246) );
  INV_X1 U18833 ( .A(n18247), .ZN(n8849) );
  AOI22_X1 U18834 ( .A1(\mem[993][7] ), .A2(n18240), .B1(n26137), .B2(
        data_in[7]), .ZN(n18247) );
  INV_X1 U18835 ( .A(n18249), .ZN(n8848) );
  AOI22_X1 U18836 ( .A1(\mem[994][0] ), .A2(n18250), .B1(n26136), .B2(
        data_in[0]), .ZN(n18249) );
  INV_X1 U18837 ( .A(n18251), .ZN(n8847) );
  AOI22_X1 U18838 ( .A1(\mem[994][1] ), .A2(n18250), .B1(n26136), .B2(
        data_in[1]), .ZN(n18251) );
  INV_X1 U18839 ( .A(n18252), .ZN(n8846) );
  AOI22_X1 U18840 ( .A1(\mem[994][2] ), .A2(n18250), .B1(n26136), .B2(
        data_in[2]), .ZN(n18252) );
  INV_X1 U18841 ( .A(n18253), .ZN(n8845) );
  AOI22_X1 U18842 ( .A1(\mem[994][3] ), .A2(n18250), .B1(n26136), .B2(
        data_in[3]), .ZN(n18253) );
  INV_X1 U18843 ( .A(n18254), .ZN(n8844) );
  AOI22_X1 U18844 ( .A1(\mem[994][4] ), .A2(n18250), .B1(n26136), .B2(
        data_in[4]), .ZN(n18254) );
  INV_X1 U18845 ( .A(n18255), .ZN(n8843) );
  AOI22_X1 U18846 ( .A1(\mem[994][5] ), .A2(n18250), .B1(n26136), .B2(
        data_in[5]), .ZN(n18255) );
  INV_X1 U18847 ( .A(n18256), .ZN(n8842) );
  AOI22_X1 U18848 ( .A1(\mem[994][6] ), .A2(n18250), .B1(n26136), .B2(
        data_in[6]), .ZN(n18256) );
  INV_X1 U18849 ( .A(n18257), .ZN(n8841) );
  AOI22_X1 U18850 ( .A1(\mem[994][7] ), .A2(n18250), .B1(n26136), .B2(
        data_in[7]), .ZN(n18257) );
  INV_X1 U18851 ( .A(n18259), .ZN(n8840) );
  AOI22_X1 U18852 ( .A1(\mem[995][0] ), .A2(n18260), .B1(n26135), .B2(
        data_in[0]), .ZN(n18259) );
  INV_X1 U18853 ( .A(n18261), .ZN(n8839) );
  AOI22_X1 U18854 ( .A1(\mem[995][1] ), .A2(n18260), .B1(n26135), .B2(
        data_in[1]), .ZN(n18261) );
  INV_X1 U18855 ( .A(n18262), .ZN(n8838) );
  AOI22_X1 U18856 ( .A1(\mem[995][2] ), .A2(n18260), .B1(n26135), .B2(
        data_in[2]), .ZN(n18262) );
  INV_X1 U18857 ( .A(n18263), .ZN(n8837) );
  AOI22_X1 U18858 ( .A1(\mem[995][3] ), .A2(n18260), .B1(n26135), .B2(
        data_in[3]), .ZN(n18263) );
  INV_X1 U18859 ( .A(n18264), .ZN(n8836) );
  AOI22_X1 U18860 ( .A1(\mem[995][4] ), .A2(n18260), .B1(n26135), .B2(
        data_in[4]), .ZN(n18264) );
  INV_X1 U18861 ( .A(n18265), .ZN(n8835) );
  AOI22_X1 U18862 ( .A1(\mem[995][5] ), .A2(n18260), .B1(n26135), .B2(
        data_in[5]), .ZN(n18265) );
  INV_X1 U18863 ( .A(n18266), .ZN(n8834) );
  AOI22_X1 U18864 ( .A1(\mem[995][6] ), .A2(n18260), .B1(n26135), .B2(
        data_in[6]), .ZN(n18266) );
  INV_X1 U18865 ( .A(n18267), .ZN(n8833) );
  AOI22_X1 U18866 ( .A1(\mem[995][7] ), .A2(n18260), .B1(n26135), .B2(
        data_in[7]), .ZN(n18267) );
  INV_X1 U18867 ( .A(n18269), .ZN(n8832) );
  AOI22_X1 U18868 ( .A1(\mem[996][0] ), .A2(n18270), .B1(n26134), .B2(
        data_in[0]), .ZN(n18269) );
  INV_X1 U18869 ( .A(n18271), .ZN(n8831) );
  AOI22_X1 U18870 ( .A1(\mem[996][1] ), .A2(n18270), .B1(n26134), .B2(
        data_in[1]), .ZN(n18271) );
  INV_X1 U18871 ( .A(n18272), .ZN(n8830) );
  AOI22_X1 U18872 ( .A1(\mem[996][2] ), .A2(n18270), .B1(n26134), .B2(
        data_in[2]), .ZN(n18272) );
  INV_X1 U18873 ( .A(n18273), .ZN(n8829) );
  AOI22_X1 U18874 ( .A1(\mem[996][3] ), .A2(n18270), .B1(n26134), .B2(
        data_in[3]), .ZN(n18273) );
  INV_X1 U18875 ( .A(n18274), .ZN(n8828) );
  AOI22_X1 U18876 ( .A1(\mem[996][4] ), .A2(n18270), .B1(n26134), .B2(
        data_in[4]), .ZN(n18274) );
  INV_X1 U18877 ( .A(n18275), .ZN(n8827) );
  AOI22_X1 U18878 ( .A1(\mem[996][5] ), .A2(n18270), .B1(n26134), .B2(
        data_in[5]), .ZN(n18275) );
  INV_X1 U18879 ( .A(n18276), .ZN(n8826) );
  AOI22_X1 U18880 ( .A1(\mem[996][6] ), .A2(n18270), .B1(n26134), .B2(
        data_in[6]), .ZN(n18276) );
  INV_X1 U18881 ( .A(n18277), .ZN(n8825) );
  AOI22_X1 U18882 ( .A1(\mem[996][7] ), .A2(n18270), .B1(n26134), .B2(
        data_in[7]), .ZN(n18277) );
  INV_X1 U18883 ( .A(n18279), .ZN(n8824) );
  AOI22_X1 U18884 ( .A1(\mem[997][0] ), .A2(n18280), .B1(n26133), .B2(
        data_in[0]), .ZN(n18279) );
  INV_X1 U18885 ( .A(n18281), .ZN(n8823) );
  AOI22_X1 U18886 ( .A1(\mem[997][1] ), .A2(n18280), .B1(n26133), .B2(
        data_in[1]), .ZN(n18281) );
  INV_X1 U18887 ( .A(n18282), .ZN(n8822) );
  AOI22_X1 U18888 ( .A1(\mem[997][2] ), .A2(n18280), .B1(n26133), .B2(
        data_in[2]), .ZN(n18282) );
  INV_X1 U18889 ( .A(n18283), .ZN(n8821) );
  AOI22_X1 U18890 ( .A1(\mem[997][3] ), .A2(n18280), .B1(n26133), .B2(
        data_in[3]), .ZN(n18283) );
  INV_X1 U18891 ( .A(n18284), .ZN(n8820) );
  AOI22_X1 U18892 ( .A1(\mem[997][4] ), .A2(n18280), .B1(n26133), .B2(
        data_in[4]), .ZN(n18284) );
  INV_X1 U18893 ( .A(n18285), .ZN(n8819) );
  AOI22_X1 U18894 ( .A1(\mem[997][5] ), .A2(n18280), .B1(n26133), .B2(
        data_in[5]), .ZN(n18285) );
  INV_X1 U18895 ( .A(n18286), .ZN(n8818) );
  AOI22_X1 U18896 ( .A1(\mem[997][6] ), .A2(n18280), .B1(n26133), .B2(
        data_in[6]), .ZN(n18286) );
  INV_X1 U18897 ( .A(n18287), .ZN(n8817) );
  AOI22_X1 U18898 ( .A1(\mem[997][7] ), .A2(n18280), .B1(n26133), .B2(
        data_in[7]), .ZN(n18287) );
  INV_X1 U18899 ( .A(n18289), .ZN(n8816) );
  AOI22_X1 U18900 ( .A1(\mem[998][0] ), .A2(n18290), .B1(n26132), .B2(
        data_in[0]), .ZN(n18289) );
  INV_X1 U18901 ( .A(n18291), .ZN(n8815) );
  AOI22_X1 U18902 ( .A1(\mem[998][1] ), .A2(n18290), .B1(n26132), .B2(
        data_in[1]), .ZN(n18291) );
  INV_X1 U18903 ( .A(n18292), .ZN(n8814) );
  AOI22_X1 U18904 ( .A1(\mem[998][2] ), .A2(n18290), .B1(n26132), .B2(
        data_in[2]), .ZN(n18292) );
  INV_X1 U18905 ( .A(n18293), .ZN(n8813) );
  AOI22_X1 U18906 ( .A1(\mem[998][3] ), .A2(n18290), .B1(n26132), .B2(
        data_in[3]), .ZN(n18293) );
  INV_X1 U18907 ( .A(n18294), .ZN(n8812) );
  AOI22_X1 U18908 ( .A1(\mem[998][4] ), .A2(n18290), .B1(n26132), .B2(
        data_in[4]), .ZN(n18294) );
  INV_X1 U18909 ( .A(n18295), .ZN(n8811) );
  AOI22_X1 U18910 ( .A1(\mem[998][5] ), .A2(n18290), .B1(n26132), .B2(
        data_in[5]), .ZN(n18295) );
  INV_X1 U18911 ( .A(n18296), .ZN(n8810) );
  AOI22_X1 U18912 ( .A1(\mem[998][6] ), .A2(n18290), .B1(n26132), .B2(
        data_in[6]), .ZN(n18296) );
  INV_X1 U18913 ( .A(n18297), .ZN(n8809) );
  AOI22_X1 U18914 ( .A1(\mem[998][7] ), .A2(n18290), .B1(n26132), .B2(
        data_in[7]), .ZN(n18297) );
  INV_X1 U18915 ( .A(n18299), .ZN(n8808) );
  AOI22_X1 U18916 ( .A1(\mem[999][0] ), .A2(n18300), .B1(n26131), .B2(
        data_in[0]), .ZN(n18299) );
  INV_X1 U18917 ( .A(n18301), .ZN(n8807) );
  AOI22_X1 U18918 ( .A1(\mem[999][1] ), .A2(n18300), .B1(n26131), .B2(
        data_in[1]), .ZN(n18301) );
  INV_X1 U18919 ( .A(n18302), .ZN(n8806) );
  AOI22_X1 U18920 ( .A1(\mem[999][2] ), .A2(n18300), .B1(n26131), .B2(
        data_in[2]), .ZN(n18302) );
  INV_X1 U18921 ( .A(n18303), .ZN(n8805) );
  AOI22_X1 U18922 ( .A1(\mem[999][3] ), .A2(n18300), .B1(n26131), .B2(
        data_in[3]), .ZN(n18303) );
  INV_X1 U18923 ( .A(n18304), .ZN(n8804) );
  AOI22_X1 U18924 ( .A1(\mem[999][4] ), .A2(n18300), .B1(n26131), .B2(
        data_in[4]), .ZN(n18304) );
  INV_X1 U18925 ( .A(n18305), .ZN(n8803) );
  AOI22_X1 U18926 ( .A1(\mem[999][5] ), .A2(n18300), .B1(n26131), .B2(
        data_in[5]), .ZN(n18305) );
  INV_X1 U18927 ( .A(n18306), .ZN(n8802) );
  AOI22_X1 U18928 ( .A1(\mem[999][6] ), .A2(n18300), .B1(n26131), .B2(
        data_in[6]), .ZN(n18306) );
  INV_X1 U18929 ( .A(n18307), .ZN(n8801) );
  AOI22_X1 U18930 ( .A1(\mem[999][7] ), .A2(n18300), .B1(n26131), .B2(
        data_in[7]), .ZN(n18307) );
  NOR2_X1 U18931 ( .A1(N26), .A2(N27), .ZN(n9544) );
  NOR2_X1 U18932 ( .A1(N21), .A2(N22), .ZN(n18238) );
  NOR2_X1 U18933 ( .A1(n27131), .A2(N27), .ZN(n11866) );
  NOR2_X1 U18934 ( .A1(n8606), .A2(N22), .ZN(n18318) );
  NOR3_X1 U18935 ( .A1(N24), .A2(N25), .A3(N23), .ZN(n9546) );
  NOR3_X1 U18936 ( .A1(N24), .A2(N25), .A3(n8607), .ZN(n9836) );
  NOR3_X1 U18937 ( .A1(N23), .A2(N25), .A3(n8608), .ZN(n10126) );
  NOR3_X1 U18938 ( .A1(n8607), .A2(N25), .A3(n8608), .ZN(n10416) );
  BUF_X1 U18939 ( .A(N25), .Z(n8177) );
  INV_X1 U18940 ( .A(N26), .ZN(n27131) );
  AND2_X1 U18941 ( .A1(N27), .A2(N26), .ZN(n16492) );
  AND2_X1 U18942 ( .A1(N27), .A2(n27131), .ZN(n14179) );
  AND2_X1 U18943 ( .A1(N22), .A2(n8606), .ZN(n18391) );
  AND2_X1 U18944 ( .A1(N22), .A2(N21), .ZN(n18464) );
  AND3_X1 U18945 ( .A1(n8607), .A2(n8608), .A3(N25), .ZN(n10706) );
  AND3_X1 U18946 ( .A1(N23), .A2(n8608), .A3(N25), .ZN(n10996) );
  AND3_X1 U18947 ( .A1(N24), .A2(n8607), .A3(N25), .ZN(n11286) );
  AND3_X1 U18948 ( .A1(N24), .A2(N23), .A3(N25), .ZN(n11576) );
  BUF_X1 U18949 ( .A(N22), .Z(n8195) );
  MUX2_X1 U18950 ( .A(\mem[1022][0] ), .B(\mem[1023][0] ), .S(n8389), .Z(n1)
         );
  MUX2_X1 U18951 ( .A(\mem[1020][0] ), .B(\mem[1021][0] ), .S(n8389), .Z(n2)
         );
  MUX2_X1 U18952 ( .A(n2), .B(n1), .S(n8318), .Z(n3) );
  MUX2_X1 U18953 ( .A(\mem[1018][0] ), .B(\mem[1019][0] ), .S(n8389), .Z(n4)
         );
  MUX2_X1 U18954 ( .A(\mem[1016][0] ), .B(\mem[1017][0] ), .S(n8389), .Z(n5)
         );
  MUX2_X1 U18955 ( .A(n5), .B(n4), .S(n8266), .Z(n6) );
  MUX2_X1 U18956 ( .A(n6), .B(n3), .S(n8226), .Z(n7) );
  MUX2_X1 U18957 ( .A(\mem[1014][0] ), .B(\mem[1015][0] ), .S(n8390), .Z(n8)
         );
  MUX2_X1 U18958 ( .A(\mem[1012][0] ), .B(\mem[1013][0] ), .S(n8390), .Z(n9)
         );
  MUX2_X1 U18959 ( .A(n9), .B(n8), .S(n8267), .Z(n10) );
  MUX2_X1 U18960 ( .A(\mem[1010][0] ), .B(\mem[1011][0] ), .S(n8390), .Z(n11)
         );
  MUX2_X1 U18961 ( .A(\mem[1008][0] ), .B(\mem[1009][0] ), .S(n8390), .Z(n12)
         );
  MUX2_X1 U18962 ( .A(n12), .B(n11), .S(n8269), .Z(n13) );
  MUX2_X1 U18963 ( .A(n13), .B(n10), .S(n8226), .Z(n14) );
  MUX2_X1 U18964 ( .A(n14), .B(n7), .S(n8214), .Z(n15) );
  MUX2_X1 U18965 ( .A(\mem[1006][0] ), .B(\mem[1007][0] ), .S(n8390), .Z(n16)
         );
  MUX2_X1 U18966 ( .A(\mem[1004][0] ), .B(\mem[1005][0] ), .S(n8390), .Z(n17)
         );
  MUX2_X1 U18967 ( .A(n17), .B(n16), .S(n8270), .Z(n18) );
  MUX2_X1 U18968 ( .A(\mem[1002][0] ), .B(\mem[1003][0] ), .S(n8390), .Z(n19)
         );
  MUX2_X1 U18969 ( .A(\mem[1000][0] ), .B(\mem[1001][0] ), .S(n8390), .Z(n20)
         );
  MUX2_X1 U18970 ( .A(n20), .B(n19), .S(n8304), .Z(n21) );
  MUX2_X1 U18971 ( .A(n21), .B(n18), .S(n8226), .Z(n22) );
  MUX2_X1 U18972 ( .A(\mem[998][0] ), .B(\mem[999][0] ), .S(n8390), .Z(n23) );
  MUX2_X1 U18973 ( .A(\mem[996][0] ), .B(\mem[997][0] ), .S(n8390), .Z(n24) );
  MUX2_X1 U18974 ( .A(n24), .B(n23), .S(n8311), .Z(n25) );
  MUX2_X1 U18975 ( .A(\mem[994][0] ), .B(\mem[995][0] ), .S(n8390), .Z(n26) );
  MUX2_X1 U18976 ( .A(\mem[992][0] ), .B(\mem[993][0] ), .S(n8390), .Z(n27) );
  MUX2_X1 U18977 ( .A(n27), .B(n26), .S(n8297), .Z(n28) );
  MUX2_X1 U18978 ( .A(n28), .B(n25), .S(n8226), .Z(n29) );
  MUX2_X1 U18979 ( .A(n29), .B(n22), .S(n8202), .Z(n30) );
  MUX2_X1 U18980 ( .A(n30), .B(n15), .S(N22), .Z(n31) );
  MUX2_X1 U18981 ( .A(\mem[990][0] ), .B(\mem[991][0] ), .S(n8391), .Z(n32) );
  MUX2_X1 U18982 ( .A(\mem[988][0] ), .B(\mem[989][0] ), .S(n8391), .Z(n33) );
  MUX2_X1 U18983 ( .A(n33), .B(n32), .S(n8314), .Z(n34) );
  MUX2_X1 U18984 ( .A(\mem[986][0] ), .B(\mem[987][0] ), .S(n8391), .Z(n35) );
  MUX2_X1 U18985 ( .A(\mem[984][0] ), .B(\mem[985][0] ), .S(n8391), .Z(n36) );
  MUX2_X1 U18986 ( .A(n36), .B(n35), .S(n8315), .Z(n37) );
  MUX2_X1 U18987 ( .A(n37), .B(n34), .S(n8227), .Z(n38) );
  MUX2_X1 U18988 ( .A(\mem[982][0] ), .B(\mem[983][0] ), .S(n8391), .Z(n39) );
  MUX2_X1 U18989 ( .A(\mem[980][0] ), .B(\mem[981][0] ), .S(n8391), .Z(n40) );
  MUX2_X1 U18990 ( .A(n40), .B(n39), .S(n8316), .Z(n41) );
  MUX2_X1 U18991 ( .A(\mem[978][0] ), .B(\mem[979][0] ), .S(n8391), .Z(n42) );
  MUX2_X1 U18992 ( .A(\mem[976][0] ), .B(\mem[977][0] ), .S(n8391), .Z(n43) );
  MUX2_X1 U18993 ( .A(n43), .B(n42), .S(n8311), .Z(n44) );
  MUX2_X1 U18994 ( .A(n44), .B(n41), .S(n8227), .Z(n45) );
  MUX2_X1 U18995 ( .A(n45), .B(n38), .S(n8203), .Z(n46) );
  MUX2_X1 U18996 ( .A(\mem[974][0] ), .B(\mem[975][0] ), .S(n8391), .Z(n47) );
  MUX2_X1 U18997 ( .A(\mem[972][0] ), .B(\mem[973][0] ), .S(n8391), .Z(n48) );
  MUX2_X1 U18998 ( .A(n48), .B(n47), .S(n8312), .Z(n49) );
  MUX2_X1 U18999 ( .A(\mem[970][0] ), .B(\mem[971][0] ), .S(n8391), .Z(n50) );
  MUX2_X1 U19000 ( .A(\mem[968][0] ), .B(\mem[969][0] ), .S(n8391), .Z(n51) );
  MUX2_X1 U19001 ( .A(n51), .B(n50), .S(n8313), .Z(n52) );
  MUX2_X1 U19002 ( .A(n52), .B(n49), .S(n8227), .Z(n53) );
  MUX2_X1 U19003 ( .A(\mem[966][0] ), .B(\mem[967][0] ), .S(n8392), .Z(n54) );
  MUX2_X1 U19004 ( .A(\mem[964][0] ), .B(\mem[965][0] ), .S(n8392), .Z(n55) );
  MUX2_X1 U19005 ( .A(n55), .B(n54), .S(n8320), .Z(n56) );
  MUX2_X1 U19006 ( .A(\mem[962][0] ), .B(\mem[963][0] ), .S(n8392), .Z(n57) );
  MUX2_X1 U19007 ( .A(\mem[960][0] ), .B(\mem[961][0] ), .S(n8392), .Z(n58) );
  MUX2_X1 U19008 ( .A(n58), .B(n57), .S(n8321), .Z(n59) );
  MUX2_X1 U19009 ( .A(n59), .B(n56), .S(n8227), .Z(n60) );
  MUX2_X1 U19010 ( .A(n60), .B(n53), .S(n8204), .Z(n61) );
  MUX2_X1 U19011 ( .A(n61), .B(n46), .S(n8195), .Z(n62) );
  MUX2_X1 U19012 ( .A(n62), .B(n31), .S(n8184), .Z(n63) );
  MUX2_X1 U19013 ( .A(\mem[958][0] ), .B(\mem[959][0] ), .S(n8392), .Z(n64) );
  MUX2_X1 U19014 ( .A(\mem[956][0] ), .B(\mem[957][0] ), .S(n8392), .Z(n65) );
  MUX2_X1 U19015 ( .A(n65), .B(n64), .S(n8322), .Z(n66) );
  MUX2_X1 U19016 ( .A(\mem[954][0] ), .B(\mem[955][0] ), .S(n8392), .Z(n67) );
  MUX2_X1 U19017 ( .A(\mem[952][0] ), .B(\mem[953][0] ), .S(n8392), .Z(n68) );
  MUX2_X1 U19018 ( .A(n68), .B(n67), .S(n8317), .Z(n69) );
  MUX2_X1 U19019 ( .A(n69), .B(n66), .S(n8227), .Z(n70) );
  MUX2_X1 U19020 ( .A(\mem[950][0] ), .B(\mem[951][0] ), .S(n8392), .Z(n71) );
  MUX2_X1 U19021 ( .A(\mem[948][0] ), .B(\mem[949][0] ), .S(n8392), .Z(n72) );
  MUX2_X1 U19022 ( .A(n72), .B(n71), .S(n8318), .Z(n73) );
  MUX2_X1 U19023 ( .A(\mem[946][0] ), .B(\mem[947][0] ), .S(n8392), .Z(n74) );
  MUX2_X1 U19024 ( .A(\mem[944][0] ), .B(\mem[945][0] ), .S(n8392), .Z(n75) );
  MUX2_X1 U19025 ( .A(n75), .B(n74), .S(n8319), .Z(n76) );
  MUX2_X1 U19026 ( .A(n76), .B(n73), .S(n8227), .Z(n77) );
  MUX2_X1 U19027 ( .A(n77), .B(n70), .S(n8205), .Z(n78) );
  MUX2_X1 U19028 ( .A(\mem[942][0] ), .B(\mem[943][0] ), .S(n8393), .Z(n79) );
  MUX2_X1 U19029 ( .A(\mem[940][0] ), .B(\mem[941][0] ), .S(n8393), .Z(n80) );
  MUX2_X1 U19030 ( .A(n80), .B(n79), .S(n8296), .Z(n81) );
  MUX2_X1 U19031 ( .A(\mem[938][0] ), .B(\mem[939][0] ), .S(n8393), .Z(n82) );
  MUX2_X1 U19032 ( .A(\mem[936][0] ), .B(\mem[937][0] ), .S(n8393), .Z(n83) );
  MUX2_X1 U19033 ( .A(n83), .B(n82), .S(n8297), .Z(n84) );
  MUX2_X1 U19034 ( .A(n84), .B(n81), .S(n8227), .Z(n85) );
  MUX2_X1 U19035 ( .A(\mem[934][0] ), .B(\mem[935][0] ), .S(n8393), .Z(n86) );
  MUX2_X1 U19036 ( .A(\mem[932][0] ), .B(\mem[933][0] ), .S(n8393), .Z(n87) );
  MUX2_X1 U19037 ( .A(n87), .B(n86), .S(n8298), .Z(n88) );
  MUX2_X1 U19038 ( .A(\mem[930][0] ), .B(\mem[931][0] ), .S(n8393), .Z(n89) );
  MUX2_X1 U19039 ( .A(\mem[928][0] ), .B(\mem[929][0] ), .S(n8393), .Z(n90) );
  MUX2_X1 U19040 ( .A(n90), .B(n89), .S(n8293), .Z(n91) );
  MUX2_X1 U19041 ( .A(n91), .B(n88), .S(n8227), .Z(n92) );
  MUX2_X1 U19042 ( .A(n92), .B(n85), .S(n8217), .Z(n93) );
  MUX2_X1 U19043 ( .A(n93), .B(n78), .S(n8189), .Z(n94) );
  MUX2_X1 U19044 ( .A(\mem[926][0] ), .B(\mem[927][0] ), .S(n8393), .Z(n95) );
  MUX2_X1 U19045 ( .A(\mem[924][0] ), .B(\mem[925][0] ), .S(n8393), .Z(n96) );
  MUX2_X1 U19046 ( .A(n96), .B(n95), .S(n8294), .Z(n97) );
  MUX2_X1 U19047 ( .A(\mem[922][0] ), .B(\mem[923][0] ), .S(n8393), .Z(n98) );
  MUX2_X1 U19048 ( .A(\mem[920][0] ), .B(\mem[921][0] ), .S(n8393), .Z(n99) );
  MUX2_X1 U19049 ( .A(n99), .B(n98), .S(n8295), .Z(n100) );
  MUX2_X1 U19050 ( .A(n100), .B(n97), .S(n8227), .Z(n101) );
  MUX2_X1 U19051 ( .A(\mem[918][0] ), .B(\mem[919][0] ), .S(n8394), .Z(n102)
         );
  MUX2_X1 U19052 ( .A(\mem[916][0] ), .B(\mem[917][0] ), .S(n8394), .Z(n103)
         );
  MUX2_X1 U19053 ( .A(n103), .B(n102), .S(n8302), .Z(n104) );
  MUX2_X1 U19054 ( .A(\mem[914][0] ), .B(\mem[915][0] ), .S(n8394), .Z(n105)
         );
  MUX2_X1 U19055 ( .A(\mem[912][0] ), .B(\mem[913][0] ), .S(n8394), .Z(n106)
         );
  MUX2_X1 U19056 ( .A(n106), .B(n105), .S(n8303), .Z(n107) );
  MUX2_X1 U19057 ( .A(n107), .B(n104), .S(n8227), .Z(n108) );
  MUX2_X1 U19058 ( .A(n108), .B(n101), .S(n8212), .Z(n109) );
  MUX2_X1 U19059 ( .A(\mem[910][0] ), .B(\mem[911][0] ), .S(n8394), .Z(n110)
         );
  MUX2_X1 U19060 ( .A(\mem[908][0] ), .B(\mem[909][0] ), .S(n8394), .Z(n111)
         );
  MUX2_X1 U19061 ( .A(n111), .B(n110), .S(n8304), .Z(n112) );
  MUX2_X1 U19062 ( .A(\mem[906][0] ), .B(\mem[907][0] ), .S(n8394), .Z(n113)
         );
  MUX2_X1 U19063 ( .A(\mem[904][0] ), .B(\mem[905][0] ), .S(n8394), .Z(n114)
         );
  MUX2_X1 U19064 ( .A(n114), .B(n113), .S(n8299), .Z(n115) );
  MUX2_X1 U19065 ( .A(n115), .B(n112), .S(n8227), .Z(n116) );
  MUX2_X1 U19066 ( .A(\mem[902][0] ), .B(\mem[903][0] ), .S(n8394), .Z(n117)
         );
  MUX2_X1 U19067 ( .A(\mem[900][0] ), .B(\mem[901][0] ), .S(n8394), .Z(n118)
         );
  MUX2_X1 U19068 ( .A(n118), .B(n117), .S(n8300), .Z(n119) );
  MUX2_X1 U19069 ( .A(\mem[898][0] ), .B(\mem[899][0] ), .S(n8394), .Z(n120)
         );
  MUX2_X1 U19070 ( .A(\mem[896][0] ), .B(\mem[897][0] ), .S(n8394), .Z(n121)
         );
  MUX2_X1 U19071 ( .A(n121), .B(n120), .S(n8301), .Z(n122) );
  MUX2_X1 U19072 ( .A(n122), .B(n119), .S(n8227), .Z(n123) );
  MUX2_X1 U19073 ( .A(n123), .B(n116), .S(n8213), .Z(n124) );
  MUX2_X1 U19074 ( .A(n124), .B(n109), .S(n8194), .Z(n125) );
  MUX2_X1 U19075 ( .A(n125), .B(n94), .S(N23), .Z(n126) );
  MUX2_X1 U19076 ( .A(n126), .B(n63), .S(n8178), .Z(n127) );
  MUX2_X1 U19077 ( .A(\mem[894][0] ), .B(\mem[895][0] ), .S(n8395), .Z(n128)
         );
  MUX2_X1 U19078 ( .A(\mem[892][0] ), .B(\mem[893][0] ), .S(n8395), .Z(n129)
         );
  MUX2_X1 U19079 ( .A(n129), .B(n128), .S(n8314), .Z(n130) );
  MUX2_X1 U19080 ( .A(\mem[890][0] ), .B(\mem[891][0] ), .S(n8395), .Z(n131)
         );
  MUX2_X1 U19081 ( .A(\mem[888][0] ), .B(\mem[889][0] ), .S(n8395), .Z(n132)
         );
  MUX2_X1 U19082 ( .A(n132), .B(n131), .S(n8350), .Z(n133) );
  MUX2_X1 U19083 ( .A(n133), .B(n130), .S(n8228), .Z(n134) );
  MUX2_X1 U19084 ( .A(\mem[886][0] ), .B(\mem[887][0] ), .S(n8395), .Z(n135)
         );
  MUX2_X1 U19085 ( .A(\mem[884][0] ), .B(\mem[885][0] ), .S(n8395), .Z(n136)
         );
  MUX2_X1 U19086 ( .A(n136), .B(n135), .S(n8323), .Z(n137) );
  MUX2_X1 U19087 ( .A(\mem[882][0] ), .B(\mem[883][0] ), .S(n8395), .Z(n138)
         );
  MUX2_X1 U19088 ( .A(\mem[880][0] ), .B(\mem[881][0] ), .S(n8395), .Z(n139)
         );
  MUX2_X1 U19089 ( .A(n139), .B(n138), .S(n8290), .Z(n140) );
  MUX2_X1 U19090 ( .A(n140), .B(n137), .S(n8228), .Z(n141) );
  MUX2_X1 U19091 ( .A(n141), .B(n134), .S(n8214), .Z(n142) );
  MUX2_X1 U19092 ( .A(\mem[878][0] ), .B(\mem[879][0] ), .S(n8395), .Z(n143)
         );
  MUX2_X1 U19093 ( .A(\mem[876][0] ), .B(\mem[877][0] ), .S(n8395), .Z(n144)
         );
  MUX2_X1 U19094 ( .A(n144), .B(n143), .S(n8284), .Z(n145) );
  MUX2_X1 U19095 ( .A(\mem[874][0] ), .B(\mem[875][0] ), .S(n8395), .Z(n146)
         );
  MUX2_X1 U19096 ( .A(\mem[872][0] ), .B(\mem[873][0] ), .S(n8395), .Z(n147)
         );
  MUX2_X1 U19097 ( .A(n147), .B(n146), .S(n8329), .Z(n148) );
  MUX2_X1 U19098 ( .A(n148), .B(n145), .S(n8228), .Z(n149) );
  MUX2_X1 U19099 ( .A(\mem[870][0] ), .B(\mem[871][0] ), .S(n8396), .Z(n150)
         );
  MUX2_X1 U19100 ( .A(\mem[868][0] ), .B(\mem[869][0] ), .S(n8396), .Z(n151)
         );
  MUX2_X1 U19101 ( .A(n151), .B(n150), .S(n8296), .Z(n152) );
  MUX2_X1 U19102 ( .A(\mem[866][0] ), .B(\mem[867][0] ), .S(n8396), .Z(n153)
         );
  MUX2_X1 U19103 ( .A(\mem[864][0] ), .B(\mem[865][0] ), .S(n8396), .Z(n154)
         );
  MUX2_X1 U19104 ( .A(n154), .B(n153), .S(n8280), .Z(n155) );
  MUX2_X1 U19105 ( .A(n155), .B(n152), .S(n8228), .Z(n156) );
  MUX2_X1 U19106 ( .A(n156), .B(n149), .S(n8215), .Z(n157) );
  MUX2_X1 U19107 ( .A(n157), .B(n142), .S(n8194), .Z(n158) );
  MUX2_X1 U19108 ( .A(\mem[862][0] ), .B(\mem[863][0] ), .S(n8396), .Z(n159)
         );
  MUX2_X1 U19109 ( .A(\mem[860][0] ), .B(\mem[861][0] ), .S(n8396), .Z(n160)
         );
  MUX2_X1 U19110 ( .A(n160), .B(n159), .S(n8284), .Z(n161) );
  MUX2_X1 U19111 ( .A(\mem[858][0] ), .B(\mem[859][0] ), .S(n8396), .Z(n162)
         );
  MUX2_X1 U19112 ( .A(\mem[856][0] ), .B(\mem[857][0] ), .S(n8396), .Z(n163)
         );
  MUX2_X1 U19113 ( .A(n163), .B(n162), .S(n8285), .Z(n164) );
  MUX2_X1 U19114 ( .A(n164), .B(n161), .S(n8228), .Z(n165) );
  MUX2_X1 U19115 ( .A(\mem[854][0] ), .B(\mem[855][0] ), .S(n8396), .Z(n166)
         );
  MUX2_X1 U19116 ( .A(\mem[852][0] ), .B(\mem[853][0] ), .S(n8396), .Z(n167)
         );
  MUX2_X1 U19117 ( .A(n167), .B(n166), .S(n8286), .Z(n168) );
  MUX2_X1 U19118 ( .A(\mem[850][0] ), .B(\mem[851][0] ), .S(n8396), .Z(n169)
         );
  MUX2_X1 U19119 ( .A(\mem[848][0] ), .B(\mem[849][0] ), .S(n8396), .Z(n170)
         );
  MUX2_X1 U19120 ( .A(n170), .B(n169), .S(n8290), .Z(n171) );
  MUX2_X1 U19121 ( .A(n171), .B(n168), .S(n8228), .Z(n172) );
  MUX2_X1 U19122 ( .A(n172), .B(n165), .S(n8211), .Z(n173) );
  MUX2_X1 U19123 ( .A(\mem[846][0] ), .B(\mem[847][0] ), .S(n8397), .Z(n174)
         );
  MUX2_X1 U19124 ( .A(\mem[844][0] ), .B(\mem[845][0] ), .S(n8397), .Z(n175)
         );
  MUX2_X1 U19125 ( .A(n175), .B(n174), .S(n8333), .Z(n176) );
  MUX2_X1 U19126 ( .A(\mem[842][0] ), .B(\mem[843][0] ), .S(n8397), .Z(n177)
         );
  MUX2_X1 U19127 ( .A(\mem[840][0] ), .B(\mem[841][0] ), .S(n8397), .Z(n178)
         );
  MUX2_X1 U19128 ( .A(n178), .B(n177), .S(n8334), .Z(n179) );
  MUX2_X1 U19129 ( .A(n179), .B(n176), .S(n8228), .Z(n180) );
  MUX2_X1 U19130 ( .A(\mem[838][0] ), .B(\mem[839][0] ), .S(n8397), .Z(n181)
         );
  MUX2_X1 U19131 ( .A(\mem[836][0] ), .B(\mem[837][0] ), .S(n8397), .Z(n182)
         );
  MUX2_X1 U19132 ( .A(n182), .B(n181), .S(n8329), .Z(n183) );
  MUX2_X1 U19133 ( .A(\mem[834][0] ), .B(\mem[835][0] ), .S(n8397), .Z(n184)
         );
  MUX2_X1 U19134 ( .A(\mem[832][0] ), .B(\mem[833][0] ), .S(n8397), .Z(n185)
         );
  MUX2_X1 U19135 ( .A(n185), .B(n184), .S(n8330), .Z(n186) );
  MUX2_X1 U19136 ( .A(n186), .B(n183), .S(n8228), .Z(n187) );
  MUX2_X1 U19137 ( .A(n187), .B(n180), .S(n8216), .Z(n188) );
  MUX2_X1 U19138 ( .A(n188), .B(n173), .S(n8186), .Z(n189) );
  MUX2_X1 U19139 ( .A(n189), .B(n158), .S(n8185), .Z(n190) );
  MUX2_X1 U19140 ( .A(\mem[830][0] ), .B(\mem[831][0] ), .S(n8397), .Z(n191)
         );
  MUX2_X1 U19141 ( .A(\mem[828][0] ), .B(\mem[829][0] ), .S(n8397), .Z(n192)
         );
  MUX2_X1 U19142 ( .A(n192), .B(n191), .S(n8331), .Z(n193) );
  MUX2_X1 U19143 ( .A(\mem[826][0] ), .B(\mem[827][0] ), .S(n8397), .Z(n194)
         );
  MUX2_X1 U19144 ( .A(\mem[824][0] ), .B(\mem[825][0] ), .S(n8397), .Z(n195)
         );
  MUX2_X1 U19145 ( .A(n195), .B(n194), .S(n8338), .Z(n196) );
  MUX2_X1 U19146 ( .A(n196), .B(n193), .S(n8228), .Z(n197) );
  MUX2_X1 U19147 ( .A(\mem[822][0] ), .B(\mem[823][0] ), .S(n8398), .Z(n198)
         );
  MUX2_X1 U19148 ( .A(\mem[820][0] ), .B(\mem[821][0] ), .S(n8398), .Z(n199)
         );
  MUX2_X1 U19149 ( .A(n199), .B(n198), .S(n8339), .Z(n200) );
  MUX2_X1 U19150 ( .A(\mem[818][0] ), .B(\mem[819][0] ), .S(n8398), .Z(n201)
         );
  MUX2_X1 U19151 ( .A(\mem[816][0] ), .B(\mem[817][0] ), .S(n8398), .Z(n202)
         );
  MUX2_X1 U19152 ( .A(n202), .B(n201), .S(n8340), .Z(n203) );
  MUX2_X1 U19153 ( .A(n203), .B(n200), .S(n8228), .Z(n204) );
  MUX2_X1 U19154 ( .A(n204), .B(n197), .S(n8217), .Z(n205) );
  MUX2_X1 U19155 ( .A(\mem[814][0] ), .B(\mem[815][0] ), .S(n8398), .Z(n206)
         );
  MUX2_X1 U19156 ( .A(\mem[812][0] ), .B(\mem[813][0] ), .S(n8398), .Z(n207)
         );
  MUX2_X1 U19157 ( .A(n207), .B(n206), .S(n8335), .Z(n208) );
  MUX2_X1 U19158 ( .A(\mem[810][0] ), .B(\mem[811][0] ), .S(n8398), .Z(n209)
         );
  MUX2_X1 U19159 ( .A(\mem[808][0] ), .B(\mem[809][0] ), .S(n8398), .Z(n210)
         );
  MUX2_X1 U19160 ( .A(n210), .B(n209), .S(n8337), .Z(n211) );
  MUX2_X1 U19161 ( .A(n211), .B(n208), .S(n8228), .Z(n212) );
  MUX2_X1 U19162 ( .A(\mem[806][0] ), .B(\mem[807][0] ), .S(n8398), .Z(n213)
         );
  MUX2_X1 U19163 ( .A(\mem[804][0] ), .B(\mem[805][0] ), .S(n8398), .Z(n214)
         );
  MUX2_X1 U19164 ( .A(n214), .B(n213), .S(N19), .Z(n215) );
  MUX2_X1 U19165 ( .A(\mem[802][0] ), .B(\mem[803][0] ), .S(n8398), .Z(n216)
         );
  MUX2_X1 U19166 ( .A(\mem[800][0] ), .B(\mem[801][0] ), .S(n8398), .Z(n217)
         );
  MUX2_X1 U19167 ( .A(n217), .B(n216), .S(n8356), .Z(n218) );
  MUX2_X1 U19168 ( .A(n218), .B(n215), .S(n8228), .Z(n219) );
  MUX2_X1 U19169 ( .A(n219), .B(n212), .S(n8218), .Z(n220) );
  MUX2_X1 U19170 ( .A(n220), .B(n205), .S(n8187), .Z(n221) );
  MUX2_X1 U19171 ( .A(\mem[798][0] ), .B(\mem[799][0] ), .S(n8399), .Z(n222)
         );
  MUX2_X1 U19172 ( .A(\mem[796][0] ), .B(\mem[797][0] ), .S(n8399), .Z(n223)
         );
  MUX2_X1 U19173 ( .A(n223), .B(n222), .S(n8343), .Z(n224) );
  MUX2_X1 U19174 ( .A(\mem[794][0] ), .B(\mem[795][0] ), .S(n8399), .Z(n225)
         );
  MUX2_X1 U19175 ( .A(\mem[792][0] ), .B(\mem[793][0] ), .S(n8399), .Z(n226)
         );
  MUX2_X1 U19176 ( .A(n226), .B(n225), .S(n8350), .Z(n227) );
  MUX2_X1 U19177 ( .A(n227), .B(n224), .S(n8229), .Z(n228) );
  MUX2_X1 U19178 ( .A(\mem[790][0] ), .B(\mem[791][0] ), .S(n8399), .Z(n229)
         );
  MUX2_X1 U19179 ( .A(\mem[788][0] ), .B(\mem[789][0] ), .S(n8399), .Z(n230)
         );
  MUX2_X1 U19180 ( .A(n230), .B(n229), .S(n8351), .Z(n231) );
  MUX2_X1 U19181 ( .A(\mem[786][0] ), .B(\mem[787][0] ), .S(n8399), .Z(n232)
         );
  MUX2_X1 U19182 ( .A(\mem[784][0] ), .B(\mem[785][0] ), .S(n8399), .Z(n233)
         );
  MUX2_X1 U19183 ( .A(n233), .B(n232), .S(n8352), .Z(n234) );
  MUX2_X1 U19184 ( .A(n234), .B(n231), .S(n8229), .Z(n235) );
  MUX2_X1 U19185 ( .A(n235), .B(n228), .S(n8207), .Z(n236) );
  MUX2_X1 U19186 ( .A(\mem[782][0] ), .B(\mem[783][0] ), .S(n8399), .Z(n237)
         );
  MUX2_X1 U19187 ( .A(\mem[780][0] ), .B(\mem[781][0] ), .S(n8399), .Z(n238)
         );
  MUX2_X1 U19188 ( .A(n238), .B(n237), .S(n8347), .Z(n239) );
  MUX2_X1 U19189 ( .A(\mem[778][0] ), .B(\mem[779][0] ), .S(n8399), .Z(n240)
         );
  MUX2_X1 U19190 ( .A(\mem[776][0] ), .B(\mem[777][0] ), .S(n8399), .Z(n241)
         );
  MUX2_X1 U19191 ( .A(n241), .B(n240), .S(n8348), .Z(n242) );
  MUX2_X1 U19192 ( .A(n242), .B(n239), .S(n8229), .Z(n243) );
  MUX2_X1 U19193 ( .A(\mem[774][0] ), .B(\mem[775][0] ), .S(n8400), .Z(n244)
         );
  MUX2_X1 U19194 ( .A(\mem[772][0] ), .B(\mem[773][0] ), .S(n8400), .Z(n245)
         );
  MUX2_X1 U19195 ( .A(n245), .B(n244), .S(n8349), .Z(n246) );
  MUX2_X1 U19196 ( .A(\mem[770][0] ), .B(\mem[771][0] ), .S(n8400), .Z(n247)
         );
  MUX2_X1 U19197 ( .A(\mem[768][0] ), .B(\mem[769][0] ), .S(n8400), .Z(n248)
         );
  MUX2_X1 U19198 ( .A(n248), .B(n247), .S(n8353), .Z(n249) );
  MUX2_X1 U19199 ( .A(n249), .B(n246), .S(n8229), .Z(n250) );
  MUX2_X1 U19200 ( .A(n250), .B(n243), .S(n8208), .Z(n251) );
  MUX2_X1 U19201 ( .A(n251), .B(n236), .S(n8188), .Z(n252) );
  MUX2_X1 U19202 ( .A(n252), .B(n221), .S(n8181), .Z(n253) );
  MUX2_X1 U19203 ( .A(n253), .B(n190), .S(n8178), .Z(n254) );
  MUX2_X1 U19204 ( .A(n254), .B(n127), .S(N25), .Z(n255) );
  MUX2_X1 U19205 ( .A(\mem[766][0] ), .B(\mem[767][0] ), .S(n8400), .Z(n256)
         );
  MUX2_X1 U19206 ( .A(\mem[764][0] ), .B(\mem[765][0] ), .S(n8400), .Z(n257)
         );
  MUX2_X1 U19207 ( .A(n257), .B(n256), .S(n8354), .Z(n258) );
  MUX2_X1 U19208 ( .A(\mem[762][0] ), .B(\mem[763][0] ), .S(n8400), .Z(n259)
         );
  MUX2_X1 U19209 ( .A(\mem[760][0] ), .B(\mem[761][0] ), .S(n8400), .Z(n260)
         );
  MUX2_X1 U19210 ( .A(n260), .B(n259), .S(n8355), .Z(n261) );
  MUX2_X1 U19211 ( .A(n261), .B(n258), .S(n8229), .Z(n262) );
  MUX2_X1 U19212 ( .A(\mem[758][0] ), .B(\mem[759][0] ), .S(n8400), .Z(n263)
         );
  MUX2_X1 U19213 ( .A(\mem[756][0] ), .B(\mem[757][0] ), .S(n8400), .Z(n264)
         );
  MUX2_X1 U19214 ( .A(n264), .B(n263), .S(n8326), .Z(n265) );
  MUX2_X1 U19215 ( .A(\mem[754][0] ), .B(\mem[755][0] ), .S(n8400), .Z(n266)
         );
  MUX2_X1 U19216 ( .A(\mem[752][0] ), .B(\mem[753][0] ), .S(n8400), .Z(n267)
         );
  MUX2_X1 U19217 ( .A(n267), .B(n266), .S(n8327), .Z(n268) );
  MUX2_X1 U19218 ( .A(n268), .B(n265), .S(n8229), .Z(n269) );
  MUX2_X1 U19219 ( .A(n269), .B(n262), .S(n8209), .Z(n270) );
  MUX2_X1 U19220 ( .A(\mem[750][0] ), .B(\mem[751][0] ), .S(n8401), .Z(n271)
         );
  MUX2_X1 U19221 ( .A(\mem[748][0] ), .B(\mem[749][0] ), .S(n8401), .Z(n272)
         );
  MUX2_X1 U19222 ( .A(n272), .B(n271), .S(n8291), .Z(n273) );
  MUX2_X1 U19223 ( .A(\mem[746][0] ), .B(\mem[747][0] ), .S(n8401), .Z(n274)
         );
  MUX2_X1 U19224 ( .A(\mem[744][0] ), .B(\mem[745][0] ), .S(n8401), .Z(n275)
         );
  MUX2_X1 U19225 ( .A(n275), .B(n274), .S(n8292), .Z(n276) );
  MUX2_X1 U19226 ( .A(n276), .B(n273), .S(n8229), .Z(n277) );
  MUX2_X1 U19227 ( .A(\mem[742][0] ), .B(\mem[743][0] ), .S(n8401), .Z(n278)
         );
  MUX2_X1 U19228 ( .A(\mem[740][0] ), .B(\mem[741][0] ), .S(n8401), .Z(n279)
         );
  MUX2_X1 U19229 ( .A(n279), .B(n278), .S(n8287), .Z(n280) );
  MUX2_X1 U19230 ( .A(\mem[738][0] ), .B(\mem[739][0] ), .S(n8401), .Z(n281)
         );
  MUX2_X1 U19231 ( .A(\mem[736][0] ), .B(\mem[737][0] ), .S(n8401), .Z(n282)
         );
  MUX2_X1 U19232 ( .A(n282), .B(n281), .S(n8288), .Z(n283) );
  MUX2_X1 U19233 ( .A(n283), .B(n280), .S(n8229), .Z(n284) );
  MUX2_X1 U19234 ( .A(n284), .B(n277), .S(n8210), .Z(n285) );
  MUX2_X1 U19235 ( .A(n285), .B(n270), .S(n8192), .Z(n286) );
  MUX2_X1 U19236 ( .A(\mem[734][0] ), .B(\mem[735][0] ), .S(n8401), .Z(n287)
         );
  MUX2_X1 U19237 ( .A(\mem[732][0] ), .B(\mem[733][0] ), .S(n8401), .Z(n288)
         );
  MUX2_X1 U19238 ( .A(n288), .B(n287), .S(n8289), .Z(n289) );
  MUX2_X1 U19239 ( .A(\mem[730][0] ), .B(\mem[731][0] ), .S(n8401), .Z(n290)
         );
  MUX2_X1 U19240 ( .A(\mem[728][0] ), .B(\mem[729][0] ), .S(n8401), .Z(n291)
         );
  MUX2_X1 U19241 ( .A(n291), .B(n290), .S(n8296), .Z(n292) );
  MUX2_X1 U19242 ( .A(n292), .B(n289), .S(n8229), .Z(n293) );
  MUX2_X1 U19243 ( .A(\mem[726][0] ), .B(\mem[727][0] ), .S(n8402), .Z(n294)
         );
  MUX2_X1 U19244 ( .A(\mem[724][0] ), .B(\mem[725][0] ), .S(n8402), .Z(n295)
         );
  MUX2_X1 U19245 ( .A(n295), .B(n294), .S(n8297), .Z(n296) );
  MUX2_X1 U19246 ( .A(\mem[722][0] ), .B(\mem[723][0] ), .S(n8402), .Z(n297)
         );
  MUX2_X1 U19247 ( .A(\mem[720][0] ), .B(\mem[721][0] ), .S(n8402), .Z(n298)
         );
  MUX2_X1 U19248 ( .A(n298), .B(n297), .S(n8298), .Z(n299) );
  MUX2_X1 U19249 ( .A(n299), .B(n296), .S(n8229), .Z(n300) );
  MUX2_X1 U19250 ( .A(n300), .B(n293), .S(n8206), .Z(n301) );
  MUX2_X1 U19251 ( .A(\mem[718][0] ), .B(\mem[719][0] ), .S(n8402), .Z(n302)
         );
  MUX2_X1 U19252 ( .A(\mem[716][0] ), .B(\mem[717][0] ), .S(n8402), .Z(n303)
         );
  MUX2_X1 U19253 ( .A(n303), .B(n302), .S(n8293), .Z(n304) );
  MUX2_X1 U19254 ( .A(\mem[714][0] ), .B(\mem[715][0] ), .S(n8402), .Z(n305)
         );
  MUX2_X1 U19255 ( .A(\mem[712][0] ), .B(\mem[713][0] ), .S(n8402), .Z(n306)
         );
  MUX2_X1 U19256 ( .A(n306), .B(n305), .S(n8294), .Z(n307) );
  MUX2_X1 U19257 ( .A(n307), .B(n304), .S(n8229), .Z(n308) );
  MUX2_X1 U19258 ( .A(\mem[710][0] ), .B(\mem[711][0] ), .S(n8402), .Z(n309)
         );
  MUX2_X1 U19259 ( .A(\mem[708][0] ), .B(\mem[709][0] ), .S(n8402), .Z(n310)
         );
  MUX2_X1 U19260 ( .A(n310), .B(n309), .S(n8295), .Z(n311) );
  MUX2_X1 U19261 ( .A(\mem[706][0] ), .B(\mem[707][0] ), .S(n8402), .Z(n312)
         );
  MUX2_X1 U19262 ( .A(\mem[704][0] ), .B(\mem[705][0] ), .S(n8402), .Z(n313)
         );
  MUX2_X1 U19263 ( .A(n313), .B(n312), .S(n8302), .Z(n314) );
  MUX2_X1 U19264 ( .A(n314), .B(n311), .S(n8229), .Z(n315) );
  MUX2_X1 U19265 ( .A(n315), .B(n308), .S(n8198), .Z(n316) );
  MUX2_X1 U19266 ( .A(n316), .B(n301), .S(n8193), .Z(n317) );
  MUX2_X1 U19267 ( .A(n317), .B(n286), .S(n8182), .Z(n318) );
  MUX2_X1 U19268 ( .A(\mem[702][0] ), .B(\mem[703][0] ), .S(n8403), .Z(n319)
         );
  MUX2_X1 U19269 ( .A(\mem[700][0] ), .B(\mem[701][0] ), .S(n8403), .Z(n320)
         );
  MUX2_X1 U19270 ( .A(n320), .B(n319), .S(n8337), .Z(n321) );
  MUX2_X1 U19271 ( .A(\mem[698][0] ), .B(\mem[699][0] ), .S(n8403), .Z(n322)
         );
  MUX2_X1 U19272 ( .A(\mem[696][0] ), .B(\mem[697][0] ), .S(n8403), .Z(n323)
         );
  MUX2_X1 U19273 ( .A(n323), .B(n322), .S(N19), .Z(n324) );
  MUX2_X1 U19274 ( .A(n324), .B(n321), .S(n8230), .Z(n325) );
  MUX2_X1 U19275 ( .A(\mem[694][0] ), .B(\mem[695][0] ), .S(n8403), .Z(n326)
         );
  MUX2_X1 U19276 ( .A(\mem[692][0] ), .B(\mem[693][0] ), .S(n8403), .Z(n327)
         );
  MUX2_X1 U19277 ( .A(n327), .B(n326), .S(n8356), .Z(n328) );
  MUX2_X1 U19278 ( .A(\mem[690][0] ), .B(\mem[691][0] ), .S(n8403), .Z(n329)
         );
  MUX2_X1 U19279 ( .A(\mem[688][0] ), .B(\mem[689][0] ), .S(n8403), .Z(n330)
         );
  MUX2_X1 U19280 ( .A(n330), .B(n329), .S(n8336), .Z(n331) );
  MUX2_X1 U19281 ( .A(n331), .B(n328), .S(n8230), .Z(n332) );
  MUX2_X1 U19282 ( .A(n332), .B(n325), .S(n8216), .Z(n333) );
  MUX2_X1 U19283 ( .A(\mem[686][0] ), .B(\mem[687][0] ), .S(n8403), .Z(n334)
         );
  MUX2_X1 U19284 ( .A(\mem[684][0] ), .B(\mem[685][0] ), .S(n8403), .Z(n335)
         );
  MUX2_X1 U19285 ( .A(n335), .B(n334), .S(n8344), .Z(n336) );
  MUX2_X1 U19286 ( .A(\mem[682][0] ), .B(\mem[683][0] ), .S(n8403), .Z(n337)
         );
  MUX2_X1 U19287 ( .A(\mem[680][0] ), .B(\mem[681][0] ), .S(n8403), .Z(n338)
         );
  MUX2_X1 U19288 ( .A(n338), .B(n337), .S(n8267), .Z(n339) );
  MUX2_X1 U19289 ( .A(n339), .B(n336), .S(n8230), .Z(n340) );
  MUX2_X1 U19290 ( .A(\mem[678][0] ), .B(\mem[679][0] ), .S(n8404), .Z(n341)
         );
  MUX2_X1 U19291 ( .A(\mem[676][0] ), .B(\mem[677][0] ), .S(n8404), .Z(n342)
         );
  MUX2_X1 U19292 ( .A(n342), .B(n341), .S(n8269), .Z(n343) );
  MUX2_X1 U19293 ( .A(\mem[674][0] ), .B(\mem[675][0] ), .S(n8404), .Z(n344)
         );
  MUX2_X1 U19294 ( .A(\mem[672][0] ), .B(\mem[673][0] ), .S(n8404), .Z(n345)
         );
  MUX2_X1 U19295 ( .A(n345), .B(n344), .S(n8273), .Z(n346) );
  MUX2_X1 U19296 ( .A(n346), .B(n343), .S(n8230), .Z(n347) );
  MUX2_X1 U19297 ( .A(n347), .B(n340), .S(n8212), .Z(n348) );
  MUX2_X1 U19298 ( .A(n348), .B(n333), .S(n8190), .Z(n349) );
  MUX2_X1 U19299 ( .A(\mem[670][0] ), .B(\mem[671][0] ), .S(n8404), .Z(n350)
         );
  MUX2_X1 U19300 ( .A(\mem[668][0] ), .B(\mem[669][0] ), .S(n8404), .Z(n351)
         );
  MUX2_X1 U19301 ( .A(n351), .B(n350), .S(n8337), .Z(n352) );
  MUX2_X1 U19302 ( .A(\mem[666][0] ), .B(\mem[667][0] ), .S(n8404), .Z(n353)
         );
  MUX2_X1 U19303 ( .A(\mem[664][0] ), .B(\mem[665][0] ), .S(n8404), .Z(n354)
         );
  MUX2_X1 U19304 ( .A(n354), .B(n353), .S(n8300), .Z(n355) );
  MUX2_X1 U19305 ( .A(n355), .B(n352), .S(n8230), .Z(n356) );
  MUX2_X1 U19306 ( .A(\mem[662][0] ), .B(\mem[663][0] ), .S(n8404), .Z(n357)
         );
  MUX2_X1 U19307 ( .A(\mem[660][0] ), .B(\mem[661][0] ), .S(n8404), .Z(n358)
         );
  MUX2_X1 U19308 ( .A(n358), .B(n357), .S(n8282), .Z(n359) );
  MUX2_X1 U19309 ( .A(\mem[658][0] ), .B(\mem[659][0] ), .S(n8404), .Z(n360)
         );
  MUX2_X1 U19310 ( .A(\mem[656][0] ), .B(\mem[657][0] ), .S(n8404), .Z(n361)
         );
  MUX2_X1 U19311 ( .A(n361), .B(n360), .S(n8281), .Z(n362) );
  MUX2_X1 U19312 ( .A(n362), .B(n359), .S(n8230), .Z(n363) );
  MUX2_X1 U19313 ( .A(n363), .B(n356), .S(n8213), .Z(n364) );
  MUX2_X1 U19314 ( .A(\mem[654][0] ), .B(\mem[655][0] ), .S(n8405), .Z(n365)
         );
  MUX2_X1 U19315 ( .A(\mem[652][0] ), .B(\mem[653][0] ), .S(n8405), .Z(n366)
         );
  MUX2_X1 U19316 ( .A(n366), .B(n365), .S(n8316), .Z(n367) );
  MUX2_X1 U19317 ( .A(\mem[650][0] ), .B(\mem[651][0] ), .S(n8405), .Z(n368)
         );
  MUX2_X1 U19318 ( .A(\mem[648][0] ), .B(\mem[649][0] ), .S(n8405), .Z(n369)
         );
  MUX2_X1 U19319 ( .A(n369), .B(n368), .S(n8326), .Z(n370) );
  MUX2_X1 U19320 ( .A(n370), .B(n367), .S(n8230), .Z(n371) );
  MUX2_X1 U19321 ( .A(\mem[646][0] ), .B(\mem[647][0] ), .S(n8405), .Z(n372)
         );
  MUX2_X1 U19322 ( .A(\mem[644][0] ), .B(\mem[645][0] ), .S(n8405), .Z(n373)
         );
  MUX2_X1 U19323 ( .A(n373), .B(n372), .S(n8322), .Z(n374) );
  MUX2_X1 U19324 ( .A(\mem[642][0] ), .B(\mem[643][0] ), .S(n8405), .Z(n375)
         );
  MUX2_X1 U19325 ( .A(\mem[640][0] ), .B(\mem[641][0] ), .S(n8405), .Z(n376)
         );
  MUX2_X1 U19326 ( .A(n376), .B(n375), .S(n8327), .Z(n377) );
  MUX2_X1 U19327 ( .A(n377), .B(n374), .S(n8230), .Z(n378) );
  MUX2_X1 U19328 ( .A(n378), .B(n371), .S(n8214), .Z(n379) );
  MUX2_X1 U19329 ( .A(n379), .B(n364), .S(n8193), .Z(n380) );
  MUX2_X1 U19330 ( .A(n380), .B(n349), .S(n8183), .Z(n381) );
  MUX2_X1 U19331 ( .A(n381), .B(n318), .S(n8178), .Z(n382) );
  MUX2_X1 U19332 ( .A(\mem[638][0] ), .B(\mem[639][0] ), .S(n8405), .Z(n383)
         );
  MUX2_X1 U19333 ( .A(\mem[636][0] ), .B(\mem[637][0] ), .S(n8405), .Z(n384)
         );
  MUX2_X1 U19334 ( .A(n384), .B(n383), .S(n8283), .Z(n385) );
  MUX2_X1 U19335 ( .A(\mem[634][0] ), .B(\mem[635][0] ), .S(n8405), .Z(n386)
         );
  MUX2_X1 U19336 ( .A(\mem[632][0] ), .B(\mem[633][0] ), .S(n8405), .Z(n387)
         );
  MUX2_X1 U19337 ( .A(n387), .B(n386), .S(n8307), .Z(n388) );
  MUX2_X1 U19338 ( .A(n388), .B(n385), .S(n8230), .Z(n389) );
  MUX2_X1 U19339 ( .A(\mem[630][0] ), .B(\mem[631][0] ), .S(n8406), .Z(n390)
         );
  MUX2_X1 U19340 ( .A(\mem[628][0] ), .B(\mem[629][0] ), .S(n8406), .Z(n391)
         );
  MUX2_X1 U19341 ( .A(n391), .B(n390), .S(n8343), .Z(n392) );
  MUX2_X1 U19342 ( .A(\mem[626][0] ), .B(\mem[627][0] ), .S(n8406), .Z(n393)
         );
  MUX2_X1 U19343 ( .A(\mem[624][0] ), .B(\mem[625][0] ), .S(n8406), .Z(n394)
         );
  MUX2_X1 U19344 ( .A(n394), .B(n393), .S(n8328), .Z(n395) );
  MUX2_X1 U19345 ( .A(n395), .B(n392), .S(n8230), .Z(n396) );
  MUX2_X1 U19346 ( .A(n396), .B(n389), .S(n8215), .Z(n397) );
  MUX2_X1 U19347 ( .A(\mem[622][0] ), .B(\mem[623][0] ), .S(n8406), .Z(n398)
         );
  MUX2_X1 U19348 ( .A(\mem[620][0] ), .B(\mem[621][0] ), .S(n8406), .Z(n399)
         );
  MUX2_X1 U19349 ( .A(n399), .B(n398), .S(n8283), .Z(n400) );
  MUX2_X1 U19350 ( .A(\mem[618][0] ), .B(\mem[619][0] ), .S(n8406), .Z(n401)
         );
  MUX2_X1 U19351 ( .A(\mem[616][0] ), .B(\mem[617][0] ), .S(n8406), .Z(n402)
         );
  MUX2_X1 U19352 ( .A(n402), .B(n401), .S(n8349), .Z(n403) );
  MUX2_X1 U19353 ( .A(n403), .B(n400), .S(n8230), .Z(n404) );
  MUX2_X1 U19354 ( .A(\mem[614][0] ), .B(\mem[615][0] ), .S(n8406), .Z(n405)
         );
  MUX2_X1 U19355 ( .A(\mem[612][0] ), .B(\mem[613][0] ), .S(n8406), .Z(n406)
         );
  MUX2_X1 U19356 ( .A(n406), .B(n405), .S(n8334), .Z(n407) );
  MUX2_X1 U19357 ( .A(\mem[610][0] ), .B(\mem[611][0] ), .S(n8406), .Z(n408)
         );
  MUX2_X1 U19358 ( .A(\mem[608][0] ), .B(\mem[609][0] ), .S(n8406), .Z(n409)
         );
  MUX2_X1 U19359 ( .A(n409), .B(n408), .S(n8289), .Z(n410) );
  MUX2_X1 U19360 ( .A(n410), .B(n407), .S(n8230), .Z(n411) );
  MUX2_X1 U19361 ( .A(n411), .B(n404), .S(n8211), .Z(n412) );
  MUX2_X1 U19362 ( .A(n412), .B(n397), .S(n8191), .Z(n413) );
  MUX2_X1 U19363 ( .A(\mem[606][0] ), .B(\mem[607][0] ), .S(n8426), .Z(n414)
         );
  MUX2_X1 U19364 ( .A(\mem[604][0] ), .B(\mem[605][0] ), .S(n8488), .Z(n415)
         );
  MUX2_X1 U19365 ( .A(n415), .B(n414), .S(n8297), .Z(n416) );
  MUX2_X1 U19366 ( .A(\mem[602][0] ), .B(\mem[603][0] ), .S(n8462), .Z(n417)
         );
  MUX2_X1 U19367 ( .A(\mem[600][0] ), .B(\mem[601][0] ), .S(n8437), .Z(n418)
         );
  MUX2_X1 U19368 ( .A(n418), .B(n417), .S(n8298), .Z(n419) );
  MUX2_X1 U19369 ( .A(n419), .B(n416), .S(n8231), .Z(n420) );
  MUX2_X1 U19370 ( .A(\mem[598][0] ), .B(\mem[599][0] ), .S(n8424), .Z(n421)
         );
  MUX2_X1 U19371 ( .A(\mem[596][0] ), .B(\mem[597][0] ), .S(n8358), .Z(n422)
         );
  MUX2_X1 U19372 ( .A(n422), .B(n421), .S(n8293), .Z(n423) );
  MUX2_X1 U19373 ( .A(\mem[594][0] ), .B(\mem[595][0] ), .S(n8529), .Z(n424)
         );
  MUX2_X1 U19374 ( .A(\mem[592][0] ), .B(\mem[593][0] ), .S(n8446), .Z(n425)
         );
  MUX2_X1 U19375 ( .A(n425), .B(n424), .S(n8294), .Z(n426) );
  MUX2_X1 U19376 ( .A(n426), .B(n423), .S(n8231), .Z(n427) );
  MUX2_X1 U19377 ( .A(n427), .B(n420), .S(n8216), .Z(n428) );
  MUX2_X1 U19378 ( .A(\mem[590][0] ), .B(\mem[591][0] ), .S(n8361), .Z(n429)
         );
  MUX2_X1 U19379 ( .A(\mem[588][0] ), .B(\mem[589][0] ), .S(n8448), .Z(n430)
         );
  MUX2_X1 U19380 ( .A(n430), .B(n429), .S(n8295), .Z(n431) );
  MUX2_X1 U19381 ( .A(\mem[586][0] ), .B(\mem[587][0] ), .S(n8452), .Z(n432)
         );
  MUX2_X1 U19382 ( .A(\mem[584][0] ), .B(\mem[585][0] ), .S(n8368), .Z(n433)
         );
  MUX2_X1 U19383 ( .A(n433), .B(n432), .S(n8302), .Z(n434) );
  MUX2_X1 U19384 ( .A(n434), .B(n431), .S(n8231), .Z(n435) );
  MUX2_X1 U19385 ( .A(\mem[582][0] ), .B(\mem[583][0] ), .S(n8463), .Z(n436)
         );
  MUX2_X1 U19386 ( .A(\mem[580][0] ), .B(\mem[581][0] ), .S(n8444), .Z(n437)
         );
  MUX2_X1 U19387 ( .A(n437), .B(n436), .S(n8303), .Z(n438) );
  MUX2_X1 U19388 ( .A(\mem[578][0] ), .B(\mem[579][0] ), .S(n8425), .Z(n439)
         );
  MUX2_X1 U19389 ( .A(\mem[576][0] ), .B(\mem[577][0] ), .S(n8358), .Z(n440)
         );
  MUX2_X1 U19390 ( .A(n440), .B(n439), .S(n8304), .Z(n441) );
  MUX2_X1 U19391 ( .A(n441), .B(n438), .S(n8231), .Z(n442) );
  MUX2_X1 U19392 ( .A(n442), .B(n435), .S(n8217), .Z(n443) );
  MUX2_X1 U19393 ( .A(n443), .B(n428), .S(N22), .Z(n444) );
  MUX2_X1 U19394 ( .A(n444), .B(n413), .S(n8184), .Z(n445) );
  MUX2_X1 U19395 ( .A(\mem[574][0] ), .B(\mem[575][0] ), .S(n8474), .Z(n446)
         );
  MUX2_X1 U19396 ( .A(\mem[572][0] ), .B(\mem[573][0] ), .S(n8367), .Z(n447)
         );
  MUX2_X1 U19397 ( .A(n447), .B(n446), .S(n8299), .Z(n448) );
  MUX2_X1 U19398 ( .A(\mem[570][0] ), .B(\mem[571][0] ), .S(n8507), .Z(n449)
         );
  MUX2_X1 U19399 ( .A(\mem[568][0] ), .B(\mem[569][0] ), .S(n8366), .Z(n450)
         );
  MUX2_X1 U19400 ( .A(n450), .B(n449), .S(n8300), .Z(n451) );
  MUX2_X1 U19401 ( .A(n451), .B(n448), .S(n8231), .Z(n452) );
  MUX2_X1 U19402 ( .A(\mem[566][0] ), .B(\mem[567][0] ), .S(n8485), .Z(n453)
         );
  MUX2_X1 U19403 ( .A(\mem[564][0] ), .B(\mem[565][0] ), .S(n8440), .Z(n454)
         );
  MUX2_X1 U19404 ( .A(n454), .B(n453), .S(n8301), .Z(n455) );
  MUX2_X1 U19405 ( .A(\mem[562][0] ), .B(\mem[563][0] ), .S(n8461), .Z(n456)
         );
  MUX2_X1 U19406 ( .A(\mem[560][0] ), .B(\mem[561][0] ), .S(n8451), .Z(n457)
         );
  MUX2_X1 U19407 ( .A(n457), .B(n456), .S(n8326), .Z(n458) );
  MUX2_X1 U19408 ( .A(n458), .B(n455), .S(n8231), .Z(n459) );
  MUX2_X1 U19409 ( .A(n459), .B(n452), .S(n8218), .Z(n460) );
  MUX2_X1 U19410 ( .A(\mem[558][0] ), .B(\mem[559][0] ), .S(n8374), .Z(n461)
         );
  MUX2_X1 U19411 ( .A(\mem[556][0] ), .B(\mem[557][0] ), .S(n8376), .Z(n462)
         );
  MUX2_X1 U19412 ( .A(n462), .B(n461), .S(n8324), .Z(n463) );
  MUX2_X1 U19413 ( .A(\mem[554][0] ), .B(\mem[555][0] ), .S(n8380), .Z(n464)
         );
  MUX2_X1 U19414 ( .A(\mem[552][0] ), .B(\mem[553][0] ), .S(n8427), .Z(n465)
         );
  MUX2_X1 U19415 ( .A(n465), .B(n464), .S(n8291), .Z(n466) );
  MUX2_X1 U19416 ( .A(n466), .B(n463), .S(n8231), .Z(n467) );
  MUX2_X1 U19417 ( .A(\mem[550][0] ), .B(\mem[551][0] ), .S(n8432), .Z(n468)
         );
  MUX2_X1 U19418 ( .A(\mem[548][0] ), .B(\mem[549][0] ), .S(n8403), .Z(n469)
         );
  MUX2_X1 U19419 ( .A(n469), .B(n468), .S(n8285), .Z(n470) );
  MUX2_X1 U19420 ( .A(\mem[546][0] ), .B(\mem[547][0] ), .S(n8492), .Z(n471)
         );
  MUX2_X1 U19421 ( .A(\mem[544][0] ), .B(\mem[545][0] ), .S(n8435), .Z(n472)
         );
  MUX2_X1 U19422 ( .A(n472), .B(n471), .S(n8330), .Z(n473) );
  MUX2_X1 U19423 ( .A(n473), .B(n470), .S(n8231), .Z(n474) );
  MUX2_X1 U19424 ( .A(n474), .B(n467), .S(n8207), .Z(n475) );
  MUX2_X1 U19425 ( .A(n475), .B(n460), .S(n8195), .Z(n476) );
  MUX2_X1 U19426 ( .A(\mem[542][0] ), .B(\mem[543][0] ), .S(n8468), .Z(n477)
         );
  MUX2_X1 U19427 ( .A(\mem[540][0] ), .B(\mem[541][0] ), .S(n8452), .Z(n478)
         );
  MUX2_X1 U19428 ( .A(n478), .B(n477), .S(n8297), .Z(n479) );
  MUX2_X1 U19429 ( .A(\mem[538][0] ), .B(\mem[539][0] ), .S(n8427), .Z(n480)
         );
  MUX2_X1 U19430 ( .A(\mem[536][0] ), .B(\mem[537][0] ), .S(n8424), .Z(n481)
         );
  MUX2_X1 U19431 ( .A(n481), .B(n480), .S(n8279), .Z(n482) );
  MUX2_X1 U19432 ( .A(n482), .B(n479), .S(n8231), .Z(n483) );
  MUX2_X1 U19433 ( .A(\mem[534][0] ), .B(\mem[535][0] ), .S(n8385), .Z(n484)
         );
  MUX2_X1 U19434 ( .A(\mem[532][0] ), .B(\mem[533][0] ), .S(n8384), .Z(n485)
         );
  MUX2_X1 U19435 ( .A(n485), .B(n484), .S(n8284), .Z(n486) );
  MUX2_X1 U19436 ( .A(\mem[530][0] ), .B(\mem[531][0] ), .S(n8383), .Z(n487)
         );
  MUX2_X1 U19437 ( .A(\mem[528][0] ), .B(\mem[529][0] ), .S(n8360), .Z(n488)
         );
  MUX2_X1 U19438 ( .A(n488), .B(n487), .S(n8285), .Z(n489) );
  MUX2_X1 U19439 ( .A(n489), .B(n486), .S(n8231), .Z(n490) );
  MUX2_X1 U19440 ( .A(n490), .B(n483), .S(n8208), .Z(n491) );
  MUX2_X1 U19441 ( .A(\mem[526][0] ), .B(\mem[527][0] ), .S(n8484), .Z(n492)
         );
  MUX2_X1 U19442 ( .A(\mem[524][0] ), .B(\mem[525][0] ), .S(n8439), .Z(n493)
         );
  MUX2_X1 U19443 ( .A(n493), .B(n492), .S(n8286), .Z(n494) );
  MUX2_X1 U19444 ( .A(\mem[522][0] ), .B(\mem[523][0] ), .S(n8460), .Z(n495)
         );
  MUX2_X1 U19445 ( .A(\mem[520][0] ), .B(\mem[521][0] ), .S(n8450), .Z(n496)
         );
  MUX2_X1 U19446 ( .A(n496), .B(n495), .S(n8290), .Z(n497) );
  MUX2_X1 U19447 ( .A(n497), .B(n494), .S(n8231), .Z(n498) );
  MUX2_X1 U19448 ( .A(\mem[518][0] ), .B(\mem[519][0] ), .S(n8455), .Z(n499)
         );
  MUX2_X1 U19449 ( .A(\mem[516][0] ), .B(\mem[517][0] ), .S(n8436), .Z(n500)
         );
  MUX2_X1 U19450 ( .A(n500), .B(n499), .S(n8291), .Z(n501) );
  MUX2_X1 U19451 ( .A(\mem[514][0] ), .B(\mem[515][0] ), .S(n8423), .Z(n502)
         );
  MUX2_X1 U19452 ( .A(\mem[512][0] ), .B(\mem[513][0] ), .S(n8358), .Z(n503)
         );
  MUX2_X1 U19453 ( .A(n503), .B(n502), .S(n8292), .Z(n504) );
  MUX2_X1 U19454 ( .A(n504), .B(n501), .S(n8231), .Z(n505) );
  MUX2_X1 U19455 ( .A(n505), .B(n498), .S(n8209), .Z(n506) );
  MUX2_X1 U19456 ( .A(n506), .B(n491), .S(N22), .Z(n507) );
  MUX2_X1 U19457 ( .A(n507), .B(n476), .S(N23), .Z(n508) );
  MUX2_X1 U19458 ( .A(n508), .B(n445), .S(n8178), .Z(n509) );
  MUX2_X1 U19459 ( .A(n509), .B(n382), .S(N25), .Z(n510) );
  MUX2_X1 U19460 ( .A(n510), .B(n255), .S(N26), .Z(n511) );
  MUX2_X1 U19461 ( .A(\mem[510][0] ), .B(\mem[511][0] ), .S(n8463), .Z(n512)
         );
  MUX2_X1 U19462 ( .A(\mem[508][0] ), .B(\mem[509][0] ), .S(n8473), .Z(n513)
         );
  MUX2_X1 U19463 ( .A(n513), .B(n512), .S(n8276), .Z(n514) );
  MUX2_X1 U19464 ( .A(\mem[506][0] ), .B(\mem[507][0] ), .S(n8423), .Z(n515)
         );
  MUX2_X1 U19465 ( .A(\mem[504][0] ), .B(\mem[505][0] ), .S(n8520), .Z(n516)
         );
  MUX2_X1 U19466 ( .A(n516), .B(n515), .S(n8319), .Z(n517) );
  MUX2_X1 U19467 ( .A(n517), .B(n514), .S(n8232), .Z(n518) );
  MUX2_X1 U19468 ( .A(\mem[502][0] ), .B(\mem[503][0] ), .S(n8467), .Z(n519)
         );
  MUX2_X1 U19469 ( .A(\mem[500][0] ), .B(\mem[501][0] ), .S(n8401), .Z(n520)
         );
  MUX2_X1 U19470 ( .A(n520), .B(n519), .S(n8266), .Z(n521) );
  MUX2_X1 U19471 ( .A(\mem[498][0] ), .B(\mem[499][0] ), .S(n8422), .Z(n522)
         );
  MUX2_X1 U19472 ( .A(\mem[496][0] ), .B(\mem[497][0] ), .S(n8452), .Z(n523)
         );
  MUX2_X1 U19473 ( .A(n523), .B(n522), .S(n8268), .Z(n524) );
  MUX2_X1 U19474 ( .A(n524), .B(n521), .S(n8232), .Z(n525) );
  MUX2_X1 U19475 ( .A(n525), .B(n518), .S(n8204), .Z(n526) );
  MUX2_X1 U19476 ( .A(\mem[494][0] ), .B(\mem[495][0] ), .S(n8398), .Z(n527)
         );
  MUX2_X1 U19477 ( .A(\mem[492][0] ), .B(\mem[493][0] ), .S(n8464), .Z(n528)
         );
  MUX2_X1 U19478 ( .A(n528), .B(n527), .S(n8269), .Z(n529) );
  MUX2_X1 U19479 ( .A(\mem[490][0] ), .B(\mem[491][0] ), .S(n8536), .Z(n530)
         );
  MUX2_X1 U19480 ( .A(\mem[488][0] ), .B(\mem[489][0] ), .S(n8507), .Z(n531)
         );
  MUX2_X1 U19481 ( .A(n531), .B(n530), .S(n8270), .Z(n532) );
  MUX2_X1 U19482 ( .A(n532), .B(n529), .S(n8232), .Z(n533) );
  MUX2_X1 U19483 ( .A(\mem[486][0] ), .B(\mem[487][0] ), .S(n8419), .Z(n534)
         );
  MUX2_X1 U19484 ( .A(\mem[484][0] ), .B(\mem[485][0] ), .S(n8375), .Z(n535)
         );
  MUX2_X1 U19485 ( .A(n535), .B(n534), .S(n8318), .Z(n536) );
  MUX2_X1 U19486 ( .A(\mem[482][0] ), .B(\mem[483][0] ), .S(n8472), .Z(n537)
         );
  MUX2_X1 U19487 ( .A(\mem[480][0] ), .B(\mem[481][0] ), .S(n8464), .Z(n538)
         );
  MUX2_X1 U19488 ( .A(n538), .B(n537), .S(n8312), .Z(n539) );
  MUX2_X1 U19489 ( .A(n539), .B(n536), .S(n8232), .Z(n540) );
  MUX2_X1 U19490 ( .A(n540), .B(n533), .S(n8206), .Z(n541) );
  MUX2_X1 U19491 ( .A(n541), .B(n526), .S(n8196), .Z(n542) );
  MUX2_X1 U19492 ( .A(\mem[478][0] ), .B(\mem[479][0] ), .S(n8402), .Z(n543)
         );
  MUX2_X1 U19493 ( .A(\mem[476][0] ), .B(\mem[477][0] ), .S(n8496), .Z(n544)
         );
  MUX2_X1 U19494 ( .A(n544), .B(n543), .S(n8298), .Z(n545) );
  MUX2_X1 U19495 ( .A(\mem[474][0] ), .B(\mem[475][0] ), .S(n8449), .Z(n546)
         );
  MUX2_X1 U19496 ( .A(\mem[472][0] ), .B(\mem[473][0] ), .S(n8415), .Z(n547)
         );
  MUX2_X1 U19497 ( .A(n547), .B(n546), .S(n8306), .Z(n548) );
  MUX2_X1 U19498 ( .A(n548), .B(n545), .S(n8232), .Z(n549) );
  MUX2_X1 U19499 ( .A(\mem[470][0] ), .B(\mem[471][0] ), .S(n8433), .Z(n550)
         );
  MUX2_X1 U19500 ( .A(\mem[468][0] ), .B(\mem[469][0] ), .S(n8396), .Z(n551)
         );
  MUX2_X1 U19501 ( .A(n551), .B(n550), .S(n8276), .Z(n552) );
  MUX2_X1 U19502 ( .A(\mem[466][0] ), .B(\mem[467][0] ), .S(n8365), .Z(n553)
         );
  MUX2_X1 U19503 ( .A(\mem[464][0] ), .B(\mem[465][0] ), .S(n8404), .Z(n554)
         );
  MUX2_X1 U19504 ( .A(n554), .B(n553), .S(n8350), .Z(n555) );
  MUX2_X1 U19505 ( .A(n555), .B(n552), .S(n8232), .Z(n556) );
  MUX2_X1 U19506 ( .A(n556), .B(n549), .S(n8205), .Z(n557) );
  MUX2_X1 U19507 ( .A(\mem[462][0] ), .B(\mem[463][0] ), .S(n8477), .Z(n558)
         );
  MUX2_X1 U19508 ( .A(\mem[460][0] ), .B(\mem[461][0] ), .S(n8514), .Z(n559)
         );
  MUX2_X1 U19509 ( .A(n559), .B(n558), .S(n8266), .Z(n560) );
  MUX2_X1 U19510 ( .A(\mem[458][0] ), .B(\mem[459][0] ), .S(n8383), .Z(n561)
         );
  MUX2_X1 U19511 ( .A(\mem[456][0] ), .B(\mem[457][0] ), .S(n8538), .Z(n562)
         );
  MUX2_X1 U19512 ( .A(n562), .B(n561), .S(n8269), .Z(n563) );
  MUX2_X1 U19513 ( .A(n563), .B(n560), .S(n8232), .Z(n564) );
  MUX2_X1 U19514 ( .A(\mem[454][0] ), .B(\mem[455][0] ), .S(n8414), .Z(n565)
         );
  MUX2_X1 U19515 ( .A(\mem[452][0] ), .B(\mem[453][0] ), .S(n8385), .Z(n566)
         );
  MUX2_X1 U19516 ( .A(n566), .B(n565), .S(n8356), .Z(n567) );
  MUX2_X1 U19517 ( .A(\mem[450][0] ), .B(\mem[451][0] ), .S(n8384), .Z(n568)
         );
  MUX2_X1 U19518 ( .A(\mem[448][0] ), .B(\mem[449][0] ), .S(n8426), .Z(n569)
         );
  MUX2_X1 U19519 ( .A(n569), .B(n568), .S(n8271), .Z(n570) );
  MUX2_X1 U19520 ( .A(n570), .B(n567), .S(n8232), .Z(n571) );
  MUX2_X1 U19521 ( .A(n571), .B(n564), .S(n8211), .Z(n572) );
  MUX2_X1 U19522 ( .A(n572), .B(n557), .S(n8191), .Z(n573) );
  MUX2_X1 U19523 ( .A(n573), .B(n542), .S(n8181), .Z(n574) );
  MUX2_X1 U19524 ( .A(\mem[446][0] ), .B(\mem[447][0] ), .S(n8432), .Z(n575)
         );
  MUX2_X1 U19525 ( .A(\mem[444][0] ), .B(\mem[445][0] ), .S(n8469), .Z(n576)
         );
  MUX2_X1 U19526 ( .A(n576), .B(n575), .S(n8349), .Z(n577) );
  MUX2_X1 U19527 ( .A(\mem[442][0] ), .B(\mem[443][0] ), .S(n8400), .Z(n578)
         );
  MUX2_X1 U19528 ( .A(\mem[440][0] ), .B(\mem[441][0] ), .S(n8367), .Z(n579)
         );
  MUX2_X1 U19529 ( .A(n579), .B(n578), .S(n8310), .Z(n580) );
  MUX2_X1 U19530 ( .A(n580), .B(n577), .S(n8232), .Z(n581) );
  MUX2_X1 U19531 ( .A(\mem[438][0] ), .B(\mem[439][0] ), .S(n8454), .Z(n582)
         );
  MUX2_X1 U19532 ( .A(\mem[436][0] ), .B(\mem[437][0] ), .S(n8435), .Z(n583)
         );
  MUX2_X1 U19533 ( .A(n583), .B(n582), .S(n8281), .Z(n584) );
  MUX2_X1 U19534 ( .A(\mem[434][0] ), .B(\mem[435][0] ), .S(n8361), .Z(n585)
         );
  MUX2_X1 U19535 ( .A(\mem[432][0] ), .B(\mem[433][0] ), .S(n8399), .Z(n586)
         );
  MUX2_X1 U19536 ( .A(n586), .B(n585), .S(n8352), .Z(n587) );
  MUX2_X1 U19537 ( .A(n587), .B(n584), .S(n8232), .Z(n588) );
  MUX2_X1 U19538 ( .A(n588), .B(n581), .S(n8198), .Z(n589) );
  MUX2_X1 U19539 ( .A(\mem[430][0] ), .B(\mem[431][0] ), .S(n8483), .Z(n590)
         );
  MUX2_X1 U19540 ( .A(\mem[428][0] ), .B(\mem[429][0] ), .S(n8418), .Z(n591)
         );
  MUX2_X1 U19541 ( .A(n591), .B(n590), .S(n8266), .Z(n592) );
  MUX2_X1 U19542 ( .A(\mem[426][0] ), .B(\mem[427][0] ), .S(n8428), .Z(n593)
         );
  MUX2_X1 U19543 ( .A(\mem[424][0] ), .B(\mem[425][0] ), .S(n8358), .Z(n594)
         );
  MUX2_X1 U19544 ( .A(n594), .B(n593), .S(n8267), .Z(n595) );
  MUX2_X1 U19545 ( .A(n595), .B(n592), .S(n8232), .Z(n596) );
  MUX2_X1 U19546 ( .A(\mem[422][0] ), .B(\mem[423][0] ), .S(n8360), .Z(n597)
         );
  MUX2_X1 U19547 ( .A(\mem[420][0] ), .B(\mem[421][0] ), .S(n8443), .Z(n598)
         );
  MUX2_X1 U19548 ( .A(n598), .B(n597), .S(n8271), .Z(n599) );
  MUX2_X1 U19549 ( .A(\mem[418][0] ), .B(\mem[419][0] ), .S(n8538), .Z(n600)
         );
  MUX2_X1 U19550 ( .A(\mem[416][0] ), .B(\mem[417][0] ), .S(n8359), .Z(n601)
         );
  MUX2_X1 U19551 ( .A(n601), .B(n600), .S(n8349), .Z(n602) );
  MUX2_X1 U19552 ( .A(n602), .B(n599), .S(n8232), .Z(n603) );
  MUX2_X1 U19553 ( .A(n603), .B(n596), .S(n8207), .Z(n604) );
  MUX2_X1 U19554 ( .A(n604), .B(n589), .S(n8194), .Z(n605) );
  MUX2_X1 U19555 ( .A(\mem[414][0] ), .B(\mem[415][0] ), .S(n8382), .Z(n606)
         );
  MUX2_X1 U19556 ( .A(\mem[412][0] ), .B(\mem[413][0] ), .S(n8381), .Z(n607)
         );
  MUX2_X1 U19557 ( .A(n607), .B(n606), .S(n8267), .Z(n608) );
  MUX2_X1 U19558 ( .A(\mem[410][0] ), .B(\mem[411][0] ), .S(n8380), .Z(n609)
         );
  MUX2_X1 U19559 ( .A(\mem[408][0] ), .B(\mem[409][0] ), .S(n8379), .Z(n610)
         );
  MUX2_X1 U19560 ( .A(n610), .B(n609), .S(n8273), .Z(n611) );
  MUX2_X1 U19561 ( .A(n611), .B(n608), .S(n8233), .Z(n612) );
  MUX2_X1 U19562 ( .A(\mem[406][0] ), .B(\mem[407][0] ), .S(n8378), .Z(n613)
         );
  MUX2_X1 U19563 ( .A(\mem[404][0] ), .B(\mem[405][0] ), .S(n8377), .Z(n614)
         );
  MUX2_X1 U19564 ( .A(n614), .B(n613), .S(N19), .Z(n615) );
  MUX2_X1 U19565 ( .A(\mem[402][0] ), .B(\mem[403][0] ), .S(n8376), .Z(n616)
         );
  MUX2_X1 U19566 ( .A(\mem[400][0] ), .B(\mem[401][0] ), .S(n8375), .Z(n617)
         );
  MUX2_X1 U19567 ( .A(n617), .B(n616), .S(n8350), .Z(n618) );
  MUX2_X1 U19568 ( .A(n618), .B(n615), .S(n8233), .Z(n619) );
  MUX2_X1 U19569 ( .A(n619), .B(n612), .S(n8201), .Z(n620) );
  MUX2_X1 U19570 ( .A(\mem[398][0] ), .B(\mem[399][0] ), .S(n8374), .Z(n621)
         );
  MUX2_X1 U19571 ( .A(\mem[396][0] ), .B(\mem[397][0] ), .S(n8438), .Z(n622)
         );
  MUX2_X1 U19572 ( .A(n622), .B(n621), .S(n8270), .Z(n623) );
  MUX2_X1 U19573 ( .A(\mem[394][0] ), .B(\mem[395][0] ), .S(n8459), .Z(n624)
         );
  MUX2_X1 U19574 ( .A(\mem[392][0] ), .B(\mem[393][0] ), .S(n8501), .Z(n625)
         );
  MUX2_X1 U19575 ( .A(n625), .B(n624), .S(n8327), .Z(n626) );
  MUX2_X1 U19576 ( .A(n626), .B(n623), .S(n8233), .Z(n627) );
  MUX2_X1 U19577 ( .A(\mem[390][0] ), .B(\mem[391][0] ), .S(n8500), .Z(n628)
         );
  MUX2_X1 U19578 ( .A(\mem[388][0] ), .B(\mem[389][0] ), .S(n8361), .Z(n629)
         );
  MUX2_X1 U19579 ( .A(n629), .B(n628), .S(n8272), .Z(n630) );
  MUX2_X1 U19580 ( .A(\mem[386][0] ), .B(\mem[387][0] ), .S(n8477), .Z(n631)
         );
  MUX2_X1 U19581 ( .A(\mem[384][0] ), .B(\mem[385][0] ), .S(n8469), .Z(n632)
         );
  MUX2_X1 U19582 ( .A(n632), .B(n631), .S(n8271), .Z(n633) );
  MUX2_X1 U19583 ( .A(n633), .B(n630), .S(n8233), .Z(n634) );
  MUX2_X1 U19584 ( .A(n634), .B(n627), .S(n8200), .Z(n635) );
  MUX2_X1 U19585 ( .A(n635), .B(n620), .S(N22), .Z(n636) );
  MUX2_X1 U19586 ( .A(n636), .B(n605), .S(n8181), .Z(n637) );
  MUX2_X1 U19587 ( .A(n637), .B(n574), .S(n8179), .Z(n638) );
  MUX2_X1 U19588 ( .A(\mem[382][0] ), .B(\mem[383][0] ), .S(n8488), .Z(n639)
         );
  MUX2_X1 U19589 ( .A(\mem[380][0] ), .B(\mem[381][0] ), .S(n8453), .Z(n640)
         );
  MUX2_X1 U19590 ( .A(n640), .B(n639), .S(n8268), .Z(n641) );
  MUX2_X1 U19591 ( .A(\mem[378][0] ), .B(\mem[379][0] ), .S(n8431), .Z(n642)
         );
  MUX2_X1 U19592 ( .A(\mem[376][0] ), .B(\mem[377][0] ), .S(n8406), .Z(n643)
         );
  MUX2_X1 U19593 ( .A(n643), .B(n642), .S(n8270), .Z(n644) );
  MUX2_X1 U19594 ( .A(n644), .B(n641), .S(n8233), .Z(n645) );
  MUX2_X1 U19595 ( .A(\mem[374][0] ), .B(\mem[375][0] ), .S(n8440), .Z(n646)
         );
  MUX2_X1 U19596 ( .A(\mem[372][0] ), .B(\mem[373][0] ), .S(n8427), .Z(n647)
         );
  MUX2_X1 U19597 ( .A(n647), .B(n646), .S(n8313), .Z(n648) );
  MUX2_X1 U19598 ( .A(\mem[370][0] ), .B(\mem[371][0] ), .S(n8358), .Z(n649)
         );
  MUX2_X1 U19599 ( .A(\mem[368][0] ), .B(\mem[369][0] ), .S(n8360), .Z(n650)
         );
  MUX2_X1 U19600 ( .A(n650), .B(n649), .S(n8285), .Z(n651) );
  MUX2_X1 U19601 ( .A(n651), .B(n648), .S(n8233), .Z(n652) );
  MUX2_X1 U19602 ( .A(n652), .B(n645), .S(n8213), .Z(n653) );
  MUX2_X1 U19603 ( .A(\mem[366][0] ), .B(\mem[367][0] ), .S(n8381), .Z(n654)
         );
  MUX2_X1 U19604 ( .A(\mem[364][0] ), .B(\mem[365][0] ), .S(n8380), .Z(n655)
         );
  MUX2_X1 U19605 ( .A(n655), .B(n654), .S(n8313), .Z(n656) );
  MUX2_X1 U19606 ( .A(\mem[362][0] ), .B(\mem[363][0] ), .S(n8379), .Z(n657)
         );
  MUX2_X1 U19607 ( .A(\mem[360][0] ), .B(\mem[361][0] ), .S(n8378), .Z(n658)
         );
  MUX2_X1 U19608 ( .A(n658), .B(n657), .S(n8282), .Z(n659) );
  MUX2_X1 U19609 ( .A(n659), .B(n656), .S(n8233), .Z(n660) );
  MUX2_X1 U19610 ( .A(\mem[358][0] ), .B(\mem[359][0] ), .S(n8377), .Z(n661)
         );
  MUX2_X1 U19611 ( .A(\mem[356][0] ), .B(\mem[357][0] ), .S(n8376), .Z(n662)
         );
  MUX2_X1 U19612 ( .A(n662), .B(n661), .S(n8282), .Z(n663) );
  MUX2_X1 U19613 ( .A(\mem[354][0] ), .B(\mem[355][0] ), .S(n8375), .Z(n664)
         );
  MUX2_X1 U19614 ( .A(\mem[352][0] ), .B(\mem[353][0] ), .S(n8466), .Z(n665)
         );
  MUX2_X1 U19615 ( .A(n665), .B(n664), .S(n8328), .Z(n666) );
  MUX2_X1 U19616 ( .A(n666), .B(n663), .S(n8233), .Z(n667) );
  MUX2_X1 U19617 ( .A(n667), .B(n660), .S(n8202), .Z(n668) );
  MUX2_X1 U19618 ( .A(n668), .B(n653), .S(n8196), .Z(n669) );
  MUX2_X1 U19619 ( .A(\mem[350][0] ), .B(\mem[351][0] ), .S(n8374), .Z(n670)
         );
  MUX2_X1 U19620 ( .A(\mem[348][0] ), .B(\mem[349][0] ), .S(n8382), .Z(n671)
         );
  MUX2_X1 U19621 ( .A(n671), .B(n670), .S(n8280), .Z(n672) );
  MUX2_X1 U19622 ( .A(\mem[346][0] ), .B(\mem[347][0] ), .S(n8464), .Z(n673)
         );
  MUX2_X1 U19623 ( .A(\mem[344][0] ), .B(\mem[345][0] ), .S(n8453), .Z(n674)
         );
  MUX2_X1 U19624 ( .A(n674), .B(n673), .S(n8279), .Z(n675) );
  MUX2_X1 U19625 ( .A(n675), .B(n672), .S(n8233), .Z(n676) );
  MUX2_X1 U19626 ( .A(\mem[342][0] ), .B(\mem[343][0] ), .S(n8363), .Z(n677)
         );
  MUX2_X1 U19627 ( .A(\mem[340][0] ), .B(\mem[341][0] ), .S(n8372), .Z(n678)
         );
  MUX2_X1 U19628 ( .A(n678), .B(n677), .S(n8331), .Z(n679) );
  MUX2_X1 U19629 ( .A(\mem[338][0] ), .B(\mem[339][0] ), .S(n8361), .Z(n680)
         );
  MUX2_X1 U19630 ( .A(\mem[336][0] ), .B(\mem[337][0] ), .S(n8499), .Z(n681)
         );
  MUX2_X1 U19631 ( .A(n681), .B(n680), .S(n8278), .Z(n682) );
  MUX2_X1 U19632 ( .A(n682), .B(n679), .S(n8233), .Z(n683) );
  MUX2_X1 U19633 ( .A(n683), .B(n676), .S(n8203), .Z(n684) );
  MUX2_X1 U19634 ( .A(\mem[334][0] ), .B(\mem[335][0] ), .S(n8465), .Z(n685)
         );
  MUX2_X1 U19635 ( .A(\mem[332][0] ), .B(\mem[333][0] ), .S(n8405), .Z(n686)
         );
  MUX2_X1 U19636 ( .A(n686), .B(n685), .S(n8277), .Z(n687) );
  MUX2_X1 U19637 ( .A(\mem[330][0] ), .B(\mem[331][0] ), .S(n8420), .Z(n688)
         );
  MUX2_X1 U19638 ( .A(\mem[328][0] ), .B(\mem[329][0] ), .S(n8450), .Z(n689)
         );
  MUX2_X1 U19639 ( .A(n689), .B(n688), .S(n8276), .Z(n690) );
  MUX2_X1 U19640 ( .A(n690), .B(n687), .S(n8233), .Z(n691) );
  MUX2_X1 U19641 ( .A(\mem[326][0] ), .B(\mem[327][0] ), .S(n8532), .Z(n692)
         );
  MUX2_X1 U19642 ( .A(\mem[324][0] ), .B(\mem[325][0] ), .S(n8462), .Z(n693)
         );
  MUX2_X1 U19643 ( .A(n693), .B(n692), .S(n8275), .Z(n694) );
  MUX2_X1 U19644 ( .A(\mem[322][0] ), .B(\mem[323][0] ), .S(n8534), .Z(n695)
         );
  MUX2_X1 U19645 ( .A(\mem[320][0] ), .B(\mem[321][0] ), .S(n8511), .Z(n696)
         );
  MUX2_X1 U19646 ( .A(n696), .B(n695), .S(n8274), .Z(n697) );
  MUX2_X1 U19647 ( .A(n697), .B(n694), .S(n8233), .Z(n698) );
  MUX2_X1 U19648 ( .A(n698), .B(n691), .S(n8204), .Z(n699) );
  MUX2_X1 U19649 ( .A(n699), .B(n684), .S(n8195), .Z(n700) );
  MUX2_X1 U19650 ( .A(n700), .B(n669), .S(n8181), .Z(n701) );
  MUX2_X1 U19651 ( .A(\mem[318][0] ), .B(\mem[319][0] ), .S(n8372), .Z(n702)
         );
  MUX2_X1 U19652 ( .A(\mem[316][0] ), .B(\mem[317][0] ), .S(n8438), .Z(n703)
         );
  MUX2_X1 U19653 ( .A(n703), .B(n702), .S(n8355), .Z(n704) );
  MUX2_X1 U19654 ( .A(\mem[314][0] ), .B(\mem[315][0] ), .S(n8456), .Z(n705)
         );
  MUX2_X1 U19655 ( .A(\mem[312][0] ), .B(\mem[313][0] ), .S(n8430), .Z(n706)
         );
  MUX2_X1 U19656 ( .A(n706), .B(n705), .S(n8356), .Z(n707) );
  MUX2_X1 U19657 ( .A(n707), .B(n704), .S(n8234), .Z(n708) );
  MUX2_X1 U19658 ( .A(\mem[310][0] ), .B(\mem[311][0] ), .S(n8455), .Z(n709)
         );
  MUX2_X1 U19659 ( .A(\mem[308][0] ), .B(\mem[309][0] ), .S(n8446), .Z(n710)
         );
  MUX2_X1 U19660 ( .A(n710), .B(n709), .S(n8275), .Z(n711) );
  MUX2_X1 U19661 ( .A(\mem[306][0] ), .B(\mem[307][0] ), .S(n8407), .Z(n712)
         );
  MUX2_X1 U19662 ( .A(\mem[304][0] ), .B(\mem[305][0] ), .S(n8410), .Z(n713)
         );
  MUX2_X1 U19663 ( .A(n713), .B(n712), .S(n8275), .Z(n714) );
  MUX2_X1 U19664 ( .A(n714), .B(n711), .S(n8234), .Z(n715) );
  MUX2_X1 U19665 ( .A(n715), .B(n708), .S(n8200), .Z(n716) );
  MUX2_X1 U19666 ( .A(\mem[302][0] ), .B(\mem[303][0] ), .S(n8398), .Z(n717)
         );
  MUX2_X1 U19667 ( .A(\mem[300][0] ), .B(\mem[301][0] ), .S(n8371), .Z(n718)
         );
  MUX2_X1 U19668 ( .A(n718), .B(n717), .S(n8290), .Z(n719) );
  MUX2_X1 U19669 ( .A(\mem[298][0] ), .B(\mem[299][0] ), .S(n8437), .Z(n720)
         );
  MUX2_X1 U19670 ( .A(\mem[296][0] ), .B(\mem[297][0] ), .S(n8377), .Z(n721)
         );
  MUX2_X1 U19671 ( .A(n721), .B(n720), .S(n8266), .Z(n722) );
  MUX2_X1 U19672 ( .A(n722), .B(n719), .S(n8234), .Z(n723) );
  MUX2_X1 U19673 ( .A(\mem[294][0] ), .B(\mem[295][0] ), .S(n8360), .Z(n724)
         );
  MUX2_X1 U19674 ( .A(\mem[292][0] ), .B(\mem[293][0] ), .S(n8415), .Z(n725)
         );
  MUX2_X1 U19675 ( .A(n725), .B(n724), .S(n8266), .Z(n726) );
  MUX2_X1 U19676 ( .A(\mem[290][0] ), .B(\mem[291][0] ), .S(n8387), .Z(n727)
         );
  MUX2_X1 U19677 ( .A(\mem[288][0] ), .B(\mem[289][0] ), .S(n8434), .Z(n728)
         );
  MUX2_X1 U19678 ( .A(n728), .B(n727), .S(n8267), .Z(n729) );
  MUX2_X1 U19679 ( .A(n729), .B(n726), .S(n8234), .Z(n730) );
  MUX2_X1 U19680 ( .A(n730), .B(n723), .S(n8200), .Z(n731) );
  MUX2_X1 U19681 ( .A(n731), .B(n716), .S(n8194), .Z(n732) );
  MUX2_X1 U19682 ( .A(\mem[286][0] ), .B(\mem[287][0] ), .S(n8369), .Z(n733)
         );
  MUX2_X1 U19683 ( .A(\mem[284][0] ), .B(\mem[285][0] ), .S(n8376), .Z(n734)
         );
  MUX2_X1 U19684 ( .A(n734), .B(n733), .S(n8268), .Z(n735) );
  MUX2_X1 U19685 ( .A(\mem[282][0] ), .B(\mem[283][0] ), .S(n8476), .Z(n736)
         );
  MUX2_X1 U19686 ( .A(\mem[280][0] ), .B(\mem[281][0] ), .S(n8462), .Z(n737)
         );
  MUX2_X1 U19687 ( .A(n737), .B(n736), .S(n8269), .Z(n738) );
  MUX2_X1 U19688 ( .A(n738), .B(n735), .S(n8234), .Z(n739) );
  MUX2_X1 U19689 ( .A(\mem[278][0] ), .B(\mem[279][0] ), .S(n8533), .Z(n740)
         );
  MUX2_X1 U19690 ( .A(\mem[276][0] ), .B(\mem[277][0] ), .S(n8361), .Z(n741)
         );
  MUX2_X1 U19691 ( .A(n741), .B(n740), .S(n8270), .Z(n742) );
  MUX2_X1 U19692 ( .A(\mem[274][0] ), .B(\mem[275][0] ), .S(n8384), .Z(n743)
         );
  MUX2_X1 U19693 ( .A(\mem[272][0] ), .B(\mem[273][0] ), .S(n8429), .Z(n744)
         );
  MUX2_X1 U19694 ( .A(n744), .B(n743), .S(n8336), .Z(n745) );
  MUX2_X1 U19695 ( .A(n745), .B(n742), .S(n8234), .Z(n746) );
  MUX2_X1 U19696 ( .A(n746), .B(n739), .S(n8212), .Z(n747) );
  MUX2_X1 U19697 ( .A(\mem[270][0] ), .B(\mem[271][0] ), .S(n8463), .Z(n748)
         );
  MUX2_X1 U19698 ( .A(\mem[268][0] ), .B(\mem[269][0] ), .S(n8383), .Z(n749)
         );
  MUX2_X1 U19699 ( .A(n749), .B(n748), .S(n8269), .Z(n750) );
  MUX2_X1 U19700 ( .A(\mem[266][0] ), .B(\mem[267][0] ), .S(n8479), .Z(n751)
         );
  MUX2_X1 U19701 ( .A(\mem[264][0] ), .B(\mem[265][0] ), .S(n8361), .Z(n752)
         );
  MUX2_X1 U19702 ( .A(n752), .B(n751), .S(n8314), .Z(n753) );
  MUX2_X1 U19703 ( .A(n753), .B(n750), .S(n8234), .Z(n754) );
  MUX2_X1 U19704 ( .A(\mem[262][0] ), .B(\mem[263][0] ), .S(n8402), .Z(n755)
         );
  MUX2_X1 U19705 ( .A(\mem[260][0] ), .B(\mem[261][0] ), .S(n8401), .Z(n756)
         );
  MUX2_X1 U19706 ( .A(n756), .B(n755), .S(n8326), .Z(n757) );
  MUX2_X1 U19707 ( .A(\mem[258][0] ), .B(\mem[259][0] ), .S(n8471), .Z(n758)
         );
  MUX2_X1 U19708 ( .A(\mem[256][0] ), .B(\mem[257][0] ), .S(n8463), .Z(n759)
         );
  MUX2_X1 U19709 ( .A(n759), .B(n758), .S(n8272), .Z(n760) );
  MUX2_X1 U19710 ( .A(n760), .B(n757), .S(n8234), .Z(n761) );
  MUX2_X1 U19711 ( .A(n761), .B(n754), .S(N21), .Z(n762) );
  MUX2_X1 U19712 ( .A(n762), .B(n747), .S(n8196), .Z(n763) );
  MUX2_X1 U19713 ( .A(n763), .B(n732), .S(n8181), .Z(n764) );
  MUX2_X1 U19714 ( .A(n764), .B(n701), .S(n8179), .Z(n765) );
  MUX2_X1 U19715 ( .A(n765), .B(n638), .S(N25), .Z(n766) );
  MUX2_X1 U19716 ( .A(\mem[254][0] ), .B(\mem[255][0] ), .S(n8408), .Z(n767)
         );
  MUX2_X1 U19717 ( .A(\mem[252][0] ), .B(\mem[253][0] ), .S(n8442), .Z(n768)
         );
  MUX2_X1 U19718 ( .A(n768), .B(n767), .S(n8271), .Z(n769) );
  MUX2_X1 U19719 ( .A(\mem[250][0] ), .B(\mem[251][0] ), .S(n8377), .Z(n770)
         );
  MUX2_X1 U19720 ( .A(\mem[248][0] ), .B(\mem[249][0] ), .S(n8434), .Z(n771)
         );
  MUX2_X1 U19721 ( .A(n771), .B(n770), .S(n8285), .Z(n772) );
  MUX2_X1 U19722 ( .A(n772), .B(n769), .S(n8234), .Z(n773) );
  MUX2_X1 U19723 ( .A(\mem[246][0] ), .B(\mem[247][0] ), .S(n8395), .Z(n774)
         );
  MUX2_X1 U19724 ( .A(\mem[244][0] ), .B(\mem[245][0] ), .S(n8366), .Z(n775)
         );
  MUX2_X1 U19725 ( .A(n775), .B(n774), .S(n8267), .Z(n776) );
  MUX2_X1 U19726 ( .A(\mem[242][0] ), .B(\mem[243][0] ), .S(n8368), .Z(n777)
         );
  MUX2_X1 U19727 ( .A(\mem[240][0] ), .B(\mem[241][0] ), .S(n8368), .Z(n778)
         );
  MUX2_X1 U19728 ( .A(n778), .B(n777), .S(n8288), .Z(n779) );
  MUX2_X1 U19729 ( .A(n779), .B(n776), .S(n8234), .Z(n780) );
  MUX2_X1 U19730 ( .A(n780), .B(n773), .S(n8199), .Z(n781) );
  MUX2_X1 U19731 ( .A(\mem[238][0] ), .B(\mem[239][0] ), .S(n8364), .Z(n782)
         );
  MUX2_X1 U19732 ( .A(\mem[236][0] ), .B(\mem[237][0] ), .S(n8385), .Z(n783)
         );
  MUX2_X1 U19733 ( .A(n783), .B(n782), .S(n8312), .Z(n784) );
  MUX2_X1 U19734 ( .A(\mem[234][0] ), .B(\mem[235][0] ), .S(n8466), .Z(n785)
         );
  MUX2_X1 U19735 ( .A(\mem[232][0] ), .B(\mem[233][0] ), .S(n8406), .Z(n786)
         );
  MUX2_X1 U19736 ( .A(n786), .B(n785), .S(n8282), .Z(n787) );
  MUX2_X1 U19737 ( .A(n787), .B(n784), .S(n8234), .Z(n788) );
  MUX2_X1 U19738 ( .A(\mem[230][0] ), .B(\mem[231][0] ), .S(n8421), .Z(n789)
         );
  MUX2_X1 U19739 ( .A(\mem[228][0] ), .B(\mem[229][0] ), .S(n8451), .Z(n790)
         );
  MUX2_X1 U19740 ( .A(n790), .B(n789), .S(n8327), .Z(n791) );
  MUX2_X1 U19741 ( .A(\mem[226][0] ), .B(\mem[227][0] ), .S(n8533), .Z(n792)
         );
  MUX2_X1 U19742 ( .A(\mem[224][0] ), .B(\mem[225][0] ), .S(n8463), .Z(n793)
         );
  MUX2_X1 U19743 ( .A(n793), .B(n792), .S(n8270), .Z(n794) );
  MUX2_X1 U19744 ( .A(n794), .B(n791), .S(n8234), .Z(n795) );
  MUX2_X1 U19745 ( .A(n795), .B(n788), .S(n8219), .Z(n796) );
  MUX2_X1 U19746 ( .A(n796), .B(n781), .S(n8195), .Z(n797) );
  MUX2_X1 U19747 ( .A(\mem[222][0] ), .B(\mem[223][0] ), .S(n8535), .Z(n798)
         );
  MUX2_X1 U19748 ( .A(\mem[220][0] ), .B(\mem[221][0] ), .S(n8378), .Z(n799)
         );
  MUX2_X1 U19749 ( .A(n799), .B(n798), .S(n8272), .Z(n800) );
  MUX2_X1 U19750 ( .A(\mem[218][0] ), .B(\mem[219][0] ), .S(n8377), .Z(n801)
         );
  MUX2_X1 U19751 ( .A(\mem[216][0] ), .B(\mem[217][0] ), .S(n8376), .Z(n802)
         );
  MUX2_X1 U19752 ( .A(n802), .B(n801), .S(n8280), .Z(n803) );
  MUX2_X1 U19753 ( .A(n803), .B(n800), .S(n8235), .Z(n804) );
  MUX2_X1 U19754 ( .A(\mem[214][0] ), .B(\mem[215][0] ), .S(n8375), .Z(n805)
         );
  MUX2_X1 U19755 ( .A(\mem[212][0] ), .B(\mem[213][0] ), .S(n8374), .Z(n806)
         );
  MUX2_X1 U19756 ( .A(n806), .B(n805), .S(n8279), .Z(n807) );
  MUX2_X1 U19757 ( .A(\mem[210][0] ), .B(\mem[211][0] ), .S(n8360), .Z(n808)
         );
  MUX2_X1 U19758 ( .A(\mem[208][0] ), .B(\mem[209][0] ), .S(n8361), .Z(n809)
         );
  MUX2_X1 U19759 ( .A(n809), .B(n808), .S(n8330), .Z(n810) );
  MUX2_X1 U19760 ( .A(n810), .B(n807), .S(n8235), .Z(n811) );
  MUX2_X1 U19761 ( .A(n811), .B(n804), .S(n8219), .Z(n812) );
  MUX2_X1 U19762 ( .A(\mem[206][0] ), .B(\mem[207][0] ), .S(n8538), .Z(n813)
         );
  MUX2_X1 U19763 ( .A(\mem[204][0] ), .B(\mem[205][0] ), .S(n8359), .Z(n814)
         );
  MUX2_X1 U19764 ( .A(n814), .B(n813), .S(n8278), .Z(n815) );
  MUX2_X1 U19765 ( .A(\mem[202][0] ), .B(\mem[203][0] ), .S(n8512), .Z(n816)
         );
  MUX2_X1 U19766 ( .A(\mem[200][0] ), .B(\mem[201][0] ), .S(n8432), .Z(n817)
         );
  MUX2_X1 U19767 ( .A(n817), .B(n816), .S(n8277), .Z(n818) );
  MUX2_X1 U19768 ( .A(n818), .B(n815), .S(n8235), .Z(n819) );
  MUX2_X1 U19769 ( .A(\mem[198][0] ), .B(\mem[199][0] ), .S(n8538), .Z(n820)
         );
  MUX2_X1 U19770 ( .A(\mem[196][0] ), .B(\mem[197][0] ), .S(n8359), .Z(n821)
         );
  MUX2_X1 U19771 ( .A(n821), .B(n820), .S(n8276), .Z(n822) );
  MUX2_X1 U19772 ( .A(\mem[194][0] ), .B(\mem[195][0] ), .S(n8360), .Z(n823)
         );
  MUX2_X1 U19773 ( .A(\mem[192][0] ), .B(\mem[193][0] ), .S(n8361), .Z(n824)
         );
  MUX2_X1 U19774 ( .A(n824), .B(n823), .S(n8275), .Z(n825) );
  MUX2_X1 U19775 ( .A(n825), .B(n822), .S(n8235), .Z(n826) );
  MUX2_X1 U19776 ( .A(n826), .B(n819), .S(n8197), .Z(n827) );
  MUX2_X1 U19777 ( .A(n827), .B(n812), .S(n8190), .Z(n828) );
  MUX2_X1 U19778 ( .A(n828), .B(n797), .S(n8181), .Z(n829) );
  MUX2_X1 U19779 ( .A(\mem[190][0] ), .B(\mem[191][0] ), .S(n8538), .Z(n830)
         );
  MUX2_X1 U19780 ( .A(\mem[188][0] ), .B(\mem[189][0] ), .S(n8359), .Z(n831)
         );
  MUX2_X1 U19781 ( .A(n831), .B(n830), .S(n8274), .Z(n832) );
  MUX2_X1 U19782 ( .A(\mem[186][0] ), .B(\mem[187][0] ), .S(n8360), .Z(n833)
         );
  MUX2_X1 U19783 ( .A(\mem[184][0] ), .B(\mem[185][0] ), .S(n8361), .Z(n834)
         );
  MUX2_X1 U19784 ( .A(n834), .B(n833), .S(n8273), .Z(n835) );
  MUX2_X1 U19785 ( .A(n835), .B(n832), .S(n8235), .Z(n836) );
  MUX2_X1 U19786 ( .A(\mem[182][0] ), .B(\mem[183][0] ), .S(n8382), .Z(n837)
         );
  MUX2_X1 U19787 ( .A(\mem[180][0] ), .B(\mem[181][0] ), .S(n8381), .Z(n838)
         );
  MUX2_X1 U19788 ( .A(n838), .B(n837), .S(n8266), .Z(n839) );
  MUX2_X1 U19789 ( .A(\mem[178][0] ), .B(\mem[179][0] ), .S(n8380), .Z(n840)
         );
  MUX2_X1 U19790 ( .A(\mem[176][0] ), .B(\mem[177][0] ), .S(n8379), .Z(n841)
         );
  MUX2_X1 U19791 ( .A(n841), .B(n840), .S(n8356), .Z(n842) );
  MUX2_X1 U19792 ( .A(n842), .B(n839), .S(n8235), .Z(n843) );
  MUX2_X1 U19793 ( .A(n843), .B(n836), .S(n8214), .Z(n844) );
  MUX2_X1 U19794 ( .A(\mem[174][0] ), .B(\mem[175][0] ), .S(n8359), .Z(n845)
         );
  MUX2_X1 U19795 ( .A(\mem[172][0] ), .B(\mem[173][0] ), .S(n8538), .Z(n846)
         );
  MUX2_X1 U19796 ( .A(n846), .B(n845), .S(n8308), .Z(n847) );
  MUX2_X1 U19797 ( .A(\mem[170][0] ), .B(\mem[171][0] ), .S(n8374), .Z(n848)
         );
  MUX2_X1 U19798 ( .A(\mem[168][0] ), .B(\mem[169][0] ), .S(n8370), .Z(n849)
         );
  MUX2_X1 U19799 ( .A(n849), .B(n848), .S(n8283), .Z(n850) );
  MUX2_X1 U19800 ( .A(n850), .B(n847), .S(n8235), .Z(n851) );
  MUX2_X1 U19801 ( .A(\mem[166][0] ), .B(\mem[167][0] ), .S(n8377), .Z(n852)
         );
  MUX2_X1 U19802 ( .A(\mem[164][0] ), .B(\mem[165][0] ), .S(n8455), .Z(n853)
         );
  MUX2_X1 U19803 ( .A(n853), .B(n852), .S(n8353), .Z(n854) );
  MUX2_X1 U19804 ( .A(\mem[162][0] ), .B(\mem[163][0] ), .S(n8389), .Z(n855)
         );
  MUX2_X1 U19805 ( .A(\mem[160][0] ), .B(\mem[161][0] ), .S(n8385), .Z(n856)
         );
  MUX2_X1 U19806 ( .A(n856), .B(n855), .S(n8354), .Z(n857) );
  MUX2_X1 U19807 ( .A(n857), .B(n854), .S(n8235), .Z(n858) );
  MUX2_X1 U19808 ( .A(n858), .B(n851), .S(n8210), .Z(n859) );
  MUX2_X1 U19809 ( .A(n859), .B(n844), .S(n8194), .Z(n860) );
  MUX2_X1 U19810 ( .A(\mem[158][0] ), .B(\mem[159][0] ), .S(n8393), .Z(n861)
         );
  MUX2_X1 U19811 ( .A(\mem[156][0] ), .B(\mem[157][0] ), .S(n8538), .Z(n862)
         );
  MUX2_X1 U19812 ( .A(n862), .B(n861), .S(n8268), .Z(n863) );
  MUX2_X1 U19813 ( .A(\mem[154][0] ), .B(\mem[155][0] ), .S(n8369), .Z(n864)
         );
  MUX2_X1 U19814 ( .A(\mem[152][0] ), .B(\mem[153][0] ), .S(n8532), .Z(n865)
         );
  MUX2_X1 U19815 ( .A(n865), .B(n864), .S(n8276), .Z(n866) );
  MUX2_X1 U19816 ( .A(n866), .B(n863), .S(n8235), .Z(n867) );
  MUX2_X1 U19817 ( .A(\mem[150][0] ), .B(\mem[151][0] ), .S(n8359), .Z(n868)
         );
  MUX2_X1 U19818 ( .A(\mem[148][0] ), .B(\mem[149][0] ), .S(n8380), .Z(n869)
         );
  MUX2_X1 U19819 ( .A(n869), .B(n868), .S(n8270), .Z(n870) );
  MUX2_X1 U19820 ( .A(\mem[146][0] ), .B(\mem[147][0] ), .S(n8359), .Z(n871)
         );
  MUX2_X1 U19821 ( .A(\mem[144][0] ), .B(\mem[145][0] ), .S(n8384), .Z(n872)
         );
  MUX2_X1 U19822 ( .A(n872), .B(n871), .S(n8274), .Z(n873) );
  MUX2_X1 U19823 ( .A(n873), .B(n870), .S(n8235), .Z(n874) );
  MUX2_X1 U19824 ( .A(n874), .B(n867), .S(n8205), .Z(n875) );
  MUX2_X1 U19825 ( .A(\mem[142][0] ), .B(\mem[143][0] ), .S(n8383), .Z(n876)
         );
  MUX2_X1 U19826 ( .A(\mem[140][0] ), .B(\mem[141][0] ), .S(n8441), .Z(n877)
         );
  MUX2_X1 U19827 ( .A(n877), .B(n876), .S(n8346), .Z(n878) );
  MUX2_X1 U19828 ( .A(\mem[138][0] ), .B(\mem[139][0] ), .S(n8417), .Z(n879)
         );
  MUX2_X1 U19829 ( .A(\mem[136][0] ), .B(\mem[137][0] ), .S(n8538), .Z(n880)
         );
  MUX2_X1 U19830 ( .A(n880), .B(n879), .S(n8325), .Z(n881) );
  MUX2_X1 U19831 ( .A(n881), .B(n878), .S(n8235), .Z(n882) );
  MUX2_X1 U19832 ( .A(\mem[134][0] ), .B(\mem[135][0] ), .S(n8359), .Z(n883)
         );
  MUX2_X1 U19833 ( .A(\mem[132][0] ), .B(\mem[133][0] ), .S(n8359), .Z(n884)
         );
  MUX2_X1 U19834 ( .A(n884), .B(n883), .S(n8272), .Z(n885) );
  MUX2_X1 U19835 ( .A(\mem[130][0] ), .B(\mem[131][0] ), .S(n8385), .Z(n886)
         );
  MUX2_X1 U19836 ( .A(\mem[128][0] ), .B(\mem[129][0] ), .S(n8417), .Z(n887)
         );
  MUX2_X1 U19837 ( .A(n887), .B(n886), .S(n8354), .Z(n888) );
  MUX2_X1 U19838 ( .A(n888), .B(n885), .S(n8235), .Z(n889) );
  MUX2_X1 U19839 ( .A(n889), .B(n882), .S(n8212), .Z(n890) );
  MUX2_X1 U19840 ( .A(n890), .B(n875), .S(n8195), .Z(n891) );
  MUX2_X1 U19841 ( .A(n891), .B(n860), .S(n8181), .Z(n892) );
  MUX2_X1 U19842 ( .A(n892), .B(n829), .S(n8179), .Z(n893) );
  MUX2_X1 U19843 ( .A(\mem[126][0] ), .B(\mem[127][0] ), .S(n8431), .Z(n894)
         );
  MUX2_X1 U19844 ( .A(\mem[124][0] ), .B(\mem[125][0] ), .S(n8416), .Z(n895)
         );
  MUX2_X1 U19845 ( .A(n895), .B(n894), .S(n8274), .Z(n896) );
  MUX2_X1 U19846 ( .A(\mem[122][0] ), .B(\mem[123][0] ), .S(n8399), .Z(n897)
         );
  MUX2_X1 U19847 ( .A(\mem[120][0] ), .B(\mem[121][0] ), .S(n8537), .Z(n898)
         );
  MUX2_X1 U19848 ( .A(n898), .B(n897), .S(n8320), .Z(n899) );
  MUX2_X1 U19849 ( .A(n899), .B(n896), .S(n8236), .Z(n900) );
  MUX2_X1 U19850 ( .A(\mem[118][0] ), .B(\mem[119][0] ), .S(n8414), .Z(n901)
         );
  MUX2_X1 U19851 ( .A(\mem[116][0] ), .B(\mem[117][0] ), .S(n8495), .Z(n902)
         );
  MUX2_X1 U19852 ( .A(n902), .B(n901), .S(n8317), .Z(n903) );
  MUX2_X1 U19853 ( .A(\mem[114][0] ), .B(\mem[115][0] ), .S(n8532), .Z(n904)
         );
  MUX2_X1 U19854 ( .A(\mem[112][0] ), .B(\mem[113][0] ), .S(n8384), .Z(n905)
         );
  MUX2_X1 U19855 ( .A(n905), .B(n904), .S(n8271), .Z(n906) );
  MUX2_X1 U19856 ( .A(n906), .B(n903), .S(n8236), .Z(n907) );
  MUX2_X1 U19857 ( .A(n907), .B(n900), .S(n8210), .Z(n908) );
  MUX2_X1 U19858 ( .A(\mem[110][0] ), .B(\mem[111][0] ), .S(n8400), .Z(n909)
         );
  MUX2_X1 U19859 ( .A(\mem[108][0] ), .B(\mem[109][0] ), .S(n8469), .Z(n910)
         );
  MUX2_X1 U19860 ( .A(n910), .B(n909), .S(n8281), .Z(n911) );
  MUX2_X1 U19861 ( .A(\mem[106][0] ), .B(\mem[107][0] ), .S(n8382), .Z(n912)
         );
  MUX2_X1 U19862 ( .A(\mem[104][0] ), .B(\mem[105][0] ), .S(n8381), .Z(n913)
         );
  MUX2_X1 U19863 ( .A(n913), .B(n912), .S(n8280), .Z(n914) );
  MUX2_X1 U19864 ( .A(n914), .B(n911), .S(n8236), .Z(n915) );
  MUX2_X1 U19865 ( .A(\mem[102][0] ), .B(\mem[103][0] ), .S(n8377), .Z(n916)
         );
  MUX2_X1 U19866 ( .A(\mem[100][0] ), .B(\mem[101][0] ), .S(n8376), .Z(n917)
         );
  MUX2_X1 U19867 ( .A(n917), .B(n916), .S(n8279), .Z(n918) );
  MUX2_X1 U19868 ( .A(\mem[98][0] ), .B(\mem[99][0] ), .S(n8375), .Z(n919) );
  MUX2_X1 U19869 ( .A(\mem[96][0] ), .B(\mem[97][0] ), .S(n8475), .Z(n920) );
  MUX2_X1 U19870 ( .A(n920), .B(n919), .S(n8289), .Z(n921) );
  MUX2_X1 U19871 ( .A(n921), .B(n918), .S(n8236), .Z(n922) );
  MUX2_X1 U19872 ( .A(n922), .B(n915), .S(n8200), .Z(n923) );
  MUX2_X1 U19873 ( .A(n923), .B(n908), .S(n8196), .Z(n924) );
  MUX2_X1 U19874 ( .A(\mem[94][0] ), .B(\mem[95][0] ), .S(n8422), .Z(n925) );
  MUX2_X1 U19875 ( .A(\mem[92][0] ), .B(\mem[93][0] ), .S(n8358), .Z(n926) );
  MUX2_X1 U19876 ( .A(n926), .B(n925), .S(n8335), .Z(n927) );
  MUX2_X1 U19877 ( .A(\mem[90][0] ), .B(\mem[91][0] ), .S(n8458), .Z(n928) );
  MUX2_X1 U19878 ( .A(\mem[88][0] ), .B(\mem[89][0] ), .S(n8517), .Z(n929) );
  MUX2_X1 U19879 ( .A(n929), .B(n928), .S(n8279), .Z(n930) );
  MUX2_X1 U19880 ( .A(n930), .B(n927), .S(n8236), .Z(n931) );
  MUX2_X1 U19881 ( .A(\mem[86][0] ), .B(\mem[87][0] ), .S(n8377), .Z(n932) );
  MUX2_X1 U19882 ( .A(\mem[84][0] ), .B(\mem[85][0] ), .S(n8487), .Z(n933) );
  MUX2_X1 U19883 ( .A(n933), .B(n932), .S(n8295), .Z(n934) );
  MUX2_X1 U19884 ( .A(\mem[82][0] ), .B(\mem[83][0] ), .S(n8430), .Z(n935) );
  MUX2_X1 U19885 ( .A(\mem[80][0] ), .B(\mem[81][0] ), .S(n8385), .Z(n936) );
  MUX2_X1 U19886 ( .A(n936), .B(n935), .S(n8293), .Z(n937) );
  MUX2_X1 U19887 ( .A(n937), .B(n934), .S(n8236), .Z(n938) );
  MUX2_X1 U19888 ( .A(n938), .B(n931), .S(n8199), .Z(n939) );
  MUX2_X1 U19889 ( .A(\mem[78][0] ), .B(\mem[79][0] ), .S(n8537), .Z(n940) );
  MUX2_X1 U19890 ( .A(\mem[76][0] ), .B(\mem[77][0] ), .S(n8380), .Z(n941) );
  MUX2_X1 U19891 ( .A(n941), .B(n940), .S(n8281), .Z(n942) );
  MUX2_X1 U19892 ( .A(\mem[74][0] ), .B(\mem[75][0] ), .S(n8384), .Z(n943) );
  MUX2_X1 U19893 ( .A(\mem[72][0] ), .B(\mem[73][0] ), .S(n8383), .Z(n944) );
  MUX2_X1 U19894 ( .A(n944), .B(n943), .S(n8284), .Z(n945) );
  MUX2_X1 U19895 ( .A(n945), .B(n942), .S(n8236), .Z(n946) );
  MUX2_X1 U19896 ( .A(\mem[70][0] ), .B(\mem[71][0] ), .S(n8413), .Z(n947) );
  MUX2_X1 U19897 ( .A(\mem[68][0] ), .B(\mem[69][0] ), .S(n8389), .Z(n948) );
  MUX2_X1 U19898 ( .A(n948), .B(n947), .S(n8334), .Z(n949) );
  MUX2_X1 U19899 ( .A(\mem[66][0] ), .B(\mem[67][0] ), .S(n8531), .Z(n950) );
  MUX2_X1 U19900 ( .A(\mem[64][0] ), .B(\mem[65][0] ), .S(n8455), .Z(n951) );
  MUX2_X1 U19901 ( .A(n951), .B(n950), .S(n8268), .Z(n952) );
  MUX2_X1 U19902 ( .A(n952), .B(n949), .S(n8236), .Z(n953) );
  MUX2_X1 U19903 ( .A(n953), .B(n946), .S(n8198), .Z(n954) );
  MUX2_X1 U19904 ( .A(n954), .B(n939), .S(n8196), .Z(n955) );
  MUX2_X1 U19905 ( .A(n955), .B(n924), .S(n8181), .Z(n956) );
  MUX2_X1 U19906 ( .A(\mem[62][0] ), .B(\mem[63][0] ), .S(n8527), .Z(n957) );
  MUX2_X1 U19907 ( .A(\mem[60][0] ), .B(\mem[61][0] ), .S(n8510), .Z(n958) );
  MUX2_X1 U19908 ( .A(n958), .B(n957), .S(n8270), .Z(n959) );
  MUX2_X1 U19909 ( .A(\mem[58][0] ), .B(\mem[59][0] ), .S(n8379), .Z(n960) );
  MUX2_X1 U19910 ( .A(\mem[56][0] ), .B(\mem[57][0] ), .S(n8378), .Z(n961) );
  MUX2_X1 U19911 ( .A(n961), .B(n960), .S(n8356), .Z(n962) );
  MUX2_X1 U19912 ( .A(n962), .B(n959), .S(n8236), .Z(n963) );
  MUX2_X1 U19913 ( .A(\mem[54][0] ), .B(\mem[55][0] ), .S(n8408), .Z(n964) );
  MUX2_X1 U19914 ( .A(\mem[52][0] ), .B(\mem[53][0] ), .S(n8517), .Z(n965) );
  MUX2_X1 U19915 ( .A(n965), .B(n964), .S(n8309), .Z(n966) );
  MUX2_X1 U19916 ( .A(\mem[50][0] ), .B(\mem[51][0] ), .S(n8399), .Z(n967) );
  MUX2_X1 U19917 ( .A(\mem[48][0] ), .B(\mem[49][0] ), .S(n8370), .Z(n968) );
  MUX2_X1 U19918 ( .A(n968), .B(n967), .S(n8348), .Z(n969) );
  MUX2_X1 U19919 ( .A(n969), .B(n966), .S(n8236), .Z(n970) );
  MUX2_X1 U19920 ( .A(n970), .B(n963), .S(n8206), .Z(n971) );
  MUX2_X1 U19921 ( .A(\mem[46][0] ), .B(\mem[47][0] ), .S(n8535), .Z(n972) );
  MUX2_X1 U19922 ( .A(\mem[44][0] ), .B(\mem[45][0] ), .S(n8525), .Z(n973) );
  MUX2_X1 U19923 ( .A(n973), .B(n972), .S(n8272), .Z(n974) );
  MUX2_X1 U19924 ( .A(\mem[42][0] ), .B(\mem[43][0] ), .S(n8360), .Z(n975) );
  MUX2_X1 U19925 ( .A(\mem[40][0] ), .B(\mem[41][0] ), .S(n8522), .Z(n976) );
  MUX2_X1 U19926 ( .A(n976), .B(n975), .S(n8266), .Z(n977) );
  MUX2_X1 U19927 ( .A(n977), .B(n974), .S(n8236), .Z(n978) );
  MUX2_X1 U19928 ( .A(\mem[38][0] ), .B(\mem[39][0] ), .S(n8469), .Z(n979) );
  MUX2_X1 U19929 ( .A(\mem[36][0] ), .B(\mem[37][0] ), .S(n8404), .Z(n980) );
  MUX2_X1 U19930 ( .A(n980), .B(n979), .S(n8273), .Z(n981) );
  MUX2_X1 U19931 ( .A(\mem[34][0] ), .B(\mem[35][0] ), .S(n8382), .Z(n982) );
  MUX2_X1 U19932 ( .A(\mem[32][0] ), .B(\mem[33][0] ), .S(n8381), .Z(n983) );
  MUX2_X1 U19933 ( .A(n983), .B(n982), .S(n8267), .Z(n984) );
  MUX2_X1 U19934 ( .A(n984), .B(n981), .S(n8236), .Z(n985) );
  MUX2_X1 U19935 ( .A(n985), .B(n978), .S(n8219), .Z(n986) );
  MUX2_X1 U19936 ( .A(n986), .B(n971), .S(n8192), .Z(n987) );
  MUX2_X1 U19937 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n8377), .Z(n988) );
  MUX2_X1 U19938 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n8376), .Z(n989) );
  MUX2_X1 U19939 ( .A(n989), .B(n988), .S(n8286), .Z(n990) );
  MUX2_X1 U19940 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n8457), .Z(n991) );
  MUX2_X1 U19941 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n8535), .Z(n992) );
  MUX2_X1 U19942 ( .A(n992), .B(n991), .S(n8269), .Z(n993) );
  MUX2_X1 U19943 ( .A(n993), .B(n990), .S(n8237), .Z(n994) );
  MUX2_X1 U19944 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n8361), .Z(n995) );
  MUX2_X1 U19945 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n8486), .Z(n996) );
  MUX2_X1 U19946 ( .A(n996), .B(n995), .S(n8356), .Z(n997) );
  MUX2_X1 U19947 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n8429), .Z(n998) );
  MUX2_X1 U19948 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n8360), .Z(n999) );
  MUX2_X1 U19949 ( .A(n999), .B(n998), .S(n8266), .Z(n1000) );
  MUX2_X1 U19950 ( .A(n1000), .B(n997), .S(n8237), .Z(n1001) );
  MUX2_X1 U19951 ( .A(n1001), .B(n994), .S(n8214), .Z(n1002) );
  MUX2_X1 U19952 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n8462), .Z(n1003) );
  MUX2_X1 U19953 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n8446), .Z(n1004) );
  MUX2_X1 U19954 ( .A(n1004), .B(n1003), .S(n8267), .Z(n1005) );
  MUX2_X1 U19955 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n8421), .Z(n1006) );
  MUX2_X1 U19956 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n8385), .Z(n1007) );
  MUX2_X1 U19957 ( .A(n1007), .B(n1006), .S(n8267), .Z(n1008) );
  MUX2_X1 U19958 ( .A(n1008), .B(n1005), .S(n8237), .Z(n1009) );
  MUX2_X1 U19959 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n8379), .Z(n1010) );
  MUX2_X1 U19960 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n8379), .Z(n1011) );
  MUX2_X1 U19961 ( .A(n1011), .B(n1010), .S(n8286), .Z(n1012) );
  MUX2_X1 U19962 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n8378), .Z(n1013) );
  MUX2_X1 U19963 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n8412), .Z(n1014) );
  MUX2_X1 U19964 ( .A(n1014), .B(n1013), .S(n8353), .Z(n1015) );
  MUX2_X1 U19965 ( .A(n1015), .B(n1012), .S(n8237), .Z(n1016) );
  MUX2_X1 U19966 ( .A(n1016), .B(n1009), .S(n8219), .Z(n1017) );
  MUX2_X1 U19967 ( .A(n1017), .B(n1002), .S(n8189), .Z(n1018) );
  MUX2_X1 U19968 ( .A(n1018), .B(n987), .S(n8181), .Z(n1019) );
  MUX2_X1 U19969 ( .A(n1019), .B(n956), .S(n8179), .Z(n1020) );
  MUX2_X1 U19970 ( .A(n1020), .B(n893), .S(n8177), .Z(n1021) );
  MUX2_X1 U19971 ( .A(n1021), .B(n766), .S(N26), .Z(n1022) );
  MUX2_X1 U19972 ( .A(n1022), .B(n511), .S(N27), .Z(N35) );
  MUX2_X1 U19973 ( .A(\mem[1022][1] ), .B(\mem[1023][1] ), .S(n8392), .Z(n1023) );
  MUX2_X1 U19974 ( .A(\mem[1020][1] ), .B(\mem[1021][1] ), .S(n8536), .Z(n1024) );
  MUX2_X1 U19975 ( .A(n1024), .B(n1023), .S(n8315), .Z(n1025) );
  MUX2_X1 U19976 ( .A(\mem[1018][1] ), .B(\mem[1019][1] ), .S(n8454), .Z(n1026) );
  MUX2_X1 U19977 ( .A(\mem[1016][1] ), .B(\mem[1017][1] ), .S(n8526), .Z(n1027) );
  MUX2_X1 U19978 ( .A(n1027), .B(n1026), .S(n8270), .Z(n1028) );
  MUX2_X1 U19979 ( .A(n1028), .B(n1025), .S(n8237), .Z(n1029) );
  MUX2_X1 U19980 ( .A(\mem[1014][1] ), .B(\mem[1015][1] ), .S(n8503), .Z(n1030) );
  MUX2_X1 U19981 ( .A(\mem[1012][1] ), .B(\mem[1013][1] ), .S(n8385), .Z(n1031) );
  MUX2_X1 U19982 ( .A(n1031), .B(n1030), .S(n8268), .Z(n1032) );
  MUX2_X1 U19983 ( .A(\mem[1010][1] ), .B(\mem[1011][1] ), .S(n8384), .Z(n1033) );
  MUX2_X1 U19984 ( .A(\mem[1008][1] ), .B(\mem[1009][1] ), .S(n8383), .Z(n1034) );
  MUX2_X1 U19985 ( .A(n1034), .B(n1033), .S(n8275), .Z(n1035) );
  MUX2_X1 U19986 ( .A(n1035), .B(n1032), .S(n8237), .Z(n1036) );
  MUX2_X1 U19987 ( .A(n1036), .B(n1029), .S(n8197), .Z(n1037) );
  MUX2_X1 U19988 ( .A(\mem[1006][1] ), .B(\mem[1007][1] ), .S(n8374), .Z(n1038) );
  MUX2_X1 U19989 ( .A(\mem[1004][1] ), .B(\mem[1005][1] ), .S(n8371), .Z(n1039) );
  MUX2_X1 U19990 ( .A(n1039), .B(n1038), .S(n8276), .Z(n1040) );
  MUX2_X1 U19991 ( .A(\mem[1002][1] ), .B(\mem[1003][1] ), .S(n8378), .Z(n1041) );
  MUX2_X1 U19992 ( .A(\mem[1000][1] ), .B(\mem[1001][1] ), .S(n8474), .Z(n1042) );
  MUX2_X1 U19993 ( .A(n1042), .B(n1041), .S(n8275), .Z(n1043) );
  MUX2_X1 U19994 ( .A(n1043), .B(n1040), .S(n8237), .Z(n1044) );
  MUX2_X1 U19995 ( .A(\mem[998][1] ), .B(\mem[999][1] ), .S(n8454), .Z(n1045)
         );
  MUX2_X1 U19996 ( .A(\mem[996][1] ), .B(\mem[997][1] ), .S(n8359), .Z(n1046)
         );
  MUX2_X1 U19997 ( .A(n1046), .B(n1045), .S(n8274), .Z(n1047) );
  MUX2_X1 U19998 ( .A(\mem[994][1] ), .B(\mem[995][1] ), .S(n8362), .Z(n1048)
         );
  MUX2_X1 U19999 ( .A(\mem[992][1] ), .B(\mem[993][1] ), .S(n8468), .Z(n1049)
         );
  MUX2_X1 U20000 ( .A(n1049), .B(n1048), .S(n8273), .Z(n1050) );
  MUX2_X1 U20001 ( .A(n1050), .B(n1047), .S(n8237), .Z(n1051) );
  MUX2_X1 U20002 ( .A(n1051), .B(n1044), .S(n8199), .Z(n1052) );
  MUX2_X1 U20003 ( .A(n1052), .B(n1037), .S(n8193), .Z(n1053) );
  MUX2_X1 U20004 ( .A(\mem[990][1] ), .B(\mem[991][1] ), .S(n8397), .Z(n1054)
         );
  MUX2_X1 U20005 ( .A(\mem[988][1] ), .B(\mem[989][1] ), .S(n8382), .Z(n1055)
         );
  MUX2_X1 U20006 ( .A(n1055), .B(n1054), .S(n8268), .Z(n1056) );
  MUX2_X1 U20007 ( .A(\mem[986][1] ), .B(\mem[987][1] ), .S(n8381), .Z(n1057)
         );
  MUX2_X1 U20008 ( .A(\mem[984][1] ), .B(\mem[985][1] ), .S(n8380), .Z(n1058)
         );
  MUX2_X1 U20009 ( .A(n1058), .B(n1057), .S(n8339), .Z(n1059) );
  MUX2_X1 U20010 ( .A(n1059), .B(n1056), .S(n8237), .Z(n1060) );
  MUX2_X1 U20011 ( .A(\mem[982][1] ), .B(\mem[983][1] ), .S(n8357), .Z(n1061)
         );
  MUX2_X1 U20012 ( .A(\mem[980][1] ), .B(\mem[981][1] ), .S(n8450), .Z(n1062)
         );
  MUX2_X1 U20013 ( .A(n1062), .B(n1061), .S(n8340), .Z(n1063) );
  MUX2_X1 U20014 ( .A(\mem[978][1] ), .B(\mem[979][1] ), .S(n8461), .Z(n1064)
         );
  MUX2_X1 U20015 ( .A(\mem[976][1] ), .B(\mem[977][1] ), .S(n8396), .Z(n1065)
         );
  MUX2_X1 U20016 ( .A(n1065), .B(n1064), .S(n8328), .Z(n1066) );
  MUX2_X1 U20017 ( .A(n1066), .B(n1063), .S(n8237), .Z(n1067) );
  MUX2_X1 U20018 ( .A(n1067), .B(n1060), .S(n8206), .Z(n1068) );
  MUX2_X1 U20019 ( .A(\mem[974][1] ), .B(\mem[975][1] ), .S(n8382), .Z(n1069)
         );
  MUX2_X1 U20020 ( .A(\mem[972][1] ), .B(\mem[973][1] ), .S(n8381), .Z(n1070)
         );
  MUX2_X1 U20021 ( .A(n1070), .B(n1069), .S(n8272), .Z(n1071) );
  MUX2_X1 U20022 ( .A(\mem[970][1] ), .B(\mem[971][1] ), .S(n8380), .Z(n1072)
         );
  MUX2_X1 U20023 ( .A(\mem[968][1] ), .B(\mem[969][1] ), .S(n8391), .Z(n1073)
         );
  MUX2_X1 U20024 ( .A(n1073), .B(n1072), .S(n8271), .Z(n1074) );
  MUX2_X1 U20025 ( .A(n1074), .B(n1071), .S(n8237), .Z(n1075) );
  MUX2_X1 U20026 ( .A(\mem[966][1] ), .B(\mem[967][1] ), .S(n8535), .Z(n1076)
         );
  MUX2_X1 U20027 ( .A(\mem[964][1] ), .B(\mem[965][1] ), .S(n8453), .Z(n1077)
         );
  MUX2_X1 U20028 ( .A(n1077), .B(n1076), .S(n8342), .Z(n1078) );
  MUX2_X1 U20029 ( .A(\mem[962][1] ), .B(\mem[963][1] ), .S(n8525), .Z(n1079)
         );
  MUX2_X1 U20030 ( .A(\mem[960][1] ), .B(\mem[961][1] ), .S(n8502), .Z(n1080)
         );
  MUX2_X1 U20031 ( .A(n1080), .B(n1079), .S(n8298), .Z(n1081) );
  MUX2_X1 U20032 ( .A(n1081), .B(n1078), .S(n8237), .Z(n1082) );
  MUX2_X1 U20033 ( .A(n1082), .B(n1075), .S(n8205), .Z(n1083) );
  MUX2_X1 U20034 ( .A(n1083), .B(n1068), .S(n8191), .Z(n1084) );
  MUX2_X1 U20035 ( .A(n1084), .B(n1053), .S(n8181), .Z(n1085) );
  MUX2_X1 U20036 ( .A(\mem[958][1] ), .B(\mem[959][1] ), .S(n8376), .Z(n1086)
         );
  MUX2_X1 U20037 ( .A(\mem[956][1] ), .B(\mem[957][1] ), .S(n8450), .Z(n1087)
         );
  MUX2_X1 U20038 ( .A(n1087), .B(n1086), .S(n8283), .Z(n1088) );
  MUX2_X1 U20039 ( .A(\mem[954][1] ), .B(\mem[955][1] ), .S(n8377), .Z(n1089)
         );
  MUX2_X1 U20040 ( .A(\mem[952][1] ), .B(\mem[953][1] ), .S(n8453), .Z(n1090)
         );
  MUX2_X1 U20041 ( .A(n1090), .B(n1089), .S(n8320), .Z(n1091) );
  MUX2_X1 U20042 ( .A(n1091), .B(n1088), .S(n8238), .Z(n1092) );
  MUX2_X1 U20043 ( .A(\mem[950][1] ), .B(\mem[951][1] ), .S(n8476), .Z(n1093)
         );
  MUX2_X1 U20044 ( .A(\mem[948][1] ), .B(\mem[949][1] ), .S(n8474), .Z(n1094)
         );
  MUX2_X1 U20045 ( .A(n1094), .B(n1093), .S(n8282), .Z(n1095) );
  MUX2_X1 U20046 ( .A(\mem[946][1] ), .B(\mem[947][1] ), .S(n8410), .Z(n1096)
         );
  MUX2_X1 U20047 ( .A(\mem[944][1] ), .B(\mem[945][1] ), .S(n8428), .Z(n1097)
         );
  MUX2_X1 U20048 ( .A(n1097), .B(n1096), .S(n8352), .Z(n1098) );
  MUX2_X1 U20049 ( .A(n1098), .B(n1095), .S(n8238), .Z(n1099) );
  MUX2_X1 U20050 ( .A(n1099), .B(n1092), .S(n8197), .Z(n1100) );
  MUX2_X1 U20051 ( .A(\mem[942][1] ), .B(\mem[943][1] ), .S(n8533), .Z(n1101)
         );
  MUX2_X1 U20052 ( .A(\mem[940][1] ), .B(\mem[941][1] ), .S(n8372), .Z(n1102)
         );
  MUX2_X1 U20053 ( .A(n1102), .B(n1101), .S(n8336), .Z(n1103) );
  MUX2_X1 U20054 ( .A(\mem[938][1] ), .B(\mem[939][1] ), .S(n8465), .Z(n1104)
         );
  MUX2_X1 U20055 ( .A(\mem[936][1] ), .B(\mem[937][1] ), .S(n8416), .Z(n1105)
         );
  MUX2_X1 U20056 ( .A(n1105), .B(n1104), .S(n8305), .Z(n1106) );
  MUX2_X1 U20057 ( .A(n1106), .B(n1103), .S(n8238), .Z(n1107) );
  MUX2_X1 U20058 ( .A(\mem[934][1] ), .B(\mem[935][1] ), .S(n8374), .Z(n1108)
         );
  MUX2_X1 U20059 ( .A(\mem[932][1] ), .B(\mem[933][1] ), .S(n8538), .Z(n1109)
         );
  MUX2_X1 U20060 ( .A(n1109), .B(n1108), .S(n8281), .Z(n1110) );
  MUX2_X1 U20061 ( .A(\mem[930][1] ), .B(\mem[931][1] ), .S(n8359), .Z(n1111)
         );
  MUX2_X1 U20062 ( .A(\mem[928][1] ), .B(\mem[929][1] ), .S(n8360), .Z(n1112)
         );
  MUX2_X1 U20063 ( .A(n1112), .B(n1111), .S(n8280), .Z(n1113) );
  MUX2_X1 U20064 ( .A(n1113), .B(n1110), .S(n8238), .Z(n1114) );
  MUX2_X1 U20065 ( .A(n1114), .B(n1107), .S(N21), .Z(n1115) );
  MUX2_X1 U20066 ( .A(n1115), .B(n1100), .S(n8189), .Z(n1116) );
  MUX2_X1 U20067 ( .A(\mem[926][1] ), .B(\mem[927][1] ), .S(n8419), .Z(n1117)
         );
  MUX2_X1 U20068 ( .A(\mem[924][1] ), .B(\mem[925][1] ), .S(n8358), .Z(n1118)
         );
  MUX2_X1 U20069 ( .A(n1118), .B(n1117), .S(n8279), .Z(n1119) );
  MUX2_X1 U20070 ( .A(\mem[922][1] ), .B(\mem[923][1] ), .S(n8361), .Z(n1120)
         );
  MUX2_X1 U20071 ( .A(\mem[920][1] ), .B(\mem[921][1] ), .S(n8439), .Z(n1121)
         );
  MUX2_X1 U20072 ( .A(n1121), .B(n1120), .S(n8338), .Z(n1122) );
  MUX2_X1 U20073 ( .A(n1122), .B(n1119), .S(n8238), .Z(n1123) );
  MUX2_X1 U20074 ( .A(\mem[918][1] ), .B(\mem[919][1] ), .S(n8372), .Z(n1124)
         );
  MUX2_X1 U20075 ( .A(\mem[916][1] ), .B(\mem[917][1] ), .S(n8474), .Z(n1125)
         );
  MUX2_X1 U20076 ( .A(n1125), .B(n1124), .S(n8278), .Z(n1126) );
  MUX2_X1 U20077 ( .A(\mem[914][1] ), .B(\mem[915][1] ), .S(n8366), .Z(n1127)
         );
  MUX2_X1 U20078 ( .A(\mem[912][1] ), .B(\mem[913][1] ), .S(n8453), .Z(n1128)
         );
  MUX2_X1 U20079 ( .A(n1128), .B(n1127), .S(n8277), .Z(n1129) );
  MUX2_X1 U20080 ( .A(n1129), .B(n1126), .S(n8238), .Z(n1130) );
  MUX2_X1 U20081 ( .A(n1130), .B(n1123), .S(n8202), .Z(n1131) );
  MUX2_X1 U20082 ( .A(\mem[910][1] ), .B(\mem[911][1] ), .S(n8374), .Z(n1132)
         );
  MUX2_X1 U20083 ( .A(\mem[908][1] ), .B(\mem[909][1] ), .S(n8539), .Z(n1133)
         );
  MUX2_X1 U20084 ( .A(n1133), .B(n1132), .S(n8279), .Z(n1134) );
  MUX2_X1 U20085 ( .A(\mem[906][1] ), .B(\mem[907][1] ), .S(n8373), .Z(n1135)
         );
  MUX2_X1 U20086 ( .A(\mem[904][1] ), .B(\mem[905][1] ), .S(n8465), .Z(n1136)
         );
  MUX2_X1 U20087 ( .A(n1136), .B(n1135), .S(n8294), .Z(n1137) );
  MUX2_X1 U20088 ( .A(n1137), .B(n1134), .S(n8238), .Z(n1138) );
  MUX2_X1 U20089 ( .A(\mem[902][1] ), .B(\mem[903][1] ), .S(n8457), .Z(n1139)
         );
  MUX2_X1 U20090 ( .A(\mem[900][1] ), .B(\mem[901][1] ), .S(n8373), .Z(n1140)
         );
  MUX2_X1 U20091 ( .A(n1140), .B(n1139), .S(n8309), .Z(n1141) );
  MUX2_X1 U20092 ( .A(\mem[898][1] ), .B(\mem[899][1] ), .S(n8526), .Z(n1142)
         );
  MUX2_X1 U20093 ( .A(\mem[896][1] ), .B(\mem[897][1] ), .S(n8466), .Z(n1143)
         );
  MUX2_X1 U20094 ( .A(n1143), .B(n1142), .S(n8274), .Z(n1144) );
  MUX2_X1 U20095 ( .A(n1144), .B(n1141), .S(n8238), .Z(n1145) );
  MUX2_X1 U20096 ( .A(n1145), .B(n1138), .S(n8219), .Z(n1146) );
  MUX2_X1 U20097 ( .A(n1146), .B(n1131), .S(n8186), .Z(n1147) );
  MUX2_X1 U20098 ( .A(n1147), .B(n1116), .S(n8181), .Z(n1148) );
  MUX2_X1 U20099 ( .A(n1148), .B(n1085), .S(n8179), .Z(n1149) );
  MUX2_X1 U20100 ( .A(\mem[894][1] ), .B(\mem[895][1] ), .S(n8369), .Z(n1150)
         );
  MUX2_X1 U20101 ( .A(\mem[892][1] ), .B(\mem[893][1] ), .S(n8409), .Z(n1151)
         );
  MUX2_X1 U20102 ( .A(n1151), .B(n1150), .S(n8273), .Z(n1152) );
  MUX2_X1 U20103 ( .A(\mem[890][1] ), .B(\mem[891][1] ), .S(n8539), .Z(n1153)
         );
  MUX2_X1 U20104 ( .A(\mem[888][1] ), .B(\mem[889][1] ), .S(n8365), .Z(n1154)
         );
  MUX2_X1 U20105 ( .A(n1154), .B(n1153), .S(n8343), .Z(n1155) );
  MUX2_X1 U20106 ( .A(n1155), .B(n1152), .S(n8238), .Z(n1156) );
  MUX2_X1 U20107 ( .A(\mem[886][1] ), .B(\mem[887][1] ), .S(n8394), .Z(n1157)
         );
  MUX2_X1 U20108 ( .A(\mem[884][1] ), .B(\mem[885][1] ), .S(n8527), .Z(n1158)
         );
  MUX2_X1 U20109 ( .A(n1158), .B(n1157), .S(n8268), .Z(n1159) );
  MUX2_X1 U20110 ( .A(\mem[882][1] ), .B(\mem[883][1] ), .S(n8457), .Z(n1160)
         );
  MUX2_X1 U20111 ( .A(\mem[880][1] ), .B(\mem[881][1] ), .S(n8529), .Z(n1161)
         );
  MUX2_X1 U20112 ( .A(n1161), .B(n1160), .S(n8270), .Z(n1162) );
  MUX2_X1 U20113 ( .A(n1162), .B(n1159), .S(n8238), .Z(n1163) );
  MUX2_X1 U20114 ( .A(n1163), .B(n1156), .S(n8200), .Z(n1164) );
  MUX2_X1 U20115 ( .A(\mem[878][1] ), .B(\mem[879][1] ), .S(n8382), .Z(n1165)
         );
  MUX2_X1 U20116 ( .A(\mem[876][1] ), .B(\mem[877][1] ), .S(n8381), .Z(n1166)
         );
  MUX2_X1 U20117 ( .A(n1166), .B(n1165), .S(n8356), .Z(n1167) );
  MUX2_X1 U20118 ( .A(\mem[874][1] ), .B(\mem[875][1] ), .S(n8380), .Z(n1168)
         );
  MUX2_X1 U20119 ( .A(\mem[872][1] ), .B(\mem[873][1] ), .S(n8379), .Z(n1169)
         );
  MUX2_X1 U20120 ( .A(n1169), .B(n1168), .S(N19), .Z(n1170) );
  MUX2_X1 U20121 ( .A(n1170), .B(n1167), .S(n8238), .Z(n1171) );
  MUX2_X1 U20122 ( .A(\mem[870][1] ), .B(\mem[871][1] ), .S(n8378), .Z(n1172)
         );
  MUX2_X1 U20123 ( .A(\mem[868][1] ), .B(\mem[869][1] ), .S(n8377), .Z(n1173)
         );
  MUX2_X1 U20124 ( .A(n1173), .B(n1172), .S(n8308), .Z(n1174) );
  MUX2_X1 U20125 ( .A(\mem[866][1] ), .B(\mem[867][1] ), .S(n8376), .Z(n1175)
         );
  MUX2_X1 U20126 ( .A(\mem[864][1] ), .B(\mem[865][1] ), .S(n8375), .Z(n1176)
         );
  MUX2_X1 U20127 ( .A(n1176), .B(n1175), .S(n8347), .Z(n1177) );
  MUX2_X1 U20128 ( .A(n1177), .B(n1174), .S(n8238), .Z(n1178) );
  MUX2_X1 U20129 ( .A(n1178), .B(n1171), .S(n8199), .Z(n1179) );
  MUX2_X1 U20130 ( .A(n1179), .B(n1164), .S(n8187), .Z(n1180) );
  MUX2_X1 U20131 ( .A(\mem[862][1] ), .B(\mem[863][1] ), .S(n8368), .Z(n1181)
         );
  MUX2_X1 U20132 ( .A(\mem[860][1] ), .B(\mem[861][1] ), .S(n8415), .Z(n1182)
         );
  MUX2_X1 U20133 ( .A(n1182), .B(n1181), .S(n8267), .Z(n1183) );
  MUX2_X1 U20134 ( .A(\mem[858][1] ), .B(\mem[859][1] ), .S(n8497), .Z(n1184)
         );
  MUX2_X1 U20135 ( .A(\mem[856][1] ), .B(\mem[857][1] ), .S(n8417), .Z(n1185)
         );
  MUX2_X1 U20136 ( .A(n1185), .B(n1184), .S(n8276), .Z(n1186) );
  MUX2_X1 U20137 ( .A(n1186), .B(n1183), .S(n8239), .Z(n1187) );
  MUX2_X1 U20138 ( .A(\mem[854][1] ), .B(\mem[855][1] ), .S(n8358), .Z(n1188)
         );
  MUX2_X1 U20139 ( .A(\mem[852][1] ), .B(\mem[853][1] ), .S(n8367), .Z(n1189)
         );
  MUX2_X1 U20140 ( .A(n1189), .B(n1188), .S(n8275), .Z(n1190) );
  MUX2_X1 U20141 ( .A(\mem[850][1] ), .B(\mem[851][1] ), .S(n8513), .Z(n1191)
         );
  MUX2_X1 U20142 ( .A(\mem[848][1] ), .B(\mem[849][1] ), .S(n8531), .Z(n1192)
         );
  MUX2_X1 U20143 ( .A(n1192), .B(n1191), .S(n8274), .Z(n1193) );
  MUX2_X1 U20144 ( .A(n1193), .B(n1190), .S(n8239), .Z(n1194) );
  MUX2_X1 U20145 ( .A(n1194), .B(n1187), .S(n8198), .Z(n1195) );
  MUX2_X1 U20146 ( .A(\mem[846][1] ), .B(\mem[847][1] ), .S(n8385), .Z(n1196)
         );
  MUX2_X1 U20147 ( .A(\mem[844][1] ), .B(\mem[845][1] ), .S(n8372), .Z(n1197)
         );
  MUX2_X1 U20148 ( .A(n1197), .B(n1196), .S(n8273), .Z(n1198) );
  MUX2_X1 U20149 ( .A(\mem[842][1] ), .B(\mem[843][1] ), .S(n8468), .Z(n1199)
         );
  MUX2_X1 U20150 ( .A(\mem[840][1] ), .B(\mem[841][1] ), .S(n8415), .Z(n1200)
         );
  MUX2_X1 U20151 ( .A(n1200), .B(n1199), .S(n8273), .Z(n1201) );
  MUX2_X1 U20152 ( .A(n1201), .B(n1198), .S(n8239), .Z(n1202) );
  MUX2_X1 U20153 ( .A(\mem[838][1] ), .B(\mem[839][1] ), .S(n8467), .Z(n1203)
         );
  MUX2_X1 U20154 ( .A(\mem[836][1] ), .B(\mem[837][1] ), .S(n8379), .Z(n1204)
         );
  MUX2_X1 U20155 ( .A(n1204), .B(n1203), .S(n8351), .Z(n1205) );
  MUX2_X1 U20156 ( .A(\mem[834][1] ), .B(\mem[835][1] ), .S(n8378), .Z(n1206)
         );
  MUX2_X1 U20157 ( .A(\mem[832][1] ), .B(\mem[833][1] ), .S(n8411), .Z(n1207)
         );
  MUX2_X1 U20158 ( .A(n1207), .B(n1206), .S(n8319), .Z(n1208) );
  MUX2_X1 U20159 ( .A(n1208), .B(n1205), .S(n8239), .Z(n1209) );
  MUX2_X1 U20160 ( .A(n1209), .B(n1202), .S(n8200), .Z(n1210) );
  MUX2_X1 U20161 ( .A(n1210), .B(n1195), .S(n8188), .Z(n1211) );
  MUX2_X1 U20162 ( .A(n1211), .B(n1180), .S(n8181), .Z(n1212) );
  MUX2_X1 U20163 ( .A(\mem[830][1] ), .B(\mem[831][1] ), .S(n8455), .Z(n1213)
         );
  MUX2_X1 U20164 ( .A(\mem[828][1] ), .B(\mem[829][1] ), .S(n8445), .Z(n1214)
         );
  MUX2_X1 U20165 ( .A(n1214), .B(n1213), .S(n8272), .Z(n1215) );
  MUX2_X1 U20166 ( .A(\mem[826][1] ), .B(\mem[827][1] ), .S(n8538), .Z(n1216)
         );
  MUX2_X1 U20167 ( .A(\mem[824][1] ), .B(\mem[825][1] ), .S(n8359), .Z(n1217)
         );
  MUX2_X1 U20168 ( .A(n1217), .B(n1216), .S(n8271), .Z(n1218) );
  MUX2_X1 U20169 ( .A(n1218), .B(n1215), .S(n8239), .Z(n1219) );
  MUX2_X1 U20170 ( .A(\mem[822][1] ), .B(\mem[823][1] ), .S(n8360), .Z(n1220)
         );
  MUX2_X1 U20171 ( .A(\mem[820][1] ), .B(\mem[821][1] ), .S(n8418), .Z(n1221)
         );
  MUX2_X1 U20172 ( .A(n1221), .B(n1220), .S(n8281), .Z(n1222) );
  MUX2_X1 U20173 ( .A(\mem[818][1] ), .B(\mem[819][1] ), .S(n8358), .Z(n1223)
         );
  MUX2_X1 U20174 ( .A(\mem[816][1] ), .B(\mem[817][1] ), .S(n8361), .Z(n1224)
         );
  MUX2_X1 U20175 ( .A(n1224), .B(n1223), .S(n8280), .Z(n1225) );
  MUX2_X1 U20176 ( .A(n1225), .B(n1222), .S(n8239), .Z(n1226) );
  MUX2_X1 U20177 ( .A(n1226), .B(n1219), .S(n8210), .Z(n1227) );
  MUX2_X1 U20178 ( .A(\mem[814][1] ), .B(\mem[815][1] ), .S(N18), .Z(n1228) );
  MUX2_X1 U20179 ( .A(\mem[812][1] ), .B(\mem[813][1] ), .S(n8358), .Z(n1229)
         );
  MUX2_X1 U20180 ( .A(n1229), .B(n1228), .S(n8269), .Z(n1230) );
  MUX2_X1 U20181 ( .A(\mem[810][1] ), .B(\mem[811][1] ), .S(n8495), .Z(n1231)
         );
  MUX2_X1 U20182 ( .A(\mem[808][1] ), .B(\mem[809][1] ), .S(n8480), .Z(n1232)
         );
  MUX2_X1 U20183 ( .A(n1232), .B(n1231), .S(n8269), .Z(n1233) );
  MUX2_X1 U20184 ( .A(n1233), .B(n1230), .S(n8239), .Z(n1234) );
  MUX2_X1 U20185 ( .A(\mem[806][1] ), .B(\mem[807][1] ), .S(n8461), .Z(n1235)
         );
  MUX2_X1 U20186 ( .A(\mem[804][1] ), .B(\mem[805][1] ), .S(n8414), .Z(n1236)
         );
  MUX2_X1 U20187 ( .A(n1236), .B(n1235), .S(n8285), .Z(n1237) );
  MUX2_X1 U20188 ( .A(\mem[802][1] ), .B(\mem[803][1] ), .S(n8528), .Z(n1238)
         );
  MUX2_X1 U20189 ( .A(\mem[800][1] ), .B(\mem[801][1] ), .S(n8382), .Z(n1239)
         );
  MUX2_X1 U20190 ( .A(n1239), .B(n1238), .S(n8284), .Z(n1240) );
  MUX2_X1 U20191 ( .A(n1240), .B(n1237), .S(n8239), .Z(n1241) );
  MUX2_X1 U20192 ( .A(n1241), .B(n1234), .S(N21), .Z(n1242) );
  MUX2_X1 U20193 ( .A(n1242), .B(n1227), .S(n8192), .Z(n1243) );
  MUX2_X1 U20194 ( .A(\mem[798][1] ), .B(\mem[799][1] ), .S(n8381), .Z(n1244)
         );
  MUX2_X1 U20195 ( .A(\mem[796][1] ), .B(\mem[797][1] ), .S(n8380), .Z(n1245)
         );
  MUX2_X1 U20196 ( .A(n1245), .B(n1244), .S(n8351), .Z(n1246) );
  MUX2_X1 U20197 ( .A(\mem[794][1] ), .B(\mem[795][1] ), .S(n8379), .Z(n1247)
         );
  MUX2_X1 U20198 ( .A(\mem[792][1] ), .B(\mem[793][1] ), .S(n8378), .Z(n1248)
         );
  MUX2_X1 U20199 ( .A(n1248), .B(n1247), .S(n8286), .Z(n1249) );
  MUX2_X1 U20200 ( .A(n1249), .B(n1246), .S(n8239), .Z(n1250) );
  MUX2_X1 U20201 ( .A(\mem[790][1] ), .B(\mem[791][1] ), .S(n8459), .Z(n1251)
         );
  MUX2_X1 U20202 ( .A(\mem[788][1] ), .B(\mem[789][1] ), .S(n8400), .Z(n1252)
         );
  MUX2_X1 U20203 ( .A(n1252), .B(n1251), .S(n8348), .Z(n1253) );
  MUX2_X1 U20204 ( .A(\mem[786][1] ), .B(\mem[787][1] ), .S(n8506), .Z(n1254)
         );
  MUX2_X1 U20205 ( .A(\mem[784][1] ), .B(\mem[785][1] ), .S(n8385), .Z(n1255)
         );
  MUX2_X1 U20206 ( .A(n1255), .B(n1254), .S(n8311), .Z(n1256) );
  MUX2_X1 U20207 ( .A(n1256), .B(n1253), .S(n8239), .Z(n1257) );
  MUX2_X1 U20208 ( .A(n1257), .B(n1250), .S(n8219), .Z(n1258) );
  MUX2_X1 U20209 ( .A(\mem[782][1] ), .B(\mem[783][1] ), .S(n8384), .Z(n1259)
         );
  MUX2_X1 U20210 ( .A(\mem[780][1] ), .B(\mem[781][1] ), .S(n8383), .Z(n1260)
         );
  MUX2_X1 U20211 ( .A(n1260), .B(n1259), .S(n8282), .Z(n1261) );
  MUX2_X1 U20212 ( .A(\mem[778][1] ), .B(\mem[779][1] ), .S(n8414), .Z(n1262)
         );
  MUX2_X1 U20213 ( .A(\mem[776][1] ), .B(\mem[777][1] ), .S(n8437), .Z(n1263)
         );
  MUX2_X1 U20214 ( .A(n1263), .B(n1262), .S(n8329), .Z(n1264) );
  MUX2_X1 U20215 ( .A(n1264), .B(n1261), .S(n8239), .Z(n1265) );
  MUX2_X1 U20216 ( .A(\mem[774][1] ), .B(\mem[775][1] ), .S(n8523), .Z(n1266)
         );
  MUX2_X1 U20217 ( .A(\mem[772][1] ), .B(\mem[773][1] ), .S(n8429), .Z(n1267)
         );
  MUX2_X1 U20218 ( .A(n1267), .B(n1266), .S(n8278), .Z(n1268) );
  MUX2_X1 U20219 ( .A(\mem[770][1] ), .B(\mem[771][1] ), .S(n8538), .Z(n1269)
         );
  MUX2_X1 U20220 ( .A(\mem[768][1] ), .B(\mem[769][1] ), .S(n8359), .Z(n1270)
         );
  MUX2_X1 U20221 ( .A(n1270), .B(n1269), .S(n8277), .Z(n1271) );
  MUX2_X1 U20222 ( .A(n1271), .B(n1268), .S(n8239), .Z(n1272) );
  MUX2_X1 U20223 ( .A(n1272), .B(n1265), .S(n8209), .Z(n1273) );
  MUX2_X1 U20224 ( .A(n1273), .B(n1258), .S(n8193), .Z(n1274) );
  MUX2_X1 U20225 ( .A(n1274), .B(n1243), .S(n8181), .Z(n1275) );
  MUX2_X1 U20226 ( .A(n1275), .B(n1212), .S(n8179), .Z(n1276) );
  MUX2_X1 U20227 ( .A(n1276), .B(n1149), .S(N25), .Z(n1277) );
  MUX2_X1 U20228 ( .A(\mem[766][1] ), .B(\mem[767][1] ), .S(n8422), .Z(n1278)
         );
  MUX2_X1 U20229 ( .A(\mem[764][1] ), .B(\mem[765][1] ), .S(n8535), .Z(n1279)
         );
  MUX2_X1 U20230 ( .A(n1279), .B(n1278), .S(n8352), .Z(n1280) );
  MUX2_X1 U20231 ( .A(\mem[762][1] ), .B(\mem[763][1] ), .S(n8402), .Z(n1281)
         );
  MUX2_X1 U20232 ( .A(\mem[760][1] ), .B(\mem[761][1] ), .S(n8534), .Z(n1282)
         );
  MUX2_X1 U20233 ( .A(n1282), .B(n1281), .S(n8271), .Z(n1283) );
  MUX2_X1 U20234 ( .A(n1283), .B(n1280), .S(n8240), .Z(n1284) );
  MUX2_X1 U20235 ( .A(\mem[758][1] ), .B(\mem[759][1] ), .S(n8387), .Z(n1285)
         );
  MUX2_X1 U20236 ( .A(\mem[756][1] ), .B(\mem[757][1] ), .S(n8365), .Z(n1286)
         );
  MUX2_X1 U20237 ( .A(n1286), .B(n1285), .S(n8281), .Z(n1287) );
  MUX2_X1 U20238 ( .A(\mem[754][1] ), .B(\mem[755][1] ), .S(N18), .Z(n1288) );
  MUX2_X1 U20239 ( .A(\mem[752][1] ), .B(\mem[753][1] ), .S(n8405), .Z(n1289)
         );
  MUX2_X1 U20240 ( .A(n1289), .B(n1288), .S(n8280), .Z(n1290) );
  MUX2_X1 U20241 ( .A(n1290), .B(n1287), .S(n8240), .Z(n1291) );
  MUX2_X1 U20242 ( .A(n1291), .B(n1284), .S(N21), .Z(n1292) );
  MUX2_X1 U20243 ( .A(\mem[750][1] ), .B(\mem[751][1] ), .S(n8526), .Z(n1293)
         );
  MUX2_X1 U20244 ( .A(\mem[748][1] ), .B(\mem[749][1] ), .S(n8516), .Z(n1294)
         );
  MUX2_X1 U20245 ( .A(n1294), .B(n1293), .S(n8279), .Z(n1295) );
  MUX2_X1 U20246 ( .A(\mem[746][1] ), .B(\mem[747][1] ), .S(n8495), .Z(n1296)
         );
  MUX2_X1 U20247 ( .A(\mem[744][1] ), .B(\mem[745][1] ), .S(n8486), .Z(n1297)
         );
  MUX2_X1 U20248 ( .A(n1297), .B(n1296), .S(n8320), .Z(n1298) );
  MUX2_X1 U20249 ( .A(n1298), .B(n1295), .S(n8240), .Z(n1299) );
  MUX2_X1 U20250 ( .A(\mem[742][1] ), .B(\mem[743][1] ), .S(n8374), .Z(n1300)
         );
  MUX2_X1 U20251 ( .A(\mem[740][1] ), .B(\mem[741][1] ), .S(n8364), .Z(n1301)
         );
  MUX2_X1 U20252 ( .A(n1301), .B(n1300), .S(n8271), .Z(n1302) );
  MUX2_X1 U20253 ( .A(\mem[738][1] ), .B(\mem[739][1] ), .S(n8381), .Z(n1303)
         );
  MUX2_X1 U20254 ( .A(\mem[736][1] ), .B(\mem[737][1] ), .S(n8470), .Z(n1304)
         );
  MUX2_X1 U20255 ( .A(n1304), .B(n1303), .S(n8268), .Z(n1305) );
  MUX2_X1 U20256 ( .A(n1305), .B(n1302), .S(n8240), .Z(n1306) );
  MUX2_X1 U20257 ( .A(n1306), .B(n1299), .S(n8202), .Z(n1307) );
  MUX2_X1 U20258 ( .A(n1307), .B(n1292), .S(N22), .Z(n1308) );
  MUX2_X1 U20259 ( .A(\mem[734][1] ), .B(\mem[735][1] ), .S(n8456), .Z(n1309)
         );
  MUX2_X1 U20260 ( .A(\mem[732][1] ), .B(\mem[733][1] ), .S(n8442), .Z(n1310)
         );
  MUX2_X1 U20261 ( .A(n1310), .B(n1309), .S(n8270), .Z(n1311) );
  MUX2_X1 U20262 ( .A(\mem[730][1] ), .B(\mem[731][1] ), .S(n8416), .Z(n1312)
         );
  MUX2_X1 U20263 ( .A(\mem[728][1] ), .B(\mem[729][1] ), .S(n8369), .Z(n1313)
         );
  MUX2_X1 U20264 ( .A(n1313), .B(n1312), .S(n8293), .Z(n1314) );
  MUX2_X1 U20265 ( .A(n1314), .B(n1311), .S(n8240), .Z(n1315) );
  MUX2_X1 U20266 ( .A(\mem[726][1] ), .B(\mem[727][1] ), .S(n8493), .Z(n1316)
         );
  MUX2_X1 U20267 ( .A(\mem[724][1] ), .B(\mem[725][1] ), .S(n8422), .Z(n1317)
         );
  MUX2_X1 U20268 ( .A(n1317), .B(n1316), .S(n8291), .Z(n1318) );
  MUX2_X1 U20269 ( .A(\mem[722][1] ), .B(\mem[723][1] ), .S(n8536), .Z(n1319)
         );
  MUX2_X1 U20270 ( .A(\mem[720][1] ), .B(\mem[721][1] ), .S(n8358), .Z(n1320)
         );
  MUX2_X1 U20271 ( .A(n1320), .B(n1319), .S(n8356), .Z(n1321) );
  MUX2_X1 U20272 ( .A(n1321), .B(n1318), .S(n8240), .Z(n1322) );
  MUX2_X1 U20273 ( .A(n1322), .B(n1315), .S(n8197), .Z(n1323) );
  MUX2_X1 U20274 ( .A(\mem[718][1] ), .B(\mem[719][1] ), .S(n8370), .Z(n1324)
         );
  MUX2_X1 U20275 ( .A(\mem[716][1] ), .B(\mem[717][1] ), .S(n8367), .Z(n1325)
         );
  MUX2_X1 U20276 ( .A(n1325), .B(n1324), .S(n8282), .Z(n1326) );
  MUX2_X1 U20277 ( .A(\mem[714][1] ), .B(\mem[715][1] ), .S(n8464), .Z(n1327)
         );
  MUX2_X1 U20278 ( .A(\mem[712][1] ), .B(\mem[713][1] ), .S(n8399), .Z(n1328)
         );
  MUX2_X1 U20279 ( .A(n1328), .B(n1327), .S(n8334), .Z(n1329) );
  MUX2_X1 U20280 ( .A(n1329), .B(n1326), .S(n8240), .Z(n1330) );
  MUX2_X1 U20281 ( .A(\mem[710][1] ), .B(\mem[711][1] ), .S(n8377), .Z(n1331)
         );
  MUX2_X1 U20282 ( .A(\mem[708][1] ), .B(\mem[709][1] ), .S(n8376), .Z(n1332)
         );
  MUX2_X1 U20283 ( .A(n1332), .B(n1331), .S(n8278), .Z(n1333) );
  MUX2_X1 U20284 ( .A(\mem[706][1] ), .B(\mem[707][1] ), .S(n8375), .Z(n1334)
         );
  MUX2_X1 U20285 ( .A(\mem[704][1] ), .B(\mem[705][1] ), .S(n8393), .Z(n1335)
         );
  MUX2_X1 U20286 ( .A(n1335), .B(n1334), .S(n8277), .Z(n1336) );
  MUX2_X1 U20287 ( .A(n1336), .B(n1333), .S(n8240), .Z(n1337) );
  MUX2_X1 U20288 ( .A(n1337), .B(n1330), .S(n8200), .Z(n1338) );
  MUX2_X1 U20289 ( .A(n1338), .B(n1323), .S(n8186), .Z(n1339) );
  MUX2_X1 U20290 ( .A(n1339), .B(n1308), .S(n8182), .Z(n1340) );
  MUX2_X1 U20291 ( .A(\mem[702][1] ), .B(\mem[703][1] ), .S(n8526), .Z(n1341)
         );
  MUX2_X1 U20292 ( .A(\mem[700][1] ), .B(\mem[701][1] ), .S(n8421), .Z(n1342)
         );
  MUX2_X1 U20293 ( .A(n1342), .B(n1341), .S(n8276), .Z(n1343) );
  MUX2_X1 U20294 ( .A(\mem[698][1] ), .B(\mem[699][1] ), .S(n8456), .Z(n1344)
         );
  MUX2_X1 U20295 ( .A(\mem[696][1] ), .B(\mem[697][1] ), .S(n8505), .Z(n1345)
         );
  MUX2_X1 U20296 ( .A(n1345), .B(n1344), .S(n8275), .Z(n1346) );
  MUX2_X1 U20297 ( .A(n1346), .B(n1343), .S(n8240), .Z(n1347) );
  MUX2_X1 U20298 ( .A(\mem[694][1] ), .B(\mem[695][1] ), .S(n8362), .Z(n1348)
         );
  MUX2_X1 U20299 ( .A(\mem[692][1] ), .B(\mem[693][1] ), .S(n8380), .Z(n1349)
         );
  MUX2_X1 U20300 ( .A(n1349), .B(n1348), .S(n8274), .Z(n1350) );
  MUX2_X1 U20301 ( .A(\mem[690][1] ), .B(\mem[691][1] ), .S(n8466), .Z(n1351)
         );
  MUX2_X1 U20302 ( .A(\mem[688][1] ), .B(\mem[689][1] ), .S(n8458), .Z(n1352)
         );
  MUX2_X1 U20303 ( .A(n1352), .B(n1351), .S(n8273), .Z(n1353) );
  MUX2_X1 U20304 ( .A(n1353), .B(n1350), .S(n8240), .Z(n1354) );
  MUX2_X1 U20305 ( .A(n1354), .B(n1347), .S(n8199), .Z(n1355) );
  MUX2_X1 U20306 ( .A(\mem[686][1] ), .B(\mem[687][1] ), .S(n8462), .Z(n1356)
         );
  MUX2_X1 U20307 ( .A(\mem[684][1] ), .B(\mem[685][1] ), .S(n8411), .Z(n1357)
         );
  MUX2_X1 U20308 ( .A(n1357), .B(n1356), .S(n8275), .Z(n1358) );
  MUX2_X1 U20309 ( .A(\mem[682][1] ), .B(\mem[683][1] ), .S(n8375), .Z(n1359)
         );
  MUX2_X1 U20310 ( .A(\mem[680][1] ), .B(\mem[681][1] ), .S(n8433), .Z(n1360)
         );
  MUX2_X1 U20311 ( .A(n1360), .B(n1359), .S(n8278), .Z(n1361) );
  MUX2_X1 U20312 ( .A(n1361), .B(n1358), .S(n8240), .Z(n1362) );
  MUX2_X1 U20313 ( .A(\mem[678][1] ), .B(\mem[679][1] ), .S(n8462), .Z(n1363)
         );
  MUX2_X1 U20314 ( .A(\mem[676][1] ), .B(\mem[677][1] ), .S(n8454), .Z(n1364)
         );
  MUX2_X1 U20315 ( .A(n1364), .B(n1363), .S(n8318), .Z(n1365) );
  MUX2_X1 U20316 ( .A(\mem[674][1] ), .B(\mem[675][1] ), .S(n8444), .Z(n1366)
         );
  MUX2_X1 U20317 ( .A(\mem[672][1] ), .B(\mem[673][1] ), .S(n8449), .Z(n1367)
         );
  MUX2_X1 U20318 ( .A(n1367), .B(n1366), .S(n8272), .Z(n1368) );
  MUX2_X1 U20319 ( .A(n1368), .B(n1365), .S(n8240), .Z(n1369) );
  MUX2_X1 U20320 ( .A(n1369), .B(n1362), .S(n8198), .Z(n1370) );
  MUX2_X1 U20321 ( .A(n1370), .B(n1355), .S(n8195), .Z(n1371) );
  MUX2_X1 U20322 ( .A(\mem[670][1] ), .B(\mem[671][1] ), .S(n8451), .Z(n1372)
         );
  MUX2_X1 U20323 ( .A(\mem[668][1] ), .B(\mem[669][1] ), .S(n8501), .Z(n1373)
         );
  MUX2_X1 U20324 ( .A(n1373), .B(n1372), .S(n8278), .Z(n1374) );
  MUX2_X1 U20325 ( .A(\mem[666][1] ), .B(\mem[667][1] ), .S(n8385), .Z(n1375)
         );
  MUX2_X1 U20326 ( .A(\mem[664][1] ), .B(\mem[665][1] ), .S(n8384), .Z(n1376)
         );
  MUX2_X1 U20327 ( .A(n1376), .B(n1375), .S(n8277), .Z(n1377) );
  MUX2_X1 U20328 ( .A(n1377), .B(n1374), .S(n8241), .Z(n1378) );
  MUX2_X1 U20329 ( .A(\mem[662][1] ), .B(\mem[663][1] ), .S(n8383), .Z(n1379)
         );
  MUX2_X1 U20330 ( .A(\mem[660][1] ), .B(\mem[661][1] ), .S(n8380), .Z(n1380)
         );
  MUX2_X1 U20331 ( .A(n1380), .B(n1379), .S(n8269), .Z(n1381) );
  MUX2_X1 U20332 ( .A(\mem[658][1] ), .B(\mem[659][1] ), .S(n8379), .Z(n1382)
         );
  MUX2_X1 U20333 ( .A(\mem[656][1] ), .B(\mem[657][1] ), .S(n8378), .Z(n1383)
         );
  MUX2_X1 U20334 ( .A(n1383), .B(n1382), .S(n8276), .Z(n1384) );
  MUX2_X1 U20335 ( .A(n1384), .B(n1381), .S(n8241), .Z(n1385) );
  MUX2_X1 U20336 ( .A(n1385), .B(n1378), .S(n8219), .Z(n1386) );
  MUX2_X1 U20337 ( .A(\mem[654][1] ), .B(\mem[655][1] ), .S(n8377), .Z(n1387)
         );
  MUX2_X1 U20338 ( .A(\mem[652][1] ), .B(\mem[653][1] ), .S(n8376), .Z(n1388)
         );
  MUX2_X1 U20339 ( .A(n1388), .B(n1387), .S(n8266), .Z(n1389) );
  MUX2_X1 U20340 ( .A(\mem[650][1] ), .B(\mem[651][1] ), .S(n8375), .Z(n1390)
         );
  MUX2_X1 U20341 ( .A(\mem[648][1] ), .B(\mem[649][1] ), .S(n8374), .Z(n1391)
         );
  MUX2_X1 U20342 ( .A(n1391), .B(n1390), .S(n8278), .Z(n1392) );
  MUX2_X1 U20343 ( .A(n1392), .B(n1389), .S(n8241), .Z(n1393) );
  MUX2_X1 U20344 ( .A(\mem[646][1] ), .B(\mem[647][1] ), .S(n8375), .Z(n1394)
         );
  MUX2_X1 U20345 ( .A(\mem[644][1] ), .B(\mem[645][1] ), .S(n8375), .Z(n1395)
         );
  MUX2_X1 U20346 ( .A(n1395), .B(n1394), .S(n8267), .Z(n1396) );
  MUX2_X1 U20347 ( .A(\mem[642][1] ), .B(\mem[643][1] ), .S(n8478), .Z(n1397)
         );
  MUX2_X1 U20348 ( .A(\mem[640][1] ), .B(\mem[641][1] ), .S(n8362), .Z(n1398)
         );
  MUX2_X1 U20349 ( .A(n1398), .B(n1397), .S(n8277), .Z(n1399) );
  MUX2_X1 U20350 ( .A(n1399), .B(n1396), .S(n8241), .Z(n1400) );
  MUX2_X1 U20351 ( .A(n1400), .B(n1393), .S(n8215), .Z(n1401) );
  MUX2_X1 U20352 ( .A(n1401), .B(n1386), .S(n8188), .Z(n1402) );
  MUX2_X1 U20353 ( .A(n1402), .B(n1371), .S(n8182), .Z(n1403) );
  MUX2_X1 U20354 ( .A(n1403), .B(n1340), .S(n8179), .Z(n1404) );
  MUX2_X1 U20355 ( .A(\mem[638][1] ), .B(\mem[639][1] ), .S(n8387), .Z(n1405)
         );
  MUX2_X1 U20356 ( .A(\mem[636][1] ), .B(\mem[637][1] ), .S(n8460), .Z(n1406)
         );
  MUX2_X1 U20357 ( .A(n1406), .B(n1405), .S(n8356), .Z(n1407) );
  MUX2_X1 U20358 ( .A(\mem[634][1] ), .B(\mem[635][1] ), .S(n8395), .Z(n1408)
         );
  MUX2_X1 U20359 ( .A(\mem[632][1] ), .B(\mem[633][1] ), .S(n8416), .Z(n1409)
         );
  MUX2_X1 U20360 ( .A(n1409), .B(n1408), .S(n8284), .Z(n1410) );
  MUX2_X1 U20361 ( .A(n1410), .B(n1407), .S(n8241), .Z(n1411) );
  MUX2_X1 U20362 ( .A(\mem[630][1] ), .B(\mem[631][1] ), .S(n8390), .Z(n1412)
         );
  MUX2_X1 U20363 ( .A(\mem[628][1] ), .B(\mem[629][1] ), .S(n8534), .Z(n1413)
         );
  MUX2_X1 U20364 ( .A(n1413), .B(n1412), .S(n8347), .Z(n1414) );
  MUX2_X1 U20365 ( .A(\mem[626][1] ), .B(\mem[627][1] ), .S(n8458), .Z(n1415)
         );
  MUX2_X1 U20366 ( .A(\mem[624][1] ), .B(\mem[625][1] ), .S(n8530), .Z(n1416)
         );
  MUX2_X1 U20367 ( .A(n1416), .B(n1415), .S(n8316), .Z(n1417) );
  MUX2_X1 U20368 ( .A(n1417), .B(n1414), .S(n8241), .Z(n1418) );
  MUX2_X1 U20369 ( .A(n1418), .B(n1411), .S(N21), .Z(n1419) );
  MUX2_X1 U20370 ( .A(\mem[622][1] ), .B(\mem[623][1] ), .S(n8537), .Z(n1420)
         );
  MUX2_X1 U20371 ( .A(\mem[620][1] ), .B(\mem[621][1] ), .S(n8539), .Z(n1421)
         );
  MUX2_X1 U20372 ( .A(n1421), .B(n1420), .S(n8268), .Z(n1422) );
  MUX2_X1 U20373 ( .A(\mem[618][1] ), .B(\mem[619][1] ), .S(n8364), .Z(n1423)
         );
  MUX2_X1 U20374 ( .A(\mem[616][1] ), .B(\mem[617][1] ), .S(n8363), .Z(n1424)
         );
  MUX2_X1 U20375 ( .A(n1424), .B(n1423), .S(n8266), .Z(n1425) );
  MUX2_X1 U20376 ( .A(n1425), .B(n1422), .S(n8241), .Z(n1426) );
  MUX2_X1 U20377 ( .A(\mem[614][1] ), .B(\mem[615][1] ), .S(n8373), .Z(n1427)
         );
  MUX2_X1 U20378 ( .A(\mem[612][1] ), .B(\mem[613][1] ), .S(n8367), .Z(n1428)
         );
  MUX2_X1 U20379 ( .A(n1428), .B(n1427), .S(n8267), .Z(n1429) );
  MUX2_X1 U20380 ( .A(\mem[610][1] ), .B(\mem[611][1] ), .S(n8366), .Z(n1430)
         );
  MUX2_X1 U20381 ( .A(\mem[608][1] ), .B(\mem[609][1] ), .S(n8373), .Z(n1431)
         );
  MUX2_X1 U20382 ( .A(n1431), .B(n1430), .S(n8279), .Z(n1432) );
  MUX2_X1 U20383 ( .A(n1432), .B(n1429), .S(n8241), .Z(n1433) );
  MUX2_X1 U20384 ( .A(n1433), .B(n1426), .S(n8197), .Z(n1434) );
  MUX2_X1 U20385 ( .A(n1434), .B(n1419), .S(n8196), .Z(n1435) );
  MUX2_X1 U20386 ( .A(\mem[606][1] ), .B(\mem[607][1] ), .S(n8363), .Z(n1436)
         );
  MUX2_X1 U20387 ( .A(\mem[604][1] ), .B(\mem[605][1] ), .S(n8371), .Z(n1437)
         );
  MUX2_X1 U20388 ( .A(n1437), .B(n1436), .S(n8269), .Z(n1438) );
  MUX2_X1 U20389 ( .A(\mem[602][1] ), .B(\mem[603][1] ), .S(n8372), .Z(n1439)
         );
  MUX2_X1 U20390 ( .A(\mem[600][1] ), .B(\mem[601][1] ), .S(n8524), .Z(n1440)
         );
  MUX2_X1 U20391 ( .A(n1440), .B(n1439), .S(n8301), .Z(n1441) );
  MUX2_X1 U20392 ( .A(n1441), .B(n1438), .S(n8241), .Z(n1442) );
  MUX2_X1 U20393 ( .A(\mem[598][1] ), .B(\mem[599][1] ), .S(n8403), .Z(n1443)
         );
  MUX2_X1 U20394 ( .A(\mem[596][1] ), .B(\mem[597][1] ), .S(n8470), .Z(n1444)
         );
  MUX2_X1 U20395 ( .A(n1444), .B(n1443), .S(n8310), .Z(n1445) );
  MUX2_X1 U20396 ( .A(\mem[594][1] ), .B(\mem[595][1] ), .S(n8360), .Z(n1446)
         );
  MUX2_X1 U20397 ( .A(\mem[592][1] ), .B(\mem[593][1] ), .S(n8361), .Z(n1447)
         );
  MUX2_X1 U20398 ( .A(n1447), .B(n1446), .S(n8281), .Z(n1448) );
  MUX2_X1 U20399 ( .A(n1448), .B(n1445), .S(n8241), .Z(n1449) );
  MUX2_X1 U20400 ( .A(n1449), .B(n1442), .S(n8210), .Z(n1450) );
  MUX2_X1 U20401 ( .A(\mem[590][1] ), .B(\mem[591][1] ), .S(n8358), .Z(n1451)
         );
  MUX2_X1 U20402 ( .A(\mem[588][1] ), .B(\mem[589][1] ), .S(n8434), .Z(n1452)
         );
  MUX2_X1 U20403 ( .A(n1452), .B(n1451), .S(n8277), .Z(n1453) );
  MUX2_X1 U20404 ( .A(\mem[586][1] ), .B(\mem[587][1] ), .S(n8482), .Z(n1454)
         );
  MUX2_X1 U20405 ( .A(\mem[584][1] ), .B(\mem[585][1] ), .S(n8376), .Z(n1455)
         );
  MUX2_X1 U20406 ( .A(n1455), .B(n1454), .S(n8276), .Z(n1456) );
  MUX2_X1 U20407 ( .A(n1456), .B(n1453), .S(n8241), .Z(n1457) );
  MUX2_X1 U20408 ( .A(\mem[582][1] ), .B(\mem[583][1] ), .S(n8455), .Z(n1458)
         );
  MUX2_X1 U20409 ( .A(\mem[580][1] ), .B(\mem[581][1] ), .S(n8368), .Z(n1459)
         );
  MUX2_X1 U20410 ( .A(n1459), .B(n1458), .S(n8321), .Z(n1460) );
  MUX2_X1 U20411 ( .A(\mem[578][1] ), .B(\mem[579][1] ), .S(n8539), .Z(n1461)
         );
  MUX2_X1 U20412 ( .A(\mem[576][1] ), .B(\mem[577][1] ), .S(n8362), .Z(n1462)
         );
  MUX2_X1 U20413 ( .A(n1462), .B(n1461), .S(n8271), .Z(n1463) );
  MUX2_X1 U20414 ( .A(n1463), .B(n1460), .S(n8241), .Z(n1464) );
  MUX2_X1 U20415 ( .A(n1464), .B(n1457), .S(n8219), .Z(n1465) );
  MUX2_X1 U20416 ( .A(n1465), .B(n1450), .S(n8187), .Z(n1466) );
  MUX2_X1 U20417 ( .A(n1466), .B(n1435), .S(n8182), .Z(n1467) );
  MUX2_X1 U20418 ( .A(\mem[574][1] ), .B(\mem[575][1] ), .S(n8385), .Z(n1468)
         );
  MUX2_X1 U20419 ( .A(\mem[572][1] ), .B(\mem[573][1] ), .S(n8384), .Z(n1469)
         );
  MUX2_X1 U20420 ( .A(n1469), .B(n1468), .S(n8339), .Z(n1470) );
  MUX2_X1 U20421 ( .A(\mem[570][1] ), .B(\mem[571][1] ), .S(n8383), .Z(n1471)
         );
  MUX2_X1 U20422 ( .A(\mem[568][1] ), .B(\mem[569][1] ), .S(n8447), .Z(n1472)
         );
  MUX2_X1 U20423 ( .A(n1472), .B(n1471), .S(n8275), .Z(n1473) );
  MUX2_X1 U20424 ( .A(n1473), .B(n1470), .S(n8242), .Z(n1474) );
  MUX2_X1 U20425 ( .A(\mem[566][1] ), .B(\mem[567][1] ), .S(N18), .Z(n1475) );
  MUX2_X1 U20426 ( .A(\mem[564][1] ), .B(\mem[565][1] ), .S(n8477), .Z(n1476)
         );
  MUX2_X1 U20427 ( .A(n1476), .B(n1475), .S(N19), .Z(n1477) );
  MUX2_X1 U20428 ( .A(\mem[562][1] ), .B(\mem[563][1] ), .S(n8458), .Z(n1478)
         );
  MUX2_X1 U20429 ( .A(\mem[560][1] ), .B(\mem[561][1] ), .S(n8436), .Z(n1479)
         );
  MUX2_X1 U20430 ( .A(n1479), .B(n1478), .S(n8356), .Z(n1480) );
  MUX2_X1 U20431 ( .A(n1480), .B(n1477), .S(n8242), .Z(n1481) );
  MUX2_X1 U20432 ( .A(n1481), .B(n1474), .S(n8203), .Z(n1482) );
  MUX2_X1 U20433 ( .A(\mem[558][1] ), .B(\mem[559][1] ), .S(n8465), .Z(n1483)
         );
  MUX2_X1 U20434 ( .A(\mem[556][1] ), .B(\mem[557][1] ), .S(n8441), .Z(n1484)
         );
  MUX2_X1 U20435 ( .A(n1484), .B(n1483), .S(n8350), .Z(n1485) );
  MUX2_X1 U20436 ( .A(\mem[554][1] ), .B(\mem[555][1] ), .S(n8538), .Z(n1486)
         );
  MUX2_X1 U20437 ( .A(\mem[552][1] ), .B(\mem[553][1] ), .S(n8359), .Z(n1487)
         );
  MUX2_X1 U20438 ( .A(n1487), .B(n1486), .S(n8274), .Z(n1488) );
  MUX2_X1 U20439 ( .A(n1488), .B(n1485), .S(n8242), .Z(n1489) );
  MUX2_X1 U20440 ( .A(\mem[550][1] ), .B(\mem[551][1] ), .S(n8386), .Z(n1490)
         );
  MUX2_X1 U20441 ( .A(\mem[548][1] ), .B(\mem[549][1] ), .S(n8361), .Z(n1491)
         );
  MUX2_X1 U20442 ( .A(n1491), .B(n1490), .S(n8280), .Z(n1492) );
  MUX2_X1 U20443 ( .A(\mem[546][1] ), .B(\mem[547][1] ), .S(n8366), .Z(n1493)
         );
  MUX2_X1 U20444 ( .A(\mem[544][1] ), .B(\mem[545][1] ), .S(n8519), .Z(n1494)
         );
  MUX2_X1 U20445 ( .A(n1494), .B(n1493), .S(n8279), .Z(n1495) );
  MUX2_X1 U20446 ( .A(n1495), .B(n1492), .S(n8242), .Z(n1496) );
  MUX2_X1 U20447 ( .A(n1496), .B(n1489), .S(n8207), .Z(n1497) );
  MUX2_X1 U20448 ( .A(n1497), .B(n1482), .S(n8196), .Z(n1498) );
  MUX2_X1 U20449 ( .A(\mem[542][1] ), .B(\mem[543][1] ), .S(n8376), .Z(n1499)
         );
  MUX2_X1 U20450 ( .A(\mem[540][1] ), .B(\mem[541][1] ), .S(n8444), .Z(n1500)
         );
  MUX2_X1 U20451 ( .A(n1500), .B(n1499), .S(n8332), .Z(n1501) );
  MUX2_X1 U20452 ( .A(\mem[538][1] ), .B(\mem[539][1] ), .S(n8514), .Z(n1502)
         );
  MUX2_X1 U20453 ( .A(\mem[536][1] ), .B(\mem[537][1] ), .S(n8505), .Z(n1503)
         );
  MUX2_X1 U20454 ( .A(n1503), .B(n1502), .S(n8278), .Z(n1504) );
  MUX2_X1 U20455 ( .A(n1504), .B(n1501), .S(n8242), .Z(n1505) );
  MUX2_X1 U20456 ( .A(\mem[534][1] ), .B(\mem[535][1] ), .S(n8485), .Z(n1506)
         );
  MUX2_X1 U20457 ( .A(\mem[532][1] ), .B(\mem[533][1] ), .S(n8417), .Z(n1507)
         );
  MUX2_X1 U20458 ( .A(n1507), .B(n1506), .S(n8272), .Z(n1508) );
  MUX2_X1 U20459 ( .A(\mem[530][1] ), .B(\mem[531][1] ), .S(n8409), .Z(n1509)
         );
  MUX2_X1 U20460 ( .A(\mem[528][1] ), .B(\mem[529][1] ), .S(n8400), .Z(n1510)
         );
  MUX2_X1 U20461 ( .A(n1510), .B(n1509), .S(n8275), .Z(n1511) );
  MUX2_X1 U20462 ( .A(n1511), .B(n1508), .S(n8242), .Z(n1512) );
  MUX2_X1 U20463 ( .A(n1512), .B(n1505), .S(n8200), .Z(n1513) );
  MUX2_X1 U20464 ( .A(\mem[526][1] ), .B(\mem[527][1] ), .S(n8537), .Z(n1514)
         );
  MUX2_X1 U20465 ( .A(\mem[524][1] ), .B(\mem[525][1] ), .S(n8434), .Z(n1515)
         );
  MUX2_X1 U20466 ( .A(n1515), .B(n1514), .S(n8277), .Z(n1516) );
  MUX2_X1 U20467 ( .A(\mem[522][1] ), .B(\mem[523][1] ), .S(n8382), .Z(n1517)
         );
  MUX2_X1 U20468 ( .A(\mem[520][1] ), .B(\mem[521][1] ), .S(n8456), .Z(n1518)
         );
  MUX2_X1 U20469 ( .A(n1518), .B(n1517), .S(n8276), .Z(n1519) );
  MUX2_X1 U20470 ( .A(n1519), .B(n1516), .S(n8242), .Z(n1520) );
  MUX2_X1 U20471 ( .A(\mem[518][1] ), .B(\mem[519][1] ), .S(n8460), .Z(n1521)
         );
  MUX2_X1 U20472 ( .A(\mem[516][1] ), .B(\mem[517][1] ), .S(n8448), .Z(n1522)
         );
  MUX2_X1 U20473 ( .A(n1522), .B(n1521), .S(n8322), .Z(n1523) );
  MUX2_X1 U20474 ( .A(\mem[514][1] ), .B(\mem[515][1] ), .S(n8520), .Z(n1524)
         );
  MUX2_X1 U20475 ( .A(\mem[512][1] ), .B(\mem[513][1] ), .S(n8538), .Z(n1525)
         );
  MUX2_X1 U20476 ( .A(n1525), .B(n1524), .S(n8271), .Z(n1526) );
  MUX2_X1 U20477 ( .A(n1526), .B(n1523), .S(n8242), .Z(n1527) );
  MUX2_X1 U20478 ( .A(n1527), .B(n1520), .S(n8199), .Z(n1528) );
  MUX2_X1 U20479 ( .A(n1528), .B(n1513), .S(n8196), .Z(n1529) );
  MUX2_X1 U20480 ( .A(n1529), .B(n1498), .S(n8182), .Z(n1530) );
  MUX2_X1 U20481 ( .A(n1530), .B(n1467), .S(n8179), .Z(n1531) );
  MUX2_X1 U20482 ( .A(n1531), .B(n1404), .S(N25), .Z(n1532) );
  MUX2_X1 U20483 ( .A(n1532), .B(n1277), .S(N26), .Z(n1533) );
  MUX2_X1 U20484 ( .A(\mem[510][1] ), .B(\mem[511][1] ), .S(n8445), .Z(n1534)
         );
  MUX2_X1 U20485 ( .A(\mem[508][1] ), .B(\mem[509][1] ), .S(n8511), .Z(n1535)
         );
  MUX2_X1 U20486 ( .A(n1535), .B(n1534), .S(n8275), .Z(n1536) );
  MUX2_X1 U20487 ( .A(\mem[506][1] ), .B(\mem[507][1] ), .S(n8402), .Z(n1537)
         );
  MUX2_X1 U20488 ( .A(\mem[504][1] ), .B(\mem[505][1] ), .S(n8518), .Z(n1538)
         );
  MUX2_X1 U20489 ( .A(n1538), .B(n1537), .S(n8273), .Z(n1539) );
  MUX2_X1 U20490 ( .A(n1539), .B(n1536), .S(n8242), .Z(n1540) );
  MUX2_X1 U20491 ( .A(\mem[502][1] ), .B(\mem[503][1] ), .S(n8370), .Z(n1541)
         );
  MUX2_X1 U20492 ( .A(\mem[500][1] ), .B(\mem[501][1] ), .S(n8369), .Z(n1542)
         );
  MUX2_X1 U20493 ( .A(n1542), .B(n1541), .S(n8282), .Z(n1543) );
  MUX2_X1 U20494 ( .A(\mem[498][1] ), .B(\mem[499][1] ), .S(n8487), .Z(n1544)
         );
  MUX2_X1 U20495 ( .A(\mem[496][1] ), .B(\mem[497][1] ), .S(n8436), .Z(n1545)
         );
  MUX2_X1 U20496 ( .A(n1545), .B(n1544), .S(n8268), .Z(n1546) );
  MUX2_X1 U20497 ( .A(n1546), .B(n1543), .S(n8242), .Z(n1547) );
  MUX2_X1 U20498 ( .A(n1547), .B(n1540), .S(n8198), .Z(n1548) );
  MUX2_X1 U20499 ( .A(\mem[494][1] ), .B(\mem[495][1] ), .S(n8473), .Z(n1549)
         );
  MUX2_X1 U20500 ( .A(\mem[492][1] ), .B(\mem[493][1] ), .S(n8411), .Z(n1550)
         );
  MUX2_X1 U20501 ( .A(n1550), .B(n1549), .S(n8314), .Z(n1551) );
  MUX2_X1 U20502 ( .A(\mem[490][1] ), .B(\mem[491][1] ), .S(n8480), .Z(n1552)
         );
  MUX2_X1 U20503 ( .A(\mem[488][1] ), .B(\mem[489][1] ), .S(n8481), .Z(n1553)
         );
  MUX2_X1 U20504 ( .A(n1553), .B(n1552), .S(n8353), .Z(n1554) );
  MUX2_X1 U20505 ( .A(n1554), .B(n1551), .S(n8242), .Z(n1555) );
  MUX2_X1 U20506 ( .A(\mem[486][1] ), .B(\mem[487][1] ), .S(n8374), .Z(n1556)
         );
  MUX2_X1 U20507 ( .A(\mem[484][1] ), .B(\mem[485][1] ), .S(n8525), .Z(n1557)
         );
  MUX2_X1 U20508 ( .A(n1557), .B(n1556), .S(n8269), .Z(n1558) );
  MUX2_X1 U20509 ( .A(\mem[482][1] ), .B(\mem[483][1] ), .S(n8384), .Z(n1559)
         );
  MUX2_X1 U20510 ( .A(\mem[480][1] ), .B(\mem[481][1] ), .S(n8534), .Z(n1560)
         );
  MUX2_X1 U20511 ( .A(n1560), .B(n1559), .S(n8270), .Z(n1561) );
  MUX2_X1 U20512 ( .A(n1561), .B(n1558), .S(n8242), .Z(n1562) );
  MUX2_X1 U20513 ( .A(n1562), .B(n1555), .S(n8208), .Z(n1563) );
  MUX2_X1 U20514 ( .A(n1563), .B(n1548), .S(n8187), .Z(n1564) );
  MUX2_X1 U20515 ( .A(\mem[478][1] ), .B(\mem[479][1] ), .S(n8516), .Z(n1565)
         );
  MUX2_X1 U20516 ( .A(\mem[476][1] ), .B(\mem[477][1] ), .S(n8450), .Z(n1566)
         );
  MUX2_X1 U20517 ( .A(n1566), .B(n1565), .S(n8343), .Z(n1567) );
  MUX2_X1 U20518 ( .A(\mem[474][1] ), .B(\mem[475][1] ), .S(n8451), .Z(n1568)
         );
  MUX2_X1 U20519 ( .A(\mem[472][1] ), .B(\mem[473][1] ), .S(n8452), .Z(n1569)
         );
  MUX2_X1 U20520 ( .A(n1569), .B(n1568), .S(n8272), .Z(n1570) );
  MUX2_X1 U20521 ( .A(n1570), .B(n1567), .S(n8243), .Z(n1571) );
  MUX2_X1 U20522 ( .A(\mem[470][1] ), .B(\mem[471][1] ), .S(n8447), .Z(n1572)
         );
  MUX2_X1 U20523 ( .A(\mem[468][1] ), .B(\mem[469][1] ), .S(n8448), .Z(n1573)
         );
  MUX2_X1 U20524 ( .A(n1573), .B(n1572), .S(n8276), .Z(n1574) );
  MUX2_X1 U20525 ( .A(\mem[466][1] ), .B(\mem[467][1] ), .S(n8449), .Z(n1575)
         );
  MUX2_X1 U20526 ( .A(\mem[464][1] ), .B(\mem[465][1] ), .S(n8456), .Z(n1576)
         );
  MUX2_X1 U20527 ( .A(n1576), .B(n1575), .S(n8266), .Z(n1577) );
  MUX2_X1 U20528 ( .A(n1577), .B(n1574), .S(n8243), .Z(n1578) );
  MUX2_X1 U20529 ( .A(n1578), .B(n1571), .S(n8197), .Z(n1579) );
  MUX2_X1 U20530 ( .A(\mem[462][1] ), .B(\mem[463][1] ), .S(n8457), .Z(n1580)
         );
  MUX2_X1 U20531 ( .A(\mem[460][1] ), .B(\mem[461][1] ), .S(n8458), .Z(n1581)
         );
  MUX2_X1 U20532 ( .A(n1581), .B(n1580), .S(n8267), .Z(n1582) );
  MUX2_X1 U20533 ( .A(\mem[458][1] ), .B(\mem[459][1] ), .S(n8453), .Z(n1583)
         );
  MUX2_X1 U20534 ( .A(\mem[456][1] ), .B(\mem[457][1] ), .S(n8454), .Z(n1584)
         );
  MUX2_X1 U20535 ( .A(n1584), .B(n1583), .S(n8280), .Z(n1585) );
  MUX2_X1 U20536 ( .A(n1585), .B(n1582), .S(n8243), .Z(n1586) );
  MUX2_X1 U20537 ( .A(\mem[454][1] ), .B(\mem[455][1] ), .S(n8489), .Z(n1587)
         );
  MUX2_X1 U20538 ( .A(\mem[452][1] ), .B(\mem[453][1] ), .S(n8438), .Z(n1588)
         );
  MUX2_X1 U20539 ( .A(n1588), .B(n1587), .S(n8345), .Z(n1589) );
  MUX2_X1 U20540 ( .A(\mem[450][1] ), .B(\mem[451][1] ), .S(n8439), .Z(n1590)
         );
  MUX2_X1 U20541 ( .A(\mem[448][1] ), .B(\mem[449][1] ), .S(n8440), .Z(n1591)
         );
  MUX2_X1 U20542 ( .A(n1591), .B(n1590), .S(n8281), .Z(n1592) );
  MUX2_X1 U20543 ( .A(n1592), .B(n1589), .S(n8243), .Z(n1593) );
  MUX2_X1 U20544 ( .A(n1593), .B(n1586), .S(n8206), .Z(n1594) );
  MUX2_X1 U20545 ( .A(n1594), .B(n1579), .S(n8195), .Z(n1595) );
  MUX2_X1 U20546 ( .A(n1595), .B(n1564), .S(n8182), .Z(n1596) );
  MUX2_X1 U20547 ( .A(\mem[446][1] ), .B(\mem[447][1] ), .S(n8435), .Z(n1597)
         );
  MUX2_X1 U20548 ( .A(\mem[444][1] ), .B(\mem[445][1] ), .S(n8436), .Z(n1598)
         );
  MUX2_X1 U20549 ( .A(n1598), .B(n1597), .S(n8277), .Z(n1599) );
  MUX2_X1 U20550 ( .A(\mem[442][1] ), .B(\mem[443][1] ), .S(n8437), .Z(n1600)
         );
  MUX2_X1 U20551 ( .A(\mem[440][1] ), .B(\mem[441][1] ), .S(n8444), .Z(n1601)
         );
  MUX2_X1 U20552 ( .A(n1601), .B(n1600), .S(n8276), .Z(n1602) );
  MUX2_X1 U20553 ( .A(n1602), .B(n1599), .S(n8243), .Z(n1603) );
  MUX2_X1 U20554 ( .A(\mem[438][1] ), .B(\mem[439][1] ), .S(n8445), .Z(n1604)
         );
  MUX2_X1 U20555 ( .A(\mem[436][1] ), .B(\mem[437][1] ), .S(n8446), .Z(n1605)
         );
  MUX2_X1 U20556 ( .A(n1605), .B(n1604), .S(n8272), .Z(n1606) );
  MUX2_X1 U20557 ( .A(\mem[434][1] ), .B(\mem[435][1] ), .S(n8441), .Z(n1607)
         );
  MUX2_X1 U20558 ( .A(\mem[432][1] ), .B(\mem[433][1] ), .S(n8442), .Z(n1608)
         );
  MUX2_X1 U20559 ( .A(n1608), .B(n1607), .S(n8271), .Z(n1609) );
  MUX2_X1 U20560 ( .A(n1609), .B(n1606), .S(n8243), .Z(n1610) );
  MUX2_X1 U20561 ( .A(n1610), .B(n1603), .S(n8219), .Z(n1611) );
  MUX2_X1 U20562 ( .A(\mem[430][1] ), .B(\mem[431][1] ), .S(n8419), .Z(n1612)
         );
  MUX2_X1 U20563 ( .A(\mem[428][1] ), .B(\mem[429][1] ), .S(n8522), .Z(n1613)
         );
  MUX2_X1 U20564 ( .A(n1613), .B(n1612), .S(n8306), .Z(n1614) );
  MUX2_X1 U20565 ( .A(\mem[426][1] ), .B(\mem[427][1] ), .S(n8504), .Z(n1615)
         );
  MUX2_X1 U20566 ( .A(\mem[424][1] ), .B(\mem[425][1] ), .S(n8425), .Z(n1616)
         );
  MUX2_X1 U20567 ( .A(n1616), .B(n1615), .S(n8270), .Z(n1617) );
  MUX2_X1 U20568 ( .A(n1617), .B(n1614), .S(n8243), .Z(n1618) );
  MUX2_X1 U20569 ( .A(\mem[422][1] ), .B(\mem[423][1] ), .S(n8461), .Z(n1619)
         );
  MUX2_X1 U20570 ( .A(\mem[420][1] ), .B(\mem[421][1] ), .S(n8394), .Z(n1620)
         );
  MUX2_X1 U20571 ( .A(n1620), .B(n1619), .S(n8309), .Z(n1621) );
  MUX2_X1 U20572 ( .A(\mem[418][1] ), .B(\mem[419][1] ), .S(n8466), .Z(n1622)
         );
  MUX2_X1 U20573 ( .A(\mem[416][1] ), .B(\mem[417][1] ), .S(n8432), .Z(n1623)
         );
  MUX2_X1 U20574 ( .A(n1623), .B(n1622), .S(n8271), .Z(n1624) );
  MUX2_X1 U20575 ( .A(n1624), .B(n1621), .S(n8243), .Z(n1625) );
  MUX2_X1 U20576 ( .A(n1625), .B(n1618), .S(n8197), .Z(n1626) );
  MUX2_X1 U20577 ( .A(n1626), .B(n1611), .S(n8190), .Z(n1627) );
  MUX2_X1 U20578 ( .A(\mem[414][1] ), .B(\mem[415][1] ), .S(n8433), .Z(n1628)
         );
  MUX2_X1 U20579 ( .A(\mem[412][1] ), .B(\mem[413][1] ), .S(n8434), .Z(n1629)
         );
  MUX2_X1 U20580 ( .A(n1629), .B(n1628), .S(N19), .Z(n1630) );
  MUX2_X1 U20581 ( .A(\mem[410][1] ), .B(\mem[411][1] ), .S(n8429), .Z(n1631)
         );
  MUX2_X1 U20582 ( .A(\mem[408][1] ), .B(\mem[409][1] ), .S(n8430), .Z(n1632)
         );
  MUX2_X1 U20583 ( .A(n1632), .B(n1631), .S(n8356), .Z(n1633) );
  MUX2_X1 U20584 ( .A(n1633), .B(n1630), .S(n8243), .Z(n1634) );
  MUX2_X1 U20585 ( .A(\mem[406][1] ), .B(\mem[407][1] ), .S(n8528), .Z(n1635)
         );
  MUX2_X1 U20586 ( .A(\mem[404][1] ), .B(\mem[405][1] ), .S(n8502), .Z(n1636)
         );
  MUX2_X1 U20587 ( .A(n1636), .B(n1635), .S(n8343), .Z(n1637) );
  MUX2_X1 U20588 ( .A(\mem[402][1] ), .B(\mem[403][1] ), .S(n8483), .Z(n1638)
         );
  MUX2_X1 U20589 ( .A(\mem[400][1] ), .B(\mem[401][1] ), .S(n8374), .Z(n1639)
         );
  MUX2_X1 U20590 ( .A(n1639), .B(n1638), .S(n8274), .Z(n1640) );
  MUX2_X1 U20591 ( .A(n1640), .B(n1637), .S(n8243), .Z(n1641) );
  MUX2_X1 U20592 ( .A(n1641), .B(n1634), .S(n8212), .Z(n1642) );
  MUX2_X1 U20593 ( .A(\mem[398][1] ), .B(\mem[399][1] ), .S(n8367), .Z(n1643)
         );
  MUX2_X1 U20594 ( .A(\mem[396][1] ), .B(\mem[397][1] ), .S(n8390), .Z(n1644)
         );
  MUX2_X1 U20595 ( .A(n1644), .B(n1643), .S(n8280), .Z(n1645) );
  MUX2_X1 U20596 ( .A(\mem[394][1] ), .B(\mem[395][1] ), .S(n8512), .Z(n1646)
         );
  MUX2_X1 U20597 ( .A(\mem[392][1] ), .B(\mem[393][1] ), .S(n8493), .Z(n1647)
         );
  MUX2_X1 U20598 ( .A(n1647), .B(n1646), .S(n8279), .Z(n1648) );
  MUX2_X1 U20599 ( .A(n1648), .B(n1645), .S(n8243), .Z(n1649) );
  MUX2_X1 U20600 ( .A(\mem[390][1] ), .B(\mem[391][1] ), .S(n8410), .Z(n1650)
         );
  MUX2_X1 U20601 ( .A(\mem[388][1] ), .B(\mem[389][1] ), .S(n8412), .Z(n1651)
         );
  MUX2_X1 U20602 ( .A(n1651), .B(n1650), .S(n8325), .Z(n1652) );
  MUX2_X1 U20603 ( .A(\mem[386][1] ), .B(\mem[387][1] ), .S(n8441), .Z(n1653)
         );
  MUX2_X1 U20604 ( .A(\mem[384][1] ), .B(\mem[385][1] ), .S(n8438), .Z(n1654)
         );
  MUX2_X1 U20605 ( .A(n1654), .B(n1653), .S(n8278), .Z(n1655) );
  MUX2_X1 U20606 ( .A(n1655), .B(n1652), .S(n8243), .Z(n1656) );
  MUX2_X1 U20607 ( .A(n1656), .B(n1649), .S(N21), .Z(n1657) );
  MUX2_X1 U20608 ( .A(n1657), .B(n1642), .S(n8189), .Z(n1658) );
  MUX2_X1 U20609 ( .A(n1658), .B(n1627), .S(n8182), .Z(n1659) );
  MUX2_X1 U20610 ( .A(n1659), .B(n1596), .S(n8179), .Z(n1660) );
  MUX2_X1 U20611 ( .A(\mem[382][1] ), .B(\mem[383][1] ), .S(n8482), .Z(n1661)
         );
  MUX2_X1 U20612 ( .A(\mem[380][1] ), .B(\mem[381][1] ), .S(n8475), .Z(n1662)
         );
  MUX2_X1 U20613 ( .A(n1662), .B(n1661), .S(n8282), .Z(n1663) );
  MUX2_X1 U20614 ( .A(\mem[378][1] ), .B(\mem[379][1] ), .S(n8476), .Z(n1664)
         );
  MUX2_X1 U20615 ( .A(\mem[376][1] ), .B(\mem[377][1] ), .S(n8471), .Z(n1665)
         );
  MUX2_X1 U20616 ( .A(n1665), .B(n1664), .S(n8275), .Z(n1666) );
  MUX2_X1 U20617 ( .A(n1666), .B(n1663), .S(n8244), .Z(n1667) );
  MUX2_X1 U20618 ( .A(\mem[374][1] ), .B(\mem[375][1] ), .S(n8472), .Z(n1668)
         );
  MUX2_X1 U20619 ( .A(\mem[372][1] ), .B(\mem[373][1] ), .S(n8473), .Z(n1669)
         );
  MUX2_X1 U20620 ( .A(n1669), .B(n1668), .S(n8273), .Z(n1670) );
  MUX2_X1 U20621 ( .A(\mem[370][1] ), .B(\mem[371][1] ), .S(n8480), .Z(n1671)
         );
  MUX2_X1 U20622 ( .A(\mem[368][1] ), .B(\mem[369][1] ), .S(n8454), .Z(n1672)
         );
  MUX2_X1 U20623 ( .A(n1672), .B(n1671), .S(n8355), .Z(n1673) );
  MUX2_X1 U20624 ( .A(n1673), .B(n1670), .S(n8244), .Z(n1674) );
  MUX2_X1 U20625 ( .A(n1674), .B(n1667), .S(n8199), .Z(n1675) );
  MUX2_X1 U20626 ( .A(\mem[366][1] ), .B(\mem[367][1] ), .S(n8359), .Z(n1676)
         );
  MUX2_X1 U20627 ( .A(\mem[364][1] ), .B(\mem[365][1] ), .S(n8373), .Z(n1677)
         );
  MUX2_X1 U20628 ( .A(n1677), .B(n1676), .S(n8329), .Z(n1678) );
  MUX2_X1 U20629 ( .A(\mem[362][1] ), .B(\mem[363][1] ), .S(n8388), .Z(n1679)
         );
  MUX2_X1 U20630 ( .A(\mem[360][1] ), .B(\mem[361][1] ), .S(n8470), .Z(n1680)
         );
  MUX2_X1 U20631 ( .A(n1680), .B(n1679), .S(n8294), .Z(n1681) );
  MUX2_X1 U20632 ( .A(n1681), .B(n1678), .S(n8244), .Z(n1682) );
  MUX2_X1 U20633 ( .A(\mem[358][1] ), .B(\mem[359][1] ), .S(n8462), .Z(n1683)
         );
  MUX2_X1 U20634 ( .A(\mem[356][1] ), .B(\mem[357][1] ), .S(n8463), .Z(n1684)
         );
  MUX2_X1 U20635 ( .A(n1684), .B(n1683), .S(n8350), .Z(n1685) );
  MUX2_X1 U20636 ( .A(\mem[354][1] ), .B(\mem[355][1] ), .S(n8464), .Z(n1686)
         );
  MUX2_X1 U20637 ( .A(\mem[352][1] ), .B(\mem[353][1] ), .S(n8459), .Z(n1687)
         );
  MUX2_X1 U20638 ( .A(n1687), .B(n1686), .S(n8307), .Z(n1688) );
  MUX2_X1 U20639 ( .A(n1688), .B(n1685), .S(n8244), .Z(n1689) );
  MUX2_X1 U20640 ( .A(n1689), .B(n1682), .S(n8209), .Z(n1690) );
  MUX2_X1 U20641 ( .A(n1690), .B(n1675), .S(n8188), .Z(n1691) );
  MUX2_X1 U20642 ( .A(\mem[350][1] ), .B(\mem[351][1] ), .S(n8460), .Z(n1692)
         );
  MUX2_X1 U20643 ( .A(\mem[348][1] ), .B(\mem[349][1] ), .S(n8461), .Z(n1693)
         );
  MUX2_X1 U20644 ( .A(n1693), .B(n1692), .S(n8282), .Z(n1694) );
  MUX2_X1 U20645 ( .A(\mem[346][1] ), .B(\mem[347][1] ), .S(n8468), .Z(n1695)
         );
  MUX2_X1 U20646 ( .A(\mem[344][1] ), .B(\mem[345][1] ), .S(n8469), .Z(n1696)
         );
  MUX2_X1 U20647 ( .A(n1696), .B(n1695), .S(n8268), .Z(n1697) );
  MUX2_X1 U20648 ( .A(n1697), .B(n1694), .S(n8244), .Z(n1698) );
  MUX2_X1 U20649 ( .A(\mem[342][1] ), .B(\mem[343][1] ), .S(n8470), .Z(n1699)
         );
  MUX2_X1 U20650 ( .A(\mem[340][1] ), .B(\mem[341][1] ), .S(n8465), .Z(n1700)
         );
  MUX2_X1 U20651 ( .A(n1700), .B(n1699), .S(n8287), .Z(n1701) );
  MUX2_X1 U20652 ( .A(\mem[338][1] ), .B(\mem[339][1] ), .S(n8466), .Z(n1702)
         );
  MUX2_X1 U20653 ( .A(\mem[336][1] ), .B(\mem[337][1] ), .S(n8467), .Z(n1703)
         );
  MUX2_X1 U20654 ( .A(n1703), .B(n1702), .S(n8269), .Z(n1704) );
  MUX2_X1 U20655 ( .A(n1704), .B(n1701), .S(n8244), .Z(n1705) );
  MUX2_X1 U20656 ( .A(n1705), .B(n1698), .S(n8200), .Z(n1706) );
  MUX2_X1 U20657 ( .A(\mem[334][1] ), .B(\mem[335][1] ), .S(n8366), .Z(n1707)
         );
  MUX2_X1 U20658 ( .A(\mem[332][1] ), .B(\mem[333][1] ), .S(n8373), .Z(n1708)
         );
  MUX2_X1 U20659 ( .A(n1708), .B(n1707), .S(n8279), .Z(n1709) );
  MUX2_X1 U20660 ( .A(\mem[330][1] ), .B(\mem[331][1] ), .S(n8363), .Z(n1710)
         );
  MUX2_X1 U20661 ( .A(\mem[328][1] ), .B(\mem[329][1] ), .S(n8372), .Z(n1711)
         );
  MUX2_X1 U20662 ( .A(n1711), .B(n1710), .S(n8279), .Z(n1712) );
  MUX2_X1 U20663 ( .A(n1712), .B(n1709), .S(n8244), .Z(n1713) );
  MUX2_X1 U20664 ( .A(\mem[326][1] ), .B(\mem[327][1] ), .S(n8371), .Z(n1714)
         );
  MUX2_X1 U20665 ( .A(\mem[324][1] ), .B(\mem[325][1] ), .S(n8370), .Z(n1715)
         );
  MUX2_X1 U20666 ( .A(n1715), .B(n1714), .S(n8269), .Z(n1716) );
  MUX2_X1 U20667 ( .A(\mem[322][1] ), .B(\mem[323][1] ), .S(n8369), .Z(n1717)
         );
  MUX2_X1 U20668 ( .A(\mem[320][1] ), .B(\mem[321][1] ), .S(n8368), .Z(n1718)
         );
  MUX2_X1 U20669 ( .A(n1718), .B(n1717), .S(n8270), .Z(n1719) );
  MUX2_X1 U20670 ( .A(n1719), .B(n1716), .S(n8244), .Z(n1720) );
  MUX2_X1 U20671 ( .A(n1720), .B(n1713), .S(n8199), .Z(n1721) );
  MUX2_X1 U20672 ( .A(n1721), .B(n1706), .S(n8195), .Z(n1722) );
  MUX2_X1 U20673 ( .A(n1722), .B(n1691), .S(n8182), .Z(n1723) );
  MUX2_X1 U20674 ( .A(\mem[318][1] ), .B(\mem[319][1] ), .S(n8367), .Z(n1724)
         );
  MUX2_X1 U20675 ( .A(\mem[316][1] ), .B(\mem[317][1] ), .S(n8364), .Z(n1725)
         );
  MUX2_X1 U20676 ( .A(n1725), .B(n1724), .S(n8332), .Z(n1726) );
  MUX2_X1 U20677 ( .A(\mem[314][1] ), .B(\mem[315][1] ), .S(n8362), .Z(n1727)
         );
  MUX2_X1 U20678 ( .A(\mem[312][1] ), .B(\mem[313][1] ), .S(n8539), .Z(n1728)
         );
  MUX2_X1 U20679 ( .A(n1728), .B(n1727), .S(n8306), .Z(n1729) );
  MUX2_X1 U20680 ( .A(n1729), .B(n1726), .S(n8244), .Z(n1730) );
  MUX2_X1 U20681 ( .A(\mem[310][1] ), .B(\mem[311][1] ), .S(n8362), .Z(n1731)
         );
  MUX2_X1 U20682 ( .A(\mem[308][1] ), .B(\mem[309][1] ), .S(n8366), .Z(n1732)
         );
  MUX2_X1 U20683 ( .A(n1732), .B(n1731), .S(n8323), .Z(n1733) );
  MUX2_X1 U20684 ( .A(\mem[306][1] ), .B(\mem[307][1] ), .S(n8373), .Z(n1734)
         );
  MUX2_X1 U20685 ( .A(\mem[304][1] ), .B(\mem[305][1] ), .S(n8363), .Z(n1735)
         );
  MUX2_X1 U20686 ( .A(n1735), .B(n1734), .S(n8322), .Z(n1736) );
  MUX2_X1 U20687 ( .A(n1736), .B(n1733), .S(n8244), .Z(n1737) );
  MUX2_X1 U20688 ( .A(n1737), .B(n1730), .S(n8198), .Z(n1738) );
  MUX2_X1 U20689 ( .A(\mem[302][1] ), .B(\mem[303][1] ), .S(n8372), .Z(n1739)
         );
  MUX2_X1 U20690 ( .A(\mem[300][1] ), .B(\mem[301][1] ), .S(n8371), .Z(n1740)
         );
  MUX2_X1 U20691 ( .A(n1740), .B(n1739), .S(n8341), .Z(n1741) );
  MUX2_X1 U20692 ( .A(\mem[298][1] ), .B(\mem[299][1] ), .S(n8370), .Z(n1742)
         );
  MUX2_X1 U20693 ( .A(\mem[296][1] ), .B(\mem[297][1] ), .S(n8369), .Z(n1743)
         );
  MUX2_X1 U20694 ( .A(n1743), .B(n1742), .S(n8288), .Z(n1744) );
  MUX2_X1 U20695 ( .A(n1744), .B(n1741), .S(n8244), .Z(n1745) );
  MUX2_X1 U20696 ( .A(\mem[294][1] ), .B(\mem[295][1] ), .S(n8368), .Z(n1746)
         );
  MUX2_X1 U20697 ( .A(\mem[292][1] ), .B(\mem[293][1] ), .S(n8367), .Z(n1747)
         );
  MUX2_X1 U20698 ( .A(n1747), .B(n1746), .S(n8333), .Z(n1748) );
  MUX2_X1 U20699 ( .A(\mem[290][1] ), .B(\mem[291][1] ), .S(n8364), .Z(n1749)
         );
  MUX2_X1 U20700 ( .A(\mem[288][1] ), .B(\mem[289][1] ), .S(n8539), .Z(n1750)
         );
  MUX2_X1 U20701 ( .A(n1750), .B(n1749), .S(n8296), .Z(n1751) );
  MUX2_X1 U20702 ( .A(n1751), .B(n1748), .S(n8244), .Z(n1752) );
  MUX2_X1 U20703 ( .A(n1752), .B(n1745), .S(n8204), .Z(n1753) );
  MUX2_X1 U20704 ( .A(n1753), .B(n1738), .S(n8192), .Z(n1754) );
  MUX2_X1 U20705 ( .A(\mem[286][1] ), .B(\mem[287][1] ), .S(n8539), .Z(n1755)
         );
  MUX2_X1 U20706 ( .A(\mem[284][1] ), .B(\mem[285][1] ), .S(n8362), .Z(n1756)
         );
  MUX2_X1 U20707 ( .A(n1756), .B(n1755), .S(n8324), .Z(n1757) );
  MUX2_X1 U20708 ( .A(\mem[282][1] ), .B(\mem[283][1] ), .S(n8366), .Z(n1758)
         );
  MUX2_X1 U20709 ( .A(\mem[280][1] ), .B(\mem[281][1] ), .S(n8373), .Z(n1759)
         );
  MUX2_X1 U20710 ( .A(n1759), .B(n1758), .S(n8344), .Z(n1760) );
  MUX2_X1 U20711 ( .A(n1760), .B(n1757), .S(n8245), .Z(n1761) );
  MUX2_X1 U20712 ( .A(\mem[278][1] ), .B(\mem[279][1] ), .S(n8363), .Z(n1762)
         );
  MUX2_X1 U20713 ( .A(\mem[276][1] ), .B(\mem[277][1] ), .S(n8372), .Z(n1763)
         );
  MUX2_X1 U20714 ( .A(n1763), .B(n1762), .S(n8345), .Z(n1764) );
  MUX2_X1 U20715 ( .A(\mem[274][1] ), .B(\mem[275][1] ), .S(n8371), .Z(n1765)
         );
  MUX2_X1 U20716 ( .A(\mem[272][1] ), .B(\mem[273][1] ), .S(n8370), .Z(n1766)
         );
  MUX2_X1 U20717 ( .A(n1766), .B(n1765), .S(n8346), .Z(n1767) );
  MUX2_X1 U20718 ( .A(n1767), .B(n1764), .S(n8245), .Z(n1768) );
  MUX2_X1 U20719 ( .A(n1768), .B(n1761), .S(n8213), .Z(n1769) );
  MUX2_X1 U20720 ( .A(\mem[270][1] ), .B(\mem[271][1] ), .S(n8369), .Z(n1770)
         );
  MUX2_X1 U20721 ( .A(\mem[268][1] ), .B(\mem[269][1] ), .S(n8368), .Z(n1771)
         );
  MUX2_X1 U20722 ( .A(n1771), .B(n1770), .S(n8341), .Z(n1772) );
  MUX2_X1 U20723 ( .A(\mem[266][1] ), .B(\mem[267][1] ), .S(n8367), .Z(n1773)
         );
  MUX2_X1 U20724 ( .A(\mem[264][1] ), .B(\mem[265][1] ), .S(n8364), .Z(n1774)
         );
  MUX2_X1 U20725 ( .A(n1774), .B(n1773), .S(n8342), .Z(n1775) );
  MUX2_X1 U20726 ( .A(n1775), .B(n1772), .S(n8245), .Z(n1776) );
  MUX2_X1 U20727 ( .A(\mem[262][1] ), .B(\mem[263][1] ), .S(n8530), .Z(n1777)
         );
  MUX2_X1 U20728 ( .A(\mem[260][1] ), .B(\mem[261][1] ), .S(n8509), .Z(n1778)
         );
  MUX2_X1 U20729 ( .A(n1778), .B(n1777), .S(n8343), .Z(n1779) );
  MUX2_X1 U20730 ( .A(\mem[258][1] ), .B(\mem[259][1] ), .S(n8499), .Z(n1780)
         );
  MUX2_X1 U20731 ( .A(\mem[256][1] ), .B(\mem[257][1] ), .S(n8419), .Z(n1781)
         );
  MUX2_X1 U20732 ( .A(n1781), .B(n1780), .S(n8350), .Z(n1782) );
  MUX2_X1 U20733 ( .A(n1782), .B(n1779), .S(n8245), .Z(n1783) );
  MUX2_X1 U20734 ( .A(n1783), .B(n1776), .S(n8219), .Z(n1784) );
  MUX2_X1 U20735 ( .A(n1784), .B(n1769), .S(n8195), .Z(n1785) );
  MUX2_X1 U20736 ( .A(n1785), .B(n1754), .S(n8182), .Z(n1786) );
  MUX2_X1 U20737 ( .A(n1786), .B(n1723), .S(n8179), .Z(n1787) );
  MUX2_X1 U20738 ( .A(n1787), .B(n1660), .S(n8177), .Z(n1788) );
  MUX2_X1 U20739 ( .A(\mem[254][1] ), .B(\mem[255][1] ), .S(n8409), .Z(n1789)
         );
  MUX2_X1 U20740 ( .A(\mem[252][1] ), .B(\mem[253][1] ), .S(n8416), .Z(n1790)
         );
  MUX2_X1 U20741 ( .A(n1790), .B(n1789), .S(n8351), .Z(n1791) );
  MUX2_X1 U20742 ( .A(\mem[250][1] ), .B(\mem[251][1] ), .S(n8410), .Z(n1792)
         );
  MUX2_X1 U20743 ( .A(\mem[248][1] ), .B(\mem[249][1] ), .S(n8407), .Z(n1793)
         );
  MUX2_X1 U20744 ( .A(n1793), .B(n1792), .S(n8352), .Z(n1794) );
  MUX2_X1 U20745 ( .A(n1794), .B(n1791), .S(n8245), .Z(n1795) );
  MUX2_X1 U20746 ( .A(\mem[246][1] ), .B(\mem[247][1] ), .S(n8408), .Z(n1796)
         );
  MUX2_X1 U20747 ( .A(\mem[244][1] ), .B(\mem[245][1] ), .S(n8474), .Z(n1797)
         );
  MUX2_X1 U20748 ( .A(n1797), .B(n1796), .S(n8347), .Z(n1798) );
  MUX2_X1 U20749 ( .A(\mem[242][1] ), .B(\mem[243][1] ), .S(n8414), .Z(n1799)
         );
  MUX2_X1 U20750 ( .A(\mem[240][1] ), .B(\mem[241][1] ), .S(n8415), .Z(n1800)
         );
  MUX2_X1 U20751 ( .A(n1800), .B(n1799), .S(n8348), .Z(n1801) );
  MUX2_X1 U20752 ( .A(n1801), .B(n1798), .S(n8245), .Z(n1802) );
  MUX2_X1 U20753 ( .A(n1802), .B(n1795), .S(n8197), .Z(n1803) );
  MUX2_X1 U20754 ( .A(\mem[238][1] ), .B(\mem[239][1] ), .S(n8367), .Z(n1804)
         );
  MUX2_X1 U20755 ( .A(\mem[236][1] ), .B(\mem[237][1] ), .S(n8366), .Z(n1805)
         );
  MUX2_X1 U20756 ( .A(n1805), .B(n1804), .S(n8278), .Z(n1806) );
  MUX2_X1 U20757 ( .A(\mem[234][1] ), .B(\mem[235][1] ), .S(n8363), .Z(n1807)
         );
  MUX2_X1 U20758 ( .A(\mem[232][1] ), .B(\mem[233][1] ), .S(n8364), .Z(n1808)
         );
  MUX2_X1 U20759 ( .A(n1808), .B(n1807), .S(n8333), .Z(n1809) );
  MUX2_X1 U20760 ( .A(n1809), .B(n1806), .S(n8245), .Z(n1810) );
  MUX2_X1 U20761 ( .A(\mem[230][1] ), .B(\mem[231][1] ), .S(n8539), .Z(n1811)
         );
  MUX2_X1 U20762 ( .A(\mem[228][1] ), .B(\mem[229][1] ), .S(n8362), .Z(n1812)
         );
  MUX2_X1 U20763 ( .A(n1812), .B(n1811), .S(n8334), .Z(n1813) );
  MUX2_X1 U20764 ( .A(\mem[226][1] ), .B(\mem[227][1] ), .S(n8373), .Z(n1814)
         );
  MUX2_X1 U20765 ( .A(\mem[224][1] ), .B(\mem[225][1] ), .S(n8372), .Z(n1815)
         );
  MUX2_X1 U20766 ( .A(n1815), .B(n1814), .S(n8329), .Z(n1816) );
  MUX2_X1 U20767 ( .A(n1816), .B(n1813), .S(n8245), .Z(n1817) );
  MUX2_X1 U20768 ( .A(n1817), .B(n1810), .S(n8198), .Z(n1818) );
  MUX2_X1 U20769 ( .A(n1818), .B(n1803), .S(n8186), .Z(n1819) );
  MUX2_X1 U20770 ( .A(\mem[222][1] ), .B(\mem[223][1] ), .S(n8371), .Z(n1820)
         );
  MUX2_X1 U20771 ( .A(\mem[220][1] ), .B(\mem[221][1] ), .S(n8370), .Z(n1821)
         );
  MUX2_X1 U20772 ( .A(n1821), .B(n1820), .S(n8330), .Z(n1822) );
  MUX2_X1 U20773 ( .A(\mem[218][1] ), .B(\mem[219][1] ), .S(n8369), .Z(n1823)
         );
  MUX2_X1 U20774 ( .A(\mem[216][1] ), .B(\mem[217][1] ), .S(n8368), .Z(n1824)
         );
  MUX2_X1 U20775 ( .A(n1824), .B(n1823), .S(n8331), .Z(n1825) );
  MUX2_X1 U20776 ( .A(n1825), .B(n1822), .S(n8245), .Z(n1826) );
  MUX2_X1 U20777 ( .A(\mem[214][1] ), .B(\mem[215][1] ), .S(n8362), .Z(n1827)
         );
  MUX2_X1 U20778 ( .A(\mem[212][1] ), .B(\mem[213][1] ), .S(n8363), .Z(n1828)
         );
  MUX2_X1 U20779 ( .A(n1828), .B(n1827), .S(n8338), .Z(n1829) );
  MUX2_X1 U20780 ( .A(\mem[210][1] ), .B(\mem[211][1] ), .S(n8364), .Z(n1830)
         );
  MUX2_X1 U20781 ( .A(\mem[208][1] ), .B(\mem[209][1] ), .S(n8539), .Z(n1831)
         );
  MUX2_X1 U20782 ( .A(n1831), .B(n1830), .S(n8339), .Z(n1832) );
  MUX2_X1 U20783 ( .A(n1832), .B(n1829), .S(n8245), .Z(n1833) );
  MUX2_X1 U20784 ( .A(n1833), .B(n1826), .S(n8198), .Z(n1834) );
  MUX2_X1 U20785 ( .A(\mem[206][1] ), .B(\mem[207][1] ), .S(n8362), .Z(n1835)
         );
  MUX2_X1 U20786 ( .A(\mem[204][1] ), .B(\mem[205][1] ), .S(n8363), .Z(n1836)
         );
  MUX2_X1 U20787 ( .A(n1836), .B(n1835), .S(n8340), .Z(n1837) );
  MUX2_X1 U20788 ( .A(\mem[202][1] ), .B(\mem[203][1] ), .S(n8364), .Z(n1838)
         );
  MUX2_X1 U20789 ( .A(\mem[200][1] ), .B(\mem[201][1] ), .S(n8373), .Z(n1839)
         );
  MUX2_X1 U20790 ( .A(n1839), .B(n1838), .S(n8335), .Z(n1840) );
  MUX2_X1 U20791 ( .A(n1840), .B(n1837), .S(n8245), .Z(n1841) );
  MUX2_X1 U20792 ( .A(\mem[198][1] ), .B(\mem[199][1] ), .S(n8372), .Z(n1842)
         );
  MUX2_X1 U20793 ( .A(\mem[196][1] ), .B(\mem[197][1] ), .S(n8371), .Z(n1843)
         );
  MUX2_X1 U20794 ( .A(n1843), .B(n1842), .S(n8336), .Z(n1844) );
  MUX2_X1 U20795 ( .A(\mem[194][1] ), .B(\mem[195][1] ), .S(n8370), .Z(n1845)
         );
  MUX2_X1 U20796 ( .A(\mem[192][1] ), .B(\mem[193][1] ), .S(n8369), .Z(n1846)
         );
  MUX2_X1 U20797 ( .A(n1846), .B(n1845), .S(n8337), .Z(n1847) );
  MUX2_X1 U20798 ( .A(n1847), .B(n1844), .S(n8245), .Z(n1848) );
  MUX2_X1 U20799 ( .A(n1848), .B(n1841), .S(n8213), .Z(n1849) );
  MUX2_X1 U20800 ( .A(n1849), .B(n1834), .S(n8195), .Z(n1850) );
  MUX2_X1 U20801 ( .A(n1850), .B(n1819), .S(n8182), .Z(n1851) );
  MUX2_X1 U20802 ( .A(\mem[190][1] ), .B(\mem[191][1] ), .S(n8368), .Z(n1852)
         );
  MUX2_X1 U20803 ( .A(\mem[188][1] ), .B(\mem[189][1] ), .S(n8367), .Z(n1853)
         );
  MUX2_X1 U20804 ( .A(n1853), .B(n1852), .S(n8292), .Z(n1854) );
  MUX2_X1 U20805 ( .A(\mem[186][1] ), .B(\mem[187][1] ), .S(n8363), .Z(n1855)
         );
  MUX2_X1 U20806 ( .A(\mem[184][1] ), .B(\mem[185][1] ), .S(n8364), .Z(n1856)
         );
  MUX2_X1 U20807 ( .A(n1856), .B(n1855), .S(n8351), .Z(n1857) );
  MUX2_X1 U20808 ( .A(n1857), .B(n1854), .S(n8246), .Z(n1858) );
  MUX2_X1 U20809 ( .A(\mem[182][1] ), .B(\mem[183][1] ), .S(n8539), .Z(n1859)
         );
  MUX2_X1 U20810 ( .A(\mem[180][1] ), .B(\mem[181][1] ), .S(n8457), .Z(n1860)
         );
  MUX2_X1 U20811 ( .A(n1860), .B(n1859), .S(n8274), .Z(n1861) );
  MUX2_X1 U20812 ( .A(\mem[178][1] ), .B(\mem[179][1] ), .S(n8435), .Z(n1862)
         );
  MUX2_X1 U20813 ( .A(\mem[176][1] ), .B(\mem[177][1] ), .S(n8408), .Z(n1863)
         );
  MUX2_X1 U20814 ( .A(n1863), .B(n1862), .S(n8272), .Z(n1864) );
  MUX2_X1 U20815 ( .A(n1864), .B(n1861), .S(n8246), .Z(n1865) );
  MUX2_X1 U20816 ( .A(n1865), .B(n1858), .S(n8197), .Z(n1866) );
  MUX2_X1 U20817 ( .A(\mem[174][1] ), .B(\mem[175][1] ), .S(n8459), .Z(n1867)
         );
  MUX2_X1 U20818 ( .A(\mem[172][1] ), .B(\mem[173][1] ), .S(n8426), .Z(n1868)
         );
  MUX2_X1 U20819 ( .A(n1868), .B(n1867), .S(n8273), .Z(n1869) );
  MUX2_X1 U20820 ( .A(\mem[170][1] ), .B(\mem[171][1] ), .S(n8378), .Z(n1870)
         );
  MUX2_X1 U20821 ( .A(\mem[168][1] ), .B(\mem[169][1] ), .S(n8452), .Z(n1871)
         );
  MUX2_X1 U20822 ( .A(n1871), .B(n1870), .S(n8281), .Z(n1872) );
  MUX2_X1 U20823 ( .A(n1872), .B(n1869), .S(n8246), .Z(n1873) );
  MUX2_X1 U20824 ( .A(\mem[166][1] ), .B(\mem[167][1] ), .S(n8428), .Z(n1874)
         );
  MUX2_X1 U20825 ( .A(\mem[164][1] ), .B(\mem[165][1] ), .S(n8423), .Z(n1875)
         );
  MUX2_X1 U20826 ( .A(n1875), .B(n1874), .S(n8266), .Z(n1876) );
  MUX2_X1 U20827 ( .A(\mem[162][1] ), .B(\mem[163][1] ), .S(n8424), .Z(n1877)
         );
  MUX2_X1 U20828 ( .A(\mem[160][1] ), .B(\mem[161][1] ), .S(n8425), .Z(n1878)
         );
  MUX2_X1 U20829 ( .A(n1878), .B(n1877), .S(n8267), .Z(n1879) );
  MUX2_X1 U20830 ( .A(n1879), .B(n1876), .S(n8246), .Z(n1880) );
  MUX2_X1 U20831 ( .A(n1880), .B(n1873), .S(n8197), .Z(n1881) );
  MUX2_X1 U20832 ( .A(n1881), .B(n1866), .S(n8193), .Z(n1882) );
  MUX2_X1 U20833 ( .A(\mem[158][1] ), .B(\mem[159][1] ), .S(n8431), .Z(n1883)
         );
  MUX2_X1 U20834 ( .A(\mem[156][1] ), .B(\mem[157][1] ), .S(n8443), .Z(n1884)
         );
  MUX2_X1 U20835 ( .A(n1884), .B(n1883), .S(n8281), .Z(n1885) );
  MUX2_X1 U20836 ( .A(\mem[154][1] ), .B(\mem[155][1] ), .S(n8481), .Z(n1886)
         );
  MUX2_X1 U20837 ( .A(\mem[152][1] ), .B(\mem[153][1] ), .S(n8482), .Z(n1887)
         );
  MUX2_X1 U20838 ( .A(n1887), .B(n1886), .S(n8278), .Z(n1888) );
  MUX2_X1 U20839 ( .A(n1888), .B(n1885), .S(n8246), .Z(n1889) );
  MUX2_X1 U20840 ( .A(\mem[150][1] ), .B(\mem[151][1] ), .S(n8477), .Z(n1890)
         );
  MUX2_X1 U20841 ( .A(\mem[148][1] ), .B(\mem[149][1] ), .S(n8478), .Z(n1891)
         );
  MUX2_X1 U20842 ( .A(n1891), .B(n1890), .S(n8268), .Z(n1892) );
  MUX2_X1 U20843 ( .A(\mem[146][1] ), .B(\mem[147][1] ), .S(n8479), .Z(n1893)
         );
  MUX2_X1 U20844 ( .A(\mem[144][1] ), .B(\mem[145][1] ), .S(n8486), .Z(n1894)
         );
  MUX2_X1 U20845 ( .A(n1894), .B(n1893), .S(n8340), .Z(n1895) );
  MUX2_X1 U20846 ( .A(n1895), .B(n1892), .S(n8246), .Z(n1896) );
  MUX2_X1 U20847 ( .A(n1896), .B(n1889), .S(n8199), .Z(n1897) );
  MUX2_X1 U20848 ( .A(\mem[142][1] ), .B(\mem[143][1] ), .S(n8416), .Z(n1898)
         );
  MUX2_X1 U20849 ( .A(\mem[140][1] ), .B(\mem[141][1] ), .S(n8411), .Z(n1899)
         );
  MUX2_X1 U20850 ( .A(n1899), .B(n1898), .S(n8282), .Z(n1900) );
  MUX2_X1 U20851 ( .A(\mem[138][1] ), .B(\mem[139][1] ), .S(n8412), .Z(n1901)
         );
  MUX2_X1 U20852 ( .A(\mem[136][1] ), .B(\mem[137][1] ), .S(n8413), .Z(n1902)
         );
  MUX2_X1 U20853 ( .A(n1902), .B(n1901), .S(n8333), .Z(n1903) );
  MUX2_X1 U20854 ( .A(n1903), .B(n1900), .S(n8246), .Z(n1904) );
  MUX2_X1 U20855 ( .A(\mem[134][1] ), .B(\mem[135][1] ), .S(n8420), .Z(n1905)
         );
  MUX2_X1 U20856 ( .A(\mem[132][1] ), .B(\mem[133][1] ), .S(n8421), .Z(n1906)
         );
  MUX2_X1 U20857 ( .A(n1906), .B(n1905), .S(n8278), .Z(n1907) );
  MUX2_X1 U20858 ( .A(\mem[130][1] ), .B(\mem[131][1] ), .S(n8422), .Z(n1908)
         );
  MUX2_X1 U20859 ( .A(\mem[128][1] ), .B(\mem[129][1] ), .S(n8417), .Z(n1909)
         );
  MUX2_X1 U20860 ( .A(n1909), .B(n1908), .S(n8277), .Z(n1910) );
  MUX2_X1 U20861 ( .A(n1910), .B(n1907), .S(n8246), .Z(n1911) );
  MUX2_X1 U20862 ( .A(n1911), .B(n1904), .S(n8198), .Z(n1912) );
  MUX2_X1 U20863 ( .A(n1912), .B(n1897), .S(n8195), .Z(n1913) );
  MUX2_X1 U20864 ( .A(n1913), .B(n1882), .S(n8182), .Z(n1914) );
  MUX2_X1 U20865 ( .A(n1914), .B(n1851), .S(n8179), .Z(n1915) );
  MUX2_X1 U20866 ( .A(\mem[126][1] ), .B(\mem[127][1] ), .S(n8418), .Z(n1916)
         );
  MUX2_X1 U20867 ( .A(\mem[124][1] ), .B(\mem[125][1] ), .S(n8419), .Z(n1917)
         );
  MUX2_X1 U20868 ( .A(n1917), .B(n1916), .S(n8268), .Z(n1918) );
  MUX2_X1 U20869 ( .A(\mem[122][1] ), .B(\mem[123][1] ), .S(n8426), .Z(n1919)
         );
  MUX2_X1 U20870 ( .A(\mem[120][1] ), .B(\mem[121][1] ), .S(n8427), .Z(n1920)
         );
  MUX2_X1 U20871 ( .A(n1920), .B(n1919), .S(n8274), .Z(n1921) );
  MUX2_X1 U20872 ( .A(n1921), .B(n1918), .S(n8246), .Z(n1922) );
  MUX2_X1 U20873 ( .A(\mem[118][1] ), .B(\mem[119][1] ), .S(n8364), .Z(n1923)
         );
  MUX2_X1 U20874 ( .A(\mem[116][1] ), .B(\mem[117][1] ), .S(n8539), .Z(n1924)
         );
  MUX2_X1 U20875 ( .A(n1924), .B(n1923), .S(n8338), .Z(n1925) );
  MUX2_X1 U20876 ( .A(\mem[114][1] ), .B(\mem[115][1] ), .S(n8362), .Z(n1926)
         );
  MUX2_X1 U20877 ( .A(\mem[112][1] ), .B(\mem[113][1] ), .S(n8372), .Z(n1927)
         );
  MUX2_X1 U20878 ( .A(n1927), .B(n1926), .S(n8269), .Z(n1928) );
  MUX2_X1 U20879 ( .A(n1928), .B(n1925), .S(n8246), .Z(n1929) );
  MUX2_X1 U20880 ( .A(n1929), .B(n1922), .S(n8218), .Z(n1930) );
  MUX2_X1 U20881 ( .A(\mem[110][1] ), .B(\mem[111][1] ), .S(n8371), .Z(n1931)
         );
  MUX2_X1 U20882 ( .A(\mem[108][1] ), .B(\mem[109][1] ), .S(n8370), .Z(n1932)
         );
  MUX2_X1 U20883 ( .A(n1932), .B(n1931), .S(n8270), .Z(n1933) );
  MUX2_X1 U20884 ( .A(\mem[106][1] ), .B(\mem[107][1] ), .S(n8369), .Z(n1934)
         );
  MUX2_X1 U20885 ( .A(\mem[104][1] ), .B(\mem[105][1] ), .S(n8368), .Z(n1935)
         );
  MUX2_X1 U20886 ( .A(n1935), .B(n1934), .S(N19), .Z(n1936) );
  MUX2_X1 U20887 ( .A(n1936), .B(n1933), .S(n8246), .Z(n1937) );
  MUX2_X1 U20888 ( .A(\mem[102][1] ), .B(\mem[103][1] ), .S(n8367), .Z(n1938)
         );
  MUX2_X1 U20889 ( .A(\mem[100][1] ), .B(\mem[101][1] ), .S(n8366), .Z(n1939)
         );
  MUX2_X1 U20890 ( .A(n1939), .B(n1938), .S(n8274), .Z(n1940) );
  MUX2_X1 U20891 ( .A(\mem[98][1] ), .B(\mem[99][1] ), .S(n8373), .Z(n1941) );
  MUX2_X1 U20892 ( .A(\mem[96][1] ), .B(\mem[97][1] ), .S(n8363), .Z(n1942) );
  MUX2_X1 U20893 ( .A(n1942), .B(n1941), .S(n8356), .Z(n1943) );
  MUX2_X1 U20894 ( .A(n1943), .B(n1940), .S(n8246), .Z(n1944) );
  MUX2_X1 U20895 ( .A(n1944), .B(n1937), .S(n8198), .Z(n1945) );
  MUX2_X1 U20896 ( .A(n1945), .B(n1930), .S(n8191), .Z(n1946) );
  MUX2_X1 U20897 ( .A(\mem[94][1] ), .B(\mem[95][1] ), .S(n8363), .Z(n1947) );
  MUX2_X1 U20898 ( .A(\mem[92][1] ), .B(\mem[93][1] ), .S(n8364), .Z(n1948) );
  MUX2_X1 U20899 ( .A(n1948), .B(n1947), .S(n8280), .Z(n1949) );
  MUX2_X1 U20900 ( .A(\mem[90][1] ), .B(\mem[91][1] ), .S(n8539), .Z(n1950) );
  MUX2_X1 U20901 ( .A(\mem[88][1] ), .B(\mem[89][1] ), .S(n8362), .Z(n1951) );
  MUX2_X1 U20902 ( .A(n1951), .B(n1950), .S(n8353), .Z(n1952) );
  MUX2_X1 U20903 ( .A(n1952), .B(n1949), .S(n8247), .Z(n1953) );
  MUX2_X1 U20904 ( .A(\mem[86][1] ), .B(\mem[87][1] ), .S(n8372), .Z(n1954) );
  MUX2_X1 U20905 ( .A(\mem[84][1] ), .B(\mem[85][1] ), .S(n8371), .Z(n1955) );
  MUX2_X1 U20906 ( .A(n1955), .B(n1954), .S(n8354), .Z(n1956) );
  MUX2_X1 U20907 ( .A(\mem[82][1] ), .B(\mem[83][1] ), .S(n8370), .Z(n1957) );
  MUX2_X1 U20908 ( .A(\mem[80][1] ), .B(\mem[81][1] ), .S(n8369), .Z(n1958) );
  MUX2_X1 U20909 ( .A(n1958), .B(n1957), .S(n8355), .Z(n1959) );
  MUX2_X1 U20910 ( .A(n1959), .B(n1956), .S(n8247), .Z(n1960) );
  MUX2_X1 U20911 ( .A(n1960), .B(n1953), .S(n8200), .Z(n1961) );
  MUX2_X1 U20912 ( .A(\mem[78][1] ), .B(\mem[79][1] ), .S(n8368), .Z(n1962) );
  MUX2_X1 U20913 ( .A(\mem[76][1] ), .B(\mem[77][1] ), .S(n8367), .Z(n1963) );
  MUX2_X1 U20914 ( .A(n1963), .B(n1962), .S(n8309), .Z(n1964) );
  MUX2_X1 U20915 ( .A(\mem[74][1] ), .B(\mem[75][1] ), .S(n8366), .Z(n1965) );
  MUX2_X1 U20916 ( .A(\mem[72][1] ), .B(\mem[73][1] ), .S(n8373), .Z(n1966) );
  MUX2_X1 U20917 ( .A(n1966), .B(n1965), .S(n8317), .Z(n1967) );
  MUX2_X1 U20918 ( .A(n1967), .B(n1964), .S(n8247), .Z(n1968) );
  MUX2_X1 U20919 ( .A(\mem[70][1] ), .B(\mem[71][1] ), .S(n8366), .Z(n1969) );
  MUX2_X1 U20920 ( .A(\mem[68][1] ), .B(\mem[69][1] ), .S(n8363), .Z(n1970) );
  MUX2_X1 U20921 ( .A(n1970), .B(n1969), .S(n8342), .Z(n1971) );
  MUX2_X1 U20922 ( .A(\mem[66][1] ), .B(\mem[67][1] ), .S(n8364), .Z(n1972) );
  MUX2_X1 U20923 ( .A(\mem[64][1] ), .B(\mem[65][1] ), .S(n8539), .Z(n1973) );
  MUX2_X1 U20924 ( .A(n1973), .B(n1972), .S(n8334), .Z(n1974) );
  MUX2_X1 U20925 ( .A(n1974), .B(n1971), .S(n8247), .Z(n1975) );
  MUX2_X1 U20926 ( .A(n1975), .B(n1968), .S(n8201), .Z(n1976) );
  MUX2_X1 U20927 ( .A(n1976), .B(n1961), .S(n8195), .Z(n1977) );
  MUX2_X1 U20928 ( .A(n1977), .B(n1946), .S(n8182), .Z(n1978) );
  MUX2_X1 U20929 ( .A(\mem[62][1] ), .B(\mem[63][1] ), .S(n8362), .Z(n1979) );
  MUX2_X1 U20930 ( .A(\mem[60][1] ), .B(\mem[61][1] ), .S(n8372), .Z(n1980) );
  MUX2_X1 U20931 ( .A(n1980), .B(n1979), .S(n8302), .Z(n1981) );
  MUX2_X1 U20932 ( .A(\mem[58][1] ), .B(\mem[59][1] ), .S(n8371), .Z(n1982) );
  MUX2_X1 U20933 ( .A(\mem[56][1] ), .B(\mem[57][1] ), .S(n8370), .Z(n1983) );
  MUX2_X1 U20934 ( .A(n1983), .B(n1982), .S(n8310), .Z(n1984) );
  MUX2_X1 U20935 ( .A(n1984), .B(n1981), .S(n8247), .Z(n1985) );
  MUX2_X1 U20936 ( .A(\mem[54][1] ), .B(\mem[55][1] ), .S(n8369), .Z(n1986) );
  MUX2_X1 U20937 ( .A(\mem[52][1] ), .B(\mem[53][1] ), .S(n8368), .Z(n1987) );
  MUX2_X1 U20938 ( .A(n1987), .B(n1986), .S(n8344), .Z(n1988) );
  MUX2_X1 U20939 ( .A(\mem[50][1] ), .B(\mem[51][1] ), .S(n8367), .Z(n1989) );
  MUX2_X1 U20940 ( .A(\mem[48][1] ), .B(\mem[49][1] ), .S(n8366), .Z(n1990) );
  MUX2_X1 U20941 ( .A(n1990), .B(n1989), .S(n8273), .Z(n1991) );
  MUX2_X1 U20942 ( .A(n1991), .B(n1988), .S(n8247), .Z(n1992) );
  MUX2_X1 U20943 ( .A(n1992), .B(n1985), .S(N21), .Z(n1993) );
  MUX2_X1 U20944 ( .A(\mem[46][1] ), .B(\mem[47][1] ), .S(n8512), .Z(n1994) );
  MUX2_X1 U20945 ( .A(\mem[44][1] ), .B(\mem[45][1] ), .S(n8507), .Z(n1995) );
  MUX2_X1 U20946 ( .A(n1995), .B(n1994), .S(n8325), .Z(n1996) );
  MUX2_X1 U20947 ( .A(\mem[42][1] ), .B(\mem[43][1] ), .S(n8508), .Z(n1997) );
  MUX2_X1 U20948 ( .A(\mem[40][1] ), .B(\mem[41][1] ), .S(n8509), .Z(n1998) );
  MUX2_X1 U20949 ( .A(n1998), .B(n1997), .S(n8323), .Z(n1999) );
  MUX2_X1 U20950 ( .A(n1999), .B(n1996), .S(n8247), .Z(n2000) );
  MUX2_X1 U20951 ( .A(\mem[38][1] ), .B(\mem[39][1] ), .S(n8516), .Z(n2001) );
  MUX2_X1 U20952 ( .A(\mem[36][1] ), .B(\mem[37][1] ), .S(n8517), .Z(n2002) );
  MUX2_X1 U20953 ( .A(n2002), .B(n2001), .S(n8303), .Z(n2003) );
  MUX2_X1 U20954 ( .A(\mem[34][1] ), .B(\mem[35][1] ), .S(n8518), .Z(n2004) );
  MUX2_X1 U20955 ( .A(\mem[32][1] ), .B(\mem[33][1] ), .S(n8513), .Z(n2005) );
  MUX2_X1 U20956 ( .A(n2005), .B(n2004), .S(n8333), .Z(n2006) );
  MUX2_X1 U20957 ( .A(n2006), .B(n2003), .S(n8247), .Z(n2007) );
  MUX2_X1 U20958 ( .A(n2007), .B(n2000), .S(n8199), .Z(n2008) );
  MUX2_X1 U20959 ( .A(n2008), .B(n1993), .S(n8196), .Z(n2009) );
  MUX2_X1 U20960 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n8514), .Z(n2010) );
  MUX2_X1 U20961 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n8515), .Z(n2011) );
  MUX2_X1 U20962 ( .A(n2011), .B(n2010), .S(n8278), .Z(n2012) );
  MUX2_X1 U20963 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n8522), .Z(n2013) );
  MUX2_X1 U20964 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n8523), .Z(n2014) );
  MUX2_X1 U20965 ( .A(n2014), .B(n2013), .S(n8349), .Z(n2015) );
  MUX2_X1 U20966 ( .A(n2015), .B(n2012), .S(n8247), .Z(n2016) );
  MUX2_X1 U20967 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n8500), .Z(n2017) );
  MUX2_X1 U20968 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n8495), .Z(n2018) );
  MUX2_X1 U20969 ( .A(n2018), .B(n2017), .S(n8334), .Z(n2019) );
  MUX2_X1 U20970 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n8496), .Z(n2020) );
  MUX2_X1 U20971 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n8497), .Z(n2021) );
  MUX2_X1 U20972 ( .A(n2021), .B(n2020), .S(n8283), .Z(n2022) );
  MUX2_X1 U20973 ( .A(n2022), .B(n2019), .S(n8247), .Z(n2023) );
  MUX2_X1 U20974 ( .A(n2023), .B(n2016), .S(n8207), .Z(n2024) );
  MUX2_X1 U20975 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n8504), .Z(n2025) );
  MUX2_X1 U20976 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n8505), .Z(n2026) );
  MUX2_X1 U20977 ( .A(n2026), .B(n2025), .S(n8320), .Z(n2027) );
  MUX2_X1 U20978 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n8506), .Z(n2028) );
  MUX2_X1 U20979 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n8501), .Z(n2029) );
  MUX2_X1 U20980 ( .A(n2029), .B(n2028), .S(n8282), .Z(n2030) );
  MUX2_X1 U20981 ( .A(n2030), .B(n2027), .S(n8247), .Z(n2031) );
  MUX2_X1 U20982 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n8502), .Z(n2032) );
  MUX2_X1 U20983 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n8503), .Z(n2033) );
  MUX2_X1 U20984 ( .A(n2033), .B(n2032), .S(n8329), .Z(n2034) );
  MUX2_X1 U20985 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n8510), .Z(n2035) );
  MUX2_X1 U20986 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n8511), .Z(n2036) );
  MUX2_X1 U20987 ( .A(n2036), .B(n2035), .S(n8296), .Z(n2037) );
  MUX2_X1 U20988 ( .A(n2037), .B(n2034), .S(n8247), .Z(n2038) );
  MUX2_X1 U20989 ( .A(n2038), .B(n2031), .S(n8197), .Z(n2039) );
  MUX2_X1 U20990 ( .A(n2039), .B(n2024), .S(n8190), .Z(n2040) );
  MUX2_X1 U20991 ( .A(n2040), .B(n2009), .S(n8182), .Z(n2041) );
  MUX2_X1 U20992 ( .A(n2041), .B(n1978), .S(n8179), .Z(n2042) );
  MUX2_X1 U20993 ( .A(n2042), .B(n1915), .S(n8177), .Z(n2043) );
  MUX2_X1 U20994 ( .A(n2043), .B(n1788), .S(N26), .Z(n2044) );
  MUX2_X1 U20995 ( .A(n2044), .B(n1533), .S(N27), .Z(N34) );
  MUX2_X1 U20996 ( .A(\mem[1022][2] ), .B(\mem[1023][2] ), .S(n8488), .Z(n2045) );
  MUX2_X1 U20997 ( .A(\mem[1020][2] ), .B(\mem[1021][2] ), .S(n8483), .Z(n2046) );
  MUX2_X1 U20998 ( .A(n2046), .B(n2045), .S(n8287), .Z(n2047) );
  MUX2_X1 U20999 ( .A(\mem[1018][2] ), .B(\mem[1019][2] ), .S(n8484), .Z(n2048) );
  MUX2_X1 U21000 ( .A(\mem[1016][2] ), .B(\mem[1017][2] ), .S(n8485), .Z(n2049) );
  MUX2_X1 U21001 ( .A(n2049), .B(n2048), .S(n8349), .Z(n2050) );
  MUX2_X1 U21002 ( .A(n2050), .B(n2047), .S(n8248), .Z(n2051) );
  MUX2_X1 U21003 ( .A(\mem[1014][2] ), .B(\mem[1015][2] ), .S(n8492), .Z(n2052) );
  MUX2_X1 U21004 ( .A(\mem[1012][2] ), .B(\mem[1013][2] ), .S(n8493), .Z(n2053) );
  MUX2_X1 U21005 ( .A(n2053), .B(n2052), .S(n8335), .Z(n2054) );
  MUX2_X1 U21006 ( .A(\mem[1010][2] ), .B(\mem[1011][2] ), .S(n8494), .Z(n2055) );
  MUX2_X1 U21007 ( .A(\mem[1008][2] ), .B(\mem[1009][2] ), .S(n8489), .Z(n2056) );
  MUX2_X1 U21008 ( .A(n2056), .B(n2055), .S(n8326), .Z(n2057) );
  MUX2_X1 U21009 ( .A(n2057), .B(n2054), .S(n8248), .Z(n2058) );
  MUX2_X1 U21010 ( .A(n2058), .B(n2051), .S(n8219), .Z(n2059) );
  MUX2_X1 U21011 ( .A(\mem[1006][2] ), .B(\mem[1007][2] ), .S(n8490), .Z(n2060) );
  MUX2_X1 U21012 ( .A(\mem[1004][2] ), .B(\mem[1005][2] ), .S(n8491), .Z(n2061) );
  MUX2_X1 U21013 ( .A(n2061), .B(n2060), .S(n8306), .Z(n2062) );
  MUX2_X1 U21014 ( .A(\mem[1002][2] ), .B(\mem[1003][2] ), .S(n8498), .Z(n2063) );
  MUX2_X1 U21015 ( .A(\mem[1000][2] ), .B(\mem[1001][2] ), .S(n8499), .Z(n2064) );
  MUX2_X1 U21016 ( .A(n2064), .B(n2063), .S(n8271), .Z(n2065) );
  MUX2_X1 U21017 ( .A(n2065), .B(n2062), .S(n8248), .Z(n2066) );
  MUX2_X1 U21018 ( .A(\mem[998][2] ), .B(\mem[999][2] ), .S(n8508), .Z(n2067)
         );
  MUX2_X1 U21019 ( .A(\mem[996][2] ), .B(\mem[997][2] ), .S(n8398), .Z(n2068)
         );
  MUX2_X1 U21020 ( .A(n2068), .B(n2067), .S(n8285), .Z(n2069) );
  MUX2_X1 U21021 ( .A(\mem[994][2] ), .B(\mem[995][2] ), .S(n8425), .Z(n2070)
         );
  MUX2_X1 U21022 ( .A(\mem[992][2] ), .B(\mem[993][2] ), .S(n8403), .Z(n2071)
         );
  MUX2_X1 U21023 ( .A(n2071), .B(n2070), .S(n8272), .Z(n2072) );
  MUX2_X1 U21024 ( .A(n2072), .B(n2069), .S(n8248), .Z(n2073) );
  MUX2_X1 U21025 ( .A(n2073), .B(n2066), .S(n8217), .Z(n2074) );
  MUX2_X1 U21026 ( .A(n2074), .B(n2059), .S(n8188), .Z(n2075) );
  MUX2_X1 U21027 ( .A(\mem[990][2] ), .B(\mem[991][2] ), .S(n8525), .Z(n2076)
         );
  MUX2_X1 U21028 ( .A(\mem[988][2] ), .B(\mem[989][2] ), .S(n8449), .Z(n2077)
         );
  MUX2_X1 U21029 ( .A(n2077), .B(n2076), .S(n8267), .Z(n2078) );
  MUX2_X1 U21030 ( .A(\mem[986][2] ), .B(\mem[987][2] ), .S(n8521), .Z(n2079)
         );
  MUX2_X1 U21031 ( .A(\mem[984][2] ), .B(\mem[985][2] ), .S(n8504), .Z(n2080)
         );
  MUX2_X1 U21032 ( .A(n2080), .B(n2079), .S(n8306), .Z(n2081) );
  MUX2_X1 U21033 ( .A(n2081), .B(n2078), .S(n8248), .Z(n2082) );
  MUX2_X1 U21034 ( .A(\mem[982][2] ), .B(\mem[983][2] ), .S(n8385), .Z(n2083)
         );
  MUX2_X1 U21035 ( .A(\mem[980][2] ), .B(\mem[981][2] ), .S(n8384), .Z(n2084)
         );
  MUX2_X1 U21036 ( .A(n2084), .B(n2083), .S(n8342), .Z(n2085) );
  MUX2_X1 U21037 ( .A(\mem[978][2] ), .B(\mem[979][2] ), .S(n8383), .Z(n2086)
         );
  MUX2_X1 U21038 ( .A(\mem[976][2] ), .B(\mem[977][2] ), .S(n8382), .Z(n2087)
         );
  MUX2_X1 U21039 ( .A(n2087), .B(n2086), .S(n8266), .Z(n2088) );
  MUX2_X1 U21040 ( .A(n2088), .B(n2085), .S(n8248), .Z(n2089) );
  MUX2_X1 U21041 ( .A(n2089), .B(n2082), .S(n8219), .Z(n2090) );
  MUX2_X1 U21042 ( .A(\mem[974][2] ), .B(\mem[975][2] ), .S(n8380), .Z(n2091)
         );
  MUX2_X1 U21043 ( .A(\mem[972][2] ), .B(\mem[973][2] ), .S(n8535), .Z(n2092)
         );
  MUX2_X1 U21044 ( .A(n2092), .B(n2091), .S(n8296), .Z(n2093) );
  MUX2_X1 U21045 ( .A(\mem[970][2] ), .B(\mem[971][2] ), .S(n8524), .Z(n2094)
         );
  MUX2_X1 U21046 ( .A(\mem[968][2] ), .B(\mem[969][2] ), .S(n8429), .Z(n2095)
         );
  MUX2_X1 U21047 ( .A(n2095), .B(n2094), .S(n8297), .Z(n2096) );
  MUX2_X1 U21048 ( .A(n2096), .B(n2093), .S(n8248), .Z(n2097) );
  MUX2_X1 U21049 ( .A(\mem[966][2] ), .B(\mem[967][2] ), .S(n8460), .Z(n2098)
         );
  MUX2_X1 U21050 ( .A(\mem[964][2] ), .B(\mem[965][2] ), .S(n8416), .Z(n2099)
         );
  MUX2_X1 U21051 ( .A(n2099), .B(n2098), .S(n8298), .Z(n2100) );
  MUX2_X1 U21052 ( .A(\mem[962][2] ), .B(\mem[963][2] ), .S(n8370), .Z(n2101)
         );
  MUX2_X1 U21053 ( .A(\mem[960][2] ), .B(\mem[961][2] ), .S(n8463), .Z(n2102)
         );
  MUX2_X1 U21054 ( .A(n2102), .B(n2101), .S(n8293), .Z(n2103) );
  MUX2_X1 U21055 ( .A(n2103), .B(n2100), .S(n8248), .Z(n2104) );
  MUX2_X1 U21056 ( .A(n2104), .B(n2097), .S(n8197), .Z(n2105) );
  MUX2_X1 U21057 ( .A(n2105), .B(n2090), .S(n8190), .Z(n2106) );
  MUX2_X1 U21058 ( .A(n2106), .B(n2075), .S(n8183), .Z(n2107) );
  MUX2_X1 U21059 ( .A(\mem[958][2] ), .B(\mem[959][2] ), .S(n8493), .Z(n2108)
         );
  MUX2_X1 U21060 ( .A(\mem[956][2] ), .B(\mem[957][2] ), .S(n8449), .Z(n2109)
         );
  MUX2_X1 U21061 ( .A(n2109), .B(n2108), .S(n8294), .Z(n2110) );
  MUX2_X1 U21062 ( .A(\mem[954][2] ), .B(\mem[955][2] ), .S(n8459), .Z(n2111)
         );
  MUX2_X1 U21063 ( .A(\mem[952][2] ), .B(\mem[953][2] ), .S(n8421), .Z(n2112)
         );
  MUX2_X1 U21064 ( .A(n2112), .B(n2111), .S(n8295), .Z(n2113) );
  MUX2_X1 U21065 ( .A(n2113), .B(n2110), .S(n8248), .Z(n2114) );
  MUX2_X1 U21066 ( .A(\mem[950][2] ), .B(\mem[951][2] ), .S(n8519), .Z(n2115)
         );
  MUX2_X1 U21067 ( .A(\mem[948][2] ), .B(\mem[949][2] ), .S(n8520), .Z(n2116)
         );
  MUX2_X1 U21068 ( .A(n2116), .B(n2115), .S(n8302), .Z(n2117) );
  MUX2_X1 U21069 ( .A(\mem[946][2] ), .B(\mem[947][2] ), .S(n8521), .Z(n2118)
         );
  MUX2_X1 U21070 ( .A(\mem[944][2] ), .B(\mem[945][2] ), .S(n8528), .Z(n2119)
         );
  MUX2_X1 U21071 ( .A(n2119), .B(n2118), .S(n8303), .Z(n2120) );
  MUX2_X1 U21072 ( .A(n2120), .B(n2117), .S(n8248), .Z(n2121) );
  MUX2_X1 U21073 ( .A(n2121), .B(n2114), .S(n8200), .Z(n2122) );
  MUX2_X1 U21074 ( .A(\mem[942][2] ), .B(\mem[943][2] ), .S(n8529), .Z(n2123)
         );
  MUX2_X1 U21075 ( .A(\mem[940][2] ), .B(\mem[941][2] ), .S(n8530), .Z(n2124)
         );
  MUX2_X1 U21076 ( .A(n2124), .B(n2123), .S(n8304), .Z(n2125) );
  MUX2_X1 U21077 ( .A(\mem[938][2] ), .B(\mem[939][2] ), .S(n8371), .Z(n2126)
         );
  MUX2_X1 U21078 ( .A(\mem[936][2] ), .B(\mem[937][2] ), .S(n8366), .Z(n2127)
         );
  MUX2_X1 U21079 ( .A(n2127), .B(n2126), .S(n8299), .Z(n2128) );
  MUX2_X1 U21080 ( .A(n2128), .B(n2125), .S(n8248), .Z(n2129) );
  MUX2_X1 U21081 ( .A(\mem[934][2] ), .B(\mem[935][2] ), .S(n8410), .Z(n2130)
         );
  MUX2_X1 U21082 ( .A(\mem[932][2] ), .B(\mem[933][2] ), .S(n8427), .Z(n2131)
         );
  MUX2_X1 U21083 ( .A(n2131), .B(n2130), .S(n8300), .Z(n2132) );
  MUX2_X1 U21084 ( .A(\mem[930][2] ), .B(\mem[931][2] ), .S(n8361), .Z(n2133)
         );
  MUX2_X1 U21085 ( .A(\mem[928][2] ), .B(\mem[929][2] ), .S(N18), .Z(n2134) );
  MUX2_X1 U21086 ( .A(n2134), .B(n2133), .S(n8301), .Z(n2135) );
  MUX2_X1 U21087 ( .A(n2135), .B(n2132), .S(n8248), .Z(n2136) );
  MUX2_X1 U21088 ( .A(n2136), .B(n2129), .S(n8197), .Z(n2137) );
  MUX2_X1 U21089 ( .A(n2137), .B(n2122), .S(n8186), .Z(n2138) );
  MUX2_X1 U21090 ( .A(\mem[926][2] ), .B(\mem[927][2] ), .S(n8481), .Z(n2139)
         );
  MUX2_X1 U21091 ( .A(\mem[924][2] ), .B(\mem[925][2] ), .S(n8509), .Z(n2140)
         );
  MUX2_X1 U21092 ( .A(n2140), .B(n2139), .S(n8323), .Z(n2141) );
  MUX2_X1 U21093 ( .A(\mem[922][2] ), .B(\mem[923][2] ), .S(n8494), .Z(n2142)
         );
  MUX2_X1 U21094 ( .A(\mem[920][2] ), .B(\mem[921][2] ), .S(n8409), .Z(n2143)
         );
  MUX2_X1 U21095 ( .A(n2143), .B(n2142), .S(n8310), .Z(n2144) );
  MUX2_X1 U21096 ( .A(n2144), .B(n2141), .S(n8249), .Z(n2145) );
  MUX2_X1 U21097 ( .A(\mem[918][2] ), .B(\mem[919][2] ), .S(n8415), .Z(n2146)
         );
  MUX2_X1 U21098 ( .A(\mem[916][2] ), .B(\mem[917][2] ), .S(n8410), .Z(n2147)
         );
  MUX2_X1 U21099 ( .A(n2147), .B(n2146), .S(n8305), .Z(n2148) );
  MUX2_X1 U21100 ( .A(\mem[914][2] ), .B(\mem[915][2] ), .S(n8407), .Z(n2149)
         );
  MUX2_X1 U21101 ( .A(\mem[912][2] ), .B(\mem[913][2] ), .S(n8408), .Z(n2150)
         );
  MUX2_X1 U21102 ( .A(n2150), .B(n2149), .S(n8306), .Z(n2151) );
  MUX2_X1 U21103 ( .A(n2151), .B(n2148), .S(n8249), .Z(n2152) );
  MUX2_X1 U21104 ( .A(n2152), .B(n2145), .S(n8218), .Z(n2153) );
  MUX2_X1 U21105 ( .A(\mem[910][2] ), .B(\mem[911][2] ), .S(n8467), .Z(n2154)
         );
  MUX2_X1 U21106 ( .A(\mem[908][2] ), .B(\mem[909][2] ), .S(n8414), .Z(n2155)
         );
  MUX2_X1 U21107 ( .A(n2155), .B(n2154), .S(n8307), .Z(n2156) );
  MUX2_X1 U21108 ( .A(\mem[906][2] ), .B(\mem[907][2] ), .S(n8415), .Z(n2157)
         );
  MUX2_X1 U21109 ( .A(\mem[904][2] ), .B(\mem[905][2] ), .S(n8416), .Z(n2158)
         );
  MUX2_X1 U21110 ( .A(n2158), .B(n2157), .S(n8314), .Z(n2159) );
  MUX2_X1 U21111 ( .A(n2159), .B(n2156), .S(n8249), .Z(n2160) );
  MUX2_X1 U21112 ( .A(\mem[902][2] ), .B(\mem[903][2] ), .S(n8411), .Z(n2161)
         );
  MUX2_X1 U21113 ( .A(\mem[900][2] ), .B(\mem[901][2] ), .S(n8468), .Z(n2162)
         );
  MUX2_X1 U21114 ( .A(n2162), .B(n2161), .S(n8315), .Z(n2163) );
  MUX2_X1 U21115 ( .A(\mem[898][2] ), .B(\mem[899][2] ), .S(n8431), .Z(n2164)
         );
  MUX2_X1 U21116 ( .A(\mem[896][2] ), .B(\mem[897][2] ), .S(n8433), .Z(n2165)
         );
  MUX2_X1 U21117 ( .A(n2165), .B(n2164), .S(n8316), .Z(n2166) );
  MUX2_X1 U21118 ( .A(n2166), .B(n2163), .S(n8249), .Z(n2167) );
  MUX2_X1 U21119 ( .A(n2167), .B(n2160), .S(n8219), .Z(n2168) );
  MUX2_X1 U21120 ( .A(n2168), .B(n2153), .S(n8191), .Z(n2169) );
  MUX2_X1 U21121 ( .A(n2169), .B(n2138), .S(n8183), .Z(n2170) );
  MUX2_X1 U21122 ( .A(n2170), .B(n2107), .S(n8180), .Z(n2171) );
  MUX2_X1 U21123 ( .A(\mem[894][2] ), .B(\mem[895][2] ), .S(n8370), .Z(n2172)
         );
  MUX2_X1 U21124 ( .A(\mem[892][2] ), .B(\mem[893][2] ), .S(n8460), .Z(n2173)
         );
  MUX2_X1 U21125 ( .A(n2173), .B(n2172), .S(n8311), .Z(n2174) );
  MUX2_X1 U21126 ( .A(\mem[890][2] ), .B(\mem[891][2] ), .S(n8467), .Z(n2175)
         );
  MUX2_X1 U21127 ( .A(\mem[888][2] ), .B(\mem[889][2] ), .S(n8445), .Z(n2176)
         );
  MUX2_X1 U21128 ( .A(n2176), .B(n2175), .S(n8312), .Z(n2177) );
  MUX2_X1 U21129 ( .A(n2177), .B(n2174), .S(n8249), .Z(n2178) );
  MUX2_X1 U21130 ( .A(\mem[886][2] ), .B(\mem[887][2] ), .S(n8531), .Z(n2179)
         );
  MUX2_X1 U21131 ( .A(\mem[884][2] ), .B(\mem[885][2] ), .S(n8357), .Z(n2180)
         );
  MUX2_X1 U21132 ( .A(n2180), .B(n2179), .S(n8313), .Z(n2181) );
  MUX2_X1 U21133 ( .A(\mem[882][2] ), .B(\mem[883][2] ), .S(n8365), .Z(n2182)
         );
  MUX2_X1 U21134 ( .A(\mem[880][2] ), .B(\mem[881][2] ), .S(n8406), .Z(n2183)
         );
  MUX2_X1 U21135 ( .A(n2183), .B(n2182), .S(n8320), .Z(n2184) );
  MUX2_X1 U21136 ( .A(n2184), .B(n2181), .S(n8249), .Z(n2185) );
  MUX2_X1 U21137 ( .A(n2185), .B(n2178), .S(n8197), .Z(n2186) );
  MUX2_X1 U21138 ( .A(\mem[878][2] ), .B(\mem[879][2] ), .S(n8537), .Z(n2187)
         );
  MUX2_X1 U21139 ( .A(\mem[876][2] ), .B(\mem[877][2] ), .S(n8469), .Z(n2188)
         );
  MUX2_X1 U21140 ( .A(n2188), .B(n2187), .S(n8290), .Z(n2189) );
  MUX2_X1 U21141 ( .A(\mem[874][2] ), .B(\mem[875][2] ), .S(n8451), .Z(n2190)
         );
  MUX2_X1 U21142 ( .A(\mem[872][2] ), .B(\mem[873][2] ), .S(n8521), .Z(n2191)
         );
  MUX2_X1 U21143 ( .A(n2191), .B(n2190), .S(n8319), .Z(n2192) );
  MUX2_X1 U21144 ( .A(n2192), .B(n2189), .S(n8249), .Z(n2193) );
  MUX2_X1 U21145 ( .A(\mem[870][2] ), .B(\mem[871][2] ), .S(n8501), .Z(n2194)
         );
  MUX2_X1 U21146 ( .A(\mem[868][2] ), .B(\mem[869][2] ), .S(n8488), .Z(n2195)
         );
  MUX2_X1 U21147 ( .A(n2195), .B(n2194), .S(N19), .Z(n2196) );
  MUX2_X1 U21148 ( .A(\mem[866][2] ), .B(\mem[867][2] ), .S(n8375), .Z(n2197)
         );
  MUX2_X1 U21149 ( .A(\mem[864][2] ), .B(\mem[865][2] ), .S(n8370), .Z(n2198)
         );
  MUX2_X1 U21150 ( .A(n2198), .B(n2197), .S(n8332), .Z(n2199) );
  MUX2_X1 U21151 ( .A(n2199), .B(n2196), .S(n8249), .Z(n2200) );
  MUX2_X1 U21152 ( .A(n2200), .B(n2193), .S(N21), .Z(n2201) );
  MUX2_X1 U21153 ( .A(n2201), .B(n2186), .S(N22), .Z(n2202) );
  MUX2_X1 U21154 ( .A(\mem[862][2] ), .B(\mem[863][2] ), .S(n8393), .Z(n2203)
         );
  MUX2_X1 U21155 ( .A(\mem[860][2] ), .B(\mem[861][2] ), .S(n8511), .Z(n2204)
         );
  MUX2_X1 U21156 ( .A(n2204), .B(n2203), .S(n8342), .Z(n2205) );
  MUX2_X1 U21157 ( .A(\mem[858][2] ), .B(\mem[859][2] ), .S(n8492), .Z(n2206)
         );
  MUX2_X1 U21158 ( .A(\mem[856][2] ), .B(\mem[857][2] ), .S(n8409), .Z(n2207)
         );
  MUX2_X1 U21159 ( .A(n2207), .B(n2206), .S(n8307), .Z(n2208) );
  MUX2_X1 U21160 ( .A(n2208), .B(n2205), .S(n8249), .Z(n2209) );
  MUX2_X1 U21161 ( .A(\mem[854][2] ), .B(\mem[855][2] ), .S(n8437), .Z(n2210)
         );
  MUX2_X1 U21162 ( .A(\mem[852][2] ), .B(\mem[853][2] ), .S(n8444), .Z(n2211)
         );
  MUX2_X1 U21163 ( .A(n2211), .B(n2210), .S(n8289), .Z(n2212) );
  MUX2_X1 U21164 ( .A(\mem[850][2] ), .B(\mem[851][2] ), .S(n8445), .Z(n2213)
         );
  MUX2_X1 U21165 ( .A(\mem[848][2] ), .B(\mem[849][2] ), .S(n8446), .Z(n2214)
         );
  MUX2_X1 U21166 ( .A(n2214), .B(n2213), .S(n8283), .Z(n2215) );
  MUX2_X1 U21167 ( .A(n2215), .B(n2212), .S(n8249), .Z(n2216) );
  MUX2_X1 U21168 ( .A(n2216), .B(n2209), .S(n8197), .Z(n2217) );
  MUX2_X1 U21169 ( .A(\mem[846][2] ), .B(\mem[847][2] ), .S(n8441), .Z(n2218)
         );
  MUX2_X1 U21170 ( .A(\mem[844][2] ), .B(\mem[845][2] ), .S(n8442), .Z(n2219)
         );
  MUX2_X1 U21171 ( .A(n2219), .B(n2218), .S(n8272), .Z(n2220) );
  MUX2_X1 U21172 ( .A(\mem[842][2] ), .B(\mem[843][2] ), .S(n8443), .Z(n2221)
         );
  MUX2_X1 U21173 ( .A(\mem[840][2] ), .B(\mem[841][2] ), .S(n8450), .Z(n2222)
         );
  MUX2_X1 U21174 ( .A(n2222), .B(n2221), .S(n8332), .Z(n2223) );
  MUX2_X1 U21175 ( .A(n2223), .B(n2220), .S(n8249), .Z(n2224) );
  MUX2_X1 U21176 ( .A(\mem[838][2] ), .B(\mem[839][2] ), .S(n8451), .Z(n2225)
         );
  MUX2_X1 U21177 ( .A(\mem[836][2] ), .B(\mem[837][2] ), .S(n8452), .Z(n2226)
         );
  MUX2_X1 U21178 ( .A(n2226), .B(n2225), .S(n8308), .Z(n2227) );
  MUX2_X1 U21179 ( .A(\mem[834][2] ), .B(\mem[835][2] ), .S(n8447), .Z(n2228)
         );
  MUX2_X1 U21180 ( .A(\mem[832][2] ), .B(\mem[833][2] ), .S(n8448), .Z(n2229)
         );
  MUX2_X1 U21181 ( .A(n2229), .B(n2228), .S(n8309), .Z(n2230) );
  MUX2_X1 U21182 ( .A(n2230), .B(n2227), .S(n8249), .Z(n2231) );
  MUX2_X1 U21183 ( .A(n2231), .B(n2224), .S(n8207), .Z(n2232) );
  MUX2_X1 U21184 ( .A(n2232), .B(n2217), .S(n8196), .Z(n2233) );
  MUX2_X1 U21185 ( .A(n2233), .B(n2202), .S(n8183), .Z(n2234) );
  MUX2_X1 U21186 ( .A(\mem[830][2] ), .B(\mem[831][2] ), .S(n8424), .Z(n2235)
         );
  MUX2_X1 U21187 ( .A(\mem[828][2] ), .B(\mem[829][2] ), .S(n8425), .Z(n2236)
         );
  MUX2_X1 U21188 ( .A(n2236), .B(n2235), .S(n8324), .Z(n2237) );
  MUX2_X1 U21189 ( .A(\mem[826][2] ), .B(\mem[827][2] ), .S(n8432), .Z(n2238)
         );
  MUX2_X1 U21190 ( .A(\mem[824][2] ), .B(\mem[825][2] ), .S(n8433), .Z(n2239)
         );
  MUX2_X1 U21191 ( .A(n2239), .B(n2238), .S(n8308), .Z(n2240) );
  MUX2_X1 U21192 ( .A(n2240), .B(n2237), .S(n8250), .Z(n2241) );
  MUX2_X1 U21193 ( .A(\mem[822][2] ), .B(\mem[823][2] ), .S(n8434), .Z(n2242)
         );
  MUX2_X1 U21194 ( .A(\mem[820][2] ), .B(\mem[821][2] ), .S(n8429), .Z(n2243)
         );
  MUX2_X1 U21195 ( .A(n2243), .B(n2242), .S(n8335), .Z(n2244) );
  MUX2_X1 U21196 ( .A(\mem[818][2] ), .B(\mem[819][2] ), .S(n8430), .Z(n2245)
         );
  MUX2_X1 U21197 ( .A(\mem[816][2] ), .B(\mem[817][2] ), .S(n8431), .Z(n2246)
         );
  MUX2_X1 U21198 ( .A(n2246), .B(n2245), .S(n8302), .Z(n2247) );
  MUX2_X1 U21199 ( .A(n2247), .B(n2244), .S(n8250), .Z(n2248) );
  MUX2_X1 U21200 ( .A(n2248), .B(n2241), .S(n8198), .Z(n2249) );
  MUX2_X1 U21201 ( .A(\mem[814][2] ), .B(\mem[815][2] ), .S(n8438), .Z(n2250)
         );
  MUX2_X1 U21202 ( .A(\mem[812][2] ), .B(\mem[813][2] ), .S(n8439), .Z(n2251)
         );
  MUX2_X1 U21203 ( .A(n2251), .B(n2250), .S(n8267), .Z(n2252) );
  MUX2_X1 U21204 ( .A(\mem[810][2] ), .B(\mem[811][2] ), .S(n8440), .Z(n2253)
         );
  MUX2_X1 U21205 ( .A(\mem[808][2] ), .B(\mem[809][2] ), .S(n8435), .Z(n2254)
         );
  MUX2_X1 U21206 ( .A(n2254), .B(n2253), .S(n8284), .Z(n2255) );
  MUX2_X1 U21207 ( .A(n2255), .B(n2252), .S(n8250), .Z(n2256) );
  MUX2_X1 U21208 ( .A(\mem[806][2] ), .B(\mem[807][2] ), .S(n8412), .Z(n2257)
         );
  MUX2_X1 U21209 ( .A(\mem[804][2] ), .B(\mem[805][2] ), .S(n8413), .Z(n2258)
         );
  MUX2_X1 U21210 ( .A(n2258), .B(n2257), .S(n8285), .Z(n2259) );
  MUX2_X1 U21211 ( .A(\mem[802][2] ), .B(\mem[803][2] ), .S(n8420), .Z(n2260)
         );
  MUX2_X1 U21212 ( .A(\mem[800][2] ), .B(\mem[801][2] ), .S(n8421), .Z(n2261)
         );
  MUX2_X1 U21213 ( .A(n2261), .B(n2260), .S(n8286), .Z(n2262) );
  MUX2_X1 U21214 ( .A(n2262), .B(n2259), .S(n8250), .Z(n2263) );
  MUX2_X1 U21215 ( .A(n2263), .B(n2256), .S(n8211), .Z(n2264) );
  MUX2_X1 U21216 ( .A(n2264), .B(n2249), .S(n8195), .Z(n2265) );
  MUX2_X1 U21217 ( .A(\mem[798][2] ), .B(\mem[799][2] ), .S(n8422), .Z(n2266)
         );
  MUX2_X1 U21218 ( .A(\mem[796][2] ), .B(\mem[797][2] ), .S(n8417), .Z(n2267)
         );
  MUX2_X1 U21219 ( .A(n2267), .B(n2266), .S(n8349), .Z(n2268) );
  MUX2_X1 U21220 ( .A(\mem[794][2] ), .B(\mem[795][2] ), .S(n8418), .Z(n2269)
         );
  MUX2_X1 U21221 ( .A(\mem[792][2] ), .B(\mem[793][2] ), .S(n8419), .Z(n2270)
         );
  MUX2_X1 U21222 ( .A(n2270), .B(n2269), .S(n8296), .Z(n2271) );
  MUX2_X1 U21223 ( .A(n2271), .B(n2268), .S(n8250), .Z(n2272) );
  MUX2_X1 U21224 ( .A(\mem[790][2] ), .B(\mem[791][2] ), .S(n8426), .Z(n2273)
         );
  MUX2_X1 U21225 ( .A(\mem[788][2] ), .B(\mem[789][2] ), .S(n8427), .Z(n2274)
         );
  MUX2_X1 U21226 ( .A(n2274), .B(n2273), .S(n8351), .Z(n2275) );
  MUX2_X1 U21227 ( .A(\mem[786][2] ), .B(\mem[787][2] ), .S(n8428), .Z(n2276)
         );
  MUX2_X1 U21228 ( .A(\mem[784][2] ), .B(\mem[785][2] ), .S(n8423), .Z(n2277)
         );
  MUX2_X1 U21229 ( .A(n2277), .B(n2276), .S(n8277), .Z(n2278) );
  MUX2_X1 U21230 ( .A(n2278), .B(n2275), .S(n8250), .Z(n2279) );
  MUX2_X1 U21231 ( .A(n2279), .B(n2272), .S(n8212), .Z(n2280) );
  MUX2_X1 U21232 ( .A(\mem[782][2] ), .B(\mem[783][2] ), .S(n8359), .Z(n2281)
         );
  MUX2_X1 U21233 ( .A(\mem[780][2] ), .B(\mem[781][2] ), .S(n8378), .Z(n2282)
         );
  MUX2_X1 U21234 ( .A(n2282), .B(n2281), .S(n8289), .Z(n2283) );
  MUX2_X1 U21235 ( .A(\mem[778][2] ), .B(\mem[779][2] ), .S(N18), .Z(n2284) );
  MUX2_X1 U21236 ( .A(\mem[776][2] ), .B(\mem[777][2] ), .S(n8408), .Z(n2285)
         );
  MUX2_X1 U21237 ( .A(n2285), .B(n2284), .S(n8281), .Z(n2286) );
  MUX2_X1 U21238 ( .A(n2286), .B(n2283), .S(n8250), .Z(n2287) );
  MUX2_X1 U21239 ( .A(\mem[774][2] ), .B(\mem[775][2] ), .S(n8367), .Z(n2288)
         );
  MUX2_X1 U21240 ( .A(\mem[772][2] ), .B(\mem[773][2] ), .S(n8453), .Z(n2289)
         );
  MUX2_X1 U21241 ( .A(n2289), .B(n2288), .S(n8274), .Z(n2290) );
  MUX2_X1 U21242 ( .A(\mem[770][2] ), .B(\mem[771][2] ), .S(n8402), .Z(n2291)
         );
  MUX2_X1 U21243 ( .A(\mem[768][2] ), .B(\mem[769][2] ), .S(n8418), .Z(n2292)
         );
  MUX2_X1 U21244 ( .A(n2292), .B(n2291), .S(n8354), .Z(n2293) );
  MUX2_X1 U21245 ( .A(n2293), .B(n2290), .S(n8250), .Z(n2294) );
  MUX2_X1 U21246 ( .A(n2294), .B(n2287), .S(n8214), .Z(n2295) );
  MUX2_X1 U21247 ( .A(n2295), .B(n2280), .S(n8192), .Z(n2296) );
  MUX2_X1 U21248 ( .A(n2296), .B(n2265), .S(n8183), .Z(n2297) );
  MUX2_X1 U21249 ( .A(n2297), .B(n2234), .S(n8178), .Z(n2298) );
  MUX2_X1 U21250 ( .A(n2298), .B(n2171), .S(n8177), .Z(n2299) );
  MUX2_X1 U21251 ( .A(\mem[766][2] ), .B(\mem[767][2] ), .S(n8464), .Z(n2300)
         );
  MUX2_X1 U21252 ( .A(\mem[764][2] ), .B(\mem[765][2] ), .S(n8414), .Z(n2301)
         );
  MUX2_X1 U21253 ( .A(n2301), .B(n2300), .S(n8342), .Z(n2302) );
  MUX2_X1 U21254 ( .A(\mem[762][2] ), .B(\mem[763][2] ), .S(n8413), .Z(n2303)
         );
  MUX2_X1 U21255 ( .A(\mem[760][2] ), .B(\mem[761][2] ), .S(n8403), .Z(n2304)
         );
  MUX2_X1 U21256 ( .A(n2304), .B(n2303), .S(n8305), .Z(n2305) );
  MUX2_X1 U21257 ( .A(n2305), .B(n2302), .S(n8250), .Z(n2306) );
  MUX2_X1 U21258 ( .A(\mem[758][2] ), .B(\mem[759][2] ), .S(n8404), .Z(n2307)
         );
  MUX2_X1 U21259 ( .A(\mem[756][2] ), .B(\mem[757][2] ), .S(n8525), .Z(n2308)
         );
  MUX2_X1 U21260 ( .A(n2308), .B(n2307), .S(n8282), .Z(n2309) );
  MUX2_X1 U21261 ( .A(\mem[754][2] ), .B(\mem[755][2] ), .S(n8509), .Z(n2310)
         );
  MUX2_X1 U21262 ( .A(\mem[752][2] ), .B(\mem[753][2] ), .S(n8500), .Z(n2311)
         );
  MUX2_X1 U21263 ( .A(n2311), .B(n2310), .S(n8321), .Z(n2312) );
  MUX2_X1 U21264 ( .A(n2312), .B(n2309), .S(n8250), .Z(n2313) );
  MUX2_X1 U21265 ( .A(n2313), .B(n2306), .S(n8201), .Z(n2314) );
  MUX2_X1 U21266 ( .A(\mem[750][2] ), .B(\mem[751][2] ), .S(n8425), .Z(n2315)
         );
  MUX2_X1 U21267 ( .A(\mem[748][2] ), .B(\mem[749][2] ), .S(n8414), .Z(n2316)
         );
  MUX2_X1 U21268 ( .A(n2316), .B(n2315), .S(n8300), .Z(n2317) );
  MUX2_X1 U21269 ( .A(\mem[746][2] ), .B(\mem[747][2] ), .S(n8529), .Z(n2318)
         );
  MUX2_X1 U21270 ( .A(\mem[744][2] ), .B(\mem[745][2] ), .S(n8508), .Z(n2319)
         );
  MUX2_X1 U21271 ( .A(n2319), .B(n2318), .S(n8344), .Z(n2320) );
  MUX2_X1 U21272 ( .A(n2320), .B(n2317), .S(n8250), .Z(n2321) );
  MUX2_X1 U21273 ( .A(\mem[742][2] ), .B(\mem[743][2] ), .S(n8498), .Z(n2322)
         );
  MUX2_X1 U21274 ( .A(\mem[740][2] ), .B(\mem[741][2] ), .S(n8482), .Z(n2323)
         );
  MUX2_X1 U21275 ( .A(n2323), .B(n2322), .S(n8281), .Z(n2324) );
  MUX2_X1 U21276 ( .A(\mem[738][2] ), .B(\mem[739][2] ), .S(n8500), .Z(n2325)
         );
  MUX2_X1 U21277 ( .A(\mem[736][2] ), .B(\mem[737][2] ), .S(n8450), .Z(n2326)
         );
  MUX2_X1 U21278 ( .A(n2326), .B(n2325), .S(n8280), .Z(n2327) );
  MUX2_X1 U21279 ( .A(n2327), .B(n2324), .S(n8250), .Z(n2328) );
  MUX2_X1 U21280 ( .A(n2328), .B(n2321), .S(n8211), .Z(n2329) );
  MUX2_X1 U21281 ( .A(n2329), .B(n2314), .S(n8193), .Z(n2330) );
  MUX2_X1 U21282 ( .A(\mem[734][2] ), .B(\mem[735][2] ), .S(n8452), .Z(n2331)
         );
  MUX2_X1 U21283 ( .A(\mem[732][2] ), .B(\mem[733][2] ), .S(n8529), .Z(n2332)
         );
  MUX2_X1 U21284 ( .A(n2332), .B(n2331), .S(n8356), .Z(n2333) );
  MUX2_X1 U21285 ( .A(\mem[730][2] ), .B(\mem[731][2] ), .S(n8479), .Z(n2334)
         );
  MUX2_X1 U21286 ( .A(\mem[728][2] ), .B(\mem[729][2] ), .S(n8401), .Z(n2335)
         );
  MUX2_X1 U21287 ( .A(n2335), .B(n2334), .S(n8342), .Z(n2336) );
  MUX2_X1 U21288 ( .A(n2336), .B(n2333), .S(n8251), .Z(n2337) );
  MUX2_X1 U21289 ( .A(\mem[726][2] ), .B(\mem[727][2] ), .S(n8389), .Z(n2338)
         );
  MUX2_X1 U21290 ( .A(\mem[724][2] ), .B(\mem[725][2] ), .S(n8357), .Z(n2339)
         );
  MUX2_X1 U21291 ( .A(n2339), .B(n2338), .S(n8341), .Z(n2340) );
  MUX2_X1 U21292 ( .A(\mem[722][2] ), .B(\mem[723][2] ), .S(n8402), .Z(n2341)
         );
  MUX2_X1 U21293 ( .A(\mem[720][2] ), .B(\mem[721][2] ), .S(n8534), .Z(n2342)
         );
  MUX2_X1 U21294 ( .A(n2342), .B(n2341), .S(n8266), .Z(n2343) );
  MUX2_X1 U21295 ( .A(n2343), .B(n2340), .S(n8251), .Z(n2344) );
  MUX2_X1 U21296 ( .A(n2344), .B(n2337), .S(n8212), .Z(n2345) );
  MUX2_X1 U21297 ( .A(\mem[718][2] ), .B(\mem[719][2] ), .S(n8401), .Z(n2346)
         );
  MUX2_X1 U21298 ( .A(\mem[716][2] ), .B(\mem[717][2] ), .S(n8357), .Z(n2347)
         );
  MUX2_X1 U21299 ( .A(n2347), .B(n2346), .S(n8267), .Z(n2348) );
  MUX2_X1 U21300 ( .A(\mem[714][2] ), .B(\mem[715][2] ), .S(n8365), .Z(n2349)
         );
  MUX2_X1 U21301 ( .A(\mem[712][2] ), .B(\mem[713][2] ), .S(n8386), .Z(n2350)
         );
  MUX2_X1 U21302 ( .A(n2350), .B(n2349), .S(n8277), .Z(n2351) );
  MUX2_X1 U21303 ( .A(n2351), .B(n2348), .S(n8251), .Z(n2352) );
  MUX2_X1 U21304 ( .A(\mem[710][2] ), .B(\mem[711][2] ), .S(n8526), .Z(n2353)
         );
  MUX2_X1 U21305 ( .A(\mem[708][2] ), .B(\mem[709][2] ), .S(n8527), .Z(n2354)
         );
  MUX2_X1 U21306 ( .A(n2354), .B(n2353), .S(n8295), .Z(n2355) );
  MUX2_X1 U21307 ( .A(\mem[706][2] ), .B(\mem[707][2] ), .S(n8433), .Z(n2356)
         );
  MUX2_X1 U21308 ( .A(\mem[704][2] ), .B(\mem[705][2] ), .S(n8420), .Z(n2357)
         );
  MUX2_X1 U21309 ( .A(n2357), .B(n2356), .S(n8332), .Z(n2358) );
  MUX2_X1 U21310 ( .A(n2358), .B(n2355), .S(n8251), .Z(n2359) );
  MUX2_X1 U21311 ( .A(n2359), .B(n2352), .S(n8202), .Z(n2360) );
  MUX2_X1 U21312 ( .A(n2360), .B(n2345), .S(n8189), .Z(n2361) );
  MUX2_X1 U21313 ( .A(n2361), .B(n2330), .S(n8183), .Z(n2362) );
  MUX2_X1 U21314 ( .A(\mem[702][2] ), .B(\mem[703][2] ), .S(n8358), .Z(n2363)
         );
  MUX2_X1 U21315 ( .A(\mem[700][2] ), .B(\mem[701][2] ), .S(n8538), .Z(n2364)
         );
  MUX2_X1 U21316 ( .A(n2364), .B(n2363), .S(n8290), .Z(n2365) );
  MUX2_X1 U21317 ( .A(\mem[698][2] ), .B(\mem[699][2] ), .S(n8359), .Z(n2366)
         );
  MUX2_X1 U21318 ( .A(\mem[696][2] ), .B(\mem[697][2] ), .S(n8360), .Z(n2367)
         );
  MUX2_X1 U21319 ( .A(n2367), .B(n2366), .S(n8291), .Z(n2368) );
  MUX2_X1 U21320 ( .A(n2368), .B(n2365), .S(n8251), .Z(n2369) );
  MUX2_X1 U21321 ( .A(\mem[694][2] ), .B(\mem[695][2] ), .S(n8361), .Z(n2370)
         );
  MUX2_X1 U21322 ( .A(\mem[692][2] ), .B(\mem[693][2] ), .S(n8362), .Z(n2371)
         );
  MUX2_X1 U21323 ( .A(n2371), .B(n2370), .S(n8292), .Z(n2372) );
  MUX2_X1 U21324 ( .A(\mem[690][2] ), .B(\mem[691][2] ), .S(n8407), .Z(n2373)
         );
  MUX2_X1 U21325 ( .A(\mem[688][2] ), .B(\mem[689][2] ), .S(n8538), .Z(n2374)
         );
  MUX2_X1 U21326 ( .A(n2374), .B(n2373), .S(n8287), .Z(n2375) );
  MUX2_X1 U21327 ( .A(n2375), .B(n2372), .S(n8251), .Z(n2376) );
  MUX2_X1 U21328 ( .A(n2376), .B(n2369), .S(n8203), .Z(n2377) );
  MUX2_X1 U21329 ( .A(\mem[686][2] ), .B(\mem[687][2] ), .S(n8383), .Z(n2378)
         );
  MUX2_X1 U21330 ( .A(\mem[684][2] ), .B(\mem[685][2] ), .S(n8373), .Z(n2379)
         );
  MUX2_X1 U21331 ( .A(n2379), .B(n2378), .S(n8297), .Z(n2380) );
  MUX2_X1 U21332 ( .A(\mem[682][2] ), .B(\mem[683][2] ), .S(n8371), .Z(n2381)
         );
  MUX2_X1 U21333 ( .A(\mem[680][2] ), .B(\mem[681][2] ), .S(n8370), .Z(n2382)
         );
  MUX2_X1 U21334 ( .A(n2382), .B(n2381), .S(n8298), .Z(n2383) );
  MUX2_X1 U21335 ( .A(n2383), .B(n2380), .S(n8251), .Z(n2384) );
  MUX2_X1 U21336 ( .A(\mem[678][2] ), .B(\mem[679][2] ), .S(n8376), .Z(n2385)
         );
  MUX2_X1 U21337 ( .A(\mem[676][2] ), .B(\mem[677][2] ), .S(n8382), .Z(n2386)
         );
  MUX2_X1 U21338 ( .A(n2386), .B(n2385), .S(n8293), .Z(n2387) );
  MUX2_X1 U21339 ( .A(\mem[674][2] ), .B(\mem[675][2] ), .S(n8381), .Z(n2388)
         );
  MUX2_X1 U21340 ( .A(\mem[672][2] ), .B(\mem[673][2] ), .S(n8380), .Z(n2389)
         );
  MUX2_X1 U21341 ( .A(n2389), .B(n2388), .S(n8294), .Z(n2390) );
  MUX2_X1 U21342 ( .A(n2390), .B(n2387), .S(n8251), .Z(n2391) );
  MUX2_X1 U21343 ( .A(n2391), .B(n2384), .S(n8204), .Z(n2392) );
  MUX2_X1 U21344 ( .A(n2392), .B(n2377), .S(n8187), .Z(n2393) );
  MUX2_X1 U21345 ( .A(\mem[670][2] ), .B(\mem[671][2] ), .S(n8379), .Z(n2394)
         );
  MUX2_X1 U21346 ( .A(\mem[668][2] ), .B(\mem[669][2] ), .S(n8378), .Z(n2395)
         );
  MUX2_X1 U21347 ( .A(n2395), .B(n2394), .S(n8295), .Z(n2396) );
  MUX2_X1 U21348 ( .A(\mem[666][2] ), .B(\mem[667][2] ), .S(n8372), .Z(n2397)
         );
  MUX2_X1 U21349 ( .A(\mem[664][2] ), .B(\mem[665][2] ), .S(n8538), .Z(n2398)
         );
  MUX2_X1 U21350 ( .A(n2398), .B(n2397), .S(n8302), .Z(n2399) );
  MUX2_X1 U21351 ( .A(n2399), .B(n2396), .S(n8251), .Z(n2400) );
  MUX2_X1 U21352 ( .A(\mem[662][2] ), .B(\mem[663][2] ), .S(n8516), .Z(n2401)
         );
  MUX2_X1 U21353 ( .A(\mem[660][2] ), .B(\mem[661][2] ), .S(n8499), .Z(n2402)
         );
  MUX2_X1 U21354 ( .A(n2402), .B(n2401), .S(n8303), .Z(n2403) );
  MUX2_X1 U21355 ( .A(\mem[658][2] ), .B(\mem[659][2] ), .S(n8482), .Z(n2404)
         );
  MUX2_X1 U21356 ( .A(\mem[656][2] ), .B(\mem[657][2] ), .S(n8445), .Z(n2405)
         );
  MUX2_X1 U21357 ( .A(n2405), .B(n2404), .S(n8304), .Z(n2406) );
  MUX2_X1 U21358 ( .A(n2406), .B(n2403), .S(n8251), .Z(n2407) );
  MUX2_X1 U21359 ( .A(n2407), .B(n2400), .S(n8205), .Z(n2408) );
  MUX2_X1 U21360 ( .A(\mem[654][2] ), .B(\mem[655][2] ), .S(n8530), .Z(n2409)
         );
  MUX2_X1 U21361 ( .A(\mem[652][2] ), .B(\mem[653][2] ), .S(n8389), .Z(n2410)
         );
  MUX2_X1 U21362 ( .A(n2410), .B(n2409), .S(n8299), .Z(n2411) );
  MUX2_X1 U21363 ( .A(\mem[650][2] ), .B(\mem[651][2] ), .S(n8412), .Z(n2412)
         );
  MUX2_X1 U21364 ( .A(\mem[648][2] ), .B(\mem[649][2] ), .S(n8423), .Z(n2413)
         );
  MUX2_X1 U21365 ( .A(n2413), .B(n2412), .S(n8300), .Z(n2414) );
  MUX2_X1 U21366 ( .A(n2414), .B(n2411), .S(n8251), .Z(n2415) );
  MUX2_X1 U21367 ( .A(\mem[646][2] ), .B(\mem[647][2] ), .S(n8387), .Z(n2416)
         );
  MUX2_X1 U21368 ( .A(\mem[644][2] ), .B(\mem[645][2] ), .S(n8436), .Z(n2417)
         );
  MUX2_X1 U21369 ( .A(n2417), .B(n2416), .S(n8301), .Z(n2418) );
  MUX2_X1 U21370 ( .A(\mem[642][2] ), .B(\mem[643][2] ), .S(n8498), .Z(n2419)
         );
  MUX2_X1 U21371 ( .A(\mem[640][2] ), .B(\mem[641][2] ), .S(n8524), .Z(n2420)
         );
  MUX2_X1 U21372 ( .A(n2420), .B(n2419), .S(N19), .Z(n2421) );
  MUX2_X1 U21373 ( .A(n2421), .B(n2418), .S(n8251), .Z(n2422) );
  MUX2_X1 U21374 ( .A(n2422), .B(n2415), .S(n8206), .Z(n2423) );
  MUX2_X1 U21375 ( .A(n2423), .B(n2408), .S(n8188), .Z(n2424) );
  MUX2_X1 U21376 ( .A(n2424), .B(n2393), .S(n8183), .Z(n2425) );
  MUX2_X1 U21377 ( .A(n2425), .B(n2362), .S(N24), .Z(n2426) );
  MUX2_X1 U21378 ( .A(\mem[638][2] ), .B(\mem[639][2] ), .S(n8527), .Z(n2427)
         );
  MUX2_X1 U21379 ( .A(\mem[636][2] ), .B(\mem[637][2] ), .S(n8513), .Z(n2428)
         );
  MUX2_X1 U21380 ( .A(n2428), .B(n2427), .S(n8268), .Z(n2429) );
  MUX2_X1 U21381 ( .A(\mem[634][2] ), .B(\mem[635][2] ), .S(n8504), .Z(n2430)
         );
  MUX2_X1 U21382 ( .A(\mem[632][2] ), .B(\mem[633][2] ), .S(n8484), .Z(n2431)
         );
  MUX2_X1 U21383 ( .A(n2431), .B(n2430), .S(n8288), .Z(n2432) );
  MUX2_X1 U21384 ( .A(n2432), .B(n2429), .S(n8252), .Z(n2433) );
  MUX2_X1 U21385 ( .A(\mem[630][2] ), .B(\mem[631][2] ), .S(n8422), .Z(n2434)
         );
  MUX2_X1 U21386 ( .A(\mem[628][2] ), .B(\mem[629][2] ), .S(n8485), .Z(n2435)
         );
  MUX2_X1 U21387 ( .A(n2435), .B(n2434), .S(n8328), .Z(n2436) );
  MUX2_X1 U21388 ( .A(\mem[626][2] ), .B(\mem[627][2] ), .S(n8527), .Z(n2437)
         );
  MUX2_X1 U21389 ( .A(\mem[624][2] ), .B(\mem[625][2] ), .S(n8465), .Z(n2438)
         );
  MUX2_X1 U21390 ( .A(n2438), .B(n2437), .S(n8302), .Z(n2439) );
  MUX2_X1 U21391 ( .A(n2439), .B(n2436), .S(n8252), .Z(n2440) );
  MUX2_X1 U21392 ( .A(n2440), .B(n2433), .S(n8206), .Z(n2441) );
  MUX2_X1 U21393 ( .A(\mem[622][2] ), .B(\mem[623][2] ), .S(n8376), .Z(n2442)
         );
  MUX2_X1 U21394 ( .A(\mem[620][2] ), .B(\mem[621][2] ), .S(n8475), .Z(n2443)
         );
  MUX2_X1 U21395 ( .A(n2443), .B(n2442), .S(n8348), .Z(n2444) );
  MUX2_X1 U21396 ( .A(\mem[618][2] ), .B(\mem[619][2] ), .S(n8454), .Z(n2445)
         );
  MUX2_X1 U21397 ( .A(\mem[616][2] ), .B(\mem[617][2] ), .S(n8418), .Z(n2446)
         );
  MUX2_X1 U21398 ( .A(n2446), .B(n2445), .S(n8280), .Z(n2447) );
  MUX2_X1 U21399 ( .A(n2447), .B(n2444), .S(n8252), .Z(n2448) );
  MUX2_X1 U21400 ( .A(\mem[614][2] ), .B(\mem[615][2] ), .S(n8446), .Z(n2449)
         );
  MUX2_X1 U21401 ( .A(\mem[612][2] ), .B(\mem[613][2] ), .S(n8441), .Z(n2450)
         );
  MUX2_X1 U21402 ( .A(n2450), .B(n2449), .S(n8348), .Z(n2451) );
  MUX2_X1 U21403 ( .A(\mem[610][2] ), .B(\mem[611][2] ), .S(n8442), .Z(n2452)
         );
  MUX2_X1 U21404 ( .A(\mem[608][2] ), .B(\mem[609][2] ), .S(n8443), .Z(n2453)
         );
  MUX2_X1 U21405 ( .A(n2453), .B(n2452), .S(n8333), .Z(n2454) );
  MUX2_X1 U21406 ( .A(n2454), .B(n2451), .S(n8252), .Z(n2455) );
  MUX2_X1 U21407 ( .A(n2455), .B(n2448), .S(N21), .Z(n2456) );
  MUX2_X1 U21408 ( .A(n2456), .B(n2441), .S(N22), .Z(n2457) );
  MUX2_X1 U21409 ( .A(\mem[606][2] ), .B(\mem[607][2] ), .S(n8450), .Z(n2458)
         );
  MUX2_X1 U21410 ( .A(\mem[604][2] ), .B(\mem[605][2] ), .S(n8451), .Z(n2459)
         );
  MUX2_X1 U21411 ( .A(n2459), .B(n2458), .S(n8283), .Z(n2460) );
  MUX2_X1 U21412 ( .A(\mem[602][2] ), .B(\mem[603][2] ), .S(n8452), .Z(n2461)
         );
  MUX2_X1 U21413 ( .A(\mem[600][2] ), .B(\mem[601][2] ), .S(n8447), .Z(n2462)
         );
  MUX2_X1 U21414 ( .A(n2462), .B(n2461), .S(n8313), .Z(n2463) );
  MUX2_X1 U21415 ( .A(n2463), .B(n2460), .S(n8252), .Z(n2464) );
  MUX2_X1 U21416 ( .A(\mem[598][2] ), .B(\mem[599][2] ), .S(n8448), .Z(n2465)
         );
  MUX2_X1 U21417 ( .A(\mem[596][2] ), .B(\mem[597][2] ), .S(n8449), .Z(n2466)
         );
  MUX2_X1 U21418 ( .A(n2466), .B(n2465), .S(n8349), .Z(n2467) );
  MUX2_X1 U21419 ( .A(\mem[594][2] ), .B(\mem[595][2] ), .S(n8456), .Z(n2468)
         );
  MUX2_X1 U21420 ( .A(\mem[592][2] ), .B(\mem[593][2] ), .S(n8457), .Z(n2469)
         );
  MUX2_X1 U21421 ( .A(n2469), .B(n2468), .S(n8334), .Z(n2470) );
  MUX2_X1 U21422 ( .A(n2470), .B(n2467), .S(n8252), .Z(n2471) );
  MUX2_X1 U21423 ( .A(n2471), .B(n2464), .S(n8198), .Z(n2472) );
  MUX2_X1 U21424 ( .A(\mem[590][2] ), .B(\mem[591][2] ), .S(n8512), .Z(n2473)
         );
  MUX2_X1 U21425 ( .A(\mem[588][2] ), .B(\mem[589][2] ), .S(n8507), .Z(n2474)
         );
  MUX2_X1 U21426 ( .A(n2474), .B(n2473), .S(n8270), .Z(n2475) );
  MUX2_X1 U21427 ( .A(\mem[586][2] ), .B(\mem[587][2] ), .S(n8508), .Z(n2476)
         );
  MUX2_X1 U21428 ( .A(\mem[584][2] ), .B(\mem[585][2] ), .S(n8509), .Z(n2477)
         );
  MUX2_X1 U21429 ( .A(n2477), .B(n2476), .S(n8289), .Z(n2478) );
  MUX2_X1 U21430 ( .A(n2478), .B(n2475), .S(n8252), .Z(n2479) );
  MUX2_X1 U21431 ( .A(\mem[582][2] ), .B(\mem[583][2] ), .S(n8516), .Z(n2480)
         );
  MUX2_X1 U21432 ( .A(\mem[580][2] ), .B(\mem[581][2] ), .S(n8517), .Z(n2481)
         );
  MUX2_X1 U21433 ( .A(n2481), .B(n2480), .S(n8289), .Z(n2482) );
  MUX2_X1 U21434 ( .A(\mem[578][2] ), .B(\mem[579][2] ), .S(n8518), .Z(n2483)
         );
  MUX2_X1 U21435 ( .A(\mem[576][2] ), .B(\mem[577][2] ), .S(n8513), .Z(n2484)
         );
  MUX2_X1 U21436 ( .A(n2484), .B(n2483), .S(n8290), .Z(n2485) );
  MUX2_X1 U21437 ( .A(n2485), .B(n2482), .S(n8252), .Z(n2486) );
  MUX2_X1 U21438 ( .A(n2486), .B(n2479), .S(n8201), .Z(n2487) );
  MUX2_X1 U21439 ( .A(n2487), .B(n2472), .S(N22), .Z(n2488) );
  MUX2_X1 U21440 ( .A(n2488), .B(n2457), .S(n8183), .Z(n2489) );
  MUX2_X1 U21441 ( .A(\mem[574][2] ), .B(\mem[575][2] ), .S(n8514), .Z(n2490)
         );
  MUX2_X1 U21442 ( .A(\mem[572][2] ), .B(\mem[573][2] ), .S(n8515), .Z(n2491)
         );
  MUX2_X1 U21443 ( .A(n2491), .B(n2490), .S(n8348), .Z(n2492) );
  MUX2_X1 U21444 ( .A(\mem[570][2] ), .B(\mem[571][2] ), .S(n8522), .Z(n2493)
         );
  MUX2_X1 U21445 ( .A(\mem[568][2] ), .B(\mem[569][2] ), .S(n8523), .Z(n2494)
         );
  MUX2_X1 U21446 ( .A(n2494), .B(n2493), .S(n8340), .Z(n2495) );
  MUX2_X1 U21447 ( .A(n2495), .B(n2492), .S(n8252), .Z(n2496) );
  MUX2_X1 U21448 ( .A(\mem[566][2] ), .B(\mem[567][2] ), .S(n8461), .Z(n2497)
         );
  MUX2_X1 U21449 ( .A(\mem[564][2] ), .B(\mem[565][2] ), .S(n8468), .Z(n2498)
         );
  MUX2_X1 U21450 ( .A(n2498), .B(n2497), .S(n8319), .Z(n2499) );
  MUX2_X1 U21451 ( .A(\mem[562][2] ), .B(\mem[563][2] ), .S(n8469), .Z(n2500)
         );
  MUX2_X1 U21452 ( .A(\mem[560][2] ), .B(\mem[561][2] ), .S(n8530), .Z(n2501)
         );
  MUX2_X1 U21453 ( .A(n2501), .B(n2500), .S(n8305), .Z(n2502) );
  MUX2_X1 U21454 ( .A(n2502), .B(n2499), .S(n8252), .Z(n2503) );
  MUX2_X1 U21455 ( .A(n2503), .B(n2496), .S(n8199), .Z(n2504) );
  MUX2_X1 U21456 ( .A(\mem[558][2] ), .B(\mem[559][2] ), .S(n8459), .Z(n2505)
         );
  MUX2_X1 U21457 ( .A(\mem[556][2] ), .B(\mem[557][2] ), .S(n8374), .Z(n2506)
         );
  MUX2_X1 U21458 ( .A(n2506), .B(n2505), .S(n8315), .Z(n2507) );
  MUX2_X1 U21459 ( .A(\mem[554][2] ), .B(\mem[555][2] ), .S(n8494), .Z(n2508)
         );
  MUX2_X1 U21460 ( .A(\mem[552][2] ), .B(\mem[553][2] ), .S(N18), .Z(n2509) );
  MUX2_X1 U21461 ( .A(n2509), .B(n2508), .S(n8269), .Z(n2510) );
  MUX2_X1 U21462 ( .A(n2510), .B(n2507), .S(n8252), .Z(n2511) );
  MUX2_X1 U21463 ( .A(\mem[550][2] ), .B(\mem[551][2] ), .S(n8377), .Z(n2512)
         );
  MUX2_X1 U21464 ( .A(\mem[548][2] ), .B(\mem[549][2] ), .S(n8418), .Z(n2513)
         );
  MUX2_X1 U21465 ( .A(n2513), .B(n2512), .S(n8305), .Z(n2514) );
  MUX2_X1 U21466 ( .A(\mem[546][2] ), .B(\mem[547][2] ), .S(n8534), .Z(n2515)
         );
  MUX2_X1 U21467 ( .A(\mem[544][2] ), .B(\mem[545][2] ), .S(n8528), .Z(n2516)
         );
  MUX2_X1 U21468 ( .A(n2516), .B(n2515), .S(n8303), .Z(n2517) );
  MUX2_X1 U21469 ( .A(n2517), .B(n2514), .S(n8252), .Z(n2518) );
  MUX2_X1 U21470 ( .A(n2518), .B(n2511), .S(n8200), .Z(n2519) );
  MUX2_X1 U21471 ( .A(n2519), .B(n2504), .S(N22), .Z(n2520) );
  MUX2_X1 U21472 ( .A(\mem[542][2] ), .B(\mem[543][2] ), .S(n8491), .Z(n2521)
         );
  MUX2_X1 U21473 ( .A(\mem[540][2] ), .B(\mem[541][2] ), .S(n8498), .Z(n2522)
         );
  MUX2_X1 U21474 ( .A(n2522), .B(n2521), .S(n8279), .Z(n2523) );
  MUX2_X1 U21475 ( .A(\mem[538][2] ), .B(\mem[539][2] ), .S(n8499), .Z(n2524)
         );
  MUX2_X1 U21476 ( .A(\mem[536][2] ), .B(\mem[537][2] ), .S(n8500), .Z(n2525)
         );
  MUX2_X1 U21477 ( .A(n2525), .B(n2524), .S(n8323), .Z(n2526) );
  MUX2_X1 U21478 ( .A(n2526), .B(n2523), .S(n8253), .Z(n2527) );
  MUX2_X1 U21479 ( .A(\mem[534][2] ), .B(\mem[535][2] ), .S(n8495), .Z(n2528)
         );
  MUX2_X1 U21480 ( .A(\mem[532][2] ), .B(\mem[533][2] ), .S(n8496), .Z(n2529)
         );
  MUX2_X1 U21481 ( .A(n2529), .B(n2528), .S(n8278), .Z(n2530) );
  MUX2_X1 U21482 ( .A(\mem[530][2] ), .B(\mem[531][2] ), .S(n8497), .Z(n2531)
         );
  MUX2_X1 U21483 ( .A(\mem[528][2] ), .B(\mem[529][2] ), .S(n8504), .Z(n2532)
         );
  MUX2_X1 U21484 ( .A(n2532), .B(n2531), .S(n8277), .Z(n2533) );
  MUX2_X1 U21485 ( .A(n2533), .B(n2530), .S(n8253), .Z(n2534) );
  MUX2_X1 U21486 ( .A(n2534), .B(n2527), .S(n8198), .Z(n2535) );
  MUX2_X1 U21487 ( .A(\mem[526][2] ), .B(\mem[527][2] ), .S(n8505), .Z(n2536)
         );
  MUX2_X1 U21488 ( .A(\mem[524][2] ), .B(\mem[525][2] ), .S(n8506), .Z(n2537)
         );
  MUX2_X1 U21489 ( .A(n2537), .B(n2536), .S(n8276), .Z(n2538) );
  MUX2_X1 U21490 ( .A(\mem[522][2] ), .B(\mem[523][2] ), .S(n8501), .Z(n2539)
         );
  MUX2_X1 U21491 ( .A(\mem[520][2] ), .B(\mem[521][2] ), .S(n8502), .Z(n2540)
         );
  MUX2_X1 U21492 ( .A(n2540), .B(n2539), .S(n8272), .Z(n2541) );
  MUX2_X1 U21493 ( .A(n2541), .B(n2538), .S(n8253), .Z(n2542) );
  MUX2_X1 U21494 ( .A(\mem[518][2] ), .B(\mem[519][2] ), .S(n8515), .Z(n2543)
         );
  MUX2_X1 U21495 ( .A(\mem[516][2] ), .B(\mem[517][2] ), .S(n8497), .Z(n2544)
         );
  MUX2_X1 U21496 ( .A(n2544), .B(n2543), .S(n8271), .Z(n2545) );
  MUX2_X1 U21497 ( .A(\mem[514][2] ), .B(\mem[515][2] ), .S(n8424), .Z(n2546)
         );
  MUX2_X1 U21498 ( .A(\mem[512][2] ), .B(\mem[513][2] ), .S(n8408), .Z(n2547)
         );
  MUX2_X1 U21499 ( .A(n2547), .B(n2546), .S(n8275), .Z(n2548) );
  MUX2_X1 U21500 ( .A(n2548), .B(n2545), .S(n8253), .Z(n2549) );
  MUX2_X1 U21501 ( .A(n2549), .B(n2542), .S(n8208), .Z(n2550) );
  MUX2_X1 U21502 ( .A(n2550), .B(n2535), .S(n8196), .Z(n2551) );
  MUX2_X1 U21503 ( .A(n2551), .B(n2520), .S(n8183), .Z(n2552) );
  MUX2_X1 U21504 ( .A(n2552), .B(n2489), .S(n8179), .Z(n2553) );
  MUX2_X1 U21505 ( .A(n2553), .B(n2426), .S(n8177), .Z(n2554) );
  MUX2_X1 U21506 ( .A(n2554), .B(n2299), .S(N26), .Z(n2555) );
  MUX2_X1 U21507 ( .A(\mem[510][2] ), .B(\mem[511][2] ), .S(n8426), .Z(n2556)
         );
  MUX2_X1 U21508 ( .A(\mem[508][2] ), .B(\mem[509][2] ), .S(n8465), .Z(n2557)
         );
  MUX2_X1 U21509 ( .A(n2557), .B(n2556), .S(n8273), .Z(n2558) );
  MUX2_X1 U21510 ( .A(\mem[506][2] ), .B(\mem[507][2] ), .S(n8464), .Z(n2559)
         );
  MUX2_X1 U21511 ( .A(\mem[504][2] ), .B(\mem[505][2] ), .S(n8503), .Z(n2560)
         );
  MUX2_X1 U21512 ( .A(n2560), .B(n2559), .S(n8268), .Z(n2561) );
  MUX2_X1 U21513 ( .A(n2561), .B(n2558), .S(n8253), .Z(n2562) );
  MUX2_X1 U21514 ( .A(\mem[502][2] ), .B(\mem[503][2] ), .S(n8497), .Z(n2563)
         );
  MUX2_X1 U21515 ( .A(\mem[500][2] ), .B(\mem[501][2] ), .S(n8510), .Z(n2564)
         );
  MUX2_X1 U21516 ( .A(n2564), .B(n2563), .S(n8347), .Z(n2565) );
  MUX2_X1 U21517 ( .A(\mem[498][2] ), .B(\mem[499][2] ), .S(n8489), .Z(n2566)
         );
  MUX2_X1 U21518 ( .A(\mem[496][2] ), .B(\mem[497][2] ), .S(n8490), .Z(n2567)
         );
  MUX2_X1 U21519 ( .A(n2567), .B(n2566), .S(n8269), .Z(n2568) );
  MUX2_X1 U21520 ( .A(n2568), .B(n2565), .S(n8253), .Z(n2569) );
  MUX2_X1 U21521 ( .A(n2569), .B(n2562), .S(n8208), .Z(n2570) );
  MUX2_X1 U21522 ( .A(\mem[494][2] ), .B(\mem[495][2] ), .S(n8363), .Z(n2571)
         );
  MUX2_X1 U21523 ( .A(\mem[492][2] ), .B(\mem[493][2] ), .S(n8407), .Z(n2572)
         );
  MUX2_X1 U21524 ( .A(n2572), .B(n2571), .S(n8327), .Z(n2573) );
  MUX2_X1 U21525 ( .A(\mem[490][2] ), .B(\mem[491][2] ), .S(n8458), .Z(n2574)
         );
  MUX2_X1 U21526 ( .A(\mem[488][2] ), .B(\mem[489][2] ), .S(n8434), .Z(n2575)
         );
  MUX2_X1 U21527 ( .A(n2575), .B(n2574), .S(n8328), .Z(n2576) );
  MUX2_X1 U21528 ( .A(n2576), .B(n2573), .S(n8253), .Z(n2577) );
  MUX2_X1 U21529 ( .A(\mem[486][2] ), .B(\mem[487][2] ), .S(n8429), .Z(n2578)
         );
  MUX2_X1 U21530 ( .A(\mem[484][2] ), .B(\mem[485][2] ), .S(n8412), .Z(n2579)
         );
  MUX2_X1 U21531 ( .A(n2579), .B(n2578), .S(n8323), .Z(n2580) );
  MUX2_X1 U21532 ( .A(\mem[482][2] ), .B(\mem[483][2] ), .S(n8406), .Z(n2581)
         );
  MUX2_X1 U21533 ( .A(\mem[480][2] ), .B(\mem[481][2] ), .S(n8357), .Z(n2582)
         );
  MUX2_X1 U21534 ( .A(n2582), .B(n2581), .S(n8324), .Z(n2583) );
  MUX2_X1 U21535 ( .A(n2583), .B(n2580), .S(n8253), .Z(n2584) );
  MUX2_X1 U21536 ( .A(n2584), .B(n2577), .S(N21), .Z(n2585) );
  MUX2_X1 U21537 ( .A(n2585), .B(n2570), .S(n8194), .Z(n2586) );
  MUX2_X1 U21538 ( .A(\mem[478][2] ), .B(\mem[479][2] ), .S(n8537), .Z(n2587)
         );
  MUX2_X1 U21539 ( .A(\mem[476][2] ), .B(\mem[477][2] ), .S(n8401), .Z(n2588)
         );
  MUX2_X1 U21540 ( .A(n2588), .B(n2587), .S(n8325), .Z(n2589) );
  MUX2_X1 U21541 ( .A(\mem[474][2] ), .B(\mem[475][2] ), .S(n8357), .Z(n2590)
         );
  MUX2_X1 U21542 ( .A(\mem[472][2] ), .B(\mem[473][2] ), .S(n8406), .Z(n2591)
         );
  MUX2_X1 U21543 ( .A(n2591), .B(n2590), .S(n8333), .Z(n2592) );
  MUX2_X1 U21544 ( .A(n2592), .B(n2589), .S(n8253), .Z(n2593) );
  MUX2_X1 U21545 ( .A(\mem[470][2] ), .B(\mem[471][2] ), .S(n8413), .Z(n2594)
         );
  MUX2_X1 U21546 ( .A(\mem[468][2] ), .B(\mem[469][2] ), .S(n8451), .Z(n2595)
         );
  MUX2_X1 U21547 ( .A(n2595), .B(n2594), .S(n8334), .Z(n2596) );
  MUX2_X1 U21548 ( .A(\mem[466][2] ), .B(\mem[467][2] ), .S(n8440), .Z(n2597)
         );
  MUX2_X1 U21549 ( .A(\mem[464][2] ), .B(\mem[465][2] ), .S(n8407), .Z(n2598)
         );
  MUX2_X1 U21550 ( .A(n2598), .B(n2597), .S(n8329), .Z(n2599) );
  MUX2_X1 U21551 ( .A(n2599), .B(n2596), .S(n8253), .Z(n2600) );
  MUX2_X1 U21552 ( .A(n2600), .B(n2593), .S(n8199), .Z(n2601) );
  MUX2_X1 U21553 ( .A(\mem[462][2] ), .B(\mem[463][2] ), .S(n8478), .Z(n2602)
         );
  MUX2_X1 U21554 ( .A(\mem[460][2] ), .B(\mem[461][2] ), .S(n8359), .Z(n2603)
         );
  MUX2_X1 U21555 ( .A(n2603), .B(n2602), .S(n8330), .Z(n2604) );
  MUX2_X1 U21556 ( .A(\mem[458][2] ), .B(\mem[459][2] ), .S(n8360), .Z(n2605)
         );
  MUX2_X1 U21557 ( .A(\mem[456][2] ), .B(\mem[457][2] ), .S(n8539), .Z(n2606)
         );
  MUX2_X1 U21558 ( .A(n2606), .B(n2605), .S(n8331), .Z(n2607) );
  MUX2_X1 U21559 ( .A(n2607), .B(n2604), .S(n8253), .Z(n2608) );
  MUX2_X1 U21560 ( .A(\mem[454][2] ), .B(\mem[455][2] ), .S(n8362), .Z(n2609)
         );
  MUX2_X1 U21561 ( .A(\mem[452][2] ), .B(\mem[453][2] ), .S(n8358), .Z(n2610)
         );
  MUX2_X1 U21562 ( .A(n2610), .B(n2609), .S(n8338), .Z(n2611) );
  MUX2_X1 U21563 ( .A(\mem[450][2] ), .B(\mem[451][2] ), .S(n8432), .Z(n2612)
         );
  MUX2_X1 U21564 ( .A(\mem[448][2] ), .B(\mem[449][2] ), .S(n8364), .Z(n2613)
         );
  MUX2_X1 U21565 ( .A(n2613), .B(n2612), .S(n8339), .Z(n2614) );
  MUX2_X1 U21566 ( .A(n2614), .B(n2611), .S(n8253), .Z(n2615) );
  MUX2_X1 U21567 ( .A(n2615), .B(n2608), .S(n8219), .Z(n2616) );
  MUX2_X1 U21568 ( .A(n2616), .B(n2601), .S(n8192), .Z(n2617) );
  MUX2_X1 U21569 ( .A(n2617), .B(n2586), .S(n8183), .Z(n2618) );
  MUX2_X1 U21570 ( .A(\mem[446][2] ), .B(\mem[447][2] ), .S(n8520), .Z(n2619)
         );
  MUX2_X1 U21571 ( .A(\mem[444][2] ), .B(\mem[445][2] ), .S(n8521), .Z(n2620)
         );
  MUX2_X1 U21572 ( .A(n2620), .B(n2619), .S(n8307), .Z(n2621) );
  MUX2_X1 U21573 ( .A(\mem[442][2] ), .B(\mem[443][2] ), .S(n8528), .Z(n2622)
         );
  MUX2_X1 U21574 ( .A(\mem[440][2] ), .B(\mem[441][2] ), .S(n8529), .Z(n2623)
         );
  MUX2_X1 U21575 ( .A(n2623), .B(n2622), .S(n8314), .Z(n2624) );
  MUX2_X1 U21576 ( .A(n2624), .B(n2621), .S(n8254), .Z(n2625) );
  MUX2_X1 U21577 ( .A(\mem[438][2] ), .B(\mem[439][2] ), .S(n8530), .Z(n2626)
         );
  MUX2_X1 U21578 ( .A(\mem[436][2] ), .B(\mem[437][2] ), .S(n8525), .Z(n2627)
         );
  MUX2_X1 U21579 ( .A(n2627), .B(n2626), .S(n8315), .Z(n2628) );
  MUX2_X1 U21580 ( .A(\mem[434][2] ), .B(\mem[435][2] ), .S(n8375), .Z(n2629)
         );
  MUX2_X1 U21581 ( .A(\mem[432][2] ), .B(\mem[433][2] ), .S(n8374), .Z(n2630)
         );
  MUX2_X1 U21582 ( .A(n2630), .B(n2629), .S(n8316), .Z(n2631) );
  MUX2_X1 U21583 ( .A(n2631), .B(n2628), .S(n8254), .Z(n2632) );
  MUX2_X1 U21584 ( .A(n2632), .B(n2625), .S(n8219), .Z(n2633) );
  MUX2_X1 U21585 ( .A(\mem[430][2] ), .B(\mem[431][2] ), .S(n8369), .Z(n2634)
         );
  MUX2_X1 U21586 ( .A(\mem[428][2] ), .B(\mem[429][2] ), .S(n8368), .Z(n2635)
         );
  MUX2_X1 U21587 ( .A(n2635), .B(n2634), .S(n8311), .Z(n2636) );
  MUX2_X1 U21588 ( .A(\mem[426][2] ), .B(\mem[427][2] ), .S(n8385), .Z(n2637)
         );
  MUX2_X1 U21589 ( .A(\mem[424][2] ), .B(\mem[425][2] ), .S(n8367), .Z(n2638)
         );
  MUX2_X1 U21590 ( .A(n2638), .B(n2637), .S(n8312), .Z(n2639) );
  MUX2_X1 U21591 ( .A(n2639), .B(n2636), .S(n8254), .Z(n2640) );
  MUX2_X1 U21592 ( .A(\mem[422][2] ), .B(\mem[423][2] ), .S(n8527), .Z(n2641)
         );
  MUX2_X1 U21593 ( .A(\mem[420][2] ), .B(\mem[421][2] ), .S(n8509), .Z(n2642)
         );
  MUX2_X1 U21594 ( .A(n2642), .B(n2641), .S(n8313), .Z(n2643) );
  MUX2_X1 U21595 ( .A(\mem[418][2] ), .B(\mem[419][2] ), .S(n8498), .Z(n2644)
         );
  MUX2_X1 U21596 ( .A(\mem[416][2] ), .B(\mem[417][2] ), .S(n8481), .Z(n2645)
         );
  MUX2_X1 U21597 ( .A(n2645), .B(n2644), .S(n8320), .Z(n2646) );
  MUX2_X1 U21598 ( .A(n2646), .B(n2643), .S(n8254), .Z(n2647) );
  MUX2_X1 U21599 ( .A(n2647), .B(n2640), .S(n8212), .Z(n2648) );
  MUX2_X1 U21600 ( .A(n2648), .B(n2633), .S(n8195), .Z(n2649) );
  MUX2_X1 U21601 ( .A(\mem[414][2] ), .B(\mem[415][2] ), .S(n8444), .Z(n2650)
         );
  MUX2_X1 U21602 ( .A(\mem[412][2] ), .B(\mem[413][2] ), .S(n8406), .Z(n2651)
         );
  MUX2_X1 U21603 ( .A(n2651), .B(n2650), .S(n8321), .Z(n2652) );
  MUX2_X1 U21604 ( .A(\mem[410][2] ), .B(\mem[411][2] ), .S(n8392), .Z(n2653)
         );
  MUX2_X1 U21605 ( .A(\mem[408][2] ), .B(\mem[409][2] ), .S(n8419), .Z(n2654)
         );
  MUX2_X1 U21606 ( .A(n2654), .B(n2653), .S(n8322), .Z(n2655) );
  MUX2_X1 U21607 ( .A(n2655), .B(n2652), .S(n8254), .Z(n2656) );
  MUX2_X1 U21608 ( .A(\mem[406][2] ), .B(\mem[407][2] ), .S(n8464), .Z(n2657)
         );
  MUX2_X1 U21609 ( .A(\mem[404][2] ), .B(\mem[405][2] ), .S(n8439), .Z(n2658)
         );
  MUX2_X1 U21610 ( .A(n2658), .B(n2657), .S(n8317), .Z(n2659) );
  MUX2_X1 U21611 ( .A(\mem[402][2] ), .B(\mem[403][2] ), .S(n8518), .Z(n2660)
         );
  MUX2_X1 U21612 ( .A(\mem[400][2] ), .B(\mem[401][2] ), .S(n8378), .Z(n2661)
         );
  MUX2_X1 U21613 ( .A(n2661), .B(n2660), .S(n8318), .Z(n2662) );
  MUX2_X1 U21614 ( .A(n2662), .B(n2659), .S(n8254), .Z(n2663) );
  MUX2_X1 U21615 ( .A(n2663), .B(n2656), .S(n8201), .Z(n2664) );
  MUX2_X1 U21616 ( .A(\mem[398][2] ), .B(\mem[399][2] ), .S(n8443), .Z(n2665)
         );
  MUX2_X1 U21617 ( .A(\mem[396][2] ), .B(\mem[397][2] ), .S(n8433), .Z(n2666)
         );
  MUX2_X1 U21618 ( .A(n2666), .B(n2665), .S(n8286), .Z(n2667) );
  MUX2_X1 U21619 ( .A(\mem[394][2] ), .B(\mem[395][2] ), .S(n8538), .Z(n2668)
         );
  MUX2_X1 U21620 ( .A(\mem[392][2] ), .B(\mem[393][2] ), .S(n8470), .Z(n2669)
         );
  MUX2_X1 U21621 ( .A(n2669), .B(n2668), .S(n8307), .Z(n2670) );
  MUX2_X1 U21622 ( .A(n2670), .B(n2667), .S(n8254), .Z(n2671) );
  MUX2_X1 U21623 ( .A(\mem[390][2] ), .B(\mem[391][2] ), .S(n8374), .Z(n2672)
         );
  MUX2_X1 U21624 ( .A(\mem[388][2] ), .B(\mem[389][2] ), .S(n8470), .Z(n2673)
         );
  MUX2_X1 U21625 ( .A(n2673), .B(n2672), .S(n8355), .Z(n2674) );
  MUX2_X1 U21626 ( .A(\mem[386][2] ), .B(\mem[387][2] ), .S(n8368), .Z(n2675)
         );
  MUX2_X1 U21627 ( .A(\mem[384][2] ), .B(\mem[385][2] ), .S(n8388), .Z(n2676)
         );
  MUX2_X1 U21628 ( .A(n2676), .B(n2675), .S(n8325), .Z(n2677) );
  MUX2_X1 U21629 ( .A(n2677), .B(n2674), .S(n8254), .Z(n2678) );
  MUX2_X1 U21630 ( .A(n2678), .B(n2671), .S(n8199), .Z(n2679) );
  MUX2_X1 U21631 ( .A(n2679), .B(n2664), .S(n8189), .Z(n2680) );
  MUX2_X1 U21632 ( .A(n2680), .B(n2649), .S(n8183), .Z(n2681) );
  MUX2_X1 U21633 ( .A(n2681), .B(n2618), .S(n8180), .Z(n2682) );
  MUX2_X1 U21634 ( .A(\mem[382][2] ), .B(\mem[383][2] ), .S(n8401), .Z(n2683)
         );
  MUX2_X1 U21635 ( .A(\mem[380][2] ), .B(\mem[381][2] ), .S(n8417), .Z(n2684)
         );
  MUX2_X1 U21636 ( .A(n2684), .B(n2683), .S(n8341), .Z(n2685) );
  MUX2_X1 U21637 ( .A(\mem[378][2] ), .B(\mem[379][2] ), .S(n8409), .Z(n2686)
         );
  MUX2_X1 U21638 ( .A(\mem[376][2] ), .B(\mem[377][2] ), .S(n8398), .Z(n2687)
         );
  MUX2_X1 U21639 ( .A(n2687), .B(n2686), .S(n8306), .Z(n2688) );
  MUX2_X1 U21640 ( .A(n2688), .B(n2685), .S(n8254), .Z(n2689) );
  MUX2_X1 U21641 ( .A(\mem[374][2] ), .B(\mem[375][2] ), .S(n8388), .Z(n2690)
         );
  MUX2_X1 U21642 ( .A(\mem[372][2] ), .B(\mem[373][2] ), .S(n8447), .Z(n2691)
         );
  MUX2_X1 U21643 ( .A(n2691), .B(n2690), .S(n8288), .Z(n2692) );
  MUX2_X1 U21644 ( .A(\mem[370][2] ), .B(\mem[371][2] ), .S(n8397), .Z(n2693)
         );
  MUX2_X1 U21645 ( .A(\mem[368][2] ), .B(\mem[369][2] ), .S(n8530), .Z(n2694)
         );
  MUX2_X1 U21646 ( .A(n2694), .B(n2693), .S(n8328), .Z(n2695) );
  MUX2_X1 U21647 ( .A(n2695), .B(n2692), .S(n8254), .Z(n2696) );
  MUX2_X1 U21648 ( .A(n2696), .B(n2689), .S(n8217), .Z(n2697) );
  MUX2_X1 U21649 ( .A(\mem[366][2] ), .B(\mem[367][2] ), .S(n8508), .Z(n2698)
         );
  MUX2_X1 U21650 ( .A(\mem[364][2] ), .B(\mem[365][2] ), .S(n8499), .Z(n2699)
         );
  MUX2_X1 U21651 ( .A(n2699), .B(n2698), .S(n8276), .Z(n2700) );
  MUX2_X1 U21652 ( .A(\mem[362][2] ), .B(\mem[363][2] ), .S(n8424), .Z(n2701)
         );
  MUX2_X1 U21653 ( .A(\mem[360][2] ), .B(\mem[361][2] ), .S(n8486), .Z(n2702)
         );
  MUX2_X1 U21654 ( .A(n2702), .B(n2701), .S(n8308), .Z(n2703) );
  MUX2_X1 U21655 ( .A(n2703), .B(n2700), .S(n8254), .Z(n2704) );
  MUX2_X1 U21656 ( .A(\mem[358][2] ), .B(\mem[359][2] ), .S(n8528), .Z(n2705)
         );
  MUX2_X1 U21657 ( .A(\mem[356][2] ), .B(\mem[357][2] ), .S(n8507), .Z(n2706)
         );
  MUX2_X1 U21658 ( .A(n2706), .B(n2705), .S(n8309), .Z(n2707) );
  MUX2_X1 U21659 ( .A(\mem[354][2] ), .B(\mem[355][2] ), .S(n8491), .Z(n2708)
         );
  MUX2_X1 U21660 ( .A(\mem[352][2] ), .B(\mem[353][2] ), .S(n8481), .Z(n2709)
         );
  MUX2_X1 U21661 ( .A(n2709), .B(n2708), .S(n8310), .Z(n2710) );
  MUX2_X1 U21662 ( .A(n2710), .B(n2707), .S(n8254), .Z(n2711) );
  MUX2_X1 U21663 ( .A(n2711), .B(n2704), .S(n8200), .Z(n2712) );
  MUX2_X1 U21664 ( .A(n2712), .B(n2697), .S(n8194), .Z(n2713) );
  MUX2_X1 U21665 ( .A(\mem[350][2] ), .B(\mem[351][2] ), .S(n8506), .Z(n2714)
         );
  MUX2_X1 U21666 ( .A(\mem[348][2] ), .B(\mem[349][2] ), .S(n8501), .Z(n2715)
         );
  MUX2_X1 U21667 ( .A(n2715), .B(n2714), .S(n8343), .Z(n2716) );
  MUX2_X1 U21668 ( .A(\mem[346][2] ), .B(\mem[347][2] ), .S(n8502), .Z(n2717)
         );
  MUX2_X1 U21669 ( .A(\mem[344][2] ), .B(\mem[345][2] ), .S(n8503), .Z(n2718)
         );
  MUX2_X1 U21670 ( .A(n2718), .B(n2717), .S(n8277), .Z(n2719) );
  MUX2_X1 U21671 ( .A(n2719), .B(n2716), .S(n8255), .Z(n2720) );
  MUX2_X1 U21672 ( .A(\mem[342][2] ), .B(\mem[343][2] ), .S(n8510), .Z(n2721)
         );
  MUX2_X1 U21673 ( .A(\mem[340][2] ), .B(\mem[341][2] ), .S(n8511), .Z(n2722)
         );
  MUX2_X1 U21674 ( .A(n2722), .B(n2721), .S(n8308), .Z(n2723) );
  MUX2_X1 U21675 ( .A(\mem[338][2] ), .B(\mem[339][2] ), .S(n8512), .Z(n2724)
         );
  MUX2_X1 U21676 ( .A(\mem[336][2] ), .B(\mem[337][2] ), .S(n8507), .Z(n2725)
         );
  MUX2_X1 U21677 ( .A(n2725), .B(n2724), .S(n8309), .Z(n2726) );
  MUX2_X1 U21678 ( .A(n2726), .B(n2723), .S(n8255), .Z(n2727) );
  MUX2_X1 U21679 ( .A(n2727), .B(n2720), .S(n8213), .Z(n2728) );
  MUX2_X1 U21680 ( .A(\mem[334][2] ), .B(\mem[335][2] ), .S(n8508), .Z(n2729)
         );
  MUX2_X1 U21681 ( .A(\mem[332][2] ), .B(\mem[333][2] ), .S(n8509), .Z(n2730)
         );
  MUX2_X1 U21682 ( .A(n2730), .B(n2729), .S(n8310), .Z(n2731) );
  MUX2_X1 U21683 ( .A(\mem[330][2] ), .B(\mem[331][2] ), .S(n8516), .Z(n2732)
         );
  MUX2_X1 U21684 ( .A(\mem[328][2] ), .B(\mem[329][2] ), .S(n8517), .Z(n2733)
         );
  MUX2_X1 U21685 ( .A(n2733), .B(n2732), .S(n8305), .Z(n2734) );
  MUX2_X1 U21686 ( .A(n2734), .B(n2731), .S(n8255), .Z(n2735) );
  MUX2_X1 U21687 ( .A(\mem[326][2] ), .B(\mem[327][2] ), .S(n8492), .Z(n2736)
         );
  MUX2_X1 U21688 ( .A(\mem[324][2] ), .B(\mem[325][2] ), .S(n8493), .Z(n2737)
         );
  MUX2_X1 U21689 ( .A(n2737), .B(n2736), .S(n8306), .Z(n2738) );
  MUX2_X1 U21690 ( .A(\mem[322][2] ), .B(\mem[323][2] ), .S(n8494), .Z(n2739)
         );
  MUX2_X1 U21691 ( .A(\mem[320][2] ), .B(\mem[321][2] ), .S(n8489), .Z(n2740)
         );
  MUX2_X1 U21692 ( .A(n2740), .B(n2739), .S(n8307), .Z(n2741) );
  MUX2_X1 U21693 ( .A(n2741), .B(n2738), .S(n8255), .Z(n2742) );
  MUX2_X1 U21694 ( .A(n2742), .B(n2735), .S(n8205), .Z(n2743) );
  MUX2_X1 U21695 ( .A(n2743), .B(n2728), .S(N22), .Z(n2744) );
  MUX2_X1 U21696 ( .A(n2744), .B(n2713), .S(n8183), .Z(n2745) );
  MUX2_X1 U21697 ( .A(\mem[318][2] ), .B(\mem[319][2] ), .S(n8490), .Z(n2746)
         );
  MUX2_X1 U21698 ( .A(\mem[316][2] ), .B(\mem[317][2] ), .S(n8491), .Z(n2747)
         );
  MUX2_X1 U21699 ( .A(n2747), .B(n2746), .S(n8314), .Z(n2748) );
  MUX2_X1 U21700 ( .A(\mem[314][2] ), .B(\mem[315][2] ), .S(n8498), .Z(n2749)
         );
  MUX2_X1 U21701 ( .A(\mem[312][2] ), .B(\mem[313][2] ), .S(n8499), .Z(n2750)
         );
  MUX2_X1 U21702 ( .A(n2750), .B(n2749), .S(n8315), .Z(n2751) );
  MUX2_X1 U21703 ( .A(n2751), .B(n2748), .S(n8255), .Z(n2752) );
  MUX2_X1 U21704 ( .A(\mem[310][2] ), .B(\mem[311][2] ), .S(n8500), .Z(n2753)
         );
  MUX2_X1 U21705 ( .A(\mem[308][2] ), .B(\mem[309][2] ), .S(n8495), .Z(n2754)
         );
  MUX2_X1 U21706 ( .A(n2754), .B(n2753), .S(n8316), .Z(n2755) );
  MUX2_X1 U21707 ( .A(\mem[306][2] ), .B(\mem[307][2] ), .S(n8496), .Z(n2756)
         );
  MUX2_X1 U21708 ( .A(\mem[304][2] ), .B(\mem[305][2] ), .S(n8497), .Z(n2757)
         );
  MUX2_X1 U21709 ( .A(n2757), .B(n2756), .S(n8311), .Z(n2758) );
  MUX2_X1 U21710 ( .A(n2758), .B(n2755), .S(n8255), .Z(n2759) );
  MUX2_X1 U21711 ( .A(n2759), .B(n2752), .S(n8213), .Z(n2760) );
  MUX2_X1 U21712 ( .A(\mem[302][2] ), .B(\mem[303][2] ), .S(n8418), .Z(n2761)
         );
  MUX2_X1 U21713 ( .A(\mem[300][2] ), .B(\mem[301][2] ), .S(n8419), .Z(n2762)
         );
  MUX2_X1 U21714 ( .A(n2762), .B(n2761), .S(n8353), .Z(n2763) );
  MUX2_X1 U21715 ( .A(\mem[298][2] ), .B(\mem[299][2] ), .S(n8426), .Z(n2764)
         );
  MUX2_X1 U21716 ( .A(\mem[296][2] ), .B(\mem[297][2] ), .S(n8427), .Z(n2765)
         );
  MUX2_X1 U21717 ( .A(n2765), .B(n2764), .S(n8354), .Z(n2766) );
  MUX2_X1 U21718 ( .A(n2766), .B(n2763), .S(n8255), .Z(n2767) );
  MUX2_X1 U21719 ( .A(\mem[294][2] ), .B(\mem[295][2] ), .S(n8428), .Z(n2768)
         );
  MUX2_X1 U21720 ( .A(\mem[292][2] ), .B(\mem[293][2] ), .S(n8423), .Z(n2769)
         );
  MUX2_X1 U21721 ( .A(n2769), .B(n2768), .S(n8355), .Z(n2770) );
  MUX2_X1 U21722 ( .A(\mem[290][2] ), .B(\mem[291][2] ), .S(n8424), .Z(n2771)
         );
  MUX2_X1 U21723 ( .A(\mem[288][2] ), .B(\mem[289][2] ), .S(n8425), .Z(n2772)
         );
  MUX2_X1 U21724 ( .A(n2772), .B(n2771), .S(n8291), .Z(n2773) );
  MUX2_X1 U21725 ( .A(n2773), .B(n2770), .S(n8255), .Z(n2774) );
  MUX2_X1 U21726 ( .A(n2774), .B(n2767), .S(n8209), .Z(n2775) );
  MUX2_X1 U21727 ( .A(n2775), .B(n2760), .S(n8193), .Z(n2776) );
  MUX2_X1 U21728 ( .A(\mem[286][2] ), .B(\mem[287][2] ), .S(n8486), .Z(n2777)
         );
  MUX2_X1 U21729 ( .A(\mem[284][2] ), .B(\mem[285][2] ), .S(n8487), .Z(n2778)
         );
  MUX2_X1 U21730 ( .A(n2778), .B(n2777), .S(n8292), .Z(n2779) );
  MUX2_X1 U21731 ( .A(\mem[282][2] ), .B(\mem[283][2] ), .S(n8488), .Z(n2780)
         );
  MUX2_X1 U21732 ( .A(\mem[280][2] ), .B(\mem[281][2] ), .S(n8483), .Z(n2781)
         );
  MUX2_X1 U21733 ( .A(n2781), .B(n2780), .S(n8287), .Z(n2782) );
  MUX2_X1 U21734 ( .A(n2782), .B(n2779), .S(n8255), .Z(n2783) );
  MUX2_X1 U21735 ( .A(\mem[278][2] ), .B(\mem[279][2] ), .S(n8455), .Z(n2784)
         );
  MUX2_X1 U21736 ( .A(\mem[276][2] ), .B(\mem[277][2] ), .S(n8532), .Z(n2785)
         );
  MUX2_X1 U21737 ( .A(n2785), .B(n2784), .S(n8288), .Z(n2786) );
  MUX2_X1 U21738 ( .A(\mem[274][2] ), .B(\mem[275][2] ), .S(n8407), .Z(n2787)
         );
  MUX2_X1 U21739 ( .A(\mem[272][2] ), .B(\mem[273][2] ), .S(n8401), .Z(n2788)
         );
  MUX2_X1 U21740 ( .A(n2788), .B(n2787), .S(n8289), .Z(n2789) );
  MUX2_X1 U21741 ( .A(n2789), .B(n2786), .S(n8255), .Z(n2790) );
  MUX2_X1 U21742 ( .A(n2790), .B(n2783), .S(n8216), .Z(n2791) );
  MUX2_X1 U21743 ( .A(\mem[270][2] ), .B(\mem[271][2] ), .S(n8529), .Z(n2792)
         );
  MUX2_X1 U21744 ( .A(\mem[268][2] ), .B(\mem[269][2] ), .S(n8447), .Z(n2793)
         );
  MUX2_X1 U21745 ( .A(n2793), .B(n2792), .S(N19), .Z(n2794) );
  MUX2_X1 U21746 ( .A(\mem[266][2] ), .B(\mem[267][2] ), .S(n8519), .Z(n2795)
         );
  MUX2_X1 U21747 ( .A(\mem[264][2] ), .B(\mem[265][2] ), .S(n8496), .Z(n2796)
         );
  MUX2_X1 U21748 ( .A(n2796), .B(n2795), .S(n8356), .Z(n2797) );
  MUX2_X1 U21749 ( .A(n2797), .B(n2794), .S(n8255), .Z(n2798) );
  MUX2_X1 U21750 ( .A(\mem[262][2] ), .B(\mem[263][2] ), .S(n8385), .Z(n2799)
         );
  MUX2_X1 U21751 ( .A(\mem[260][2] ), .B(\mem[261][2] ), .S(n8384), .Z(n2800)
         );
  MUX2_X1 U21752 ( .A(n2800), .B(n2799), .S(n8341), .Z(n2801) );
  MUX2_X1 U21753 ( .A(\mem[258][2] ), .B(\mem[259][2] ), .S(n8383), .Z(n2802)
         );
  MUX2_X1 U21754 ( .A(\mem[256][2] ), .B(\mem[257][2] ), .S(n8373), .Z(n2803)
         );
  MUX2_X1 U21755 ( .A(n2803), .B(n2802), .S(n8266), .Z(n2804) );
  MUX2_X1 U21756 ( .A(n2804), .B(n2801), .S(n8255), .Z(n2805) );
  MUX2_X1 U21757 ( .A(n2805), .B(n2798), .S(n8198), .Z(n2806) );
  MUX2_X1 U21758 ( .A(n2806), .B(n2791), .S(n8196), .Z(n2807) );
  MUX2_X1 U21759 ( .A(n2807), .B(n2776), .S(n8183), .Z(n2808) );
  MUX2_X1 U21760 ( .A(n2808), .B(n2745), .S(n8178), .Z(n2809) );
  MUX2_X1 U21761 ( .A(n2809), .B(n2682), .S(n8177), .Z(n2810) );
  MUX2_X1 U21762 ( .A(\mem[254][2] ), .B(\mem[255][2] ), .S(n8437), .Z(n2811)
         );
  MUX2_X1 U21763 ( .A(\mem[252][2] ), .B(\mem[253][2] ), .S(n8411), .Z(n2812)
         );
  MUX2_X1 U21764 ( .A(n2812), .B(n2811), .S(n8336), .Z(n2813) );
  MUX2_X1 U21765 ( .A(\mem[250][2] ), .B(\mem[251][2] ), .S(n8412), .Z(n2814)
         );
  MUX2_X1 U21766 ( .A(\mem[248][2] ), .B(\mem[249][2] ), .S(n8413), .Z(n2815)
         );
  MUX2_X1 U21767 ( .A(n2815), .B(n2814), .S(n8337), .Z(n2816) );
  MUX2_X1 U21768 ( .A(n2816), .B(n2813), .S(n8256), .Z(n2817) );
  MUX2_X1 U21769 ( .A(\mem[246][2] ), .B(\mem[247][2] ), .S(n8420), .Z(n2818)
         );
  MUX2_X1 U21770 ( .A(\mem[244][2] ), .B(\mem[245][2] ), .S(n8410), .Z(n2819)
         );
  MUX2_X1 U21771 ( .A(n2819), .B(n2818), .S(n8344), .Z(n2820) );
  MUX2_X1 U21772 ( .A(\mem[242][2] ), .B(\mem[243][2] ), .S(N18), .Z(n2821) );
  MUX2_X1 U21773 ( .A(\mem[240][2] ), .B(\mem[241][2] ), .S(n8381), .Z(n2822)
         );
  MUX2_X1 U21774 ( .A(n2822), .B(n2821), .S(n8345), .Z(n2823) );
  MUX2_X1 U21775 ( .A(n2823), .B(n2820), .S(n8256), .Z(n2824) );
  MUX2_X1 U21776 ( .A(n2824), .B(n2817), .S(n8217), .Z(n2825) );
  MUX2_X1 U21777 ( .A(\mem[238][2] ), .B(\mem[239][2] ), .S(n8391), .Z(n2826)
         );
  MUX2_X1 U21778 ( .A(\mem[236][2] ), .B(\mem[237][2] ), .S(n8357), .Z(n2827)
         );
  MUX2_X1 U21779 ( .A(n2827), .B(n2826), .S(n8346), .Z(n2828) );
  MUX2_X1 U21780 ( .A(\mem[234][2] ), .B(\mem[235][2] ), .S(n8406), .Z(n2829)
         );
  MUX2_X1 U21781 ( .A(\mem[232][2] ), .B(\mem[233][2] ), .S(n8415), .Z(n2830)
         );
  MUX2_X1 U21782 ( .A(n2830), .B(n2829), .S(n8341), .Z(n2831) );
  MUX2_X1 U21783 ( .A(n2831), .B(n2828), .S(n8256), .Z(n2832) );
  MUX2_X1 U21784 ( .A(\mem[230][2] ), .B(\mem[231][2] ), .S(n8515), .Z(n2833)
         );
  MUX2_X1 U21785 ( .A(\mem[228][2] ), .B(\mem[229][2] ), .S(n8522), .Z(n2834)
         );
  MUX2_X1 U21786 ( .A(n2834), .B(n2833), .S(n8342), .Z(n2835) );
  MUX2_X1 U21787 ( .A(\mem[226][2] ), .B(\mem[227][2] ), .S(n8523), .Z(n2836)
         );
  MUX2_X1 U21788 ( .A(\mem[224][2] ), .B(\mem[225][2] ), .S(n8524), .Z(n2837)
         );
  MUX2_X1 U21789 ( .A(n2837), .B(n2836), .S(n8343), .Z(n2838) );
  MUX2_X1 U21790 ( .A(n2838), .B(n2835), .S(n8256), .Z(n2839) );
  MUX2_X1 U21791 ( .A(n2839), .B(n2832), .S(n8218), .Z(n2840) );
  MUX2_X1 U21792 ( .A(n2840), .B(n2825), .S(n8187), .Z(n2841) );
  MUX2_X1 U21793 ( .A(\mem[222][2] ), .B(\mem[223][2] ), .S(n8519), .Z(n2842)
         );
  MUX2_X1 U21794 ( .A(\mem[220][2] ), .B(\mem[221][2] ), .S(n8520), .Z(n2843)
         );
  MUX2_X1 U21795 ( .A(n2843), .B(n2842), .S(n8350), .Z(n2844) );
  MUX2_X1 U21796 ( .A(\mem[218][2] ), .B(\mem[219][2] ), .S(n8521), .Z(n2845)
         );
  MUX2_X1 U21797 ( .A(\mem[216][2] ), .B(\mem[217][2] ), .S(n8528), .Z(n2846)
         );
  MUX2_X1 U21798 ( .A(n2846), .B(n2845), .S(n8351), .Z(n2847) );
  MUX2_X1 U21799 ( .A(n2847), .B(n2844), .S(n8256), .Z(n2848) );
  MUX2_X1 U21800 ( .A(\mem[214][2] ), .B(\mem[215][2] ), .S(n8529), .Z(n2849)
         );
  MUX2_X1 U21801 ( .A(\mem[212][2] ), .B(\mem[213][2] ), .S(n8530), .Z(n2850)
         );
  MUX2_X1 U21802 ( .A(n2850), .B(n2849), .S(n8352), .Z(n2851) );
  MUX2_X1 U21803 ( .A(\mem[210][2] ), .B(\mem[211][2] ), .S(n8525), .Z(n2852)
         );
  MUX2_X1 U21804 ( .A(\mem[208][2] ), .B(\mem[209][2] ), .S(n8526), .Z(n2853)
         );
  MUX2_X1 U21805 ( .A(n2853), .B(n2852), .S(n8347), .Z(n2854) );
  MUX2_X1 U21806 ( .A(n2854), .B(n2851), .S(n8256), .Z(n2855) );
  MUX2_X1 U21807 ( .A(n2855), .B(n2848), .S(n8210), .Z(n2856) );
  MUX2_X1 U21808 ( .A(\mem[206][2] ), .B(\mem[207][2] ), .S(n8374), .Z(n2857)
         );
  MUX2_X1 U21809 ( .A(\mem[204][2] ), .B(\mem[205][2] ), .S(n8358), .Z(n2858)
         );
  MUX2_X1 U21810 ( .A(n2858), .B(n2857), .S(n8309), .Z(n2859) );
  MUX2_X1 U21811 ( .A(\mem[202][2] ), .B(\mem[203][2] ), .S(n8360), .Z(n2860)
         );
  MUX2_X1 U21812 ( .A(\mem[200][2] ), .B(\mem[201][2] ), .S(n8361), .Z(n2861)
         );
  MUX2_X1 U21813 ( .A(n2861), .B(n2860), .S(n8291), .Z(n2862) );
  MUX2_X1 U21814 ( .A(n2862), .B(n2859), .S(n8256), .Z(n2863) );
  MUX2_X1 U21815 ( .A(\mem[198][2] ), .B(\mem[199][2] ), .S(n8539), .Z(n2864)
         );
  MUX2_X1 U21816 ( .A(\mem[196][2] ), .B(\mem[197][2] ), .S(n8362), .Z(n2865)
         );
  MUX2_X1 U21817 ( .A(n2865), .B(n2864), .S(n8283), .Z(n2866) );
  MUX2_X1 U21818 ( .A(\mem[194][2] ), .B(\mem[195][2] ), .S(n8363), .Z(n2867)
         );
  MUX2_X1 U21819 ( .A(\mem[192][2] ), .B(\mem[193][2] ), .S(n8364), .Z(n2868)
         );
  MUX2_X1 U21820 ( .A(n2868), .B(n2867), .S(n8279), .Z(n2869) );
  MUX2_X1 U21821 ( .A(n2869), .B(n2866), .S(n8256), .Z(n2870) );
  MUX2_X1 U21822 ( .A(n2870), .B(n2863), .S(n8210), .Z(n2871) );
  MUX2_X1 U21823 ( .A(n2871), .B(n2856), .S(n8196), .Z(n2872) );
  MUX2_X1 U21824 ( .A(n2872), .B(n2841), .S(n8184), .Z(n2873) );
  MUX2_X1 U21825 ( .A(\mem[190][2] ), .B(\mem[191][2] ), .S(n8425), .Z(n2874)
         );
  MUX2_X1 U21826 ( .A(\mem[188][2] ), .B(\mem[189][2] ), .S(n8412), .Z(n2875)
         );
  MUX2_X1 U21827 ( .A(n2875), .B(n2874), .S(n8311), .Z(n2876) );
  MUX2_X1 U21828 ( .A(\mem[186][2] ), .B(\mem[187][2] ), .S(n8413), .Z(n2877)
         );
  MUX2_X1 U21829 ( .A(\mem[184][2] ), .B(\mem[185][2] ), .S(n8420), .Z(n2878)
         );
  MUX2_X1 U21830 ( .A(n2878), .B(n2877), .S(n8296), .Z(n2879) );
  MUX2_X1 U21831 ( .A(n2879), .B(n2876), .S(n8256), .Z(n2880) );
  MUX2_X1 U21832 ( .A(\mem[182][2] ), .B(\mem[183][2] ), .S(n8471), .Z(n2881)
         );
  MUX2_X1 U21833 ( .A(\mem[180][2] ), .B(\mem[181][2] ), .S(n8472), .Z(n2882)
         );
  MUX2_X1 U21834 ( .A(n2882), .B(n2881), .S(n8268), .Z(n2883) );
  MUX2_X1 U21835 ( .A(\mem[178][2] ), .B(\mem[179][2] ), .S(n8473), .Z(n2884)
         );
  MUX2_X1 U21836 ( .A(\mem[176][2] ), .B(\mem[177][2] ), .S(n8480), .Z(n2885)
         );
  MUX2_X1 U21837 ( .A(n2885), .B(n2884), .S(n8293), .Z(n2886) );
  MUX2_X1 U21838 ( .A(n2886), .B(n2883), .S(n8256), .Z(n2887) );
  MUX2_X1 U21839 ( .A(n2887), .B(n2880), .S(n8203), .Z(n2888) );
  MUX2_X1 U21840 ( .A(\mem[174][2] ), .B(\mem[175][2] ), .S(n8481), .Z(n2889)
         );
  MUX2_X1 U21841 ( .A(\mem[172][2] ), .B(\mem[173][2] ), .S(n8482), .Z(n2890)
         );
  MUX2_X1 U21842 ( .A(n2890), .B(n2889), .S(n8307), .Z(n2891) );
  MUX2_X1 U21843 ( .A(\mem[170][2] ), .B(\mem[171][2] ), .S(n8477), .Z(n2892)
         );
  MUX2_X1 U21844 ( .A(\mem[168][2] ), .B(\mem[169][2] ), .S(n8478), .Z(n2893)
         );
  MUX2_X1 U21845 ( .A(n2893), .B(n2892), .S(n8345), .Z(n2894) );
  MUX2_X1 U21846 ( .A(n2894), .B(n2891), .S(n8256), .Z(n2895) );
  MUX2_X1 U21847 ( .A(\mem[166][2] ), .B(\mem[167][2] ), .S(n8479), .Z(n2896)
         );
  MUX2_X1 U21848 ( .A(\mem[164][2] ), .B(\mem[165][2] ), .S(n8382), .Z(n2897)
         );
  MUX2_X1 U21849 ( .A(n2897), .B(n2896), .S(n8292), .Z(n2898) );
  MUX2_X1 U21850 ( .A(\mem[162][2] ), .B(\mem[163][2] ), .S(n8379), .Z(n2899)
         );
  MUX2_X1 U21851 ( .A(\mem[160][2] ), .B(\mem[161][2] ), .S(n8378), .Z(n2900)
         );
  MUX2_X1 U21852 ( .A(n2900), .B(n2899), .S(n8287), .Z(n2901) );
  MUX2_X1 U21853 ( .A(n2901), .B(n2898), .S(n8256), .Z(n2902) );
  MUX2_X1 U21854 ( .A(n2902), .B(n2895), .S(n8210), .Z(n2903) );
  MUX2_X1 U21855 ( .A(n2903), .B(n2888), .S(n8195), .Z(n2904) );
  MUX2_X1 U21856 ( .A(\mem[158][2] ), .B(\mem[159][2] ), .S(n8462), .Z(n2905)
         );
  MUX2_X1 U21857 ( .A(\mem[156][2] ), .B(\mem[157][2] ), .S(n8463), .Z(n2906)
         );
  MUX2_X1 U21858 ( .A(n2906), .B(n2905), .S(N19), .Z(n2907) );
  MUX2_X1 U21859 ( .A(\mem[154][2] ), .B(\mem[155][2] ), .S(n8464), .Z(n2908)
         );
  MUX2_X1 U21860 ( .A(\mem[152][2] ), .B(\mem[153][2] ), .S(n8459), .Z(n2909)
         );
  MUX2_X1 U21861 ( .A(n2909), .B(n2908), .S(n8346), .Z(n2910) );
  MUX2_X1 U21862 ( .A(n2910), .B(n2907), .S(n8257), .Z(n2911) );
  MUX2_X1 U21863 ( .A(\mem[150][2] ), .B(\mem[151][2] ), .S(n8460), .Z(n2912)
         );
  MUX2_X1 U21864 ( .A(\mem[148][2] ), .B(\mem[149][2] ), .S(n8461), .Z(n2913)
         );
  MUX2_X1 U21865 ( .A(n2913), .B(n2912), .S(n8323), .Z(n2914) );
  MUX2_X1 U21866 ( .A(\mem[146][2] ), .B(\mem[147][2] ), .S(n8468), .Z(n2915)
         );
  MUX2_X1 U21867 ( .A(\mem[144][2] ), .B(\mem[145][2] ), .S(n8469), .Z(n2916)
         );
  MUX2_X1 U21868 ( .A(n2916), .B(n2915), .S(n8291), .Z(n2917) );
  MUX2_X1 U21869 ( .A(n2917), .B(n2914), .S(n8257), .Z(n2918) );
  MUX2_X1 U21870 ( .A(n2918), .B(n2911), .S(n8201), .Z(n2919) );
  MUX2_X1 U21871 ( .A(\mem[142][2] ), .B(\mem[143][2] ), .S(n8470), .Z(n2920)
         );
  MUX2_X1 U21872 ( .A(\mem[140][2] ), .B(\mem[141][2] ), .S(n8465), .Z(n2921)
         );
  MUX2_X1 U21873 ( .A(n2921), .B(n2920), .S(n8292), .Z(n2922) );
  MUX2_X1 U21874 ( .A(\mem[138][2] ), .B(\mem[139][2] ), .S(n8466), .Z(n2923)
         );
  MUX2_X1 U21875 ( .A(\mem[136][2] ), .B(\mem[137][2] ), .S(n8467), .Z(n2924)
         );
  MUX2_X1 U21876 ( .A(n2924), .B(n2923), .S(n8287), .Z(n2925) );
  MUX2_X1 U21877 ( .A(n2925), .B(n2922), .S(n8257), .Z(n2926) );
  MUX2_X1 U21878 ( .A(\mem[134][2] ), .B(\mem[135][2] ), .S(n8416), .Z(n2927)
         );
  MUX2_X1 U21879 ( .A(\mem[132][2] ), .B(\mem[133][2] ), .S(n8361), .Z(n2928)
         );
  MUX2_X1 U21880 ( .A(n2928), .B(n2927), .S(n8288), .Z(n2929) );
  MUX2_X1 U21881 ( .A(\mem[130][2] ), .B(\mem[131][2] ), .S(n8430), .Z(n2930)
         );
  MUX2_X1 U21882 ( .A(\mem[128][2] ), .B(\mem[129][2] ), .S(n8432), .Z(n2931)
         );
  MUX2_X1 U21883 ( .A(n2931), .B(n2930), .S(n8289), .Z(n2932) );
  MUX2_X1 U21884 ( .A(n2932), .B(n2929), .S(n8257), .Z(n2933) );
  MUX2_X1 U21885 ( .A(n2933), .B(n2926), .S(n8200), .Z(n2934) );
  MUX2_X1 U21886 ( .A(n2934), .B(n2919), .S(n8195), .Z(n2935) );
  MUX2_X1 U21887 ( .A(n2935), .B(n2904), .S(n8184), .Z(n2936) );
  MUX2_X1 U21888 ( .A(n2936), .B(n2873), .S(N24), .Z(n2937) );
  MUX2_X1 U21889 ( .A(\mem[126][2] ), .B(\mem[127][2] ), .S(n8371), .Z(n2938)
         );
  MUX2_X1 U21890 ( .A(\mem[124][2] ), .B(\mem[125][2] ), .S(n8459), .Z(n2939)
         );
  MUX2_X1 U21891 ( .A(n2939), .B(n2938), .S(n8296), .Z(n2940) );
  MUX2_X1 U21892 ( .A(\mem[122][2] ), .B(\mem[123][2] ), .S(n8466), .Z(n2941)
         );
  MUX2_X1 U21893 ( .A(\mem[120][2] ), .B(\mem[121][2] ), .S(n8444), .Z(n2942)
         );
  MUX2_X1 U21894 ( .A(n2942), .B(n2941), .S(n8297), .Z(n2943) );
  MUX2_X1 U21895 ( .A(n2943), .B(n2940), .S(n8257), .Z(n2944) );
  MUX2_X1 U21896 ( .A(\mem[118][2] ), .B(\mem[119][2] ), .S(n8536), .Z(n2945)
         );
  MUX2_X1 U21897 ( .A(\mem[116][2] ), .B(\mem[117][2] ), .S(n8364), .Z(n2946)
         );
  MUX2_X1 U21898 ( .A(n2946), .B(n2945), .S(n8298), .Z(n2947) );
  MUX2_X1 U21899 ( .A(\mem[114][2] ), .B(\mem[115][2] ), .S(n8367), .Z(n2948)
         );
  MUX2_X1 U21900 ( .A(\mem[112][2] ), .B(\mem[113][2] ), .S(n8405), .Z(n2949)
         );
  MUX2_X1 U21901 ( .A(n2949), .B(n2948), .S(n8293), .Z(n2950) );
  MUX2_X1 U21902 ( .A(n2950), .B(n2947), .S(n8257), .Z(n2951) );
  MUX2_X1 U21903 ( .A(n2951), .B(n2944), .S(n8218), .Z(n2952) );
  MUX2_X1 U21904 ( .A(\mem[110][2] ), .B(\mem[111][2] ), .S(n8358), .Z(n2953)
         );
  MUX2_X1 U21905 ( .A(\mem[108][2] ), .B(\mem[109][2] ), .S(n8375), .Z(n2954)
         );
  MUX2_X1 U21906 ( .A(n2954), .B(n2953), .S(n8321), .Z(n2955) );
  MUX2_X1 U21907 ( .A(\mem[106][2] ), .B(\mem[107][2] ), .S(n8394), .Z(n2956)
         );
  MUX2_X1 U21908 ( .A(\mem[104][2] ), .B(\mem[105][2] ), .S(n8468), .Z(n2957)
         );
  MUX2_X1 U21909 ( .A(n2957), .B(n2956), .S(n8277), .Z(n2958) );
  MUX2_X1 U21910 ( .A(n2958), .B(n2955), .S(n8257), .Z(n2959) );
  MUX2_X1 U21911 ( .A(\mem[102][2] ), .B(\mem[103][2] ), .S(n8450), .Z(n2960)
         );
  MUX2_X1 U21912 ( .A(\mem[100][2] ), .B(\mem[101][2] ), .S(n8520), .Z(n2961)
         );
  MUX2_X1 U21913 ( .A(n2961), .B(n2960), .S(n8276), .Z(n2962) );
  MUX2_X1 U21914 ( .A(\mem[98][2] ), .B(\mem[99][2] ), .S(n8506), .Z(n2963) );
  MUX2_X1 U21915 ( .A(\mem[96][2] ), .B(\mem[97][2] ), .S(n8487), .Z(n2964) );
  MUX2_X1 U21916 ( .A(n2964), .B(n2963), .S(n8294), .Z(n2965) );
  MUX2_X1 U21917 ( .A(n2965), .B(n2962), .S(n8257), .Z(n2966) );
  MUX2_X1 U21918 ( .A(n2966), .B(n2959), .S(n8202), .Z(n2967) );
  MUX2_X1 U21919 ( .A(n2967), .B(n2952), .S(n8190), .Z(n2968) );
  MUX2_X1 U21920 ( .A(\mem[94][2] ), .B(\mem[95][2] ), .S(n8376), .Z(n2969) );
  MUX2_X1 U21921 ( .A(\mem[92][2] ), .B(\mem[93][2] ), .S(n8373), .Z(n2970) );
  MUX2_X1 U21922 ( .A(n2970), .B(n2969), .S(n8308), .Z(n2971) );
  MUX2_X1 U21923 ( .A(\mem[90][2] ), .B(\mem[91][2] ), .S(n8403), .Z(n2972) );
  MUX2_X1 U21924 ( .A(\mem[88][2] ), .B(\mem[89][2] ), .S(n8510), .Z(n2973) );
  MUX2_X1 U21925 ( .A(n2973), .B(n2972), .S(n8313), .Z(n2974) );
  MUX2_X1 U21926 ( .A(n2974), .B(n2971), .S(n8257), .Z(n2975) );
  MUX2_X1 U21927 ( .A(\mem[86][2] ), .B(\mem[87][2] ), .S(n8467), .Z(n2976) );
  MUX2_X1 U21928 ( .A(\mem[84][2] ), .B(\mem[85][2] ), .S(n8474), .Z(n2977) );
  MUX2_X1 U21929 ( .A(n2977), .B(n2976), .S(n8275), .Z(n2978) );
  MUX2_X1 U21930 ( .A(\mem[82][2] ), .B(\mem[83][2] ), .S(n8475), .Z(n2979) );
  MUX2_X1 U21931 ( .A(\mem[80][2] ), .B(\mem[81][2] ), .S(n8476), .Z(n2980) );
  MUX2_X1 U21932 ( .A(n2980), .B(n2979), .S(n8283), .Z(n2981) );
  MUX2_X1 U21933 ( .A(n2981), .B(n2978), .S(n8257), .Z(n2982) );
  MUX2_X1 U21934 ( .A(n2982), .B(n2975), .S(n8203), .Z(n2983) );
  MUX2_X1 U21935 ( .A(\mem[78][2] ), .B(\mem[79][2] ), .S(n8471), .Z(n2984) );
  MUX2_X1 U21936 ( .A(\mem[76][2] ), .B(\mem[77][2] ), .S(n8472), .Z(n2985) );
  MUX2_X1 U21937 ( .A(n2985), .B(n2984), .S(n8342), .Z(n2986) );
  MUX2_X1 U21938 ( .A(\mem[74][2] ), .B(\mem[75][2] ), .S(n8473), .Z(n2987) );
  MUX2_X1 U21939 ( .A(\mem[72][2] ), .B(\mem[73][2] ), .S(n8480), .Z(n2988) );
  MUX2_X1 U21940 ( .A(n2988), .B(n2987), .S(n8333), .Z(n2989) );
  MUX2_X1 U21941 ( .A(n2989), .B(n2986), .S(n8257), .Z(n2990) );
  MUX2_X1 U21942 ( .A(\mem[70][2] ), .B(\mem[71][2] ), .S(n8481), .Z(n2991) );
  MUX2_X1 U21943 ( .A(\mem[68][2] ), .B(\mem[69][2] ), .S(n8482), .Z(n2992) );
  MUX2_X1 U21944 ( .A(n2992), .B(n2991), .S(n8312), .Z(n2993) );
  MUX2_X1 U21945 ( .A(\mem[66][2] ), .B(\mem[67][2] ), .S(n8477), .Z(n2994) );
  MUX2_X1 U21946 ( .A(\mem[64][2] ), .B(\mem[65][2] ), .S(n8478), .Z(n2995) );
  MUX2_X1 U21947 ( .A(n2995), .B(n2994), .S(n8297), .Z(n2996) );
  MUX2_X1 U21948 ( .A(n2996), .B(n2993), .S(n8257), .Z(n2997) );
  MUX2_X1 U21949 ( .A(n2997), .B(n2990), .S(n8204), .Z(n2998) );
  MUX2_X1 U21950 ( .A(n2998), .B(n2983), .S(n8196), .Z(n2999) );
  MUX2_X1 U21951 ( .A(n2999), .B(n2968), .S(n8184), .Z(n3000) );
  MUX2_X1 U21952 ( .A(\mem[62][2] ), .B(\mem[63][2] ), .S(n8403), .Z(n3001) );
  MUX2_X1 U21953 ( .A(\mem[60][2] ), .B(\mem[61][2] ), .S(n8393), .Z(n3002) );
  MUX2_X1 U21954 ( .A(n3002), .B(n3001), .S(n8312), .Z(n3003) );
  MUX2_X1 U21955 ( .A(\mem[58][2] ), .B(\mem[59][2] ), .S(n8394), .Z(n3004) );
  MUX2_X1 U21956 ( .A(\mem[56][2] ), .B(\mem[57][2] ), .S(n8390), .Z(n3005) );
  MUX2_X1 U21957 ( .A(n3005), .B(n3004), .S(n8327), .Z(n3006) );
  MUX2_X1 U21958 ( .A(n3006), .B(n3003), .S(n8258), .Z(n3007) );
  MUX2_X1 U21959 ( .A(\mem[54][2] ), .B(\mem[55][2] ), .S(n8391), .Z(n3008) );
  MUX2_X1 U21960 ( .A(\mem[52][2] ), .B(\mem[53][2] ), .S(n8392), .Z(n3009) );
  MUX2_X1 U21961 ( .A(n3009), .B(n3008), .S(n8295), .Z(n3010) );
  MUX2_X1 U21962 ( .A(\mem[50][2] ), .B(\mem[51][2] ), .S(n8389), .Z(n3011) );
  MUX2_X1 U21963 ( .A(\mem[48][2] ), .B(\mem[49][2] ), .S(n8537), .Z(n3012) );
  MUX2_X1 U21964 ( .A(n3012), .B(n3011), .S(n8282), .Z(n3013) );
  MUX2_X1 U21965 ( .A(n3013), .B(n3010), .S(n8258), .Z(n3014) );
  MUX2_X1 U21966 ( .A(n3014), .B(n3007), .S(n8214), .Z(n3015) );
  MUX2_X1 U21967 ( .A(\mem[46][2] ), .B(\mem[47][2] ), .S(n8388), .Z(n3016) );
  MUX2_X1 U21968 ( .A(\mem[44][2] ), .B(\mem[45][2] ), .S(n8386), .Z(n3017) );
  MUX2_X1 U21969 ( .A(n3017), .B(n3016), .S(n8281), .Z(n3018) );
  MUX2_X1 U21970 ( .A(\mem[42][2] ), .B(\mem[43][2] ), .S(n8365), .Z(n3019) );
  MUX2_X1 U21971 ( .A(\mem[40][2] ), .B(\mem[41][2] ), .S(n8387), .Z(n3020) );
  MUX2_X1 U21972 ( .A(n3020), .B(n3019), .S(n8347), .Z(n3021) );
  MUX2_X1 U21973 ( .A(n3021), .B(n3018), .S(n8258), .Z(n3022) );
  MUX2_X1 U21974 ( .A(\mem[38][2] ), .B(\mem[39][2] ), .S(n8388), .Z(n3023) );
  MUX2_X1 U21975 ( .A(\mem[36][2] ), .B(\mem[37][2] ), .S(n8365), .Z(n3024) );
  MUX2_X1 U21976 ( .A(n3024), .B(n3023), .S(n8332), .Z(n3025) );
  MUX2_X1 U21977 ( .A(\mem[34][2] ), .B(\mem[35][2] ), .S(n8387), .Z(n3026) );
  MUX2_X1 U21978 ( .A(\mem[32][2] ), .B(\mem[33][2] ), .S(n8386), .Z(n3027) );
  MUX2_X1 U21979 ( .A(n3027), .B(n3026), .S(n8283), .Z(n3028) );
  MUX2_X1 U21980 ( .A(n3028), .B(n3025), .S(n8258), .Z(n3029) );
  MUX2_X1 U21981 ( .A(n3029), .B(n3022), .S(n8215), .Z(n3030) );
  MUX2_X1 U21982 ( .A(n3030), .B(n3015), .S(N22), .Z(n3031) );
  MUX2_X1 U21983 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n8357), .Z(n3032) );
  MUX2_X1 U21984 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n8389), .Z(n3033) );
  MUX2_X1 U21985 ( .A(n3033), .B(n3032), .S(n8312), .Z(n3034) );
  MUX2_X1 U21986 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n8388), .Z(n3035) );
  MUX2_X1 U21987 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n8365), .Z(n3036) );
  MUX2_X1 U21988 ( .A(n3036), .B(n3035), .S(n8348), .Z(n3037) );
  MUX2_X1 U21989 ( .A(n3037), .B(n3034), .S(n8258), .Z(n3038) );
  MUX2_X1 U21990 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n8387), .Z(n3039) );
  MUX2_X1 U21991 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n8386), .Z(n3040) );
  MUX2_X1 U21992 ( .A(n3040), .B(n3039), .S(n8333), .Z(n3041) );
  MUX2_X1 U21993 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n8537), .Z(n3042) );
  MUX2_X1 U21994 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n8357), .Z(n3043) );
  MUX2_X1 U21995 ( .A(n3043), .B(n3042), .S(n8288), .Z(n3044) );
  MUX2_X1 U21996 ( .A(n3044), .B(n3041), .S(n8258), .Z(n3045) );
  MUX2_X1 U21997 ( .A(n3045), .B(n3038), .S(n8211), .Z(n3046) );
  MUX2_X1 U21998 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n8357), .Z(n3047) );
  MUX2_X1 U21999 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n8537), .Z(n3048) );
  MUX2_X1 U22000 ( .A(n3048), .B(n3047), .S(n8327), .Z(n3049) );
  MUX2_X1 U22001 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n8388), .Z(n3050) );
  MUX2_X1 U22002 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n8365), .Z(n3051) );
  MUX2_X1 U22003 ( .A(n3051), .B(n3050), .S(n8299), .Z(n3052) );
  MUX2_X1 U22004 ( .A(n3052), .B(n3049), .S(n8258), .Z(n3053) );
  MUX2_X1 U22005 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n8387), .Z(n3054) );
  MUX2_X1 U22006 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n8386), .Z(n3055) );
  MUX2_X1 U22007 ( .A(n3055), .B(n3054), .S(n8310), .Z(n3056) );
  MUX2_X1 U22008 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n8357), .Z(n3057) );
  MUX2_X1 U22009 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n8389), .Z(n3058) );
  MUX2_X1 U22010 ( .A(n3058), .B(n3057), .S(n8280), .Z(n3059) );
  MUX2_X1 U22011 ( .A(n3059), .B(n3056), .S(n8258), .Z(n3060) );
  MUX2_X1 U22012 ( .A(n3060), .B(n3053), .S(n8216), .Z(n3061) );
  MUX2_X1 U22013 ( .A(n3061), .B(n3046), .S(n8190), .Z(n3062) );
  MUX2_X1 U22014 ( .A(n3062), .B(n3031), .S(n8184), .Z(n3063) );
  MUX2_X1 U22015 ( .A(n3063), .B(n3000), .S(n8179), .Z(n3064) );
  MUX2_X1 U22016 ( .A(n3064), .B(n2937), .S(n8177), .Z(n3065) );
  MUX2_X1 U22017 ( .A(n3065), .B(n2810), .S(N26), .Z(n3066) );
  MUX2_X1 U22018 ( .A(n3066), .B(n2555), .S(N27), .Z(N33) );
  MUX2_X1 U22019 ( .A(\mem[1022][3] ), .B(\mem[1023][3] ), .S(n8537), .Z(n3067) );
  MUX2_X1 U22020 ( .A(\mem[1020][3] ), .B(\mem[1021][3] ), .S(n8388), .Z(n3068) );
  MUX2_X1 U22021 ( .A(n3068), .B(n3067), .S(n8279), .Z(n3069) );
  MUX2_X1 U22022 ( .A(\mem[1018][3] ), .B(\mem[1019][3] ), .S(n8365), .Z(n3070) );
  MUX2_X1 U22023 ( .A(\mem[1016][3] ), .B(\mem[1017][3] ), .S(n8387), .Z(n3071) );
  MUX2_X1 U22024 ( .A(n3071), .B(n3070), .S(n8277), .Z(n3072) );
  MUX2_X1 U22025 ( .A(n3072), .B(n3069), .S(n8258), .Z(n3073) );
  MUX2_X1 U22026 ( .A(\mem[1014][3] ), .B(\mem[1015][3] ), .S(n8363), .Z(n3074) );
  MUX2_X1 U22027 ( .A(\mem[1012][3] ), .B(\mem[1013][3] ), .S(n8406), .Z(n3075) );
  MUX2_X1 U22028 ( .A(n3075), .B(n3074), .S(n8276), .Z(n3076) );
  MUX2_X1 U22029 ( .A(\mem[1010][3] ), .B(\mem[1011][3] ), .S(n8469), .Z(n3077) );
  MUX2_X1 U22030 ( .A(\mem[1008][3] ), .B(\mem[1009][3] ), .S(n8404), .Z(n3078) );
  MUX2_X1 U22031 ( .A(n3078), .B(n3077), .S(n8271), .Z(n3079) );
  MUX2_X1 U22032 ( .A(n3079), .B(n3076), .S(n8258), .Z(n3080) );
  MUX2_X1 U22033 ( .A(n3080), .B(n3073), .S(n8217), .Z(n3081) );
  MUX2_X1 U22034 ( .A(\mem[1006][3] ), .B(\mem[1007][3] ), .S(n8483), .Z(n3082) );
  MUX2_X1 U22035 ( .A(\mem[1004][3] ), .B(\mem[1005][3] ), .S(n8411), .Z(n3083) );
  MUX2_X1 U22036 ( .A(n3083), .B(n3082), .S(n8268), .Z(n3084) );
  MUX2_X1 U22037 ( .A(\mem[1002][3] ), .B(\mem[1003][3] ), .S(n8401), .Z(n3085) );
  MUX2_X1 U22038 ( .A(\mem[1000][3] ), .B(\mem[1001][3] ), .S(n8526), .Z(n3086) );
  MUX2_X1 U22039 ( .A(n3086), .B(n3085), .S(n8270), .Z(n3087) );
  MUX2_X1 U22040 ( .A(n3087), .B(n3084), .S(n8258), .Z(n3088) );
  MUX2_X1 U22041 ( .A(\mem[998][3] ), .B(\mem[999][3] ), .S(n8508), .Z(n3089)
         );
  MUX2_X1 U22042 ( .A(\mem[996][3] ), .B(\mem[997][3] ), .S(n8491), .Z(n3090)
         );
  MUX2_X1 U22043 ( .A(n3090), .B(n3089), .S(n8311), .Z(n3091) );
  MUX2_X1 U22044 ( .A(\mem[994][3] ), .B(\mem[995][3] ), .S(n8480), .Z(n3092)
         );
  MUX2_X1 U22045 ( .A(\mem[992][3] ), .B(\mem[993][3] ), .S(n8437), .Z(n3093)
         );
  MUX2_X1 U22046 ( .A(n3093), .B(n3092), .S(n8280), .Z(n3094) );
  MUX2_X1 U22047 ( .A(n3094), .B(n3091), .S(n8258), .Z(n3095) );
  MUX2_X1 U22048 ( .A(n3095), .B(n3088), .S(n8218), .Z(n3096) );
  MUX2_X1 U22049 ( .A(n3096), .B(n3081), .S(n8188), .Z(n3097) );
  MUX2_X1 U22050 ( .A(\mem[990][3] ), .B(\mem[991][3] ), .S(n8376), .Z(n3098)
         );
  MUX2_X1 U22051 ( .A(\mem[988][3] ), .B(\mem[989][3] ), .S(n8469), .Z(n3099)
         );
  MUX2_X1 U22052 ( .A(n3099), .B(n3098), .S(n8290), .Z(n3100) );
  MUX2_X1 U22053 ( .A(\mem[986][3] ), .B(\mem[987][3] ), .S(n8357), .Z(n3101)
         );
  MUX2_X1 U22054 ( .A(\mem[984][3] ), .B(\mem[985][3] ), .S(n8391), .Z(n3102)
         );
  MUX2_X1 U22055 ( .A(n3102), .B(n3101), .S(n8324), .Z(n3103) );
  MUX2_X1 U22056 ( .A(n3103), .B(n3100), .S(n8259), .Z(n3104) );
  MUX2_X1 U22057 ( .A(\mem[982][3] ), .B(\mem[983][3] ), .S(n8512), .Z(n3105)
         );
  MUX2_X1 U22058 ( .A(\mem[980][3] ), .B(\mem[981][3] ), .S(n8490), .Z(n3106)
         );
  MUX2_X1 U22059 ( .A(n3106), .B(n3105), .S(n8282), .Z(n3107) );
  MUX2_X1 U22060 ( .A(\mem[978][3] ), .B(\mem[979][3] ), .S(n8480), .Z(n3108)
         );
  MUX2_X1 U22061 ( .A(\mem[976][3] ), .B(\mem[977][3] ), .S(n8421), .Z(n3109)
         );
  MUX2_X1 U22062 ( .A(n3109), .B(n3108), .S(n8281), .Z(n3110) );
  MUX2_X1 U22063 ( .A(n3110), .B(n3107), .S(n8259), .Z(n3111) );
  MUX2_X1 U22064 ( .A(n3111), .B(n3104), .S(n8201), .Z(n3112) );
  MUX2_X1 U22065 ( .A(\mem[974][3] ), .B(\mem[975][3] ), .S(n8442), .Z(n3113)
         );
  MUX2_X1 U22066 ( .A(\mem[972][3] ), .B(\mem[973][3] ), .S(n8474), .Z(n3114)
         );
  MUX2_X1 U22067 ( .A(n3114), .B(n3113), .S(n8341), .Z(n3115) );
  MUX2_X1 U22068 ( .A(\mem[970][3] ), .B(\mem[971][3] ), .S(n8388), .Z(n3116)
         );
  MUX2_X1 U22069 ( .A(\mem[968][3] ), .B(\mem[969][3] ), .S(n8390), .Z(n3117)
         );
  MUX2_X1 U22070 ( .A(n3117), .B(n3116), .S(n8310), .Z(n3118) );
  MUX2_X1 U22071 ( .A(n3118), .B(n3115), .S(n8259), .Z(n3119) );
  MUX2_X1 U22072 ( .A(\mem[966][3] ), .B(\mem[967][3] ), .S(n8445), .Z(n3120)
         );
  MUX2_X1 U22073 ( .A(\mem[964][3] ), .B(\mem[965][3] ), .S(n8405), .Z(n3121)
         );
  MUX2_X1 U22074 ( .A(n3121), .B(n3120), .S(n8282), .Z(n3122) );
  MUX2_X1 U22075 ( .A(\mem[962][3] ), .B(\mem[963][3] ), .S(n8386), .Z(n3123)
         );
  MUX2_X1 U22076 ( .A(\mem[960][3] ), .B(\mem[961][3] ), .S(n8537), .Z(n3124)
         );
  MUX2_X1 U22077 ( .A(n3124), .B(n3123), .S(n8328), .Z(n3125) );
  MUX2_X1 U22078 ( .A(n3125), .B(n3122), .S(n8259), .Z(n3126) );
  MUX2_X1 U22079 ( .A(n3126), .B(n3119), .S(n8203), .Z(n3127) );
  MUX2_X1 U22080 ( .A(n3127), .B(n3112), .S(n8194), .Z(n3128) );
  MUX2_X1 U22081 ( .A(n3128), .B(n3097), .S(n8184), .Z(n3129) );
  MUX2_X1 U22082 ( .A(\mem[958][3] ), .B(\mem[959][3] ), .S(n8406), .Z(n3130)
         );
  MUX2_X1 U22083 ( .A(\mem[956][3] ), .B(\mem[957][3] ), .S(n8404), .Z(n3131)
         );
  MUX2_X1 U22084 ( .A(n3131), .B(n3130), .S(n8278), .Z(n3132) );
  MUX2_X1 U22085 ( .A(\mem[954][3] ), .B(\mem[955][3] ), .S(n8405), .Z(n3133)
         );
  MUX2_X1 U22086 ( .A(\mem[952][3] ), .B(\mem[953][3] ), .S(n8365), .Z(n3134)
         );
  MUX2_X1 U22087 ( .A(n3134), .B(n3133), .S(n8275), .Z(n3135) );
  MUX2_X1 U22088 ( .A(n3135), .B(n3132), .S(n8259), .Z(n3136) );
  MUX2_X1 U22089 ( .A(\mem[950][3] ), .B(\mem[951][3] ), .S(n8388), .Z(n3137)
         );
  MUX2_X1 U22090 ( .A(\mem[948][3] ), .B(\mem[949][3] ), .S(n8389), .Z(n3138)
         );
  MUX2_X1 U22091 ( .A(n3138), .B(n3137), .S(n8274), .Z(n3139) );
  MUX2_X1 U22092 ( .A(\mem[946][3] ), .B(\mem[947][3] ), .S(n8438), .Z(n3140)
         );
  MUX2_X1 U22093 ( .A(\mem[944][3] ), .B(\mem[945][3] ), .S(n8381), .Z(n3141)
         );
  MUX2_X1 U22094 ( .A(n3141), .B(n3140), .S(n8273), .Z(n3142) );
  MUX2_X1 U22095 ( .A(n3142), .B(n3139), .S(n8259), .Z(n3143) );
  MUX2_X1 U22096 ( .A(n3143), .B(n3136), .S(n8206), .Z(n3144) );
  MUX2_X1 U22097 ( .A(\mem[942][3] ), .B(\mem[943][3] ), .S(n8535), .Z(n3145)
         );
  MUX2_X1 U22098 ( .A(\mem[940][3] ), .B(\mem[941][3] ), .S(n8536), .Z(n3146)
         );
  MUX2_X1 U22099 ( .A(n3146), .B(n3145), .S(n8329), .Z(n3147) );
  MUX2_X1 U22100 ( .A(\mem[938][3] ), .B(\mem[939][3] ), .S(n8531), .Z(n3148)
         );
  MUX2_X1 U22101 ( .A(\mem[936][3] ), .B(\mem[937][3] ), .S(n8532), .Z(n3149)
         );
  MUX2_X1 U22102 ( .A(n3149), .B(n3148), .S(n8330), .Z(n3150) );
  MUX2_X1 U22103 ( .A(n3150), .B(n3147), .S(n8259), .Z(n3151) );
  MUX2_X1 U22104 ( .A(\mem[934][3] ), .B(\mem[935][3] ), .S(n8533), .Z(n3152)
         );
  MUX2_X1 U22105 ( .A(\mem[932][3] ), .B(\mem[933][3] ), .S(n8398), .Z(n3153)
         );
  MUX2_X1 U22106 ( .A(n3153), .B(n3152), .S(n8331), .Z(n3154) );
  MUX2_X1 U22107 ( .A(\mem[930][3] ), .B(\mem[931][3] ), .S(n8399), .Z(n3155)
         );
  MUX2_X1 U22108 ( .A(\mem[928][3] ), .B(\mem[929][3] ), .S(n8400), .Z(n3156)
         );
  MUX2_X1 U22109 ( .A(n3156), .B(n3155), .S(n8338), .Z(n3157) );
  MUX2_X1 U22110 ( .A(n3157), .B(n3154), .S(n8259), .Z(n3158) );
  MUX2_X1 U22111 ( .A(n3158), .B(n3151), .S(n8202), .Z(n3159) );
  MUX2_X1 U22112 ( .A(n3159), .B(n3144), .S(n8189), .Z(n3160) );
  MUX2_X1 U22113 ( .A(\mem[926][3] ), .B(\mem[927][3] ), .S(n8395), .Z(n3161)
         );
  MUX2_X1 U22114 ( .A(\mem[924][3] ), .B(\mem[925][3] ), .S(n8396), .Z(n3162)
         );
  MUX2_X1 U22115 ( .A(n3162), .B(n3161), .S(n8339), .Z(n3163) );
  MUX2_X1 U22116 ( .A(\mem[922][3] ), .B(\mem[923][3] ), .S(n8397), .Z(n3164)
         );
  MUX2_X1 U22117 ( .A(\mem[920][3] ), .B(\mem[921][3] ), .S(n8404), .Z(n3165)
         );
  MUX2_X1 U22118 ( .A(n3165), .B(n3164), .S(n8340), .Z(n3166) );
  MUX2_X1 U22119 ( .A(n3166), .B(n3163), .S(n8259), .Z(n3167) );
  MUX2_X1 U22120 ( .A(\mem[918][3] ), .B(\mem[919][3] ), .S(n8357), .Z(n3168)
         );
  MUX2_X1 U22121 ( .A(\mem[916][3] ), .B(\mem[917][3] ), .S(n8389), .Z(n3169)
         );
  MUX2_X1 U22122 ( .A(n3169), .B(n3168), .S(n8335), .Z(n3170) );
  MUX2_X1 U22123 ( .A(\mem[914][3] ), .B(\mem[915][3] ), .S(n8537), .Z(n3171)
         );
  MUX2_X1 U22124 ( .A(\mem[912][3] ), .B(\mem[913][3] ), .S(n8388), .Z(n3172)
         );
  MUX2_X1 U22125 ( .A(n3172), .B(n3171), .S(n8336), .Z(n3173) );
  MUX2_X1 U22126 ( .A(n3173), .B(n3170), .S(n8259), .Z(n3174) );
  MUX2_X1 U22127 ( .A(n3174), .B(n3167), .S(n8203), .Z(n3175) );
  MUX2_X1 U22128 ( .A(\mem[910][3] ), .B(\mem[911][3] ), .S(n8386), .Z(n3176)
         );
  MUX2_X1 U22129 ( .A(\mem[908][3] ), .B(\mem[909][3] ), .S(n8365), .Z(n3177)
         );
  MUX2_X1 U22130 ( .A(n3177), .B(n3176), .S(n8337), .Z(n3178) );
  MUX2_X1 U22131 ( .A(\mem[906][3] ), .B(\mem[907][3] ), .S(n8387), .Z(n3179)
         );
  MUX2_X1 U22132 ( .A(\mem[904][3] ), .B(\mem[905][3] ), .S(n8357), .Z(n3180)
         );
  MUX2_X1 U22133 ( .A(n3180), .B(n3179), .S(n8344), .Z(n3181) );
  MUX2_X1 U22134 ( .A(n3181), .B(n3178), .S(n8259), .Z(n3182) );
  MUX2_X1 U22135 ( .A(\mem[902][3] ), .B(\mem[903][3] ), .S(n8389), .Z(n3183)
         );
  MUX2_X1 U22136 ( .A(\mem[900][3] ), .B(\mem[901][3] ), .S(n8537), .Z(n3184)
         );
  MUX2_X1 U22137 ( .A(n3184), .B(n3183), .S(n8345), .Z(n3185) );
  MUX2_X1 U22138 ( .A(\mem[898][3] ), .B(\mem[899][3] ), .S(n8388), .Z(n3186)
         );
  MUX2_X1 U22139 ( .A(\mem[896][3] ), .B(\mem[897][3] ), .S(n8386), .Z(n3187)
         );
  MUX2_X1 U22140 ( .A(n3187), .B(n3186), .S(n8346), .Z(n3188) );
  MUX2_X1 U22141 ( .A(n3188), .B(n3185), .S(n8259), .Z(n3189) );
  MUX2_X1 U22142 ( .A(n3189), .B(n3182), .S(n8204), .Z(n3190) );
  MUX2_X1 U22143 ( .A(n3190), .B(n3175), .S(n8195), .Z(n3191) );
  MUX2_X1 U22144 ( .A(n3191), .B(n3160), .S(n8184), .Z(n3192) );
  MUX2_X1 U22145 ( .A(n3192), .B(n3129), .S(n8180), .Z(n3193) );
  MUX2_X1 U22146 ( .A(\mem[894][3] ), .B(\mem[895][3] ), .S(n8387), .Z(n3194)
         );
  MUX2_X1 U22147 ( .A(\mem[892][3] ), .B(\mem[893][3] ), .S(n8537), .Z(n3195)
         );
  MUX2_X1 U22148 ( .A(n3195), .B(n3194), .S(n8303), .Z(n3196) );
  MUX2_X1 U22149 ( .A(\mem[890][3] ), .B(\mem[891][3] ), .S(n8357), .Z(n3197)
         );
  MUX2_X1 U22150 ( .A(\mem[888][3] ), .B(\mem[889][3] ), .S(n8389), .Z(n3198)
         );
  MUX2_X1 U22151 ( .A(n3198), .B(n3197), .S(n8304), .Z(n3199) );
  MUX2_X1 U22152 ( .A(n3199), .B(n3196), .S(n8260), .Z(n3200) );
  MUX2_X1 U22153 ( .A(\mem[886][3] ), .B(\mem[887][3] ), .S(n8388), .Z(n3201)
         );
  MUX2_X1 U22154 ( .A(\mem[884][3] ), .B(\mem[885][3] ), .S(n8537), .Z(n3202)
         );
  MUX2_X1 U22155 ( .A(n3202), .B(n3201), .S(n8299), .Z(n3203) );
  MUX2_X1 U22156 ( .A(\mem[882][3] ), .B(\mem[883][3] ), .S(n8386), .Z(n3204)
         );
  MUX2_X1 U22157 ( .A(\mem[880][3] ), .B(\mem[881][3] ), .S(n8365), .Z(n3205)
         );
  MUX2_X1 U22158 ( .A(n3205), .B(n3204), .S(n8300), .Z(n3206) );
  MUX2_X1 U22159 ( .A(n3206), .B(n3203), .S(n8260), .Z(n3207) );
  MUX2_X1 U22160 ( .A(n3207), .B(n3200), .S(n8208), .Z(n3208) );
  MUX2_X1 U22161 ( .A(\mem[878][3] ), .B(\mem[879][3] ), .S(n8387), .Z(n3209)
         );
  MUX2_X1 U22162 ( .A(\mem[876][3] ), .B(\mem[877][3] ), .S(n8357), .Z(n3210)
         );
  MUX2_X1 U22163 ( .A(n3210), .B(n3209), .S(n8301), .Z(n3211) );
  MUX2_X1 U22164 ( .A(\mem[874][3] ), .B(\mem[875][3] ), .S(n8389), .Z(n3212)
         );
  MUX2_X1 U22165 ( .A(\mem[872][3] ), .B(\mem[873][3] ), .S(n8537), .Z(n3213)
         );
  MUX2_X1 U22166 ( .A(n3213), .B(n3212), .S(n8326), .Z(n3214) );
  MUX2_X1 U22167 ( .A(n3214), .B(n3211), .S(n8260), .Z(n3215) );
  MUX2_X1 U22168 ( .A(\mem[870][3] ), .B(\mem[871][3] ), .S(n8393), .Z(n3216)
         );
  MUX2_X1 U22169 ( .A(\mem[868][3] ), .B(\mem[869][3] ), .S(n8394), .Z(n3217)
         );
  MUX2_X1 U22170 ( .A(n3217), .B(n3216), .S(n8327), .Z(n3218) );
  MUX2_X1 U22171 ( .A(\mem[866][3] ), .B(\mem[867][3] ), .S(n8390), .Z(n3219)
         );
  MUX2_X1 U22172 ( .A(\mem[864][3] ), .B(\mem[865][3] ), .S(n8391), .Z(n3220)
         );
  MUX2_X1 U22173 ( .A(n3220), .B(n3219), .S(n8328), .Z(n3221) );
  MUX2_X1 U22174 ( .A(n3221), .B(n3218), .S(n8260), .Z(n3222) );
  MUX2_X1 U22175 ( .A(n3222), .B(n3215), .S(N21), .Z(n3223) );
  MUX2_X1 U22176 ( .A(n3223), .B(n3208), .S(n8186), .Z(n3224) );
  MUX2_X1 U22177 ( .A(\mem[862][3] ), .B(\mem[863][3] ), .S(n8392), .Z(n3225)
         );
  MUX2_X1 U22178 ( .A(\mem[860][3] ), .B(\mem[861][3] ), .S(n8389), .Z(n3226)
         );
  MUX2_X1 U22179 ( .A(n3226), .B(n3225), .S(n8323), .Z(n3227) );
  MUX2_X1 U22180 ( .A(\mem[858][3] ), .B(\mem[859][3] ), .S(n8397), .Z(n3228)
         );
  MUX2_X1 U22181 ( .A(\mem[856][3] ), .B(\mem[857][3] ), .S(n8537), .Z(n3229)
         );
  MUX2_X1 U22182 ( .A(n3229), .B(n3228), .S(n8324), .Z(n3230) );
  MUX2_X1 U22183 ( .A(n3230), .B(n3227), .S(n8260), .Z(n3231) );
  MUX2_X1 U22184 ( .A(\mem[854][3] ), .B(\mem[855][3] ), .S(n8388), .Z(n3232)
         );
  MUX2_X1 U22185 ( .A(\mem[852][3] ), .B(\mem[853][3] ), .S(n8386), .Z(n3233)
         );
  MUX2_X1 U22186 ( .A(n3233), .B(n3232), .S(n8325), .Z(n3234) );
  MUX2_X1 U22187 ( .A(\mem[850][3] ), .B(\mem[851][3] ), .S(n8365), .Z(n3235)
         );
  MUX2_X1 U22188 ( .A(\mem[848][3] ), .B(\mem[849][3] ), .S(n8387), .Z(n3236)
         );
  MUX2_X1 U22189 ( .A(n3236), .B(n3235), .S(n8332), .Z(n3237) );
  MUX2_X1 U22190 ( .A(n3237), .B(n3234), .S(n8260), .Z(n3238) );
  MUX2_X1 U22191 ( .A(n3238), .B(n3231), .S(n8198), .Z(n3239) );
  MUX2_X1 U22192 ( .A(\mem[846][3] ), .B(\mem[847][3] ), .S(n8536), .Z(n3240)
         );
  MUX2_X1 U22193 ( .A(\mem[844][3] ), .B(\mem[845][3] ), .S(n8531), .Z(n3241)
         );
  MUX2_X1 U22194 ( .A(n3241), .B(n3240), .S(n8305), .Z(n3242) );
  MUX2_X1 U22195 ( .A(\mem[842][3] ), .B(\mem[843][3] ), .S(n8532), .Z(n3243)
         );
  MUX2_X1 U22196 ( .A(\mem[840][3] ), .B(\mem[841][3] ), .S(n8533), .Z(n3244)
         );
  MUX2_X1 U22197 ( .A(n3244), .B(n3243), .S(n8311), .Z(n3245) );
  MUX2_X1 U22198 ( .A(n3245), .B(n3242), .S(n8260), .Z(n3246) );
  MUX2_X1 U22199 ( .A(\mem[838][3] ), .B(\mem[839][3] ), .S(n8398), .Z(n3247)
         );
  MUX2_X1 U22200 ( .A(\mem[836][3] ), .B(\mem[837][3] ), .S(n8399), .Z(n3248)
         );
  MUX2_X1 U22201 ( .A(n3248), .B(n3247), .S(n8312), .Z(n3249) );
  MUX2_X1 U22202 ( .A(\mem[834][3] ), .B(\mem[835][3] ), .S(n8400), .Z(n3250)
         );
  MUX2_X1 U22203 ( .A(\mem[832][3] ), .B(\mem[833][3] ), .S(n8395), .Z(n3251)
         );
  MUX2_X1 U22204 ( .A(n3251), .B(n3250), .S(n8313), .Z(n3252) );
  MUX2_X1 U22205 ( .A(n3252), .B(n3249), .S(n8260), .Z(n3253) );
  MUX2_X1 U22206 ( .A(n3253), .B(n3246), .S(n8200), .Z(n3254) );
  MUX2_X1 U22207 ( .A(n3254), .B(n3239), .S(n8196), .Z(n3255) );
  MUX2_X1 U22208 ( .A(n3255), .B(n3224), .S(n8184), .Z(n3256) );
  MUX2_X1 U22209 ( .A(\mem[830][3] ), .B(\mem[831][3] ), .S(n8396), .Z(n3257)
         );
  MUX2_X1 U22210 ( .A(\mem[828][3] ), .B(\mem[829][3] ), .S(n8397), .Z(n3258)
         );
  MUX2_X1 U22211 ( .A(n3258), .B(n3257), .S(n8320), .Z(n3259) );
  MUX2_X1 U22212 ( .A(\mem[826][3] ), .B(\mem[827][3] ), .S(n8404), .Z(n3260)
         );
  MUX2_X1 U22213 ( .A(\mem[824][3] ), .B(\mem[825][3] ), .S(n8405), .Z(n3261)
         );
  MUX2_X1 U22214 ( .A(n3261), .B(n3260), .S(n8321), .Z(n3262) );
  MUX2_X1 U22215 ( .A(n3262), .B(n3259), .S(n8260), .Z(n3263) );
  MUX2_X1 U22216 ( .A(\mem[822][3] ), .B(\mem[823][3] ), .S(n8403), .Z(n3264)
         );
  MUX2_X1 U22217 ( .A(\mem[820][3] ), .B(\mem[821][3] ), .S(n8393), .Z(n3265)
         );
  MUX2_X1 U22218 ( .A(n3265), .B(n3264), .S(n8322), .Z(n3266) );
  MUX2_X1 U22219 ( .A(\mem[818][3] ), .B(\mem[819][3] ), .S(n8394), .Z(n3267)
         );
  MUX2_X1 U22220 ( .A(\mem[816][3] ), .B(\mem[817][3] ), .S(n8390), .Z(n3268)
         );
  MUX2_X1 U22221 ( .A(n3268), .B(n3267), .S(n8317), .Z(n3269) );
  MUX2_X1 U22222 ( .A(n3269), .B(n3266), .S(n8260), .Z(n3270) );
  MUX2_X1 U22223 ( .A(n3270), .B(n3263), .S(n8199), .Z(n3271) );
  MUX2_X1 U22224 ( .A(\mem[814][3] ), .B(\mem[815][3] ), .S(n8391), .Z(n3272)
         );
  MUX2_X1 U22225 ( .A(\mem[812][3] ), .B(\mem[813][3] ), .S(n8392), .Z(n3273)
         );
  MUX2_X1 U22226 ( .A(n3273), .B(n3272), .S(n8318), .Z(n3274) );
  MUX2_X1 U22227 ( .A(\mem[810][3] ), .B(\mem[811][3] ), .S(n8389), .Z(n3275)
         );
  MUX2_X1 U22228 ( .A(\mem[808][3] ), .B(\mem[809][3] ), .S(n8537), .Z(n3276)
         );
  MUX2_X1 U22229 ( .A(n3276), .B(n3275), .S(n8319), .Z(n3277) );
  MUX2_X1 U22230 ( .A(n3277), .B(n3274), .S(n8260), .Z(n3278) );
  MUX2_X1 U22231 ( .A(\mem[806][3] ), .B(\mem[807][3] ), .S(n8388), .Z(n3279)
         );
  MUX2_X1 U22232 ( .A(\mem[804][3] ), .B(\mem[805][3] ), .S(n8386), .Z(n3280)
         );
  MUX2_X1 U22233 ( .A(n3280), .B(n3279), .S(n8326), .Z(n3281) );
  MUX2_X1 U22234 ( .A(\mem[802][3] ), .B(\mem[803][3] ), .S(n8365), .Z(n3282)
         );
  MUX2_X1 U22235 ( .A(\mem[800][3] ), .B(\mem[801][3] ), .S(n8387), .Z(n3283)
         );
  MUX2_X1 U22236 ( .A(n3283), .B(n3282), .S(n8327), .Z(n3284) );
  MUX2_X1 U22237 ( .A(n3284), .B(n3281), .S(n8260), .Z(n3285) );
  MUX2_X1 U22238 ( .A(n3285), .B(n3278), .S(n8200), .Z(n3286) );
  MUX2_X1 U22239 ( .A(n3286), .B(n3271), .S(n8195), .Z(n3287) );
  MUX2_X1 U22240 ( .A(\mem[798][3] ), .B(\mem[799][3] ), .S(n8517), .Z(n3288)
         );
  MUX2_X1 U22241 ( .A(\mem[796][3] ), .B(\mem[797][3] ), .S(n8518), .Z(n3289)
         );
  MUX2_X1 U22242 ( .A(n3289), .B(n3288), .S(n8282), .Z(n3290) );
  MUX2_X1 U22243 ( .A(\mem[794][3] ), .B(\mem[795][3] ), .S(n8513), .Z(n3291)
         );
  MUX2_X1 U22244 ( .A(\mem[792][3] ), .B(\mem[793][3] ), .S(n8514), .Z(n3292)
         );
  MUX2_X1 U22245 ( .A(n3292), .B(n3291), .S(n8304), .Z(n3293) );
  MUX2_X1 U22246 ( .A(n3293), .B(n3290), .S(n8261), .Z(n3294) );
  MUX2_X1 U22247 ( .A(\mem[790][3] ), .B(\mem[791][3] ), .S(n8515), .Z(n3295)
         );
  MUX2_X1 U22248 ( .A(\mem[788][3] ), .B(\mem[789][3] ), .S(n8522), .Z(n3296)
         );
  MUX2_X1 U22249 ( .A(n3296), .B(n3295), .S(n8292), .Z(n3297) );
  MUX2_X1 U22250 ( .A(\mem[786][3] ), .B(\mem[787][3] ), .S(n8523), .Z(n3298)
         );
  MUX2_X1 U22251 ( .A(\mem[784][3] ), .B(\mem[785][3] ), .S(n8524), .Z(n3299)
         );
  MUX2_X1 U22252 ( .A(n3299), .B(n3298), .S(n8281), .Z(n3300) );
  MUX2_X1 U22253 ( .A(n3300), .B(n3297), .S(n8261), .Z(n3301) );
  MUX2_X1 U22254 ( .A(n3301), .B(n3294), .S(n8199), .Z(n3302) );
  MUX2_X1 U22255 ( .A(\mem[782][3] ), .B(\mem[783][3] ), .S(n8519), .Z(n3303)
         );
  MUX2_X1 U22256 ( .A(\mem[780][3] ), .B(\mem[781][3] ), .S(n8520), .Z(n3304)
         );
  MUX2_X1 U22257 ( .A(n3304), .B(n3303), .S(n8280), .Z(n3305) );
  MUX2_X1 U22258 ( .A(\mem[778][3] ), .B(\mem[779][3] ), .S(n8521), .Z(n3306)
         );
  MUX2_X1 U22259 ( .A(\mem[776][3] ), .B(\mem[777][3] ), .S(n8528), .Z(n3307)
         );
  MUX2_X1 U22260 ( .A(n3307), .B(n3306), .S(n8279), .Z(n3308) );
  MUX2_X1 U22261 ( .A(n3308), .B(n3305), .S(n8261), .Z(n3309) );
  MUX2_X1 U22262 ( .A(\mem[774][3] ), .B(\mem[775][3] ), .S(n8496), .Z(n3310)
         );
  MUX2_X1 U22263 ( .A(\mem[772][3] ), .B(\mem[773][3] ), .S(n8497), .Z(n3311)
         );
  MUX2_X1 U22264 ( .A(n3311), .B(n3310), .S(n8275), .Z(n3312) );
  MUX2_X1 U22265 ( .A(\mem[770][3] ), .B(\mem[771][3] ), .S(n8504), .Z(n3313)
         );
  MUX2_X1 U22266 ( .A(\mem[768][3] ), .B(\mem[769][3] ), .S(n8505), .Z(n3314)
         );
  MUX2_X1 U22267 ( .A(n3314), .B(n3313), .S(n8274), .Z(n3315) );
  MUX2_X1 U22268 ( .A(n3315), .B(n3312), .S(n8261), .Z(n3316) );
  MUX2_X1 U22269 ( .A(n3316), .B(n3309), .S(n8219), .Z(n3317) );
  MUX2_X1 U22270 ( .A(n3317), .B(n3302), .S(n8186), .Z(n3318) );
  MUX2_X1 U22271 ( .A(n3318), .B(n3287), .S(n8184), .Z(n3319) );
  MUX2_X1 U22272 ( .A(n3319), .B(n3256), .S(n8178), .Z(n3320) );
  MUX2_X1 U22273 ( .A(n3320), .B(n3193), .S(n8177), .Z(n3321) );
  MUX2_X1 U22274 ( .A(\mem[766][3] ), .B(\mem[767][3] ), .S(n8506), .Z(n3322)
         );
  MUX2_X1 U22275 ( .A(\mem[764][3] ), .B(\mem[765][3] ), .S(n8501), .Z(n3323)
         );
  MUX2_X1 U22276 ( .A(n3323), .B(n3322), .S(n8273), .Z(n3324) );
  MUX2_X1 U22277 ( .A(\mem[762][3] ), .B(\mem[763][3] ), .S(n8502), .Z(n3325)
         );
  MUX2_X1 U22278 ( .A(\mem[760][3] ), .B(\mem[761][3] ), .S(n8503), .Z(n3326)
         );
  MUX2_X1 U22279 ( .A(n3326), .B(n3325), .S(n8272), .Z(n3327) );
  MUX2_X1 U22280 ( .A(n3327), .B(n3324), .S(n8261), .Z(n3328) );
  MUX2_X1 U22281 ( .A(\mem[758][3] ), .B(\mem[759][3] ), .S(n8510), .Z(n3329)
         );
  MUX2_X1 U22282 ( .A(\mem[756][3] ), .B(\mem[757][3] ), .S(n8511), .Z(n3330)
         );
  MUX2_X1 U22283 ( .A(n3330), .B(n3329), .S(n8271), .Z(n3331) );
  MUX2_X1 U22284 ( .A(\mem[754][3] ), .B(\mem[755][3] ), .S(n8512), .Z(n3332)
         );
  MUX2_X1 U22285 ( .A(\mem[752][3] ), .B(\mem[753][3] ), .S(n8507), .Z(n3333)
         );
  MUX2_X1 U22286 ( .A(n3333), .B(n3332), .S(n8278), .Z(n3334) );
  MUX2_X1 U22287 ( .A(n3334), .B(n3331), .S(n8261), .Z(n3335) );
  MUX2_X1 U22288 ( .A(n3335), .B(n3328), .S(n8197), .Z(n3336) );
  MUX2_X1 U22289 ( .A(\mem[750][3] ), .B(\mem[751][3] ), .S(n8487), .Z(n3337)
         );
  MUX2_X1 U22290 ( .A(\mem[748][3] ), .B(\mem[749][3] ), .S(n8488), .Z(n3338)
         );
  MUX2_X1 U22291 ( .A(n3338), .B(n3337), .S(n8318), .Z(n3339) );
  MUX2_X1 U22292 ( .A(\mem[746][3] ), .B(\mem[747][3] ), .S(n8483), .Z(n3340)
         );
  MUX2_X1 U22293 ( .A(\mem[744][3] ), .B(\mem[745][3] ), .S(n8484), .Z(n3341)
         );
  MUX2_X1 U22294 ( .A(n3341), .B(n3340), .S(n8319), .Z(n3342) );
  MUX2_X1 U22295 ( .A(n3342), .B(n3339), .S(n8261), .Z(n3343) );
  MUX2_X1 U22296 ( .A(\mem[742][3] ), .B(\mem[743][3] ), .S(n8485), .Z(n3344)
         );
  MUX2_X1 U22297 ( .A(\mem[740][3] ), .B(\mem[741][3] ), .S(n8492), .Z(n3345)
         );
  MUX2_X1 U22298 ( .A(n3345), .B(n3344), .S(n8346), .Z(n3346) );
  MUX2_X1 U22299 ( .A(\mem[738][3] ), .B(\mem[739][3] ), .S(n8493), .Z(n3347)
         );
  MUX2_X1 U22300 ( .A(\mem[736][3] ), .B(\mem[737][3] ), .S(n8494), .Z(n3348)
         );
  MUX2_X1 U22301 ( .A(n3348), .B(n3347), .S(n8305), .Z(n3349) );
  MUX2_X1 U22302 ( .A(n3349), .B(n3346), .S(n8261), .Z(n3350) );
  MUX2_X1 U22303 ( .A(n3350), .B(n3343), .S(n8204), .Z(n3351) );
  MUX2_X1 U22304 ( .A(n3351), .B(n3336), .S(n8189), .Z(n3352) );
  MUX2_X1 U22305 ( .A(\mem[734][3] ), .B(\mem[735][3] ), .S(n8489), .Z(n3353)
         );
  MUX2_X1 U22306 ( .A(\mem[732][3] ), .B(\mem[733][3] ), .S(n8490), .Z(n3354)
         );
  MUX2_X1 U22307 ( .A(n3354), .B(n3353), .S(N19), .Z(n3355) );
  MUX2_X1 U22308 ( .A(\mem[730][3] ), .B(\mem[731][3] ), .S(n8491), .Z(n3356)
         );
  MUX2_X1 U22309 ( .A(\mem[728][3] ), .B(\mem[729][3] ), .S(n8498), .Z(n3357)
         );
  MUX2_X1 U22310 ( .A(n3357), .B(n3356), .S(n8356), .Z(n3358) );
  MUX2_X1 U22311 ( .A(n3358), .B(n3355), .S(n8261), .Z(n3359) );
  MUX2_X1 U22312 ( .A(\mem[726][3] ), .B(\mem[727][3] ), .S(n8448), .Z(n3360)
         );
  MUX2_X1 U22313 ( .A(\mem[724][3] ), .B(\mem[725][3] ), .S(n8392), .Z(n3361)
         );
  MUX2_X1 U22314 ( .A(n3361), .B(n3360), .S(n8346), .Z(n3362) );
  MUX2_X1 U22315 ( .A(\mem[722][3] ), .B(\mem[723][3] ), .S(n8507), .Z(n3363)
         );
  MUX2_X1 U22316 ( .A(\mem[720][3] ), .B(\mem[721][3] ), .S(n8492), .Z(n3364)
         );
  MUX2_X1 U22317 ( .A(n3364), .B(n3363), .S(n8325), .Z(n3365) );
  MUX2_X1 U22318 ( .A(n3365), .B(n3362), .S(n8261), .Z(n3366) );
  MUX2_X1 U22319 ( .A(n3366), .B(n3359), .S(n8207), .Z(n3367) );
  MUX2_X1 U22320 ( .A(\mem[718][3] ), .B(\mem[719][3] ), .S(n8409), .Z(n3368)
         );
  MUX2_X1 U22321 ( .A(\mem[716][3] ), .B(\mem[717][3] ), .S(n8459), .Z(n3369)
         );
  MUX2_X1 U22322 ( .A(n3369), .B(n3368), .S(n8267), .Z(n3370) );
  MUX2_X1 U22323 ( .A(\mem[714][3] ), .B(\mem[715][3] ), .S(n8428), .Z(n3371)
         );
  MUX2_X1 U22324 ( .A(\mem[712][3] ), .B(\mem[713][3] ), .S(n8423), .Z(n3372)
         );
  MUX2_X1 U22325 ( .A(n3372), .B(n3371), .S(n8266), .Z(n3373) );
  MUX2_X1 U22326 ( .A(n3373), .B(n3370), .S(n8261), .Z(n3374) );
  MUX2_X1 U22327 ( .A(\mem[710][3] ), .B(\mem[711][3] ), .S(n8537), .Z(n3375)
         );
  MUX2_X1 U22328 ( .A(\mem[708][3] ), .B(\mem[709][3] ), .S(n8388), .Z(n3376)
         );
  MUX2_X1 U22329 ( .A(n3376), .B(n3375), .S(n8324), .Z(n3377) );
  MUX2_X1 U22330 ( .A(\mem[706][3] ), .B(\mem[707][3] ), .S(n8379), .Z(n3378)
         );
  MUX2_X1 U22331 ( .A(\mem[704][3] ), .B(\mem[705][3] ), .S(n8410), .Z(n3379)
         );
  MUX2_X1 U22332 ( .A(n3379), .B(n3378), .S(n8299), .Z(n3380) );
  MUX2_X1 U22333 ( .A(n3380), .B(n3377), .S(n8261), .Z(n3381) );
  MUX2_X1 U22334 ( .A(n3381), .B(n3374), .S(n8208), .Z(n3382) );
  MUX2_X1 U22335 ( .A(n3382), .B(n3367), .S(n8195), .Z(n3383) );
  MUX2_X1 U22336 ( .A(n3383), .B(n3352), .S(n8184), .Z(n3384) );
  MUX2_X1 U22337 ( .A(\mem[702][3] ), .B(\mem[703][3] ), .S(n8406), .Z(n3385)
         );
  MUX2_X1 U22338 ( .A(\mem[700][3] ), .B(\mem[701][3] ), .S(n8401), .Z(n3386)
         );
  MUX2_X1 U22339 ( .A(n3386), .B(n3385), .S(n8343), .Z(n3387) );
  MUX2_X1 U22340 ( .A(\mem[698][3] ), .B(\mem[699][3] ), .S(n8402), .Z(n3388)
         );
  MUX2_X1 U22341 ( .A(\mem[696][3] ), .B(\mem[697][3] ), .S(n8403), .Z(n3389)
         );
  MUX2_X1 U22342 ( .A(n3389), .B(n3388), .S(n8350), .Z(n3390) );
  MUX2_X1 U22343 ( .A(n3390), .B(n3387), .S(n8221), .Z(n3391) );
  MUX2_X1 U22344 ( .A(\mem[694][3] ), .B(\mem[695][3] ), .S(n8393), .Z(n3392)
         );
  MUX2_X1 U22345 ( .A(\mem[692][3] ), .B(\mem[693][3] ), .S(n8394), .Z(n3393)
         );
  MUX2_X1 U22346 ( .A(n3393), .B(n3392), .S(n8351), .Z(n3394) );
  MUX2_X1 U22347 ( .A(\mem[690][3] ), .B(\mem[691][3] ), .S(n8390), .Z(n3395)
         );
  MUX2_X1 U22348 ( .A(\mem[688][3] ), .B(\mem[689][3] ), .S(n8391), .Z(n3396)
         );
  MUX2_X1 U22349 ( .A(n3396), .B(n3395), .S(n8352), .Z(n3397) );
  MUX2_X1 U22350 ( .A(n3397), .B(n3394), .S(n8263), .Z(n3398) );
  MUX2_X1 U22351 ( .A(n3398), .B(n3391), .S(n8214), .Z(n3399) );
  MUX2_X1 U22352 ( .A(\mem[686][3] ), .B(\mem[687][3] ), .S(n8392), .Z(n3400)
         );
  MUX2_X1 U22353 ( .A(\mem[684][3] ), .B(\mem[685][3] ), .S(n8389), .Z(n3401)
         );
  MUX2_X1 U22354 ( .A(n3401), .B(n3400), .S(n8347), .Z(n3402) );
  MUX2_X1 U22355 ( .A(\mem[682][3] ), .B(\mem[683][3] ), .S(n8430), .Z(n3403)
         );
  MUX2_X1 U22356 ( .A(\mem[680][3] ), .B(\mem[681][3] ), .S(n8431), .Z(n3404)
         );
  MUX2_X1 U22357 ( .A(n3404), .B(n3403), .S(n8348), .Z(n3405) );
  MUX2_X1 U22358 ( .A(n3405), .B(n3402), .S(n8265), .Z(n3406) );
  MUX2_X1 U22359 ( .A(\mem[678][3] ), .B(\mem[679][3] ), .S(n8527), .Z(n3407)
         );
  MUX2_X1 U22360 ( .A(\mem[676][3] ), .B(\mem[677][3] ), .S(n8534), .Z(n3408)
         );
  MUX2_X1 U22361 ( .A(n3408), .B(n3407), .S(n8349), .Z(n3409) );
  MUX2_X1 U22362 ( .A(\mem[674][3] ), .B(\mem[675][3] ), .S(n8535), .Z(n3410)
         );
  MUX2_X1 U22363 ( .A(\mem[672][3] ), .B(\mem[673][3] ), .S(n8536), .Z(n3411)
         );
  MUX2_X1 U22364 ( .A(n3411), .B(n3410), .S(n8353), .Z(n3412) );
  MUX2_X1 U22365 ( .A(n3412), .B(n3409), .S(n8264), .Z(n3413) );
  MUX2_X1 U22366 ( .A(n3413), .B(n3406), .S(n8215), .Z(n3414) );
  MUX2_X1 U22367 ( .A(n3414), .B(n3399), .S(n8187), .Z(n3415) );
  MUX2_X1 U22368 ( .A(\mem[670][3] ), .B(\mem[671][3] ), .S(n8531), .Z(n3416)
         );
  MUX2_X1 U22369 ( .A(\mem[668][3] ), .B(\mem[669][3] ), .S(n8532), .Z(n3417)
         );
  MUX2_X1 U22370 ( .A(n3417), .B(n3416), .S(n8354), .Z(n3418) );
  MUX2_X1 U22371 ( .A(\mem[666][3] ), .B(\mem[667][3] ), .S(n8533), .Z(n3419)
         );
  MUX2_X1 U22372 ( .A(\mem[664][3] ), .B(\mem[665][3] ), .S(n8398), .Z(n3420)
         );
  MUX2_X1 U22373 ( .A(n3420), .B(n3419), .S(n8355), .Z(n3421) );
  MUX2_X1 U22374 ( .A(n3421), .B(n3418), .S(n8238), .Z(n3422) );
  MUX2_X1 U22375 ( .A(\mem[662][3] ), .B(\mem[663][3] ), .S(n8399), .Z(n3423)
         );
  MUX2_X1 U22376 ( .A(\mem[660][3] ), .B(\mem[661][3] ), .S(n8400), .Z(n3424)
         );
  MUX2_X1 U22377 ( .A(n3424), .B(n3423), .S(n8313), .Z(n3425) );
  MUX2_X1 U22378 ( .A(\mem[658][3] ), .B(\mem[659][3] ), .S(n8395), .Z(n3426)
         );
  MUX2_X1 U22379 ( .A(\mem[656][3] ), .B(\mem[657][3] ), .S(n8396), .Z(n3427)
         );
  MUX2_X1 U22380 ( .A(n3427), .B(n3426), .S(n8320), .Z(n3428) );
  MUX2_X1 U22381 ( .A(n3428), .B(n3425), .S(n8222), .Z(n3429) );
  MUX2_X1 U22382 ( .A(n3429), .B(n3422), .S(n8211), .Z(n3430) );
  MUX2_X1 U22383 ( .A(\mem[654][3] ), .B(\mem[655][3] ), .S(n8500), .Z(n3431)
         );
  MUX2_X1 U22384 ( .A(\mem[652][3] ), .B(\mem[653][3] ), .S(n8495), .Z(n3432)
         );
  MUX2_X1 U22385 ( .A(n3432), .B(n3431), .S(n8351), .Z(n3433) );
  MUX2_X1 U22386 ( .A(\mem[650][3] ), .B(\mem[651][3] ), .S(n8496), .Z(n3434)
         );
  MUX2_X1 U22387 ( .A(\mem[648][3] ), .B(\mem[649][3] ), .S(n8497), .Z(n3435)
         );
  MUX2_X1 U22388 ( .A(n3435), .B(n3434), .S(n8352), .Z(n3436) );
  MUX2_X1 U22389 ( .A(n3436), .B(n3433), .S(n8225), .Z(n3437) );
  MUX2_X1 U22390 ( .A(\mem[646][3] ), .B(\mem[647][3] ), .S(n8504), .Z(n3438)
         );
  MUX2_X1 U22391 ( .A(\mem[644][3] ), .B(\mem[645][3] ), .S(n8505), .Z(n3439)
         );
  MUX2_X1 U22392 ( .A(n3439), .B(n3438), .S(n8347), .Z(n3440) );
  MUX2_X1 U22393 ( .A(\mem[642][3] ), .B(\mem[643][3] ), .S(n8506), .Z(n3441)
         );
  MUX2_X1 U22394 ( .A(\mem[640][3] ), .B(\mem[641][3] ), .S(n8501), .Z(n3442)
         );
  MUX2_X1 U22395 ( .A(n3442), .B(n3441), .S(n8348), .Z(n3443) );
  MUX2_X1 U22396 ( .A(n3443), .B(n3440), .S(n8256), .Z(n3444) );
  MUX2_X1 U22397 ( .A(n3444), .B(n3437), .S(n8216), .Z(n3445) );
  MUX2_X1 U22398 ( .A(n3445), .B(n3430), .S(n8191), .Z(n3446) );
  MUX2_X1 U22399 ( .A(n3446), .B(n3415), .S(n8184), .Z(n3447) );
  MUX2_X1 U22400 ( .A(n3447), .B(n3384), .S(N24), .Z(n3448) );
  MUX2_X1 U22401 ( .A(\mem[638][3] ), .B(\mem[639][3] ), .S(n8502), .Z(n3449)
         );
  MUX2_X1 U22402 ( .A(\mem[636][3] ), .B(\mem[637][3] ), .S(n8503), .Z(n3450)
         );
  MUX2_X1 U22403 ( .A(n3450), .B(n3449), .S(n8349), .Z(n3451) );
  MUX2_X1 U22404 ( .A(\mem[634][3] ), .B(\mem[635][3] ), .S(n8510), .Z(n3452)
         );
  MUX2_X1 U22405 ( .A(\mem[632][3] ), .B(\mem[633][3] ), .S(n8511), .Z(n3453)
         );
  MUX2_X1 U22406 ( .A(n3453), .B(n3452), .S(n8353), .Z(n3454) );
  MUX2_X1 U22407 ( .A(n3454), .B(n3451), .S(n8254), .Z(n3455) );
  MUX2_X1 U22408 ( .A(\mem[630][3] ), .B(\mem[631][3] ), .S(n8478), .Z(n3456)
         );
  MUX2_X1 U22409 ( .A(\mem[628][3] ), .B(\mem[629][3] ), .S(n8479), .Z(n3457)
         );
  MUX2_X1 U22410 ( .A(n3457), .B(n3456), .S(n8354), .Z(n3458) );
  MUX2_X1 U22411 ( .A(\mem[626][3] ), .B(\mem[627][3] ), .S(n8486), .Z(n3459)
         );
  MUX2_X1 U22412 ( .A(\mem[624][3] ), .B(\mem[625][3] ), .S(n8487), .Z(n3460)
         );
  MUX2_X1 U22413 ( .A(n3460), .B(n3459), .S(n8355), .Z(n3461) );
  MUX2_X1 U22414 ( .A(n3461), .B(n3458), .S(n8260), .Z(n3462) );
  MUX2_X1 U22415 ( .A(n3462), .B(n3455), .S(n8217), .Z(n3463) );
  MUX2_X1 U22416 ( .A(\mem[622][3] ), .B(\mem[623][3] ), .S(n8488), .Z(n3464)
         );
  MUX2_X1 U22417 ( .A(\mem[620][3] ), .B(\mem[621][3] ), .S(n8483), .Z(n3465)
         );
  MUX2_X1 U22418 ( .A(n3465), .B(n3464), .S(N19), .Z(n3466) );
  MUX2_X1 U22419 ( .A(\mem[618][3] ), .B(\mem[619][3] ), .S(n8484), .Z(n3467)
         );
  MUX2_X1 U22420 ( .A(\mem[616][3] ), .B(\mem[617][3] ), .S(n8485), .Z(n3468)
         );
  MUX2_X1 U22421 ( .A(n3468), .B(n3467), .S(n8356), .Z(n3469) );
  MUX2_X1 U22422 ( .A(n3469), .B(n3466), .S(n8224), .Z(n3470) );
  MUX2_X1 U22423 ( .A(\mem[614][3] ), .B(\mem[615][3] ), .S(n8492), .Z(n3471)
         );
  MUX2_X1 U22424 ( .A(\mem[612][3] ), .B(\mem[613][3] ), .S(n8493), .Z(n3472)
         );
  MUX2_X1 U22425 ( .A(n3472), .B(n3471), .S(n8345), .Z(n3473) );
  MUX2_X1 U22426 ( .A(\mem[610][3] ), .B(\mem[611][3] ), .S(n8494), .Z(n3474)
         );
  MUX2_X1 U22427 ( .A(\mem[608][3] ), .B(\mem[609][3] ), .S(n8489), .Z(n3475)
         );
  MUX2_X1 U22428 ( .A(n3475), .B(n3474), .S(n8267), .Z(n3476) );
  MUX2_X1 U22429 ( .A(n3476), .B(n3473), .S(n8223), .Z(n3477) );
  MUX2_X1 U22430 ( .A(n3477), .B(n3470), .S(n8218), .Z(n3478) );
  MUX2_X1 U22431 ( .A(n3478), .B(n3463), .S(n8196), .Z(n3479) );
  MUX2_X1 U22432 ( .A(\mem[606][3] ), .B(\mem[607][3] ), .S(n8462), .Z(n3480)
         );
  MUX2_X1 U22433 ( .A(\mem[604][3] ), .B(\mem[605][3] ), .S(n8535), .Z(n3481)
         );
  MUX2_X1 U22434 ( .A(n3481), .B(n3480), .S(n8330), .Z(n3482) );
  MUX2_X1 U22435 ( .A(\mem[602][3] ), .B(\mem[603][3] ), .S(n8468), .Z(n3483)
         );
  MUX2_X1 U22436 ( .A(\mem[600][3] ), .B(\mem[601][3] ), .S(n8465), .Z(n3484)
         );
  MUX2_X1 U22437 ( .A(n3484), .B(n3483), .S(n8331), .Z(n3485) );
  MUX2_X1 U22438 ( .A(n3485), .B(n3482), .S(n8229), .Z(n3486) );
  MUX2_X1 U22439 ( .A(\mem[598][3] ), .B(\mem[599][3] ), .S(n8466), .Z(n3487)
         );
  MUX2_X1 U22440 ( .A(\mem[596][3] ), .B(\mem[597][3] ), .S(n8467), .Z(n3488)
         );
  MUX2_X1 U22441 ( .A(n3488), .B(n3487), .S(n8338), .Z(n3489) );
  MUX2_X1 U22442 ( .A(\mem[594][3] ), .B(\mem[595][3] ), .S(n8474), .Z(n3490)
         );
  MUX2_X1 U22443 ( .A(\mem[592][3] ), .B(\mem[593][3] ), .S(n8475), .Z(n3491)
         );
  MUX2_X1 U22444 ( .A(n3491), .B(n3490), .S(n8339), .Z(n3492) );
  MUX2_X1 U22445 ( .A(n3492), .B(n3489), .S(n8220), .Z(n3493) );
  MUX2_X1 U22446 ( .A(n3493), .B(n3486), .S(n8205), .Z(n3494) );
  MUX2_X1 U22447 ( .A(\mem[590][3] ), .B(\mem[591][3] ), .S(n8476), .Z(n3495)
         );
  MUX2_X1 U22448 ( .A(\mem[588][3] ), .B(\mem[589][3] ), .S(n8471), .Z(n3496)
         );
  MUX2_X1 U22449 ( .A(n3496), .B(n3495), .S(n8340), .Z(n3497) );
  MUX2_X1 U22450 ( .A(\mem[586][3] ), .B(\mem[587][3] ), .S(n8472), .Z(n3498)
         );
  MUX2_X1 U22451 ( .A(\mem[584][3] ), .B(\mem[585][3] ), .S(n8473), .Z(n3499)
         );
  MUX2_X1 U22452 ( .A(n3499), .B(n3498), .S(n8335), .Z(n3500) );
  MUX2_X1 U22453 ( .A(n3500), .B(n3497), .S(n8224), .Z(n3501) );
  MUX2_X1 U22454 ( .A(\mem[582][3] ), .B(\mem[583][3] ), .S(N18), .Z(n3502) );
  MUX2_X1 U22455 ( .A(\mem[580][3] ), .B(\mem[581][3] ), .S(n8461), .Z(n3503)
         );
  MUX2_X1 U22456 ( .A(n3503), .B(n3502), .S(n8336), .Z(n3504) );
  MUX2_X1 U22457 ( .A(\mem[578][3] ), .B(\mem[579][3] ), .S(n8443), .Z(n3505)
         );
  MUX2_X1 U22458 ( .A(\mem[576][3] ), .B(\mem[577][3] ), .S(n8519), .Z(n3506)
         );
  MUX2_X1 U22459 ( .A(n3506), .B(n3505), .S(n8337), .Z(n3507) );
  MUX2_X1 U22460 ( .A(n3507), .B(n3504), .S(n8223), .Z(n3508) );
  MUX2_X1 U22461 ( .A(n3508), .B(n3501), .S(n8209), .Z(n3509) );
  MUX2_X1 U22462 ( .A(n3509), .B(n3494), .S(N22), .Z(n3510) );
  MUX2_X1 U22463 ( .A(n3510), .B(n3479), .S(n8184), .Z(n3511) );
  MUX2_X1 U22464 ( .A(\mem[574][3] ), .B(\mem[575][3] ), .S(n8505), .Z(n3512)
         );
  MUX2_X1 U22465 ( .A(\mem[572][3] ), .B(\mem[573][3] ), .S(n8486), .Z(n3513)
         );
  MUX2_X1 U22466 ( .A(n3513), .B(n3512), .S(n8344), .Z(n3514) );
  MUX2_X1 U22467 ( .A(\mem[570][3] ), .B(\mem[571][3] ), .S(n8383), .Z(n3515)
         );
  MUX2_X1 U22468 ( .A(\mem[568][3] ), .B(\mem[569][3] ), .S(n8380), .Z(n3516)
         );
  MUX2_X1 U22469 ( .A(n3516), .B(n3515), .S(n8345), .Z(n3517) );
  MUX2_X1 U22470 ( .A(n3517), .B(n3514), .S(n8225), .Z(n3518) );
  MUX2_X1 U22471 ( .A(\mem[566][3] ), .B(\mem[567][3] ), .S(n8402), .Z(n3519)
         );
  MUX2_X1 U22472 ( .A(\mem[564][3] ), .B(\mem[565][3] ), .S(n8503), .Z(n3520)
         );
  MUX2_X1 U22473 ( .A(n3520), .B(n3519), .S(n8346), .Z(n3521) );
  MUX2_X1 U22474 ( .A(\mem[562][3] ), .B(\mem[563][3] ), .S(n8484), .Z(n3522)
         );
  MUX2_X1 U22475 ( .A(\mem[560][3] ), .B(\mem[561][3] ), .S(n8486), .Z(n3523)
         );
  MUX2_X1 U22476 ( .A(n3523), .B(n3522), .S(n8341), .Z(n3524) );
  MUX2_X1 U22477 ( .A(n3524), .B(n3521), .S(n8265), .Z(n3525) );
  MUX2_X1 U22478 ( .A(n3525), .B(n3518), .S(n8201), .Z(n3526) );
  MUX2_X1 U22479 ( .A(\mem[558][3] ), .B(\mem[559][3] ), .S(n8525), .Z(n3527)
         );
  MUX2_X1 U22480 ( .A(\mem[556][3] ), .B(\mem[557][3] ), .S(n8526), .Z(n3528)
         );
  MUX2_X1 U22481 ( .A(n3528), .B(n3527), .S(n8321), .Z(n3529) );
  MUX2_X1 U22482 ( .A(\mem[554][3] ), .B(\mem[555][3] ), .S(n8527), .Z(n3530)
         );
  MUX2_X1 U22483 ( .A(\mem[552][3] ), .B(\mem[553][3] ), .S(n8534), .Z(n3531)
         );
  MUX2_X1 U22484 ( .A(n3531), .B(n3530), .S(n8322), .Z(n3532) );
  MUX2_X1 U22485 ( .A(n3532), .B(n3529), .S(n8231), .Z(n3533) );
  MUX2_X1 U22486 ( .A(\mem[550][3] ), .B(\mem[551][3] ), .S(n8535), .Z(n3534)
         );
  MUX2_X1 U22487 ( .A(\mem[548][3] ), .B(\mem[549][3] ), .S(n8536), .Z(n3535)
         );
  MUX2_X1 U22488 ( .A(n3535), .B(n3534), .S(n8317), .Z(n3536) );
  MUX2_X1 U22489 ( .A(\mem[546][3] ), .B(\mem[547][3] ), .S(n8531), .Z(n3537)
         );
  MUX2_X1 U22490 ( .A(\mem[544][3] ), .B(\mem[545][3] ), .S(n8532), .Z(n3538)
         );
  MUX2_X1 U22491 ( .A(n3538), .B(n3537), .S(n8318), .Z(n3539) );
  MUX2_X1 U22492 ( .A(n3539), .B(n3536), .S(n8222), .Z(n3540) );
  MUX2_X1 U22493 ( .A(n3540), .B(n3533), .S(n8205), .Z(n3541) );
  MUX2_X1 U22494 ( .A(n3541), .B(n3526), .S(N22), .Z(n3542) );
  MUX2_X1 U22495 ( .A(\mem[542][3] ), .B(\mem[543][3] ), .S(n8533), .Z(n3543)
         );
  MUX2_X1 U22496 ( .A(\mem[540][3] ), .B(\mem[541][3] ), .S(n8398), .Z(n3544)
         );
  MUX2_X1 U22497 ( .A(n3544), .B(n3543), .S(n8319), .Z(n3545) );
  MUX2_X1 U22498 ( .A(\mem[538][3] ), .B(\mem[539][3] ), .S(n8399), .Z(n3546)
         );
  MUX2_X1 U22499 ( .A(\mem[536][3] ), .B(\mem[537][3] ), .S(n8400), .Z(n3547)
         );
  MUX2_X1 U22500 ( .A(n3547), .B(n3546), .S(n8326), .Z(n3548) );
  MUX2_X1 U22501 ( .A(n3548), .B(n3545), .S(n8221), .Z(n3549) );
  MUX2_X1 U22502 ( .A(\mem[534][3] ), .B(\mem[535][3] ), .S(n8516), .Z(n3550)
         );
  MUX2_X1 U22503 ( .A(\mem[532][3] ), .B(\mem[533][3] ), .S(n8517), .Z(n3551)
         );
  MUX2_X1 U22504 ( .A(n3551), .B(n3550), .S(n8327), .Z(n3552) );
  MUX2_X1 U22505 ( .A(\mem[530][3] ), .B(\mem[531][3] ), .S(n8518), .Z(n3553)
         );
  MUX2_X1 U22506 ( .A(\mem[528][3] ), .B(\mem[529][3] ), .S(n8513), .Z(n3554)
         );
  MUX2_X1 U22507 ( .A(n3554), .B(n3553), .S(n8328), .Z(n3555) );
  MUX2_X1 U22508 ( .A(n3555), .B(n3552), .S(n8255), .Z(n3556) );
  MUX2_X1 U22509 ( .A(n3556), .B(n3549), .S(n8216), .Z(n3557) );
  MUX2_X1 U22510 ( .A(\mem[526][3] ), .B(\mem[527][3] ), .S(n8514), .Z(n3558)
         );
  MUX2_X1 U22511 ( .A(\mem[524][3] ), .B(\mem[525][3] ), .S(n8515), .Z(n3559)
         );
  MUX2_X1 U22512 ( .A(n3559), .B(n3558), .S(n8323), .Z(n3560) );
  MUX2_X1 U22513 ( .A(\mem[522][3] ), .B(\mem[523][3] ), .S(n8522), .Z(n3561)
         );
  MUX2_X1 U22514 ( .A(\mem[520][3] ), .B(\mem[521][3] ), .S(n8523), .Z(n3562)
         );
  MUX2_X1 U22515 ( .A(n3562), .B(n3561), .S(n8324), .Z(n3563) );
  MUX2_X1 U22516 ( .A(n3563), .B(n3560), .S(n8226), .Z(n3564) );
  MUX2_X1 U22517 ( .A(\mem[518][3] ), .B(\mem[519][3] ), .S(n8524), .Z(n3565)
         );
  MUX2_X1 U22518 ( .A(\mem[516][3] ), .B(\mem[517][3] ), .S(n8519), .Z(n3566)
         );
  MUX2_X1 U22519 ( .A(n3566), .B(n3565), .S(n8325), .Z(n3567) );
  MUX2_X1 U22520 ( .A(\mem[514][3] ), .B(\mem[515][3] ), .S(n8520), .Z(n3568)
         );
  MUX2_X1 U22521 ( .A(\mem[512][3] ), .B(\mem[513][3] ), .S(n8521), .Z(n3569)
         );
  MUX2_X1 U22522 ( .A(n3569), .B(n3568), .S(n8332), .Z(n3570) );
  MUX2_X1 U22523 ( .A(n3570), .B(n3567), .S(n8220), .Z(n3571) );
  MUX2_X1 U22524 ( .A(n3571), .B(n3564), .S(n8202), .Z(n3572) );
  MUX2_X1 U22525 ( .A(n3572), .B(n3557), .S(n8191), .Z(n3573) );
  MUX2_X1 U22526 ( .A(n3573), .B(n3542), .S(n8184), .Z(n3574) );
  MUX2_X1 U22527 ( .A(n3574), .B(n3511), .S(n8179), .Z(n3575) );
  MUX2_X1 U22528 ( .A(n3575), .B(n3448), .S(n8177), .Z(n3576) );
  MUX2_X1 U22529 ( .A(n3576), .B(n3321), .S(N26), .Z(n3577) );
  MUX2_X1 U22530 ( .A(\mem[510][3] ), .B(\mem[511][3] ), .S(n8379), .Z(n3578)
         );
  MUX2_X1 U22531 ( .A(\mem[508][3] ), .B(\mem[509][3] ), .S(n8454), .Z(n3579)
         );
  MUX2_X1 U22532 ( .A(n3579), .B(n3578), .S(n8291), .Z(n3580) );
  MUX2_X1 U22533 ( .A(\mem[506][3] ), .B(\mem[507][3] ), .S(n8531), .Z(n3581)
         );
  MUX2_X1 U22534 ( .A(\mem[504][3] ), .B(\mem[505][3] ), .S(n8375), .Z(n3582)
         );
  MUX2_X1 U22535 ( .A(n3582), .B(n3581), .S(n8287), .Z(n3583) );
  MUX2_X1 U22536 ( .A(n3583), .B(n3580), .S(n8250), .Z(n3584) );
  MUX2_X1 U22537 ( .A(\mem[502][3] ), .B(\mem[503][3] ), .S(n8374), .Z(n3585)
         );
  MUX2_X1 U22538 ( .A(\mem[500][3] ), .B(\mem[501][3] ), .S(n8373), .Z(n3586)
         );
  MUX2_X1 U22539 ( .A(n3586), .B(n3585), .S(n8288), .Z(n3587) );
  MUX2_X1 U22540 ( .A(\mem[498][3] ), .B(\mem[499][3] ), .S(n8369), .Z(n3588)
         );
  MUX2_X1 U22541 ( .A(\mem[496][3] ), .B(\mem[497][3] ), .S(n8368), .Z(n3589)
         );
  MUX2_X1 U22542 ( .A(n3589), .B(n3588), .S(n8289), .Z(n3590) );
  MUX2_X1 U22543 ( .A(n3590), .B(n3587), .S(n8226), .Z(n3591) );
  MUX2_X1 U22544 ( .A(n3591), .B(n3584), .S(N21), .Z(n3592) );
  MUX2_X1 U22545 ( .A(\mem[494][3] ), .B(\mem[495][3] ), .S(n8387), .Z(n3593)
         );
  MUX2_X1 U22546 ( .A(\mem[492][3] ), .B(\mem[493][3] ), .S(n8386), .Z(n3594)
         );
  MUX2_X1 U22547 ( .A(n3594), .B(n3593), .S(n8296), .Z(n3595) );
  MUX2_X1 U22548 ( .A(\mem[490][3] ), .B(\mem[491][3] ), .S(n8383), .Z(n3596)
         );
  MUX2_X1 U22549 ( .A(\mem[488][3] ), .B(\mem[489][3] ), .S(n8411), .Z(n3597)
         );
  MUX2_X1 U22550 ( .A(n3597), .B(n3596), .S(n8297), .Z(n3598) );
  MUX2_X1 U22551 ( .A(n3598), .B(n3595), .S(n8222), .Z(n3599) );
  MUX2_X1 U22552 ( .A(\mem[486][3] ), .B(\mem[487][3] ), .S(n8435), .Z(n3600)
         );
  MUX2_X1 U22553 ( .A(\mem[484][3] ), .B(\mem[485][3] ), .S(n8527), .Z(n3601)
         );
  MUX2_X1 U22554 ( .A(n3601), .B(n3600), .S(n8298), .Z(n3602) );
  MUX2_X1 U22555 ( .A(\mem[482][3] ), .B(\mem[483][3] ), .S(n8538), .Z(n3603)
         );
  MUX2_X1 U22556 ( .A(\mem[480][3] ), .B(\mem[481][3] ), .S(n8372), .Z(n3604)
         );
  MUX2_X1 U22557 ( .A(n3604), .B(n3603), .S(n8293), .Z(n3605) );
  MUX2_X1 U22558 ( .A(n3605), .B(n3602), .S(n8220), .Z(n3606) );
  MUX2_X1 U22559 ( .A(n3606), .B(n3599), .S(n8199), .Z(n3607) );
  MUX2_X1 U22560 ( .A(n3607), .B(n3592), .S(n8186), .Z(n3608) );
  MUX2_X1 U22561 ( .A(\mem[478][3] ), .B(\mem[479][3] ), .S(n8396), .Z(n3609)
         );
  MUX2_X1 U22562 ( .A(\mem[476][3] ), .B(\mem[477][3] ), .S(n8390), .Z(n3610)
         );
  MUX2_X1 U22563 ( .A(n3610), .B(n3609), .S(n8294), .Z(n3611) );
  MUX2_X1 U22564 ( .A(\mem[474][3] ), .B(\mem[475][3] ), .S(n8511), .Z(n3612)
         );
  MUX2_X1 U22565 ( .A(\mem[472][3] ), .B(\mem[473][3] ), .S(n8484), .Z(n3613)
         );
  MUX2_X1 U22566 ( .A(n3613), .B(n3612), .S(n8295), .Z(n3614) );
  MUX2_X1 U22567 ( .A(n3614), .B(n3611), .S(n8263), .Z(n3615) );
  MUX2_X1 U22568 ( .A(\mem[470][3] ), .B(\mem[471][3] ), .S(n8409), .Z(n3616)
         );
  MUX2_X1 U22569 ( .A(\mem[468][3] ), .B(\mem[469][3] ), .S(n8463), .Z(n3617)
         );
  MUX2_X1 U22570 ( .A(n3617), .B(n3616), .S(n8302), .Z(n3618) );
  MUX2_X1 U22571 ( .A(\mem[466][3] ), .B(\mem[467][3] ), .S(n8410), .Z(n3619)
         );
  MUX2_X1 U22572 ( .A(\mem[464][3] ), .B(\mem[465][3] ), .S(n8407), .Z(n3620)
         );
  MUX2_X1 U22573 ( .A(n3620), .B(n3619), .S(n8303), .Z(n3621) );
  MUX2_X1 U22574 ( .A(n3621), .B(n3618), .S(n8265), .Z(n3622) );
  MUX2_X1 U22575 ( .A(n3622), .B(n3615), .S(n8198), .Z(n3623) );
  MUX2_X1 U22576 ( .A(\mem[462][3] ), .B(\mem[463][3] ), .S(n8360), .Z(n3624)
         );
  MUX2_X1 U22577 ( .A(\mem[460][3] ), .B(\mem[461][3] ), .S(n8377), .Z(n3625)
         );
  MUX2_X1 U22578 ( .A(n3625), .B(n3624), .S(n8272), .Z(n3626) );
  MUX2_X1 U22579 ( .A(\mem[458][3] ), .B(\mem[459][3] ), .S(n8479), .Z(n3627)
         );
  MUX2_X1 U22580 ( .A(\mem[456][3] ), .B(\mem[457][3] ), .S(n8460), .Z(n3628)
         );
  MUX2_X1 U22581 ( .A(n3628), .B(n3627), .S(n8271), .Z(n3629) );
  MUX2_X1 U22582 ( .A(n3629), .B(n3626), .S(n8264), .Z(n3630) );
  MUX2_X1 U22583 ( .A(\mem[454][3] ), .B(\mem[455][3] ), .S(n8442), .Z(n3631)
         );
  MUX2_X1 U22584 ( .A(\mem[452][3] ), .B(\mem[453][3] ), .S(n8524), .Z(n3632)
         );
  MUX2_X1 U22585 ( .A(n3632), .B(n3631), .S(n8345), .Z(n3633) );
  MUX2_X1 U22586 ( .A(\mem[450][3] ), .B(\mem[451][3] ), .S(n8504), .Z(n3634)
         );
  MUX2_X1 U22587 ( .A(\mem[448][3] ), .B(\mem[449][3] ), .S(n8515), .Z(n3635)
         );
  MUX2_X1 U22588 ( .A(n3635), .B(n3634), .S(n8282), .Z(n3636) );
  MUX2_X1 U22589 ( .A(n3636), .B(n3633), .S(n8239), .Z(n3637) );
  MUX2_X1 U22590 ( .A(n3637), .B(n3630), .S(n8200), .Z(n3638) );
  MUX2_X1 U22591 ( .A(n3638), .B(n3623), .S(n8186), .Z(n3639) );
  MUX2_X1 U22592 ( .A(n3639), .B(n3608), .S(n8181), .Z(n3640) );
  MUX2_X1 U22593 ( .A(\mem[446][3] ), .B(\mem[447][3] ), .S(n8384), .Z(n3641)
         );
  MUX2_X1 U22594 ( .A(\mem[444][3] ), .B(\mem[445][3] ), .S(n8388), .Z(n3642)
         );
  MUX2_X1 U22595 ( .A(n3642), .B(n3641), .S(n8308), .Z(n3643) );
  MUX2_X1 U22596 ( .A(\mem[442][3] ), .B(\mem[443][3] ), .S(n8401), .Z(n3644)
         );
  MUX2_X1 U22597 ( .A(\mem[440][3] ), .B(\mem[441][3] ), .S(n8502), .Z(n3645)
         );
  MUX2_X1 U22598 ( .A(n3645), .B(n3644), .S(n8266), .Z(n3646) );
  MUX2_X1 U22599 ( .A(n3646), .B(n3643), .S(n8221), .Z(n3647) );
  MUX2_X1 U22600 ( .A(\mem[438][3] ), .B(\mem[439][3] ), .S(n8452), .Z(n3648)
         );
  MUX2_X1 U22601 ( .A(\mem[436][3] ), .B(\mem[437][3] ), .S(n8447), .Z(n3649)
         );
  MUX2_X1 U22602 ( .A(n3649), .B(n3648), .S(n8268), .Z(n3650) );
  MUX2_X1 U22603 ( .A(\mem[434][3] ), .B(\mem[435][3] ), .S(n8448), .Z(n3651)
         );
  MUX2_X1 U22604 ( .A(\mem[432][3] ), .B(\mem[433][3] ), .S(n8449), .Z(n3652)
         );
  MUX2_X1 U22605 ( .A(n3652), .B(n3651), .S(n8269), .Z(n3653) );
  MUX2_X1 U22606 ( .A(n3653), .B(n3650), .S(n8225), .Z(n3654) );
  MUX2_X1 U22607 ( .A(n3654), .B(n3647), .S(n8217), .Z(n3655) );
  MUX2_X1 U22608 ( .A(\mem[430][3] ), .B(\mem[431][3] ), .S(n8456), .Z(n3656)
         );
  MUX2_X1 U22609 ( .A(\mem[428][3] ), .B(\mem[429][3] ), .S(n8457), .Z(n3657)
         );
  MUX2_X1 U22610 ( .A(n3657), .B(n3656), .S(n8270), .Z(n3658) );
  MUX2_X1 U22611 ( .A(\mem[426][3] ), .B(\mem[427][3] ), .S(n8458), .Z(n3659)
         );
  MUX2_X1 U22612 ( .A(\mem[424][3] ), .B(\mem[425][3] ), .S(n8453), .Z(n3660)
         );
  MUX2_X1 U22613 ( .A(n3660), .B(n3659), .S(n8326), .Z(n3661) );
  MUX2_X1 U22614 ( .A(n3661), .B(n3658), .S(n8265), .Z(n3662) );
  MUX2_X1 U22615 ( .A(\mem[422][3] ), .B(\mem[423][3] ), .S(n8454), .Z(n3663)
         );
  MUX2_X1 U22616 ( .A(\mem[420][3] ), .B(\mem[421][3] ), .S(n8455), .Z(n3664)
         );
  MUX2_X1 U22617 ( .A(n3664), .B(n3663), .S(n8328), .Z(n3665) );
  MUX2_X1 U22618 ( .A(\mem[418][3] ), .B(\mem[419][3] ), .S(n8462), .Z(n3666)
         );
  MUX2_X1 U22619 ( .A(\mem[416][3] ), .B(\mem[417][3] ), .S(n8463), .Z(n3667)
         );
  MUX2_X1 U22620 ( .A(n3667), .B(n3666), .S(n8290), .Z(n3668) );
  MUX2_X1 U22621 ( .A(n3668), .B(n3665), .S(n8223), .Z(n3669) );
  MUX2_X1 U22622 ( .A(n3669), .B(n3662), .S(N21), .Z(n3670) );
  MUX2_X1 U22623 ( .A(n3670), .B(n3655), .S(n8186), .Z(n3671) );
  MUX2_X1 U22624 ( .A(\mem[414][3] ), .B(\mem[415][3] ), .S(n8430), .Z(n3672)
         );
  MUX2_X1 U22625 ( .A(\mem[412][3] ), .B(\mem[413][3] ), .S(n8431), .Z(n3673)
         );
  MUX2_X1 U22626 ( .A(n3673), .B(n3672), .S(n8307), .Z(n3674) );
  MUX2_X1 U22627 ( .A(\mem[410][3] ), .B(\mem[411][3] ), .S(n8438), .Z(n3675)
         );
  MUX2_X1 U22628 ( .A(\mem[408][3] ), .B(\mem[409][3] ), .S(n8439), .Z(n3676)
         );
  MUX2_X1 U22629 ( .A(n3676), .B(n3675), .S(n8314), .Z(n3677) );
  MUX2_X1 U22630 ( .A(n3677), .B(n3674), .S(n8220), .Z(n3678) );
  MUX2_X1 U22631 ( .A(\mem[406][3] ), .B(\mem[407][3] ), .S(n8440), .Z(n3679)
         );
  MUX2_X1 U22632 ( .A(\mem[404][3] ), .B(\mem[405][3] ), .S(n8435), .Z(n3680)
         );
  MUX2_X1 U22633 ( .A(n3680), .B(n3679), .S(n8315), .Z(n3681) );
  MUX2_X1 U22634 ( .A(\mem[402][3] ), .B(\mem[403][3] ), .S(n8436), .Z(n3682)
         );
  MUX2_X1 U22635 ( .A(\mem[400][3] ), .B(\mem[401][3] ), .S(n8437), .Z(n3683)
         );
  MUX2_X1 U22636 ( .A(n3683), .B(n3682), .S(n8316), .Z(n3684) );
  MUX2_X1 U22637 ( .A(n3684), .B(n3681), .S(n8221), .Z(n3685) );
  MUX2_X1 U22638 ( .A(n3685), .B(n3678), .S(n8219), .Z(n3686) );
  MUX2_X1 U22639 ( .A(\mem[398][3] ), .B(\mem[399][3] ), .S(n8444), .Z(n3687)
         );
  MUX2_X1 U22640 ( .A(\mem[396][3] ), .B(\mem[397][3] ), .S(n8445), .Z(n3688)
         );
  MUX2_X1 U22641 ( .A(n3688), .B(n3687), .S(n8273), .Z(n3689) );
  MUX2_X1 U22642 ( .A(\mem[394][3] ), .B(\mem[395][3] ), .S(n8446), .Z(n3690)
         );
  MUX2_X1 U22643 ( .A(\mem[392][3] ), .B(\mem[393][3] ), .S(n8441), .Z(n3691)
         );
  MUX2_X1 U22644 ( .A(n3691), .B(n3690), .S(n8308), .Z(n3692) );
  MUX2_X1 U22645 ( .A(n3692), .B(n3689), .S(n8228), .Z(n3693) );
  MUX2_X1 U22646 ( .A(\mem[390][3] ), .B(\mem[391][3] ), .S(n8464), .Z(n3694)
         );
  MUX2_X1 U22647 ( .A(\mem[388][3] ), .B(\mem[389][3] ), .S(n8539), .Z(n3695)
         );
  MUX2_X1 U22648 ( .A(n3695), .B(n3694), .S(n8281), .Z(n3696) );
  MUX2_X1 U22649 ( .A(\mem[386][3] ), .B(\mem[387][3] ), .S(n8362), .Z(n3697)
         );
  MUX2_X1 U22650 ( .A(\mem[384][3] ), .B(\mem[385][3] ), .S(n8363), .Z(n3698)
         );
  MUX2_X1 U22651 ( .A(n3698), .B(n3697), .S(n8280), .Z(n3699) );
  MUX2_X1 U22652 ( .A(n3699), .B(n3696), .S(n8253), .Z(n3700) );
  MUX2_X1 U22653 ( .A(n3700), .B(n3693), .S(n8197), .Z(n3701) );
  MUX2_X1 U22654 ( .A(n3701), .B(n3686), .S(n8186), .Z(n3702) );
  MUX2_X1 U22655 ( .A(n3702), .B(n3671), .S(n8184), .Z(n3703) );
  MUX2_X1 U22656 ( .A(n3703), .B(n3640), .S(N24), .Z(n3704) );
  MUX2_X1 U22657 ( .A(\mem[382][3] ), .B(\mem[383][3] ), .S(n8364), .Z(n3705)
         );
  MUX2_X1 U22658 ( .A(\mem[380][3] ), .B(\mem[381][3] ), .S(n8357), .Z(n3706)
         );
  MUX2_X1 U22659 ( .A(n3706), .B(n3705), .S(n8279), .Z(n3707) );
  MUX2_X1 U22660 ( .A(\mem[378][3] ), .B(\mem[379][3] ), .S(n8424), .Z(n3708)
         );
  MUX2_X1 U22661 ( .A(\mem[376][3] ), .B(\mem[377][3] ), .S(n8358), .Z(n3709)
         );
  MUX2_X1 U22662 ( .A(n3709), .B(n3708), .S(n8278), .Z(n3710) );
  MUX2_X1 U22663 ( .A(n3710), .B(n3707), .S(n8220), .Z(n3711) );
  MUX2_X1 U22664 ( .A(\mem[374][3] ), .B(\mem[375][3] ), .S(n8443), .Z(n3712)
         );
  MUX2_X1 U22665 ( .A(\mem[372][3] ), .B(\mem[373][3] ), .S(n8360), .Z(n3713)
         );
  MUX2_X1 U22666 ( .A(n3713), .B(n3712), .S(n8277), .Z(n3714) );
  MUX2_X1 U22667 ( .A(\mem[370][3] ), .B(\mem[371][3] ), .S(n8395), .Z(n3715)
         );
  MUX2_X1 U22668 ( .A(\mem[368][3] ), .B(\mem[369][3] ), .S(n8432), .Z(n3716)
         );
  MUX2_X1 U22669 ( .A(n3716), .B(n3715), .S(n8276), .Z(n3717) );
  MUX2_X1 U22670 ( .A(n3717), .B(n3714), .S(n8226), .Z(n3718) );
  MUX2_X1 U22671 ( .A(n3718), .B(n3711), .S(n8215), .Z(n3719) );
  MUX2_X1 U22672 ( .A(\mem[366][3] ), .B(\mem[367][3] ), .S(n8426), .Z(n3720)
         );
  MUX2_X1 U22673 ( .A(\mem[364][3] ), .B(\mem[365][3] ), .S(n8427), .Z(n3721)
         );
  MUX2_X1 U22674 ( .A(n3721), .B(n3720), .S(n8267), .Z(n3722) );
  MUX2_X1 U22675 ( .A(\mem[362][3] ), .B(\mem[363][3] ), .S(n8428), .Z(n3723)
         );
  MUX2_X1 U22676 ( .A(\mem[360][3] ), .B(\mem[361][3] ), .S(n8374), .Z(n3724)
         );
  MUX2_X1 U22677 ( .A(n3724), .B(n3723), .S(n8306), .Z(n3725) );
  MUX2_X1 U22678 ( .A(n3725), .B(n3722), .S(n8224), .Z(n3726) );
  MUX2_X1 U22679 ( .A(\mem[358][3] ), .B(\mem[359][3] ), .S(n8370), .Z(n3727)
         );
  MUX2_X1 U22680 ( .A(\mem[356][3] ), .B(\mem[357][3] ), .S(n8537), .Z(n3728)
         );
  MUX2_X1 U22681 ( .A(n3728), .B(n3727), .S(n8344), .Z(n3729) );
  MUX2_X1 U22682 ( .A(\mem[354][3] ), .B(\mem[355][3] ), .S(n8424), .Z(n3730)
         );
  MUX2_X1 U22683 ( .A(\mem[352][3] ), .B(\mem[353][3] ), .S(n8425), .Z(n3731)
         );
  MUX2_X1 U22684 ( .A(n3731), .B(n3730), .S(n8278), .Z(n3732) );
  MUX2_X1 U22685 ( .A(n3732), .B(n3729), .S(n8225), .Z(n3733) );
  MUX2_X1 U22686 ( .A(n3733), .B(n3726), .S(n8207), .Z(n3734) );
  MUX2_X1 U22687 ( .A(n3734), .B(n3719), .S(n8186), .Z(n3735) );
  MUX2_X1 U22688 ( .A(\mem[350][3] ), .B(\mem[351][3] ), .S(n8396), .Z(n3736)
         );
  MUX2_X1 U22689 ( .A(\mem[348][3] ), .B(\mem[349][3] ), .S(n8397), .Z(n3737)
         );
  MUX2_X1 U22690 ( .A(n3737), .B(n3736), .S(n8344), .Z(n3738) );
  MUX2_X1 U22691 ( .A(\mem[346][3] ), .B(\mem[347][3] ), .S(n8404), .Z(n3739)
         );
  MUX2_X1 U22692 ( .A(\mem[344][3] ), .B(\mem[345][3] ), .S(n8405), .Z(n3740)
         );
  MUX2_X1 U22693 ( .A(n3740), .B(n3739), .S(n8301), .Z(n3741) );
  MUX2_X1 U22694 ( .A(n3741), .B(n3738), .S(n8263), .Z(n3742) );
  MUX2_X1 U22695 ( .A(\mem[342][3] ), .B(\mem[343][3] ), .S(n8407), .Z(n3743)
         );
  MUX2_X1 U22696 ( .A(\mem[340][3] ), .B(\mem[341][3] ), .S(n8408), .Z(n3744)
         );
  MUX2_X1 U22697 ( .A(n3744), .B(n3743), .S(n8282), .Z(n3745) );
  MUX2_X1 U22698 ( .A(\mem[338][3] ), .B(\mem[339][3] ), .S(n8470), .Z(n3746)
         );
  MUX2_X1 U22699 ( .A(\mem[336][3] ), .B(\mem[337][3] ), .S(n8414), .Z(n3747)
         );
  MUX2_X1 U22700 ( .A(n3747), .B(n3746), .S(n8281), .Z(n3748) );
  MUX2_X1 U22701 ( .A(n3748), .B(n3745), .S(n8265), .Z(n3749) );
  MUX2_X1 U22702 ( .A(n3749), .B(n3742), .S(n8208), .Z(n3750) );
  MUX2_X1 U22703 ( .A(\mem[334][3] ), .B(\mem[335][3] ), .S(n8415), .Z(n3751)
         );
  MUX2_X1 U22704 ( .A(\mem[332][3] ), .B(\mem[333][3] ), .S(n8416), .Z(n3752)
         );
  MUX2_X1 U22705 ( .A(n3752), .B(n3751), .S(n8280), .Z(n3753) );
  MUX2_X1 U22706 ( .A(\mem[330][3] ), .B(\mem[331][3] ), .S(n8411), .Z(n3754)
         );
  MUX2_X1 U22707 ( .A(\mem[328][3] ), .B(\mem[329][3] ), .S(n8412), .Z(n3755)
         );
  MUX2_X1 U22708 ( .A(n3755), .B(n3754), .S(n8279), .Z(n3756) );
  MUX2_X1 U22709 ( .A(n3756), .B(n3753), .S(n8264), .Z(n3757) );
  MUX2_X1 U22710 ( .A(\mem[326][3] ), .B(\mem[327][3] ), .S(n8413), .Z(n3758)
         );
  MUX2_X1 U22711 ( .A(\mem[324][3] ), .B(\mem[325][3] ), .S(n8420), .Z(n3759)
         );
  MUX2_X1 U22712 ( .A(n3759), .B(n3758), .S(n8275), .Z(n3760) );
  MUX2_X1 U22713 ( .A(\mem[322][3] ), .B(\mem[323][3] ), .S(n8421), .Z(n3761)
         );
  MUX2_X1 U22714 ( .A(\mem[320][3] ), .B(\mem[321][3] ), .S(n8422), .Z(n3762)
         );
  MUX2_X1 U22715 ( .A(n3762), .B(n3761), .S(n8274), .Z(n3763) );
  MUX2_X1 U22716 ( .A(n3763), .B(n3760), .S(n8242), .Z(n3764) );
  MUX2_X1 U22717 ( .A(n3764), .B(n3757), .S(n8209), .Z(n3765) );
  MUX2_X1 U22718 ( .A(n3765), .B(n3750), .S(n8186), .Z(n3766) );
  MUX2_X1 U22719 ( .A(n3766), .B(n3735), .S(n8185), .Z(n3767) );
  MUX2_X1 U22720 ( .A(\mem[318][3] ), .B(\mem[319][3] ), .S(n8434), .Z(n3768)
         );
  MUX2_X1 U22721 ( .A(\mem[316][3] ), .B(\mem[317][3] ), .S(n8364), .Z(n3769)
         );
  MUX2_X1 U22722 ( .A(n3769), .B(n3768), .S(n8343), .Z(n3770) );
  MUX2_X1 U22723 ( .A(\mem[314][3] ), .B(\mem[315][3] ), .S(n8373), .Z(n3771)
         );
  MUX2_X1 U22724 ( .A(\mem[312][3] ), .B(\mem[313][3] ), .S(n8532), .Z(n3772)
         );
  MUX2_X1 U22725 ( .A(n3772), .B(n3771), .S(n8350), .Z(n3773) );
  MUX2_X1 U22726 ( .A(n3773), .B(n3770), .S(n8265), .Z(n3774) );
  MUX2_X1 U22727 ( .A(\mem[310][3] ), .B(\mem[311][3] ), .S(n8470), .Z(n3775)
         );
  MUX2_X1 U22728 ( .A(\mem[308][3] ), .B(\mem[309][3] ), .S(n8436), .Z(n3776)
         );
  MUX2_X1 U22729 ( .A(n3776), .B(n3775), .S(n8351), .Z(n3777) );
  MUX2_X1 U22730 ( .A(\mem[306][3] ), .B(\mem[307][3] ), .S(n8534), .Z(n3778)
         );
  MUX2_X1 U22731 ( .A(\mem[304][3] ), .B(\mem[305][3] ), .S(n8539), .Z(n3779)
         );
  MUX2_X1 U22732 ( .A(n3779), .B(n3778), .S(n8352), .Z(n3780) );
  MUX2_X1 U22733 ( .A(n3780), .B(n3777), .S(n8264), .Z(n3781) );
  MUX2_X1 U22734 ( .A(n3781), .B(n3774), .S(n8211), .Z(n3782) );
  MUX2_X1 U22735 ( .A(\mem[302][3] ), .B(\mem[303][3] ), .S(n8371), .Z(n3783)
         );
  MUX2_X1 U22736 ( .A(\mem[300][3] ), .B(\mem[301][3] ), .S(n8397), .Z(n3784)
         );
  MUX2_X1 U22737 ( .A(n3784), .B(n3783), .S(n8347), .Z(n3785) );
  MUX2_X1 U22738 ( .A(\mem[298][3] ), .B(\mem[299][3] ), .S(n8512), .Z(n3786)
         );
  MUX2_X1 U22739 ( .A(\mem[296][3] ), .B(\mem[297][3] ), .S(n8485), .Z(n3787)
         );
  MUX2_X1 U22740 ( .A(n3787), .B(n3786), .S(n8348), .Z(n3788) );
  MUX2_X1 U22741 ( .A(n3788), .B(n3785), .S(n8243), .Z(n3789) );
  MUX2_X1 U22742 ( .A(\mem[294][3] ), .B(\mem[295][3] ), .S(n8365), .Z(n3790)
         );
  MUX2_X1 U22743 ( .A(\mem[292][3] ), .B(\mem[293][3] ), .S(n8387), .Z(n3791)
         );
  MUX2_X1 U22744 ( .A(n3791), .B(n3790), .S(n8349), .Z(n3792) );
  MUX2_X1 U22745 ( .A(\mem[290][3] ), .B(\mem[291][3] ), .S(n8386), .Z(n3793)
         );
  MUX2_X1 U22746 ( .A(\mem[288][3] ), .B(\mem[289][3] ), .S(n8382), .Z(n3794)
         );
  MUX2_X1 U22747 ( .A(n3794), .B(n3793), .S(n8353), .Z(n3795) );
  MUX2_X1 U22748 ( .A(n3795), .B(n3792), .S(n8224), .Z(n3796) );
  MUX2_X1 U22749 ( .A(n3796), .B(n3789), .S(N21), .Z(n3797) );
  MUX2_X1 U22750 ( .A(n3797), .B(n3782), .S(n8186), .Z(n3798) );
  MUX2_X1 U22751 ( .A(\mem[286][3] ), .B(\mem[287][3] ), .S(n8381), .Z(n3799)
         );
  MUX2_X1 U22752 ( .A(\mem[284][3] ), .B(\mem[285][3] ), .S(n8380), .Z(n3800)
         );
  MUX2_X1 U22753 ( .A(n3800), .B(n3799), .S(n8354), .Z(n3801) );
  MUX2_X1 U22754 ( .A(\mem[282][3] ), .B(\mem[283][3] ), .S(n8379), .Z(n3802)
         );
  MUX2_X1 U22755 ( .A(\mem[280][3] ), .B(\mem[281][3] ), .S(n8378), .Z(n3803)
         );
  MUX2_X1 U22756 ( .A(n3803), .B(n3802), .S(n8355), .Z(n3804) );
  MUX2_X1 U22757 ( .A(n3804), .B(n3801), .S(n8226), .Z(n3805) );
  MUX2_X1 U22758 ( .A(\mem[278][3] ), .B(\mem[279][3] ), .S(n8377), .Z(n3806)
         );
  MUX2_X1 U22759 ( .A(\mem[276][3] ), .B(\mem[277][3] ), .S(n8382), .Z(n3807)
         );
  MUX2_X1 U22760 ( .A(n3807), .B(n3806), .S(n8315), .Z(n3808) );
  MUX2_X1 U22761 ( .A(\mem[274][3] ), .B(\mem[275][3] ), .S(n8536), .Z(n3809)
         );
  MUX2_X1 U22762 ( .A(\mem[272][3] ), .B(\mem[273][3] ), .S(n8375), .Z(n3810)
         );
  MUX2_X1 U22763 ( .A(n3810), .B(n3809), .S(n8316), .Z(n3811) );
  MUX2_X1 U22764 ( .A(n3811), .B(n3808), .S(n8241), .Z(n3812) );
  MUX2_X1 U22765 ( .A(n3812), .B(n3805), .S(n8198), .Z(n3813) );
  MUX2_X1 U22766 ( .A(\mem[270][3] ), .B(\mem[271][3] ), .S(n8455), .Z(n3814)
         );
  MUX2_X1 U22767 ( .A(\mem[268][3] ), .B(\mem[269][3] ), .S(n8405), .Z(n3815)
         );
  MUX2_X1 U22768 ( .A(n3815), .B(n3814), .S(n8332), .Z(n3816) );
  MUX2_X1 U22769 ( .A(\mem[266][3] ), .B(\mem[267][3] ), .S(n8521), .Z(n3817)
         );
  MUX2_X1 U22770 ( .A(\mem[264][3] ), .B(\mem[265][3] ), .S(n8451), .Z(n3818)
         );
  MUX2_X1 U22771 ( .A(n3818), .B(n3817), .S(n8333), .Z(n3819) );
  MUX2_X1 U22772 ( .A(n3819), .B(n3816), .S(n8224), .Z(n3820) );
  MUX2_X1 U22773 ( .A(\mem[262][3] ), .B(\mem[263][3] ), .S(n8523), .Z(n3821)
         );
  MUX2_X1 U22774 ( .A(\mem[260][3] ), .B(\mem[261][3] ), .S(n8500), .Z(n3822)
         );
  MUX2_X1 U22775 ( .A(n3822), .B(n3821), .S(n8334), .Z(n3823) );
  MUX2_X1 U22776 ( .A(\mem[258][3] ), .B(\mem[259][3] ), .S(n8385), .Z(n3824)
         );
  MUX2_X1 U22777 ( .A(\mem[256][3] ), .B(\mem[257][3] ), .S(n8384), .Z(n3825)
         );
  MUX2_X1 U22778 ( .A(n3825), .B(n3824), .S(n8329), .Z(n3826) );
  MUX2_X1 U22779 ( .A(n3826), .B(n3823), .S(n8223), .Z(n3827) );
  MUX2_X1 U22780 ( .A(n3827), .B(n3820), .S(n8200), .Z(n3828) );
  MUX2_X1 U22781 ( .A(n3828), .B(n3813), .S(n8186), .Z(n3829) );
  MUX2_X1 U22782 ( .A(n3829), .B(n3798), .S(N23), .Z(n3830) );
  MUX2_X1 U22783 ( .A(n3830), .B(n3767), .S(n8180), .Z(n3831) );
  MUX2_X1 U22784 ( .A(n3831), .B(n3704), .S(n8177), .Z(n3832) );
  MUX2_X1 U22785 ( .A(\mem[254][3] ), .B(\mem[255][3] ), .S(n8383), .Z(n3833)
         );
  MUX2_X1 U22786 ( .A(\mem[252][3] ), .B(\mem[253][3] ), .S(n8373), .Z(n3834)
         );
  MUX2_X1 U22787 ( .A(n3834), .B(n3833), .S(n8330), .Z(n3835) );
  MUX2_X1 U22788 ( .A(\mem[250][3] ), .B(\mem[251][3] ), .S(n8372), .Z(n3836)
         );
  MUX2_X1 U22789 ( .A(\mem[248][3] ), .B(\mem[249][3] ), .S(n8371), .Z(n3837)
         );
  MUX2_X1 U22790 ( .A(n3837), .B(n3836), .S(n8331), .Z(n3838) );
  MUX2_X1 U22791 ( .A(n3838), .B(n3835), .S(n8263), .Z(n3839) );
  MUX2_X1 U22792 ( .A(\mem[246][3] ), .B(\mem[247][3] ), .S(n8393), .Z(n3840)
         );
  MUX2_X1 U22793 ( .A(\mem[244][3] ), .B(\mem[245][3] ), .S(n8394), .Z(n3841)
         );
  MUX2_X1 U22794 ( .A(n3841), .B(n3840), .S(n8338), .Z(n3842) );
  MUX2_X1 U22795 ( .A(\mem[242][3] ), .B(\mem[243][3] ), .S(n8390), .Z(n3843)
         );
  MUX2_X1 U22796 ( .A(\mem[240][3] ), .B(\mem[241][3] ), .S(n8391), .Z(n3844)
         );
  MUX2_X1 U22797 ( .A(n3844), .B(n3843), .S(n8339), .Z(n3845) );
  MUX2_X1 U22798 ( .A(n3845), .B(n3842), .S(n8224), .Z(n3846) );
  MUX2_X1 U22799 ( .A(n3846), .B(n3839), .S(n8199), .Z(n3847) );
  MUX2_X1 U22800 ( .A(\mem[238][3] ), .B(\mem[239][3] ), .S(n8392), .Z(n3848)
         );
  MUX2_X1 U22801 ( .A(\mem[236][3] ), .B(\mem[237][3] ), .S(n8389), .Z(n3849)
         );
  MUX2_X1 U22802 ( .A(n3849), .B(n3848), .S(n8340), .Z(n3850) );
  MUX2_X1 U22803 ( .A(\mem[234][3] ), .B(\mem[235][3] ), .S(n8386), .Z(n3851)
         );
  MUX2_X1 U22804 ( .A(\mem[232][3] ), .B(\mem[233][3] ), .S(N18), .Z(n3852) );
  MUX2_X1 U22805 ( .A(n3852), .B(n3851), .S(n8335), .Z(n3853) );
  MUX2_X1 U22806 ( .A(n3853), .B(n3850), .S(n8222), .Z(n3854) );
  MUX2_X1 U22807 ( .A(\mem[230][3] ), .B(\mem[231][3] ), .S(n8423), .Z(n3855)
         );
  MUX2_X1 U22808 ( .A(\mem[228][3] ), .B(\mem[229][3] ), .S(n8417), .Z(n3856)
         );
  MUX2_X1 U22809 ( .A(n3856), .B(n3855), .S(n8336), .Z(n3857) );
  MUX2_X1 U22810 ( .A(\mem[226][3] ), .B(\mem[227][3] ), .S(n8470), .Z(n3858)
         );
  MUX2_X1 U22811 ( .A(\mem[224][3] ), .B(\mem[225][3] ), .S(n8423), .Z(n3859)
         );
  MUX2_X1 U22812 ( .A(n3859), .B(n3858), .S(n8337), .Z(n3860) );
  MUX2_X1 U22813 ( .A(n3860), .B(n3857), .S(n8222), .Z(n3861) );
  MUX2_X1 U22814 ( .A(n3861), .B(n3854), .S(n8215), .Z(n3862) );
  MUX2_X1 U22815 ( .A(n3862), .B(n3847), .S(n8186), .Z(n3863) );
  MUX2_X1 U22816 ( .A(\mem[222][3] ), .B(\mem[223][3] ), .S(n8518), .Z(n3864)
         );
  MUX2_X1 U22817 ( .A(\mem[220][3] ), .B(\mem[221][3] ), .S(n8513), .Z(n3865)
         );
  MUX2_X1 U22818 ( .A(n3865), .B(n3864), .S(n8294), .Z(n3866) );
  MUX2_X1 U22819 ( .A(\mem[218][3] ), .B(\mem[219][3] ), .S(n8514), .Z(n3867)
         );
  MUX2_X1 U22820 ( .A(\mem[216][3] ), .B(\mem[217][3] ), .S(n8515), .Z(n3868)
         );
  MUX2_X1 U22821 ( .A(n3868), .B(n3867), .S(n8295), .Z(n3869) );
  MUX2_X1 U22822 ( .A(n3869), .B(n3866), .S(n8223), .Z(n3870) );
  MUX2_X1 U22823 ( .A(\mem[214][3] ), .B(\mem[215][3] ), .S(n8522), .Z(n3871)
         );
  MUX2_X1 U22824 ( .A(\mem[212][3] ), .B(\mem[213][3] ), .S(n8523), .Z(n3872)
         );
  MUX2_X1 U22825 ( .A(n3872), .B(n3871), .S(n8302), .Z(n3873) );
  MUX2_X1 U22826 ( .A(\mem[210][3] ), .B(\mem[211][3] ), .S(n8524), .Z(n3874)
         );
  MUX2_X1 U22827 ( .A(\mem[208][3] ), .B(\mem[209][3] ), .S(n8519), .Z(n3875)
         );
  MUX2_X1 U22828 ( .A(n3875), .B(n3874), .S(n8303), .Z(n3876) );
  MUX2_X1 U22829 ( .A(n3876), .B(n3873), .S(n8264), .Z(n3877) );
  MUX2_X1 U22830 ( .A(n3877), .B(n3870), .S(n8219), .Z(n3878) );
  MUX2_X1 U22831 ( .A(\mem[206][3] ), .B(\mem[207][3] ), .S(n8520), .Z(n3879)
         );
  MUX2_X1 U22832 ( .A(\mem[204][3] ), .B(\mem[205][3] ), .S(n8521), .Z(n3880)
         );
  MUX2_X1 U22833 ( .A(n3880), .B(n3879), .S(n8304), .Z(n3881) );
  MUX2_X1 U22834 ( .A(\mem[202][3] ), .B(\mem[203][3] ), .S(n8528), .Z(n3882)
         );
  MUX2_X1 U22835 ( .A(\mem[200][3] ), .B(\mem[201][3] ), .S(n8529), .Z(n3883)
         );
  MUX2_X1 U22836 ( .A(n3883), .B(n3882), .S(n8299), .Z(n3884) );
  MUX2_X1 U22837 ( .A(n3884), .B(n3881), .S(n8222), .Z(n3885) );
  MUX2_X1 U22838 ( .A(\mem[198][3] ), .B(\mem[199][3] ), .S(n8495), .Z(n3886)
         );
  MUX2_X1 U22839 ( .A(\mem[196][3] ), .B(\mem[197][3] ), .S(n8496), .Z(n3887)
         );
  MUX2_X1 U22840 ( .A(n3887), .B(n3886), .S(n8300), .Z(n3888) );
  MUX2_X1 U22841 ( .A(\mem[194][3] ), .B(\mem[195][3] ), .S(n8497), .Z(n3889)
         );
  MUX2_X1 U22842 ( .A(\mem[192][3] ), .B(\mem[193][3] ), .S(n8504), .Z(n3890)
         );
  MUX2_X1 U22843 ( .A(n3890), .B(n3889), .S(n8301), .Z(n3891) );
  MUX2_X1 U22844 ( .A(n3891), .B(n3888), .S(n8221), .Z(n3892) );
  MUX2_X1 U22845 ( .A(n3892), .B(n3885), .S(n8197), .Z(n3893) );
  MUX2_X1 U22846 ( .A(n3893), .B(n3878), .S(n8186), .Z(n3894) );
  MUX2_X1 U22847 ( .A(n3894), .B(n3863), .S(n8182), .Z(n3895) );
  MUX2_X1 U22848 ( .A(\mem[190][3] ), .B(\mem[191][3] ), .S(n8505), .Z(n3896)
         );
  MUX2_X1 U22849 ( .A(\mem[188][3] ), .B(\mem[189][3] ), .S(n8506), .Z(n3897)
         );
  MUX2_X1 U22850 ( .A(n3897), .B(n3896), .S(n8287), .Z(n3898) );
  MUX2_X1 U22851 ( .A(\mem[186][3] ), .B(\mem[187][3] ), .S(n8501), .Z(n3899)
         );
  MUX2_X1 U22852 ( .A(\mem[184][3] ), .B(\mem[185][3] ), .S(n8502), .Z(n3900)
         );
  MUX2_X1 U22853 ( .A(n3900), .B(n3899), .S(n8323), .Z(n3901) );
  MUX2_X1 U22854 ( .A(n3901), .B(n3898), .S(n8222), .Z(n3902) );
  MUX2_X1 U22855 ( .A(\mem[182][3] ), .B(\mem[183][3] ), .S(n8503), .Z(n3903)
         );
  MUX2_X1 U22856 ( .A(\mem[180][3] ), .B(\mem[181][3] ), .S(n8510), .Z(n3904)
         );
  MUX2_X1 U22857 ( .A(n3904), .B(n3903), .S(n8273), .Z(n3905) );
  MUX2_X1 U22858 ( .A(\mem[178][3] ), .B(\mem[179][3] ), .S(n8511), .Z(n3906)
         );
  MUX2_X1 U22859 ( .A(\mem[176][3] ), .B(\mem[177][3] ), .S(n8512), .Z(n3907)
         );
  MUX2_X1 U22860 ( .A(n3907), .B(n3906), .S(n8284), .Z(n3908) );
  MUX2_X1 U22861 ( .A(n3908), .B(n3905), .S(n8221), .Z(n3909) );
  MUX2_X1 U22862 ( .A(n3909), .B(n3902), .S(n8201), .Z(n3910) );
  MUX2_X1 U22863 ( .A(\mem[174][3] ), .B(\mem[175][3] ), .S(n8478), .Z(n3911)
         );
  MUX2_X1 U22864 ( .A(\mem[172][3] ), .B(\mem[173][3] ), .S(n8479), .Z(n3912)
         );
  MUX2_X1 U22865 ( .A(n3912), .B(n3911), .S(n8266), .Z(n3913) );
  MUX2_X1 U22866 ( .A(\mem[170][3] ), .B(\mem[171][3] ), .S(n8486), .Z(n3914)
         );
  MUX2_X1 U22867 ( .A(\mem[168][3] ), .B(\mem[169][3] ), .S(n8487), .Z(n3915)
         );
  MUX2_X1 U22868 ( .A(n3915), .B(n3914), .S(n8280), .Z(n3916) );
  MUX2_X1 U22869 ( .A(n3916), .B(n3913), .S(n8254), .Z(n3917) );
  MUX2_X1 U22870 ( .A(\mem[166][3] ), .B(\mem[167][3] ), .S(n8488), .Z(n3918)
         );
  MUX2_X1 U22871 ( .A(\mem[164][3] ), .B(\mem[165][3] ), .S(n8483), .Z(n3919)
         );
  MUX2_X1 U22872 ( .A(n3919), .B(n3918), .S(n8314), .Z(n3920) );
  MUX2_X1 U22873 ( .A(\mem[162][3] ), .B(\mem[163][3] ), .S(n8484), .Z(n3921)
         );
  MUX2_X1 U22874 ( .A(\mem[160][3] ), .B(\mem[161][3] ), .S(n8485), .Z(n3922)
         );
  MUX2_X1 U22875 ( .A(n3922), .B(n3921), .S(n8315), .Z(n3923) );
  MUX2_X1 U22876 ( .A(n3923), .B(n3920), .S(n8226), .Z(n3924) );
  MUX2_X1 U22877 ( .A(n3924), .B(n3917), .S(n8202), .Z(n3925) );
  MUX2_X1 U22878 ( .A(n3925), .B(n3910), .S(n8186), .Z(n3926) );
  MUX2_X1 U22879 ( .A(\mem[158][3] ), .B(\mem[159][3] ), .S(n8492), .Z(n3927)
         );
  MUX2_X1 U22880 ( .A(\mem[156][3] ), .B(\mem[157][3] ), .S(n8493), .Z(n3928)
         );
  MUX2_X1 U22881 ( .A(n3928), .B(n3927), .S(n8316), .Z(n3929) );
  MUX2_X1 U22882 ( .A(\mem[154][3] ), .B(\mem[155][3] ), .S(n8494), .Z(n3930)
         );
  MUX2_X1 U22883 ( .A(\mem[152][3] ), .B(\mem[153][3] ), .S(n8489), .Z(n3931)
         );
  MUX2_X1 U22884 ( .A(n3931), .B(n3930), .S(n8311), .Z(n3932) );
  MUX2_X1 U22885 ( .A(n3932), .B(n3929), .S(n8220), .Z(n3933) );
  MUX2_X1 U22886 ( .A(\mem[150][3] ), .B(\mem[151][3] ), .S(n8475), .Z(n3934)
         );
  MUX2_X1 U22887 ( .A(\mem[148][3] ), .B(\mem[149][3] ), .S(n8366), .Z(n3935)
         );
  MUX2_X1 U22888 ( .A(n3935), .B(n3934), .S(n8312), .Z(n3936) );
  MUX2_X1 U22889 ( .A(\mem[146][3] ), .B(\mem[147][3] ), .S(n8420), .Z(n3937)
         );
  MUX2_X1 U22890 ( .A(\mem[144][3] ), .B(\mem[145][3] ), .S(n8381), .Z(n3938)
         );
  MUX2_X1 U22891 ( .A(n3938), .B(n3937), .S(n8313), .Z(n3939) );
  MUX2_X1 U22892 ( .A(n3939), .B(n3936), .S(n8254), .Z(n3940) );
  MUX2_X1 U22893 ( .A(n3940), .B(n3933), .S(n8203), .Z(n3941) );
  MUX2_X1 U22894 ( .A(\mem[142][3] ), .B(\mem[143][3] ), .S(N18), .Z(n3942) );
  MUX2_X1 U22895 ( .A(\mem[140][3] ), .B(\mem[141][3] ), .S(n8433), .Z(n3943)
         );
  MUX2_X1 U22896 ( .A(n3943), .B(n3942), .S(n8320), .Z(n3944) );
  MUX2_X1 U22897 ( .A(\mem[138][3] ), .B(\mem[139][3] ), .S(n8475), .Z(n3945)
         );
  MUX2_X1 U22898 ( .A(\mem[136][3] ), .B(\mem[137][3] ), .S(n8476), .Z(n3946)
         );
  MUX2_X1 U22899 ( .A(n3946), .B(n3945), .S(n8321), .Z(n3947) );
  MUX2_X1 U22900 ( .A(n3947), .B(n3944), .S(n8225), .Z(n3948) );
  MUX2_X1 U22901 ( .A(\mem[134][3] ), .B(\mem[135][3] ), .S(n8471), .Z(n3949)
         );
  MUX2_X1 U22902 ( .A(\mem[132][3] ), .B(\mem[133][3] ), .S(n8472), .Z(n3950)
         );
  MUX2_X1 U22903 ( .A(n3950), .B(n3949), .S(n8322), .Z(n3951) );
  MUX2_X1 U22904 ( .A(\mem[130][3] ), .B(\mem[131][3] ), .S(n8363), .Z(n3952)
         );
  MUX2_X1 U22905 ( .A(\mem[128][3] ), .B(\mem[129][3] ), .S(n8537), .Z(n3953)
         );
  MUX2_X1 U22906 ( .A(n3953), .B(n3952), .S(n8317), .Z(n3954) );
  MUX2_X1 U22907 ( .A(n3954), .B(n3951), .S(n8263), .Z(n3955) );
  MUX2_X1 U22908 ( .A(n3955), .B(n3948), .S(n8204), .Z(n3956) );
  MUX2_X1 U22909 ( .A(n3956), .B(n3941), .S(n8186), .Z(n3957) );
  MUX2_X1 U22910 ( .A(n3957), .B(n3926), .S(n8182), .Z(n3958) );
  MUX2_X1 U22911 ( .A(n3958), .B(n3895), .S(n8180), .Z(n3959) );
  MUX2_X1 U22912 ( .A(\mem[126][3] ), .B(\mem[127][3] ), .S(n8394), .Z(n3960)
         );
  MUX2_X1 U22913 ( .A(\mem[124][3] ), .B(\mem[125][3] ), .S(n8390), .Z(n3961)
         );
  MUX2_X1 U22914 ( .A(n3961), .B(n3960), .S(n8324), .Z(n3962) );
  MUX2_X1 U22915 ( .A(\mem[122][3] ), .B(\mem[123][3] ), .S(n8391), .Z(n3963)
         );
  MUX2_X1 U22916 ( .A(\mem[120][3] ), .B(\mem[121][3] ), .S(n8392), .Z(n3964)
         );
  MUX2_X1 U22917 ( .A(n3964), .B(n3963), .S(n8316), .Z(n3965) );
  MUX2_X1 U22918 ( .A(n3965), .B(n3962), .S(n8253), .Z(n3966) );
  MUX2_X1 U22919 ( .A(\mem[118][3] ), .B(\mem[119][3] ), .S(n8389), .Z(n3967)
         );
  MUX2_X1 U22920 ( .A(\mem[116][3] ), .B(\mem[117][3] ), .S(n8402), .Z(n3968)
         );
  MUX2_X1 U22921 ( .A(n3968), .B(n3967), .S(n8352), .Z(n3969) );
  MUX2_X1 U22922 ( .A(\mem[114][3] ), .B(\mem[115][3] ), .S(n8499), .Z(n3970)
         );
  MUX2_X1 U22923 ( .A(\mem[112][3] ), .B(\mem[113][3] ), .S(n8403), .Z(n3971)
         );
  MUX2_X1 U22924 ( .A(n3971), .B(n3970), .S(n8325), .Z(n3972) );
  MUX2_X1 U22925 ( .A(n3972), .B(n3969), .S(n8237), .Z(n3973) );
  MUX2_X1 U22926 ( .A(n3973), .B(n3966), .S(n8213), .Z(n3974) );
  MUX2_X1 U22927 ( .A(\mem[110][3] ), .B(\mem[111][3] ), .S(n8393), .Z(n3975)
         );
  MUX2_X1 U22928 ( .A(\mem[108][3] ), .B(\mem[109][3] ), .S(n8432), .Z(n3976)
         );
  MUX2_X1 U22929 ( .A(n3976), .B(n3975), .S(n8292), .Z(n3977) );
  MUX2_X1 U22930 ( .A(\mem[106][3] ), .B(\mem[107][3] ), .S(n8461), .Z(n3978)
         );
  MUX2_X1 U22931 ( .A(\mem[104][3] ), .B(\mem[105][3] ), .S(n8414), .Z(n3979)
         );
  MUX2_X1 U22932 ( .A(n3979), .B(n3978), .S(n8286), .Z(n3980) );
  MUX2_X1 U22933 ( .A(n3980), .B(n3977), .S(n8225), .Z(n3981) );
  MUX2_X1 U22934 ( .A(\mem[102][3] ), .B(\mem[103][3] ), .S(n8536), .Z(n3982)
         );
  MUX2_X1 U22935 ( .A(\mem[100][3] ), .B(\mem[101][3] ), .S(n8531), .Z(n3983)
         );
  MUX2_X1 U22936 ( .A(n3983), .B(n3982), .S(n8331), .Z(n3984) );
  MUX2_X1 U22937 ( .A(\mem[98][3] ), .B(\mem[99][3] ), .S(n8532), .Z(n3985) );
  MUX2_X1 U22938 ( .A(\mem[96][3] ), .B(\mem[97][3] ), .S(n8533), .Z(n3986) );
  MUX2_X1 U22939 ( .A(n3986), .B(n3985), .S(n8298), .Z(n3987) );
  MUX2_X1 U22940 ( .A(n3987), .B(n3984), .S(n8242), .Z(n3988) );
  MUX2_X1 U22941 ( .A(n3988), .B(n3981), .S(n8219), .Z(n3989) );
  MUX2_X1 U22942 ( .A(n3989), .B(n3974), .S(n8187), .Z(n3990) );
  MUX2_X1 U22943 ( .A(\mem[94][3] ), .B(\mem[95][3] ), .S(n8398), .Z(n3991) );
  MUX2_X1 U22944 ( .A(\mem[92][3] ), .B(\mem[93][3] ), .S(n8399), .Z(n3992) );
  MUX2_X1 U22945 ( .A(n3992), .B(n3991), .S(n8274), .Z(n3993) );
  MUX2_X1 U22946 ( .A(\mem[90][3] ), .B(\mem[91][3] ), .S(n8400), .Z(n3994) );
  MUX2_X1 U22947 ( .A(\mem[88][3] ), .B(\mem[89][3] ), .S(n8395), .Z(n3995) );
  MUX2_X1 U22948 ( .A(n3995), .B(n3994), .S(n8284), .Z(n3996) );
  MUX2_X1 U22949 ( .A(n3996), .B(n3993), .S(n8259), .Z(n3997) );
  MUX2_X1 U22950 ( .A(\mem[86][3] ), .B(\mem[87][3] ), .S(n8396), .Z(n3998) );
  MUX2_X1 U22951 ( .A(\mem[84][3] ), .B(\mem[85][3] ), .S(n8397), .Z(n3999) );
  MUX2_X1 U22952 ( .A(n3999), .B(n3998), .S(n8285), .Z(n4000) );
  MUX2_X1 U22953 ( .A(\mem[82][3] ), .B(\mem[83][3] ), .S(n8404), .Z(n4001) );
  MUX2_X1 U22954 ( .A(\mem[80][3] ), .B(\mem[81][3] ), .S(n8405), .Z(n4002) );
  MUX2_X1 U22955 ( .A(n4002), .B(n4001), .S(n8286), .Z(n4003) );
  MUX2_X1 U22956 ( .A(n4003), .B(n4000), .S(n8229), .Z(n4004) );
  MUX2_X1 U22957 ( .A(n4004), .B(n3997), .S(n8197), .Z(n4005) );
  MUX2_X1 U22958 ( .A(\mem[78][3] ), .B(\mem[79][3] ), .S(n8446), .Z(n4006) );
  MUX2_X1 U22959 ( .A(\mem[76][3] ), .B(\mem[77][3] ), .S(n8522), .Z(n4007) );
  MUX2_X1 U22960 ( .A(n4007), .B(n4006), .S(n8277), .Z(n4008) );
  MUX2_X1 U22961 ( .A(\mem[74][3] ), .B(\mem[75][3] ), .S(n8496), .Z(n4009) );
  MUX2_X1 U22962 ( .A(\mem[72][3] ), .B(\mem[73][3] ), .S(n8361), .Z(n4010) );
  MUX2_X1 U22963 ( .A(n4010), .B(n4009), .S(n8274), .Z(n4011) );
  MUX2_X1 U22964 ( .A(n4011), .B(n4008), .S(n8228), .Z(n4012) );
  MUX2_X1 U22965 ( .A(\mem[70][3] ), .B(\mem[71][3] ), .S(n8491), .Z(n4013) );
  MUX2_X1 U22966 ( .A(\mem[68][3] ), .B(\mem[69][3] ), .S(n8460), .Z(n4014) );
  MUX2_X1 U22967 ( .A(n4014), .B(n4013), .S(n8273), .Z(n4015) );
  MUX2_X1 U22968 ( .A(\mem[66][3] ), .B(\mem[67][3] ), .S(n8405), .Z(n4016) );
  MUX2_X1 U22969 ( .A(\mem[64][3] ), .B(\mem[65][3] ), .S(n8506), .Z(n4017) );
  MUX2_X1 U22970 ( .A(n4017), .B(n4016), .S(n8272), .Z(n4018) );
  MUX2_X1 U22971 ( .A(n4018), .B(n4015), .S(n8236), .Z(n4019) );
  MUX2_X1 U22972 ( .A(n4019), .B(n4012), .S(n8207), .Z(n4020) );
  MUX2_X1 U22973 ( .A(n4020), .B(n4005), .S(n8187), .Z(n4021) );
  MUX2_X1 U22974 ( .A(n4021), .B(n3990), .S(n8182), .Z(n4022) );
  MUX2_X1 U22975 ( .A(\mem[62][3] ), .B(\mem[63][3] ), .S(n8487), .Z(n4023) );
  MUX2_X1 U22976 ( .A(\mem[60][3] ), .B(\mem[61][3] ), .S(n8431), .Z(n4024) );
  MUX2_X1 U22977 ( .A(n4024), .B(n4023), .S(n8271), .Z(n4025) );
  MUX2_X1 U22978 ( .A(\mem[58][3] ), .B(\mem[59][3] ), .S(n8408), .Z(n4026) );
  MUX2_X1 U22979 ( .A(\mem[56][3] ), .B(\mem[57][3] ), .S(n8455), .Z(n4027) );
  MUX2_X1 U22980 ( .A(n4027), .B(n4026), .S(n8266), .Z(n4028) );
  MUX2_X1 U22981 ( .A(n4028), .B(n4025), .S(n8245), .Z(n4029) );
  MUX2_X1 U22982 ( .A(\mem[54][3] ), .B(\mem[55][3] ), .S(n8538), .Z(n4030) );
  MUX2_X1 U22983 ( .A(\mem[52][3] ), .B(\mem[53][3] ), .S(N18), .Z(n4031) );
  MUX2_X1 U22984 ( .A(n4031), .B(n4030), .S(n8267), .Z(n4032) );
  MUX2_X1 U22985 ( .A(\mem[50][3] ), .B(\mem[51][3] ), .S(n8428), .Z(n4033) );
  MUX2_X1 U22986 ( .A(\mem[48][3] ), .B(\mem[49][3] ), .S(n8415), .Z(n4034) );
  MUX2_X1 U22987 ( .A(n4034), .B(n4033), .S(n8268), .Z(n4035) );
  MUX2_X1 U22988 ( .A(n4035), .B(n4032), .S(n8248), .Z(n4036) );
  MUX2_X1 U22989 ( .A(n4036), .B(n4029), .S(n8208), .Z(n4037) );
  MUX2_X1 U22990 ( .A(\mem[46][3] ), .B(\mem[47][3] ), .S(n8358), .Z(n4038) );
  MUX2_X1 U22991 ( .A(\mem[44][3] ), .B(\mem[45][3] ), .S(n8539), .Z(n4039) );
  MUX2_X1 U22992 ( .A(n4039), .B(n4038), .S(n8269), .Z(n4040) );
  MUX2_X1 U22993 ( .A(\mem[42][3] ), .B(\mem[43][3] ), .S(n8362), .Z(n4041) );
  MUX2_X1 U22994 ( .A(\mem[40][3] ), .B(\mem[41][3] ), .S(n8363), .Z(n4042) );
  MUX2_X1 U22995 ( .A(n4042), .B(n4041), .S(n8356), .Z(n4043) );
  MUX2_X1 U22996 ( .A(n4043), .B(n4040), .S(n8221), .Z(n4044) );
  MUX2_X1 U22997 ( .A(\mem[38][3] ), .B(\mem[39][3] ), .S(n8364), .Z(n4045) );
  MUX2_X1 U22998 ( .A(\mem[36][3] ), .B(\mem[37][3] ), .S(n8357), .Z(n4046) );
  MUX2_X1 U22999 ( .A(n4046), .B(n4045), .S(n8270), .Z(n4047) );
  MUX2_X1 U23000 ( .A(\mem[34][3] ), .B(\mem[35][3] ), .S(n8359), .Z(n4048) );
  MUX2_X1 U23001 ( .A(\mem[32][3] ), .B(\mem[33][3] ), .S(n8360), .Z(n4049) );
  MUX2_X1 U23002 ( .A(n4049), .B(n4048), .S(n8336), .Z(n4050) );
  MUX2_X1 U23003 ( .A(n4050), .B(n4047), .S(n8238), .Z(n4051) );
  MUX2_X1 U23004 ( .A(n4051), .B(n4044), .S(n8209), .Z(n4052) );
  MUX2_X1 U23005 ( .A(n4052), .B(n4037), .S(n8187), .Z(n4053) );
  MUX2_X1 U23006 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n8426), .Z(n4054) );
  MUX2_X1 U23007 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n8427), .Z(n4055) );
  MUX2_X1 U23008 ( .A(n4055), .B(n4054), .S(n8353), .Z(n4056) );
  MUX2_X1 U23009 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n8428), .Z(n4057) );
  MUX2_X1 U23010 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n8424), .Z(n4058) );
  MUX2_X1 U23011 ( .A(n4058), .B(n4057), .S(n8354), .Z(n4059) );
  MUX2_X1 U23012 ( .A(n4059), .B(n4056), .S(n8238), .Z(n4060) );
  MUX2_X1 U23013 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n8425), .Z(n4061) );
  MUX2_X1 U23014 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n8375), .Z(n4062) );
  MUX2_X1 U23015 ( .A(n4062), .B(n4061), .S(n8355), .Z(n4063) );
  MUX2_X1 U23016 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n8409), .Z(n4064) );
  MUX2_X1 U23017 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n8404), .Z(n4065) );
  MUX2_X1 U23018 ( .A(n4065), .B(n4064), .S(N19), .Z(n4066) );
  MUX2_X1 U23019 ( .A(n4066), .B(n4063), .S(n8263), .Z(n4067) );
  MUX2_X1 U23020 ( .A(n4067), .B(n4060), .S(n8210), .Z(n4068) );
  MUX2_X1 U23021 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n8384), .Z(n4069) );
  MUX2_X1 U23022 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n8383), .Z(n4070) );
  MUX2_X1 U23023 ( .A(n4070), .B(n4069), .S(n8356), .Z(n4071) );
  MUX2_X1 U23024 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n8371), .Z(n4072) );
  MUX2_X1 U23025 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n8369), .Z(n4073) );
  MUX2_X1 U23026 ( .A(n4073), .B(n4072), .S(n8269), .Z(n4074) );
  MUX2_X1 U23027 ( .A(n4074), .B(n4071), .S(n8237), .Z(n4075) );
  MUX2_X1 U23028 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n8441), .Z(n4076) );
  MUX2_X1 U23029 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n8442), .Z(n4077) );
  MUX2_X1 U23030 ( .A(n4077), .B(n4076), .S(n8317), .Z(n4078) );
  MUX2_X1 U23031 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n8443), .Z(n4079) );
  MUX2_X1 U23032 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n8450), .Z(n4080) );
  MUX2_X1 U23033 ( .A(n4080), .B(n4079), .S(n8321), .Z(n4081) );
  MUX2_X1 U23034 ( .A(n4081), .B(n4078), .S(n8265), .Z(n4082) );
  MUX2_X1 U23035 ( .A(n4082), .B(n4075), .S(n8206), .Z(n4083) );
  MUX2_X1 U23036 ( .A(n4083), .B(n4068), .S(n8187), .Z(n4084) );
  MUX2_X1 U23037 ( .A(n4084), .B(n4053), .S(n8183), .Z(n4085) );
  MUX2_X1 U23038 ( .A(n4085), .B(n4022), .S(n8178), .Z(n4086) );
  MUX2_X1 U23039 ( .A(n4086), .B(n3959), .S(n8177), .Z(n4087) );
  MUX2_X1 U23040 ( .A(n4087), .B(n3832), .S(N26), .Z(n4088) );
  MUX2_X1 U23041 ( .A(n4088), .B(n3577), .S(N27), .Z(N32) );
  MUX2_X1 U23042 ( .A(\mem[1022][4] ), .B(\mem[1023][4] ), .S(n8451), .Z(n4089) );
  MUX2_X1 U23043 ( .A(\mem[1020][4] ), .B(\mem[1021][4] ), .S(n8452), .Z(n4090) );
  MUX2_X1 U23044 ( .A(n4090), .B(n4089), .S(n8322), .Z(n4091) );
  MUX2_X1 U23045 ( .A(\mem[1018][4] ), .B(\mem[1019][4] ), .S(n8447), .Z(n4092) );
  MUX2_X1 U23046 ( .A(\mem[1016][4] ), .B(\mem[1017][4] ), .S(n8448), .Z(n4093) );
  MUX2_X1 U23047 ( .A(n4093), .B(n4092), .S(n8317), .Z(n4094) );
  MUX2_X1 U23048 ( .A(n4094), .B(n4091), .S(n8230), .Z(n4095) );
  MUX2_X1 U23049 ( .A(\mem[1014][4] ), .B(\mem[1015][4] ), .S(n8449), .Z(n4096) );
  MUX2_X1 U23050 ( .A(\mem[1012][4] ), .B(\mem[1013][4] ), .S(n8456), .Z(n4097) );
  MUX2_X1 U23051 ( .A(n4097), .B(n4096), .S(n8318), .Z(n4098) );
  MUX2_X1 U23052 ( .A(\mem[1010][4] ), .B(\mem[1011][4] ), .S(n8457), .Z(n4099) );
  MUX2_X1 U23053 ( .A(\mem[1008][4] ), .B(\mem[1009][4] ), .S(n8458), .Z(n4100) );
  MUX2_X1 U23054 ( .A(n4100), .B(n4099), .S(n8319), .Z(n4101) );
  MUX2_X1 U23055 ( .A(n4101), .B(n4098), .S(n8235), .Z(n4102) );
  MUX2_X1 U23056 ( .A(n4102), .B(n4095), .S(n8212), .Z(n4103) );
  MUX2_X1 U23057 ( .A(\mem[1006][4] ), .B(\mem[1007][4] ), .S(n8490), .Z(n4104) );
  MUX2_X1 U23058 ( .A(\mem[1004][4] ), .B(\mem[1005][4] ), .S(n8432), .Z(n4105) );
  MUX2_X1 U23059 ( .A(n4105), .B(n4104), .S(n8329), .Z(n4106) );
  MUX2_X1 U23060 ( .A(\mem[1002][4] ), .B(\mem[1003][4] ), .S(n8433), .Z(n4107) );
  MUX2_X1 U23061 ( .A(\mem[1000][4] ), .B(\mem[1001][4] ), .S(n8434), .Z(n4108) );
  MUX2_X1 U23062 ( .A(n4108), .B(n4107), .S(n8330), .Z(n4109) );
  MUX2_X1 U23063 ( .A(n4109), .B(n4106), .S(n8237), .Z(n4110) );
  MUX2_X1 U23064 ( .A(\mem[998][4] ), .B(\mem[999][4] ), .S(n8429), .Z(n4111)
         );
  MUX2_X1 U23065 ( .A(\mem[996][4] ), .B(\mem[997][4] ), .S(n8430), .Z(n4112)
         );
  MUX2_X1 U23066 ( .A(n4112), .B(n4111), .S(n8331), .Z(n4113) );
  MUX2_X1 U23067 ( .A(\mem[994][4] ), .B(\mem[995][4] ), .S(n8431), .Z(n4114)
         );
  MUX2_X1 U23068 ( .A(\mem[992][4] ), .B(\mem[993][4] ), .S(n8438), .Z(n4115)
         );
  MUX2_X1 U23069 ( .A(n4115), .B(n4114), .S(n8338), .Z(n4116) );
  MUX2_X1 U23070 ( .A(n4116), .B(n4113), .S(n8252), .Z(n4117) );
  MUX2_X1 U23071 ( .A(n4117), .B(n4110), .S(n8213), .Z(n4118) );
  MUX2_X1 U23072 ( .A(n4118), .B(n4103), .S(n8187), .Z(n4119) );
  MUX2_X1 U23073 ( .A(\mem[990][4] ), .B(\mem[991][4] ), .S(n8439), .Z(n4120)
         );
  MUX2_X1 U23074 ( .A(\mem[988][4] ), .B(\mem[989][4] ), .S(n8440), .Z(n4121)
         );
  MUX2_X1 U23075 ( .A(n4121), .B(n4120), .S(n8339), .Z(n4122) );
  MUX2_X1 U23076 ( .A(\mem[986][4] ), .B(\mem[987][4] ), .S(n8435), .Z(n4123)
         );
  MUX2_X1 U23077 ( .A(\mem[984][4] ), .B(\mem[985][4] ), .S(n8436), .Z(n4124)
         );
  MUX2_X1 U23078 ( .A(n4124), .B(n4123), .S(n8340), .Z(n4125) );
  MUX2_X1 U23079 ( .A(n4125), .B(n4122), .S(n8262), .Z(n4126) );
  MUX2_X1 U23080 ( .A(\mem[982][4] ), .B(\mem[983][4] ), .S(n8433), .Z(n4127)
         );
  MUX2_X1 U23081 ( .A(\mem[980][4] ), .B(\mem[981][4] ), .S(n8434), .Z(n4128)
         );
  MUX2_X1 U23082 ( .A(n4128), .B(n4127), .S(n8335), .Z(n4129) );
  MUX2_X1 U23083 ( .A(\mem[978][4] ), .B(\mem[979][4] ), .S(n8429), .Z(n4130)
         );
  MUX2_X1 U23084 ( .A(\mem[976][4] ), .B(\mem[977][4] ), .S(n8430), .Z(n4131)
         );
  MUX2_X1 U23085 ( .A(n4131), .B(n4130), .S(n8337), .Z(n4132) );
  MUX2_X1 U23086 ( .A(n4132), .B(n4129), .S(n8247), .Z(n4133) );
  MUX2_X1 U23087 ( .A(n4133), .B(n4126), .S(n8214), .Z(n4134) );
  MUX2_X1 U23088 ( .A(\mem[974][4] ), .B(\mem[975][4] ), .S(n8431), .Z(n4135)
         );
  MUX2_X1 U23089 ( .A(\mem[972][4] ), .B(\mem[973][4] ), .S(n8438), .Z(n4136)
         );
  MUX2_X1 U23090 ( .A(n4136), .B(n4135), .S(n8345), .Z(n4137) );
  MUX2_X1 U23091 ( .A(\mem[970][4] ), .B(\mem[971][4] ), .S(n8439), .Z(n4138)
         );
  MUX2_X1 U23092 ( .A(\mem[968][4] ), .B(\mem[969][4] ), .S(n8440), .Z(n4139)
         );
  MUX2_X1 U23093 ( .A(n4139), .B(n4138), .S(n8346), .Z(n4140) );
  MUX2_X1 U23094 ( .A(n4140), .B(n4137), .S(n8248), .Z(n4141) );
  MUX2_X1 U23095 ( .A(\mem[966][4] ), .B(\mem[967][4] ), .S(n8435), .Z(n4142)
         );
  MUX2_X1 U23096 ( .A(\mem[964][4] ), .B(\mem[965][4] ), .S(n8436), .Z(n4143)
         );
  MUX2_X1 U23097 ( .A(n4143), .B(n4142), .S(n8341), .Z(n4144) );
  MUX2_X1 U23098 ( .A(\mem[962][4] ), .B(\mem[963][4] ), .S(n8437), .Z(n4145)
         );
  MUX2_X1 U23099 ( .A(\mem[960][4] ), .B(\mem[961][4] ), .S(n8444), .Z(n4146)
         );
  MUX2_X1 U23100 ( .A(n4146), .B(n4145), .S(n8342), .Z(n4147) );
  MUX2_X1 U23101 ( .A(n4147), .B(n4144), .S(n8257), .Z(n4148) );
  MUX2_X1 U23102 ( .A(n4148), .B(n4141), .S(n8215), .Z(n4149) );
  MUX2_X1 U23103 ( .A(n4149), .B(n4134), .S(n8187), .Z(n4150) );
  MUX2_X1 U23104 ( .A(n4150), .B(n4119), .S(n8181), .Z(n4151) );
  MUX2_X1 U23105 ( .A(\mem[958][4] ), .B(\mem[959][4] ), .S(n8414), .Z(n4152)
         );
  MUX2_X1 U23106 ( .A(\mem[956][4] ), .B(\mem[957][4] ), .S(n8415), .Z(n4153)
         );
  MUX2_X1 U23107 ( .A(n4153), .B(n4152), .S(n8324), .Z(n4154) );
  MUX2_X1 U23108 ( .A(\mem[954][4] ), .B(\mem[955][4] ), .S(n8416), .Z(n4155)
         );
  MUX2_X1 U23109 ( .A(\mem[952][4] ), .B(\mem[953][4] ), .S(n8411), .Z(n4156)
         );
  MUX2_X1 U23110 ( .A(n4156), .B(n4155), .S(n8325), .Z(n4157) );
  MUX2_X1 U23111 ( .A(n4157), .B(n4154), .S(n8240), .Z(n4158) );
  MUX2_X1 U23112 ( .A(\mem[950][4] ), .B(\mem[951][4] ), .S(n8412), .Z(n4159)
         );
  MUX2_X1 U23113 ( .A(\mem[948][4] ), .B(\mem[949][4] ), .S(n8413), .Z(n4160)
         );
  MUX2_X1 U23114 ( .A(n4160), .B(n4159), .S(n8332), .Z(n4161) );
  MUX2_X1 U23115 ( .A(\mem[946][4] ), .B(\mem[947][4] ), .S(n8420), .Z(n4162)
         );
  MUX2_X1 U23116 ( .A(\mem[944][4] ), .B(\mem[945][4] ), .S(n8421), .Z(n4163)
         );
  MUX2_X1 U23117 ( .A(n4163), .B(n4162), .S(n8333), .Z(n4164) );
  MUX2_X1 U23118 ( .A(n4164), .B(n4161), .S(n8265), .Z(n4165) );
  MUX2_X1 U23119 ( .A(n4165), .B(n4158), .S(n8209), .Z(n4166) );
  MUX2_X1 U23120 ( .A(\mem[942][4] ), .B(\mem[943][4] ), .S(n8422), .Z(n4167)
         );
  MUX2_X1 U23121 ( .A(\mem[940][4] ), .B(\mem[941][4] ), .S(n8417), .Z(n4168)
         );
  MUX2_X1 U23122 ( .A(n4168), .B(n4167), .S(n8334), .Z(n4169) );
  MUX2_X1 U23123 ( .A(\mem[938][4] ), .B(\mem[939][4] ), .S(n8418), .Z(n4170)
         );
  MUX2_X1 U23124 ( .A(\mem[936][4] ), .B(\mem[937][4] ), .S(n8419), .Z(n4171)
         );
  MUX2_X1 U23125 ( .A(n4171), .B(n4170), .S(n8329), .Z(n4172) );
  MUX2_X1 U23126 ( .A(n4172), .B(n4169), .S(n8232), .Z(n4173) );
  MUX2_X1 U23127 ( .A(\mem[934][4] ), .B(\mem[935][4] ), .S(n8375), .Z(n4174)
         );
  MUX2_X1 U23128 ( .A(\mem[932][4] ), .B(\mem[933][4] ), .S(n8397), .Z(n4175)
         );
  MUX2_X1 U23129 ( .A(n4175), .B(n4174), .S(n8330), .Z(n4176) );
  MUX2_X1 U23130 ( .A(\mem[930][4] ), .B(\mem[931][4] ), .S(n8468), .Z(n4177)
         );
  MUX2_X1 U23131 ( .A(\mem[928][4] ), .B(\mem[929][4] ), .S(n8440), .Z(n4178)
         );
  MUX2_X1 U23132 ( .A(n4178), .B(n4177), .S(n8331), .Z(n4179) );
  MUX2_X1 U23133 ( .A(n4179), .B(n4176), .S(n8225), .Z(n4180) );
  MUX2_X1 U23134 ( .A(n4180), .B(n4173), .S(n8210), .Z(n4181) );
  MUX2_X1 U23135 ( .A(n4181), .B(n4166), .S(n8187), .Z(n4182) );
  MUX2_X1 U23136 ( .A(\mem[926][4] ), .B(\mem[927][4] ), .S(n8526), .Z(n4183)
         );
  MUX2_X1 U23137 ( .A(\mem[924][4] ), .B(\mem[925][4] ), .S(n8362), .Z(n4184)
         );
  MUX2_X1 U23138 ( .A(n4184), .B(n4183), .S(n8338), .Z(n4185) );
  MUX2_X1 U23139 ( .A(\mem[922][4] ), .B(\mem[923][4] ), .S(n8366), .Z(n4186)
         );
  MUX2_X1 U23140 ( .A(\mem[920][4] ), .B(\mem[921][4] ), .S(n8395), .Z(n4187)
         );
  MUX2_X1 U23141 ( .A(n4187), .B(n4186), .S(n8339), .Z(n4188) );
  MUX2_X1 U23142 ( .A(n4188), .B(n4185), .S(n8223), .Z(n4189) );
  MUX2_X1 U23143 ( .A(\mem[918][4] ), .B(\mem[919][4] ), .S(n8394), .Z(n4190)
         );
  MUX2_X1 U23144 ( .A(\mem[916][4] ), .B(\mem[917][4] ), .S(n8510), .Z(n4191)
         );
  MUX2_X1 U23145 ( .A(n4191), .B(n4190), .S(n8340), .Z(n4192) );
  MUX2_X1 U23146 ( .A(\mem[914][4] ), .B(\mem[915][4] ), .S(n8483), .Z(n4193)
         );
  MUX2_X1 U23147 ( .A(\mem[912][4] ), .B(\mem[913][4] ), .S(n8409), .Z(n4194)
         );
  MUX2_X1 U23148 ( .A(n4194), .B(n4193), .S(n8335), .Z(n4195) );
  MUX2_X1 U23149 ( .A(n4195), .B(n4192), .S(n8262), .Z(n4196) );
  MUX2_X1 U23150 ( .A(n4196), .B(n4189), .S(n8206), .Z(n4197) );
  MUX2_X1 U23151 ( .A(\mem[910][4] ), .B(\mem[911][4] ), .S(n8467), .Z(n4198)
         );
  MUX2_X1 U23152 ( .A(\mem[908][4] ), .B(\mem[909][4] ), .S(n8474), .Z(n4199)
         );
  MUX2_X1 U23153 ( .A(n4199), .B(n4198), .S(n8304), .Z(n4200) );
  MUX2_X1 U23154 ( .A(\mem[906][4] ), .B(\mem[907][4] ), .S(n8475), .Z(n4201)
         );
  MUX2_X1 U23155 ( .A(\mem[904][4] ), .B(\mem[905][4] ), .S(n8476), .Z(n4202)
         );
  MUX2_X1 U23156 ( .A(n4202), .B(n4201), .S(n8299), .Z(n4203) );
  MUX2_X1 U23157 ( .A(n4203), .B(n4200), .S(n8223), .Z(n4204) );
  MUX2_X1 U23158 ( .A(\mem[902][4] ), .B(\mem[903][4] ), .S(n8471), .Z(n4205)
         );
  MUX2_X1 U23159 ( .A(\mem[900][4] ), .B(\mem[901][4] ), .S(n8472), .Z(n4206)
         );
  MUX2_X1 U23160 ( .A(n4206), .B(n4205), .S(n8300), .Z(n4207) );
  MUX2_X1 U23161 ( .A(\mem[898][4] ), .B(\mem[899][4] ), .S(n8473), .Z(n4208)
         );
  MUX2_X1 U23162 ( .A(\mem[896][4] ), .B(\mem[897][4] ), .S(n8480), .Z(n4209)
         );
  MUX2_X1 U23163 ( .A(n4209), .B(n4208), .S(n8301), .Z(n4210) );
  MUX2_X1 U23164 ( .A(n4210), .B(n4207), .S(n8222), .Z(n4211) );
  MUX2_X1 U23165 ( .A(n4211), .B(n4204), .S(n8215), .Z(n4212) );
  MUX2_X1 U23166 ( .A(n4212), .B(n4197), .S(n8187), .Z(n4213) );
  MUX2_X1 U23167 ( .A(n4213), .B(n4182), .S(n8182), .Z(n4214) );
  MUX2_X1 U23168 ( .A(n4214), .B(n4151), .S(N24), .Z(n4215) );
  MUX2_X1 U23169 ( .A(\mem[894][4] ), .B(\mem[895][4] ), .S(n8481), .Z(n4216)
         );
  MUX2_X1 U23170 ( .A(\mem[892][4] ), .B(\mem[893][4] ), .S(n8482), .Z(n4217)
         );
  MUX2_X1 U23171 ( .A(n4217), .B(n4216), .S(n8308), .Z(n4218) );
  MUX2_X1 U23172 ( .A(\mem[890][4] ), .B(\mem[891][4] ), .S(n8477), .Z(n4219)
         );
  MUX2_X1 U23173 ( .A(\mem[888][4] ), .B(\mem[889][4] ), .S(n8478), .Z(n4220)
         );
  MUX2_X1 U23174 ( .A(n4220), .B(n4219), .S(n8309), .Z(n4221) );
  MUX2_X1 U23175 ( .A(n4221), .B(n4218), .S(n8221), .Z(n4222) );
  MUX2_X1 U23176 ( .A(\mem[886][4] ), .B(\mem[887][4] ), .S(n8523), .Z(n4223)
         );
  MUX2_X1 U23177 ( .A(\mem[884][4] ), .B(\mem[885][4] ), .S(n8524), .Z(n4224)
         );
  MUX2_X1 U23178 ( .A(n4224), .B(n4223), .S(n8310), .Z(n4225) );
  MUX2_X1 U23179 ( .A(\mem[882][4] ), .B(\mem[883][4] ), .S(n8519), .Z(n4226)
         );
  MUX2_X1 U23180 ( .A(\mem[880][4] ), .B(\mem[881][4] ), .S(n8520), .Z(n4227)
         );
  MUX2_X1 U23181 ( .A(n4227), .B(n4226), .S(n8305), .Z(n4228) );
  MUX2_X1 U23182 ( .A(n4228), .B(n4225), .S(n8256), .Z(n4229) );
  MUX2_X1 U23183 ( .A(n4229), .B(n4222), .S(n8211), .Z(n4230) );
  MUX2_X1 U23184 ( .A(\mem[878][4] ), .B(\mem[879][4] ), .S(n8521), .Z(n4231)
         );
  MUX2_X1 U23185 ( .A(\mem[876][4] ), .B(\mem[877][4] ), .S(n8528), .Z(n4232)
         );
  MUX2_X1 U23186 ( .A(n4232), .B(n4231), .S(n8306), .Z(n4233) );
  MUX2_X1 U23187 ( .A(\mem[874][4] ), .B(\mem[875][4] ), .S(n8529), .Z(n4234)
         );
  MUX2_X1 U23188 ( .A(\mem[872][4] ), .B(\mem[873][4] ), .S(n8530), .Z(n4235)
         );
  MUX2_X1 U23189 ( .A(n4235), .B(n4234), .S(n8307), .Z(n4236) );
  MUX2_X1 U23190 ( .A(n4236), .B(n4233), .S(n8224), .Z(n4237) );
  MUX2_X1 U23191 ( .A(\mem[870][4] ), .B(\mem[871][4] ), .S(n8525), .Z(n4238)
         );
  MUX2_X1 U23192 ( .A(\mem[868][4] ), .B(\mem[869][4] ), .S(n8526), .Z(n4239)
         );
  MUX2_X1 U23193 ( .A(n4239), .B(n4238), .S(n8314), .Z(n4240) );
  MUX2_X1 U23194 ( .A(\mem[866][4] ), .B(\mem[867][4] ), .S(n8527), .Z(n4241)
         );
  MUX2_X1 U23195 ( .A(\mem[864][4] ), .B(\mem[865][4] ), .S(n8534), .Z(n4242)
         );
  MUX2_X1 U23196 ( .A(n4242), .B(n4241), .S(n8315), .Z(n4243) );
  MUX2_X1 U23197 ( .A(n4243), .B(n4240), .S(n8259), .Z(n4244) );
  MUX2_X1 U23198 ( .A(n4244), .B(n4237), .S(n8216), .Z(n4245) );
  MUX2_X1 U23199 ( .A(n4245), .B(n4230), .S(n8187), .Z(n4246) );
  MUX2_X1 U23200 ( .A(\mem[862][4] ), .B(\mem[863][4] ), .S(n8505), .Z(n4247)
         );
  MUX2_X1 U23201 ( .A(\mem[860][4] ), .B(\mem[861][4] ), .S(n8506), .Z(n4248)
         );
  MUX2_X1 U23202 ( .A(n4248), .B(n4247), .S(n8288), .Z(n4249) );
  MUX2_X1 U23203 ( .A(\mem[858][4] ), .B(\mem[859][4] ), .S(n8501), .Z(n4250)
         );
  MUX2_X1 U23204 ( .A(\mem[856][4] ), .B(\mem[857][4] ), .S(n8502), .Z(n4251)
         );
  MUX2_X1 U23205 ( .A(n4251), .B(n4250), .S(n8276), .Z(n4252) );
  MUX2_X1 U23206 ( .A(n4252), .B(n4249), .S(n8222), .Z(n4253) );
  MUX2_X1 U23207 ( .A(\mem[854][4] ), .B(\mem[855][4] ), .S(n8503), .Z(n4254)
         );
  MUX2_X1 U23208 ( .A(\mem[852][4] ), .B(\mem[853][4] ), .S(n8510), .Z(n4255)
         );
  MUX2_X1 U23209 ( .A(n4255), .B(n4254), .S(n8284), .Z(n4256) );
  MUX2_X1 U23210 ( .A(\mem[850][4] ), .B(\mem[851][4] ), .S(n8511), .Z(n4257)
         );
  MUX2_X1 U23211 ( .A(\mem[848][4] ), .B(\mem[849][4] ), .S(n8512), .Z(n4258)
         );
  MUX2_X1 U23212 ( .A(n4258), .B(n4257), .S(n8285), .Z(n4259) );
  MUX2_X1 U23213 ( .A(n4259), .B(n4256), .S(n8264), .Z(n4260) );
  MUX2_X1 U23214 ( .A(n4260), .B(n4253), .S(n8217), .Z(n4261) );
  MUX2_X1 U23215 ( .A(\mem[846][4] ), .B(\mem[847][4] ), .S(n8507), .Z(n4262)
         );
  MUX2_X1 U23216 ( .A(\mem[844][4] ), .B(\mem[845][4] ), .S(n8508), .Z(n4263)
         );
  MUX2_X1 U23217 ( .A(n4263), .B(n4262), .S(n8286), .Z(n4264) );
  MUX2_X1 U23218 ( .A(\mem[842][4] ), .B(\mem[843][4] ), .S(n8509), .Z(n4265)
         );
  MUX2_X1 U23219 ( .A(\mem[840][4] ), .B(\mem[841][4] ), .S(n8516), .Z(n4266)
         );
  MUX2_X1 U23220 ( .A(n4266), .B(n4265), .S(n8290), .Z(n4267) );
  MUX2_X1 U23221 ( .A(n4267), .B(n4264), .S(n8225), .Z(n4268) );
  MUX2_X1 U23222 ( .A(\mem[838][4] ), .B(\mem[839][4] ), .S(n8486), .Z(n4269)
         );
  MUX2_X1 U23223 ( .A(\mem[836][4] ), .B(\mem[837][4] ), .S(n8487), .Z(n4270)
         );
  MUX2_X1 U23224 ( .A(n4270), .B(n4269), .S(n8291), .Z(n4271) );
  MUX2_X1 U23225 ( .A(\mem[834][4] ), .B(\mem[835][4] ), .S(n8488), .Z(n4272)
         );
  MUX2_X1 U23226 ( .A(\mem[832][4] ), .B(\mem[833][4] ), .S(n8483), .Z(n4273)
         );
  MUX2_X1 U23227 ( .A(n4273), .B(n4272), .S(n8292), .Z(n4274) );
  MUX2_X1 U23228 ( .A(n4274), .B(n4271), .S(n8221), .Z(n4275) );
  MUX2_X1 U23229 ( .A(n4275), .B(n4268), .S(n8218), .Z(n4276) );
  MUX2_X1 U23230 ( .A(n4276), .B(n4261), .S(n8187), .Z(n4277) );
  MUX2_X1 U23231 ( .A(n4277), .B(n4246), .S(n8183), .Z(n4278) );
  MUX2_X1 U23232 ( .A(\mem[830][4] ), .B(\mem[831][4] ), .S(n8484), .Z(n4279)
         );
  MUX2_X1 U23233 ( .A(\mem[828][4] ), .B(\mem[829][4] ), .S(n8485), .Z(n4280)
         );
  MUX2_X1 U23234 ( .A(n4280), .B(n4279), .S(n8287), .Z(n4281) );
  MUX2_X1 U23235 ( .A(\mem[826][4] ), .B(\mem[827][4] ), .S(n8492), .Z(n4282)
         );
  MUX2_X1 U23236 ( .A(\mem[824][4] ), .B(\mem[825][4] ), .S(n8493), .Z(n4283)
         );
  MUX2_X1 U23237 ( .A(n4283), .B(n4282), .S(n8288), .Z(n4284) );
  MUX2_X1 U23238 ( .A(n4284), .B(n4281), .S(n8243), .Z(n4285) );
  MUX2_X1 U23239 ( .A(\mem[822][4] ), .B(\mem[823][4] ), .S(n8494), .Z(n4286)
         );
  MUX2_X1 U23240 ( .A(\mem[820][4] ), .B(\mem[821][4] ), .S(n8489), .Z(n4287)
         );
  MUX2_X1 U23241 ( .A(n4287), .B(n4286), .S(n8289), .Z(n4288) );
  MUX2_X1 U23242 ( .A(\mem[818][4] ), .B(\mem[819][4] ), .S(n8490), .Z(n4289)
         );
  MUX2_X1 U23243 ( .A(\mem[816][4] ), .B(\mem[817][4] ), .S(n8491), .Z(n4290)
         );
  MUX2_X1 U23244 ( .A(n4290), .B(n4289), .S(n8296), .Z(n4291) );
  MUX2_X1 U23245 ( .A(n4291), .B(n4288), .S(n8257), .Z(n4292) );
  MUX2_X1 U23246 ( .A(n4292), .B(n4285), .S(N21), .Z(n4293) );
  MUX2_X1 U23247 ( .A(\mem[814][4] ), .B(\mem[815][4] ), .S(n8446), .Z(n4294)
         );
  MUX2_X1 U23248 ( .A(\mem[812][4] ), .B(\mem[813][4] ), .S(n8519), .Z(n4295)
         );
  MUX2_X1 U23249 ( .A(n4295), .B(n4294), .S(n8330), .Z(n4296) );
  MUX2_X1 U23250 ( .A(\mem[810][4] ), .B(\mem[811][4] ), .S(n8443), .Z(n4297)
         );
  MUX2_X1 U23251 ( .A(\mem[808][4] ), .B(\mem[809][4] ), .S(n8515), .Z(n4298)
         );
  MUX2_X1 U23252 ( .A(n4298), .B(n4297), .S(n8331), .Z(n4299) );
  MUX2_X1 U23253 ( .A(n4299), .B(n4296), .S(n8258), .Z(n4300) );
  MUX2_X1 U23254 ( .A(\mem[806][4] ), .B(\mem[807][4] ), .S(n8498), .Z(n4301)
         );
  MUX2_X1 U23255 ( .A(\mem[804][4] ), .B(\mem[805][4] ), .S(n8385), .Z(n4302)
         );
  MUX2_X1 U23256 ( .A(n4302), .B(n4301), .S(n8338), .Z(n4303) );
  MUX2_X1 U23257 ( .A(\mem[802][4] ), .B(\mem[803][4] ), .S(n8384), .Z(n4304)
         );
  MUX2_X1 U23258 ( .A(\mem[800][4] ), .B(\mem[801][4] ), .S(n8383), .Z(n4305)
         );
  MUX2_X1 U23259 ( .A(n4305), .B(n4304), .S(n8339), .Z(n4306) );
  MUX2_X1 U23260 ( .A(n4306), .B(n4303), .S(n8224), .Z(n4307) );
  MUX2_X1 U23261 ( .A(n4307), .B(n4300), .S(n8216), .Z(n4308) );
  MUX2_X1 U23262 ( .A(n4308), .B(n4293), .S(n8187), .Z(n4309) );
  MUX2_X1 U23263 ( .A(\mem[798][4] ), .B(\mem[799][4] ), .S(n8382), .Z(n4310)
         );
  MUX2_X1 U23264 ( .A(\mem[796][4] ), .B(\mem[797][4] ), .S(n8381), .Z(n4311)
         );
  MUX2_X1 U23265 ( .A(n4311), .B(n4310), .S(n8340), .Z(n4312) );
  MUX2_X1 U23266 ( .A(\mem[794][4] ), .B(\mem[795][4] ), .S(n8380), .Z(n4313)
         );
  MUX2_X1 U23267 ( .A(\mem[792][4] ), .B(\mem[793][4] ), .S(n8379), .Z(n4314)
         );
  MUX2_X1 U23268 ( .A(n4314), .B(n4313), .S(n8335), .Z(n4315) );
  MUX2_X1 U23269 ( .A(n4315), .B(n4312), .S(n8223), .Z(n4316) );
  MUX2_X1 U23270 ( .A(\mem[790][4] ), .B(\mem[791][4] ), .S(n8465), .Z(n4317)
         );
  MUX2_X1 U23271 ( .A(\mem[788][4] ), .B(\mem[789][4] ), .S(n8466), .Z(n4318)
         );
  MUX2_X1 U23272 ( .A(n4318), .B(n4317), .S(n8336), .Z(n4319) );
  MUX2_X1 U23273 ( .A(\mem[786][4] ), .B(\mem[787][4] ), .S(n8467), .Z(n4320)
         );
  MUX2_X1 U23274 ( .A(\mem[784][4] ), .B(\mem[785][4] ), .S(n8474), .Z(n4321)
         );
  MUX2_X1 U23275 ( .A(n4321), .B(n4320), .S(n8337), .Z(n4322) );
  MUX2_X1 U23276 ( .A(n4322), .B(n4319), .S(n8224), .Z(n4323) );
  MUX2_X1 U23277 ( .A(n4323), .B(n4316), .S(n8200), .Z(n4324) );
  MUX2_X1 U23278 ( .A(\mem[782][4] ), .B(\mem[783][4] ), .S(n8476), .Z(n4325)
         );
  MUX2_X1 U23279 ( .A(\mem[780][4] ), .B(\mem[781][4] ), .S(n8471), .Z(n4326)
         );
  MUX2_X1 U23280 ( .A(n4326), .B(n4325), .S(n8344), .Z(n4327) );
  MUX2_X1 U23281 ( .A(\mem[778][4] ), .B(\mem[779][4] ), .S(n8472), .Z(n4328)
         );
  MUX2_X1 U23282 ( .A(\mem[776][4] ), .B(\mem[777][4] ), .S(n8473), .Z(n4329)
         );
  MUX2_X1 U23283 ( .A(n4329), .B(n4328), .S(n8345), .Z(n4330) );
  MUX2_X1 U23284 ( .A(n4330), .B(n4327), .S(n8264), .Z(n4331) );
  MUX2_X1 U23285 ( .A(\mem[774][4] ), .B(\mem[775][4] ), .S(n8480), .Z(n4332)
         );
  MUX2_X1 U23286 ( .A(\mem[772][4] ), .B(\mem[773][4] ), .S(n8481), .Z(n4333)
         );
  MUX2_X1 U23287 ( .A(n4333), .B(n4332), .S(n8346), .Z(n4334) );
  MUX2_X1 U23288 ( .A(\mem[770][4] ), .B(\mem[771][4] ), .S(n8482), .Z(n4335)
         );
  MUX2_X1 U23289 ( .A(\mem[768][4] ), .B(\mem[769][4] ), .S(n8477), .Z(n4336)
         );
  MUX2_X1 U23290 ( .A(n4336), .B(n4335), .S(n8341), .Z(n4337) );
  MUX2_X1 U23291 ( .A(n4337), .B(n4334), .S(n8257), .Z(n4338) );
  MUX2_X1 U23292 ( .A(n4338), .B(n4331), .S(n8199), .Z(n4339) );
  MUX2_X1 U23293 ( .A(n4339), .B(n4324), .S(n8187), .Z(n4340) );
  MUX2_X1 U23294 ( .A(n4340), .B(n4309), .S(n8184), .Z(n4341) );
  MUX2_X1 U23295 ( .A(n4341), .B(n4278), .S(n8179), .Z(n4342) );
  MUX2_X1 U23296 ( .A(n4342), .B(n4215), .S(n8177), .Z(n4343) );
  MUX2_X1 U23297 ( .A(\mem[766][4] ), .B(\mem[767][4] ), .S(n8447), .Z(n4344)
         );
  MUX2_X1 U23298 ( .A(\mem[764][4] ), .B(\mem[765][4] ), .S(n8448), .Z(n4345)
         );
  MUX2_X1 U23299 ( .A(n4345), .B(n4344), .S(n8297), .Z(n4346) );
  MUX2_X1 U23300 ( .A(\mem[762][4] ), .B(\mem[763][4] ), .S(n8449), .Z(n4347)
         );
  MUX2_X1 U23301 ( .A(\mem[760][4] ), .B(\mem[761][4] ), .S(n8456), .Z(n4348)
         );
  MUX2_X1 U23302 ( .A(n4348), .B(n4347), .S(n8298), .Z(n4349) );
  MUX2_X1 U23303 ( .A(n4349), .B(n4346), .S(n8251), .Z(n4350) );
  MUX2_X1 U23304 ( .A(\mem[758][4] ), .B(\mem[759][4] ), .S(n8457), .Z(n4351)
         );
  MUX2_X1 U23305 ( .A(\mem[756][4] ), .B(\mem[757][4] ), .S(n8458), .Z(n4352)
         );
  MUX2_X1 U23306 ( .A(n4352), .B(n4351), .S(n8293), .Z(n4353) );
  MUX2_X1 U23307 ( .A(\mem[754][4] ), .B(\mem[755][4] ), .S(n8453), .Z(n4354)
         );
  MUX2_X1 U23308 ( .A(\mem[752][4] ), .B(\mem[753][4] ), .S(n8454), .Z(n4355)
         );
  MUX2_X1 U23309 ( .A(n4355), .B(n4354), .S(n8294), .Z(n4356) );
  MUX2_X1 U23310 ( .A(n4356), .B(n4353), .S(n8240), .Z(n4357) );
  MUX2_X1 U23311 ( .A(n4357), .B(n4350), .S(n8201), .Z(n4358) );
  MUX2_X1 U23312 ( .A(\mem[750][4] ), .B(\mem[751][4] ), .S(n8455), .Z(n4359)
         );
  MUX2_X1 U23313 ( .A(\mem[748][4] ), .B(\mem[749][4] ), .S(n8462), .Z(n4360)
         );
  MUX2_X1 U23314 ( .A(n4360), .B(n4359), .S(n8295), .Z(n4361) );
  MUX2_X1 U23315 ( .A(\mem[746][4] ), .B(\mem[747][4] ), .S(n8463), .Z(n4362)
         );
  MUX2_X1 U23316 ( .A(\mem[744][4] ), .B(\mem[745][4] ), .S(n8464), .Z(n4363)
         );
  MUX2_X1 U23317 ( .A(n4363), .B(n4362), .S(n8302), .Z(n4364) );
  MUX2_X1 U23318 ( .A(n4364), .B(n4361), .S(n8265), .Z(n4365) );
  MUX2_X1 U23319 ( .A(\mem[742][4] ), .B(\mem[743][4] ), .S(n8473), .Z(n4366)
         );
  MUX2_X1 U23320 ( .A(\mem[740][4] ), .B(\mem[741][4] ), .S(n8539), .Z(n4367)
         );
  MUX2_X1 U23321 ( .A(n4367), .B(n4366), .S(n8303), .Z(n4368) );
  MUX2_X1 U23322 ( .A(\mem[738][4] ), .B(\mem[739][4] ), .S(n8384), .Z(n4369)
         );
  MUX2_X1 U23323 ( .A(\mem[736][4] ), .B(\mem[737][4] ), .S(n8396), .Z(n4370)
         );
  MUX2_X1 U23324 ( .A(n4370), .B(n4369), .S(n8304), .Z(n4371) );
  MUX2_X1 U23325 ( .A(n4371), .B(n4368), .S(n8263), .Z(n4372) );
  MUX2_X1 U23326 ( .A(n4372), .B(n4365), .S(n8201), .Z(n4373) );
  MUX2_X1 U23327 ( .A(n4373), .B(n4358), .S(n8188), .Z(n4374) );
  MUX2_X1 U23328 ( .A(\mem[734][4] ), .B(\mem[735][4] ), .S(n8461), .Z(n4375)
         );
  MUX2_X1 U23329 ( .A(\mem[732][4] ), .B(\mem[733][4] ), .S(n8439), .Z(n4376)
         );
  MUX2_X1 U23330 ( .A(n4376), .B(n4375), .S(n8299), .Z(n4377) );
  MUX2_X1 U23331 ( .A(\mem[730][4] ), .B(\mem[731][4] ), .S(n8525), .Z(n4378)
         );
  MUX2_X1 U23332 ( .A(\mem[728][4] ), .B(\mem[729][4] ), .S(n8361), .Z(n4379)
         );
  MUX2_X1 U23333 ( .A(n4379), .B(n4378), .S(n8300), .Z(n4380) );
  MUX2_X1 U23334 ( .A(n4380), .B(n4377), .S(n8265), .Z(n4381) );
  MUX2_X1 U23335 ( .A(\mem[726][4] ), .B(\mem[727][4] ), .S(n8370), .Z(n4382)
         );
  MUX2_X1 U23336 ( .A(\mem[724][4] ), .B(\mem[725][4] ), .S(n8400), .Z(n4383)
         );
  MUX2_X1 U23337 ( .A(n4383), .B(n4382), .S(n8301), .Z(n4384) );
  MUX2_X1 U23338 ( .A(\mem[722][4] ), .B(\mem[723][4] ), .S(n8393), .Z(n4385)
         );
  MUX2_X1 U23339 ( .A(\mem[720][4] ), .B(\mem[721][4] ), .S(n8503), .Z(n4386)
         );
  MUX2_X1 U23340 ( .A(n4386), .B(n4385), .S(n8326), .Z(n4387) );
  MUX2_X1 U23341 ( .A(n4387), .B(n4384), .S(n8264), .Z(n4388) );
  MUX2_X1 U23342 ( .A(n4388), .B(n4381), .S(n8201), .Z(n4389) );
  MUX2_X1 U23343 ( .A(\mem[718][4] ), .B(\mem[719][4] ), .S(n8361), .Z(n4390)
         );
  MUX2_X1 U23344 ( .A(\mem[716][4] ), .B(\mem[717][4] ), .S(n8539), .Z(n4391)
         );
  MUX2_X1 U23345 ( .A(n4391), .B(n4390), .S(n8309), .Z(n4392) );
  MUX2_X1 U23346 ( .A(\mem[714][4] ), .B(\mem[715][4] ), .S(n8362), .Z(n4393)
         );
  MUX2_X1 U23347 ( .A(\mem[712][4] ), .B(\mem[713][4] ), .S(n8363), .Z(n4394)
         );
  MUX2_X1 U23348 ( .A(n4394), .B(n4393), .S(n8310), .Z(n4395) );
  MUX2_X1 U23349 ( .A(n4395), .B(n4392), .S(n8252), .Z(n4396) );
  MUX2_X1 U23350 ( .A(\mem[710][4] ), .B(\mem[711][4] ), .S(n8364), .Z(n4397)
         );
  MUX2_X1 U23351 ( .A(\mem[708][4] ), .B(\mem[709][4] ), .S(n8479), .Z(n4398)
         );
  MUX2_X1 U23352 ( .A(n4398), .B(n4397), .S(n8305), .Z(n4399) );
  MUX2_X1 U23353 ( .A(\mem[706][4] ), .B(\mem[707][4] ), .S(n8488), .Z(n4400)
         );
  MUX2_X1 U23354 ( .A(\mem[704][4] ), .B(\mem[705][4] ), .S(n8447), .Z(n4401)
         );
  MUX2_X1 U23355 ( .A(n4401), .B(n4400), .S(n8306), .Z(n4402) );
  MUX2_X1 U23356 ( .A(n4402), .B(n4399), .S(n8230), .Z(n4403) );
  MUX2_X1 U23357 ( .A(n4403), .B(n4396), .S(n8201), .Z(n4404) );
  MUX2_X1 U23358 ( .A(n4404), .B(n4389), .S(n8188), .Z(n4405) );
  MUX2_X1 U23359 ( .A(n4405), .B(n4374), .S(n8184), .Z(n4406) );
  MUX2_X1 U23360 ( .A(\mem[702][4] ), .B(\mem[703][4] ), .S(n8448), .Z(n4407)
         );
  MUX2_X1 U23361 ( .A(\mem[700][4] ), .B(\mem[701][4] ), .S(n8358), .Z(n4408)
         );
  MUX2_X1 U23362 ( .A(n4408), .B(n4407), .S(n8307), .Z(n4409) );
  MUX2_X1 U23363 ( .A(\mem[698][4] ), .B(\mem[699][4] ), .S(n8514), .Z(n4410)
         );
  MUX2_X1 U23364 ( .A(\mem[696][4] ), .B(\mem[697][4] ), .S(n8456), .Z(n4411)
         );
  MUX2_X1 U23365 ( .A(n4411), .B(n4410), .S(n8314), .Z(n4412) );
  MUX2_X1 U23366 ( .A(n4412), .B(n4409), .S(n8264), .Z(n4413) );
  MUX2_X1 U23367 ( .A(\mem[694][4] ), .B(\mem[695][4] ), .S(n8372), .Z(n4414)
         );
  MUX2_X1 U23368 ( .A(\mem[692][4] ), .B(\mem[693][4] ), .S(n8371), .Z(n4415)
         );
  MUX2_X1 U23369 ( .A(n4415), .B(n4414), .S(n8315), .Z(n4416) );
  MUX2_X1 U23370 ( .A(\mem[690][4] ), .B(\mem[691][4] ), .S(n8370), .Z(n4417)
         );
  MUX2_X1 U23371 ( .A(\mem[688][4] ), .B(\mem[689][4] ), .S(n8369), .Z(n4418)
         );
  MUX2_X1 U23372 ( .A(n4418), .B(n4417), .S(n8316), .Z(n4419) );
  MUX2_X1 U23373 ( .A(n4419), .B(n4416), .S(n8221), .Z(n4420) );
  MUX2_X1 U23374 ( .A(n4420), .B(n4413), .S(n8201), .Z(n4421) );
  MUX2_X1 U23375 ( .A(\mem[686][4] ), .B(\mem[687][4] ), .S(n8368), .Z(n4422)
         );
  MUX2_X1 U23376 ( .A(\mem[684][4] ), .B(\mem[685][4] ), .S(n8367), .Z(n4423)
         );
  MUX2_X1 U23377 ( .A(n4423), .B(n4422), .S(n8311), .Z(n4424) );
  MUX2_X1 U23378 ( .A(\mem[682][4] ), .B(\mem[683][4] ), .S(n8366), .Z(n4425)
         );
  MUX2_X1 U23379 ( .A(\mem[680][4] ), .B(\mem[681][4] ), .S(n8365), .Z(n4426)
         );
  MUX2_X1 U23380 ( .A(n4426), .B(n4425), .S(n8312), .Z(n4427) );
  MUX2_X1 U23381 ( .A(n4427), .B(n4424), .S(n8263), .Z(n4428) );
  MUX2_X1 U23382 ( .A(\mem[678][4] ), .B(\mem[679][4] ), .S(n8387), .Z(n4429)
         );
  MUX2_X1 U23383 ( .A(\mem[676][4] ), .B(\mem[677][4] ), .S(n8386), .Z(n4430)
         );
  MUX2_X1 U23384 ( .A(n4430), .B(n4429), .S(n8313), .Z(n4431) );
  MUX2_X1 U23385 ( .A(\mem[674][4] ), .B(\mem[675][4] ), .S(n8445), .Z(n4432)
         );
  MUX2_X1 U23386 ( .A(\mem[672][4] ), .B(\mem[673][4] ), .S(n8357), .Z(n4433)
         );
  MUX2_X1 U23387 ( .A(n4433), .B(n4432), .S(n8320), .Z(n4434) );
  MUX2_X1 U23388 ( .A(n4434), .B(n4431), .S(n8265), .Z(n4435) );
  MUX2_X1 U23389 ( .A(n4435), .B(n4428), .S(n8201), .Z(n4436) );
  MUX2_X1 U23390 ( .A(n4436), .B(n4421), .S(n8188), .Z(n4437) );
  MUX2_X1 U23391 ( .A(\mem[670][4] ), .B(\mem[671][4] ), .S(n8382), .Z(n4438)
         );
  MUX2_X1 U23392 ( .A(\mem[668][4] ), .B(\mem[669][4] ), .S(n8381), .Z(n4439)
         );
  MUX2_X1 U23393 ( .A(n4439), .B(n4438), .S(n8283), .Z(n4440) );
  MUX2_X1 U23394 ( .A(\mem[666][4] ), .B(\mem[667][4] ), .S(n8449), .Z(n4441)
         );
  MUX2_X1 U23395 ( .A(\mem[664][4] ), .B(\mem[665][4] ), .S(n8359), .Z(n4442)
         );
  MUX2_X1 U23396 ( .A(n4442), .B(n4441), .S(n8283), .Z(n4443) );
  MUX2_X1 U23397 ( .A(n4443), .B(n4440), .S(n8220), .Z(n4444) );
  MUX2_X1 U23398 ( .A(\mem[662][4] ), .B(\mem[663][4] ), .S(n8538), .Z(n4445)
         );
  MUX2_X1 U23399 ( .A(\mem[660][4] ), .B(\mem[661][4] ), .S(n8539), .Z(n4446)
         );
  MUX2_X1 U23400 ( .A(n4446), .B(n4445), .S(n8283), .Z(n4447) );
  MUX2_X1 U23401 ( .A(\mem[658][4] ), .B(\mem[659][4] ), .S(n8362), .Z(n4448)
         );
  MUX2_X1 U23402 ( .A(\mem[656][4] ), .B(\mem[657][4] ), .S(n8363), .Z(n4449)
         );
  MUX2_X1 U23403 ( .A(n4449), .B(n4448), .S(n8283), .Z(n4450) );
  MUX2_X1 U23404 ( .A(n4450), .B(n4447), .S(n8236), .Z(n4451) );
  MUX2_X1 U23405 ( .A(n4451), .B(n4444), .S(n8201), .Z(n4452) );
  MUX2_X1 U23406 ( .A(\mem[654][4] ), .B(\mem[655][4] ), .S(n8364), .Z(n4453)
         );
  MUX2_X1 U23407 ( .A(\mem[652][4] ), .B(\mem[653][4] ), .S(n8357), .Z(n4454)
         );
  MUX2_X1 U23408 ( .A(n4454), .B(n4453), .S(n8283), .Z(n4455) );
  MUX2_X1 U23409 ( .A(\mem[650][4] ), .B(\mem[651][4] ), .S(n8360), .Z(n4456)
         );
  MUX2_X1 U23410 ( .A(\mem[648][4] ), .B(\mem[649][4] ), .S(n8459), .Z(n4457)
         );
  MUX2_X1 U23411 ( .A(n4457), .B(n4456), .S(n8283), .Z(n4458) );
  MUX2_X1 U23412 ( .A(n4458), .B(n4455), .S(n8237), .Z(n4459) );
  MUX2_X1 U23413 ( .A(\mem[646][4] ), .B(\mem[647][4] ), .S(n8366), .Z(n4460)
         );
  MUX2_X1 U23414 ( .A(\mem[644][4] ), .B(\mem[645][4] ), .S(n8387), .Z(n4461)
         );
  MUX2_X1 U23415 ( .A(n4461), .B(n4460), .S(n8283), .Z(n4462) );
  MUX2_X1 U23416 ( .A(\mem[642][4] ), .B(\mem[643][4] ), .S(n8372), .Z(n4463)
         );
  MUX2_X1 U23417 ( .A(\mem[640][4] ), .B(\mem[641][4] ), .S(n8371), .Z(n4464)
         );
  MUX2_X1 U23418 ( .A(n4464), .B(n4463), .S(n8283), .Z(n4465) );
  MUX2_X1 U23419 ( .A(n4465), .B(n4462), .S(n8232), .Z(n4466) );
  MUX2_X1 U23420 ( .A(n4466), .B(n4459), .S(n8201), .Z(n4467) );
  MUX2_X1 U23421 ( .A(n4467), .B(n4452), .S(n8188), .Z(n4468) );
  MUX2_X1 U23422 ( .A(n4468), .B(n4437), .S(N23), .Z(n4469) );
  MUX2_X1 U23423 ( .A(n4469), .B(n4406), .S(n8178), .Z(n4470) );
  MUX2_X1 U23424 ( .A(\mem[638][4] ), .B(\mem[639][4] ), .S(n8369), .Z(n4471)
         );
  MUX2_X1 U23425 ( .A(\mem[636][4] ), .B(\mem[637][4] ), .S(n8368), .Z(n4472)
         );
  MUX2_X1 U23426 ( .A(n4472), .B(n4471), .S(n8283), .Z(n4473) );
  MUX2_X1 U23427 ( .A(\mem[634][4] ), .B(\mem[635][4] ), .S(n8365), .Z(n4474)
         );
  MUX2_X1 U23428 ( .A(\mem[632][4] ), .B(\mem[633][4] ), .S(n8386), .Z(n4475)
         );
  MUX2_X1 U23429 ( .A(n4475), .B(n4474), .S(n8283), .Z(n4476) );
  MUX2_X1 U23430 ( .A(n4476), .B(n4473), .S(n8233), .Z(n4477) );
  MUX2_X1 U23431 ( .A(\mem[630][4] ), .B(\mem[631][4] ), .S(n8379), .Z(n4478)
         );
  MUX2_X1 U23432 ( .A(\mem[628][4] ), .B(\mem[629][4] ), .S(n8378), .Z(n4479)
         );
  MUX2_X1 U23433 ( .A(n4479), .B(n4478), .S(n8283), .Z(n4480) );
  MUX2_X1 U23434 ( .A(\mem[626][4] ), .B(\mem[627][4] ), .S(n8377), .Z(n4481)
         );
  MUX2_X1 U23435 ( .A(\mem[624][4] ), .B(\mem[625][4] ), .S(n8442), .Z(n4482)
         );
  MUX2_X1 U23436 ( .A(n4482), .B(n4481), .S(n8283), .Z(n4483) );
  MUX2_X1 U23437 ( .A(n4483), .B(n4480), .S(n8234), .Z(n4484) );
  MUX2_X1 U23438 ( .A(n4484), .B(n4477), .S(n8201), .Z(n4485) );
  MUX2_X1 U23439 ( .A(\mem[622][4] ), .B(\mem[623][4] ), .S(n8391), .Z(n4486)
         );
  MUX2_X1 U23440 ( .A(\mem[620][4] ), .B(\mem[621][4] ), .S(n8392), .Z(n4487)
         );
  MUX2_X1 U23441 ( .A(n4487), .B(n4486), .S(n8322), .Z(n4488) );
  MUX2_X1 U23442 ( .A(\mem[618][4] ), .B(\mem[619][4] ), .S(n8389), .Z(n4489)
         );
  MUX2_X1 U23443 ( .A(\mem[616][4] ), .B(\mem[617][4] ), .S(n8441), .Z(n4490)
         );
  MUX2_X1 U23444 ( .A(n4490), .B(n4489), .S(n8317), .Z(n4491) );
  MUX2_X1 U23445 ( .A(n4491), .B(n4488), .S(n8241), .Z(n4492) );
  MUX2_X1 U23446 ( .A(\mem[614][4] ), .B(\mem[615][4] ), .S(n8457), .Z(n4493)
         );
  MUX2_X1 U23447 ( .A(\mem[612][4] ), .B(\mem[613][4] ), .S(N18), .Z(n4494) );
  MUX2_X1 U23448 ( .A(n4494), .B(n4493), .S(n8318), .Z(n4495) );
  MUX2_X1 U23449 ( .A(\mem[610][4] ), .B(\mem[611][4] ), .S(n8446), .Z(n4496)
         );
  MUX2_X1 U23450 ( .A(\mem[608][4] ), .B(\mem[609][4] ), .S(n8400), .Z(n4497)
         );
  MUX2_X1 U23451 ( .A(n4497), .B(n4496), .S(n8319), .Z(n4498) );
  MUX2_X1 U23452 ( .A(n4498), .B(n4495), .S(n8242), .Z(n4499) );
  MUX2_X1 U23453 ( .A(n4499), .B(n4492), .S(n8201), .Z(n4500) );
  MUX2_X1 U23454 ( .A(n4500), .B(n4485), .S(n8188), .Z(n4501) );
  MUX2_X1 U23455 ( .A(\mem[606][4] ), .B(\mem[607][4] ), .S(n8395), .Z(n4502)
         );
  MUX2_X1 U23456 ( .A(\mem[604][4] ), .B(\mem[605][4] ), .S(n8396), .Z(n4503)
         );
  MUX2_X1 U23457 ( .A(n4503), .B(n4502), .S(N19), .Z(n4504) );
  MUX2_X1 U23458 ( .A(\mem[602][4] ), .B(\mem[603][4] ), .S(n8397), .Z(n4505)
         );
  MUX2_X1 U23459 ( .A(\mem[600][4] ), .B(\mem[601][4] ), .S(n8459), .Z(n4506)
         );
  MUX2_X1 U23460 ( .A(n4506), .B(n4505), .S(n8356), .Z(n4507) );
  MUX2_X1 U23461 ( .A(n4507), .B(n4504), .S(n8243), .Z(n4508) );
  MUX2_X1 U23462 ( .A(\mem[598][4] ), .B(\mem[599][4] ), .S(n8529), .Z(n4509)
         );
  MUX2_X1 U23463 ( .A(\mem[596][4] ), .B(\mem[597][4] ), .S(n8530), .Z(n4510)
         );
  MUX2_X1 U23464 ( .A(n4510), .B(n4509), .S(n8270), .Z(n4511) );
  MUX2_X1 U23465 ( .A(\mem[594][4] ), .B(\mem[595][4] ), .S(n8525), .Z(n4512)
         );
  MUX2_X1 U23466 ( .A(\mem[592][4] ), .B(\mem[593][4] ), .S(n8526), .Z(n4513)
         );
  MUX2_X1 U23467 ( .A(n4513), .B(n4512), .S(n8321), .Z(n4514) );
  MUX2_X1 U23468 ( .A(n4514), .B(n4511), .S(n8238), .Z(n4515) );
  MUX2_X1 U23469 ( .A(n4515), .B(n4508), .S(n8201), .Z(n4516) );
  MUX2_X1 U23470 ( .A(\mem[590][4] ), .B(\mem[591][4] ), .S(n8527), .Z(n4517)
         );
  MUX2_X1 U23471 ( .A(\mem[588][4] ), .B(\mem[589][4] ), .S(n8534), .Z(n4518)
         );
  MUX2_X1 U23472 ( .A(n4518), .B(n4517), .S(n8326), .Z(n4519) );
  MUX2_X1 U23473 ( .A(\mem[586][4] ), .B(\mem[587][4] ), .S(n8535), .Z(n4520)
         );
  MUX2_X1 U23474 ( .A(\mem[584][4] ), .B(\mem[585][4] ), .S(n8536), .Z(n4521)
         );
  MUX2_X1 U23475 ( .A(n4521), .B(n4520), .S(n8281), .Z(n4522) );
  MUX2_X1 U23476 ( .A(n4522), .B(n4519), .S(n8239), .Z(n4523) );
  MUX2_X1 U23477 ( .A(\mem[582][4] ), .B(\mem[583][4] ), .S(n8531), .Z(n4524)
         );
  MUX2_X1 U23478 ( .A(\mem[580][4] ), .B(\mem[581][4] ), .S(n8532), .Z(n4525)
         );
  MUX2_X1 U23479 ( .A(n4525), .B(n4524), .S(n8275), .Z(n4526) );
  MUX2_X1 U23480 ( .A(\mem[578][4] ), .B(\mem[579][4] ), .S(n8533), .Z(n4527)
         );
  MUX2_X1 U23481 ( .A(\mem[576][4] ), .B(\mem[577][4] ), .S(n8398), .Z(n4528)
         );
  MUX2_X1 U23482 ( .A(n4528), .B(n4527), .S(n8272), .Z(n4529) );
  MUX2_X1 U23483 ( .A(n4529), .B(n4526), .S(n8240), .Z(n4530) );
  MUX2_X1 U23484 ( .A(n4530), .B(n4523), .S(n8201), .Z(n4531) );
  MUX2_X1 U23485 ( .A(n4531), .B(n4516), .S(n8188), .Z(n4532) );
  MUX2_X1 U23486 ( .A(n4532), .B(n4501), .S(n8185), .Z(n4533) );
  MUX2_X1 U23487 ( .A(\mem[574][4] ), .B(\mem[575][4] ), .S(n8503), .Z(n4534)
         );
  MUX2_X1 U23488 ( .A(\mem[572][4] ), .B(\mem[573][4] ), .S(n8510), .Z(n4535)
         );
  MUX2_X1 U23489 ( .A(n4535), .B(n4534), .S(n8282), .Z(n4536) );
  MUX2_X1 U23490 ( .A(\mem[570][4] ), .B(\mem[571][4] ), .S(n8511), .Z(n4537)
         );
  MUX2_X1 U23491 ( .A(\mem[568][4] ), .B(\mem[569][4] ), .S(n8512), .Z(n4538)
         );
  MUX2_X1 U23492 ( .A(n4538), .B(n4537), .S(n8282), .Z(n4539) );
  MUX2_X1 U23493 ( .A(n4539), .B(n4536), .S(N20), .Z(n4540) );
  MUX2_X1 U23494 ( .A(\mem[566][4] ), .B(\mem[567][4] ), .S(n8507), .Z(n4541)
         );
  MUX2_X1 U23495 ( .A(\mem[564][4] ), .B(\mem[565][4] ), .S(n8508), .Z(n4542)
         );
  MUX2_X1 U23496 ( .A(n4542), .B(n4541), .S(n8284), .Z(n4543) );
  MUX2_X1 U23497 ( .A(\mem[562][4] ), .B(\mem[563][4] ), .S(n8509), .Z(n4544)
         );
  MUX2_X1 U23498 ( .A(\mem[560][4] ), .B(\mem[561][4] ), .S(n8516), .Z(n4545)
         );
  MUX2_X1 U23499 ( .A(n4545), .B(n4544), .S(n8285), .Z(n4546) );
  MUX2_X1 U23500 ( .A(n4546), .B(n4543), .S(n8225), .Z(n4547) );
  MUX2_X1 U23501 ( .A(n4547), .B(n4540), .S(n8216), .Z(n4548) );
  MUX2_X1 U23502 ( .A(\mem[558][4] ), .B(\mem[559][4] ), .S(n8517), .Z(n4549)
         );
  MUX2_X1 U23503 ( .A(\mem[556][4] ), .B(\mem[557][4] ), .S(n8518), .Z(n4550)
         );
  MUX2_X1 U23504 ( .A(n4550), .B(n4549), .S(n8286), .Z(n4551) );
  MUX2_X1 U23505 ( .A(\mem[554][4] ), .B(\mem[555][4] ), .S(n8513), .Z(n4552)
         );
  MUX2_X1 U23506 ( .A(\mem[552][4] ), .B(\mem[553][4] ), .S(n8514), .Z(n4553)
         );
  MUX2_X1 U23507 ( .A(n4553), .B(n4552), .S(n8353), .Z(n4554) );
  MUX2_X1 U23508 ( .A(n4554), .B(n4551), .S(n8253), .Z(n4555) );
  MUX2_X1 U23509 ( .A(\mem[550][4] ), .B(\mem[551][4] ), .S(n8484), .Z(n4556)
         );
  MUX2_X1 U23510 ( .A(\mem[548][4] ), .B(\mem[549][4] ), .S(n8485), .Z(n4557)
         );
  MUX2_X1 U23511 ( .A(n4557), .B(n4556), .S(n8354), .Z(n4558) );
  MUX2_X1 U23512 ( .A(\mem[546][4] ), .B(\mem[547][4] ), .S(n8492), .Z(n4559)
         );
  MUX2_X1 U23513 ( .A(\mem[544][4] ), .B(\mem[545][4] ), .S(n8493), .Z(n4560)
         );
  MUX2_X1 U23514 ( .A(n4560), .B(n4559), .S(n8355), .Z(n4561) );
  MUX2_X1 U23515 ( .A(n4561), .B(n4558), .S(n8228), .Z(n4562) );
  MUX2_X1 U23516 ( .A(n4562), .B(n4555), .S(n8219), .Z(n4563) );
  MUX2_X1 U23517 ( .A(n4563), .B(n4548), .S(n8188), .Z(n4564) );
  MUX2_X1 U23518 ( .A(\mem[542][4] ), .B(\mem[543][4] ), .S(n8494), .Z(n4565)
         );
  MUX2_X1 U23519 ( .A(\mem[540][4] ), .B(\mem[541][4] ), .S(n8489), .Z(n4566)
         );
  MUX2_X1 U23520 ( .A(n4566), .B(n4565), .S(n8308), .Z(n4567) );
  MUX2_X1 U23521 ( .A(\mem[538][4] ), .B(\mem[539][4] ), .S(n8490), .Z(n4568)
         );
  MUX2_X1 U23522 ( .A(\mem[536][4] ), .B(\mem[537][4] ), .S(n8491), .Z(n4569)
         );
  MUX2_X1 U23523 ( .A(n4569), .B(n4568), .S(n8309), .Z(n4570) );
  MUX2_X1 U23524 ( .A(n4570), .B(n4567), .S(n8258), .Z(n4571) );
  MUX2_X1 U23525 ( .A(\mem[534][4] ), .B(\mem[535][4] ), .S(n8498), .Z(n4572)
         );
  MUX2_X1 U23526 ( .A(\mem[532][4] ), .B(\mem[533][4] ), .S(n8499), .Z(n4573)
         );
  MUX2_X1 U23527 ( .A(n4573), .B(n4572), .S(n8310), .Z(n4574) );
  MUX2_X1 U23528 ( .A(\mem[530][4] ), .B(\mem[531][4] ), .S(n8500), .Z(n4575)
         );
  MUX2_X1 U23529 ( .A(\mem[528][4] ), .B(\mem[529][4] ), .S(n8495), .Z(n4576)
         );
  MUX2_X1 U23530 ( .A(n4576), .B(n4575), .S(n8305), .Z(n4577) );
  MUX2_X1 U23531 ( .A(n4577), .B(n4574), .S(n8224), .Z(n4578) );
  MUX2_X1 U23532 ( .A(n4578), .B(n4571), .S(n8197), .Z(n4579) );
  MUX2_X1 U23533 ( .A(\mem[526][4] ), .B(\mem[527][4] ), .S(n8413), .Z(n4580)
         );
  MUX2_X1 U23534 ( .A(\mem[524][4] ), .B(\mem[525][4] ), .S(n8420), .Z(n4581)
         );
  MUX2_X1 U23535 ( .A(n4581), .B(n4580), .S(n8284), .Z(n4582) );
  MUX2_X1 U23536 ( .A(\mem[522][4] ), .B(\mem[523][4] ), .S(n8421), .Z(n4583)
         );
  MUX2_X1 U23537 ( .A(\mem[520][4] ), .B(\mem[521][4] ), .S(n8422), .Z(n4584)
         );
  MUX2_X1 U23538 ( .A(n4584), .B(n4583), .S(n8284), .Z(n4585) );
  MUX2_X1 U23539 ( .A(n4585), .B(n4582), .S(n8223), .Z(n4586) );
  MUX2_X1 U23540 ( .A(\mem[518][4] ), .B(\mem[519][4] ), .S(n8417), .Z(n4587)
         );
  MUX2_X1 U23541 ( .A(\mem[516][4] ), .B(\mem[517][4] ), .S(n8418), .Z(n4588)
         );
  MUX2_X1 U23542 ( .A(n4588), .B(n4587), .S(n8284), .Z(n4589) );
  MUX2_X1 U23543 ( .A(\mem[514][4] ), .B(\mem[515][4] ), .S(n8419), .Z(n4590)
         );
  MUX2_X1 U23544 ( .A(\mem[512][4] ), .B(\mem[513][4] ), .S(n8426), .Z(n4591)
         );
  MUX2_X1 U23545 ( .A(n4591), .B(n4590), .S(n8284), .Z(n4592) );
  MUX2_X1 U23546 ( .A(n4592), .B(n4589), .S(n8231), .Z(n4593) );
  MUX2_X1 U23547 ( .A(n4593), .B(n4586), .S(n8201), .Z(n4594) );
  MUX2_X1 U23548 ( .A(n4594), .B(n4579), .S(n8188), .Z(n4595) );
  MUX2_X1 U23549 ( .A(n4595), .B(n4564), .S(N23), .Z(n4596) );
  MUX2_X1 U23550 ( .A(n4596), .B(n4533), .S(n8180), .Z(n4597) );
  MUX2_X1 U23551 ( .A(n4597), .B(n4470), .S(n8177), .Z(n4598) );
  MUX2_X1 U23552 ( .A(n4598), .B(n4343), .S(N26), .Z(n4599) );
  MUX2_X1 U23553 ( .A(\mem[510][4] ), .B(\mem[511][4] ), .S(n8427), .Z(n4600)
         );
  MUX2_X1 U23554 ( .A(\mem[508][4] ), .B(\mem[509][4] ), .S(n8428), .Z(n4601)
         );
  MUX2_X1 U23555 ( .A(n4601), .B(n4600), .S(n8284), .Z(n4602) );
  MUX2_X1 U23556 ( .A(\mem[506][4] ), .B(\mem[507][4] ), .S(n8423), .Z(n4603)
         );
  MUX2_X1 U23557 ( .A(\mem[504][4] ), .B(\mem[505][4] ), .S(n8424), .Z(n4604)
         );
  MUX2_X1 U23558 ( .A(n4604), .B(n4603), .S(n8284), .Z(n4605) );
  MUX2_X1 U23559 ( .A(n4605), .B(n4602), .S(n8220), .Z(n4606) );
  MUX2_X1 U23560 ( .A(\mem[502][4] ), .B(\mem[503][4] ), .S(n8425), .Z(n4607)
         );
  MUX2_X1 U23561 ( .A(\mem[500][4] ), .B(\mem[501][4] ), .S(n8438), .Z(n4608)
         );
  MUX2_X1 U23562 ( .A(n4608), .B(n4607), .S(n8284), .Z(n4609) );
  MUX2_X1 U23563 ( .A(\mem[498][4] ), .B(\mem[499][4] ), .S(n8530), .Z(n4610)
         );
  MUX2_X1 U23564 ( .A(\mem[496][4] ), .B(\mem[497][4] ), .S(n8489), .Z(n4611)
         );
  MUX2_X1 U23565 ( .A(n4611), .B(n4610), .S(n8284), .Z(n4612) );
  MUX2_X1 U23566 ( .A(n4612), .B(n4609), .S(n8222), .Z(n4613) );
  MUX2_X1 U23567 ( .A(n4613), .B(n4606), .S(n8202), .Z(n4614) );
  MUX2_X1 U23568 ( .A(\mem[494][4] ), .B(\mem[495][4] ), .S(n8376), .Z(n4615)
         );
  MUX2_X1 U23569 ( .A(\mem[492][4] ), .B(\mem[493][4] ), .S(n8399), .Z(n4616)
         );
  MUX2_X1 U23570 ( .A(n4616), .B(n4615), .S(n8284), .Z(n4617) );
  MUX2_X1 U23571 ( .A(\mem[490][4] ), .B(\mem[491][4] ), .S(n8533), .Z(n4618)
         );
  MUX2_X1 U23572 ( .A(\mem[488][4] ), .B(\mem[489][4] ), .S(n8502), .Z(n4619)
         );
  MUX2_X1 U23573 ( .A(n4619), .B(n4618), .S(n8284), .Z(n4620) );
  MUX2_X1 U23574 ( .A(n4620), .B(n4617), .S(n8221), .Z(n4621) );
  MUX2_X1 U23575 ( .A(\mem[486][4] ), .B(\mem[487][4] ), .S(n8487), .Z(n4622)
         );
  MUX2_X1 U23576 ( .A(\mem[484][4] ), .B(\mem[485][4] ), .S(n8409), .Z(n4623)
         );
  MUX2_X1 U23577 ( .A(n4623), .B(n4622), .S(n8284), .Z(n4624) );
  MUX2_X1 U23578 ( .A(\mem[482][4] ), .B(\mem[483][4] ), .S(n8454), .Z(n4625)
         );
  MUX2_X1 U23579 ( .A(\mem[480][4] ), .B(\mem[481][4] ), .S(n8410), .Z(n4626)
         );
  MUX2_X1 U23580 ( .A(n4626), .B(n4625), .S(n8284), .Z(n4627) );
  MUX2_X1 U23581 ( .A(n4627), .B(n4624), .S(n8245), .Z(n4628) );
  MUX2_X1 U23582 ( .A(n4628), .B(n4621), .S(n8203), .Z(n4629) );
  MUX2_X1 U23583 ( .A(n4629), .B(n4614), .S(n8188), .Z(n4630) );
  MUX2_X1 U23584 ( .A(\mem[478][4] ), .B(\mem[479][4] ), .S(n8439), .Z(n4631)
         );
  MUX2_X1 U23585 ( .A(\mem[476][4] ), .B(\mem[477][4] ), .S(n8440), .Z(n4632)
         );
  MUX2_X1 U23586 ( .A(n4632), .B(n4631), .S(n8285), .Z(n4633) );
  MUX2_X1 U23587 ( .A(\mem[474][4] ), .B(\mem[475][4] ), .S(n8435), .Z(n4634)
         );
  MUX2_X1 U23588 ( .A(\mem[472][4] ), .B(\mem[473][4] ), .S(n8436), .Z(n4635)
         );
  MUX2_X1 U23589 ( .A(n4635), .B(n4634), .S(n8285), .Z(n4636) );
  MUX2_X1 U23590 ( .A(n4636), .B(n4633), .S(n8224), .Z(n4637) );
  MUX2_X1 U23591 ( .A(\mem[470][4] ), .B(\mem[471][4] ), .S(n8437), .Z(n4638)
         );
  MUX2_X1 U23592 ( .A(\mem[468][4] ), .B(\mem[469][4] ), .S(n8444), .Z(n4639)
         );
  MUX2_X1 U23593 ( .A(n4639), .B(n4638), .S(n8285), .Z(n4640) );
  MUX2_X1 U23594 ( .A(\mem[466][4] ), .B(\mem[467][4] ), .S(n8445), .Z(n4641)
         );
  MUX2_X1 U23595 ( .A(\mem[464][4] ), .B(\mem[465][4] ), .S(n8441), .Z(n4642)
         );
  MUX2_X1 U23596 ( .A(n4642), .B(n4641), .S(n8285), .Z(n4643) );
  MUX2_X1 U23597 ( .A(n4643), .B(n4640), .S(n8229), .Z(n4644) );
  MUX2_X1 U23598 ( .A(n4644), .B(n4637), .S(n8204), .Z(n4645) );
  MUX2_X1 U23599 ( .A(\mem[462][4] ), .B(\mem[463][4] ), .S(n8442), .Z(n4646)
         );
  MUX2_X1 U23600 ( .A(\mem[460][4] ), .B(\mem[461][4] ), .S(n8443), .Z(n4647)
         );
  MUX2_X1 U23601 ( .A(n4647), .B(n4646), .S(n8285), .Z(n4648) );
  MUX2_X1 U23602 ( .A(\mem[458][4] ), .B(\mem[459][4] ), .S(n8458), .Z(n4649)
         );
  MUX2_X1 U23603 ( .A(\mem[456][4] ), .B(\mem[457][4] ), .S(n8453), .Z(n4650)
         );
  MUX2_X1 U23604 ( .A(n4650), .B(n4649), .S(n8285), .Z(n4651) );
  MUX2_X1 U23605 ( .A(n4651), .B(n4648), .S(n8265), .Z(n4652) );
  MUX2_X1 U23606 ( .A(\mem[454][4] ), .B(\mem[455][4] ), .S(n8507), .Z(n4653)
         );
  MUX2_X1 U23607 ( .A(\mem[452][4] ), .B(\mem[453][4] ), .S(n8508), .Z(n4654)
         );
  MUX2_X1 U23608 ( .A(n4654), .B(n4653), .S(n8285), .Z(n4655) );
  MUX2_X1 U23609 ( .A(\mem[450][4] ), .B(\mem[451][4] ), .S(n8509), .Z(n4656)
         );
  MUX2_X1 U23610 ( .A(\mem[448][4] ), .B(\mem[449][4] ), .S(n8516), .Z(n4657)
         );
  MUX2_X1 U23611 ( .A(n4657), .B(n4656), .S(n8285), .Z(n4658) );
  MUX2_X1 U23612 ( .A(n4658), .B(n4655), .S(n8263), .Z(n4659) );
  MUX2_X1 U23613 ( .A(n4659), .B(n4652), .S(n8205), .Z(n4660) );
  MUX2_X1 U23614 ( .A(n4660), .B(n4645), .S(n8188), .Z(n4661) );
  MUX2_X1 U23615 ( .A(n4661), .B(n4630), .S(n8185), .Z(n4662) );
  MUX2_X1 U23616 ( .A(\mem[446][4] ), .B(\mem[447][4] ), .S(n8517), .Z(n4663)
         );
  MUX2_X1 U23617 ( .A(\mem[444][4] ), .B(\mem[445][4] ), .S(n8518), .Z(n4664)
         );
  MUX2_X1 U23618 ( .A(n4664), .B(n4663), .S(n8285), .Z(n4665) );
  MUX2_X1 U23619 ( .A(\mem[442][4] ), .B(\mem[443][4] ), .S(n8513), .Z(n4666)
         );
  MUX2_X1 U23620 ( .A(\mem[440][4] ), .B(\mem[441][4] ), .S(n8514), .Z(n4667)
         );
  MUX2_X1 U23621 ( .A(n4667), .B(n4666), .S(n8285), .Z(n4668) );
  MUX2_X1 U23622 ( .A(n4668), .B(n4665), .S(n8246), .Z(n4669) );
  MUX2_X1 U23623 ( .A(\mem[438][4] ), .B(\mem[439][4] ), .S(n8515), .Z(n4670)
         );
  MUX2_X1 U23624 ( .A(\mem[436][4] ), .B(\mem[437][4] ), .S(n8522), .Z(n4671)
         );
  MUX2_X1 U23625 ( .A(n4671), .B(n4670), .S(n8285), .Z(n4672) );
  MUX2_X1 U23626 ( .A(\mem[434][4] ), .B(\mem[435][4] ), .S(n8523), .Z(n4673)
         );
  MUX2_X1 U23627 ( .A(\mem[432][4] ), .B(\mem[433][4] ), .S(n8524), .Z(n4674)
         );
  MUX2_X1 U23628 ( .A(n4674), .B(n4673), .S(n8285), .Z(n4675) );
  MUX2_X1 U23629 ( .A(n4675), .B(n4672), .S(n8220), .Z(n4676) );
  MUX2_X1 U23630 ( .A(n4676), .B(n4669), .S(n8205), .Z(n4677) );
  MUX2_X1 U23631 ( .A(\mem[430][4] ), .B(\mem[431][4] ), .S(n8494), .Z(n4678)
         );
  MUX2_X1 U23632 ( .A(\mem[428][4] ), .B(\mem[429][4] ), .S(n8489), .Z(n4679)
         );
  MUX2_X1 U23633 ( .A(n4679), .B(n4678), .S(n8286), .Z(n4680) );
  MUX2_X1 U23634 ( .A(\mem[426][4] ), .B(\mem[427][4] ), .S(n8490), .Z(n4681)
         );
  MUX2_X1 U23635 ( .A(\mem[424][4] ), .B(\mem[425][4] ), .S(n8491), .Z(n4682)
         );
  MUX2_X1 U23636 ( .A(n4682), .B(n4681), .S(n8286), .Z(n4683) );
  MUX2_X1 U23637 ( .A(n4683), .B(n4680), .S(n8226), .Z(n4684) );
  MUX2_X1 U23638 ( .A(\mem[422][4] ), .B(\mem[423][4] ), .S(n8498), .Z(n4685)
         );
  MUX2_X1 U23639 ( .A(\mem[420][4] ), .B(\mem[421][4] ), .S(n8499), .Z(n4686)
         );
  MUX2_X1 U23640 ( .A(n4686), .B(n4685), .S(n8286), .Z(n4687) );
  MUX2_X1 U23641 ( .A(\mem[418][4] ), .B(\mem[419][4] ), .S(n8500), .Z(n4688)
         );
  MUX2_X1 U23642 ( .A(\mem[416][4] ), .B(\mem[417][4] ), .S(n8495), .Z(n4689)
         );
  MUX2_X1 U23643 ( .A(n4689), .B(n4688), .S(n8286), .Z(n4690) );
  MUX2_X1 U23644 ( .A(n4690), .B(n4687), .S(n8220), .Z(n4691) );
  MUX2_X1 U23645 ( .A(n4691), .B(n4684), .S(n8207), .Z(n4692) );
  MUX2_X1 U23646 ( .A(n4692), .B(n4677), .S(n8188), .Z(n4693) );
  MUX2_X1 U23647 ( .A(\mem[414][4] ), .B(\mem[415][4] ), .S(n8496), .Z(n4694)
         );
  MUX2_X1 U23648 ( .A(\mem[412][4] ), .B(\mem[413][4] ), .S(n8497), .Z(n4695)
         );
  MUX2_X1 U23649 ( .A(n4695), .B(n4694), .S(n8286), .Z(n4696) );
  MUX2_X1 U23650 ( .A(\mem[410][4] ), .B(\mem[411][4] ), .S(n8504), .Z(n4697)
         );
  MUX2_X1 U23651 ( .A(\mem[408][4] ), .B(\mem[409][4] ), .S(n8505), .Z(n4698)
         );
  MUX2_X1 U23652 ( .A(n4698), .B(n4697), .S(n8286), .Z(n4699) );
  MUX2_X1 U23653 ( .A(n4699), .B(n4696), .S(n8264), .Z(n4700) );
  MUX2_X1 U23654 ( .A(\mem[406][4] ), .B(\mem[407][4] ), .S(n8407), .Z(n4701)
         );
  MUX2_X1 U23655 ( .A(\mem[404][4] ), .B(\mem[405][4] ), .S(n8408), .Z(n4702)
         );
  MUX2_X1 U23656 ( .A(n4702), .B(n4701), .S(n8286), .Z(n4703) );
  MUX2_X1 U23657 ( .A(\mem[402][4] ), .B(\mem[403][4] ), .S(n8423), .Z(n4704)
         );
  MUX2_X1 U23658 ( .A(\mem[400][4] ), .B(\mem[401][4] ), .S(n8470), .Z(n4705)
         );
  MUX2_X1 U23659 ( .A(n4705), .B(n4704), .S(n8286), .Z(n4706) );
  MUX2_X1 U23660 ( .A(n4706), .B(n4703), .S(n8265), .Z(n4707) );
  MUX2_X1 U23661 ( .A(n4707), .B(n4700), .S(n8208), .Z(n4708) );
  MUX2_X1 U23662 ( .A(\mem[398][4] ), .B(\mem[399][4] ), .S(n8465), .Z(n4709)
         );
  MUX2_X1 U23663 ( .A(\mem[396][4] ), .B(\mem[397][4] ), .S(n8466), .Z(n4710)
         );
  MUX2_X1 U23664 ( .A(n4710), .B(n4709), .S(n8286), .Z(n4711) );
  MUX2_X1 U23665 ( .A(\mem[394][4] ), .B(\mem[395][4] ), .S(n8467), .Z(n4712)
         );
  MUX2_X1 U23666 ( .A(\mem[392][4] ), .B(\mem[393][4] ), .S(n8474), .Z(n4713)
         );
  MUX2_X1 U23667 ( .A(n4713), .B(n4712), .S(n8286), .Z(n4714) );
  MUX2_X1 U23668 ( .A(n4714), .B(n4711), .S(n8241), .Z(n4715) );
  MUX2_X1 U23669 ( .A(\mem[390][4] ), .B(\mem[391][4] ), .S(n8475), .Z(n4716)
         );
  MUX2_X1 U23670 ( .A(\mem[388][4] ), .B(\mem[389][4] ), .S(n8476), .Z(n4717)
         );
  MUX2_X1 U23671 ( .A(n4717), .B(n4716), .S(n8286), .Z(n4718) );
  MUX2_X1 U23672 ( .A(\mem[386][4] ), .B(\mem[387][4] ), .S(n8471), .Z(n4719)
         );
  MUX2_X1 U23673 ( .A(\mem[384][4] ), .B(\mem[385][4] ), .S(n8472), .Z(n4720)
         );
  MUX2_X1 U23674 ( .A(n4720), .B(n4719), .S(n8286), .Z(n4721) );
  MUX2_X1 U23675 ( .A(n4721), .B(n4718), .S(n8225), .Z(n4722) );
  MUX2_X1 U23676 ( .A(n4722), .B(n4715), .S(n8209), .Z(n4723) );
  MUX2_X1 U23677 ( .A(n4723), .B(n4708), .S(n8188), .Z(n4724) );
  MUX2_X1 U23678 ( .A(n4724), .B(n4693), .S(n8181), .Z(n4725) );
  MUX2_X1 U23679 ( .A(n4725), .B(n4662), .S(n8178), .Z(n4726) );
  MUX2_X1 U23680 ( .A(\mem[382][4] ), .B(\mem[383][4] ), .S(n8475), .Z(n4727)
         );
  MUX2_X1 U23681 ( .A(\mem[380][4] ), .B(\mem[381][4] ), .S(n8476), .Z(n4728)
         );
  MUX2_X1 U23682 ( .A(n4728), .B(n4727), .S(n8336), .Z(n4729) );
  MUX2_X1 U23683 ( .A(\mem[378][4] ), .B(\mem[379][4] ), .S(n8471), .Z(n4730)
         );
  MUX2_X1 U23684 ( .A(\mem[376][4] ), .B(\mem[377][4] ), .S(n8472), .Z(n4731)
         );
  MUX2_X1 U23685 ( .A(n4731), .B(n4730), .S(n8337), .Z(n4732) );
  MUX2_X1 U23686 ( .A(n4732), .B(n4729), .S(n8264), .Z(n4733) );
  MUX2_X1 U23687 ( .A(\mem[374][4] ), .B(\mem[375][4] ), .S(n8473), .Z(n4734)
         );
  MUX2_X1 U23688 ( .A(\mem[372][4] ), .B(\mem[373][4] ), .S(n8480), .Z(n4735)
         );
  MUX2_X1 U23689 ( .A(n4735), .B(n4734), .S(n8344), .Z(n4736) );
  MUX2_X1 U23690 ( .A(\mem[370][4] ), .B(\mem[371][4] ), .S(n8481), .Z(n4737)
         );
  MUX2_X1 U23691 ( .A(\mem[368][4] ), .B(\mem[369][4] ), .S(n8482), .Z(n4738)
         );
  MUX2_X1 U23692 ( .A(n4738), .B(n4737), .S(n8345), .Z(n4739) );
  MUX2_X1 U23693 ( .A(n4739), .B(n4736), .S(n8256), .Z(n4740) );
  MUX2_X1 U23694 ( .A(n4740), .B(n4733), .S(n8218), .Z(n4741) );
  MUX2_X1 U23695 ( .A(\mem[366][4] ), .B(\mem[367][4] ), .S(n8477), .Z(n4742)
         );
  MUX2_X1 U23696 ( .A(\mem[364][4] ), .B(\mem[365][4] ), .S(n8478), .Z(n4743)
         );
  MUX2_X1 U23697 ( .A(n4743), .B(n4742), .S(n8346), .Z(n4744) );
  MUX2_X1 U23698 ( .A(\mem[362][4] ), .B(\mem[363][4] ), .S(n8479), .Z(n4745)
         );
  MUX2_X1 U23699 ( .A(\mem[360][4] ), .B(\mem[361][4] ), .S(n8395), .Z(n4746)
         );
  MUX2_X1 U23700 ( .A(n4746), .B(n4745), .S(n8341), .Z(n4747) );
  MUX2_X1 U23701 ( .A(n4747), .B(n4744), .S(n8257), .Z(n4748) );
  MUX2_X1 U23702 ( .A(\mem[358][4] ), .B(\mem[359][4] ), .S(n8441), .Z(n4749)
         );
  MUX2_X1 U23703 ( .A(\mem[356][4] ), .B(\mem[357][4] ), .S(n8442), .Z(n4750)
         );
  MUX2_X1 U23704 ( .A(n4750), .B(n4749), .S(n8342), .Z(n4751) );
  MUX2_X1 U23705 ( .A(\mem[354][4] ), .B(\mem[355][4] ), .S(n8443), .Z(n4752)
         );
  MUX2_X1 U23706 ( .A(\mem[352][4] ), .B(\mem[353][4] ), .S(n8450), .Z(n4753)
         );
  MUX2_X1 U23707 ( .A(n4753), .B(n4752), .S(n8343), .Z(n4754) );
  MUX2_X1 U23708 ( .A(n4754), .B(n4751), .S(n8258), .Z(n4755) );
  MUX2_X1 U23709 ( .A(n4755), .B(n4748), .S(n8212), .Z(n4756) );
  MUX2_X1 U23710 ( .A(n4756), .B(n4741), .S(n8196), .Z(n4757) );
  MUX2_X1 U23711 ( .A(\mem[350][4] ), .B(\mem[351][4] ), .S(n8451), .Z(n4758)
         );
  MUX2_X1 U23712 ( .A(\mem[348][4] ), .B(\mem[349][4] ), .S(n8452), .Z(n4759)
         );
  MUX2_X1 U23713 ( .A(n4759), .B(n4758), .S(n8350), .Z(n4760) );
  MUX2_X1 U23714 ( .A(\mem[346][4] ), .B(\mem[347][4] ), .S(n8447), .Z(n4761)
         );
  MUX2_X1 U23715 ( .A(\mem[344][4] ), .B(\mem[345][4] ), .S(n8448), .Z(n4762)
         );
  MUX2_X1 U23716 ( .A(n4762), .B(n4761), .S(n8351), .Z(n4763) );
  MUX2_X1 U23717 ( .A(n4763), .B(n4760), .S(N20), .Z(n4764) );
  MUX2_X1 U23718 ( .A(\mem[342][4] ), .B(\mem[343][4] ), .S(n8449), .Z(n4765)
         );
  MUX2_X1 U23719 ( .A(\mem[340][4] ), .B(\mem[341][4] ), .S(n8456), .Z(n4766)
         );
  MUX2_X1 U23720 ( .A(n4766), .B(n4765), .S(n8352), .Z(n4767) );
  MUX2_X1 U23721 ( .A(\mem[338][4] ), .B(\mem[339][4] ), .S(n8457), .Z(n4768)
         );
  MUX2_X1 U23722 ( .A(\mem[336][4] ), .B(\mem[337][4] ), .S(n8458), .Z(n4769)
         );
  MUX2_X1 U23723 ( .A(n4769), .B(n4768), .S(n8347), .Z(n4770) );
  MUX2_X1 U23724 ( .A(n4770), .B(n4767), .S(n8238), .Z(n4771) );
  MUX2_X1 U23725 ( .A(n4771), .B(n4764), .S(n8213), .Z(n4772) );
  MUX2_X1 U23726 ( .A(\mem[334][4] ), .B(\mem[335][4] ), .S(n8533), .Z(n4773)
         );
  MUX2_X1 U23727 ( .A(\mem[332][4] ), .B(\mem[333][4] ), .S(n8398), .Z(n4774)
         );
  MUX2_X1 U23728 ( .A(n4774), .B(n4773), .S(n8303), .Z(n4775) );
  MUX2_X1 U23729 ( .A(\mem[330][4] ), .B(\mem[331][4] ), .S(n8399), .Z(n4776)
         );
  MUX2_X1 U23730 ( .A(\mem[328][4] ), .B(\mem[329][4] ), .S(n8395), .Z(n4777)
         );
  MUX2_X1 U23731 ( .A(n4777), .B(n4776), .S(n8304), .Z(n4778) );
  MUX2_X1 U23732 ( .A(n4778), .B(n4775), .S(n8263), .Z(n4779) );
  MUX2_X1 U23733 ( .A(\mem[326][4] ), .B(\mem[327][4] ), .S(n8396), .Z(n4780)
         );
  MUX2_X1 U23734 ( .A(\mem[324][4] ), .B(\mem[325][4] ), .S(n8397), .Z(n4781)
         );
  MUX2_X1 U23735 ( .A(n4781), .B(n4780), .S(n8299), .Z(n4782) );
  MUX2_X1 U23736 ( .A(\mem[322][4] ), .B(\mem[323][4] ), .S(n8404), .Z(n4783)
         );
  MUX2_X1 U23737 ( .A(\mem[320][4] ), .B(\mem[321][4] ), .S(n8405), .Z(n4784)
         );
  MUX2_X1 U23738 ( .A(n4784), .B(n4783), .S(n8300), .Z(n4785) );
  MUX2_X1 U23739 ( .A(n4785), .B(n4782), .S(n8264), .Z(n4786) );
  MUX2_X1 U23740 ( .A(n4786), .B(n4779), .S(n8214), .Z(n4787) );
  MUX2_X1 U23741 ( .A(n4787), .B(n4772), .S(n8196), .Z(n4788) );
  MUX2_X1 U23742 ( .A(n4788), .B(n4757), .S(N23), .Z(n4789) );
  MUX2_X1 U23743 ( .A(\mem[318][4] ), .B(\mem[319][4] ), .S(n8406), .Z(n4790)
         );
  MUX2_X1 U23744 ( .A(\mem[316][4] ), .B(\mem[317][4] ), .S(n8401), .Z(n4791)
         );
  MUX2_X1 U23745 ( .A(n4791), .B(n4790), .S(n8301), .Z(n4792) );
  MUX2_X1 U23746 ( .A(\mem[314][4] ), .B(\mem[315][4] ), .S(n8402), .Z(n4793)
         );
  MUX2_X1 U23747 ( .A(\mem[312][4] ), .B(\mem[313][4] ), .S(n8403), .Z(n4794)
         );
  MUX2_X1 U23748 ( .A(n4794), .B(n4793), .S(N19), .Z(n4795) );
  MUX2_X1 U23749 ( .A(n4795), .B(n4792), .S(n8246), .Z(n4796) );
  MUX2_X1 U23750 ( .A(\mem[310][4] ), .B(\mem[311][4] ), .S(n8429), .Z(n4797)
         );
  MUX2_X1 U23751 ( .A(\mem[308][4] ), .B(\mem[309][4] ), .S(n8430), .Z(n4798)
         );
  MUX2_X1 U23752 ( .A(n4798), .B(n4797), .S(n8327), .Z(n4799) );
  MUX2_X1 U23753 ( .A(\mem[306][4] ), .B(\mem[307][4] ), .S(n8431), .Z(n4800)
         );
  MUX2_X1 U23754 ( .A(\mem[304][4] ), .B(\mem[305][4] ), .S(n8438), .Z(n4801)
         );
  MUX2_X1 U23755 ( .A(n4801), .B(n4800), .S(n8328), .Z(n4802) );
  MUX2_X1 U23756 ( .A(n4802), .B(n4799), .S(n8243), .Z(n4803) );
  MUX2_X1 U23757 ( .A(n4803), .B(n4796), .S(n8211), .Z(n4804) );
  MUX2_X1 U23758 ( .A(\mem[302][4] ), .B(\mem[303][4] ), .S(n8439), .Z(n4805)
         );
  MUX2_X1 U23759 ( .A(\mem[300][4] ), .B(\mem[301][4] ), .S(n8440), .Z(n4806)
         );
  MUX2_X1 U23760 ( .A(n4806), .B(n4805), .S(n8323), .Z(n4807) );
  MUX2_X1 U23761 ( .A(\mem[298][4] ), .B(\mem[299][4] ), .S(n8435), .Z(n4808)
         );
  MUX2_X1 U23762 ( .A(\mem[296][4] ), .B(\mem[297][4] ), .S(n8436), .Z(n4809)
         );
  MUX2_X1 U23763 ( .A(n4809), .B(n4808), .S(n8324), .Z(n4810) );
  MUX2_X1 U23764 ( .A(n4810), .B(n4807), .S(n8249), .Z(n4811) );
  MUX2_X1 U23765 ( .A(\mem[294][4] ), .B(\mem[295][4] ), .S(n8437), .Z(n4812)
         );
  MUX2_X1 U23766 ( .A(\mem[292][4] ), .B(\mem[293][4] ), .S(n8444), .Z(n4813)
         );
  MUX2_X1 U23767 ( .A(n4813), .B(n4812), .S(n8325), .Z(n4814) );
  MUX2_X1 U23768 ( .A(\mem[290][4] ), .B(\mem[291][4] ), .S(n8445), .Z(n4815)
         );
  MUX2_X1 U23769 ( .A(\mem[288][4] ), .B(\mem[289][4] ), .S(n8446), .Z(n4816)
         );
  MUX2_X1 U23770 ( .A(n4816), .B(n4815), .S(n8332), .Z(n4817) );
  MUX2_X1 U23771 ( .A(n4817), .B(n4814), .S(n8236), .Z(n4818) );
  MUX2_X1 U23772 ( .A(n4818), .B(n4811), .S(N21), .Z(n4819) );
  MUX2_X1 U23773 ( .A(n4819), .B(n4804), .S(n8189), .Z(n4820) );
  MUX2_X1 U23774 ( .A(\mem[286][4] ), .B(\mem[287][4] ), .S(n8368), .Z(n4821)
         );
  MUX2_X1 U23775 ( .A(\mem[284][4] ), .B(\mem[285][4] ), .S(n8367), .Z(n4822)
         );
  MUX2_X1 U23776 ( .A(n4822), .B(n4821), .S(n8266), .Z(n4823) );
  MUX2_X1 U23777 ( .A(\mem[282][4] ), .B(\mem[283][4] ), .S(n8366), .Z(n4824)
         );
  MUX2_X1 U23778 ( .A(\mem[280][4] ), .B(\mem[281][4] ), .S(n8365), .Z(n4825)
         );
  MUX2_X1 U23779 ( .A(n4825), .B(n4824), .S(n8268), .Z(n4826) );
  MUX2_X1 U23780 ( .A(n4826), .B(n4823), .S(n8263), .Z(n4827) );
  MUX2_X1 U23781 ( .A(\mem[278][4] ), .B(\mem[279][4] ), .S(n8386), .Z(n4828)
         );
  MUX2_X1 U23782 ( .A(\mem[276][4] ), .B(\mem[277][4] ), .S(n8531), .Z(n4829)
         );
  MUX2_X1 U23783 ( .A(n4829), .B(n4828), .S(n8269), .Z(n4830) );
  MUX2_X1 U23784 ( .A(\mem[274][4] ), .B(\mem[275][4] ), .S(n8357), .Z(n4831)
         );
  MUX2_X1 U23785 ( .A(\mem[272][4] ), .B(\mem[273][4] ), .S(n8538), .Z(n4832)
         );
  MUX2_X1 U23786 ( .A(n4832), .B(n4831), .S(n8322), .Z(n4833) );
  MUX2_X1 U23787 ( .A(n4833), .B(n4830), .S(n8220), .Z(n4834) );
  MUX2_X1 U23788 ( .A(n4834), .B(n4827), .S(n8198), .Z(n4835) );
  MUX2_X1 U23789 ( .A(\mem[270][4] ), .B(\mem[271][4] ), .S(n8359), .Z(n4836)
         );
  MUX2_X1 U23790 ( .A(\mem[268][4] ), .B(\mem[269][4] ), .S(n8360), .Z(n4837)
         );
  MUX2_X1 U23791 ( .A(n4837), .B(n4836), .S(n8317), .Z(n4838) );
  MUX2_X1 U23792 ( .A(\mem[266][4] ), .B(\mem[267][4] ), .S(n8461), .Z(n4839)
         );
  MUX2_X1 U23793 ( .A(\mem[264][4] ), .B(\mem[265][4] ), .S(n8358), .Z(n4840)
         );
  MUX2_X1 U23794 ( .A(n4840), .B(n4839), .S(n8318), .Z(n4841) );
  MUX2_X1 U23795 ( .A(n4841), .B(n4838), .S(n8264), .Z(n4842) );
  MUX2_X1 U23796 ( .A(\mem[262][4] ), .B(\mem[263][4] ), .S(n8388), .Z(n4843)
         );
  MUX2_X1 U23797 ( .A(\mem[260][4] ), .B(\mem[261][4] ), .S(n8382), .Z(n4844)
         );
  MUX2_X1 U23798 ( .A(n4844), .B(n4843), .S(n8319), .Z(n4845) );
  MUX2_X1 U23799 ( .A(\mem[258][4] ), .B(\mem[259][4] ), .S(n8378), .Z(n4846)
         );
  MUX2_X1 U23800 ( .A(\mem[256][4] ), .B(\mem[257][4] ), .S(n8377), .Z(n4847)
         );
  MUX2_X1 U23801 ( .A(n4847), .B(n4846), .S(n8283), .Z(n4848) );
  MUX2_X1 U23802 ( .A(n4848), .B(n4845), .S(n8265), .Z(n4849) );
  MUX2_X1 U23803 ( .A(n4849), .B(n4842), .S(n8199), .Z(n4850) );
  MUX2_X1 U23804 ( .A(n4850), .B(n4835), .S(n8186), .Z(n4851) );
  MUX2_X1 U23805 ( .A(n4851), .B(n4820), .S(N23), .Z(n4852) );
  MUX2_X1 U23806 ( .A(n4852), .B(n4789), .S(N24), .Z(n4853) );
  MUX2_X1 U23807 ( .A(n4853), .B(n4726), .S(n8177), .Z(n4854) );
  MUX2_X1 U23808 ( .A(\mem[254][4] ), .B(\mem[255][4] ), .S(n8490), .Z(n4855)
         );
  MUX2_X1 U23809 ( .A(\mem[252][4] ), .B(\mem[253][4] ), .S(n8385), .Z(n4856)
         );
  MUX2_X1 U23810 ( .A(n4856), .B(n4855), .S(n8290), .Z(n4857) );
  MUX2_X1 U23811 ( .A(\mem[250][4] ), .B(\mem[251][4] ), .S(n8383), .Z(n4858)
         );
  MUX2_X1 U23812 ( .A(\mem[248][4] ), .B(\mem[249][4] ), .S(n8376), .Z(n4859)
         );
  MUX2_X1 U23813 ( .A(n4859), .B(n4858), .S(n8291), .Z(n4860) );
  MUX2_X1 U23814 ( .A(n4860), .B(n4857), .S(n8233), .Z(n4861) );
  MUX2_X1 U23815 ( .A(\mem[246][4] ), .B(\mem[247][4] ), .S(n8387), .Z(n4862)
         );
  MUX2_X1 U23816 ( .A(\mem[244][4] ), .B(\mem[245][4] ), .S(n8381), .Z(n4863)
         );
  MUX2_X1 U23817 ( .A(n4863), .B(n4862), .S(n8292), .Z(n4864) );
  MUX2_X1 U23818 ( .A(\mem[242][4] ), .B(\mem[243][4] ), .S(n8380), .Z(n4865)
         );
  MUX2_X1 U23819 ( .A(\mem[240][4] ), .B(\mem[241][4] ), .S(n8379), .Z(n4866)
         );
  MUX2_X1 U23820 ( .A(n4866), .B(n4865), .S(n8287), .Z(n4867) );
  MUX2_X1 U23821 ( .A(n4867), .B(n4864), .S(N20), .Z(n4868) );
  MUX2_X1 U23822 ( .A(n4868), .B(n4861), .S(n8200), .Z(n4869) );
  MUX2_X1 U23823 ( .A(\mem[238][4] ), .B(\mem[239][4] ), .S(n8477), .Z(n4870)
         );
  MUX2_X1 U23824 ( .A(\mem[236][4] ), .B(\mem[237][4] ), .S(n8478), .Z(n4871)
         );
  MUX2_X1 U23825 ( .A(n4871), .B(n4870), .S(n8287), .Z(n4872) );
  MUX2_X1 U23826 ( .A(\mem[234][4] ), .B(\mem[235][4] ), .S(n8479), .Z(n4873)
         );
  MUX2_X1 U23827 ( .A(\mem[232][4] ), .B(\mem[233][4] ), .S(N18), .Z(n4874) );
  MUX2_X1 U23828 ( .A(n4874), .B(n4873), .S(n8287), .Z(n4875) );
  MUX2_X1 U23829 ( .A(n4875), .B(n4872), .S(n8249), .Z(n4876) );
  MUX2_X1 U23830 ( .A(\mem[230][4] ), .B(\mem[231][4] ), .S(n8430), .Z(n4877)
         );
  MUX2_X1 U23831 ( .A(\mem[228][4] ), .B(\mem[229][4] ), .S(n8468), .Z(n4878)
         );
  MUX2_X1 U23832 ( .A(n4878), .B(n4877), .S(n8287), .Z(n4879) );
  MUX2_X1 U23833 ( .A(\mem[226][4] ), .B(\mem[227][4] ), .S(n8460), .Z(n4880)
         );
  MUX2_X1 U23834 ( .A(\mem[224][4] ), .B(\mem[225][4] ), .S(n8469), .Z(n4881)
         );
  MUX2_X1 U23835 ( .A(n4881), .B(n4880), .S(n8287), .Z(n4882) );
  MUX2_X1 U23836 ( .A(n4882), .B(n4879), .S(n8225), .Z(n4883) );
  MUX2_X1 U23837 ( .A(n4883), .B(n4876), .S(n8215), .Z(n4884) );
  MUX2_X1 U23838 ( .A(n4884), .B(n4869), .S(n8187), .Z(n4885) );
  MUX2_X1 U23839 ( .A(\mem[222][4] ), .B(\mem[223][4] ), .S(n8537), .Z(n4886)
         );
  MUX2_X1 U23840 ( .A(\mem[220][4] ), .B(\mem[221][4] ), .S(n8388), .Z(n4887)
         );
  MUX2_X1 U23841 ( .A(n4887), .B(n4886), .S(n8287), .Z(n4888) );
  MUX2_X1 U23842 ( .A(\mem[218][4] ), .B(\mem[219][4] ), .S(n8369), .Z(n4889)
         );
  MUX2_X1 U23843 ( .A(\mem[216][4] ), .B(\mem[217][4] ), .S(n8373), .Z(n4890)
         );
  MUX2_X1 U23844 ( .A(n4890), .B(n4889), .S(n8287), .Z(n4891) );
  MUX2_X1 U23845 ( .A(n4891), .B(n4888), .S(n8224), .Z(n4892) );
  MUX2_X1 U23846 ( .A(\mem[214][4] ), .B(\mem[215][4] ), .S(n8517), .Z(n4893)
         );
  MUX2_X1 U23847 ( .A(\mem[212][4] ), .B(\mem[213][4] ), .S(n8518), .Z(n4894)
         );
  MUX2_X1 U23848 ( .A(n4894), .B(n4893), .S(n8287), .Z(n4895) );
  MUX2_X1 U23849 ( .A(\mem[210][4] ), .B(\mem[211][4] ), .S(n8513), .Z(n4896)
         );
  MUX2_X1 U23850 ( .A(\mem[208][4] ), .B(\mem[209][4] ), .S(n8514), .Z(n4897)
         );
  MUX2_X1 U23851 ( .A(n4897), .B(n4896), .S(n8287), .Z(n4898) );
  MUX2_X1 U23852 ( .A(n4898), .B(n4895), .S(n8223), .Z(n4899) );
  MUX2_X1 U23853 ( .A(n4899), .B(n4892), .S(n8219), .Z(n4900) );
  MUX2_X1 U23854 ( .A(\mem[206][4] ), .B(\mem[207][4] ), .S(n8515), .Z(n4901)
         );
  MUX2_X1 U23855 ( .A(\mem[204][4] ), .B(\mem[205][4] ), .S(n8522), .Z(n4902)
         );
  MUX2_X1 U23856 ( .A(n4902), .B(n4901), .S(n8287), .Z(n4903) );
  MUX2_X1 U23857 ( .A(\mem[202][4] ), .B(\mem[203][4] ), .S(n8523), .Z(n4904)
         );
  MUX2_X1 U23858 ( .A(\mem[200][4] ), .B(\mem[201][4] ), .S(n8524), .Z(n4905)
         );
  MUX2_X1 U23859 ( .A(n4905), .B(n4904), .S(n8287), .Z(n4906) );
  MUX2_X1 U23860 ( .A(n4906), .B(n4903), .S(N20), .Z(n4907) );
  MUX2_X1 U23861 ( .A(\mem[198][4] ), .B(\mem[199][4] ), .S(n8519), .Z(n4908)
         );
  MUX2_X1 U23862 ( .A(\mem[196][4] ), .B(\mem[197][4] ), .S(n8520), .Z(n4909)
         );
  MUX2_X1 U23863 ( .A(n4909), .B(n4908), .S(n8287), .Z(n4910) );
  MUX2_X1 U23864 ( .A(\mem[194][4] ), .B(\mem[195][4] ), .S(n8521), .Z(n4911)
         );
  MUX2_X1 U23865 ( .A(\mem[192][4] ), .B(\mem[193][4] ), .S(n8528), .Z(n4912)
         );
  MUX2_X1 U23866 ( .A(n4912), .B(n4911), .S(n8287), .Z(n4913) );
  MUX2_X1 U23867 ( .A(n4913), .B(n4910), .S(n8228), .Z(n4914) );
  MUX2_X1 U23868 ( .A(n4914), .B(n4907), .S(n8197), .Z(n4915) );
  MUX2_X1 U23869 ( .A(n4915), .B(n4900), .S(n8188), .Z(n4916) );
  MUX2_X1 U23870 ( .A(n4916), .B(n4885), .S(n8182), .Z(n4917) );
  MUX2_X1 U23871 ( .A(\mem[190][4] ), .B(\mem[191][4] ), .S(n8490), .Z(n4918)
         );
  MUX2_X1 U23872 ( .A(\mem[188][4] ), .B(\mem[189][4] ), .S(n8491), .Z(n4919)
         );
  MUX2_X1 U23873 ( .A(n4919), .B(n4918), .S(n8288), .Z(n4920) );
  MUX2_X1 U23874 ( .A(\mem[186][4] ), .B(\mem[187][4] ), .S(n8498), .Z(n4921)
         );
  MUX2_X1 U23875 ( .A(\mem[184][4] ), .B(\mem[185][4] ), .S(n8499), .Z(n4922)
         );
  MUX2_X1 U23876 ( .A(n4922), .B(n4921), .S(n8288), .Z(n4923) );
  MUX2_X1 U23877 ( .A(n4923), .B(n4920), .S(n8263), .Z(n4924) );
  MUX2_X1 U23878 ( .A(\mem[182][4] ), .B(\mem[183][4] ), .S(n8500), .Z(n4925)
         );
  MUX2_X1 U23879 ( .A(\mem[180][4] ), .B(\mem[181][4] ), .S(n8495), .Z(n4926)
         );
  MUX2_X1 U23880 ( .A(n4926), .B(n4925), .S(n8288), .Z(n4927) );
  MUX2_X1 U23881 ( .A(\mem[178][4] ), .B(\mem[179][4] ), .S(n8496), .Z(n4928)
         );
  MUX2_X1 U23882 ( .A(\mem[176][4] ), .B(\mem[177][4] ), .S(n8497), .Z(n4929)
         );
  MUX2_X1 U23883 ( .A(n4929), .B(n4928), .S(n8288), .Z(n4930) );
  MUX2_X1 U23884 ( .A(n4930), .B(n4927), .S(n8226), .Z(n4931) );
  MUX2_X1 U23885 ( .A(n4931), .B(n4924), .S(n8202), .Z(n4932) );
  MUX2_X1 U23886 ( .A(\mem[174][4] ), .B(\mem[175][4] ), .S(n8504), .Z(n4933)
         );
  MUX2_X1 U23887 ( .A(\mem[172][4] ), .B(\mem[173][4] ), .S(n8505), .Z(n4934)
         );
  MUX2_X1 U23888 ( .A(n4934), .B(n4933), .S(n8288), .Z(n4935) );
  MUX2_X1 U23889 ( .A(\mem[170][4] ), .B(\mem[171][4] ), .S(n8506), .Z(n4936)
         );
  MUX2_X1 U23890 ( .A(\mem[168][4] ), .B(\mem[169][4] ), .S(n8501), .Z(n4937)
         );
  MUX2_X1 U23891 ( .A(n4937), .B(n4936), .S(n8288), .Z(n4938) );
  MUX2_X1 U23892 ( .A(n4938), .B(n4935), .S(n8225), .Z(n4939) );
  MUX2_X1 U23893 ( .A(\mem[166][4] ), .B(\mem[167][4] ), .S(n8360), .Z(n4940)
         );
  MUX2_X1 U23894 ( .A(\mem[164][4] ), .B(\mem[165][4] ), .S(n8358), .Z(n4941)
         );
  MUX2_X1 U23895 ( .A(n4941), .B(n4940), .S(n8288), .Z(n4942) );
  MUX2_X1 U23896 ( .A(\mem[162][4] ), .B(\mem[163][4] ), .S(n8453), .Z(n4943)
         );
  MUX2_X1 U23897 ( .A(\mem[160][4] ), .B(\mem[161][4] ), .S(n8486), .Z(n4944)
         );
  MUX2_X1 U23898 ( .A(n4944), .B(n4943), .S(n8288), .Z(n4945) );
  MUX2_X1 U23899 ( .A(n4945), .B(n4942), .S(n8222), .Z(n4946) );
  MUX2_X1 U23900 ( .A(n4946), .B(n4939), .S(n8202), .Z(n4947) );
  MUX2_X1 U23901 ( .A(n4947), .B(n4932), .S(n8192), .Z(n4948) );
  MUX2_X1 U23902 ( .A(\mem[158][4] ), .B(\mem[159][4] ), .S(n8487), .Z(n4949)
         );
  MUX2_X1 U23903 ( .A(\mem[156][4] ), .B(\mem[157][4] ), .S(n8488), .Z(n4950)
         );
  MUX2_X1 U23904 ( .A(n4950), .B(n4949), .S(n8288), .Z(n4951) );
  MUX2_X1 U23905 ( .A(\mem[154][4] ), .B(\mem[155][4] ), .S(n8483), .Z(n4952)
         );
  MUX2_X1 U23906 ( .A(\mem[152][4] ), .B(\mem[153][4] ), .S(n8484), .Z(n4953)
         );
  MUX2_X1 U23907 ( .A(n4953), .B(n4952), .S(n8288), .Z(n4954) );
  MUX2_X1 U23908 ( .A(n4954), .B(n4951), .S(n8221), .Z(n4955) );
  MUX2_X1 U23909 ( .A(\mem[150][4] ), .B(\mem[151][4] ), .S(n8485), .Z(n4956)
         );
  MUX2_X1 U23910 ( .A(\mem[148][4] ), .B(\mem[149][4] ), .S(n8492), .Z(n4957)
         );
  MUX2_X1 U23911 ( .A(n4957), .B(n4956), .S(n8288), .Z(n4958) );
  MUX2_X1 U23912 ( .A(\mem[146][4] ), .B(\mem[147][4] ), .S(n8493), .Z(n4959)
         );
  MUX2_X1 U23913 ( .A(\mem[144][4] ), .B(\mem[145][4] ), .S(n8494), .Z(n4960)
         );
  MUX2_X1 U23914 ( .A(n4960), .B(n4959), .S(n8288), .Z(n4961) );
  MUX2_X1 U23915 ( .A(n4961), .B(n4958), .S(n8226), .Z(n4962) );
  MUX2_X1 U23916 ( .A(n4962), .B(n4955), .S(n8202), .Z(n4963) );
  MUX2_X1 U23917 ( .A(\mem[142][4] ), .B(\mem[143][4] ), .S(n8386), .Z(n4964)
         );
  MUX2_X1 U23918 ( .A(\mem[140][4] ), .B(\mem[141][4] ), .S(n8382), .Z(n4965)
         );
  MUX2_X1 U23919 ( .A(n4965), .B(n4964), .S(n8289), .Z(n4966) );
  MUX2_X1 U23920 ( .A(\mem[138][4] ), .B(\mem[139][4] ), .S(n8381), .Z(n4967)
         );
  MUX2_X1 U23921 ( .A(\mem[136][4] ), .B(\mem[137][4] ), .S(n8380), .Z(n4968)
         );
  MUX2_X1 U23922 ( .A(n4968), .B(n4967), .S(n8289), .Z(n4969) );
  MUX2_X1 U23923 ( .A(n4969), .B(n4966), .S(n8227), .Z(n4970) );
  MUX2_X1 U23924 ( .A(\mem[134][4] ), .B(\mem[135][4] ), .S(n8379), .Z(n4971)
         );
  MUX2_X1 U23925 ( .A(\mem[132][4] ), .B(\mem[133][4] ), .S(n8378), .Z(n4972)
         );
  MUX2_X1 U23926 ( .A(n4972), .B(n4971), .S(n8289), .Z(n4973) );
  MUX2_X1 U23927 ( .A(\mem[130][4] ), .B(\mem[131][4] ), .S(n8377), .Z(n4974)
         );
  MUX2_X1 U23928 ( .A(\mem[128][4] ), .B(\mem[129][4] ), .S(n8385), .Z(n4975)
         );
  MUX2_X1 U23929 ( .A(n4975), .B(n4974), .S(n8289), .Z(n4976) );
  MUX2_X1 U23930 ( .A(n4976), .B(n4973), .S(n8258), .Z(n4977) );
  MUX2_X1 U23931 ( .A(n4977), .B(n4970), .S(n8202), .Z(n4978) );
  MUX2_X1 U23932 ( .A(n4978), .B(n4963), .S(n8193), .Z(n4979) );
  MUX2_X1 U23933 ( .A(n4979), .B(n4948), .S(n8185), .Z(n4980) );
  MUX2_X1 U23934 ( .A(n4980), .B(n4917), .S(n8179), .Z(n4981) );
  MUX2_X1 U23935 ( .A(\mem[126][4] ), .B(\mem[127][4] ), .S(n8384), .Z(n4982)
         );
  MUX2_X1 U23936 ( .A(\mem[124][4] ), .B(\mem[125][4] ), .S(n8383), .Z(n4983)
         );
  MUX2_X1 U23937 ( .A(n4983), .B(n4982), .S(n8289), .Z(n4984) );
  MUX2_X1 U23938 ( .A(\mem[122][4] ), .B(\mem[123][4] ), .S(n8375), .Z(n4985)
         );
  MUX2_X1 U23939 ( .A(\mem[120][4] ), .B(\mem[121][4] ), .S(n8374), .Z(n4986)
         );
  MUX2_X1 U23940 ( .A(n4986), .B(n4985), .S(n8289), .Z(n4987) );
  MUX2_X1 U23941 ( .A(n4987), .B(n4984), .S(n8263), .Z(n4988) );
  MUX2_X1 U23942 ( .A(\mem[118][4] ), .B(\mem[119][4] ), .S(n8402), .Z(n4989)
         );
  MUX2_X1 U23943 ( .A(\mem[116][4] ), .B(\mem[117][4] ), .S(n8403), .Z(n4990)
         );
  MUX2_X1 U23944 ( .A(n4990), .B(n4989), .S(n8289), .Z(n4991) );
  MUX2_X1 U23945 ( .A(\mem[114][4] ), .B(\mem[115][4] ), .S(n8393), .Z(n4992)
         );
  MUX2_X1 U23946 ( .A(\mem[112][4] ), .B(\mem[113][4] ), .S(n8394), .Z(n4993)
         );
  MUX2_X1 U23947 ( .A(n4993), .B(n4992), .S(n8289), .Z(n4994) );
  MUX2_X1 U23948 ( .A(n4994), .B(n4991), .S(n8244), .Z(n4995) );
  MUX2_X1 U23949 ( .A(n4995), .B(n4988), .S(n8202), .Z(n4996) );
  MUX2_X1 U23950 ( .A(\mem[110][4] ), .B(\mem[111][4] ), .S(n8390), .Z(n4997)
         );
  MUX2_X1 U23951 ( .A(\mem[108][4] ), .B(\mem[109][4] ), .S(n8391), .Z(n4998)
         );
  MUX2_X1 U23952 ( .A(n4998), .B(n4997), .S(n8289), .Z(n4999) );
  MUX2_X1 U23953 ( .A(\mem[106][4] ), .B(\mem[107][4] ), .S(n8392), .Z(n5000)
         );
  MUX2_X1 U23954 ( .A(\mem[104][4] ), .B(\mem[105][4] ), .S(n8389), .Z(n5001)
         );
  MUX2_X1 U23955 ( .A(n5001), .B(n5000), .S(n8289), .Z(n5002) );
  MUX2_X1 U23956 ( .A(n5002), .B(n4999), .S(n8226), .Z(n5003) );
  MUX2_X1 U23957 ( .A(\mem[102][4] ), .B(\mem[103][4] ), .S(n8432), .Z(n5004)
         );
  MUX2_X1 U23958 ( .A(\mem[100][4] ), .B(\mem[101][4] ), .S(n8433), .Z(n5005)
         );
  MUX2_X1 U23959 ( .A(n5005), .B(n5004), .S(n8289), .Z(n5006) );
  MUX2_X1 U23960 ( .A(\mem[98][4] ), .B(\mem[99][4] ), .S(n8434), .Z(n5007) );
  MUX2_X1 U23961 ( .A(\mem[96][4] ), .B(\mem[97][4] ), .S(n8429), .Z(n5008) );
  MUX2_X1 U23962 ( .A(n5008), .B(n5007), .S(n8289), .Z(n5009) );
  MUX2_X1 U23963 ( .A(n5009), .B(n5006), .S(N20), .Z(n5010) );
  MUX2_X1 U23964 ( .A(n5010), .B(n5003), .S(n8202), .Z(n5011) );
  MUX2_X1 U23965 ( .A(n5011), .B(n4996), .S(n8190), .Z(n5012) );
  MUX2_X1 U23966 ( .A(\mem[94][4] ), .B(\mem[95][4] ), .S(n8407), .Z(n5013) );
  MUX2_X1 U23967 ( .A(\mem[92][4] ), .B(\mem[93][4] ), .S(n8407), .Z(n5014) );
  MUX2_X1 U23968 ( .A(n5014), .B(n5013), .S(n8290), .Z(n5015) );
  MUX2_X1 U23969 ( .A(\mem[90][4] ), .B(\mem[91][4] ), .S(n8407), .Z(n5016) );
  MUX2_X1 U23970 ( .A(\mem[88][4] ), .B(\mem[89][4] ), .S(n8407), .Z(n5017) );
  MUX2_X1 U23971 ( .A(n5017), .B(n5016), .S(n8290), .Z(n5018) );
  MUX2_X1 U23972 ( .A(n5018), .B(n5015), .S(n8263), .Z(n5019) );
  MUX2_X1 U23973 ( .A(\mem[86][4] ), .B(\mem[87][4] ), .S(n8407), .Z(n5020) );
  MUX2_X1 U23974 ( .A(\mem[84][4] ), .B(\mem[85][4] ), .S(n8407), .Z(n5021) );
  MUX2_X1 U23975 ( .A(n5021), .B(n5020), .S(n8290), .Z(n5022) );
  MUX2_X1 U23976 ( .A(\mem[82][4] ), .B(\mem[83][4] ), .S(n8407), .Z(n5023) );
  MUX2_X1 U23977 ( .A(\mem[80][4] ), .B(\mem[81][4] ), .S(n8407), .Z(n5024) );
  MUX2_X1 U23978 ( .A(n5024), .B(n5023), .S(n8290), .Z(n5025) );
  MUX2_X1 U23979 ( .A(n5025), .B(n5022), .S(n8226), .Z(n5026) );
  MUX2_X1 U23980 ( .A(n5026), .B(n5019), .S(n8202), .Z(n5027) );
  MUX2_X1 U23981 ( .A(\mem[78][4] ), .B(\mem[79][4] ), .S(n8407), .Z(n5028) );
  MUX2_X1 U23982 ( .A(\mem[76][4] ), .B(\mem[77][4] ), .S(n8407), .Z(n5029) );
  MUX2_X1 U23983 ( .A(n5029), .B(n5028), .S(n8290), .Z(n5030) );
  MUX2_X1 U23984 ( .A(\mem[74][4] ), .B(\mem[75][4] ), .S(n8407), .Z(n5031) );
  MUX2_X1 U23985 ( .A(\mem[72][4] ), .B(\mem[73][4] ), .S(n8407), .Z(n5032) );
  MUX2_X1 U23986 ( .A(n5032), .B(n5031), .S(n8290), .Z(n5033) );
  MUX2_X1 U23987 ( .A(n5033), .B(n5030), .S(n8226), .Z(n5034) );
  MUX2_X1 U23988 ( .A(\mem[70][4] ), .B(\mem[71][4] ), .S(n8408), .Z(n5035) );
  MUX2_X1 U23989 ( .A(\mem[68][4] ), .B(\mem[69][4] ), .S(n8408), .Z(n5036) );
  MUX2_X1 U23990 ( .A(n5036), .B(n5035), .S(n8290), .Z(n5037) );
  MUX2_X1 U23991 ( .A(\mem[66][4] ), .B(\mem[67][4] ), .S(n8408), .Z(n5038) );
  MUX2_X1 U23992 ( .A(\mem[64][4] ), .B(\mem[65][4] ), .S(n8408), .Z(n5039) );
  MUX2_X1 U23993 ( .A(n5039), .B(n5038), .S(n8290), .Z(n5040) );
  MUX2_X1 U23994 ( .A(n5040), .B(n5037), .S(N20), .Z(n5041) );
  MUX2_X1 U23995 ( .A(n5041), .B(n5034), .S(n8202), .Z(n5042) );
  MUX2_X1 U23996 ( .A(n5042), .B(n5027), .S(n8186), .Z(n5043) );
  MUX2_X1 U23997 ( .A(n5043), .B(n5012), .S(n8185), .Z(n5044) );
  MUX2_X1 U23998 ( .A(\mem[62][4] ), .B(\mem[63][4] ), .S(n8408), .Z(n5045) );
  MUX2_X1 U23999 ( .A(\mem[60][4] ), .B(\mem[61][4] ), .S(n8408), .Z(n5046) );
  MUX2_X1 U24000 ( .A(n5046), .B(n5045), .S(n8290), .Z(n5047) );
  MUX2_X1 U24001 ( .A(\mem[58][4] ), .B(\mem[59][4] ), .S(n8408), .Z(n5048) );
  MUX2_X1 U24002 ( .A(\mem[56][4] ), .B(\mem[57][4] ), .S(n8408), .Z(n5049) );
  MUX2_X1 U24003 ( .A(n5049), .B(n5048), .S(n8290), .Z(n5050) );
  MUX2_X1 U24004 ( .A(n5050), .B(n5047), .S(n8220), .Z(n5051) );
  MUX2_X1 U24005 ( .A(\mem[54][4] ), .B(\mem[55][4] ), .S(n8408), .Z(n5052) );
  MUX2_X1 U24006 ( .A(\mem[52][4] ), .B(\mem[53][4] ), .S(n8408), .Z(n5053) );
  MUX2_X1 U24007 ( .A(n5053), .B(n5052), .S(n8290), .Z(n5054) );
  MUX2_X1 U24008 ( .A(\mem[50][4] ), .B(\mem[51][4] ), .S(n8408), .Z(n5055) );
  MUX2_X1 U24009 ( .A(\mem[48][4] ), .B(\mem[49][4] ), .S(n8408), .Z(n5056) );
  MUX2_X1 U24010 ( .A(n5056), .B(n5055), .S(n8290), .Z(n5057) );
  MUX2_X1 U24011 ( .A(n5057), .B(n5054), .S(n8264), .Z(n5058) );
  MUX2_X1 U24012 ( .A(n5058), .B(n5051), .S(n8202), .Z(n5059) );
  MUX2_X1 U24013 ( .A(\mem[46][4] ), .B(\mem[47][4] ), .S(n8475), .Z(n5060) );
  MUX2_X1 U24014 ( .A(\mem[44][4] ), .B(\mem[45][4] ), .S(n8476), .Z(n5061) );
  MUX2_X1 U24015 ( .A(n5061), .B(n5060), .S(n8291), .Z(n5062) );
  MUX2_X1 U24016 ( .A(\mem[42][4] ), .B(\mem[43][4] ), .S(n8471), .Z(n5063) );
  MUX2_X1 U24017 ( .A(\mem[40][4] ), .B(\mem[41][4] ), .S(n8472), .Z(n5064) );
  MUX2_X1 U24018 ( .A(n5064), .B(n5063), .S(n8291), .Z(n5065) );
  MUX2_X1 U24019 ( .A(n5065), .B(n5062), .S(n8265), .Z(n5066) );
  MUX2_X1 U24020 ( .A(\mem[38][4] ), .B(\mem[39][4] ), .S(n8473), .Z(n5067) );
  MUX2_X1 U24021 ( .A(\mem[36][4] ), .B(\mem[37][4] ), .S(n8480), .Z(n5068) );
  MUX2_X1 U24022 ( .A(n5068), .B(n5067), .S(n8291), .Z(n5069) );
  MUX2_X1 U24023 ( .A(\mem[34][4] ), .B(\mem[35][4] ), .S(n8481), .Z(n5070) );
  MUX2_X1 U24024 ( .A(\mem[32][4] ), .B(\mem[33][4] ), .S(n8482), .Z(n5071) );
  MUX2_X1 U24025 ( .A(n5071), .B(n5070), .S(n8291), .Z(n5072) );
  MUX2_X1 U24026 ( .A(n5072), .B(n5069), .S(n8234), .Z(n5073) );
  MUX2_X1 U24027 ( .A(n5073), .B(n5066), .S(n8202), .Z(n5074) );
  MUX2_X1 U24028 ( .A(n5074), .B(n5059), .S(n8191), .Z(n5075) );
  MUX2_X1 U24029 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n8477), .Z(n5076) );
  MUX2_X1 U24030 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n8478), .Z(n5077) );
  MUX2_X1 U24031 ( .A(n5077), .B(n5076), .S(n8291), .Z(n5078) );
  MUX2_X1 U24032 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n8479), .Z(n5079) );
  MUX2_X1 U24033 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n8410), .Z(n5080) );
  MUX2_X1 U24034 ( .A(n5080), .B(n5079), .S(n8291), .Z(n5081) );
  MUX2_X1 U24035 ( .A(n5081), .B(n5078), .S(n8223), .Z(n5082) );
  MUX2_X1 U24036 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n8409), .Z(n5083) );
  MUX2_X1 U24037 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n8409), .Z(n5084) );
  MUX2_X1 U24038 ( .A(n5084), .B(n5083), .S(n8291), .Z(n5085) );
  MUX2_X1 U24039 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n8409), .Z(n5086) );
  MUX2_X1 U24040 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n8409), .Z(n5087) );
  MUX2_X1 U24041 ( .A(n5087), .B(n5086), .S(n8291), .Z(n5088) );
  MUX2_X1 U24042 ( .A(n5088), .B(n5085), .S(n8225), .Z(n5089) );
  MUX2_X1 U24043 ( .A(n5089), .B(n5082), .S(n8202), .Z(n5090) );
  MUX2_X1 U24044 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n8409), .Z(n5091) );
  MUX2_X1 U24045 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n8409), .Z(n5092) );
  MUX2_X1 U24046 ( .A(n5092), .B(n5091), .S(n8291), .Z(n5093) );
  MUX2_X1 U24047 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n8409), .Z(n5094) );
  MUX2_X1 U24048 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n8409), .Z(n5095) );
  MUX2_X1 U24049 ( .A(n5095), .B(n5094), .S(n8291), .Z(n5096) );
  MUX2_X1 U24050 ( .A(n5096), .B(n5093), .S(n8224), .Z(n5097) );
  MUX2_X1 U24051 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n8409), .Z(n5098) );
  MUX2_X1 U24052 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n8409), .Z(n5099) );
  MUX2_X1 U24053 ( .A(n5099), .B(n5098), .S(n8291), .Z(n5100) );
  MUX2_X1 U24054 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n8409), .Z(n5101) );
  MUX2_X1 U24055 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n8409), .Z(n5102) );
  MUX2_X1 U24056 ( .A(n5102), .B(n5101), .S(n8291), .Z(n5103) );
  MUX2_X1 U24057 ( .A(n5103), .B(n5100), .S(n8223), .Z(n5104) );
  MUX2_X1 U24058 ( .A(n5104), .B(n5097), .S(n8202), .Z(n5105) );
  MUX2_X1 U24059 ( .A(n5105), .B(n5090), .S(N22), .Z(n5106) );
  MUX2_X1 U24060 ( .A(n5106), .B(n5075), .S(N23), .Z(n5107) );
  MUX2_X1 U24061 ( .A(n5107), .B(n5044), .S(N24), .Z(n5108) );
  MUX2_X1 U24062 ( .A(n5108), .B(n4981), .S(n8177), .Z(n5109) );
  MUX2_X1 U24063 ( .A(n5109), .B(n4854), .S(N26), .Z(n5110) );
  MUX2_X1 U24064 ( .A(n5110), .B(n4599), .S(N27), .Z(N31) );
  MUX2_X1 U24065 ( .A(\mem[1022][5] ), .B(\mem[1023][5] ), .S(n8411), .Z(n5111) );
  MUX2_X1 U24066 ( .A(\mem[1020][5] ), .B(\mem[1021][5] ), .S(n8412), .Z(n5112) );
  MUX2_X1 U24067 ( .A(n5112), .B(n5111), .S(n8292), .Z(n5113) );
  MUX2_X1 U24068 ( .A(\mem[1018][5] ), .B(\mem[1019][5] ), .S(n8413), .Z(n5114) );
  MUX2_X1 U24069 ( .A(\mem[1016][5] ), .B(\mem[1017][5] ), .S(n8420), .Z(n5115) );
  MUX2_X1 U24070 ( .A(n5115), .B(n5114), .S(n8292), .Z(n5116) );
  MUX2_X1 U24071 ( .A(n5116), .B(n5113), .S(n8263), .Z(n5117) );
  MUX2_X1 U24072 ( .A(\mem[1014][5] ), .B(\mem[1015][5] ), .S(n8421), .Z(n5118) );
  MUX2_X1 U24073 ( .A(\mem[1012][5] ), .B(\mem[1013][5] ), .S(n8422), .Z(n5119) );
  MUX2_X1 U24074 ( .A(n5119), .B(n5118), .S(n8292), .Z(n5120) );
  MUX2_X1 U24075 ( .A(\mem[1010][5] ), .B(\mem[1011][5] ), .S(n8417), .Z(n5121) );
  MUX2_X1 U24076 ( .A(\mem[1008][5] ), .B(\mem[1009][5] ), .S(n8418), .Z(n5122) );
  MUX2_X1 U24077 ( .A(n5122), .B(n5121), .S(n8292), .Z(n5123) );
  MUX2_X1 U24078 ( .A(n5123), .B(n5120), .S(n8260), .Z(n5124) );
  MUX2_X1 U24079 ( .A(n5124), .B(n5117), .S(n8203), .Z(n5125) );
  MUX2_X1 U24080 ( .A(\mem[1006][5] ), .B(\mem[1007][5] ), .S(n8419), .Z(n5126) );
  MUX2_X1 U24081 ( .A(\mem[1004][5] ), .B(\mem[1005][5] ), .S(n8426), .Z(n5127) );
  MUX2_X1 U24082 ( .A(n5127), .B(n5126), .S(n8292), .Z(n5128) );
  MUX2_X1 U24083 ( .A(\mem[1002][5] ), .B(\mem[1003][5] ), .S(n8427), .Z(n5129) );
  MUX2_X1 U24084 ( .A(\mem[1000][5] ), .B(\mem[1001][5] ), .S(n8428), .Z(n5130) );
  MUX2_X1 U24085 ( .A(n5130), .B(n5129), .S(n8292), .Z(n5131) );
  MUX2_X1 U24086 ( .A(n5131), .B(n5128), .S(n8239), .Z(n5132) );
  MUX2_X1 U24087 ( .A(\mem[998][5] ), .B(\mem[999][5] ), .S(n8410), .Z(n5133)
         );
  MUX2_X1 U24088 ( .A(\mem[996][5] ), .B(\mem[997][5] ), .S(n8410), .Z(n5134)
         );
  MUX2_X1 U24089 ( .A(n5134), .B(n5133), .S(n8292), .Z(n5135) );
  MUX2_X1 U24090 ( .A(\mem[994][5] ), .B(\mem[995][5] ), .S(n8410), .Z(n5136)
         );
  MUX2_X1 U24091 ( .A(\mem[992][5] ), .B(\mem[993][5] ), .S(n8410), .Z(n5137)
         );
  MUX2_X1 U24092 ( .A(n5137), .B(n5136), .S(n8292), .Z(n5138) );
  MUX2_X1 U24093 ( .A(n5138), .B(n5135), .S(n8265), .Z(n5139) );
  MUX2_X1 U24094 ( .A(n5139), .B(n5132), .S(n8203), .Z(n5140) );
  MUX2_X1 U24095 ( .A(n5140), .B(n5125), .S(n8189), .Z(n5141) );
  MUX2_X1 U24096 ( .A(\mem[990][5] ), .B(\mem[991][5] ), .S(n8410), .Z(n5142)
         );
  MUX2_X1 U24097 ( .A(\mem[988][5] ), .B(\mem[989][5] ), .S(n8410), .Z(n5143)
         );
  MUX2_X1 U24098 ( .A(n5143), .B(n5142), .S(n8292), .Z(n5144) );
  MUX2_X1 U24099 ( .A(\mem[986][5] ), .B(\mem[987][5] ), .S(n8410), .Z(n5145)
         );
  MUX2_X1 U24100 ( .A(\mem[984][5] ), .B(\mem[985][5] ), .S(n8410), .Z(n5146)
         );
  MUX2_X1 U24101 ( .A(n5146), .B(n5145), .S(n8292), .Z(n5147) );
  MUX2_X1 U24102 ( .A(n5147), .B(n5144), .S(n8253), .Z(n5148) );
  MUX2_X1 U24103 ( .A(\mem[982][5] ), .B(\mem[983][5] ), .S(n8410), .Z(n5149)
         );
  MUX2_X1 U24104 ( .A(\mem[980][5] ), .B(\mem[981][5] ), .S(n8410), .Z(n5150)
         );
  MUX2_X1 U24105 ( .A(n5150), .B(n5149), .S(n8292), .Z(n5151) );
  MUX2_X1 U24106 ( .A(\mem[978][5] ), .B(\mem[979][5] ), .S(n8410), .Z(n5152)
         );
  MUX2_X1 U24107 ( .A(\mem[976][5] ), .B(\mem[977][5] ), .S(n8410), .Z(n5153)
         );
  MUX2_X1 U24108 ( .A(n5153), .B(n5152), .S(n8292), .Z(n5154) );
  MUX2_X1 U24109 ( .A(n5154), .B(n5151), .S(n8238), .Z(n5155) );
  MUX2_X1 U24110 ( .A(n5155), .B(n5148), .S(n8203), .Z(n5156) );
  MUX2_X1 U24111 ( .A(\mem[974][5] ), .B(\mem[975][5] ), .S(n8411), .Z(n5157)
         );
  MUX2_X1 U24112 ( .A(\mem[972][5] ), .B(\mem[973][5] ), .S(n8411), .Z(n5158)
         );
  MUX2_X1 U24113 ( .A(n5158), .B(n5157), .S(n8293), .Z(n5159) );
  MUX2_X1 U24114 ( .A(\mem[970][5] ), .B(\mem[971][5] ), .S(n8411), .Z(n5160)
         );
  MUX2_X1 U24115 ( .A(\mem[968][5] ), .B(\mem[969][5] ), .S(n8411), .Z(n5161)
         );
  MUX2_X1 U24116 ( .A(n5161), .B(n5160), .S(n8293), .Z(n5162) );
  MUX2_X1 U24117 ( .A(n5162), .B(n5159), .S(n8244), .Z(n5163) );
  MUX2_X1 U24118 ( .A(\mem[966][5] ), .B(\mem[967][5] ), .S(n8411), .Z(n5164)
         );
  MUX2_X1 U24119 ( .A(\mem[964][5] ), .B(\mem[965][5] ), .S(n8411), .Z(n5165)
         );
  MUX2_X1 U24120 ( .A(n5165), .B(n5164), .S(n8293), .Z(n5166) );
  MUX2_X1 U24121 ( .A(\mem[962][5] ), .B(\mem[963][5] ), .S(n8411), .Z(n5167)
         );
  MUX2_X1 U24122 ( .A(\mem[960][5] ), .B(\mem[961][5] ), .S(n8411), .Z(n5168)
         );
  MUX2_X1 U24123 ( .A(n5168), .B(n5167), .S(n8293), .Z(n5169) );
  MUX2_X1 U24124 ( .A(n5169), .B(n5166), .S(n8237), .Z(n5170) );
  MUX2_X1 U24125 ( .A(n5170), .B(n5163), .S(n8203), .Z(n5171) );
  MUX2_X1 U24126 ( .A(n5171), .B(n5156), .S(n8186), .Z(n5172) );
  MUX2_X1 U24127 ( .A(n5172), .B(n5141), .S(n8185), .Z(n5173) );
  MUX2_X1 U24128 ( .A(\mem[958][5] ), .B(\mem[959][5] ), .S(n8411), .Z(n5174)
         );
  MUX2_X1 U24129 ( .A(\mem[956][5] ), .B(\mem[957][5] ), .S(n8411), .Z(n5175)
         );
  MUX2_X1 U24130 ( .A(n5175), .B(n5174), .S(n8293), .Z(n5176) );
  MUX2_X1 U24131 ( .A(\mem[954][5] ), .B(\mem[955][5] ), .S(n8411), .Z(n5177)
         );
  MUX2_X1 U24132 ( .A(\mem[952][5] ), .B(\mem[953][5] ), .S(n8411), .Z(n5178)
         );
  MUX2_X1 U24133 ( .A(n5178), .B(n5177), .S(n8293), .Z(n5179) );
  MUX2_X1 U24134 ( .A(n5179), .B(n5176), .S(n8247), .Z(n5180) );
  MUX2_X1 U24135 ( .A(\mem[950][5] ), .B(\mem[951][5] ), .S(n8412), .Z(n5181)
         );
  MUX2_X1 U24136 ( .A(\mem[948][5] ), .B(\mem[949][5] ), .S(n8412), .Z(n5182)
         );
  MUX2_X1 U24137 ( .A(n5182), .B(n5181), .S(n8293), .Z(n5183) );
  MUX2_X1 U24138 ( .A(\mem[946][5] ), .B(\mem[947][5] ), .S(n8412), .Z(n5184)
         );
  MUX2_X1 U24139 ( .A(\mem[944][5] ), .B(\mem[945][5] ), .S(n8412), .Z(n5185)
         );
  MUX2_X1 U24140 ( .A(n5185), .B(n5184), .S(n8293), .Z(n5186) );
  MUX2_X1 U24141 ( .A(n5186), .B(n5183), .S(n8243), .Z(n5187) );
  MUX2_X1 U24142 ( .A(n5187), .B(n5180), .S(n8203), .Z(n5188) );
  MUX2_X1 U24143 ( .A(\mem[942][5] ), .B(\mem[943][5] ), .S(n8412), .Z(n5189)
         );
  MUX2_X1 U24144 ( .A(\mem[940][5] ), .B(\mem[941][5] ), .S(n8412), .Z(n5190)
         );
  MUX2_X1 U24145 ( .A(n5190), .B(n5189), .S(n8293), .Z(n5191) );
  MUX2_X1 U24146 ( .A(\mem[938][5] ), .B(\mem[939][5] ), .S(n8412), .Z(n5192)
         );
  MUX2_X1 U24147 ( .A(\mem[936][5] ), .B(\mem[937][5] ), .S(n8412), .Z(n5193)
         );
  MUX2_X1 U24148 ( .A(n5193), .B(n5192), .S(n8293), .Z(n5194) );
  MUX2_X1 U24149 ( .A(n5194), .B(n5191), .S(n8225), .Z(n5195) );
  MUX2_X1 U24150 ( .A(\mem[934][5] ), .B(\mem[935][5] ), .S(n8412), .Z(n5196)
         );
  MUX2_X1 U24151 ( .A(\mem[932][5] ), .B(\mem[933][5] ), .S(n8412), .Z(n5197)
         );
  MUX2_X1 U24152 ( .A(n5197), .B(n5196), .S(n8293), .Z(n5198) );
  MUX2_X1 U24153 ( .A(\mem[930][5] ), .B(\mem[931][5] ), .S(n8412), .Z(n5199)
         );
  MUX2_X1 U24154 ( .A(\mem[928][5] ), .B(\mem[929][5] ), .S(n8412), .Z(n5200)
         );
  MUX2_X1 U24155 ( .A(n5200), .B(n5199), .S(n8293), .Z(n5201) );
  MUX2_X1 U24156 ( .A(n5201), .B(n5198), .S(n8261), .Z(n5202) );
  MUX2_X1 U24157 ( .A(n5202), .B(n5195), .S(n8203), .Z(n5203) );
  MUX2_X1 U24158 ( .A(n5203), .B(n5188), .S(n8187), .Z(n5204) );
  MUX2_X1 U24159 ( .A(\mem[926][5] ), .B(\mem[927][5] ), .S(n8413), .Z(n5205)
         );
  MUX2_X1 U24160 ( .A(\mem[924][5] ), .B(\mem[925][5] ), .S(n8413), .Z(n5206)
         );
  MUX2_X1 U24161 ( .A(n5206), .B(n5205), .S(n8294), .Z(n5207) );
  MUX2_X1 U24162 ( .A(\mem[922][5] ), .B(\mem[923][5] ), .S(n8413), .Z(n5208)
         );
  MUX2_X1 U24163 ( .A(\mem[920][5] ), .B(\mem[921][5] ), .S(n8413), .Z(n5209)
         );
  MUX2_X1 U24164 ( .A(n5209), .B(n5208), .S(n8294), .Z(n5210) );
  MUX2_X1 U24165 ( .A(n5210), .B(n5207), .S(n8255), .Z(n5211) );
  MUX2_X1 U24166 ( .A(\mem[918][5] ), .B(\mem[919][5] ), .S(n8413), .Z(n5212)
         );
  MUX2_X1 U24167 ( .A(\mem[916][5] ), .B(\mem[917][5] ), .S(n8413), .Z(n5213)
         );
  MUX2_X1 U24168 ( .A(n5213), .B(n5212), .S(n8294), .Z(n5214) );
  MUX2_X1 U24169 ( .A(\mem[914][5] ), .B(\mem[915][5] ), .S(n8413), .Z(n5215)
         );
  MUX2_X1 U24170 ( .A(\mem[912][5] ), .B(\mem[913][5] ), .S(n8413), .Z(n5216)
         );
  MUX2_X1 U24171 ( .A(n5216), .B(n5215), .S(n8294), .Z(n5217) );
  MUX2_X1 U24172 ( .A(n5217), .B(n5214), .S(n8250), .Z(n5218) );
  MUX2_X1 U24173 ( .A(n5218), .B(n5211), .S(n8203), .Z(n5219) );
  MUX2_X1 U24174 ( .A(\mem[910][5] ), .B(\mem[911][5] ), .S(n8413), .Z(n5220)
         );
  MUX2_X1 U24175 ( .A(\mem[908][5] ), .B(\mem[909][5] ), .S(n8413), .Z(n5221)
         );
  MUX2_X1 U24176 ( .A(n5221), .B(n5220), .S(n8294), .Z(n5222) );
  MUX2_X1 U24177 ( .A(\mem[906][5] ), .B(\mem[907][5] ), .S(n8413), .Z(n5223)
         );
  MUX2_X1 U24178 ( .A(\mem[904][5] ), .B(\mem[905][5] ), .S(n8413), .Z(n5224)
         );
  MUX2_X1 U24179 ( .A(n5224), .B(n5223), .S(n8294), .Z(n5225) );
  MUX2_X1 U24180 ( .A(n5225), .B(n5222), .S(n8251), .Z(n5226) );
  MUX2_X1 U24181 ( .A(\mem[902][5] ), .B(\mem[903][5] ), .S(n8414), .Z(n5227)
         );
  MUX2_X1 U24182 ( .A(\mem[900][5] ), .B(\mem[901][5] ), .S(n8414), .Z(n5228)
         );
  MUX2_X1 U24183 ( .A(n5228), .B(n5227), .S(n8294), .Z(n5229) );
  MUX2_X1 U24184 ( .A(\mem[898][5] ), .B(\mem[899][5] ), .S(n8414), .Z(n5230)
         );
  MUX2_X1 U24185 ( .A(\mem[896][5] ), .B(\mem[897][5] ), .S(n8414), .Z(n5231)
         );
  MUX2_X1 U24186 ( .A(n5231), .B(n5230), .S(n8294), .Z(n5232) );
  MUX2_X1 U24187 ( .A(n5232), .B(n5229), .S(n8252), .Z(n5233) );
  MUX2_X1 U24188 ( .A(n5233), .B(n5226), .S(n8203), .Z(n5234) );
  MUX2_X1 U24189 ( .A(n5234), .B(n5219), .S(n8188), .Z(n5235) );
  MUX2_X1 U24190 ( .A(n5235), .B(n5204), .S(n8181), .Z(n5236) );
  MUX2_X1 U24191 ( .A(n5236), .B(n5173), .S(n8178), .Z(n5237) );
  MUX2_X1 U24192 ( .A(\mem[894][5] ), .B(\mem[895][5] ), .S(n8414), .Z(n5238)
         );
  MUX2_X1 U24193 ( .A(\mem[892][5] ), .B(\mem[893][5] ), .S(n8414), .Z(n5239)
         );
  MUX2_X1 U24194 ( .A(n5239), .B(n5238), .S(n8294), .Z(n5240) );
  MUX2_X1 U24195 ( .A(\mem[890][5] ), .B(\mem[891][5] ), .S(n8414), .Z(n5241)
         );
  MUX2_X1 U24196 ( .A(\mem[888][5] ), .B(\mem[889][5] ), .S(n8414), .Z(n5242)
         );
  MUX2_X1 U24197 ( .A(n5242), .B(n5241), .S(n8294), .Z(n5243) );
  MUX2_X1 U24198 ( .A(n5243), .B(n5240), .S(n8259), .Z(n5244) );
  MUX2_X1 U24199 ( .A(\mem[886][5] ), .B(\mem[887][5] ), .S(n8414), .Z(n5245)
         );
  MUX2_X1 U24200 ( .A(\mem[884][5] ), .B(\mem[885][5] ), .S(n8414), .Z(n5246)
         );
  MUX2_X1 U24201 ( .A(n5246), .B(n5245), .S(n8294), .Z(n5247) );
  MUX2_X1 U24202 ( .A(\mem[882][5] ), .B(\mem[883][5] ), .S(n8414), .Z(n5248)
         );
  MUX2_X1 U24203 ( .A(\mem[880][5] ), .B(\mem[881][5] ), .S(n8414), .Z(n5249)
         );
  MUX2_X1 U24204 ( .A(n5249), .B(n5248), .S(n8294), .Z(n5250) );
  MUX2_X1 U24205 ( .A(n5250), .B(n5247), .S(n8260), .Z(n5251) );
  MUX2_X1 U24206 ( .A(n5251), .B(n5244), .S(n8203), .Z(n5252) );
  MUX2_X1 U24207 ( .A(\mem[878][5] ), .B(\mem[879][5] ), .S(n8415), .Z(n5253)
         );
  MUX2_X1 U24208 ( .A(\mem[876][5] ), .B(\mem[877][5] ), .S(n8415), .Z(n5254)
         );
  MUX2_X1 U24209 ( .A(n5254), .B(n5253), .S(n8295), .Z(n5255) );
  MUX2_X1 U24210 ( .A(\mem[874][5] ), .B(\mem[875][5] ), .S(n8415), .Z(n5256)
         );
  MUX2_X1 U24211 ( .A(\mem[872][5] ), .B(\mem[873][5] ), .S(n8415), .Z(n5257)
         );
  MUX2_X1 U24212 ( .A(n5257), .B(n5256), .S(n8295), .Z(n5258) );
  MUX2_X1 U24213 ( .A(n5258), .B(n5255), .S(n8261), .Z(n5259) );
  MUX2_X1 U24214 ( .A(\mem[870][5] ), .B(\mem[871][5] ), .S(n8415), .Z(n5260)
         );
  MUX2_X1 U24215 ( .A(\mem[868][5] ), .B(\mem[869][5] ), .S(n8415), .Z(n5261)
         );
  MUX2_X1 U24216 ( .A(n5261), .B(n5260), .S(n8295), .Z(n5262) );
  MUX2_X1 U24217 ( .A(\mem[866][5] ), .B(\mem[867][5] ), .S(n8415), .Z(n5263)
         );
  MUX2_X1 U24218 ( .A(\mem[864][5] ), .B(\mem[865][5] ), .S(n8415), .Z(n5264)
         );
  MUX2_X1 U24219 ( .A(n5264), .B(n5263), .S(n8295), .Z(n5265) );
  MUX2_X1 U24220 ( .A(n5265), .B(n5262), .S(n8256), .Z(n5266) );
  MUX2_X1 U24221 ( .A(n5266), .B(n5259), .S(n8203), .Z(n5267) );
  MUX2_X1 U24222 ( .A(n5267), .B(n5252), .S(n8192), .Z(n5268) );
  MUX2_X1 U24223 ( .A(\mem[862][5] ), .B(\mem[863][5] ), .S(n8415), .Z(n5269)
         );
  MUX2_X1 U24224 ( .A(\mem[860][5] ), .B(\mem[861][5] ), .S(n8415), .Z(n5270)
         );
  MUX2_X1 U24225 ( .A(n5270), .B(n5269), .S(n8295), .Z(n5271) );
  MUX2_X1 U24226 ( .A(\mem[858][5] ), .B(\mem[859][5] ), .S(n8415), .Z(n5272)
         );
  MUX2_X1 U24227 ( .A(\mem[856][5] ), .B(\mem[857][5] ), .S(n8415), .Z(n5273)
         );
  MUX2_X1 U24228 ( .A(n5273), .B(n5272), .S(n8295), .Z(n5274) );
  MUX2_X1 U24229 ( .A(n5274), .B(n5271), .S(n8257), .Z(n5275) );
  MUX2_X1 U24230 ( .A(\mem[854][5] ), .B(\mem[855][5] ), .S(n8416), .Z(n5276)
         );
  MUX2_X1 U24231 ( .A(\mem[852][5] ), .B(\mem[853][5] ), .S(n8416), .Z(n5277)
         );
  MUX2_X1 U24232 ( .A(n5277), .B(n5276), .S(n8295), .Z(n5278) );
  MUX2_X1 U24233 ( .A(\mem[850][5] ), .B(\mem[851][5] ), .S(n8416), .Z(n5279)
         );
  MUX2_X1 U24234 ( .A(\mem[848][5] ), .B(\mem[849][5] ), .S(n8416), .Z(n5280)
         );
  MUX2_X1 U24235 ( .A(n5280), .B(n5279), .S(n8295), .Z(n5281) );
  MUX2_X1 U24236 ( .A(n5281), .B(n5278), .S(n8258), .Z(n5282) );
  MUX2_X1 U24237 ( .A(n5282), .B(n5275), .S(n8203), .Z(n5283) );
  MUX2_X1 U24238 ( .A(\mem[846][5] ), .B(\mem[847][5] ), .S(n8416), .Z(n5284)
         );
  MUX2_X1 U24239 ( .A(\mem[844][5] ), .B(\mem[845][5] ), .S(n8416), .Z(n5285)
         );
  MUX2_X1 U24240 ( .A(n5285), .B(n5284), .S(n8295), .Z(n5286) );
  MUX2_X1 U24241 ( .A(\mem[842][5] ), .B(\mem[843][5] ), .S(n8416), .Z(n5287)
         );
  MUX2_X1 U24242 ( .A(\mem[840][5] ), .B(\mem[841][5] ), .S(n8416), .Z(n5288)
         );
  MUX2_X1 U24243 ( .A(n5288), .B(n5287), .S(n8295), .Z(n5289) );
  MUX2_X1 U24244 ( .A(n5289), .B(n5286), .S(N20), .Z(n5290) );
  MUX2_X1 U24245 ( .A(\mem[838][5] ), .B(\mem[839][5] ), .S(n8416), .Z(n5291)
         );
  MUX2_X1 U24246 ( .A(\mem[836][5] ), .B(\mem[837][5] ), .S(n8416), .Z(n5292)
         );
  MUX2_X1 U24247 ( .A(n5292), .B(n5291), .S(n8295), .Z(n5293) );
  MUX2_X1 U24248 ( .A(\mem[834][5] ), .B(\mem[835][5] ), .S(n8416), .Z(n5294)
         );
  MUX2_X1 U24249 ( .A(\mem[832][5] ), .B(\mem[833][5] ), .S(n8416), .Z(n5295)
         );
  MUX2_X1 U24250 ( .A(n5295), .B(n5294), .S(n8295), .Z(n5296) );
  MUX2_X1 U24251 ( .A(n5296), .B(n5293), .S(n8264), .Z(n5297) );
  MUX2_X1 U24252 ( .A(n5297), .B(n5290), .S(n8203), .Z(n5298) );
  MUX2_X1 U24253 ( .A(n5298), .B(n5283), .S(n8193), .Z(n5299) );
  MUX2_X1 U24254 ( .A(n5299), .B(n5268), .S(n8185), .Z(n5300) );
  MUX2_X1 U24255 ( .A(\mem[830][5] ), .B(\mem[831][5] ), .S(n8417), .Z(n5301)
         );
  MUX2_X1 U24256 ( .A(\mem[828][5] ), .B(\mem[829][5] ), .S(n8417), .Z(n5302)
         );
  MUX2_X1 U24257 ( .A(n5302), .B(n5301), .S(n8296), .Z(n5303) );
  MUX2_X1 U24258 ( .A(\mem[826][5] ), .B(\mem[827][5] ), .S(n8417), .Z(n5304)
         );
  MUX2_X1 U24259 ( .A(\mem[824][5] ), .B(\mem[825][5] ), .S(n8417), .Z(n5305)
         );
  MUX2_X1 U24260 ( .A(n5305), .B(n5304), .S(n8296), .Z(n5306) );
  MUX2_X1 U24261 ( .A(n5306), .B(n5303), .S(n8264), .Z(n5307) );
  MUX2_X1 U24262 ( .A(\mem[822][5] ), .B(\mem[823][5] ), .S(n8417), .Z(n5308)
         );
  MUX2_X1 U24263 ( .A(\mem[820][5] ), .B(\mem[821][5] ), .S(n8417), .Z(n5309)
         );
  MUX2_X1 U24264 ( .A(n5309), .B(n5308), .S(n8296), .Z(n5310) );
  MUX2_X1 U24265 ( .A(\mem[818][5] ), .B(\mem[819][5] ), .S(n8417), .Z(n5311)
         );
  MUX2_X1 U24266 ( .A(\mem[816][5] ), .B(\mem[817][5] ), .S(n8417), .Z(n5312)
         );
  MUX2_X1 U24267 ( .A(n5312), .B(n5311), .S(n8296), .Z(n5313) );
  MUX2_X1 U24268 ( .A(n5313), .B(n5310), .S(n8261), .Z(n5314) );
  MUX2_X1 U24269 ( .A(n5314), .B(n5307), .S(n8204), .Z(n5315) );
  MUX2_X1 U24270 ( .A(\mem[814][5] ), .B(\mem[815][5] ), .S(n8417), .Z(n5316)
         );
  MUX2_X1 U24271 ( .A(\mem[812][5] ), .B(\mem[813][5] ), .S(n8417), .Z(n5317)
         );
  MUX2_X1 U24272 ( .A(n5317), .B(n5316), .S(n8296), .Z(n5318) );
  MUX2_X1 U24273 ( .A(\mem[810][5] ), .B(\mem[811][5] ), .S(n8417), .Z(n5319)
         );
  MUX2_X1 U24274 ( .A(\mem[808][5] ), .B(\mem[809][5] ), .S(n8417), .Z(n5320)
         );
  MUX2_X1 U24275 ( .A(n5320), .B(n5319), .S(n8296), .Z(n5321) );
  MUX2_X1 U24276 ( .A(n5321), .B(n5318), .S(n8259), .Z(n5322) );
  MUX2_X1 U24277 ( .A(\mem[806][5] ), .B(\mem[807][5] ), .S(n8418), .Z(n5323)
         );
  MUX2_X1 U24278 ( .A(\mem[804][5] ), .B(\mem[805][5] ), .S(n8418), .Z(n5324)
         );
  MUX2_X1 U24279 ( .A(n5324), .B(n5323), .S(n8296), .Z(n5325) );
  MUX2_X1 U24280 ( .A(\mem[802][5] ), .B(\mem[803][5] ), .S(n8418), .Z(n5326)
         );
  MUX2_X1 U24281 ( .A(\mem[800][5] ), .B(\mem[801][5] ), .S(n8418), .Z(n5327)
         );
  MUX2_X1 U24282 ( .A(n5327), .B(n5326), .S(n8296), .Z(n5328) );
  MUX2_X1 U24283 ( .A(n5328), .B(n5325), .S(n8262), .Z(n5329) );
  MUX2_X1 U24284 ( .A(n5329), .B(n5322), .S(n8204), .Z(n5330) );
  MUX2_X1 U24285 ( .A(n5330), .B(n5315), .S(n8190), .Z(n5331) );
  MUX2_X1 U24286 ( .A(\mem[798][5] ), .B(\mem[799][5] ), .S(n8418), .Z(n5332)
         );
  MUX2_X1 U24287 ( .A(\mem[796][5] ), .B(\mem[797][5] ), .S(n8418), .Z(n5333)
         );
  MUX2_X1 U24288 ( .A(n5333), .B(n5332), .S(n8296), .Z(n5334) );
  MUX2_X1 U24289 ( .A(\mem[794][5] ), .B(\mem[795][5] ), .S(n8418), .Z(n5335)
         );
  MUX2_X1 U24290 ( .A(\mem[792][5] ), .B(\mem[793][5] ), .S(n8418), .Z(n5336)
         );
  MUX2_X1 U24291 ( .A(n5336), .B(n5335), .S(n8296), .Z(n5337) );
  MUX2_X1 U24292 ( .A(n5337), .B(n5334), .S(n8247), .Z(n5338) );
  MUX2_X1 U24293 ( .A(\mem[790][5] ), .B(\mem[791][5] ), .S(n8418), .Z(n5339)
         );
  MUX2_X1 U24294 ( .A(\mem[788][5] ), .B(\mem[789][5] ), .S(n8418), .Z(n5340)
         );
  MUX2_X1 U24295 ( .A(n5340), .B(n5339), .S(n8296), .Z(n5341) );
  MUX2_X1 U24296 ( .A(\mem[786][5] ), .B(\mem[787][5] ), .S(n8418), .Z(n5342)
         );
  MUX2_X1 U24297 ( .A(\mem[784][5] ), .B(\mem[785][5] ), .S(n8418), .Z(n5343)
         );
  MUX2_X1 U24298 ( .A(n5343), .B(n5342), .S(n8296), .Z(n5344) );
  MUX2_X1 U24299 ( .A(n5344), .B(n5341), .S(n8248), .Z(n5345) );
  MUX2_X1 U24300 ( .A(n5345), .B(n5338), .S(n8204), .Z(n5346) );
  MUX2_X1 U24301 ( .A(\mem[782][5] ), .B(\mem[783][5] ), .S(n8419), .Z(n5347)
         );
  MUX2_X1 U24302 ( .A(\mem[780][5] ), .B(\mem[781][5] ), .S(n8419), .Z(n5348)
         );
  MUX2_X1 U24303 ( .A(n5348), .B(n5347), .S(n8297), .Z(n5349) );
  MUX2_X1 U24304 ( .A(\mem[778][5] ), .B(\mem[779][5] ), .S(n8419), .Z(n5350)
         );
  MUX2_X1 U24305 ( .A(\mem[776][5] ), .B(\mem[777][5] ), .S(n8419), .Z(n5351)
         );
  MUX2_X1 U24306 ( .A(n5351), .B(n5350), .S(n8297), .Z(n5352) );
  MUX2_X1 U24307 ( .A(n5352), .B(n5349), .S(n8249), .Z(n5353) );
  MUX2_X1 U24308 ( .A(\mem[774][5] ), .B(\mem[775][5] ), .S(n8419), .Z(n5354)
         );
  MUX2_X1 U24309 ( .A(\mem[772][5] ), .B(\mem[773][5] ), .S(n8419), .Z(n5355)
         );
  MUX2_X1 U24310 ( .A(n5355), .B(n5354), .S(n8297), .Z(n5356) );
  MUX2_X1 U24311 ( .A(\mem[770][5] ), .B(\mem[771][5] ), .S(n8419), .Z(n5357)
         );
  MUX2_X1 U24312 ( .A(\mem[768][5] ), .B(\mem[769][5] ), .S(n8419), .Z(n5358)
         );
  MUX2_X1 U24313 ( .A(n5358), .B(n5357), .S(n8297), .Z(n5359) );
  MUX2_X1 U24314 ( .A(n5359), .B(n5356), .S(n8244), .Z(n5360) );
  MUX2_X1 U24315 ( .A(n5360), .B(n5353), .S(n8204), .Z(n5361) );
  MUX2_X1 U24316 ( .A(n5361), .B(n5346), .S(n8192), .Z(n5362) );
  MUX2_X1 U24317 ( .A(n5362), .B(n5331), .S(n8182), .Z(n5363) );
  MUX2_X1 U24318 ( .A(n5363), .B(n5300), .S(n8178), .Z(n5364) );
  MUX2_X1 U24319 ( .A(n5364), .B(n5237), .S(N25), .Z(n5365) );
  MUX2_X1 U24320 ( .A(\mem[766][5] ), .B(\mem[767][5] ), .S(n8419), .Z(n5366)
         );
  MUX2_X1 U24321 ( .A(\mem[764][5] ), .B(\mem[765][5] ), .S(n8419), .Z(n5367)
         );
  MUX2_X1 U24322 ( .A(n5367), .B(n5366), .S(n8297), .Z(n5368) );
  MUX2_X1 U24323 ( .A(\mem[762][5] ), .B(\mem[763][5] ), .S(n8419), .Z(n5369)
         );
  MUX2_X1 U24324 ( .A(\mem[760][5] ), .B(\mem[761][5] ), .S(n8419), .Z(n5370)
         );
  MUX2_X1 U24325 ( .A(n5370), .B(n5369), .S(n8297), .Z(n5371) );
  MUX2_X1 U24326 ( .A(n5371), .B(n5368), .S(n8245), .Z(n5372) );
  MUX2_X1 U24327 ( .A(\mem[758][5] ), .B(\mem[759][5] ), .S(n8420), .Z(n5373)
         );
  MUX2_X1 U24328 ( .A(\mem[756][5] ), .B(\mem[757][5] ), .S(n8420), .Z(n5374)
         );
  MUX2_X1 U24329 ( .A(n5374), .B(n5373), .S(n8297), .Z(n5375) );
  MUX2_X1 U24330 ( .A(\mem[754][5] ), .B(\mem[755][5] ), .S(n8420), .Z(n5376)
         );
  MUX2_X1 U24331 ( .A(\mem[752][5] ), .B(\mem[753][5] ), .S(n8420), .Z(n5377)
         );
  MUX2_X1 U24332 ( .A(n5377), .B(n5376), .S(n8297), .Z(n5378) );
  MUX2_X1 U24333 ( .A(n5378), .B(n5375), .S(n8246), .Z(n5379) );
  MUX2_X1 U24334 ( .A(n5379), .B(n5372), .S(n8204), .Z(n5380) );
  MUX2_X1 U24335 ( .A(\mem[750][5] ), .B(\mem[751][5] ), .S(n8420), .Z(n5381)
         );
  MUX2_X1 U24336 ( .A(\mem[748][5] ), .B(\mem[749][5] ), .S(n8420), .Z(n5382)
         );
  MUX2_X1 U24337 ( .A(n5382), .B(n5381), .S(n8297), .Z(n5383) );
  MUX2_X1 U24338 ( .A(\mem[746][5] ), .B(\mem[747][5] ), .S(n8420), .Z(n5384)
         );
  MUX2_X1 U24339 ( .A(\mem[744][5] ), .B(\mem[745][5] ), .S(n8420), .Z(n5385)
         );
  MUX2_X1 U24340 ( .A(n5385), .B(n5384), .S(n8297), .Z(n5386) );
  MUX2_X1 U24341 ( .A(n5386), .B(n5383), .S(n8253), .Z(n5387) );
  MUX2_X1 U24342 ( .A(\mem[742][5] ), .B(\mem[743][5] ), .S(n8420), .Z(n5388)
         );
  MUX2_X1 U24343 ( .A(\mem[740][5] ), .B(\mem[741][5] ), .S(n8420), .Z(n5389)
         );
  MUX2_X1 U24344 ( .A(n5389), .B(n5388), .S(n8297), .Z(n5390) );
  MUX2_X1 U24345 ( .A(\mem[738][5] ), .B(\mem[739][5] ), .S(n8420), .Z(n5391)
         );
  MUX2_X1 U24346 ( .A(\mem[736][5] ), .B(\mem[737][5] ), .S(n8420), .Z(n5392)
         );
  MUX2_X1 U24347 ( .A(n5392), .B(n5391), .S(n8297), .Z(n5393) );
  MUX2_X1 U24348 ( .A(n5393), .B(n5390), .S(n8254), .Z(n5394) );
  MUX2_X1 U24349 ( .A(n5394), .B(n5387), .S(n8204), .Z(n5395) );
  MUX2_X1 U24350 ( .A(n5395), .B(n5380), .S(n8191), .Z(n5396) );
  MUX2_X1 U24351 ( .A(\mem[734][5] ), .B(\mem[735][5] ), .S(n8421), .Z(n5397)
         );
  MUX2_X1 U24352 ( .A(\mem[732][5] ), .B(\mem[733][5] ), .S(n8421), .Z(n5398)
         );
  MUX2_X1 U24353 ( .A(n5398), .B(n5397), .S(n8298), .Z(n5399) );
  MUX2_X1 U24354 ( .A(\mem[730][5] ), .B(\mem[731][5] ), .S(n8421), .Z(n5400)
         );
  MUX2_X1 U24355 ( .A(\mem[728][5] ), .B(\mem[729][5] ), .S(n8421), .Z(n5401)
         );
  MUX2_X1 U24356 ( .A(n5401), .B(n5400), .S(n8298), .Z(n5402) );
  MUX2_X1 U24357 ( .A(n5402), .B(n5399), .S(n8232), .Z(n5403) );
  MUX2_X1 U24358 ( .A(\mem[726][5] ), .B(\mem[727][5] ), .S(n8421), .Z(n5404)
         );
  MUX2_X1 U24359 ( .A(\mem[724][5] ), .B(\mem[725][5] ), .S(n8421), .Z(n5405)
         );
  MUX2_X1 U24360 ( .A(n5405), .B(n5404), .S(n8298), .Z(n5406) );
  MUX2_X1 U24361 ( .A(\mem[722][5] ), .B(\mem[723][5] ), .S(n8421), .Z(n5407)
         );
  MUX2_X1 U24362 ( .A(\mem[720][5] ), .B(\mem[721][5] ), .S(n8421), .Z(n5408)
         );
  MUX2_X1 U24363 ( .A(n5408), .B(n5407), .S(n8298), .Z(n5409) );
  MUX2_X1 U24364 ( .A(n5409), .B(n5406), .S(n8233), .Z(n5410) );
  MUX2_X1 U24365 ( .A(n5410), .B(n5403), .S(n8204), .Z(n5411) );
  MUX2_X1 U24366 ( .A(\mem[718][5] ), .B(\mem[719][5] ), .S(n8421), .Z(n5412)
         );
  MUX2_X1 U24367 ( .A(\mem[716][5] ), .B(\mem[717][5] ), .S(n8421), .Z(n5413)
         );
  MUX2_X1 U24368 ( .A(n5413), .B(n5412), .S(n8298), .Z(n5414) );
  MUX2_X1 U24369 ( .A(\mem[714][5] ), .B(\mem[715][5] ), .S(n8421), .Z(n5415)
         );
  MUX2_X1 U24370 ( .A(\mem[712][5] ), .B(\mem[713][5] ), .S(n8421), .Z(n5416)
         );
  MUX2_X1 U24371 ( .A(n5416), .B(n5415), .S(n8298), .Z(n5417) );
  MUX2_X1 U24372 ( .A(n5417), .B(n5414), .S(n8234), .Z(n5418) );
  MUX2_X1 U24373 ( .A(\mem[710][5] ), .B(\mem[711][5] ), .S(n8422), .Z(n5419)
         );
  MUX2_X1 U24374 ( .A(\mem[708][5] ), .B(\mem[709][5] ), .S(n8422), .Z(n5420)
         );
  MUX2_X1 U24375 ( .A(n5420), .B(n5419), .S(n8298), .Z(n5421) );
  MUX2_X1 U24376 ( .A(\mem[706][5] ), .B(\mem[707][5] ), .S(n8422), .Z(n5422)
         );
  MUX2_X1 U24377 ( .A(\mem[704][5] ), .B(\mem[705][5] ), .S(n8422), .Z(n5423)
         );
  MUX2_X1 U24378 ( .A(n5423), .B(n5422), .S(n8298), .Z(n5424) );
  MUX2_X1 U24379 ( .A(n5424), .B(n5421), .S(n8241), .Z(n5425) );
  MUX2_X1 U24380 ( .A(n5425), .B(n5418), .S(n8204), .Z(n5426) );
  MUX2_X1 U24381 ( .A(n5426), .B(n5411), .S(N22), .Z(n5427) );
  MUX2_X1 U24382 ( .A(n5427), .B(n5396), .S(n8185), .Z(n5428) );
  MUX2_X1 U24383 ( .A(\mem[702][5] ), .B(\mem[703][5] ), .S(n8422), .Z(n5429)
         );
  MUX2_X1 U24384 ( .A(\mem[700][5] ), .B(\mem[701][5] ), .S(n8422), .Z(n5430)
         );
  MUX2_X1 U24385 ( .A(n5430), .B(n5429), .S(n8298), .Z(n5431) );
  MUX2_X1 U24386 ( .A(\mem[698][5] ), .B(\mem[699][5] ), .S(n8422), .Z(n5432)
         );
  MUX2_X1 U24387 ( .A(\mem[696][5] ), .B(\mem[697][5] ), .S(n8422), .Z(n5433)
         );
  MUX2_X1 U24388 ( .A(n5433), .B(n5432), .S(n8298), .Z(n5434) );
  MUX2_X1 U24389 ( .A(n5434), .B(n5431), .S(n8242), .Z(n5435) );
  MUX2_X1 U24390 ( .A(\mem[694][5] ), .B(\mem[695][5] ), .S(n8422), .Z(n5436)
         );
  MUX2_X1 U24391 ( .A(\mem[692][5] ), .B(\mem[693][5] ), .S(n8422), .Z(n5437)
         );
  MUX2_X1 U24392 ( .A(n5437), .B(n5436), .S(n8298), .Z(n5438) );
  MUX2_X1 U24393 ( .A(\mem[690][5] ), .B(\mem[691][5] ), .S(n8422), .Z(n5439)
         );
  MUX2_X1 U24394 ( .A(\mem[688][5] ), .B(\mem[689][5] ), .S(n8422), .Z(n5440)
         );
  MUX2_X1 U24395 ( .A(n5440), .B(n5439), .S(n8298), .Z(n5441) );
  MUX2_X1 U24396 ( .A(n5441), .B(n5438), .S(n8243), .Z(n5442) );
  MUX2_X1 U24397 ( .A(n5442), .B(n5435), .S(n8204), .Z(n5443) );
  MUX2_X1 U24398 ( .A(\mem[686][5] ), .B(\mem[687][5] ), .S(n8423), .Z(n5444)
         );
  MUX2_X1 U24399 ( .A(\mem[684][5] ), .B(\mem[685][5] ), .S(n8423), .Z(n5445)
         );
  MUX2_X1 U24400 ( .A(n5445), .B(n5444), .S(n8299), .Z(n5446) );
  MUX2_X1 U24401 ( .A(\mem[682][5] ), .B(\mem[683][5] ), .S(n8423), .Z(n5447)
         );
  MUX2_X1 U24402 ( .A(\mem[680][5] ), .B(\mem[681][5] ), .S(n8423), .Z(n5448)
         );
  MUX2_X1 U24403 ( .A(n5448), .B(n5447), .S(n8299), .Z(n5449) );
  MUX2_X1 U24404 ( .A(n5449), .B(n5446), .S(n8238), .Z(n5450) );
  MUX2_X1 U24405 ( .A(\mem[678][5] ), .B(\mem[679][5] ), .S(n8423), .Z(n5451)
         );
  MUX2_X1 U24406 ( .A(\mem[676][5] ), .B(\mem[677][5] ), .S(n8423), .Z(n5452)
         );
  MUX2_X1 U24407 ( .A(n5452), .B(n5451), .S(n8299), .Z(n5453) );
  MUX2_X1 U24408 ( .A(\mem[674][5] ), .B(\mem[675][5] ), .S(n8423), .Z(n5454)
         );
  MUX2_X1 U24409 ( .A(\mem[672][5] ), .B(\mem[673][5] ), .S(n8423), .Z(n5455)
         );
  MUX2_X1 U24410 ( .A(n5455), .B(n5454), .S(n8299), .Z(n5456) );
  MUX2_X1 U24411 ( .A(n5456), .B(n5453), .S(n8239), .Z(n5457) );
  MUX2_X1 U24412 ( .A(n5457), .B(n5450), .S(n8204), .Z(n5458) );
  MUX2_X1 U24413 ( .A(n5458), .B(n5443), .S(n8194), .Z(n5459) );
  MUX2_X1 U24414 ( .A(\mem[670][5] ), .B(\mem[671][5] ), .S(n8423), .Z(n5460)
         );
  MUX2_X1 U24415 ( .A(\mem[668][5] ), .B(\mem[669][5] ), .S(n8423), .Z(n5461)
         );
  MUX2_X1 U24416 ( .A(n5461), .B(n5460), .S(n8299), .Z(n5462) );
  MUX2_X1 U24417 ( .A(\mem[666][5] ), .B(\mem[667][5] ), .S(n8423), .Z(n5463)
         );
  MUX2_X1 U24418 ( .A(\mem[664][5] ), .B(\mem[665][5] ), .S(n8423), .Z(n5464)
         );
  MUX2_X1 U24419 ( .A(n5464), .B(n5463), .S(n8299), .Z(n5465) );
  MUX2_X1 U24420 ( .A(n5465), .B(n5462), .S(n8240), .Z(n5466) );
  MUX2_X1 U24421 ( .A(\mem[662][5] ), .B(\mem[663][5] ), .S(n8424), .Z(n5467)
         );
  MUX2_X1 U24422 ( .A(\mem[660][5] ), .B(\mem[661][5] ), .S(n8424), .Z(n5468)
         );
  MUX2_X1 U24423 ( .A(n5468), .B(n5467), .S(n8299), .Z(n5469) );
  MUX2_X1 U24424 ( .A(\mem[658][5] ), .B(\mem[659][5] ), .S(n8424), .Z(n5470)
         );
  MUX2_X1 U24425 ( .A(\mem[656][5] ), .B(\mem[657][5] ), .S(n8424), .Z(n5471)
         );
  MUX2_X1 U24426 ( .A(n5471), .B(n5470), .S(n8299), .Z(n5472) );
  MUX2_X1 U24427 ( .A(n5472), .B(n5469), .S(n8230), .Z(n5473) );
  MUX2_X1 U24428 ( .A(n5473), .B(n5466), .S(n8204), .Z(n5474) );
  MUX2_X1 U24429 ( .A(\mem[654][5] ), .B(\mem[655][5] ), .S(n8424), .Z(n5475)
         );
  MUX2_X1 U24430 ( .A(\mem[652][5] ), .B(\mem[653][5] ), .S(n8424), .Z(n5476)
         );
  MUX2_X1 U24431 ( .A(n5476), .B(n5475), .S(n8299), .Z(n5477) );
  MUX2_X1 U24432 ( .A(\mem[650][5] ), .B(\mem[651][5] ), .S(n8424), .Z(n5478)
         );
  MUX2_X1 U24433 ( .A(\mem[648][5] ), .B(\mem[649][5] ), .S(n8424), .Z(n5479)
         );
  MUX2_X1 U24434 ( .A(n5479), .B(n5478), .S(n8299), .Z(n5480) );
  MUX2_X1 U24435 ( .A(n5480), .B(n5477), .S(n8231), .Z(n5481) );
  MUX2_X1 U24436 ( .A(\mem[646][5] ), .B(\mem[647][5] ), .S(n8424), .Z(n5482)
         );
  MUX2_X1 U24437 ( .A(\mem[644][5] ), .B(\mem[645][5] ), .S(n8424), .Z(n5483)
         );
  MUX2_X1 U24438 ( .A(n5483), .B(n5482), .S(n8299), .Z(n5484) );
  MUX2_X1 U24439 ( .A(\mem[642][5] ), .B(\mem[643][5] ), .S(n8424), .Z(n5485)
         );
  MUX2_X1 U24440 ( .A(\mem[640][5] ), .B(\mem[641][5] ), .S(n8424), .Z(n5486)
         );
  MUX2_X1 U24441 ( .A(n5486), .B(n5485), .S(n8299), .Z(n5487) );
  MUX2_X1 U24442 ( .A(n5487), .B(n5484), .S(n8227), .Z(n5488) );
  MUX2_X1 U24443 ( .A(n5488), .B(n5481), .S(n8204), .Z(n5489) );
  MUX2_X1 U24444 ( .A(n5489), .B(n5474), .S(n8195), .Z(n5490) );
  MUX2_X1 U24445 ( .A(n5490), .B(n5459), .S(n8183), .Z(n5491) );
  MUX2_X1 U24446 ( .A(n5491), .B(n5428), .S(n8178), .Z(n5492) );
  MUX2_X1 U24447 ( .A(\mem[638][5] ), .B(\mem[639][5] ), .S(n8425), .Z(n5493)
         );
  MUX2_X1 U24448 ( .A(\mem[636][5] ), .B(\mem[637][5] ), .S(n8425), .Z(n5494)
         );
  MUX2_X1 U24449 ( .A(n5494), .B(n5493), .S(n8300), .Z(n5495) );
  MUX2_X1 U24450 ( .A(\mem[634][5] ), .B(\mem[635][5] ), .S(n8425), .Z(n5496)
         );
  MUX2_X1 U24451 ( .A(\mem[632][5] ), .B(\mem[633][5] ), .S(n8425), .Z(n5497)
         );
  MUX2_X1 U24452 ( .A(n5497), .B(n5496), .S(n8300), .Z(n5498) );
  MUX2_X1 U24453 ( .A(n5498), .B(n5495), .S(n8236), .Z(n5499) );
  MUX2_X1 U24454 ( .A(\mem[630][5] ), .B(\mem[631][5] ), .S(n8425), .Z(n5500)
         );
  MUX2_X1 U24455 ( .A(\mem[628][5] ), .B(\mem[629][5] ), .S(n8425), .Z(n5501)
         );
  MUX2_X1 U24456 ( .A(n5501), .B(n5500), .S(n8300), .Z(n5502) );
  MUX2_X1 U24457 ( .A(\mem[626][5] ), .B(\mem[627][5] ), .S(n8425), .Z(n5503)
         );
  MUX2_X1 U24458 ( .A(\mem[624][5] ), .B(\mem[625][5] ), .S(n8425), .Z(n5504)
         );
  MUX2_X1 U24459 ( .A(n5504), .B(n5503), .S(n8300), .Z(n5505) );
  MUX2_X1 U24460 ( .A(n5505), .B(n5502), .S(n8261), .Z(n5506) );
  MUX2_X1 U24461 ( .A(n5506), .B(n5499), .S(n8205), .Z(n5507) );
  MUX2_X1 U24462 ( .A(\mem[622][5] ), .B(\mem[623][5] ), .S(n8425), .Z(n5508)
         );
  MUX2_X1 U24463 ( .A(\mem[620][5] ), .B(\mem[621][5] ), .S(n8425), .Z(n5509)
         );
  MUX2_X1 U24464 ( .A(n5509), .B(n5508), .S(n8300), .Z(n5510) );
  MUX2_X1 U24465 ( .A(\mem[618][5] ), .B(\mem[619][5] ), .S(n8425), .Z(n5511)
         );
  MUX2_X1 U24466 ( .A(\mem[616][5] ), .B(\mem[617][5] ), .S(n8425), .Z(n5512)
         );
  MUX2_X1 U24467 ( .A(n5512), .B(n5511), .S(n8300), .Z(n5513) );
  MUX2_X1 U24468 ( .A(n5513), .B(n5510), .S(n8235), .Z(n5514) );
  MUX2_X1 U24469 ( .A(\mem[614][5] ), .B(\mem[615][5] ), .S(n8426), .Z(n5515)
         );
  MUX2_X1 U24470 ( .A(\mem[612][5] ), .B(\mem[613][5] ), .S(n8426), .Z(n5516)
         );
  MUX2_X1 U24471 ( .A(n5516), .B(n5515), .S(n8300), .Z(n5517) );
  MUX2_X1 U24472 ( .A(\mem[610][5] ), .B(\mem[611][5] ), .S(n8426), .Z(n5518)
         );
  MUX2_X1 U24473 ( .A(\mem[608][5] ), .B(\mem[609][5] ), .S(n8426), .Z(n5519)
         );
  MUX2_X1 U24474 ( .A(n5519), .B(n5518), .S(n8300), .Z(n5520) );
  MUX2_X1 U24475 ( .A(n5520), .B(n5517), .S(n8252), .Z(n5521) );
  MUX2_X1 U24476 ( .A(n5521), .B(n5514), .S(n8205), .Z(n5522) );
  MUX2_X1 U24477 ( .A(n5522), .B(n5507), .S(n8189), .Z(n5523) );
  MUX2_X1 U24478 ( .A(\mem[606][5] ), .B(\mem[607][5] ), .S(n8426), .Z(n5524)
         );
  MUX2_X1 U24479 ( .A(\mem[604][5] ), .B(\mem[605][5] ), .S(n8426), .Z(n5525)
         );
  MUX2_X1 U24480 ( .A(n5525), .B(n5524), .S(n8300), .Z(n5526) );
  MUX2_X1 U24481 ( .A(\mem[602][5] ), .B(\mem[603][5] ), .S(n8426), .Z(n5527)
         );
  MUX2_X1 U24482 ( .A(\mem[600][5] ), .B(\mem[601][5] ), .S(n8426), .Z(n5528)
         );
  MUX2_X1 U24483 ( .A(n5528), .B(n5527), .S(n8300), .Z(n5529) );
  MUX2_X1 U24484 ( .A(n5529), .B(n5526), .S(n8228), .Z(n5530) );
  MUX2_X1 U24485 ( .A(\mem[598][5] ), .B(\mem[599][5] ), .S(n8426), .Z(n5531)
         );
  MUX2_X1 U24486 ( .A(\mem[596][5] ), .B(\mem[597][5] ), .S(n8426), .Z(n5532)
         );
  MUX2_X1 U24487 ( .A(n5532), .B(n5531), .S(n8300), .Z(n5533) );
  MUX2_X1 U24488 ( .A(\mem[594][5] ), .B(\mem[595][5] ), .S(n8426), .Z(n5534)
         );
  MUX2_X1 U24489 ( .A(\mem[592][5] ), .B(\mem[593][5] ), .S(n8426), .Z(n5535)
         );
  MUX2_X1 U24490 ( .A(n5535), .B(n5534), .S(n8300), .Z(n5536) );
  MUX2_X1 U24491 ( .A(n5536), .B(n5533), .S(n8227), .Z(n5537) );
  MUX2_X1 U24492 ( .A(n5537), .B(n5530), .S(n8205), .Z(n5538) );
  MUX2_X1 U24493 ( .A(\mem[590][5] ), .B(\mem[591][5] ), .S(n8427), .Z(n5539)
         );
  MUX2_X1 U24494 ( .A(\mem[588][5] ), .B(\mem[589][5] ), .S(n8427), .Z(n5540)
         );
  MUX2_X1 U24495 ( .A(n5540), .B(n5539), .S(n8301), .Z(n5541) );
  MUX2_X1 U24496 ( .A(\mem[586][5] ), .B(\mem[587][5] ), .S(n8427), .Z(n5542)
         );
  MUX2_X1 U24497 ( .A(\mem[584][5] ), .B(\mem[585][5] ), .S(n8427), .Z(n5543)
         );
  MUX2_X1 U24498 ( .A(n5543), .B(n5542), .S(n8301), .Z(n5544) );
  MUX2_X1 U24499 ( .A(n5544), .B(n5541), .S(n8235), .Z(n5545) );
  MUX2_X1 U24500 ( .A(\mem[582][5] ), .B(\mem[583][5] ), .S(n8427), .Z(n5546)
         );
  MUX2_X1 U24501 ( .A(\mem[580][5] ), .B(\mem[581][5] ), .S(n8427), .Z(n5547)
         );
  MUX2_X1 U24502 ( .A(n5547), .B(n5546), .S(n8301), .Z(n5548) );
  MUX2_X1 U24503 ( .A(\mem[578][5] ), .B(\mem[579][5] ), .S(n8427), .Z(n5549)
         );
  MUX2_X1 U24504 ( .A(\mem[576][5] ), .B(\mem[577][5] ), .S(n8427), .Z(n5550)
         );
  MUX2_X1 U24505 ( .A(n5550), .B(n5549), .S(n8301), .Z(n5551) );
  MUX2_X1 U24506 ( .A(n5551), .B(n5548), .S(n8264), .Z(n5552) );
  MUX2_X1 U24507 ( .A(n5552), .B(n5545), .S(n8205), .Z(n5553) );
  MUX2_X1 U24508 ( .A(n5553), .B(n5538), .S(n8189), .Z(n5554) );
  MUX2_X1 U24509 ( .A(n5554), .B(n5523), .S(n8185), .Z(n5555) );
  MUX2_X1 U24510 ( .A(\mem[574][5] ), .B(\mem[575][5] ), .S(n8427), .Z(n5556)
         );
  MUX2_X1 U24511 ( .A(\mem[572][5] ), .B(\mem[573][5] ), .S(n8427), .Z(n5557)
         );
  MUX2_X1 U24512 ( .A(n5557), .B(n5556), .S(n8301), .Z(n5558) );
  MUX2_X1 U24513 ( .A(\mem[570][5] ), .B(\mem[571][5] ), .S(n8427), .Z(n5559)
         );
  MUX2_X1 U24514 ( .A(\mem[568][5] ), .B(\mem[569][5] ), .S(n8427), .Z(n5560)
         );
  MUX2_X1 U24515 ( .A(n5560), .B(n5559), .S(n8301), .Z(n5561) );
  MUX2_X1 U24516 ( .A(n5561), .B(n5558), .S(n8247), .Z(n5562) );
  MUX2_X1 U24517 ( .A(\mem[566][5] ), .B(\mem[567][5] ), .S(n8428), .Z(n5563)
         );
  MUX2_X1 U24518 ( .A(\mem[564][5] ), .B(\mem[565][5] ), .S(n8428), .Z(n5564)
         );
  MUX2_X1 U24519 ( .A(n5564), .B(n5563), .S(n8301), .Z(n5565) );
  MUX2_X1 U24520 ( .A(\mem[562][5] ), .B(\mem[563][5] ), .S(n8428), .Z(n5566)
         );
  MUX2_X1 U24521 ( .A(\mem[560][5] ), .B(\mem[561][5] ), .S(n8428), .Z(n5567)
         );
  MUX2_X1 U24522 ( .A(n5567), .B(n5566), .S(n8301), .Z(n5568) );
  MUX2_X1 U24523 ( .A(n5568), .B(n5565), .S(n8222), .Z(n5569) );
  MUX2_X1 U24524 ( .A(n5569), .B(n5562), .S(n8205), .Z(n5570) );
  MUX2_X1 U24525 ( .A(\mem[558][5] ), .B(\mem[559][5] ), .S(n8428), .Z(n5571)
         );
  MUX2_X1 U24526 ( .A(\mem[556][5] ), .B(\mem[557][5] ), .S(n8428), .Z(n5572)
         );
  MUX2_X1 U24527 ( .A(n5572), .B(n5571), .S(n8301), .Z(n5573) );
  MUX2_X1 U24528 ( .A(\mem[554][5] ), .B(\mem[555][5] ), .S(n8428), .Z(n5574)
         );
  MUX2_X1 U24529 ( .A(\mem[552][5] ), .B(\mem[553][5] ), .S(n8428), .Z(n5575)
         );
  MUX2_X1 U24530 ( .A(n5575), .B(n5574), .S(n8301), .Z(n5576) );
  MUX2_X1 U24531 ( .A(n5576), .B(n5573), .S(n8243), .Z(n5577) );
  MUX2_X1 U24532 ( .A(\mem[550][5] ), .B(\mem[551][5] ), .S(n8428), .Z(n5578)
         );
  MUX2_X1 U24533 ( .A(\mem[548][5] ), .B(\mem[549][5] ), .S(n8428), .Z(n5579)
         );
  MUX2_X1 U24534 ( .A(n5579), .B(n5578), .S(n8301), .Z(n5580) );
  MUX2_X1 U24535 ( .A(\mem[546][5] ), .B(\mem[547][5] ), .S(n8428), .Z(n5581)
         );
  MUX2_X1 U24536 ( .A(\mem[544][5] ), .B(\mem[545][5] ), .S(n8428), .Z(n5582)
         );
  MUX2_X1 U24537 ( .A(n5582), .B(n5581), .S(n8301), .Z(n5583) );
  MUX2_X1 U24538 ( .A(n5583), .B(n5580), .S(n8235), .Z(n5584) );
  MUX2_X1 U24539 ( .A(n5584), .B(n5577), .S(n8205), .Z(n5585) );
  MUX2_X1 U24540 ( .A(n5585), .B(n5570), .S(n8189), .Z(n5586) );
  MUX2_X1 U24541 ( .A(\mem[542][5] ), .B(\mem[543][5] ), .S(n8429), .Z(n5587)
         );
  MUX2_X1 U24542 ( .A(\mem[540][5] ), .B(\mem[541][5] ), .S(n8429), .Z(n5588)
         );
  MUX2_X1 U24543 ( .A(n5588), .B(n5587), .S(n8302), .Z(n5589) );
  MUX2_X1 U24544 ( .A(\mem[538][5] ), .B(\mem[539][5] ), .S(n8429), .Z(n5590)
         );
  MUX2_X1 U24545 ( .A(\mem[536][5] ), .B(\mem[537][5] ), .S(n8429), .Z(n5591)
         );
  MUX2_X1 U24546 ( .A(n5591), .B(n5590), .S(n8302), .Z(n5592) );
  MUX2_X1 U24547 ( .A(n5592), .B(n5589), .S(n8224), .Z(n5593) );
  MUX2_X1 U24548 ( .A(\mem[534][5] ), .B(\mem[535][5] ), .S(n8429), .Z(n5594)
         );
  MUX2_X1 U24549 ( .A(\mem[532][5] ), .B(\mem[533][5] ), .S(n8429), .Z(n5595)
         );
  MUX2_X1 U24550 ( .A(n5595), .B(n5594), .S(n8302), .Z(n5596) );
  MUX2_X1 U24551 ( .A(\mem[530][5] ), .B(\mem[531][5] ), .S(n8429), .Z(n5597)
         );
  MUX2_X1 U24552 ( .A(\mem[528][5] ), .B(\mem[529][5] ), .S(n8429), .Z(n5598)
         );
  MUX2_X1 U24553 ( .A(n5598), .B(n5597), .S(n8302), .Z(n5599) );
  MUX2_X1 U24554 ( .A(n5599), .B(n5596), .S(n8223), .Z(n5600) );
  MUX2_X1 U24555 ( .A(n5600), .B(n5593), .S(n8205), .Z(n5601) );
  MUX2_X1 U24556 ( .A(\mem[526][5] ), .B(\mem[527][5] ), .S(n8429), .Z(n5602)
         );
  MUX2_X1 U24557 ( .A(\mem[524][5] ), .B(\mem[525][5] ), .S(n8429), .Z(n5603)
         );
  MUX2_X1 U24558 ( .A(n5603), .B(n5602), .S(n8302), .Z(n5604) );
  MUX2_X1 U24559 ( .A(\mem[522][5] ), .B(\mem[523][5] ), .S(n8429), .Z(n5605)
         );
  MUX2_X1 U24560 ( .A(\mem[520][5] ), .B(\mem[521][5] ), .S(n8429), .Z(n5606)
         );
  MUX2_X1 U24561 ( .A(n5606), .B(n5605), .S(n8302), .Z(n5607) );
  MUX2_X1 U24562 ( .A(n5607), .B(n5604), .S(n8236), .Z(n5608) );
  MUX2_X1 U24563 ( .A(\mem[518][5] ), .B(\mem[519][5] ), .S(n8430), .Z(n5609)
         );
  MUX2_X1 U24564 ( .A(\mem[516][5] ), .B(\mem[517][5] ), .S(n8430), .Z(n5610)
         );
  MUX2_X1 U24565 ( .A(n5610), .B(n5609), .S(n8302), .Z(n5611) );
  MUX2_X1 U24566 ( .A(\mem[514][5] ), .B(\mem[515][5] ), .S(n8430), .Z(n5612)
         );
  MUX2_X1 U24567 ( .A(\mem[512][5] ), .B(\mem[513][5] ), .S(n8430), .Z(n5613)
         );
  MUX2_X1 U24568 ( .A(n5613), .B(n5612), .S(n8302), .Z(n5614) );
  MUX2_X1 U24569 ( .A(n5614), .B(n5611), .S(n8263), .Z(n5615) );
  MUX2_X1 U24570 ( .A(n5615), .B(n5608), .S(n8205), .Z(n5616) );
  MUX2_X1 U24571 ( .A(n5616), .B(n5601), .S(n8189), .Z(n5617) );
  MUX2_X1 U24572 ( .A(n5617), .B(n5586), .S(n8184), .Z(n5618) );
  MUX2_X1 U24573 ( .A(n5618), .B(n5555), .S(n8178), .Z(n5619) );
  MUX2_X1 U24574 ( .A(n5619), .B(n5492), .S(n8177), .Z(n5620) );
  MUX2_X1 U24575 ( .A(n5620), .B(n5365), .S(N26), .Z(n5621) );
  MUX2_X1 U24576 ( .A(\mem[510][5] ), .B(\mem[511][5] ), .S(n8430), .Z(n5622)
         );
  MUX2_X1 U24577 ( .A(\mem[508][5] ), .B(\mem[509][5] ), .S(n8430), .Z(n5623)
         );
  MUX2_X1 U24578 ( .A(n5623), .B(n5622), .S(n8302), .Z(n5624) );
  MUX2_X1 U24579 ( .A(\mem[506][5] ), .B(\mem[507][5] ), .S(n8430), .Z(n5625)
         );
  MUX2_X1 U24580 ( .A(\mem[504][5] ), .B(\mem[505][5] ), .S(n8430), .Z(n5626)
         );
  MUX2_X1 U24581 ( .A(n5626), .B(n5625), .S(n8302), .Z(n5627) );
  MUX2_X1 U24582 ( .A(n5627), .B(n5624), .S(n8222), .Z(n5628) );
  MUX2_X1 U24583 ( .A(\mem[502][5] ), .B(\mem[503][5] ), .S(n8430), .Z(n5629)
         );
  MUX2_X1 U24584 ( .A(\mem[500][5] ), .B(\mem[501][5] ), .S(n8430), .Z(n5630)
         );
  MUX2_X1 U24585 ( .A(n5630), .B(n5629), .S(n8302), .Z(n5631) );
  MUX2_X1 U24586 ( .A(\mem[498][5] ), .B(\mem[499][5] ), .S(n8430), .Z(n5632)
         );
  MUX2_X1 U24587 ( .A(\mem[496][5] ), .B(\mem[497][5] ), .S(n8430), .Z(n5633)
         );
  MUX2_X1 U24588 ( .A(n5633), .B(n5632), .S(n8302), .Z(n5634) );
  MUX2_X1 U24589 ( .A(n5634), .B(n5631), .S(n8221), .Z(n5635) );
  MUX2_X1 U24590 ( .A(n5635), .B(n5628), .S(n8205), .Z(n5636) );
  MUX2_X1 U24591 ( .A(\mem[494][5] ), .B(\mem[495][5] ), .S(n8431), .Z(n5637)
         );
  MUX2_X1 U24592 ( .A(\mem[492][5] ), .B(\mem[493][5] ), .S(n8431), .Z(n5638)
         );
  MUX2_X1 U24593 ( .A(n5638), .B(n5637), .S(n8303), .Z(n5639) );
  MUX2_X1 U24594 ( .A(\mem[490][5] ), .B(\mem[491][5] ), .S(n8431), .Z(n5640)
         );
  MUX2_X1 U24595 ( .A(\mem[488][5] ), .B(\mem[489][5] ), .S(n8431), .Z(n5641)
         );
  MUX2_X1 U24596 ( .A(n5641), .B(n5640), .S(n8303), .Z(n5642) );
  MUX2_X1 U24597 ( .A(n5642), .B(n5639), .S(n8220), .Z(n5643) );
  MUX2_X1 U24598 ( .A(\mem[486][5] ), .B(\mem[487][5] ), .S(n8431), .Z(n5644)
         );
  MUX2_X1 U24599 ( .A(\mem[484][5] ), .B(\mem[485][5] ), .S(n8431), .Z(n5645)
         );
  MUX2_X1 U24600 ( .A(n5645), .B(n5644), .S(n8303), .Z(n5646) );
  MUX2_X1 U24601 ( .A(\mem[482][5] ), .B(\mem[483][5] ), .S(n8431), .Z(n5647)
         );
  MUX2_X1 U24602 ( .A(\mem[480][5] ), .B(\mem[481][5] ), .S(n8431), .Z(n5648)
         );
  MUX2_X1 U24603 ( .A(n5648), .B(n5647), .S(n8303), .Z(n5649) );
  MUX2_X1 U24604 ( .A(n5649), .B(n5646), .S(n8236), .Z(n5650) );
  MUX2_X1 U24605 ( .A(n5650), .B(n5643), .S(n8205), .Z(n5651) );
  MUX2_X1 U24606 ( .A(n5651), .B(n5636), .S(n8189), .Z(n5652) );
  MUX2_X1 U24607 ( .A(\mem[478][5] ), .B(\mem[479][5] ), .S(n8431), .Z(n5653)
         );
  MUX2_X1 U24608 ( .A(\mem[476][5] ), .B(\mem[477][5] ), .S(n8431), .Z(n5654)
         );
  MUX2_X1 U24609 ( .A(n5654), .B(n5653), .S(n8303), .Z(n5655) );
  MUX2_X1 U24610 ( .A(\mem[474][5] ), .B(\mem[475][5] ), .S(n8431), .Z(n5656)
         );
  MUX2_X1 U24611 ( .A(\mem[472][5] ), .B(\mem[473][5] ), .S(n8431), .Z(n5657)
         );
  MUX2_X1 U24612 ( .A(n5657), .B(n5656), .S(n8303), .Z(n5658) );
  MUX2_X1 U24613 ( .A(n5658), .B(n5655), .S(n8258), .Z(n5659) );
  MUX2_X1 U24614 ( .A(\mem[470][5] ), .B(\mem[471][5] ), .S(n8432), .Z(n5660)
         );
  MUX2_X1 U24615 ( .A(\mem[468][5] ), .B(\mem[469][5] ), .S(n8432), .Z(n5661)
         );
  MUX2_X1 U24616 ( .A(n5661), .B(n5660), .S(n8303), .Z(n5662) );
  MUX2_X1 U24617 ( .A(\mem[466][5] ), .B(\mem[467][5] ), .S(n8432), .Z(n5663)
         );
  MUX2_X1 U24618 ( .A(\mem[464][5] ), .B(\mem[465][5] ), .S(n8432), .Z(n5664)
         );
  MUX2_X1 U24619 ( .A(n5664), .B(n5663), .S(n8303), .Z(n5665) );
  MUX2_X1 U24620 ( .A(n5665), .B(n5662), .S(n8228), .Z(n5666) );
  MUX2_X1 U24621 ( .A(n5666), .B(n5659), .S(n8205), .Z(n5667) );
  MUX2_X1 U24622 ( .A(\mem[462][5] ), .B(\mem[463][5] ), .S(n8432), .Z(n5668)
         );
  MUX2_X1 U24623 ( .A(\mem[460][5] ), .B(\mem[461][5] ), .S(n8432), .Z(n5669)
         );
  MUX2_X1 U24624 ( .A(n5669), .B(n5668), .S(n8303), .Z(n5670) );
  MUX2_X1 U24625 ( .A(\mem[458][5] ), .B(\mem[459][5] ), .S(n8432), .Z(n5671)
         );
  MUX2_X1 U24626 ( .A(\mem[456][5] ), .B(\mem[457][5] ), .S(n8432), .Z(n5672)
         );
  MUX2_X1 U24627 ( .A(n5672), .B(n5671), .S(n8303), .Z(n5673) );
  MUX2_X1 U24628 ( .A(n5673), .B(n5670), .S(n8236), .Z(n5674) );
  MUX2_X1 U24629 ( .A(\mem[454][5] ), .B(\mem[455][5] ), .S(n8432), .Z(n5675)
         );
  MUX2_X1 U24630 ( .A(\mem[452][5] ), .B(\mem[453][5] ), .S(n8432), .Z(n5676)
         );
  MUX2_X1 U24631 ( .A(n5676), .B(n5675), .S(n8303), .Z(n5677) );
  MUX2_X1 U24632 ( .A(\mem[450][5] ), .B(\mem[451][5] ), .S(n8432), .Z(n5678)
         );
  MUX2_X1 U24633 ( .A(\mem[448][5] ), .B(\mem[449][5] ), .S(n8432), .Z(n5679)
         );
  MUX2_X1 U24634 ( .A(n5679), .B(n5678), .S(n8303), .Z(n5680) );
  MUX2_X1 U24635 ( .A(n5680), .B(n5677), .S(n8221), .Z(n5681) );
  MUX2_X1 U24636 ( .A(n5681), .B(n5674), .S(n8205), .Z(n5682) );
  MUX2_X1 U24637 ( .A(n5682), .B(n5667), .S(n8189), .Z(n5683) );
  MUX2_X1 U24638 ( .A(n5683), .B(n5652), .S(n8185), .Z(n5684) );
  MUX2_X1 U24639 ( .A(\mem[446][5] ), .B(\mem[447][5] ), .S(n8433), .Z(n5685)
         );
  MUX2_X1 U24640 ( .A(\mem[444][5] ), .B(\mem[445][5] ), .S(n8433), .Z(n5686)
         );
  MUX2_X1 U24641 ( .A(n5686), .B(n5685), .S(n8304), .Z(n5687) );
  MUX2_X1 U24642 ( .A(\mem[442][5] ), .B(\mem[443][5] ), .S(n8433), .Z(n5688)
         );
  MUX2_X1 U24643 ( .A(\mem[440][5] ), .B(\mem[441][5] ), .S(n8433), .Z(n5689)
         );
  MUX2_X1 U24644 ( .A(n5689), .B(n5688), .S(n8304), .Z(n5690) );
  MUX2_X1 U24645 ( .A(n5690), .B(n5687), .S(n8261), .Z(n5691) );
  MUX2_X1 U24646 ( .A(\mem[438][5] ), .B(\mem[439][5] ), .S(n8433), .Z(n5692)
         );
  MUX2_X1 U24647 ( .A(\mem[436][5] ), .B(\mem[437][5] ), .S(n8433), .Z(n5693)
         );
  MUX2_X1 U24648 ( .A(n5693), .B(n5692), .S(n8304), .Z(n5694) );
  MUX2_X1 U24649 ( .A(\mem[434][5] ), .B(\mem[435][5] ), .S(n8433), .Z(n5695)
         );
  MUX2_X1 U24650 ( .A(\mem[432][5] ), .B(\mem[433][5] ), .S(n8433), .Z(n5696)
         );
  MUX2_X1 U24651 ( .A(n5696), .B(n5695), .S(n8304), .Z(n5697) );
  MUX2_X1 U24652 ( .A(n5697), .B(n5694), .S(n8224), .Z(n5698) );
  MUX2_X1 U24653 ( .A(n5698), .B(n5691), .S(n8206), .Z(n5699) );
  MUX2_X1 U24654 ( .A(\mem[430][5] ), .B(\mem[431][5] ), .S(n8433), .Z(n5700)
         );
  MUX2_X1 U24655 ( .A(\mem[428][5] ), .B(\mem[429][5] ), .S(n8433), .Z(n5701)
         );
  MUX2_X1 U24656 ( .A(n5701), .B(n5700), .S(n8304), .Z(n5702) );
  MUX2_X1 U24657 ( .A(\mem[426][5] ), .B(\mem[427][5] ), .S(n8433), .Z(n5703)
         );
  MUX2_X1 U24658 ( .A(\mem[424][5] ), .B(\mem[425][5] ), .S(n8433), .Z(n5704)
         );
  MUX2_X1 U24659 ( .A(n5704), .B(n5703), .S(n8304), .Z(n5705) );
  MUX2_X1 U24660 ( .A(n5705), .B(n5702), .S(n8262), .Z(n5706) );
  MUX2_X1 U24661 ( .A(\mem[422][5] ), .B(\mem[423][5] ), .S(n8434), .Z(n5707)
         );
  MUX2_X1 U24662 ( .A(\mem[420][5] ), .B(\mem[421][5] ), .S(n8434), .Z(n5708)
         );
  MUX2_X1 U24663 ( .A(n5708), .B(n5707), .S(n8304), .Z(n5709) );
  MUX2_X1 U24664 ( .A(\mem[418][5] ), .B(\mem[419][5] ), .S(n8434), .Z(n5710)
         );
  MUX2_X1 U24665 ( .A(\mem[416][5] ), .B(\mem[417][5] ), .S(n8434), .Z(n5711)
         );
  MUX2_X1 U24666 ( .A(n5711), .B(n5710), .S(n8304), .Z(n5712) );
  MUX2_X1 U24667 ( .A(n5712), .B(n5709), .S(n8251), .Z(n5713) );
  MUX2_X1 U24668 ( .A(n5713), .B(n5706), .S(n8206), .Z(n5714) );
  MUX2_X1 U24669 ( .A(n5714), .B(n5699), .S(n8189), .Z(n5715) );
  MUX2_X1 U24670 ( .A(\mem[414][5] ), .B(\mem[415][5] ), .S(n8434), .Z(n5716)
         );
  MUX2_X1 U24671 ( .A(\mem[412][5] ), .B(\mem[413][5] ), .S(n8434), .Z(n5717)
         );
  MUX2_X1 U24672 ( .A(n5717), .B(n5716), .S(n8304), .Z(n5718) );
  MUX2_X1 U24673 ( .A(\mem[410][5] ), .B(\mem[411][5] ), .S(n8434), .Z(n5719)
         );
  MUX2_X1 U24674 ( .A(\mem[408][5] ), .B(\mem[409][5] ), .S(n8434), .Z(n5720)
         );
  MUX2_X1 U24675 ( .A(n5720), .B(n5719), .S(n8304), .Z(n5721) );
  MUX2_X1 U24676 ( .A(n5721), .B(n5718), .S(n8262), .Z(n5722) );
  MUX2_X1 U24677 ( .A(\mem[406][5] ), .B(\mem[407][5] ), .S(n8434), .Z(n5723)
         );
  MUX2_X1 U24678 ( .A(\mem[404][5] ), .B(\mem[405][5] ), .S(n8434), .Z(n5724)
         );
  MUX2_X1 U24679 ( .A(n5724), .B(n5723), .S(n8304), .Z(n5725) );
  MUX2_X1 U24680 ( .A(\mem[402][5] ), .B(\mem[403][5] ), .S(n8434), .Z(n5726)
         );
  MUX2_X1 U24681 ( .A(\mem[400][5] ), .B(\mem[401][5] ), .S(n8434), .Z(n5727)
         );
  MUX2_X1 U24682 ( .A(n5727), .B(n5726), .S(n8304), .Z(n5728) );
  MUX2_X1 U24683 ( .A(n5728), .B(n5725), .S(n8222), .Z(n5729) );
  MUX2_X1 U24684 ( .A(n5729), .B(n5722), .S(n8206), .Z(n5730) );
  MUX2_X1 U24685 ( .A(\mem[398][5] ), .B(\mem[399][5] ), .S(n8435), .Z(n5731)
         );
  MUX2_X1 U24686 ( .A(\mem[396][5] ), .B(\mem[397][5] ), .S(n8435), .Z(n5732)
         );
  MUX2_X1 U24687 ( .A(n5732), .B(n5731), .S(n8305), .Z(n5733) );
  MUX2_X1 U24688 ( .A(\mem[394][5] ), .B(\mem[395][5] ), .S(n8435), .Z(n5734)
         );
  MUX2_X1 U24689 ( .A(\mem[392][5] ), .B(\mem[393][5] ), .S(n8435), .Z(n5735)
         );
  MUX2_X1 U24690 ( .A(n5735), .B(n5734), .S(n8305), .Z(n5736) );
  MUX2_X1 U24691 ( .A(n5736), .B(n5733), .S(n8225), .Z(n5737) );
  MUX2_X1 U24692 ( .A(\mem[390][5] ), .B(\mem[391][5] ), .S(n8435), .Z(n5738)
         );
  MUX2_X1 U24693 ( .A(\mem[388][5] ), .B(\mem[389][5] ), .S(n8435), .Z(n5739)
         );
  MUX2_X1 U24694 ( .A(n5739), .B(n5738), .S(n8305), .Z(n5740) );
  MUX2_X1 U24695 ( .A(\mem[386][5] ), .B(\mem[387][5] ), .S(n8435), .Z(n5741)
         );
  MUX2_X1 U24696 ( .A(\mem[384][5] ), .B(\mem[385][5] ), .S(n8435), .Z(n5742)
         );
  MUX2_X1 U24697 ( .A(n5742), .B(n5741), .S(n8305), .Z(n5743) );
  MUX2_X1 U24698 ( .A(n5743), .B(n5740), .S(n8234), .Z(n5744) );
  MUX2_X1 U24699 ( .A(n5744), .B(n5737), .S(n8206), .Z(n5745) );
  MUX2_X1 U24700 ( .A(n5745), .B(n5730), .S(n8189), .Z(n5746) );
  MUX2_X1 U24701 ( .A(n5746), .B(n5715), .S(n8183), .Z(n5747) );
  MUX2_X1 U24702 ( .A(n5747), .B(n5684), .S(n8178), .Z(n5748) );
  MUX2_X1 U24703 ( .A(\mem[382][5] ), .B(\mem[383][5] ), .S(n8435), .Z(n5749)
         );
  MUX2_X1 U24704 ( .A(\mem[380][5] ), .B(\mem[381][5] ), .S(n8435), .Z(n5750)
         );
  MUX2_X1 U24705 ( .A(n5750), .B(n5749), .S(n8305), .Z(n5751) );
  MUX2_X1 U24706 ( .A(\mem[378][5] ), .B(\mem[379][5] ), .S(n8435), .Z(n5752)
         );
  MUX2_X1 U24707 ( .A(\mem[376][5] ), .B(\mem[377][5] ), .S(n8435), .Z(n5753)
         );
  MUX2_X1 U24708 ( .A(n5753), .B(n5752), .S(n8305), .Z(n5754) );
  MUX2_X1 U24709 ( .A(n5754), .B(n5751), .S(n8242), .Z(n5755) );
  MUX2_X1 U24710 ( .A(\mem[374][5] ), .B(\mem[375][5] ), .S(n8436), .Z(n5756)
         );
  MUX2_X1 U24711 ( .A(\mem[372][5] ), .B(\mem[373][5] ), .S(n8436), .Z(n5757)
         );
  MUX2_X1 U24712 ( .A(n5757), .B(n5756), .S(n8305), .Z(n5758) );
  MUX2_X1 U24713 ( .A(\mem[370][5] ), .B(\mem[371][5] ), .S(n8436), .Z(n5759)
         );
  MUX2_X1 U24714 ( .A(\mem[368][5] ), .B(\mem[369][5] ), .S(n8436), .Z(n5760)
         );
  MUX2_X1 U24715 ( .A(n5760), .B(n5759), .S(n8305), .Z(n5761) );
  MUX2_X1 U24716 ( .A(n5761), .B(n5758), .S(n8248), .Z(n5762) );
  MUX2_X1 U24717 ( .A(n5762), .B(n5755), .S(n8206), .Z(n5763) );
  MUX2_X1 U24718 ( .A(\mem[366][5] ), .B(\mem[367][5] ), .S(n8436), .Z(n5764)
         );
  MUX2_X1 U24719 ( .A(\mem[364][5] ), .B(\mem[365][5] ), .S(n8436), .Z(n5765)
         );
  MUX2_X1 U24720 ( .A(n5765), .B(n5764), .S(n8305), .Z(n5766) );
  MUX2_X1 U24721 ( .A(\mem[362][5] ), .B(\mem[363][5] ), .S(n8436), .Z(n5767)
         );
  MUX2_X1 U24722 ( .A(\mem[360][5] ), .B(\mem[361][5] ), .S(n8436), .Z(n5768)
         );
  MUX2_X1 U24723 ( .A(n5768), .B(n5767), .S(n8305), .Z(n5769) );
  MUX2_X1 U24724 ( .A(n5769), .B(n5766), .S(N20), .Z(n5770) );
  MUX2_X1 U24725 ( .A(\mem[358][5] ), .B(\mem[359][5] ), .S(n8436), .Z(n5771)
         );
  MUX2_X1 U24726 ( .A(\mem[356][5] ), .B(\mem[357][5] ), .S(n8436), .Z(n5772)
         );
  MUX2_X1 U24727 ( .A(n5772), .B(n5771), .S(n8305), .Z(n5773) );
  MUX2_X1 U24728 ( .A(\mem[354][5] ), .B(\mem[355][5] ), .S(n8436), .Z(n5774)
         );
  MUX2_X1 U24729 ( .A(\mem[352][5] ), .B(\mem[353][5] ), .S(n8436), .Z(n5775)
         );
  MUX2_X1 U24730 ( .A(n5775), .B(n5774), .S(n8305), .Z(n5776) );
  MUX2_X1 U24731 ( .A(n5776), .B(n5773), .S(n8263), .Z(n5777) );
  MUX2_X1 U24732 ( .A(n5777), .B(n5770), .S(n8206), .Z(n5778) );
  MUX2_X1 U24733 ( .A(n5778), .B(n5763), .S(n8189), .Z(n5779) );
  MUX2_X1 U24734 ( .A(\mem[350][5] ), .B(\mem[351][5] ), .S(n8437), .Z(n5780)
         );
  MUX2_X1 U24735 ( .A(\mem[348][5] ), .B(\mem[349][5] ), .S(n8437), .Z(n5781)
         );
  MUX2_X1 U24736 ( .A(n5781), .B(n5780), .S(n8306), .Z(n5782) );
  MUX2_X1 U24737 ( .A(\mem[346][5] ), .B(\mem[347][5] ), .S(n8437), .Z(n5783)
         );
  MUX2_X1 U24738 ( .A(\mem[344][5] ), .B(\mem[345][5] ), .S(n8437), .Z(n5784)
         );
  MUX2_X1 U24739 ( .A(n5784), .B(n5783), .S(n8306), .Z(n5785) );
  MUX2_X1 U24740 ( .A(n5785), .B(n5782), .S(n8260), .Z(n5786) );
  MUX2_X1 U24741 ( .A(\mem[342][5] ), .B(\mem[343][5] ), .S(n8437), .Z(n5787)
         );
  MUX2_X1 U24742 ( .A(\mem[340][5] ), .B(\mem[341][5] ), .S(n8437), .Z(n5788)
         );
  MUX2_X1 U24743 ( .A(n5788), .B(n5787), .S(n8306), .Z(n5789) );
  MUX2_X1 U24744 ( .A(\mem[338][5] ), .B(\mem[339][5] ), .S(n8437), .Z(n5790)
         );
  MUX2_X1 U24745 ( .A(\mem[336][5] ), .B(\mem[337][5] ), .S(n8437), .Z(n5791)
         );
  MUX2_X1 U24746 ( .A(n5791), .B(n5790), .S(n8306), .Z(n5792) );
  MUX2_X1 U24747 ( .A(n5792), .B(n5789), .S(n8252), .Z(n5793) );
  MUX2_X1 U24748 ( .A(n5793), .B(n5786), .S(n8206), .Z(n5794) );
  MUX2_X1 U24749 ( .A(\mem[334][5] ), .B(\mem[335][5] ), .S(n8437), .Z(n5795)
         );
  MUX2_X1 U24750 ( .A(\mem[332][5] ), .B(\mem[333][5] ), .S(n8437), .Z(n5796)
         );
  MUX2_X1 U24751 ( .A(n5796), .B(n5795), .S(n8306), .Z(n5797) );
  MUX2_X1 U24752 ( .A(\mem[330][5] ), .B(\mem[331][5] ), .S(n8437), .Z(n5798)
         );
  MUX2_X1 U24753 ( .A(\mem[328][5] ), .B(\mem[329][5] ), .S(n8437), .Z(n5799)
         );
  MUX2_X1 U24754 ( .A(n5799), .B(n5798), .S(n8306), .Z(n5800) );
  MUX2_X1 U24755 ( .A(n5800), .B(n5797), .S(n8259), .Z(n5801) );
  MUX2_X1 U24756 ( .A(\mem[326][5] ), .B(\mem[327][5] ), .S(n8438), .Z(n5802)
         );
  MUX2_X1 U24757 ( .A(\mem[324][5] ), .B(\mem[325][5] ), .S(n8438), .Z(n5803)
         );
  MUX2_X1 U24758 ( .A(n5803), .B(n5802), .S(n8306), .Z(n5804) );
  MUX2_X1 U24759 ( .A(\mem[322][5] ), .B(\mem[323][5] ), .S(n8438), .Z(n5805)
         );
  MUX2_X1 U24760 ( .A(\mem[320][5] ), .B(\mem[321][5] ), .S(n8438), .Z(n5806)
         );
  MUX2_X1 U24761 ( .A(n5806), .B(n5805), .S(n8306), .Z(n5807) );
  MUX2_X1 U24762 ( .A(n5807), .B(n5804), .S(n8260), .Z(n5808) );
  MUX2_X1 U24763 ( .A(n5808), .B(n5801), .S(n8206), .Z(n5809) );
  MUX2_X1 U24764 ( .A(n5809), .B(n5794), .S(n8189), .Z(n5810) );
  MUX2_X1 U24765 ( .A(n5810), .B(n5779), .S(N23), .Z(n5811) );
  MUX2_X1 U24766 ( .A(\mem[318][5] ), .B(\mem[319][5] ), .S(n8438), .Z(n5812)
         );
  MUX2_X1 U24767 ( .A(\mem[316][5] ), .B(\mem[317][5] ), .S(n8438), .Z(n5813)
         );
  MUX2_X1 U24768 ( .A(n5813), .B(n5812), .S(n8306), .Z(n5814) );
  MUX2_X1 U24769 ( .A(\mem[314][5] ), .B(\mem[315][5] ), .S(n8438), .Z(n5815)
         );
  MUX2_X1 U24770 ( .A(\mem[312][5] ), .B(\mem[313][5] ), .S(n8438), .Z(n5816)
         );
  MUX2_X1 U24771 ( .A(n5816), .B(n5815), .S(n8306), .Z(n5817) );
  MUX2_X1 U24772 ( .A(n5817), .B(n5814), .S(n8226), .Z(n5818) );
  MUX2_X1 U24773 ( .A(\mem[310][5] ), .B(\mem[311][5] ), .S(n8438), .Z(n5819)
         );
  MUX2_X1 U24774 ( .A(\mem[308][5] ), .B(\mem[309][5] ), .S(n8438), .Z(n5820)
         );
  MUX2_X1 U24775 ( .A(n5820), .B(n5819), .S(n8306), .Z(n5821) );
  MUX2_X1 U24776 ( .A(\mem[306][5] ), .B(\mem[307][5] ), .S(n8438), .Z(n5822)
         );
  MUX2_X1 U24777 ( .A(\mem[304][5] ), .B(\mem[305][5] ), .S(n8438), .Z(n5823)
         );
  MUX2_X1 U24778 ( .A(n5823), .B(n5822), .S(n8306), .Z(n5824) );
  MUX2_X1 U24779 ( .A(n5824), .B(n5821), .S(n8223), .Z(n5825) );
  MUX2_X1 U24780 ( .A(n5825), .B(n5818), .S(n8206), .Z(n5826) );
  MUX2_X1 U24781 ( .A(\mem[302][5] ), .B(\mem[303][5] ), .S(n8439), .Z(n5827)
         );
  MUX2_X1 U24782 ( .A(\mem[300][5] ), .B(\mem[301][5] ), .S(n8439), .Z(n5828)
         );
  MUX2_X1 U24783 ( .A(n5828), .B(n5827), .S(n8307), .Z(n5829) );
  MUX2_X1 U24784 ( .A(\mem[298][5] ), .B(\mem[299][5] ), .S(n8439), .Z(n5830)
         );
  MUX2_X1 U24785 ( .A(\mem[296][5] ), .B(\mem[297][5] ), .S(n8439), .Z(n5831)
         );
  MUX2_X1 U24786 ( .A(n5831), .B(n5830), .S(n8307), .Z(n5832) );
  MUX2_X1 U24787 ( .A(n5832), .B(n5829), .S(n8242), .Z(n5833) );
  MUX2_X1 U24788 ( .A(\mem[294][5] ), .B(\mem[295][5] ), .S(n8439), .Z(n5834)
         );
  MUX2_X1 U24789 ( .A(\mem[292][5] ), .B(\mem[293][5] ), .S(n8439), .Z(n5835)
         );
  MUX2_X1 U24790 ( .A(n5835), .B(n5834), .S(n8307), .Z(n5836) );
  MUX2_X1 U24791 ( .A(\mem[290][5] ), .B(\mem[291][5] ), .S(n8439), .Z(n5837)
         );
  MUX2_X1 U24792 ( .A(\mem[288][5] ), .B(\mem[289][5] ), .S(n8439), .Z(n5838)
         );
  MUX2_X1 U24793 ( .A(n5838), .B(n5837), .S(n8307), .Z(n5839) );
  MUX2_X1 U24794 ( .A(n5839), .B(n5836), .S(n8256), .Z(n5840) );
  MUX2_X1 U24795 ( .A(n5840), .B(n5833), .S(n8206), .Z(n5841) );
  MUX2_X1 U24796 ( .A(n5841), .B(n5826), .S(n8189), .Z(n5842) );
  MUX2_X1 U24797 ( .A(\mem[286][5] ), .B(\mem[287][5] ), .S(n8439), .Z(n5843)
         );
  MUX2_X1 U24798 ( .A(\mem[284][5] ), .B(\mem[285][5] ), .S(n8439), .Z(n5844)
         );
  MUX2_X1 U24799 ( .A(n5844), .B(n5843), .S(n8307), .Z(n5845) );
  MUX2_X1 U24800 ( .A(\mem[282][5] ), .B(\mem[283][5] ), .S(n8439), .Z(n5846)
         );
  MUX2_X1 U24801 ( .A(\mem[280][5] ), .B(\mem[281][5] ), .S(n8439), .Z(n5847)
         );
  MUX2_X1 U24802 ( .A(n5847), .B(n5846), .S(n8307), .Z(n5848) );
  MUX2_X1 U24803 ( .A(n5848), .B(n5845), .S(n8257), .Z(n5849) );
  MUX2_X1 U24804 ( .A(\mem[278][5] ), .B(\mem[279][5] ), .S(n8440), .Z(n5850)
         );
  MUX2_X1 U24805 ( .A(\mem[276][5] ), .B(\mem[277][5] ), .S(n8440), .Z(n5851)
         );
  MUX2_X1 U24806 ( .A(n5851), .B(n5850), .S(n8307), .Z(n5852) );
  MUX2_X1 U24807 ( .A(\mem[274][5] ), .B(\mem[275][5] ), .S(n8440), .Z(n5853)
         );
  MUX2_X1 U24808 ( .A(\mem[272][5] ), .B(\mem[273][5] ), .S(n8440), .Z(n5854)
         );
  MUX2_X1 U24809 ( .A(n5854), .B(n5853), .S(n8307), .Z(n5855) );
  MUX2_X1 U24810 ( .A(n5855), .B(n5852), .S(n8258), .Z(n5856) );
  MUX2_X1 U24811 ( .A(n5856), .B(n5849), .S(n8206), .Z(n5857) );
  MUX2_X1 U24812 ( .A(\mem[270][5] ), .B(\mem[271][5] ), .S(n8440), .Z(n5858)
         );
  MUX2_X1 U24813 ( .A(\mem[268][5] ), .B(\mem[269][5] ), .S(n8440), .Z(n5859)
         );
  MUX2_X1 U24814 ( .A(n5859), .B(n5858), .S(n8307), .Z(n5860) );
  MUX2_X1 U24815 ( .A(\mem[266][5] ), .B(\mem[267][5] ), .S(n8440), .Z(n5861)
         );
  MUX2_X1 U24816 ( .A(\mem[264][5] ), .B(\mem[265][5] ), .S(n8440), .Z(n5862)
         );
  MUX2_X1 U24817 ( .A(n5862), .B(n5861), .S(n8307), .Z(n5863) );
  MUX2_X1 U24818 ( .A(n5863), .B(n5860), .S(n8243), .Z(n5864) );
  MUX2_X1 U24819 ( .A(\mem[262][5] ), .B(\mem[263][5] ), .S(n8440), .Z(n5865)
         );
  MUX2_X1 U24820 ( .A(\mem[260][5] ), .B(\mem[261][5] ), .S(n8440), .Z(n5866)
         );
  MUX2_X1 U24821 ( .A(n5866), .B(n5865), .S(n8307), .Z(n5867) );
  MUX2_X1 U24822 ( .A(\mem[258][5] ), .B(\mem[259][5] ), .S(n8440), .Z(n5868)
         );
  MUX2_X1 U24823 ( .A(\mem[256][5] ), .B(\mem[257][5] ), .S(n8440), .Z(n5869)
         );
  MUX2_X1 U24824 ( .A(n5869), .B(n5868), .S(n8307), .Z(n5870) );
  MUX2_X1 U24825 ( .A(n5870), .B(n5867), .S(n8264), .Z(n5871) );
  MUX2_X1 U24826 ( .A(n5871), .B(n5864), .S(n8206), .Z(n5872) );
  MUX2_X1 U24827 ( .A(n5872), .B(n5857), .S(n8189), .Z(n5873) );
  MUX2_X1 U24828 ( .A(n5873), .B(n5842), .S(n8185), .Z(n5874) );
  MUX2_X1 U24829 ( .A(n5874), .B(n5811), .S(n8178), .Z(n5875) );
  MUX2_X1 U24830 ( .A(n5875), .B(n5748), .S(N25), .Z(n5876) );
  MUX2_X1 U24831 ( .A(\mem[254][5] ), .B(\mem[255][5] ), .S(n8441), .Z(n5877)
         );
  MUX2_X1 U24832 ( .A(\mem[252][5] ), .B(\mem[253][5] ), .S(n8441), .Z(n5878)
         );
  MUX2_X1 U24833 ( .A(n5878), .B(n5877), .S(n8308), .Z(n5879) );
  MUX2_X1 U24834 ( .A(\mem[250][5] ), .B(\mem[251][5] ), .S(n8441), .Z(n5880)
         );
  MUX2_X1 U24835 ( .A(\mem[248][5] ), .B(\mem[249][5] ), .S(n8441), .Z(n5881)
         );
  MUX2_X1 U24836 ( .A(n5881), .B(n5880), .S(n8308), .Z(n5882) );
  MUX2_X1 U24837 ( .A(n5882), .B(n5879), .S(n8226), .Z(n5883) );
  MUX2_X1 U24838 ( .A(\mem[246][5] ), .B(\mem[247][5] ), .S(n8441), .Z(n5884)
         );
  MUX2_X1 U24839 ( .A(\mem[244][5] ), .B(\mem[245][5] ), .S(n8441), .Z(n5885)
         );
  MUX2_X1 U24840 ( .A(n5885), .B(n5884), .S(n8308), .Z(n5886) );
  MUX2_X1 U24841 ( .A(\mem[242][5] ), .B(\mem[243][5] ), .S(n8441), .Z(n5887)
         );
  MUX2_X1 U24842 ( .A(\mem[240][5] ), .B(\mem[241][5] ), .S(n8441), .Z(n5888)
         );
  MUX2_X1 U24843 ( .A(n5888), .B(n5887), .S(n8308), .Z(n5889) );
  MUX2_X1 U24844 ( .A(n5889), .B(n5886), .S(n8247), .Z(n5890) );
  MUX2_X1 U24845 ( .A(n5890), .B(n5883), .S(n8207), .Z(n5891) );
  MUX2_X1 U24846 ( .A(\mem[238][5] ), .B(\mem[239][5] ), .S(n8441), .Z(n5892)
         );
  MUX2_X1 U24847 ( .A(\mem[236][5] ), .B(\mem[237][5] ), .S(n8441), .Z(n5893)
         );
  MUX2_X1 U24848 ( .A(n5893), .B(n5892), .S(n8308), .Z(n5894) );
  MUX2_X1 U24849 ( .A(\mem[234][5] ), .B(\mem[235][5] ), .S(n8441), .Z(n5895)
         );
  MUX2_X1 U24850 ( .A(\mem[232][5] ), .B(\mem[233][5] ), .S(n8441), .Z(n5896)
         );
  MUX2_X1 U24851 ( .A(n5896), .B(n5895), .S(n8308), .Z(n5897) );
  MUX2_X1 U24852 ( .A(n5897), .B(n5894), .S(n8248), .Z(n5898) );
  MUX2_X1 U24853 ( .A(\mem[230][5] ), .B(\mem[231][5] ), .S(n8442), .Z(n5899)
         );
  MUX2_X1 U24854 ( .A(\mem[228][5] ), .B(\mem[229][5] ), .S(n8442), .Z(n5900)
         );
  MUX2_X1 U24855 ( .A(n5900), .B(n5899), .S(n8308), .Z(n5901) );
  MUX2_X1 U24856 ( .A(\mem[226][5] ), .B(\mem[227][5] ), .S(n8442), .Z(n5902)
         );
  MUX2_X1 U24857 ( .A(\mem[224][5] ), .B(\mem[225][5] ), .S(n8442), .Z(n5903)
         );
  MUX2_X1 U24858 ( .A(n5903), .B(n5902), .S(n8308), .Z(n5904) );
  MUX2_X1 U24859 ( .A(n5904), .B(n5901), .S(n8249), .Z(n5905) );
  MUX2_X1 U24860 ( .A(n5905), .B(n5898), .S(n8207), .Z(n5906) );
  MUX2_X1 U24861 ( .A(n5906), .B(n5891), .S(n8190), .Z(n5907) );
  MUX2_X1 U24862 ( .A(\mem[222][5] ), .B(\mem[223][5] ), .S(n8442), .Z(n5908)
         );
  MUX2_X1 U24863 ( .A(\mem[220][5] ), .B(\mem[221][5] ), .S(n8442), .Z(n5909)
         );
  MUX2_X1 U24864 ( .A(n5909), .B(n5908), .S(n8308), .Z(n5910) );
  MUX2_X1 U24865 ( .A(\mem[218][5] ), .B(\mem[219][5] ), .S(n8442), .Z(n5911)
         );
  MUX2_X1 U24866 ( .A(\mem[216][5] ), .B(\mem[217][5] ), .S(n8442), .Z(n5912)
         );
  MUX2_X1 U24867 ( .A(n5912), .B(n5911), .S(n8308), .Z(n5913) );
  MUX2_X1 U24868 ( .A(n5913), .B(n5910), .S(n8244), .Z(n5914) );
  MUX2_X1 U24869 ( .A(\mem[214][5] ), .B(\mem[215][5] ), .S(n8442), .Z(n5915)
         );
  MUX2_X1 U24870 ( .A(\mem[212][5] ), .B(\mem[213][5] ), .S(n8442), .Z(n5916)
         );
  MUX2_X1 U24871 ( .A(n5916), .B(n5915), .S(n8308), .Z(n5917) );
  MUX2_X1 U24872 ( .A(\mem[210][5] ), .B(\mem[211][5] ), .S(n8442), .Z(n5918)
         );
  MUX2_X1 U24873 ( .A(\mem[208][5] ), .B(\mem[209][5] ), .S(n8442), .Z(n5919)
         );
  MUX2_X1 U24874 ( .A(n5919), .B(n5918), .S(n8308), .Z(n5920) );
  MUX2_X1 U24875 ( .A(n5920), .B(n5917), .S(n8245), .Z(n5921) );
  MUX2_X1 U24876 ( .A(n5921), .B(n5914), .S(n8207), .Z(n5922) );
  MUX2_X1 U24877 ( .A(\mem[206][5] ), .B(\mem[207][5] ), .S(n8443), .Z(n5923)
         );
  MUX2_X1 U24878 ( .A(\mem[204][5] ), .B(\mem[205][5] ), .S(n8443), .Z(n5924)
         );
  MUX2_X1 U24879 ( .A(n5924), .B(n5923), .S(n8309), .Z(n5925) );
  MUX2_X1 U24880 ( .A(\mem[202][5] ), .B(\mem[203][5] ), .S(n8443), .Z(n5926)
         );
  MUX2_X1 U24881 ( .A(\mem[200][5] ), .B(\mem[201][5] ), .S(n8443), .Z(n5927)
         );
  MUX2_X1 U24882 ( .A(n5927), .B(n5926), .S(n8309), .Z(n5928) );
  MUX2_X1 U24883 ( .A(n5928), .B(n5925), .S(n8246), .Z(n5929) );
  MUX2_X1 U24884 ( .A(\mem[198][5] ), .B(\mem[199][5] ), .S(n8443), .Z(n5930)
         );
  MUX2_X1 U24885 ( .A(\mem[196][5] ), .B(\mem[197][5] ), .S(n8443), .Z(n5931)
         );
  MUX2_X1 U24886 ( .A(n5931), .B(n5930), .S(n8309), .Z(n5932) );
  MUX2_X1 U24887 ( .A(\mem[194][5] ), .B(\mem[195][5] ), .S(n8443), .Z(n5933)
         );
  MUX2_X1 U24888 ( .A(\mem[192][5] ), .B(\mem[193][5] ), .S(n8443), .Z(n5934)
         );
  MUX2_X1 U24889 ( .A(n5934), .B(n5933), .S(n8309), .Z(n5935) );
  MUX2_X1 U24890 ( .A(n5935), .B(n5932), .S(n8253), .Z(n5936) );
  MUX2_X1 U24891 ( .A(n5936), .B(n5929), .S(n8207), .Z(n5937) );
  MUX2_X1 U24892 ( .A(n5937), .B(n5922), .S(n8190), .Z(n5938) );
  MUX2_X1 U24893 ( .A(n5938), .B(n5907), .S(n8183), .Z(n5939) );
  MUX2_X1 U24894 ( .A(\mem[190][5] ), .B(\mem[191][5] ), .S(n8443), .Z(n5940)
         );
  MUX2_X1 U24895 ( .A(\mem[188][5] ), .B(\mem[189][5] ), .S(n8443), .Z(n5941)
         );
  MUX2_X1 U24896 ( .A(n5941), .B(n5940), .S(n8309), .Z(n5942) );
  MUX2_X1 U24897 ( .A(\mem[186][5] ), .B(\mem[187][5] ), .S(n8443), .Z(n5943)
         );
  MUX2_X1 U24898 ( .A(\mem[184][5] ), .B(\mem[185][5] ), .S(n8443), .Z(n5944)
         );
  MUX2_X1 U24899 ( .A(n5944), .B(n5943), .S(n8309), .Z(n5945) );
  MUX2_X1 U24900 ( .A(n5945), .B(n5942), .S(n8254), .Z(n5946) );
  MUX2_X1 U24901 ( .A(\mem[182][5] ), .B(\mem[183][5] ), .S(n8444), .Z(n5947)
         );
  MUX2_X1 U24902 ( .A(\mem[180][5] ), .B(\mem[181][5] ), .S(n8444), .Z(n5948)
         );
  MUX2_X1 U24903 ( .A(n5948), .B(n5947), .S(n8309), .Z(n5949) );
  MUX2_X1 U24904 ( .A(\mem[178][5] ), .B(\mem[179][5] ), .S(n8444), .Z(n5950)
         );
  MUX2_X1 U24905 ( .A(\mem[176][5] ), .B(\mem[177][5] ), .S(n8444), .Z(n5951)
         );
  MUX2_X1 U24906 ( .A(n5951), .B(n5950), .S(n8309), .Z(n5952) );
  MUX2_X1 U24907 ( .A(n5952), .B(n5949), .S(n8255), .Z(n5953) );
  MUX2_X1 U24908 ( .A(n5953), .B(n5946), .S(n8207), .Z(n5954) );
  MUX2_X1 U24909 ( .A(\mem[174][5] ), .B(\mem[175][5] ), .S(n8444), .Z(n5955)
         );
  MUX2_X1 U24910 ( .A(\mem[172][5] ), .B(\mem[173][5] ), .S(n8444), .Z(n5956)
         );
  MUX2_X1 U24911 ( .A(n5956), .B(n5955), .S(n8309), .Z(n5957) );
  MUX2_X1 U24912 ( .A(\mem[170][5] ), .B(\mem[171][5] ), .S(n8444), .Z(n5958)
         );
  MUX2_X1 U24913 ( .A(\mem[168][5] ), .B(\mem[169][5] ), .S(n8444), .Z(n5959)
         );
  MUX2_X1 U24914 ( .A(n5959), .B(n5958), .S(n8309), .Z(n5960) );
  MUX2_X1 U24915 ( .A(n5960), .B(n5957), .S(n8250), .Z(n5961) );
  MUX2_X1 U24916 ( .A(\mem[166][5] ), .B(\mem[167][5] ), .S(n8444), .Z(n5962)
         );
  MUX2_X1 U24917 ( .A(\mem[164][5] ), .B(\mem[165][5] ), .S(n8444), .Z(n5963)
         );
  MUX2_X1 U24918 ( .A(n5963), .B(n5962), .S(n8309), .Z(n5964) );
  MUX2_X1 U24919 ( .A(\mem[162][5] ), .B(\mem[163][5] ), .S(n8444), .Z(n5965)
         );
  MUX2_X1 U24920 ( .A(\mem[160][5] ), .B(\mem[161][5] ), .S(n8444), .Z(n5966)
         );
  MUX2_X1 U24921 ( .A(n5966), .B(n5965), .S(n8309), .Z(n5967) );
  MUX2_X1 U24922 ( .A(n5967), .B(n5964), .S(n8251), .Z(n5968) );
  MUX2_X1 U24923 ( .A(n5968), .B(n5961), .S(n8207), .Z(n5969) );
  MUX2_X1 U24924 ( .A(n5969), .B(n5954), .S(n8190), .Z(n5970) );
  MUX2_X1 U24925 ( .A(\mem[158][5] ), .B(\mem[159][5] ), .S(n8445), .Z(n5971)
         );
  MUX2_X1 U24926 ( .A(\mem[156][5] ), .B(\mem[157][5] ), .S(n8445), .Z(n5972)
         );
  MUX2_X1 U24927 ( .A(n5972), .B(n5971), .S(n8310), .Z(n5973) );
  MUX2_X1 U24928 ( .A(\mem[154][5] ), .B(\mem[155][5] ), .S(n8445), .Z(n5974)
         );
  MUX2_X1 U24929 ( .A(\mem[152][5] ), .B(\mem[153][5] ), .S(n8445), .Z(n5975)
         );
  MUX2_X1 U24930 ( .A(n5975), .B(n5974), .S(n8310), .Z(n5976) );
  MUX2_X1 U24931 ( .A(n5976), .B(n5973), .S(n8224), .Z(n5977) );
  MUX2_X1 U24932 ( .A(\mem[150][5] ), .B(\mem[151][5] ), .S(n8445), .Z(n5978)
         );
  MUX2_X1 U24933 ( .A(\mem[148][5] ), .B(\mem[149][5] ), .S(n8445), .Z(n5979)
         );
  MUX2_X1 U24934 ( .A(n5979), .B(n5978), .S(n8310), .Z(n5980) );
  MUX2_X1 U24935 ( .A(\mem[146][5] ), .B(\mem[147][5] ), .S(n8445), .Z(n5981)
         );
  MUX2_X1 U24936 ( .A(\mem[144][5] ), .B(\mem[145][5] ), .S(n8445), .Z(n5982)
         );
  MUX2_X1 U24937 ( .A(n5982), .B(n5981), .S(n8310), .Z(n5983) );
  MUX2_X1 U24938 ( .A(n5983), .B(n5980), .S(n8241), .Z(n5984) );
  MUX2_X1 U24939 ( .A(n5984), .B(n5977), .S(n8207), .Z(n5985) );
  MUX2_X1 U24940 ( .A(\mem[142][5] ), .B(\mem[143][5] ), .S(n8445), .Z(n5986)
         );
  MUX2_X1 U24941 ( .A(\mem[140][5] ), .B(\mem[141][5] ), .S(n8445), .Z(n5987)
         );
  MUX2_X1 U24942 ( .A(n5987), .B(n5986), .S(n8310), .Z(n5988) );
  MUX2_X1 U24943 ( .A(\mem[138][5] ), .B(\mem[139][5] ), .S(n8445), .Z(n5989)
         );
  MUX2_X1 U24944 ( .A(\mem[136][5] ), .B(\mem[137][5] ), .S(n8445), .Z(n5990)
         );
  MUX2_X1 U24945 ( .A(n5990), .B(n5989), .S(n8310), .Z(n5991) );
  MUX2_X1 U24946 ( .A(n5991), .B(n5988), .S(n8220), .Z(n5992) );
  MUX2_X1 U24947 ( .A(\mem[134][5] ), .B(\mem[135][5] ), .S(n8446), .Z(n5993)
         );
  MUX2_X1 U24948 ( .A(\mem[132][5] ), .B(\mem[133][5] ), .S(n8446), .Z(n5994)
         );
  MUX2_X1 U24949 ( .A(n5994), .B(n5993), .S(n8310), .Z(n5995) );
  MUX2_X1 U24950 ( .A(\mem[130][5] ), .B(\mem[131][5] ), .S(n8446), .Z(n5996)
         );
  MUX2_X1 U24951 ( .A(\mem[128][5] ), .B(\mem[129][5] ), .S(n8446), .Z(n5997)
         );
  MUX2_X1 U24952 ( .A(n5997), .B(n5996), .S(n8310), .Z(n5998) );
  MUX2_X1 U24953 ( .A(n5998), .B(n5995), .S(n8239), .Z(n5999) );
  MUX2_X1 U24954 ( .A(n5999), .B(n5992), .S(n8207), .Z(n6000) );
  MUX2_X1 U24955 ( .A(n6000), .B(n5985), .S(n8190), .Z(n6001) );
  MUX2_X1 U24956 ( .A(n6001), .B(n5970), .S(n8184), .Z(n6002) );
  MUX2_X1 U24957 ( .A(n6002), .B(n5939), .S(N24), .Z(n6003) );
  MUX2_X1 U24958 ( .A(\mem[126][5] ), .B(\mem[127][5] ), .S(n8446), .Z(n6004)
         );
  MUX2_X1 U24959 ( .A(\mem[124][5] ), .B(\mem[125][5] ), .S(n8446), .Z(n6005)
         );
  MUX2_X1 U24960 ( .A(n6005), .B(n6004), .S(n8310), .Z(n6006) );
  MUX2_X1 U24961 ( .A(\mem[122][5] ), .B(\mem[123][5] ), .S(n8446), .Z(n6007)
         );
  MUX2_X1 U24962 ( .A(\mem[120][5] ), .B(\mem[121][5] ), .S(n8446), .Z(n6008)
         );
  MUX2_X1 U24963 ( .A(n6008), .B(n6007), .S(n8310), .Z(n6009) );
  MUX2_X1 U24964 ( .A(n6009), .B(n6006), .S(n8241), .Z(n6010) );
  MUX2_X1 U24965 ( .A(\mem[118][5] ), .B(\mem[119][5] ), .S(n8446), .Z(n6011)
         );
  MUX2_X1 U24966 ( .A(\mem[116][5] ), .B(\mem[117][5] ), .S(n8446), .Z(n6012)
         );
  MUX2_X1 U24967 ( .A(n6012), .B(n6011), .S(n8310), .Z(n6013) );
  MUX2_X1 U24968 ( .A(\mem[114][5] ), .B(\mem[115][5] ), .S(n8446), .Z(n6014)
         );
  MUX2_X1 U24969 ( .A(\mem[112][5] ), .B(\mem[113][5] ), .S(n8446), .Z(n6015)
         );
  MUX2_X1 U24970 ( .A(n6015), .B(n6014), .S(n8310), .Z(n6016) );
  MUX2_X1 U24971 ( .A(n6016), .B(n6013), .S(n8247), .Z(n6017) );
  MUX2_X1 U24972 ( .A(n6017), .B(n6010), .S(n8207), .Z(n6018) );
  MUX2_X1 U24973 ( .A(\mem[110][5] ), .B(\mem[111][5] ), .S(n8447), .Z(n6019)
         );
  MUX2_X1 U24974 ( .A(\mem[108][5] ), .B(\mem[109][5] ), .S(n8447), .Z(n6020)
         );
  MUX2_X1 U24975 ( .A(n6020), .B(n6019), .S(n8311), .Z(n6021) );
  MUX2_X1 U24976 ( .A(\mem[106][5] ), .B(\mem[107][5] ), .S(n8447), .Z(n6022)
         );
  MUX2_X1 U24977 ( .A(\mem[104][5] ), .B(\mem[105][5] ), .S(n8447), .Z(n6023)
         );
  MUX2_X1 U24978 ( .A(n6023), .B(n6022), .S(n8311), .Z(n6024) );
  MUX2_X1 U24979 ( .A(n6024), .B(n6021), .S(N20), .Z(n6025) );
  MUX2_X1 U24980 ( .A(\mem[102][5] ), .B(\mem[103][5] ), .S(n8447), .Z(n6026)
         );
  MUX2_X1 U24981 ( .A(\mem[100][5] ), .B(\mem[101][5] ), .S(n8447), .Z(n6027)
         );
  MUX2_X1 U24982 ( .A(n6027), .B(n6026), .S(n8311), .Z(n6028) );
  MUX2_X1 U24983 ( .A(\mem[98][5] ), .B(\mem[99][5] ), .S(n8447), .Z(n6029) );
  MUX2_X1 U24984 ( .A(\mem[96][5] ), .B(\mem[97][5] ), .S(n8447), .Z(n6030) );
  MUX2_X1 U24985 ( .A(n6030), .B(n6029), .S(n8311), .Z(n6031) );
  MUX2_X1 U24986 ( .A(n6031), .B(n6028), .S(n8263), .Z(n6032) );
  MUX2_X1 U24987 ( .A(n6032), .B(n6025), .S(n8207), .Z(n6033) );
  MUX2_X1 U24988 ( .A(n6033), .B(n6018), .S(n8190), .Z(n6034) );
  MUX2_X1 U24989 ( .A(\mem[94][5] ), .B(\mem[95][5] ), .S(n8447), .Z(n6035) );
  MUX2_X1 U24990 ( .A(\mem[92][5] ), .B(\mem[93][5] ), .S(n8447), .Z(n6036) );
  MUX2_X1 U24991 ( .A(n6036), .B(n6035), .S(n8311), .Z(n6037) );
  MUX2_X1 U24992 ( .A(\mem[90][5] ), .B(\mem[91][5] ), .S(n8447), .Z(n6038) );
  MUX2_X1 U24993 ( .A(\mem[88][5] ), .B(\mem[89][5] ), .S(n8447), .Z(n6039) );
  MUX2_X1 U24994 ( .A(n6039), .B(n6038), .S(n8311), .Z(n6040) );
  MUX2_X1 U24995 ( .A(n6040), .B(n6037), .S(n8242), .Z(n6041) );
  MUX2_X1 U24996 ( .A(\mem[86][5] ), .B(\mem[87][5] ), .S(n8448), .Z(n6042) );
  MUX2_X1 U24997 ( .A(\mem[84][5] ), .B(\mem[85][5] ), .S(n8448), .Z(n6043) );
  MUX2_X1 U24998 ( .A(n6043), .B(n6042), .S(n8311), .Z(n6044) );
  MUX2_X1 U24999 ( .A(\mem[82][5] ), .B(\mem[83][5] ), .S(n8448), .Z(n6045) );
  MUX2_X1 U25000 ( .A(\mem[80][5] ), .B(\mem[81][5] ), .S(n8448), .Z(n6046) );
  MUX2_X1 U25001 ( .A(n6046), .B(n6045), .S(n8311), .Z(n6047) );
  MUX2_X1 U25002 ( .A(n6047), .B(n6044), .S(n8264), .Z(n6048) );
  MUX2_X1 U25003 ( .A(n6048), .B(n6041), .S(n8207), .Z(n6049) );
  MUX2_X1 U25004 ( .A(\mem[78][5] ), .B(\mem[79][5] ), .S(n8448), .Z(n6050) );
  MUX2_X1 U25005 ( .A(\mem[76][5] ), .B(\mem[77][5] ), .S(n8448), .Z(n6051) );
  MUX2_X1 U25006 ( .A(n6051), .B(n6050), .S(n8311), .Z(n6052) );
  MUX2_X1 U25007 ( .A(\mem[74][5] ), .B(\mem[75][5] ), .S(n8448), .Z(n6053) );
  MUX2_X1 U25008 ( .A(\mem[72][5] ), .B(\mem[73][5] ), .S(n8448), .Z(n6054) );
  MUX2_X1 U25009 ( .A(n6054), .B(n6053), .S(n8311), .Z(n6055) );
  MUX2_X1 U25010 ( .A(n6055), .B(n6052), .S(n8250), .Z(n6056) );
  MUX2_X1 U25011 ( .A(\mem[70][5] ), .B(\mem[71][5] ), .S(n8448), .Z(n6057) );
  MUX2_X1 U25012 ( .A(\mem[68][5] ), .B(\mem[69][5] ), .S(n8448), .Z(n6058) );
  MUX2_X1 U25013 ( .A(n6058), .B(n6057), .S(n8311), .Z(n6059) );
  MUX2_X1 U25014 ( .A(\mem[66][5] ), .B(\mem[67][5] ), .S(n8448), .Z(n6060) );
  MUX2_X1 U25015 ( .A(\mem[64][5] ), .B(\mem[65][5] ), .S(n8448), .Z(n6061) );
  MUX2_X1 U25016 ( .A(n6061), .B(n6060), .S(n8311), .Z(n6062) );
  MUX2_X1 U25017 ( .A(n6062), .B(n6059), .S(n8262), .Z(n6063) );
  MUX2_X1 U25018 ( .A(n6063), .B(n6056), .S(n8207), .Z(n6064) );
  MUX2_X1 U25019 ( .A(n6064), .B(n6049), .S(n8190), .Z(n6065) );
  MUX2_X1 U25020 ( .A(n6065), .B(n6034), .S(N23), .Z(n6066) );
  MUX2_X1 U25021 ( .A(\mem[62][5] ), .B(\mem[63][5] ), .S(n8449), .Z(n6067) );
  MUX2_X1 U25022 ( .A(\mem[60][5] ), .B(\mem[61][5] ), .S(n8449), .Z(n6068) );
  MUX2_X1 U25023 ( .A(n6068), .B(n6067), .S(n8312), .Z(n6069) );
  MUX2_X1 U25024 ( .A(\mem[58][5] ), .B(\mem[59][5] ), .S(n8449), .Z(n6070) );
  MUX2_X1 U25025 ( .A(\mem[56][5] ), .B(\mem[57][5] ), .S(n8449), .Z(n6071) );
  MUX2_X1 U25026 ( .A(n6071), .B(n6070), .S(n8312), .Z(n6072) );
  MUX2_X1 U25027 ( .A(n6072), .B(n6069), .S(n8232), .Z(n6073) );
  MUX2_X1 U25028 ( .A(\mem[54][5] ), .B(\mem[55][5] ), .S(n8449), .Z(n6074) );
  MUX2_X1 U25029 ( .A(\mem[52][5] ), .B(\mem[53][5] ), .S(n8449), .Z(n6075) );
  MUX2_X1 U25030 ( .A(n6075), .B(n6074), .S(n8312), .Z(n6076) );
  MUX2_X1 U25031 ( .A(\mem[50][5] ), .B(\mem[51][5] ), .S(n8449), .Z(n6077) );
  MUX2_X1 U25032 ( .A(\mem[48][5] ), .B(\mem[49][5] ), .S(n8449), .Z(n6078) );
  MUX2_X1 U25033 ( .A(n6078), .B(n6077), .S(n8312), .Z(n6079) );
  MUX2_X1 U25034 ( .A(n6079), .B(n6076), .S(n8233), .Z(n6080) );
  MUX2_X1 U25035 ( .A(n6080), .B(n6073), .S(n8208), .Z(n6081) );
  MUX2_X1 U25036 ( .A(\mem[46][5] ), .B(\mem[47][5] ), .S(n8449), .Z(n6082) );
  MUX2_X1 U25037 ( .A(\mem[44][5] ), .B(\mem[45][5] ), .S(n8449), .Z(n6083) );
  MUX2_X1 U25038 ( .A(n6083), .B(n6082), .S(n8312), .Z(n6084) );
  MUX2_X1 U25039 ( .A(\mem[42][5] ), .B(\mem[43][5] ), .S(n8449), .Z(n6085) );
  MUX2_X1 U25040 ( .A(\mem[40][5] ), .B(\mem[41][5] ), .S(n8449), .Z(n6086) );
  MUX2_X1 U25041 ( .A(n6086), .B(n6085), .S(n8312), .Z(n6087) );
  MUX2_X1 U25042 ( .A(n6087), .B(n6084), .S(n8234), .Z(n6088) );
  MUX2_X1 U25043 ( .A(\mem[38][5] ), .B(\mem[39][5] ), .S(n8450), .Z(n6089) );
  MUX2_X1 U25044 ( .A(\mem[36][5] ), .B(\mem[37][5] ), .S(n8450), .Z(n6090) );
  MUX2_X1 U25045 ( .A(n6090), .B(n6089), .S(n8312), .Z(n6091) );
  MUX2_X1 U25046 ( .A(\mem[34][5] ), .B(\mem[35][5] ), .S(n8450), .Z(n6092) );
  MUX2_X1 U25047 ( .A(\mem[32][5] ), .B(\mem[33][5] ), .S(n8450), .Z(n6093) );
  MUX2_X1 U25048 ( .A(n6093), .B(n6092), .S(n8312), .Z(n6094) );
  MUX2_X1 U25049 ( .A(n6094), .B(n6091), .S(n8241), .Z(n6095) );
  MUX2_X1 U25050 ( .A(n6095), .B(n6088), .S(n8208), .Z(n6096) );
  MUX2_X1 U25051 ( .A(n6096), .B(n6081), .S(n8190), .Z(n6097) );
  MUX2_X1 U25052 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n8450), .Z(n6098) );
  MUX2_X1 U25053 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n8450), .Z(n6099) );
  MUX2_X1 U25054 ( .A(n6099), .B(n6098), .S(n8312), .Z(n6100) );
  MUX2_X1 U25055 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n8450), .Z(n6101) );
  MUX2_X1 U25056 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n8450), .Z(n6102) );
  MUX2_X1 U25057 ( .A(n6102), .B(n6101), .S(n8312), .Z(n6103) );
  MUX2_X1 U25058 ( .A(n6103), .B(n6100), .S(n8242), .Z(n6104) );
  MUX2_X1 U25059 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n8450), .Z(n6105) );
  MUX2_X1 U25060 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n8450), .Z(n6106) );
  MUX2_X1 U25061 ( .A(n6106), .B(n6105), .S(n8312), .Z(n6107) );
  MUX2_X1 U25062 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n8450), .Z(n6108) );
  MUX2_X1 U25063 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n8450), .Z(n6109) );
  MUX2_X1 U25064 ( .A(n6109), .B(n6108), .S(n8312), .Z(n6110) );
  MUX2_X1 U25065 ( .A(n6110), .B(n6107), .S(n8243), .Z(n6111) );
  MUX2_X1 U25066 ( .A(n6111), .B(n6104), .S(n8208), .Z(n6112) );
  MUX2_X1 U25067 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n8451), .Z(n6113) );
  MUX2_X1 U25068 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n8451), .Z(n6114) );
  MUX2_X1 U25069 ( .A(n6114), .B(n6113), .S(n8313), .Z(n6115) );
  MUX2_X1 U25070 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n8451), .Z(n6116) );
  MUX2_X1 U25071 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n8451), .Z(n6117) );
  MUX2_X1 U25072 ( .A(n6117), .B(n6116), .S(n8313), .Z(n6118) );
  MUX2_X1 U25073 ( .A(n6118), .B(n6115), .S(n8238), .Z(n6119) );
  MUX2_X1 U25074 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n8451), .Z(n6120) );
  MUX2_X1 U25075 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n8451), .Z(n6121) );
  MUX2_X1 U25076 ( .A(n6121), .B(n6120), .S(n8313), .Z(n6122) );
  MUX2_X1 U25077 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n8451), .Z(n6123) );
  MUX2_X1 U25078 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n8451), .Z(n6124) );
  MUX2_X1 U25079 ( .A(n6124), .B(n6123), .S(n8313), .Z(n6125) );
  MUX2_X1 U25080 ( .A(n6125), .B(n6122), .S(n8239), .Z(n6126) );
  MUX2_X1 U25081 ( .A(n6126), .B(n6119), .S(n8208), .Z(n6127) );
  MUX2_X1 U25082 ( .A(n6127), .B(n6112), .S(n8190), .Z(n6128) );
  MUX2_X1 U25083 ( .A(n6128), .B(n6097), .S(n8183), .Z(n6129) );
  MUX2_X1 U25084 ( .A(n6129), .B(n6066), .S(n8178), .Z(n6130) );
  MUX2_X1 U25085 ( .A(n6130), .B(n6003), .S(n8177), .Z(n6131) );
  MUX2_X1 U25086 ( .A(n6131), .B(n5876), .S(N26), .Z(n6132) );
  MUX2_X1 U25087 ( .A(n6132), .B(n5621), .S(N27), .Z(N30) );
  MUX2_X1 U25088 ( .A(\mem[1022][6] ), .B(\mem[1023][6] ), .S(n8451), .Z(n6133) );
  MUX2_X1 U25089 ( .A(\mem[1020][6] ), .B(\mem[1021][6] ), .S(n8451), .Z(n6134) );
  MUX2_X1 U25090 ( .A(n6134), .B(n6133), .S(n8313), .Z(n6135) );
  MUX2_X1 U25091 ( .A(\mem[1018][6] ), .B(\mem[1019][6] ), .S(n8451), .Z(n6136) );
  MUX2_X1 U25092 ( .A(\mem[1016][6] ), .B(\mem[1017][6] ), .S(n8451), .Z(n6137) );
  MUX2_X1 U25093 ( .A(n6137), .B(n6136), .S(n8313), .Z(n6138) );
  MUX2_X1 U25094 ( .A(n6138), .B(n6135), .S(n8240), .Z(n6139) );
  MUX2_X1 U25095 ( .A(\mem[1014][6] ), .B(\mem[1015][6] ), .S(n8452), .Z(n6140) );
  MUX2_X1 U25096 ( .A(\mem[1012][6] ), .B(\mem[1013][6] ), .S(n8452), .Z(n6141) );
  MUX2_X1 U25097 ( .A(n6141), .B(n6140), .S(n8313), .Z(n6142) );
  MUX2_X1 U25098 ( .A(\mem[1010][6] ), .B(\mem[1011][6] ), .S(n8452), .Z(n6143) );
  MUX2_X1 U25099 ( .A(\mem[1008][6] ), .B(\mem[1009][6] ), .S(n8452), .Z(n6144) );
  MUX2_X1 U25100 ( .A(n6144), .B(n6143), .S(n8313), .Z(n6145) );
  MUX2_X1 U25101 ( .A(n6145), .B(n6142), .S(n8230), .Z(n6146) );
  MUX2_X1 U25102 ( .A(n6146), .B(n6139), .S(n8208), .Z(n6147) );
  MUX2_X1 U25103 ( .A(\mem[1006][6] ), .B(\mem[1007][6] ), .S(n8452), .Z(n6148) );
  MUX2_X1 U25104 ( .A(\mem[1004][6] ), .B(\mem[1005][6] ), .S(n8452), .Z(n6149) );
  MUX2_X1 U25105 ( .A(n6149), .B(n6148), .S(n8313), .Z(n6150) );
  MUX2_X1 U25106 ( .A(\mem[1002][6] ), .B(\mem[1003][6] ), .S(n8452), .Z(n6151) );
  MUX2_X1 U25107 ( .A(\mem[1000][6] ), .B(\mem[1001][6] ), .S(n8452), .Z(n6152) );
  MUX2_X1 U25108 ( .A(n6152), .B(n6151), .S(n8313), .Z(n6153) );
  MUX2_X1 U25109 ( .A(n6153), .B(n6150), .S(n8231), .Z(n6154) );
  MUX2_X1 U25110 ( .A(\mem[998][6] ), .B(\mem[999][6] ), .S(n8452), .Z(n6155)
         );
  MUX2_X1 U25111 ( .A(\mem[996][6] ), .B(\mem[997][6] ), .S(n8452), .Z(n6156)
         );
  MUX2_X1 U25112 ( .A(n6156), .B(n6155), .S(n8313), .Z(n6157) );
  MUX2_X1 U25113 ( .A(\mem[994][6] ), .B(\mem[995][6] ), .S(n8452), .Z(n6158)
         );
  MUX2_X1 U25114 ( .A(\mem[992][6] ), .B(\mem[993][6] ), .S(n8452), .Z(n6159)
         );
  MUX2_X1 U25115 ( .A(n6159), .B(n6158), .S(n8313), .Z(n6160) );
  MUX2_X1 U25116 ( .A(n6160), .B(n6157), .S(n8227), .Z(n6161) );
  MUX2_X1 U25117 ( .A(n6161), .B(n6154), .S(n8208), .Z(n6162) );
  MUX2_X1 U25118 ( .A(n6162), .B(n6147), .S(n8190), .Z(n6163) );
  MUX2_X1 U25119 ( .A(\mem[990][6] ), .B(\mem[991][6] ), .S(n8453), .Z(n6164)
         );
  MUX2_X1 U25120 ( .A(\mem[988][6] ), .B(\mem[989][6] ), .S(n8453), .Z(n6165)
         );
  MUX2_X1 U25121 ( .A(n6165), .B(n6164), .S(n8314), .Z(n6166) );
  MUX2_X1 U25122 ( .A(\mem[986][6] ), .B(\mem[987][6] ), .S(n8453), .Z(n6167)
         );
  MUX2_X1 U25123 ( .A(\mem[984][6] ), .B(\mem[985][6] ), .S(n8453), .Z(n6168)
         );
  MUX2_X1 U25124 ( .A(n6168), .B(n6167), .S(n8314), .Z(n6169) );
  MUX2_X1 U25125 ( .A(n6169), .B(n6166), .S(n8244), .Z(n6170) );
  MUX2_X1 U25126 ( .A(\mem[982][6] ), .B(\mem[983][6] ), .S(n8453), .Z(n6171)
         );
  MUX2_X1 U25127 ( .A(\mem[980][6] ), .B(\mem[981][6] ), .S(n8453), .Z(n6172)
         );
  MUX2_X1 U25128 ( .A(n6172), .B(n6171), .S(n8314), .Z(n6173) );
  MUX2_X1 U25129 ( .A(\mem[978][6] ), .B(\mem[979][6] ), .S(n8453), .Z(n6174)
         );
  MUX2_X1 U25130 ( .A(\mem[976][6] ), .B(\mem[977][6] ), .S(n8453), .Z(n6175)
         );
  MUX2_X1 U25131 ( .A(n6175), .B(n6174), .S(n8314), .Z(n6176) );
  MUX2_X1 U25132 ( .A(n6176), .B(n6173), .S(n8224), .Z(n6177) );
  MUX2_X1 U25133 ( .A(n6177), .B(n6170), .S(n8208), .Z(n6178) );
  MUX2_X1 U25134 ( .A(\mem[974][6] ), .B(\mem[975][6] ), .S(n8453), .Z(n6179)
         );
  MUX2_X1 U25135 ( .A(\mem[972][6] ), .B(\mem[973][6] ), .S(n8453), .Z(n6180)
         );
  MUX2_X1 U25136 ( .A(n6180), .B(n6179), .S(n8314), .Z(n6181) );
  MUX2_X1 U25137 ( .A(\mem[970][6] ), .B(\mem[971][6] ), .S(n8453), .Z(n6182)
         );
  MUX2_X1 U25138 ( .A(\mem[968][6] ), .B(\mem[969][6] ), .S(n8453), .Z(n6183)
         );
  MUX2_X1 U25139 ( .A(n6183), .B(n6182), .S(n8314), .Z(n6184) );
  MUX2_X1 U25140 ( .A(n6184), .B(n6181), .S(n8223), .Z(n6185) );
  MUX2_X1 U25141 ( .A(\mem[966][6] ), .B(\mem[967][6] ), .S(n8454), .Z(n6186)
         );
  MUX2_X1 U25142 ( .A(\mem[964][6] ), .B(\mem[965][6] ), .S(n8454), .Z(n6187)
         );
  MUX2_X1 U25143 ( .A(n6187), .B(n6186), .S(n8314), .Z(n6188) );
  MUX2_X1 U25144 ( .A(\mem[962][6] ), .B(\mem[963][6] ), .S(n8454), .Z(n6189)
         );
  MUX2_X1 U25145 ( .A(\mem[960][6] ), .B(\mem[961][6] ), .S(n8454), .Z(n6190)
         );
  MUX2_X1 U25146 ( .A(n6190), .B(n6189), .S(n8314), .Z(n6191) );
  MUX2_X1 U25147 ( .A(n6191), .B(n6188), .S(n8222), .Z(n6192) );
  MUX2_X1 U25148 ( .A(n6192), .B(n6185), .S(n8208), .Z(n6193) );
  MUX2_X1 U25149 ( .A(n6193), .B(n6178), .S(n8190), .Z(n6194) );
  MUX2_X1 U25150 ( .A(n6194), .B(n6163), .S(n8185), .Z(n6195) );
  MUX2_X1 U25151 ( .A(\mem[958][6] ), .B(\mem[959][6] ), .S(n8454), .Z(n6196)
         );
  MUX2_X1 U25152 ( .A(\mem[956][6] ), .B(\mem[957][6] ), .S(n8454), .Z(n6197)
         );
  MUX2_X1 U25153 ( .A(n6197), .B(n6196), .S(n8314), .Z(n6198) );
  MUX2_X1 U25154 ( .A(\mem[954][6] ), .B(\mem[955][6] ), .S(n8454), .Z(n6199)
         );
  MUX2_X1 U25155 ( .A(\mem[952][6] ), .B(\mem[953][6] ), .S(n8454), .Z(n6200)
         );
  MUX2_X1 U25156 ( .A(n6200), .B(n6199), .S(n8314), .Z(n6201) );
  MUX2_X1 U25157 ( .A(n6201), .B(n6198), .S(n8221), .Z(n6202) );
  MUX2_X1 U25158 ( .A(\mem[950][6] ), .B(\mem[951][6] ), .S(n8454), .Z(n6203)
         );
  MUX2_X1 U25159 ( .A(\mem[948][6] ), .B(\mem[949][6] ), .S(n8454), .Z(n6204)
         );
  MUX2_X1 U25160 ( .A(n6204), .B(n6203), .S(n8314), .Z(n6205) );
  MUX2_X1 U25161 ( .A(\mem[946][6] ), .B(\mem[947][6] ), .S(n8454), .Z(n6206)
         );
  MUX2_X1 U25162 ( .A(\mem[944][6] ), .B(\mem[945][6] ), .S(n8454), .Z(n6207)
         );
  MUX2_X1 U25163 ( .A(n6207), .B(n6206), .S(n8314), .Z(n6208) );
  MUX2_X1 U25164 ( .A(n6208), .B(n6205), .S(n8220), .Z(n6209) );
  MUX2_X1 U25165 ( .A(n6209), .B(n6202), .S(n8208), .Z(n6210) );
  MUX2_X1 U25166 ( .A(\mem[942][6] ), .B(\mem[943][6] ), .S(n8455), .Z(n6211)
         );
  MUX2_X1 U25167 ( .A(\mem[940][6] ), .B(\mem[941][6] ), .S(n8455), .Z(n6212)
         );
  MUX2_X1 U25168 ( .A(n6212), .B(n6211), .S(n8315), .Z(n6213) );
  MUX2_X1 U25169 ( .A(\mem[938][6] ), .B(\mem[939][6] ), .S(n8455), .Z(n6214)
         );
  MUX2_X1 U25170 ( .A(\mem[936][6] ), .B(\mem[937][6] ), .S(n8455), .Z(n6215)
         );
  MUX2_X1 U25171 ( .A(n6215), .B(n6214), .S(n8315), .Z(n6216) );
  MUX2_X1 U25172 ( .A(n6216), .B(n6213), .S(n8251), .Z(n6217) );
  MUX2_X1 U25173 ( .A(\mem[934][6] ), .B(\mem[935][6] ), .S(n8455), .Z(n6218)
         );
  MUX2_X1 U25174 ( .A(\mem[932][6] ), .B(\mem[933][6] ), .S(n8455), .Z(n6219)
         );
  MUX2_X1 U25175 ( .A(n6219), .B(n6218), .S(n8315), .Z(n6220) );
  MUX2_X1 U25176 ( .A(\mem[930][6] ), .B(\mem[931][6] ), .S(n8455), .Z(n6221)
         );
  MUX2_X1 U25177 ( .A(\mem[928][6] ), .B(\mem[929][6] ), .S(n8455), .Z(n6222)
         );
  MUX2_X1 U25178 ( .A(n6222), .B(n6221), .S(n8315), .Z(n6223) );
  MUX2_X1 U25179 ( .A(n6223), .B(n6220), .S(n8231), .Z(n6224) );
  MUX2_X1 U25180 ( .A(n6224), .B(n6217), .S(n8208), .Z(n6225) );
  MUX2_X1 U25181 ( .A(n6225), .B(n6210), .S(n8190), .Z(n6226) );
  MUX2_X1 U25182 ( .A(\mem[926][6] ), .B(\mem[927][6] ), .S(n8455), .Z(n6227)
         );
  MUX2_X1 U25183 ( .A(\mem[924][6] ), .B(\mem[925][6] ), .S(n8455), .Z(n6228)
         );
  MUX2_X1 U25184 ( .A(n6228), .B(n6227), .S(n8315), .Z(n6229) );
  MUX2_X1 U25185 ( .A(\mem[922][6] ), .B(\mem[923][6] ), .S(n8455), .Z(n6230)
         );
  MUX2_X1 U25186 ( .A(\mem[920][6] ), .B(\mem[921][6] ), .S(n8455), .Z(n6231)
         );
  MUX2_X1 U25187 ( .A(n6231), .B(n6230), .S(n8315), .Z(n6232) );
  MUX2_X1 U25188 ( .A(n6232), .B(n6229), .S(n8235), .Z(n6233) );
  MUX2_X1 U25189 ( .A(\mem[918][6] ), .B(\mem[919][6] ), .S(n8456), .Z(n6234)
         );
  MUX2_X1 U25190 ( .A(\mem[916][6] ), .B(\mem[917][6] ), .S(n8456), .Z(n6235)
         );
  MUX2_X1 U25191 ( .A(n6235), .B(n6234), .S(n8315), .Z(n6236) );
  MUX2_X1 U25192 ( .A(\mem[914][6] ), .B(\mem[915][6] ), .S(n8456), .Z(n6237)
         );
  MUX2_X1 U25193 ( .A(\mem[912][6] ), .B(\mem[913][6] ), .S(n8456), .Z(n6238)
         );
  MUX2_X1 U25194 ( .A(n6238), .B(n6237), .S(n8315), .Z(n6239) );
  MUX2_X1 U25195 ( .A(n6239), .B(n6236), .S(n8265), .Z(n6240) );
  MUX2_X1 U25196 ( .A(n6240), .B(n6233), .S(n8208), .Z(n6241) );
  MUX2_X1 U25197 ( .A(\mem[910][6] ), .B(\mem[911][6] ), .S(n8456), .Z(n6242)
         );
  MUX2_X1 U25198 ( .A(\mem[908][6] ), .B(\mem[909][6] ), .S(n8456), .Z(n6243)
         );
  MUX2_X1 U25199 ( .A(n6243), .B(n6242), .S(n8315), .Z(n6244) );
  MUX2_X1 U25200 ( .A(\mem[906][6] ), .B(\mem[907][6] ), .S(n8456), .Z(n6245)
         );
  MUX2_X1 U25201 ( .A(\mem[904][6] ), .B(\mem[905][6] ), .S(n8456), .Z(n6246)
         );
  MUX2_X1 U25202 ( .A(n6246), .B(n6245), .S(n8315), .Z(n6247) );
  MUX2_X1 U25203 ( .A(n6247), .B(n6244), .S(n8246), .Z(n6248) );
  MUX2_X1 U25204 ( .A(\mem[902][6] ), .B(\mem[903][6] ), .S(n8456), .Z(n6249)
         );
  MUX2_X1 U25205 ( .A(\mem[900][6] ), .B(\mem[901][6] ), .S(n8456), .Z(n6250)
         );
  MUX2_X1 U25206 ( .A(n6250), .B(n6249), .S(n8315), .Z(n6251) );
  MUX2_X1 U25207 ( .A(\mem[898][6] ), .B(\mem[899][6] ), .S(n8456), .Z(n6252)
         );
  MUX2_X1 U25208 ( .A(\mem[896][6] ), .B(\mem[897][6] ), .S(n8456), .Z(n6253)
         );
  MUX2_X1 U25209 ( .A(n6253), .B(n6252), .S(n8315), .Z(n6254) );
  MUX2_X1 U25210 ( .A(n6254), .B(n6251), .S(n8235), .Z(n6255) );
  MUX2_X1 U25211 ( .A(n6255), .B(n6248), .S(n8208), .Z(n6256) );
  MUX2_X1 U25212 ( .A(n6256), .B(n6241), .S(n8190), .Z(n6257) );
  MUX2_X1 U25213 ( .A(n6257), .B(n6226), .S(N23), .Z(n6258) );
  MUX2_X1 U25214 ( .A(n6258), .B(n6195), .S(N24), .Z(n6259) );
  MUX2_X1 U25215 ( .A(\mem[894][6] ), .B(\mem[895][6] ), .S(n8457), .Z(n6260)
         );
  MUX2_X1 U25216 ( .A(\mem[892][6] ), .B(\mem[893][6] ), .S(n8457), .Z(n6261)
         );
  MUX2_X1 U25217 ( .A(n6261), .B(n6260), .S(n8316), .Z(n6262) );
  MUX2_X1 U25218 ( .A(\mem[890][6] ), .B(\mem[891][6] ), .S(n8457), .Z(n6263)
         );
  MUX2_X1 U25219 ( .A(\mem[888][6] ), .B(\mem[889][6] ), .S(n8457), .Z(n6264)
         );
  MUX2_X1 U25220 ( .A(n6264), .B(n6263), .S(n8316), .Z(n6265) );
  MUX2_X1 U25221 ( .A(n6265), .B(n6262), .S(n8249), .Z(n6266) );
  MUX2_X1 U25222 ( .A(\mem[886][6] ), .B(\mem[887][6] ), .S(n8457), .Z(n6267)
         );
  MUX2_X1 U25223 ( .A(\mem[884][6] ), .B(\mem[885][6] ), .S(n8457), .Z(n6268)
         );
  MUX2_X1 U25224 ( .A(n6268), .B(n6267), .S(n8316), .Z(n6269) );
  MUX2_X1 U25225 ( .A(\mem[882][6] ), .B(\mem[883][6] ), .S(n8457), .Z(n6270)
         );
  MUX2_X1 U25226 ( .A(\mem[880][6] ), .B(\mem[881][6] ), .S(n8457), .Z(n6271)
         );
  MUX2_X1 U25227 ( .A(n6271), .B(n6270), .S(n8316), .Z(n6272) );
  MUX2_X1 U25228 ( .A(n6272), .B(n6269), .S(n8244), .Z(n6273) );
  MUX2_X1 U25229 ( .A(n6273), .B(n6266), .S(n8209), .Z(n6274) );
  MUX2_X1 U25230 ( .A(\mem[878][6] ), .B(\mem[879][6] ), .S(n8457), .Z(n6275)
         );
  MUX2_X1 U25231 ( .A(\mem[876][6] ), .B(\mem[877][6] ), .S(n8457), .Z(n6276)
         );
  MUX2_X1 U25232 ( .A(n6276), .B(n6275), .S(n8316), .Z(n6277) );
  MUX2_X1 U25233 ( .A(\mem[874][6] ), .B(\mem[875][6] ), .S(n8457), .Z(n6278)
         );
  MUX2_X1 U25234 ( .A(\mem[872][6] ), .B(\mem[873][6] ), .S(n8457), .Z(n6279)
         );
  MUX2_X1 U25235 ( .A(n6279), .B(n6278), .S(n8316), .Z(n6280) );
  MUX2_X1 U25236 ( .A(n6280), .B(n6277), .S(n8245), .Z(n6281) );
  MUX2_X1 U25237 ( .A(\mem[870][6] ), .B(\mem[871][6] ), .S(n8458), .Z(n6282)
         );
  MUX2_X1 U25238 ( .A(\mem[868][6] ), .B(\mem[869][6] ), .S(n8458), .Z(n6283)
         );
  MUX2_X1 U25239 ( .A(n6283), .B(n6282), .S(n8316), .Z(n6284) );
  MUX2_X1 U25240 ( .A(\mem[866][6] ), .B(\mem[867][6] ), .S(n8458), .Z(n6285)
         );
  MUX2_X1 U25241 ( .A(\mem[864][6] ), .B(\mem[865][6] ), .S(n8458), .Z(n6286)
         );
  MUX2_X1 U25242 ( .A(n6286), .B(n6285), .S(n8316), .Z(n6287) );
  MUX2_X1 U25243 ( .A(n6287), .B(n6284), .S(n8246), .Z(n6288) );
  MUX2_X1 U25244 ( .A(n6288), .B(n6281), .S(n8209), .Z(n6289) );
  MUX2_X1 U25245 ( .A(n6289), .B(n6274), .S(n8187), .Z(n6290) );
  MUX2_X1 U25246 ( .A(\mem[862][6] ), .B(\mem[863][6] ), .S(n8458), .Z(n6291)
         );
  MUX2_X1 U25247 ( .A(\mem[860][6] ), .B(\mem[861][6] ), .S(n8458), .Z(n6292)
         );
  MUX2_X1 U25248 ( .A(n6292), .B(n6291), .S(n8316), .Z(n6293) );
  MUX2_X1 U25249 ( .A(\mem[858][6] ), .B(\mem[859][6] ), .S(n8458), .Z(n6294)
         );
  MUX2_X1 U25250 ( .A(\mem[856][6] ), .B(\mem[857][6] ), .S(n8458), .Z(n6295)
         );
  MUX2_X1 U25251 ( .A(n6295), .B(n6294), .S(n8316), .Z(n6296) );
  MUX2_X1 U25252 ( .A(n6296), .B(n6293), .S(n8253), .Z(n6297) );
  MUX2_X1 U25253 ( .A(\mem[854][6] ), .B(\mem[855][6] ), .S(n8458), .Z(n6298)
         );
  MUX2_X1 U25254 ( .A(\mem[852][6] ), .B(\mem[853][6] ), .S(n8458), .Z(n6299)
         );
  MUX2_X1 U25255 ( .A(n6299), .B(n6298), .S(n8316), .Z(n6300) );
  MUX2_X1 U25256 ( .A(\mem[850][6] ), .B(\mem[851][6] ), .S(n8458), .Z(n6301)
         );
  MUX2_X1 U25257 ( .A(\mem[848][6] ), .B(\mem[849][6] ), .S(n8458), .Z(n6302)
         );
  MUX2_X1 U25258 ( .A(n6302), .B(n6301), .S(n8316), .Z(n6303) );
  MUX2_X1 U25259 ( .A(n6303), .B(n6300), .S(n8254), .Z(n6304) );
  MUX2_X1 U25260 ( .A(n6304), .B(n6297), .S(n8209), .Z(n6305) );
  MUX2_X1 U25261 ( .A(\mem[846][6] ), .B(\mem[847][6] ), .S(n8459), .Z(n6306)
         );
  MUX2_X1 U25262 ( .A(\mem[844][6] ), .B(\mem[845][6] ), .S(n8459), .Z(n6307)
         );
  MUX2_X1 U25263 ( .A(n6307), .B(n6306), .S(n8317), .Z(n6308) );
  MUX2_X1 U25264 ( .A(\mem[842][6] ), .B(\mem[843][6] ), .S(n8459), .Z(n6309)
         );
  MUX2_X1 U25265 ( .A(\mem[840][6] ), .B(\mem[841][6] ), .S(n8459), .Z(n6310)
         );
  MUX2_X1 U25266 ( .A(n6310), .B(n6309), .S(n8317), .Z(n6311) );
  MUX2_X1 U25267 ( .A(n6311), .B(n6308), .S(n8255), .Z(n6312) );
  MUX2_X1 U25268 ( .A(\mem[838][6] ), .B(\mem[839][6] ), .S(n8459), .Z(n6313)
         );
  MUX2_X1 U25269 ( .A(\mem[836][6] ), .B(\mem[837][6] ), .S(n8459), .Z(n6314)
         );
  MUX2_X1 U25270 ( .A(n6314), .B(n6313), .S(n8317), .Z(n6315) );
  MUX2_X1 U25271 ( .A(\mem[834][6] ), .B(\mem[835][6] ), .S(n8459), .Z(n6316)
         );
  MUX2_X1 U25272 ( .A(\mem[832][6] ), .B(\mem[833][6] ), .S(n8459), .Z(n6317)
         );
  MUX2_X1 U25273 ( .A(n6317), .B(n6316), .S(n8317), .Z(n6318) );
  MUX2_X1 U25274 ( .A(n6318), .B(n6315), .S(n8250), .Z(n6319) );
  MUX2_X1 U25275 ( .A(n6319), .B(n6312), .S(n8209), .Z(n6320) );
  MUX2_X1 U25276 ( .A(n6320), .B(n6305), .S(n8188), .Z(n6321) );
  MUX2_X1 U25277 ( .A(n6321), .B(n6290), .S(n8181), .Z(n6322) );
  MUX2_X1 U25278 ( .A(\mem[830][6] ), .B(\mem[831][6] ), .S(n8459), .Z(n6323)
         );
  MUX2_X1 U25279 ( .A(\mem[828][6] ), .B(\mem[829][6] ), .S(n8459), .Z(n6324)
         );
  MUX2_X1 U25280 ( .A(n6324), .B(n6323), .S(n8317), .Z(n6325) );
  MUX2_X1 U25281 ( .A(\mem[826][6] ), .B(\mem[827][6] ), .S(n8459), .Z(n6326)
         );
  MUX2_X1 U25282 ( .A(\mem[824][6] ), .B(\mem[825][6] ), .S(n8459), .Z(n6327)
         );
  MUX2_X1 U25283 ( .A(n6327), .B(n6326), .S(n8317), .Z(n6328) );
  MUX2_X1 U25284 ( .A(n6328), .B(n6325), .S(n8251), .Z(n6329) );
  MUX2_X1 U25285 ( .A(\mem[822][6] ), .B(\mem[823][6] ), .S(n8460), .Z(n6330)
         );
  MUX2_X1 U25286 ( .A(\mem[820][6] ), .B(\mem[821][6] ), .S(n8460), .Z(n6331)
         );
  MUX2_X1 U25287 ( .A(n6331), .B(n6330), .S(n8317), .Z(n6332) );
  MUX2_X1 U25288 ( .A(\mem[818][6] ), .B(\mem[819][6] ), .S(n8460), .Z(n6333)
         );
  MUX2_X1 U25289 ( .A(\mem[816][6] ), .B(\mem[817][6] ), .S(n8460), .Z(n6334)
         );
  MUX2_X1 U25290 ( .A(n6334), .B(n6333), .S(n8317), .Z(n6335) );
  MUX2_X1 U25291 ( .A(n6335), .B(n6332), .S(n8252), .Z(n6336) );
  MUX2_X1 U25292 ( .A(n6336), .B(n6329), .S(n8209), .Z(n6337) );
  MUX2_X1 U25293 ( .A(\mem[814][6] ), .B(\mem[815][6] ), .S(n8460), .Z(n6338)
         );
  MUX2_X1 U25294 ( .A(\mem[812][6] ), .B(\mem[813][6] ), .S(n8460), .Z(n6339)
         );
  MUX2_X1 U25295 ( .A(n6339), .B(n6338), .S(n8317), .Z(n6340) );
  MUX2_X1 U25296 ( .A(\mem[810][6] ), .B(\mem[811][6] ), .S(n8460), .Z(n6341)
         );
  MUX2_X1 U25297 ( .A(\mem[808][6] ), .B(\mem[809][6] ), .S(n8460), .Z(n6342)
         );
  MUX2_X1 U25298 ( .A(n6342), .B(n6341), .S(n8317), .Z(n6343) );
  MUX2_X1 U25299 ( .A(n6343), .B(n6340), .S(n8259), .Z(n6344) );
  MUX2_X1 U25300 ( .A(\mem[806][6] ), .B(\mem[807][6] ), .S(n8460), .Z(n6345)
         );
  MUX2_X1 U25301 ( .A(\mem[804][6] ), .B(\mem[805][6] ), .S(n8460), .Z(n6346)
         );
  MUX2_X1 U25302 ( .A(n6346), .B(n6345), .S(n8317), .Z(n6347) );
  MUX2_X1 U25303 ( .A(\mem[802][6] ), .B(\mem[803][6] ), .S(n8460), .Z(n6348)
         );
  MUX2_X1 U25304 ( .A(\mem[800][6] ), .B(\mem[801][6] ), .S(n8460), .Z(n6349)
         );
  MUX2_X1 U25305 ( .A(n6349), .B(n6348), .S(n8317), .Z(n6350) );
  MUX2_X1 U25306 ( .A(n6350), .B(n6347), .S(n8260), .Z(n6351) );
  MUX2_X1 U25307 ( .A(n6351), .B(n6344), .S(n8209), .Z(n6352) );
  MUX2_X1 U25308 ( .A(n6352), .B(n6337), .S(n8194), .Z(n6353) );
  MUX2_X1 U25309 ( .A(\mem[798][6] ), .B(\mem[799][6] ), .S(n8461), .Z(n6354)
         );
  MUX2_X1 U25310 ( .A(\mem[796][6] ), .B(\mem[797][6] ), .S(n8461), .Z(n6355)
         );
  MUX2_X1 U25311 ( .A(n6355), .B(n6354), .S(n8318), .Z(n6356) );
  MUX2_X1 U25312 ( .A(\mem[794][6] ), .B(\mem[795][6] ), .S(n8461), .Z(n6357)
         );
  MUX2_X1 U25313 ( .A(\mem[792][6] ), .B(\mem[793][6] ), .S(n8461), .Z(n6358)
         );
  MUX2_X1 U25314 ( .A(n6358), .B(n6357), .S(n8318), .Z(n6359) );
  MUX2_X1 U25315 ( .A(n6359), .B(n6356), .S(n8220), .Z(n6360) );
  MUX2_X1 U25316 ( .A(\mem[790][6] ), .B(\mem[791][6] ), .S(n8461), .Z(n6361)
         );
  MUX2_X1 U25317 ( .A(\mem[788][6] ), .B(\mem[789][6] ), .S(n8461), .Z(n6362)
         );
  MUX2_X1 U25318 ( .A(n6362), .B(n6361), .S(n8318), .Z(n6363) );
  MUX2_X1 U25319 ( .A(\mem[786][6] ), .B(\mem[787][6] ), .S(n8461), .Z(n6364)
         );
  MUX2_X1 U25320 ( .A(\mem[784][6] ), .B(\mem[785][6] ), .S(n8461), .Z(n6365)
         );
  MUX2_X1 U25321 ( .A(n6365), .B(n6364), .S(n8318), .Z(n6366) );
  MUX2_X1 U25322 ( .A(n6366), .B(n6363), .S(n8226), .Z(n6367) );
  MUX2_X1 U25323 ( .A(n6367), .B(n6360), .S(n8209), .Z(n6368) );
  MUX2_X1 U25324 ( .A(\mem[782][6] ), .B(\mem[783][6] ), .S(n8461), .Z(n6369)
         );
  MUX2_X1 U25325 ( .A(\mem[780][6] ), .B(\mem[781][6] ), .S(n8461), .Z(n6370)
         );
  MUX2_X1 U25326 ( .A(n6370), .B(n6369), .S(n8318), .Z(n6371) );
  MUX2_X1 U25327 ( .A(\mem[778][6] ), .B(\mem[779][6] ), .S(n8461), .Z(n6372)
         );
  MUX2_X1 U25328 ( .A(\mem[776][6] ), .B(\mem[777][6] ), .S(n8461), .Z(n6373)
         );
  MUX2_X1 U25329 ( .A(n6373), .B(n6372), .S(n8318), .Z(n6374) );
  MUX2_X1 U25330 ( .A(n6374), .B(n6371), .S(n8240), .Z(n6375) );
  MUX2_X1 U25331 ( .A(\mem[774][6] ), .B(\mem[775][6] ), .S(n8462), .Z(n6376)
         );
  MUX2_X1 U25332 ( .A(\mem[772][6] ), .B(\mem[773][6] ), .S(n8462), .Z(n6377)
         );
  MUX2_X1 U25333 ( .A(n6377), .B(n6376), .S(n8318), .Z(n6378) );
  MUX2_X1 U25334 ( .A(\mem[770][6] ), .B(\mem[771][6] ), .S(n8462), .Z(n6379)
         );
  MUX2_X1 U25335 ( .A(\mem[768][6] ), .B(\mem[769][6] ), .S(n8462), .Z(n6380)
         );
  MUX2_X1 U25336 ( .A(n6380), .B(n6379), .S(n8318), .Z(n6381) );
  MUX2_X1 U25337 ( .A(n6381), .B(n6378), .S(n8264), .Z(n6382) );
  MUX2_X1 U25338 ( .A(n6382), .B(n6375), .S(n8209), .Z(n6383) );
  MUX2_X1 U25339 ( .A(n6383), .B(n6368), .S(n8190), .Z(n6384) );
  MUX2_X1 U25340 ( .A(n6384), .B(n6353), .S(n8182), .Z(n6385) );
  MUX2_X1 U25341 ( .A(n6385), .B(n6322), .S(n8178), .Z(n6386) );
  MUX2_X1 U25342 ( .A(n6386), .B(n6259), .S(N25), .Z(n6387) );
  MUX2_X1 U25343 ( .A(\mem[766][6] ), .B(\mem[767][6] ), .S(n8462), .Z(n6388)
         );
  MUX2_X1 U25344 ( .A(\mem[764][6] ), .B(\mem[765][6] ), .S(n8462), .Z(n6389)
         );
  MUX2_X1 U25345 ( .A(n6389), .B(n6388), .S(n8318), .Z(n6390) );
  MUX2_X1 U25346 ( .A(\mem[762][6] ), .B(\mem[763][6] ), .S(n8462), .Z(n6391)
         );
  MUX2_X1 U25347 ( .A(\mem[760][6] ), .B(\mem[761][6] ), .S(n8462), .Z(n6392)
         );
  MUX2_X1 U25348 ( .A(n6392), .B(n6391), .S(n8318), .Z(n6393) );
  MUX2_X1 U25349 ( .A(n6393), .B(n6390), .S(n8265), .Z(n6394) );
  MUX2_X1 U25350 ( .A(\mem[758][6] ), .B(\mem[759][6] ), .S(n8462), .Z(n6395)
         );
  MUX2_X1 U25351 ( .A(\mem[756][6] ), .B(\mem[757][6] ), .S(n8462), .Z(n6396)
         );
  MUX2_X1 U25352 ( .A(n6396), .B(n6395), .S(n8318), .Z(n6397) );
  MUX2_X1 U25353 ( .A(\mem[754][6] ), .B(\mem[755][6] ), .S(n8462), .Z(n6398)
         );
  MUX2_X1 U25354 ( .A(\mem[752][6] ), .B(\mem[753][6] ), .S(n8462), .Z(n6399)
         );
  MUX2_X1 U25355 ( .A(n6399), .B(n6398), .S(n8318), .Z(n6400) );
  MUX2_X1 U25356 ( .A(n6400), .B(n6397), .S(n8261), .Z(n6401) );
  MUX2_X1 U25357 ( .A(n6401), .B(n6394), .S(n8209), .Z(n6402) );
  MUX2_X1 U25358 ( .A(\mem[750][6] ), .B(\mem[751][6] ), .S(n8463), .Z(n6403)
         );
  MUX2_X1 U25359 ( .A(\mem[748][6] ), .B(\mem[749][6] ), .S(n8463), .Z(n6404)
         );
  MUX2_X1 U25360 ( .A(n6404), .B(n6403), .S(n8319), .Z(n6405) );
  MUX2_X1 U25361 ( .A(\mem[746][6] ), .B(\mem[747][6] ), .S(n8463), .Z(n6406)
         );
  MUX2_X1 U25362 ( .A(\mem[744][6] ), .B(\mem[745][6] ), .S(n8463), .Z(n6407)
         );
  MUX2_X1 U25363 ( .A(n6407), .B(n6406), .S(n8319), .Z(n6408) );
  MUX2_X1 U25364 ( .A(n6408), .B(n6405), .S(n8235), .Z(n6409) );
  MUX2_X1 U25365 ( .A(\mem[742][6] ), .B(\mem[743][6] ), .S(n8463), .Z(n6410)
         );
  MUX2_X1 U25366 ( .A(\mem[740][6] ), .B(\mem[741][6] ), .S(n8463), .Z(n6411)
         );
  MUX2_X1 U25367 ( .A(n6411), .B(n6410), .S(n8319), .Z(n6412) );
  MUX2_X1 U25368 ( .A(\mem[738][6] ), .B(\mem[739][6] ), .S(n8463), .Z(n6413)
         );
  MUX2_X1 U25369 ( .A(\mem[736][6] ), .B(\mem[737][6] ), .S(n8463), .Z(n6414)
         );
  MUX2_X1 U25370 ( .A(n6414), .B(n6413), .S(n8319), .Z(n6415) );
  MUX2_X1 U25371 ( .A(n6415), .B(n6412), .S(n8236), .Z(n6416) );
  MUX2_X1 U25372 ( .A(n6416), .B(n6409), .S(n8209), .Z(n6417) );
  MUX2_X1 U25373 ( .A(n6417), .B(n6402), .S(n8191), .Z(n6418) );
  MUX2_X1 U25374 ( .A(\mem[734][6] ), .B(\mem[735][6] ), .S(n8463), .Z(n6419)
         );
  MUX2_X1 U25375 ( .A(\mem[732][6] ), .B(\mem[733][6] ), .S(n8463), .Z(n6420)
         );
  MUX2_X1 U25376 ( .A(n6420), .B(n6419), .S(n8319), .Z(n6421) );
  MUX2_X1 U25377 ( .A(\mem[730][6] ), .B(\mem[731][6] ), .S(n8463), .Z(n6422)
         );
  MUX2_X1 U25378 ( .A(\mem[728][6] ), .B(\mem[729][6] ), .S(n8463), .Z(n6423)
         );
  MUX2_X1 U25379 ( .A(n6423), .B(n6422), .S(n8319), .Z(n6424) );
  MUX2_X1 U25380 ( .A(n6424), .B(n6421), .S(n8237), .Z(n6425) );
  MUX2_X1 U25381 ( .A(\mem[726][6] ), .B(\mem[727][6] ), .S(n8464), .Z(n6426)
         );
  MUX2_X1 U25382 ( .A(\mem[724][6] ), .B(\mem[725][6] ), .S(n8464), .Z(n6427)
         );
  MUX2_X1 U25383 ( .A(n6427), .B(n6426), .S(n8319), .Z(n6428) );
  MUX2_X1 U25384 ( .A(\mem[722][6] ), .B(\mem[723][6] ), .S(n8464), .Z(n6429)
         );
  MUX2_X1 U25385 ( .A(\mem[720][6] ), .B(\mem[721][6] ), .S(n8464), .Z(n6430)
         );
  MUX2_X1 U25386 ( .A(n6430), .B(n6429), .S(n8319), .Z(n6431) );
  MUX2_X1 U25387 ( .A(n6431), .B(n6428), .S(n8232), .Z(n6432) );
  MUX2_X1 U25388 ( .A(n6432), .B(n6425), .S(n8209), .Z(n6433) );
  MUX2_X1 U25389 ( .A(\mem[718][6] ), .B(\mem[719][6] ), .S(n8464), .Z(n6434)
         );
  MUX2_X1 U25390 ( .A(\mem[716][6] ), .B(\mem[717][6] ), .S(n8464), .Z(n6435)
         );
  MUX2_X1 U25391 ( .A(n6435), .B(n6434), .S(n8319), .Z(n6436) );
  MUX2_X1 U25392 ( .A(\mem[714][6] ), .B(\mem[715][6] ), .S(n8464), .Z(n6437)
         );
  MUX2_X1 U25393 ( .A(\mem[712][6] ), .B(\mem[713][6] ), .S(n8464), .Z(n6438)
         );
  MUX2_X1 U25394 ( .A(n6438), .B(n6437), .S(n8319), .Z(n6439) );
  MUX2_X1 U25395 ( .A(n6439), .B(n6436), .S(n8233), .Z(n6440) );
  MUX2_X1 U25396 ( .A(\mem[710][6] ), .B(\mem[711][6] ), .S(n8464), .Z(n6441)
         );
  MUX2_X1 U25397 ( .A(\mem[708][6] ), .B(\mem[709][6] ), .S(n8464), .Z(n6442)
         );
  MUX2_X1 U25398 ( .A(n6442), .B(n6441), .S(n8319), .Z(n6443) );
  MUX2_X1 U25399 ( .A(\mem[706][6] ), .B(\mem[707][6] ), .S(n8464), .Z(n6444)
         );
  MUX2_X1 U25400 ( .A(\mem[704][6] ), .B(\mem[705][6] ), .S(n8464), .Z(n6445)
         );
  MUX2_X1 U25401 ( .A(n6445), .B(n6444), .S(n8319), .Z(n6446) );
  MUX2_X1 U25402 ( .A(n6446), .B(n6443), .S(n8234), .Z(n6447) );
  MUX2_X1 U25403 ( .A(n6447), .B(n6440), .S(n8209), .Z(n6448) );
  MUX2_X1 U25404 ( .A(n6448), .B(n6433), .S(N22), .Z(n6449) );
  MUX2_X1 U25405 ( .A(n6449), .B(n6418), .S(n8183), .Z(n6450) );
  MUX2_X1 U25406 ( .A(\mem[702][6] ), .B(\mem[703][6] ), .S(n8465), .Z(n6451)
         );
  MUX2_X1 U25407 ( .A(\mem[700][6] ), .B(\mem[701][6] ), .S(n8465), .Z(n6452)
         );
  MUX2_X1 U25408 ( .A(n6452), .B(n6451), .S(n8320), .Z(n6453) );
  MUX2_X1 U25409 ( .A(\mem[698][6] ), .B(\mem[699][6] ), .S(n8465), .Z(n6454)
         );
  MUX2_X1 U25410 ( .A(\mem[696][6] ), .B(\mem[697][6] ), .S(n8465), .Z(n6455)
         );
  MUX2_X1 U25411 ( .A(n6455), .B(n6454), .S(n8320), .Z(n6456) );
  MUX2_X1 U25412 ( .A(n6456), .B(n6453), .S(n8239), .Z(n6457) );
  MUX2_X1 U25413 ( .A(\mem[694][6] ), .B(\mem[695][6] ), .S(n8465), .Z(n6458)
         );
  MUX2_X1 U25414 ( .A(\mem[692][6] ), .B(\mem[693][6] ), .S(n8465), .Z(n6459)
         );
  MUX2_X1 U25415 ( .A(n6459), .B(n6458), .S(n8320), .Z(n6460) );
  MUX2_X1 U25416 ( .A(\mem[690][6] ), .B(\mem[691][6] ), .S(n8465), .Z(n6461)
         );
  MUX2_X1 U25417 ( .A(\mem[688][6] ), .B(\mem[689][6] ), .S(n8465), .Z(n6462)
         );
  MUX2_X1 U25418 ( .A(n6462), .B(n6461), .S(n8320), .Z(n6463) );
  MUX2_X1 U25419 ( .A(n6463), .B(n6460), .S(n8240), .Z(n6464) );
  MUX2_X1 U25420 ( .A(n6464), .B(n6457), .S(n8210), .Z(n6465) );
  MUX2_X1 U25421 ( .A(\mem[686][6] ), .B(\mem[687][6] ), .S(n8465), .Z(n6466)
         );
  MUX2_X1 U25422 ( .A(\mem[684][6] ), .B(\mem[685][6] ), .S(n8465), .Z(n6467)
         );
  MUX2_X1 U25423 ( .A(n6467), .B(n6466), .S(n8320), .Z(n6468) );
  MUX2_X1 U25424 ( .A(\mem[682][6] ), .B(\mem[683][6] ), .S(n8465), .Z(n6469)
         );
  MUX2_X1 U25425 ( .A(\mem[680][6] ), .B(\mem[681][6] ), .S(n8465), .Z(n6470)
         );
  MUX2_X1 U25426 ( .A(n6470), .B(n6469), .S(n8320), .Z(n6471) );
  MUX2_X1 U25427 ( .A(n6471), .B(n6468), .S(n8230), .Z(n6472) );
  MUX2_X1 U25428 ( .A(\mem[678][6] ), .B(\mem[679][6] ), .S(n8466), .Z(n6473)
         );
  MUX2_X1 U25429 ( .A(\mem[676][6] ), .B(\mem[677][6] ), .S(n8466), .Z(n6474)
         );
  MUX2_X1 U25430 ( .A(n6474), .B(n6473), .S(n8320), .Z(n6475) );
  MUX2_X1 U25431 ( .A(\mem[674][6] ), .B(\mem[675][6] ), .S(n8466), .Z(n6476)
         );
  MUX2_X1 U25432 ( .A(\mem[672][6] ), .B(\mem[673][6] ), .S(n8466), .Z(n6477)
         );
  MUX2_X1 U25433 ( .A(n6477), .B(n6476), .S(n8320), .Z(n6478) );
  MUX2_X1 U25434 ( .A(n6478), .B(n6475), .S(n8231), .Z(n6479) );
  MUX2_X1 U25435 ( .A(n6479), .B(n6472), .S(n8210), .Z(n6480) );
  MUX2_X1 U25436 ( .A(n6480), .B(n6465), .S(n8195), .Z(n6481) );
  MUX2_X1 U25437 ( .A(\mem[670][6] ), .B(\mem[671][6] ), .S(n8466), .Z(n6482)
         );
  MUX2_X1 U25438 ( .A(\mem[668][6] ), .B(\mem[669][6] ), .S(n8466), .Z(n6483)
         );
  MUX2_X1 U25439 ( .A(n6483), .B(n6482), .S(n8320), .Z(n6484) );
  MUX2_X1 U25440 ( .A(\mem[666][6] ), .B(\mem[667][6] ), .S(n8466), .Z(n6485)
         );
  MUX2_X1 U25441 ( .A(\mem[664][6] ), .B(\mem[665][6] ), .S(n8466), .Z(n6486)
         );
  MUX2_X1 U25442 ( .A(n6486), .B(n6485), .S(n8320), .Z(n6487) );
  MUX2_X1 U25443 ( .A(n6487), .B(n6484), .S(n8227), .Z(n6488) );
  MUX2_X1 U25444 ( .A(\mem[662][6] ), .B(\mem[663][6] ), .S(n8466), .Z(n6489)
         );
  MUX2_X1 U25445 ( .A(\mem[660][6] ), .B(\mem[661][6] ), .S(n8466), .Z(n6490)
         );
  MUX2_X1 U25446 ( .A(n6490), .B(n6489), .S(n8320), .Z(n6491) );
  MUX2_X1 U25447 ( .A(\mem[658][6] ), .B(\mem[659][6] ), .S(n8466), .Z(n6492)
         );
  MUX2_X1 U25448 ( .A(\mem[656][6] ), .B(\mem[657][6] ), .S(n8466), .Z(n6493)
         );
  MUX2_X1 U25449 ( .A(n6493), .B(n6492), .S(n8320), .Z(n6494) );
  MUX2_X1 U25450 ( .A(n6494), .B(n6491), .S(n8228), .Z(n6495) );
  MUX2_X1 U25451 ( .A(n6495), .B(n6488), .S(n8210), .Z(n6496) );
  MUX2_X1 U25452 ( .A(\mem[654][6] ), .B(\mem[655][6] ), .S(n8467), .Z(n6497)
         );
  MUX2_X1 U25453 ( .A(\mem[652][6] ), .B(\mem[653][6] ), .S(n8467), .Z(n6498)
         );
  MUX2_X1 U25454 ( .A(n6498), .B(n6497), .S(n8321), .Z(n6499) );
  MUX2_X1 U25455 ( .A(\mem[650][6] ), .B(\mem[651][6] ), .S(n8467), .Z(n6500)
         );
  MUX2_X1 U25456 ( .A(\mem[648][6] ), .B(\mem[649][6] ), .S(n8467), .Z(n6501)
         );
  MUX2_X1 U25457 ( .A(n6501), .B(n6500), .S(n8321), .Z(n6502) );
  MUX2_X1 U25458 ( .A(n6502), .B(n6499), .S(n8229), .Z(n6503) );
  MUX2_X1 U25459 ( .A(\mem[646][6] ), .B(\mem[647][6] ), .S(n8467), .Z(n6504)
         );
  MUX2_X1 U25460 ( .A(\mem[644][6] ), .B(\mem[645][6] ), .S(n8467), .Z(n6505)
         );
  MUX2_X1 U25461 ( .A(n6505), .B(n6504), .S(n8321), .Z(n6506) );
  MUX2_X1 U25462 ( .A(\mem[642][6] ), .B(\mem[643][6] ), .S(n8467), .Z(n6507)
         );
  MUX2_X1 U25463 ( .A(\mem[640][6] ), .B(\mem[641][6] ), .S(n8467), .Z(n6508)
         );
  MUX2_X1 U25464 ( .A(n6508), .B(n6507), .S(n8321), .Z(n6509) );
  MUX2_X1 U25465 ( .A(n6509), .B(n6506), .S(n8226), .Z(n6510) );
  MUX2_X1 U25466 ( .A(n6510), .B(n6503), .S(n8210), .Z(n6511) );
  MUX2_X1 U25467 ( .A(n6511), .B(n6496), .S(n8192), .Z(n6512) );
  MUX2_X1 U25468 ( .A(n6512), .B(n6481), .S(n8184), .Z(n6513) );
  MUX2_X1 U25469 ( .A(n6513), .B(n6450), .S(N24), .Z(n6514) );
  MUX2_X1 U25470 ( .A(\mem[638][6] ), .B(\mem[639][6] ), .S(n8467), .Z(n6515)
         );
  MUX2_X1 U25471 ( .A(\mem[636][6] ), .B(\mem[637][6] ), .S(n8467), .Z(n6516)
         );
  MUX2_X1 U25472 ( .A(n6516), .B(n6515), .S(n8321), .Z(n6517) );
  MUX2_X1 U25473 ( .A(\mem[634][6] ), .B(\mem[635][6] ), .S(n8467), .Z(n6518)
         );
  MUX2_X1 U25474 ( .A(\mem[632][6] ), .B(\mem[633][6] ), .S(n8467), .Z(n6519)
         );
  MUX2_X1 U25475 ( .A(n6519), .B(n6518), .S(n8321), .Z(n6520) );
  MUX2_X1 U25476 ( .A(n6520), .B(n6517), .S(n8247), .Z(n6521) );
  MUX2_X1 U25477 ( .A(\mem[630][6] ), .B(\mem[631][6] ), .S(n8468), .Z(n6522)
         );
  MUX2_X1 U25478 ( .A(\mem[628][6] ), .B(\mem[629][6] ), .S(n8468), .Z(n6523)
         );
  MUX2_X1 U25479 ( .A(n6523), .B(n6522), .S(n8321), .Z(n6524) );
  MUX2_X1 U25480 ( .A(\mem[626][6] ), .B(\mem[627][6] ), .S(n8468), .Z(n6525)
         );
  MUX2_X1 U25481 ( .A(\mem[624][6] ), .B(\mem[625][6] ), .S(n8468), .Z(n6526)
         );
  MUX2_X1 U25482 ( .A(n6526), .B(n6525), .S(n8321), .Z(n6527) );
  MUX2_X1 U25483 ( .A(n6527), .B(n6524), .S(n8248), .Z(n6528) );
  MUX2_X1 U25484 ( .A(n6528), .B(n6521), .S(n8210), .Z(n6529) );
  MUX2_X1 U25485 ( .A(\mem[622][6] ), .B(\mem[623][6] ), .S(n8468), .Z(n6530)
         );
  MUX2_X1 U25486 ( .A(\mem[620][6] ), .B(\mem[621][6] ), .S(n8468), .Z(n6531)
         );
  MUX2_X1 U25487 ( .A(n6531), .B(n6530), .S(n8321), .Z(n6532) );
  MUX2_X1 U25488 ( .A(\mem[618][6] ), .B(\mem[619][6] ), .S(n8468), .Z(n6533)
         );
  MUX2_X1 U25489 ( .A(\mem[616][6] ), .B(\mem[617][6] ), .S(n8468), .Z(n6534)
         );
  MUX2_X1 U25490 ( .A(n6534), .B(n6533), .S(n8321), .Z(n6535) );
  MUX2_X1 U25491 ( .A(n6535), .B(n6532), .S(n8249), .Z(n6536) );
  MUX2_X1 U25492 ( .A(\mem[614][6] ), .B(\mem[615][6] ), .S(n8468), .Z(n6537)
         );
  MUX2_X1 U25493 ( .A(\mem[612][6] ), .B(\mem[613][6] ), .S(n8468), .Z(n6538)
         );
  MUX2_X1 U25494 ( .A(n6538), .B(n6537), .S(n8321), .Z(n6539) );
  MUX2_X1 U25495 ( .A(\mem[610][6] ), .B(\mem[611][6] ), .S(n8468), .Z(n6540)
         );
  MUX2_X1 U25496 ( .A(\mem[608][6] ), .B(\mem[609][6] ), .S(n8468), .Z(n6541)
         );
  MUX2_X1 U25497 ( .A(n6541), .B(n6540), .S(n8321), .Z(n6542) );
  MUX2_X1 U25498 ( .A(n6542), .B(n6539), .S(n8244), .Z(n6543) );
  MUX2_X1 U25499 ( .A(n6543), .B(n6536), .S(n8210), .Z(n6544) );
  MUX2_X1 U25500 ( .A(n6544), .B(n6529), .S(n8193), .Z(n6545) );
  MUX2_X1 U25501 ( .A(\mem[606][6] ), .B(\mem[607][6] ), .S(n8469), .Z(n6546)
         );
  MUX2_X1 U25502 ( .A(\mem[604][6] ), .B(\mem[605][6] ), .S(n8469), .Z(n6547)
         );
  MUX2_X1 U25503 ( .A(n6547), .B(n6546), .S(n8322), .Z(n6548) );
  MUX2_X1 U25504 ( .A(\mem[602][6] ), .B(\mem[603][6] ), .S(n8469), .Z(n6549)
         );
  MUX2_X1 U25505 ( .A(\mem[600][6] ), .B(\mem[601][6] ), .S(n8469), .Z(n6550)
         );
  MUX2_X1 U25506 ( .A(n6550), .B(n6549), .S(n8322), .Z(n6551) );
  MUX2_X1 U25507 ( .A(n6551), .B(n6548), .S(n8229), .Z(n6552) );
  MUX2_X1 U25508 ( .A(\mem[598][6] ), .B(\mem[599][6] ), .S(n8469), .Z(n6553)
         );
  MUX2_X1 U25509 ( .A(\mem[596][6] ), .B(\mem[597][6] ), .S(n8469), .Z(n6554)
         );
  MUX2_X1 U25510 ( .A(n6554), .B(n6553), .S(n8322), .Z(n6555) );
  MUX2_X1 U25511 ( .A(\mem[594][6] ), .B(\mem[595][6] ), .S(n8469), .Z(n6556)
         );
  MUX2_X1 U25512 ( .A(\mem[592][6] ), .B(\mem[593][6] ), .S(n8469), .Z(n6557)
         );
  MUX2_X1 U25513 ( .A(n6557), .B(n6556), .S(n8322), .Z(n6558) );
  MUX2_X1 U25514 ( .A(n6558), .B(n6555), .S(n8226), .Z(n6559) );
  MUX2_X1 U25515 ( .A(n6559), .B(n6552), .S(n8210), .Z(n6560) );
  MUX2_X1 U25516 ( .A(\mem[590][6] ), .B(\mem[591][6] ), .S(n8469), .Z(n6561)
         );
  MUX2_X1 U25517 ( .A(\mem[588][6] ), .B(\mem[589][6] ), .S(n8469), .Z(n6562)
         );
  MUX2_X1 U25518 ( .A(n6562), .B(n6561), .S(n8322), .Z(n6563) );
  MUX2_X1 U25519 ( .A(\mem[586][6] ), .B(\mem[587][6] ), .S(n8469), .Z(n6564)
         );
  MUX2_X1 U25520 ( .A(\mem[584][6] ), .B(\mem[585][6] ), .S(n8469), .Z(n6565)
         );
  MUX2_X1 U25521 ( .A(n6565), .B(n6564), .S(n8322), .Z(n6566) );
  MUX2_X1 U25522 ( .A(n6566), .B(n6563), .S(n8247), .Z(n6567) );
  MUX2_X1 U25523 ( .A(\mem[582][6] ), .B(\mem[583][6] ), .S(n8470), .Z(n6568)
         );
  MUX2_X1 U25524 ( .A(\mem[580][6] ), .B(\mem[581][6] ), .S(n8470), .Z(n6569)
         );
  MUX2_X1 U25525 ( .A(n6569), .B(n6568), .S(n8322), .Z(n6570) );
  MUX2_X1 U25526 ( .A(\mem[578][6] ), .B(\mem[579][6] ), .S(n8470), .Z(n6571)
         );
  MUX2_X1 U25527 ( .A(\mem[576][6] ), .B(\mem[577][6] ), .S(n8470), .Z(n6572)
         );
  MUX2_X1 U25528 ( .A(n6572), .B(n6571), .S(n8322), .Z(n6573) );
  MUX2_X1 U25529 ( .A(n6573), .B(n6570), .S(n8248), .Z(n6574) );
  MUX2_X1 U25530 ( .A(n6574), .B(n6567), .S(n8210), .Z(n6575) );
  MUX2_X1 U25531 ( .A(n6575), .B(n6560), .S(n8196), .Z(n6576) );
  MUX2_X1 U25532 ( .A(n6576), .B(n6545), .S(n8185), .Z(n6577) );
  MUX2_X1 U25533 ( .A(\mem[574][6] ), .B(\mem[575][6] ), .S(n8470), .Z(n6578)
         );
  MUX2_X1 U25534 ( .A(\mem[572][6] ), .B(\mem[573][6] ), .S(n8470), .Z(n6579)
         );
  MUX2_X1 U25535 ( .A(n6579), .B(n6578), .S(n8322), .Z(n6580) );
  MUX2_X1 U25536 ( .A(\mem[570][6] ), .B(\mem[571][6] ), .S(n8470), .Z(n6581)
         );
  MUX2_X1 U25537 ( .A(\mem[568][6] ), .B(\mem[569][6] ), .S(n8470), .Z(n6582)
         );
  MUX2_X1 U25538 ( .A(n6582), .B(n6581), .S(n8322), .Z(n6583) );
  MUX2_X1 U25539 ( .A(n6583), .B(n6580), .S(n8249), .Z(n6584) );
  MUX2_X1 U25540 ( .A(\mem[566][6] ), .B(\mem[567][6] ), .S(n8470), .Z(n6585)
         );
  MUX2_X1 U25541 ( .A(\mem[564][6] ), .B(\mem[565][6] ), .S(n8470), .Z(n6586)
         );
  MUX2_X1 U25542 ( .A(n6586), .B(n6585), .S(n8322), .Z(n6587) );
  MUX2_X1 U25543 ( .A(\mem[562][6] ), .B(\mem[563][6] ), .S(n8470), .Z(n6588)
         );
  MUX2_X1 U25544 ( .A(\mem[560][6] ), .B(\mem[561][6] ), .S(n8470), .Z(n6589)
         );
  MUX2_X1 U25545 ( .A(n6589), .B(n6588), .S(n8322), .Z(n6590) );
  MUX2_X1 U25546 ( .A(n6590), .B(n6587), .S(n8244), .Z(n6591) );
  MUX2_X1 U25547 ( .A(n6591), .B(n6584), .S(n8210), .Z(n6592) );
  MUX2_X1 U25548 ( .A(\mem[558][6] ), .B(\mem[559][6] ), .S(n8471), .Z(n6593)
         );
  MUX2_X1 U25549 ( .A(\mem[556][6] ), .B(\mem[557][6] ), .S(n8471), .Z(n6594)
         );
  MUX2_X1 U25550 ( .A(n6594), .B(n6593), .S(n8323), .Z(n6595) );
  MUX2_X1 U25551 ( .A(\mem[554][6] ), .B(\mem[555][6] ), .S(n8471), .Z(n6596)
         );
  MUX2_X1 U25552 ( .A(\mem[552][6] ), .B(\mem[553][6] ), .S(n8471), .Z(n6597)
         );
  MUX2_X1 U25553 ( .A(n6597), .B(n6596), .S(n8323), .Z(n6598) );
  MUX2_X1 U25554 ( .A(n6598), .B(n6595), .S(n8245), .Z(n6599) );
  MUX2_X1 U25555 ( .A(\mem[550][6] ), .B(\mem[551][6] ), .S(n8471), .Z(n6600)
         );
  MUX2_X1 U25556 ( .A(\mem[548][6] ), .B(\mem[549][6] ), .S(n8471), .Z(n6601)
         );
  MUX2_X1 U25557 ( .A(n6601), .B(n6600), .S(n8323), .Z(n6602) );
  MUX2_X1 U25558 ( .A(\mem[546][6] ), .B(\mem[547][6] ), .S(n8471), .Z(n6603)
         );
  MUX2_X1 U25559 ( .A(\mem[544][6] ), .B(\mem[545][6] ), .S(n8471), .Z(n6604)
         );
  MUX2_X1 U25560 ( .A(n6604), .B(n6603), .S(n8323), .Z(n6605) );
  MUX2_X1 U25561 ( .A(n6605), .B(n6602), .S(n8246), .Z(n6606) );
  MUX2_X1 U25562 ( .A(n6606), .B(n6599), .S(n8210), .Z(n6607) );
  MUX2_X1 U25563 ( .A(n6607), .B(n6592), .S(n8189), .Z(n6608) );
  MUX2_X1 U25564 ( .A(\mem[542][6] ), .B(\mem[543][6] ), .S(n8471), .Z(n6609)
         );
  MUX2_X1 U25565 ( .A(\mem[540][6] ), .B(\mem[541][6] ), .S(n8471), .Z(n6610)
         );
  MUX2_X1 U25566 ( .A(n6610), .B(n6609), .S(n8323), .Z(n6611) );
  MUX2_X1 U25567 ( .A(\mem[538][6] ), .B(\mem[539][6] ), .S(n8471), .Z(n6612)
         );
  MUX2_X1 U25568 ( .A(\mem[536][6] ), .B(\mem[537][6] ), .S(n8471), .Z(n6613)
         );
  MUX2_X1 U25569 ( .A(n6613), .B(n6612), .S(n8323), .Z(n6614) );
  MUX2_X1 U25570 ( .A(n6614), .B(n6611), .S(n8253), .Z(n6615) );
  MUX2_X1 U25571 ( .A(\mem[534][6] ), .B(\mem[535][6] ), .S(n8472), .Z(n6616)
         );
  MUX2_X1 U25572 ( .A(\mem[532][6] ), .B(\mem[533][6] ), .S(n8472), .Z(n6617)
         );
  MUX2_X1 U25573 ( .A(n6617), .B(n6616), .S(n8323), .Z(n6618) );
  MUX2_X1 U25574 ( .A(\mem[530][6] ), .B(\mem[531][6] ), .S(n8472), .Z(n6619)
         );
  MUX2_X1 U25575 ( .A(\mem[528][6] ), .B(\mem[529][6] ), .S(n8472), .Z(n6620)
         );
  MUX2_X1 U25576 ( .A(n6620), .B(n6619), .S(n8323), .Z(n6621) );
  MUX2_X1 U25577 ( .A(n6621), .B(n6618), .S(n8254), .Z(n6622) );
  MUX2_X1 U25578 ( .A(n6622), .B(n6615), .S(n8210), .Z(n6623) );
  MUX2_X1 U25579 ( .A(\mem[526][6] ), .B(\mem[527][6] ), .S(n8472), .Z(n6624)
         );
  MUX2_X1 U25580 ( .A(\mem[524][6] ), .B(\mem[525][6] ), .S(n8472), .Z(n6625)
         );
  MUX2_X1 U25581 ( .A(n6625), .B(n6624), .S(n8323), .Z(n6626) );
  MUX2_X1 U25582 ( .A(\mem[522][6] ), .B(\mem[523][6] ), .S(n8472), .Z(n6627)
         );
  MUX2_X1 U25583 ( .A(\mem[520][6] ), .B(\mem[521][6] ), .S(n8472), .Z(n6628)
         );
  MUX2_X1 U25584 ( .A(n6628), .B(n6627), .S(n8323), .Z(n6629) );
  MUX2_X1 U25585 ( .A(n6629), .B(n6626), .S(n8255), .Z(n6630) );
  MUX2_X1 U25586 ( .A(\mem[518][6] ), .B(\mem[519][6] ), .S(n8472), .Z(n6631)
         );
  MUX2_X1 U25587 ( .A(\mem[516][6] ), .B(\mem[517][6] ), .S(n8472), .Z(n6632)
         );
  MUX2_X1 U25588 ( .A(n6632), .B(n6631), .S(n8323), .Z(n6633) );
  MUX2_X1 U25589 ( .A(\mem[514][6] ), .B(\mem[515][6] ), .S(n8472), .Z(n6634)
         );
  MUX2_X1 U25590 ( .A(\mem[512][6] ), .B(\mem[513][6] ), .S(n8472), .Z(n6635)
         );
  MUX2_X1 U25591 ( .A(n6635), .B(n6634), .S(n8323), .Z(n6636) );
  MUX2_X1 U25592 ( .A(n6636), .B(n6633), .S(n8250), .Z(n6637) );
  MUX2_X1 U25593 ( .A(n6637), .B(n6630), .S(n8210), .Z(n6638) );
  MUX2_X1 U25594 ( .A(n6638), .B(n6623), .S(n8186), .Z(n6639) );
  MUX2_X1 U25595 ( .A(n6639), .B(n6608), .S(n8184), .Z(n6640) );
  MUX2_X1 U25596 ( .A(n6640), .B(n6577), .S(n8179), .Z(n6641) );
  MUX2_X1 U25597 ( .A(n6641), .B(n6514), .S(n8177), .Z(n6642) );
  MUX2_X1 U25598 ( .A(n6642), .B(n6387), .S(N26), .Z(n6643) );
  MUX2_X1 U25599 ( .A(\mem[510][6] ), .B(\mem[511][6] ), .S(n8473), .Z(n6644)
         );
  MUX2_X1 U25600 ( .A(\mem[508][6] ), .B(\mem[509][6] ), .S(n8473), .Z(n6645)
         );
  MUX2_X1 U25601 ( .A(n6645), .B(n6644), .S(n8324), .Z(n6646) );
  MUX2_X1 U25602 ( .A(\mem[506][6] ), .B(\mem[507][6] ), .S(n8473), .Z(n6647)
         );
  MUX2_X1 U25603 ( .A(\mem[504][6] ), .B(\mem[505][6] ), .S(n8473), .Z(n6648)
         );
  MUX2_X1 U25604 ( .A(n6648), .B(n6647), .S(n8324), .Z(n6649) );
  MUX2_X1 U25605 ( .A(n6649), .B(n6646), .S(n8237), .Z(n6650) );
  MUX2_X1 U25606 ( .A(\mem[502][6] ), .B(\mem[503][6] ), .S(n8473), .Z(n6651)
         );
  MUX2_X1 U25607 ( .A(\mem[500][6] ), .B(\mem[501][6] ), .S(n8473), .Z(n6652)
         );
  MUX2_X1 U25608 ( .A(n6652), .B(n6651), .S(n8324), .Z(n6653) );
  MUX2_X1 U25609 ( .A(\mem[498][6] ), .B(\mem[499][6] ), .S(n8473), .Z(n6654)
         );
  MUX2_X1 U25610 ( .A(\mem[496][6] ), .B(\mem[497][6] ), .S(n8473), .Z(n6655)
         );
  MUX2_X1 U25611 ( .A(n6655), .B(n6654), .S(n8324), .Z(n6656) );
  MUX2_X1 U25612 ( .A(n6656), .B(n6653), .S(n8232), .Z(n6657) );
  MUX2_X1 U25613 ( .A(n6657), .B(n6650), .S(n8211), .Z(n6658) );
  MUX2_X1 U25614 ( .A(\mem[494][6] ), .B(\mem[495][6] ), .S(n8473), .Z(n6659)
         );
  MUX2_X1 U25615 ( .A(\mem[492][6] ), .B(\mem[493][6] ), .S(n8473), .Z(n6660)
         );
  MUX2_X1 U25616 ( .A(n6660), .B(n6659), .S(n8324), .Z(n6661) );
  MUX2_X1 U25617 ( .A(\mem[490][6] ), .B(\mem[491][6] ), .S(n8473), .Z(n6662)
         );
  MUX2_X1 U25618 ( .A(\mem[488][6] ), .B(\mem[489][6] ), .S(n8473), .Z(n6663)
         );
  MUX2_X1 U25619 ( .A(n6663), .B(n6662), .S(n8324), .Z(n6664) );
  MUX2_X1 U25620 ( .A(n6664), .B(n6661), .S(n8233), .Z(n6665) );
  MUX2_X1 U25621 ( .A(\mem[486][6] ), .B(\mem[487][6] ), .S(n8474), .Z(n6666)
         );
  MUX2_X1 U25622 ( .A(\mem[484][6] ), .B(\mem[485][6] ), .S(n8474), .Z(n6667)
         );
  MUX2_X1 U25623 ( .A(n6667), .B(n6666), .S(n8324), .Z(n6668) );
  MUX2_X1 U25624 ( .A(\mem[482][6] ), .B(\mem[483][6] ), .S(n8474), .Z(n6669)
         );
  MUX2_X1 U25625 ( .A(\mem[480][6] ), .B(\mem[481][6] ), .S(n8474), .Z(n6670)
         );
  MUX2_X1 U25626 ( .A(n6670), .B(n6669), .S(n8324), .Z(n6671) );
  MUX2_X1 U25627 ( .A(n6671), .B(n6668), .S(n8234), .Z(n6672) );
  MUX2_X1 U25628 ( .A(n6672), .B(n6665), .S(n8211), .Z(n6673) );
  MUX2_X1 U25629 ( .A(n6673), .B(n6658), .S(n8191), .Z(n6674) );
  MUX2_X1 U25630 ( .A(\mem[478][6] ), .B(\mem[479][6] ), .S(n8474), .Z(n6675)
         );
  MUX2_X1 U25631 ( .A(\mem[476][6] ), .B(\mem[477][6] ), .S(n8474), .Z(n6676)
         );
  MUX2_X1 U25632 ( .A(n6676), .B(n6675), .S(n8324), .Z(n6677) );
  MUX2_X1 U25633 ( .A(\mem[474][6] ), .B(\mem[475][6] ), .S(n8474), .Z(n6678)
         );
  MUX2_X1 U25634 ( .A(\mem[472][6] ), .B(\mem[473][6] ), .S(n8474), .Z(n6679)
         );
  MUX2_X1 U25635 ( .A(n6679), .B(n6678), .S(n8324), .Z(n6680) );
  MUX2_X1 U25636 ( .A(n6680), .B(n6677), .S(n8241), .Z(n6681) );
  MUX2_X1 U25637 ( .A(\mem[470][6] ), .B(\mem[471][6] ), .S(n8474), .Z(n6682)
         );
  MUX2_X1 U25638 ( .A(\mem[468][6] ), .B(\mem[469][6] ), .S(n8474), .Z(n6683)
         );
  MUX2_X1 U25639 ( .A(n6683), .B(n6682), .S(n8324), .Z(n6684) );
  MUX2_X1 U25640 ( .A(\mem[466][6] ), .B(\mem[467][6] ), .S(n8474), .Z(n6685)
         );
  MUX2_X1 U25641 ( .A(\mem[464][6] ), .B(\mem[465][6] ), .S(n8474), .Z(n6686)
         );
  MUX2_X1 U25642 ( .A(n6686), .B(n6685), .S(n8324), .Z(n6687) );
  MUX2_X1 U25643 ( .A(n6687), .B(n6684), .S(n8242), .Z(n6688) );
  MUX2_X1 U25644 ( .A(n6688), .B(n6681), .S(n8211), .Z(n6689) );
  MUX2_X1 U25645 ( .A(\mem[462][6] ), .B(\mem[463][6] ), .S(n8475), .Z(n6690)
         );
  MUX2_X1 U25646 ( .A(\mem[460][6] ), .B(\mem[461][6] ), .S(n8475), .Z(n6691)
         );
  MUX2_X1 U25647 ( .A(n6691), .B(n6690), .S(n8325), .Z(n6692) );
  MUX2_X1 U25648 ( .A(\mem[458][6] ), .B(\mem[459][6] ), .S(n8475), .Z(n6693)
         );
  MUX2_X1 U25649 ( .A(\mem[456][6] ), .B(\mem[457][6] ), .S(n8475), .Z(n6694)
         );
  MUX2_X1 U25650 ( .A(n6694), .B(n6693), .S(n8325), .Z(n6695) );
  MUX2_X1 U25651 ( .A(n6695), .B(n6692), .S(n8243), .Z(n6696) );
  MUX2_X1 U25652 ( .A(\mem[454][6] ), .B(\mem[455][6] ), .S(n8475), .Z(n6697)
         );
  MUX2_X1 U25653 ( .A(\mem[452][6] ), .B(\mem[453][6] ), .S(n8475), .Z(n6698)
         );
  MUX2_X1 U25654 ( .A(n6698), .B(n6697), .S(n8325), .Z(n6699) );
  MUX2_X1 U25655 ( .A(\mem[450][6] ), .B(\mem[451][6] ), .S(n8475), .Z(n6700)
         );
  MUX2_X1 U25656 ( .A(\mem[448][6] ), .B(\mem[449][6] ), .S(n8475), .Z(n6701)
         );
  MUX2_X1 U25657 ( .A(n6701), .B(n6700), .S(n8325), .Z(n6702) );
  MUX2_X1 U25658 ( .A(n6702), .B(n6699), .S(n8238), .Z(n6703) );
  MUX2_X1 U25659 ( .A(n6703), .B(n6696), .S(n8211), .Z(n6704) );
  MUX2_X1 U25660 ( .A(n6704), .B(n6689), .S(n8191), .Z(n6705) );
  MUX2_X1 U25661 ( .A(n6705), .B(n6674), .S(n8185), .Z(n6706) );
  MUX2_X1 U25662 ( .A(\mem[446][6] ), .B(\mem[447][6] ), .S(n8475), .Z(n6707)
         );
  MUX2_X1 U25663 ( .A(\mem[444][6] ), .B(\mem[445][6] ), .S(n8475), .Z(n6708)
         );
  MUX2_X1 U25664 ( .A(n6708), .B(n6707), .S(n8325), .Z(n6709) );
  MUX2_X1 U25665 ( .A(\mem[442][6] ), .B(\mem[443][6] ), .S(n8475), .Z(n6710)
         );
  MUX2_X1 U25666 ( .A(\mem[440][6] ), .B(\mem[441][6] ), .S(n8475), .Z(n6711)
         );
  MUX2_X1 U25667 ( .A(n6711), .B(n6710), .S(n8325), .Z(n6712) );
  MUX2_X1 U25668 ( .A(n6712), .B(n6709), .S(n8239), .Z(n6713) );
  MUX2_X1 U25669 ( .A(\mem[438][6] ), .B(\mem[439][6] ), .S(n8476), .Z(n6714)
         );
  MUX2_X1 U25670 ( .A(\mem[436][6] ), .B(\mem[437][6] ), .S(n8476), .Z(n6715)
         );
  MUX2_X1 U25671 ( .A(n6715), .B(n6714), .S(n8325), .Z(n6716) );
  MUX2_X1 U25672 ( .A(\mem[434][6] ), .B(\mem[435][6] ), .S(n8476), .Z(n6717)
         );
  MUX2_X1 U25673 ( .A(\mem[432][6] ), .B(\mem[433][6] ), .S(n8476), .Z(n6718)
         );
  MUX2_X1 U25674 ( .A(n6718), .B(n6717), .S(n8325), .Z(n6719) );
  MUX2_X1 U25675 ( .A(n6719), .B(n6716), .S(n8240), .Z(n6720) );
  MUX2_X1 U25676 ( .A(n6720), .B(n6713), .S(n8211), .Z(n6721) );
  MUX2_X1 U25677 ( .A(\mem[430][6] ), .B(\mem[431][6] ), .S(n8476), .Z(n6722)
         );
  MUX2_X1 U25678 ( .A(\mem[428][6] ), .B(\mem[429][6] ), .S(n8476), .Z(n6723)
         );
  MUX2_X1 U25679 ( .A(n6723), .B(n6722), .S(n8325), .Z(n6724) );
  MUX2_X1 U25680 ( .A(\mem[426][6] ), .B(\mem[427][6] ), .S(n8476), .Z(n6725)
         );
  MUX2_X1 U25681 ( .A(\mem[424][6] ), .B(\mem[425][6] ), .S(n8476), .Z(n6726)
         );
  MUX2_X1 U25682 ( .A(n6726), .B(n6725), .S(n8325), .Z(n6727) );
  MUX2_X1 U25683 ( .A(n6727), .B(n6724), .S(n8230), .Z(n6728) );
  MUX2_X1 U25684 ( .A(\mem[422][6] ), .B(\mem[423][6] ), .S(n8476), .Z(n6729)
         );
  MUX2_X1 U25685 ( .A(\mem[420][6] ), .B(\mem[421][6] ), .S(n8476), .Z(n6730)
         );
  MUX2_X1 U25686 ( .A(n6730), .B(n6729), .S(n8325), .Z(n6731) );
  MUX2_X1 U25687 ( .A(\mem[418][6] ), .B(\mem[419][6] ), .S(n8476), .Z(n6732)
         );
  MUX2_X1 U25688 ( .A(\mem[416][6] ), .B(\mem[417][6] ), .S(n8476), .Z(n6733)
         );
  MUX2_X1 U25689 ( .A(n6733), .B(n6732), .S(n8325), .Z(n6734) );
  MUX2_X1 U25690 ( .A(n6734), .B(n6731), .S(n8231), .Z(n6735) );
  MUX2_X1 U25691 ( .A(n6735), .B(n6728), .S(n8211), .Z(n6736) );
  MUX2_X1 U25692 ( .A(n6736), .B(n6721), .S(n8191), .Z(n6737) );
  MUX2_X1 U25693 ( .A(\mem[414][6] ), .B(\mem[415][6] ), .S(n8477), .Z(n6738)
         );
  MUX2_X1 U25694 ( .A(\mem[412][6] ), .B(\mem[413][6] ), .S(n8477), .Z(n6739)
         );
  MUX2_X1 U25695 ( .A(n6739), .B(n6738), .S(n8326), .Z(n6740) );
  MUX2_X1 U25696 ( .A(\mem[410][6] ), .B(\mem[411][6] ), .S(n8477), .Z(n6741)
         );
  MUX2_X1 U25697 ( .A(\mem[408][6] ), .B(\mem[409][6] ), .S(n8477), .Z(n6742)
         );
  MUX2_X1 U25698 ( .A(n6742), .B(n6741), .S(n8326), .Z(n6743) );
  MUX2_X1 U25699 ( .A(n6743), .B(n6740), .S(n8261), .Z(n6744) );
  MUX2_X1 U25700 ( .A(\mem[406][6] ), .B(\mem[407][6] ), .S(n8477), .Z(n6745)
         );
  MUX2_X1 U25701 ( .A(\mem[404][6] ), .B(\mem[405][6] ), .S(n8477), .Z(n6746)
         );
  MUX2_X1 U25702 ( .A(n6746), .B(n6745), .S(n8326), .Z(n6747) );
  MUX2_X1 U25703 ( .A(\mem[402][6] ), .B(\mem[403][6] ), .S(n8477), .Z(n6748)
         );
  MUX2_X1 U25704 ( .A(\mem[400][6] ), .B(\mem[401][6] ), .S(n8477), .Z(n6749)
         );
  MUX2_X1 U25705 ( .A(n6749), .B(n6748), .S(n8326), .Z(n6750) );
  MUX2_X1 U25706 ( .A(n6750), .B(n6747), .S(n8225), .Z(n6751) );
  MUX2_X1 U25707 ( .A(n6751), .B(n6744), .S(n8211), .Z(n6752) );
  MUX2_X1 U25708 ( .A(\mem[398][6] ), .B(\mem[399][6] ), .S(n8477), .Z(n6753)
         );
  MUX2_X1 U25709 ( .A(\mem[396][6] ), .B(\mem[397][6] ), .S(n8477), .Z(n6754)
         );
  MUX2_X1 U25710 ( .A(n6754), .B(n6753), .S(n8326), .Z(n6755) );
  MUX2_X1 U25711 ( .A(\mem[394][6] ), .B(\mem[395][6] ), .S(n8477), .Z(n6756)
         );
  MUX2_X1 U25712 ( .A(\mem[392][6] ), .B(\mem[393][6] ), .S(n8477), .Z(n6757)
         );
  MUX2_X1 U25713 ( .A(n6757), .B(n6756), .S(n8326), .Z(n6758) );
  MUX2_X1 U25714 ( .A(n6758), .B(n6755), .S(n8249), .Z(n6759) );
  MUX2_X1 U25715 ( .A(\mem[390][6] ), .B(\mem[391][6] ), .S(n8478), .Z(n6760)
         );
  MUX2_X1 U25716 ( .A(\mem[388][6] ), .B(\mem[389][6] ), .S(n8478), .Z(n6761)
         );
  MUX2_X1 U25717 ( .A(n6761), .B(n6760), .S(n8326), .Z(n6762) );
  MUX2_X1 U25718 ( .A(\mem[386][6] ), .B(\mem[387][6] ), .S(n8478), .Z(n6763)
         );
  MUX2_X1 U25719 ( .A(\mem[384][6] ), .B(\mem[385][6] ), .S(n8478), .Z(n6764)
         );
  MUX2_X1 U25720 ( .A(n6764), .B(n6763), .S(n8326), .Z(n6765) );
  MUX2_X1 U25721 ( .A(n6765), .B(n6762), .S(n8224), .Z(n6766) );
  MUX2_X1 U25722 ( .A(n6766), .B(n6759), .S(n8211), .Z(n6767) );
  MUX2_X1 U25723 ( .A(n6767), .B(n6752), .S(n8191), .Z(n6768) );
  MUX2_X1 U25724 ( .A(n6768), .B(n6737), .S(N23), .Z(n6769) );
  MUX2_X1 U25725 ( .A(n6769), .B(n6706), .S(n8180), .Z(n6770) );
  MUX2_X1 U25726 ( .A(\mem[382][6] ), .B(\mem[383][6] ), .S(n8478), .Z(n6771)
         );
  MUX2_X1 U25727 ( .A(\mem[380][6] ), .B(\mem[381][6] ), .S(n8478), .Z(n6772)
         );
  MUX2_X1 U25728 ( .A(n6772), .B(n6771), .S(n8326), .Z(n6773) );
  MUX2_X1 U25729 ( .A(\mem[378][6] ), .B(\mem[379][6] ), .S(n8478), .Z(n6774)
         );
  MUX2_X1 U25730 ( .A(\mem[376][6] ), .B(\mem[377][6] ), .S(n8478), .Z(n6775)
         );
  MUX2_X1 U25731 ( .A(n6775), .B(n6774), .S(n8326), .Z(n6776) );
  MUX2_X1 U25732 ( .A(n6776), .B(n6773), .S(n8223), .Z(n6777) );
  MUX2_X1 U25733 ( .A(\mem[374][6] ), .B(\mem[375][6] ), .S(n8478), .Z(n6778)
         );
  MUX2_X1 U25734 ( .A(\mem[372][6] ), .B(\mem[373][6] ), .S(n8478), .Z(n6779)
         );
  MUX2_X1 U25735 ( .A(n6779), .B(n6778), .S(n8326), .Z(n6780) );
  MUX2_X1 U25736 ( .A(\mem[370][6] ), .B(\mem[371][6] ), .S(n8478), .Z(n6781)
         );
  MUX2_X1 U25737 ( .A(\mem[368][6] ), .B(\mem[369][6] ), .S(n8478), .Z(n6782)
         );
  MUX2_X1 U25738 ( .A(n6782), .B(n6781), .S(n8326), .Z(n6783) );
  MUX2_X1 U25739 ( .A(n6783), .B(n6780), .S(n8222), .Z(n6784) );
  MUX2_X1 U25740 ( .A(n6784), .B(n6777), .S(n8211), .Z(n6785) );
  MUX2_X1 U25741 ( .A(\mem[366][6] ), .B(\mem[367][6] ), .S(n8479), .Z(n6786)
         );
  MUX2_X1 U25742 ( .A(\mem[364][6] ), .B(\mem[365][6] ), .S(n8479), .Z(n6787)
         );
  MUX2_X1 U25743 ( .A(n6787), .B(n6786), .S(n8327), .Z(n6788) );
  MUX2_X1 U25744 ( .A(\mem[362][6] ), .B(\mem[363][6] ), .S(n8479), .Z(n6789)
         );
  MUX2_X1 U25745 ( .A(\mem[360][6] ), .B(\mem[361][6] ), .S(n8479), .Z(n6790)
         );
  MUX2_X1 U25746 ( .A(n6790), .B(n6789), .S(n8327), .Z(n6791) );
  MUX2_X1 U25747 ( .A(n6791), .B(n6788), .S(n8221), .Z(n6792) );
  MUX2_X1 U25748 ( .A(\mem[358][6] ), .B(\mem[359][6] ), .S(n8479), .Z(n6793)
         );
  MUX2_X1 U25749 ( .A(\mem[356][6] ), .B(\mem[357][6] ), .S(n8479), .Z(n6794)
         );
  MUX2_X1 U25750 ( .A(n6794), .B(n6793), .S(n8327), .Z(n6795) );
  MUX2_X1 U25751 ( .A(\mem[354][6] ), .B(\mem[355][6] ), .S(n8479), .Z(n6796)
         );
  MUX2_X1 U25752 ( .A(\mem[352][6] ), .B(\mem[353][6] ), .S(n8479), .Z(n6797)
         );
  MUX2_X1 U25753 ( .A(n6797), .B(n6796), .S(n8327), .Z(n6798) );
  MUX2_X1 U25754 ( .A(n6798), .B(n6795), .S(n8220), .Z(n6799) );
  MUX2_X1 U25755 ( .A(n6799), .B(n6792), .S(n8211), .Z(n6800) );
  MUX2_X1 U25756 ( .A(n6800), .B(n6785), .S(n8191), .Z(n6801) );
  MUX2_X1 U25757 ( .A(\mem[350][6] ), .B(\mem[351][6] ), .S(n8479), .Z(n6802)
         );
  MUX2_X1 U25758 ( .A(\mem[348][6] ), .B(\mem[349][6] ), .S(n8479), .Z(n6803)
         );
  MUX2_X1 U25759 ( .A(n6803), .B(n6802), .S(n8327), .Z(n6804) );
  MUX2_X1 U25760 ( .A(\mem[346][6] ), .B(\mem[347][6] ), .S(n8479), .Z(n6805)
         );
  MUX2_X1 U25761 ( .A(\mem[344][6] ), .B(\mem[345][6] ), .S(n8479), .Z(n6806)
         );
  MUX2_X1 U25762 ( .A(n6806), .B(n6805), .S(n8327), .Z(n6807) );
  MUX2_X1 U25763 ( .A(n6807), .B(n6804), .S(N20), .Z(n6808) );
  MUX2_X1 U25764 ( .A(\mem[342][6] ), .B(\mem[343][6] ), .S(n8480), .Z(n6809)
         );
  MUX2_X1 U25765 ( .A(\mem[340][6] ), .B(\mem[341][6] ), .S(n8480), .Z(n6810)
         );
  MUX2_X1 U25766 ( .A(n6810), .B(n6809), .S(n8327), .Z(n6811) );
  MUX2_X1 U25767 ( .A(\mem[338][6] ), .B(\mem[339][6] ), .S(n8480), .Z(n6812)
         );
  MUX2_X1 U25768 ( .A(\mem[336][6] ), .B(\mem[337][6] ), .S(n8480), .Z(n6813)
         );
  MUX2_X1 U25769 ( .A(n6813), .B(n6812), .S(n8327), .Z(n6814) );
  MUX2_X1 U25770 ( .A(n6814), .B(n6811), .S(n8265), .Z(n6815) );
  MUX2_X1 U25771 ( .A(n6815), .B(n6808), .S(n8211), .Z(n6816) );
  MUX2_X1 U25772 ( .A(\mem[334][6] ), .B(\mem[335][6] ), .S(n8480), .Z(n6817)
         );
  MUX2_X1 U25773 ( .A(\mem[332][6] ), .B(\mem[333][6] ), .S(n8480), .Z(n6818)
         );
  MUX2_X1 U25774 ( .A(n6818), .B(n6817), .S(n8327), .Z(n6819) );
  MUX2_X1 U25775 ( .A(\mem[330][6] ), .B(\mem[331][6] ), .S(n8480), .Z(n6820)
         );
  MUX2_X1 U25776 ( .A(\mem[328][6] ), .B(\mem[329][6] ), .S(n8480), .Z(n6821)
         );
  MUX2_X1 U25777 ( .A(n6821), .B(n6820), .S(n8327), .Z(n6822) );
  MUX2_X1 U25778 ( .A(n6822), .B(n6819), .S(n8265), .Z(n6823) );
  MUX2_X1 U25779 ( .A(\mem[326][6] ), .B(\mem[327][6] ), .S(n8480), .Z(n6824)
         );
  MUX2_X1 U25780 ( .A(\mem[324][6] ), .B(\mem[325][6] ), .S(n8480), .Z(n6825)
         );
  MUX2_X1 U25781 ( .A(n6825), .B(n6824), .S(n8327), .Z(n6826) );
  MUX2_X1 U25782 ( .A(\mem[322][6] ), .B(\mem[323][6] ), .S(n8480), .Z(n6827)
         );
  MUX2_X1 U25783 ( .A(\mem[320][6] ), .B(\mem[321][6] ), .S(n8480), .Z(n6828)
         );
  MUX2_X1 U25784 ( .A(n6828), .B(n6827), .S(n8327), .Z(n6829) );
  MUX2_X1 U25785 ( .A(n6829), .B(n6826), .S(n8225), .Z(n6830) );
  MUX2_X1 U25786 ( .A(n6830), .B(n6823), .S(n8211), .Z(n6831) );
  MUX2_X1 U25787 ( .A(n6831), .B(n6816), .S(n8191), .Z(n6832) );
  MUX2_X1 U25788 ( .A(n6832), .B(n6801), .S(n8185), .Z(n6833) );
  MUX2_X1 U25789 ( .A(\mem[318][6] ), .B(\mem[319][6] ), .S(n8481), .Z(n6834)
         );
  MUX2_X1 U25790 ( .A(\mem[316][6] ), .B(\mem[317][6] ), .S(n8481), .Z(n6835)
         );
  MUX2_X1 U25791 ( .A(n6835), .B(n6834), .S(n8328), .Z(n6836) );
  MUX2_X1 U25792 ( .A(\mem[314][6] ), .B(\mem[315][6] ), .S(n8481), .Z(n6837)
         );
  MUX2_X1 U25793 ( .A(\mem[312][6] ), .B(\mem[313][6] ), .S(n8481), .Z(n6838)
         );
  MUX2_X1 U25794 ( .A(n6838), .B(n6837), .S(n8328), .Z(n6839) );
  MUX2_X1 U25795 ( .A(n6839), .B(n6836), .S(n8254), .Z(n6840) );
  MUX2_X1 U25796 ( .A(\mem[310][6] ), .B(\mem[311][6] ), .S(n8481), .Z(n6841)
         );
  MUX2_X1 U25797 ( .A(\mem[308][6] ), .B(\mem[309][6] ), .S(n8481), .Z(n6842)
         );
  MUX2_X1 U25798 ( .A(n6842), .B(n6841), .S(n8328), .Z(n6843) );
  MUX2_X1 U25799 ( .A(\mem[306][6] ), .B(\mem[307][6] ), .S(n8481), .Z(n6844)
         );
  MUX2_X1 U25800 ( .A(\mem[304][6] ), .B(\mem[305][6] ), .S(n8481), .Z(n6845)
         );
  MUX2_X1 U25801 ( .A(n6845), .B(n6844), .S(n8328), .Z(n6846) );
  MUX2_X1 U25802 ( .A(n6846), .B(n6843), .S(n8255), .Z(n6847) );
  MUX2_X1 U25803 ( .A(n6847), .B(n6840), .S(n8212), .Z(n6848) );
  MUX2_X1 U25804 ( .A(\mem[302][6] ), .B(\mem[303][6] ), .S(n8481), .Z(n6849)
         );
  MUX2_X1 U25805 ( .A(\mem[300][6] ), .B(\mem[301][6] ), .S(n8481), .Z(n6850)
         );
  MUX2_X1 U25806 ( .A(n6850), .B(n6849), .S(n8328), .Z(n6851) );
  MUX2_X1 U25807 ( .A(\mem[298][6] ), .B(\mem[299][6] ), .S(n8481), .Z(n6852)
         );
  MUX2_X1 U25808 ( .A(\mem[296][6] ), .B(\mem[297][6] ), .S(n8481), .Z(n6853)
         );
  MUX2_X1 U25809 ( .A(n6853), .B(n6852), .S(n8328), .Z(n6854) );
  MUX2_X1 U25810 ( .A(n6854), .B(n6851), .S(n8250), .Z(n6855) );
  MUX2_X1 U25811 ( .A(\mem[294][6] ), .B(\mem[295][6] ), .S(n8482), .Z(n6856)
         );
  MUX2_X1 U25812 ( .A(\mem[292][6] ), .B(\mem[293][6] ), .S(n8482), .Z(n6857)
         );
  MUX2_X1 U25813 ( .A(n6857), .B(n6856), .S(n8328), .Z(n6858) );
  MUX2_X1 U25814 ( .A(\mem[290][6] ), .B(\mem[291][6] ), .S(n8482), .Z(n6859)
         );
  MUX2_X1 U25815 ( .A(\mem[288][6] ), .B(\mem[289][6] ), .S(n8482), .Z(n6860)
         );
  MUX2_X1 U25816 ( .A(n6860), .B(n6859), .S(n8328), .Z(n6861) );
  MUX2_X1 U25817 ( .A(n6861), .B(n6858), .S(n8251), .Z(n6862) );
  MUX2_X1 U25818 ( .A(n6862), .B(n6855), .S(n8212), .Z(n6863) );
  MUX2_X1 U25819 ( .A(n6863), .B(n6848), .S(n8191), .Z(n6864) );
  MUX2_X1 U25820 ( .A(\mem[286][6] ), .B(\mem[287][6] ), .S(n8482), .Z(n6865)
         );
  MUX2_X1 U25821 ( .A(\mem[284][6] ), .B(\mem[285][6] ), .S(n8482), .Z(n6866)
         );
  MUX2_X1 U25822 ( .A(n6866), .B(n6865), .S(n8328), .Z(n6867) );
  MUX2_X1 U25823 ( .A(\mem[282][6] ), .B(\mem[283][6] ), .S(n8482), .Z(n6868)
         );
  MUX2_X1 U25824 ( .A(\mem[280][6] ), .B(\mem[281][6] ), .S(n8482), .Z(n6869)
         );
  MUX2_X1 U25825 ( .A(n6869), .B(n6868), .S(n8328), .Z(n6870) );
  MUX2_X1 U25826 ( .A(n6870), .B(n6867), .S(n8252), .Z(n6871) );
  MUX2_X1 U25827 ( .A(\mem[278][6] ), .B(\mem[279][6] ), .S(n8482), .Z(n6872)
         );
  MUX2_X1 U25828 ( .A(\mem[276][6] ), .B(\mem[277][6] ), .S(n8482), .Z(n6873)
         );
  MUX2_X1 U25829 ( .A(n6873), .B(n6872), .S(n8328), .Z(n6874) );
  MUX2_X1 U25830 ( .A(\mem[274][6] ), .B(\mem[275][6] ), .S(n8482), .Z(n6875)
         );
  MUX2_X1 U25831 ( .A(\mem[272][6] ), .B(\mem[273][6] ), .S(n8482), .Z(n6876)
         );
  MUX2_X1 U25832 ( .A(n6876), .B(n6875), .S(n8328), .Z(n6877) );
  MUX2_X1 U25833 ( .A(n6877), .B(n6874), .S(n8259), .Z(n6878) );
  MUX2_X1 U25834 ( .A(n6878), .B(n6871), .S(n8212), .Z(n6879) );
  MUX2_X1 U25835 ( .A(\mem[270][6] ), .B(\mem[271][6] ), .S(n8483), .Z(n6880)
         );
  MUX2_X1 U25836 ( .A(\mem[268][6] ), .B(\mem[269][6] ), .S(n8483), .Z(n6881)
         );
  MUX2_X1 U25837 ( .A(n6881), .B(n6880), .S(n8329), .Z(n6882) );
  MUX2_X1 U25838 ( .A(\mem[266][6] ), .B(\mem[267][6] ), .S(n8483), .Z(n6883)
         );
  MUX2_X1 U25839 ( .A(\mem[264][6] ), .B(\mem[265][6] ), .S(n8483), .Z(n6884)
         );
  MUX2_X1 U25840 ( .A(n6884), .B(n6883), .S(n8329), .Z(n6885) );
  MUX2_X1 U25841 ( .A(n6885), .B(n6882), .S(n8260), .Z(n6886) );
  MUX2_X1 U25842 ( .A(\mem[262][6] ), .B(\mem[263][6] ), .S(n8483), .Z(n6887)
         );
  MUX2_X1 U25843 ( .A(\mem[260][6] ), .B(\mem[261][6] ), .S(n8483), .Z(n6888)
         );
  MUX2_X1 U25844 ( .A(n6888), .B(n6887), .S(n8329), .Z(n6889) );
  MUX2_X1 U25845 ( .A(\mem[258][6] ), .B(\mem[259][6] ), .S(n8483), .Z(n6890)
         );
  MUX2_X1 U25846 ( .A(\mem[256][6] ), .B(\mem[257][6] ), .S(n8483), .Z(n6891)
         );
  MUX2_X1 U25847 ( .A(n6891), .B(n6890), .S(n8329), .Z(n6892) );
  MUX2_X1 U25848 ( .A(n6892), .B(n6889), .S(n8261), .Z(n6893) );
  MUX2_X1 U25849 ( .A(n6893), .B(n6886), .S(n8212), .Z(n6894) );
  MUX2_X1 U25850 ( .A(n6894), .B(n6879), .S(n8191), .Z(n6895) );
  MUX2_X1 U25851 ( .A(n6895), .B(n6864), .S(n8181), .Z(n6896) );
  MUX2_X1 U25852 ( .A(n6896), .B(n6833), .S(n8180), .Z(n6897) );
  MUX2_X1 U25853 ( .A(n6897), .B(n6770), .S(N25), .Z(n6898) );
  MUX2_X1 U25854 ( .A(\mem[254][6] ), .B(\mem[255][6] ), .S(n8483), .Z(n6899)
         );
  MUX2_X1 U25855 ( .A(\mem[252][6] ), .B(\mem[253][6] ), .S(n8483), .Z(n6900)
         );
  MUX2_X1 U25856 ( .A(n6900), .B(n6899), .S(n8329), .Z(n6901) );
  MUX2_X1 U25857 ( .A(\mem[250][6] ), .B(\mem[251][6] ), .S(n8483), .Z(n6902)
         );
  MUX2_X1 U25858 ( .A(\mem[248][6] ), .B(\mem[249][6] ), .S(n8483), .Z(n6903)
         );
  MUX2_X1 U25859 ( .A(n6903), .B(n6902), .S(n8329), .Z(n6904) );
  MUX2_X1 U25860 ( .A(n6904), .B(n6901), .S(n8256), .Z(n6905) );
  MUX2_X1 U25861 ( .A(\mem[246][6] ), .B(\mem[247][6] ), .S(n8484), .Z(n6906)
         );
  MUX2_X1 U25862 ( .A(\mem[244][6] ), .B(\mem[245][6] ), .S(n8484), .Z(n6907)
         );
  MUX2_X1 U25863 ( .A(n6907), .B(n6906), .S(n8329), .Z(n6908) );
  MUX2_X1 U25864 ( .A(\mem[242][6] ), .B(\mem[243][6] ), .S(n8484), .Z(n6909)
         );
  MUX2_X1 U25865 ( .A(\mem[240][6] ), .B(\mem[241][6] ), .S(n8484), .Z(n6910)
         );
  MUX2_X1 U25866 ( .A(n6910), .B(n6909), .S(n8329), .Z(n6911) );
  MUX2_X1 U25867 ( .A(n6911), .B(n6908), .S(n8257), .Z(n6912) );
  MUX2_X1 U25868 ( .A(n6912), .B(n6905), .S(n8212), .Z(n6913) );
  MUX2_X1 U25869 ( .A(\mem[238][6] ), .B(\mem[239][6] ), .S(n8484), .Z(n6914)
         );
  MUX2_X1 U25870 ( .A(\mem[236][6] ), .B(\mem[237][6] ), .S(n8484), .Z(n6915)
         );
  MUX2_X1 U25871 ( .A(n6915), .B(n6914), .S(n8329), .Z(n6916) );
  MUX2_X1 U25872 ( .A(\mem[234][6] ), .B(\mem[235][6] ), .S(n8484), .Z(n6917)
         );
  MUX2_X1 U25873 ( .A(\mem[232][6] ), .B(\mem[233][6] ), .S(n8484), .Z(n6918)
         );
  MUX2_X1 U25874 ( .A(n6918), .B(n6917), .S(n8329), .Z(n6919) );
  MUX2_X1 U25875 ( .A(n6919), .B(n6916), .S(n8258), .Z(n6920) );
  MUX2_X1 U25876 ( .A(\mem[230][6] ), .B(\mem[231][6] ), .S(n8484), .Z(n6921)
         );
  MUX2_X1 U25877 ( .A(\mem[228][6] ), .B(\mem[229][6] ), .S(n8484), .Z(n6922)
         );
  MUX2_X1 U25878 ( .A(n6922), .B(n6921), .S(n8329), .Z(n6923) );
  MUX2_X1 U25879 ( .A(\mem[226][6] ), .B(\mem[227][6] ), .S(n8484), .Z(n6924)
         );
  MUX2_X1 U25880 ( .A(\mem[224][6] ), .B(\mem[225][6] ), .S(n8484), .Z(n6925)
         );
  MUX2_X1 U25881 ( .A(n6925), .B(n6924), .S(n8329), .Z(n6926) );
  MUX2_X1 U25882 ( .A(n6926), .B(n6923), .S(n8245), .Z(n6927) );
  MUX2_X1 U25883 ( .A(n6927), .B(n6920), .S(n8212), .Z(n6928) );
  MUX2_X1 U25884 ( .A(n6928), .B(n6913), .S(n8191), .Z(n6929) );
  MUX2_X1 U25885 ( .A(\mem[222][6] ), .B(\mem[223][6] ), .S(n8485), .Z(n6930)
         );
  MUX2_X1 U25886 ( .A(\mem[220][6] ), .B(\mem[221][6] ), .S(n8485), .Z(n6931)
         );
  MUX2_X1 U25887 ( .A(n6931), .B(n6930), .S(n8330), .Z(n6932) );
  MUX2_X1 U25888 ( .A(\mem[218][6] ), .B(\mem[219][6] ), .S(n8485), .Z(n6933)
         );
  MUX2_X1 U25889 ( .A(\mem[216][6] ), .B(\mem[217][6] ), .S(n8485), .Z(n6934)
         );
  MUX2_X1 U25890 ( .A(n6934), .B(n6933), .S(n8330), .Z(n6935) );
  MUX2_X1 U25891 ( .A(n6935), .B(n6932), .S(n8239), .Z(n6936) );
  MUX2_X1 U25892 ( .A(\mem[214][6] ), .B(\mem[215][6] ), .S(n8485), .Z(n6937)
         );
  MUX2_X1 U25893 ( .A(\mem[212][6] ), .B(\mem[213][6] ), .S(n8485), .Z(n6938)
         );
  MUX2_X1 U25894 ( .A(n6938), .B(n6937), .S(n8330), .Z(n6939) );
  MUX2_X1 U25895 ( .A(\mem[210][6] ), .B(\mem[211][6] ), .S(n8485), .Z(n6940)
         );
  MUX2_X1 U25896 ( .A(\mem[208][6] ), .B(\mem[209][6] ), .S(n8485), .Z(n6941)
         );
  MUX2_X1 U25897 ( .A(n6941), .B(n6940), .S(n8330), .Z(n6942) );
  MUX2_X1 U25898 ( .A(n6942), .B(n6939), .S(n8240), .Z(n6943) );
  MUX2_X1 U25899 ( .A(n6943), .B(n6936), .S(n8212), .Z(n6944) );
  MUX2_X1 U25900 ( .A(\mem[206][6] ), .B(\mem[207][6] ), .S(n8485), .Z(n6945)
         );
  MUX2_X1 U25901 ( .A(\mem[204][6] ), .B(\mem[205][6] ), .S(n8485), .Z(n6946)
         );
  MUX2_X1 U25902 ( .A(n6946), .B(n6945), .S(n8330), .Z(n6947) );
  MUX2_X1 U25903 ( .A(\mem[202][6] ), .B(\mem[203][6] ), .S(n8485), .Z(n6948)
         );
  MUX2_X1 U25904 ( .A(\mem[200][6] ), .B(\mem[201][6] ), .S(n8485), .Z(n6949)
         );
  MUX2_X1 U25905 ( .A(n6949), .B(n6948), .S(n8330), .Z(n6950) );
  MUX2_X1 U25906 ( .A(n6950), .B(n6947), .S(n8230), .Z(n6951) );
  MUX2_X1 U25907 ( .A(\mem[198][6] ), .B(\mem[199][6] ), .S(n8486), .Z(n6952)
         );
  MUX2_X1 U25908 ( .A(\mem[196][6] ), .B(\mem[197][6] ), .S(n8486), .Z(n6953)
         );
  MUX2_X1 U25909 ( .A(n6953), .B(n6952), .S(n8330), .Z(n6954) );
  MUX2_X1 U25910 ( .A(\mem[194][6] ), .B(\mem[195][6] ), .S(n8486), .Z(n6955)
         );
  MUX2_X1 U25911 ( .A(\mem[192][6] ), .B(\mem[193][6] ), .S(n8486), .Z(n6956)
         );
  MUX2_X1 U25912 ( .A(n6956), .B(n6955), .S(n8330), .Z(n6957) );
  MUX2_X1 U25913 ( .A(n6957), .B(n6954), .S(n8231), .Z(n6958) );
  MUX2_X1 U25914 ( .A(n6958), .B(n6951), .S(n8212), .Z(n6959) );
  MUX2_X1 U25915 ( .A(n6959), .B(n6944), .S(n8191), .Z(n6960) );
  MUX2_X1 U25916 ( .A(n6960), .B(n6929), .S(n8182), .Z(n6961) );
  MUX2_X1 U25917 ( .A(\mem[190][6] ), .B(\mem[191][6] ), .S(n8486), .Z(n6962)
         );
  MUX2_X1 U25918 ( .A(\mem[188][6] ), .B(\mem[189][6] ), .S(n8486), .Z(n6963)
         );
  MUX2_X1 U25919 ( .A(n6963), .B(n6962), .S(n8330), .Z(n6964) );
  MUX2_X1 U25920 ( .A(\mem[186][6] ), .B(\mem[187][6] ), .S(n8486), .Z(n6965)
         );
  MUX2_X1 U25921 ( .A(\mem[184][6] ), .B(\mem[185][6] ), .S(n8486), .Z(n6966)
         );
  MUX2_X1 U25922 ( .A(n6966), .B(n6965), .S(n8330), .Z(n6967) );
  MUX2_X1 U25923 ( .A(n6967), .B(n6964), .S(n8227), .Z(n6968) );
  MUX2_X1 U25924 ( .A(\mem[182][6] ), .B(\mem[183][6] ), .S(n8486), .Z(n6969)
         );
  MUX2_X1 U25925 ( .A(\mem[180][6] ), .B(\mem[181][6] ), .S(n8486), .Z(n6970)
         );
  MUX2_X1 U25926 ( .A(n6970), .B(n6969), .S(n8330), .Z(n6971) );
  MUX2_X1 U25927 ( .A(\mem[178][6] ), .B(\mem[179][6] ), .S(n8486), .Z(n6972)
         );
  MUX2_X1 U25928 ( .A(\mem[176][6] ), .B(\mem[177][6] ), .S(n8486), .Z(n6973)
         );
  MUX2_X1 U25929 ( .A(n6973), .B(n6972), .S(n8330), .Z(n6974) );
  MUX2_X1 U25930 ( .A(n6974), .B(n6971), .S(n8228), .Z(n6975) );
  MUX2_X1 U25931 ( .A(n6975), .B(n6968), .S(n8212), .Z(n6976) );
  MUX2_X1 U25932 ( .A(\mem[174][6] ), .B(\mem[175][6] ), .S(n8487), .Z(n6977)
         );
  MUX2_X1 U25933 ( .A(\mem[172][6] ), .B(\mem[173][6] ), .S(n8487), .Z(n6978)
         );
  MUX2_X1 U25934 ( .A(n6978), .B(n6977), .S(n8331), .Z(n6979) );
  MUX2_X1 U25935 ( .A(\mem[170][6] ), .B(\mem[171][6] ), .S(n8487), .Z(n6980)
         );
  MUX2_X1 U25936 ( .A(\mem[168][6] ), .B(\mem[169][6] ), .S(n8487), .Z(n6981)
         );
  MUX2_X1 U25937 ( .A(n6981), .B(n6980), .S(n8331), .Z(n6982) );
  MUX2_X1 U25938 ( .A(n6982), .B(n6979), .S(n8229), .Z(n6983) );
  MUX2_X1 U25939 ( .A(\mem[166][6] ), .B(\mem[167][6] ), .S(n8487), .Z(n6984)
         );
  MUX2_X1 U25940 ( .A(\mem[164][6] ), .B(\mem[165][6] ), .S(n8487), .Z(n6985)
         );
  MUX2_X1 U25941 ( .A(n6985), .B(n6984), .S(n8331), .Z(n6986) );
  MUX2_X1 U25942 ( .A(\mem[162][6] ), .B(\mem[163][6] ), .S(n8487), .Z(n6987)
         );
  MUX2_X1 U25943 ( .A(\mem[160][6] ), .B(\mem[161][6] ), .S(n8487), .Z(n6988)
         );
  MUX2_X1 U25944 ( .A(n6988), .B(n6987), .S(n8331), .Z(n6989) );
  MUX2_X1 U25945 ( .A(n6989), .B(n6986), .S(n8226), .Z(n6990) );
  MUX2_X1 U25946 ( .A(n6990), .B(n6983), .S(n8212), .Z(n6991) );
  MUX2_X1 U25947 ( .A(n6991), .B(n6976), .S(n8191), .Z(n6992) );
  MUX2_X1 U25948 ( .A(\mem[158][6] ), .B(\mem[159][6] ), .S(n8487), .Z(n6993)
         );
  MUX2_X1 U25949 ( .A(\mem[156][6] ), .B(\mem[157][6] ), .S(n8487), .Z(n6994)
         );
  MUX2_X1 U25950 ( .A(n6994), .B(n6993), .S(n8331), .Z(n6995) );
  MUX2_X1 U25951 ( .A(\mem[154][6] ), .B(\mem[155][6] ), .S(n8487), .Z(n6996)
         );
  MUX2_X1 U25952 ( .A(\mem[152][6] ), .B(\mem[153][6] ), .S(n8487), .Z(n6997)
         );
  MUX2_X1 U25953 ( .A(n6997), .B(n6996), .S(n8331), .Z(n6998) );
  MUX2_X1 U25954 ( .A(n6998), .B(n6995), .S(n8247), .Z(n6999) );
  MUX2_X1 U25955 ( .A(\mem[150][6] ), .B(\mem[151][6] ), .S(n8488), .Z(n7000)
         );
  MUX2_X1 U25956 ( .A(\mem[148][6] ), .B(\mem[149][6] ), .S(n8488), .Z(n7001)
         );
  MUX2_X1 U25957 ( .A(n7001), .B(n7000), .S(n8331), .Z(n7002) );
  MUX2_X1 U25958 ( .A(\mem[146][6] ), .B(\mem[147][6] ), .S(n8488), .Z(n7003)
         );
  MUX2_X1 U25959 ( .A(\mem[144][6] ), .B(\mem[145][6] ), .S(n8488), .Z(n7004)
         );
  MUX2_X1 U25960 ( .A(n7004), .B(n7003), .S(n8331), .Z(n7005) );
  MUX2_X1 U25961 ( .A(n7005), .B(n7002), .S(n8248), .Z(n7006) );
  MUX2_X1 U25962 ( .A(n7006), .B(n6999), .S(n8212), .Z(n7007) );
  MUX2_X1 U25963 ( .A(\mem[142][6] ), .B(\mem[143][6] ), .S(n8488), .Z(n7008)
         );
  MUX2_X1 U25964 ( .A(\mem[140][6] ), .B(\mem[141][6] ), .S(n8488), .Z(n7009)
         );
  MUX2_X1 U25965 ( .A(n7009), .B(n7008), .S(n8331), .Z(n7010) );
  MUX2_X1 U25966 ( .A(\mem[138][6] ), .B(\mem[139][6] ), .S(n8488), .Z(n7011)
         );
  MUX2_X1 U25967 ( .A(\mem[136][6] ), .B(\mem[137][6] ), .S(n8488), .Z(n7012)
         );
  MUX2_X1 U25968 ( .A(n7012), .B(n7011), .S(n8331), .Z(n7013) );
  MUX2_X1 U25969 ( .A(n7013), .B(n7010), .S(n8249), .Z(n7014) );
  MUX2_X1 U25970 ( .A(\mem[134][6] ), .B(\mem[135][6] ), .S(n8488), .Z(n7015)
         );
  MUX2_X1 U25971 ( .A(\mem[132][6] ), .B(\mem[133][6] ), .S(n8488), .Z(n7016)
         );
  MUX2_X1 U25972 ( .A(n7016), .B(n7015), .S(n8331), .Z(n7017) );
  MUX2_X1 U25973 ( .A(\mem[130][6] ), .B(\mem[131][6] ), .S(n8488), .Z(n7018)
         );
  MUX2_X1 U25974 ( .A(\mem[128][6] ), .B(\mem[129][6] ), .S(n8488), .Z(n7019)
         );
  MUX2_X1 U25975 ( .A(n7019), .B(n7018), .S(n8331), .Z(n7020) );
  MUX2_X1 U25976 ( .A(n7020), .B(n7017), .S(n8244), .Z(n7021) );
  MUX2_X1 U25977 ( .A(n7021), .B(n7014), .S(n8212), .Z(n7022) );
  MUX2_X1 U25978 ( .A(n7022), .B(n7007), .S(n8191), .Z(n7023) );
  MUX2_X1 U25979 ( .A(n7023), .B(n6992), .S(n8183), .Z(n7024) );
  MUX2_X1 U25980 ( .A(n7024), .B(n6961), .S(n8180), .Z(n7025) );
  MUX2_X1 U25981 ( .A(\mem[126][6] ), .B(\mem[127][6] ), .S(n8489), .Z(n7026)
         );
  MUX2_X1 U25982 ( .A(\mem[124][6] ), .B(\mem[125][6] ), .S(n8489), .Z(n7027)
         );
  MUX2_X1 U25983 ( .A(n7027), .B(n7026), .S(n8332), .Z(n7028) );
  MUX2_X1 U25984 ( .A(\mem[122][6] ), .B(\mem[123][6] ), .S(n8489), .Z(n7029)
         );
  MUX2_X1 U25985 ( .A(\mem[120][6] ), .B(\mem[121][6] ), .S(n8489), .Z(n7030)
         );
  MUX2_X1 U25986 ( .A(n7030), .B(n7029), .S(n8332), .Z(n7031) );
  MUX2_X1 U25987 ( .A(n7031), .B(n7028), .S(n8245), .Z(n7032) );
  MUX2_X1 U25988 ( .A(\mem[118][6] ), .B(\mem[119][6] ), .S(n8489), .Z(n7033)
         );
  MUX2_X1 U25989 ( .A(\mem[116][6] ), .B(\mem[117][6] ), .S(n8489), .Z(n7034)
         );
  MUX2_X1 U25990 ( .A(n7034), .B(n7033), .S(n8332), .Z(n7035) );
  MUX2_X1 U25991 ( .A(\mem[114][6] ), .B(\mem[115][6] ), .S(n8489), .Z(n7036)
         );
  MUX2_X1 U25992 ( .A(\mem[112][6] ), .B(\mem[113][6] ), .S(n8489), .Z(n7037)
         );
  MUX2_X1 U25993 ( .A(n7037), .B(n7036), .S(n8332), .Z(n7038) );
  MUX2_X1 U25994 ( .A(n7038), .B(n7035), .S(n8246), .Z(n7039) );
  MUX2_X1 U25995 ( .A(n7039), .B(n7032), .S(n8213), .Z(n7040) );
  MUX2_X1 U25996 ( .A(\mem[110][6] ), .B(\mem[111][6] ), .S(n8489), .Z(n7041)
         );
  MUX2_X1 U25997 ( .A(\mem[108][6] ), .B(\mem[109][6] ), .S(n8489), .Z(n7042)
         );
  MUX2_X1 U25998 ( .A(n7042), .B(n7041), .S(n8332), .Z(n7043) );
  MUX2_X1 U25999 ( .A(\mem[106][6] ), .B(\mem[107][6] ), .S(n8489), .Z(n7044)
         );
  MUX2_X1 U26000 ( .A(\mem[104][6] ), .B(\mem[105][6] ), .S(n8489), .Z(n7045)
         );
  MUX2_X1 U26001 ( .A(n7045), .B(n7044), .S(n8332), .Z(n7046) );
  MUX2_X1 U26002 ( .A(n7046), .B(n7043), .S(n8253), .Z(n7047) );
  MUX2_X1 U26003 ( .A(\mem[102][6] ), .B(\mem[103][6] ), .S(n8490), .Z(n7048)
         );
  MUX2_X1 U26004 ( .A(\mem[100][6] ), .B(\mem[101][6] ), .S(n8490), .Z(n7049)
         );
  MUX2_X1 U26005 ( .A(n7049), .B(n7048), .S(n8332), .Z(n7050) );
  MUX2_X1 U26006 ( .A(\mem[98][6] ), .B(\mem[99][6] ), .S(n8490), .Z(n7051) );
  MUX2_X1 U26007 ( .A(\mem[96][6] ), .B(\mem[97][6] ), .S(n8490), .Z(n7052) );
  MUX2_X1 U26008 ( .A(n7052), .B(n7051), .S(n8332), .Z(n7053) );
  MUX2_X1 U26009 ( .A(n7053), .B(n7050), .S(n8254), .Z(n7054) );
  MUX2_X1 U26010 ( .A(n7054), .B(n7047), .S(n8213), .Z(n7055) );
  MUX2_X1 U26011 ( .A(n7055), .B(n7040), .S(n8192), .Z(n7056) );
  MUX2_X1 U26012 ( .A(\mem[94][6] ), .B(\mem[95][6] ), .S(n8490), .Z(n7057) );
  MUX2_X1 U26013 ( .A(\mem[92][6] ), .B(\mem[93][6] ), .S(n8490), .Z(n7058) );
  MUX2_X1 U26014 ( .A(n7058), .B(n7057), .S(n8332), .Z(n7059) );
  MUX2_X1 U26015 ( .A(\mem[90][6] ), .B(\mem[91][6] ), .S(n8490), .Z(n7060) );
  MUX2_X1 U26016 ( .A(\mem[88][6] ), .B(\mem[89][6] ), .S(n8490), .Z(n7061) );
  MUX2_X1 U26017 ( .A(n7061), .B(n7060), .S(n8332), .Z(n7062) );
  MUX2_X1 U26018 ( .A(n7062), .B(n7059), .S(n8255), .Z(n7063) );
  MUX2_X1 U26019 ( .A(\mem[86][6] ), .B(\mem[87][6] ), .S(n8490), .Z(n7064) );
  MUX2_X1 U26020 ( .A(\mem[84][6] ), .B(\mem[85][6] ), .S(n8490), .Z(n7065) );
  MUX2_X1 U26021 ( .A(n7065), .B(n7064), .S(n8332), .Z(n7066) );
  MUX2_X1 U26022 ( .A(\mem[82][6] ), .B(\mem[83][6] ), .S(n8490), .Z(n7067) );
  MUX2_X1 U26023 ( .A(\mem[80][6] ), .B(\mem[81][6] ), .S(n8490), .Z(n7068) );
  MUX2_X1 U26024 ( .A(n7068), .B(n7067), .S(n8332), .Z(n7069) );
  MUX2_X1 U26025 ( .A(n7069), .B(n7066), .S(n8250), .Z(n7070) );
  MUX2_X1 U26026 ( .A(n7070), .B(n7063), .S(n8213), .Z(n7071) );
  MUX2_X1 U26027 ( .A(\mem[78][6] ), .B(\mem[79][6] ), .S(n8491), .Z(n7072) );
  MUX2_X1 U26028 ( .A(\mem[76][6] ), .B(\mem[77][6] ), .S(n8491), .Z(n7073) );
  MUX2_X1 U26029 ( .A(n7073), .B(n7072), .S(n8333), .Z(n7074) );
  MUX2_X1 U26030 ( .A(\mem[74][6] ), .B(\mem[75][6] ), .S(n8491), .Z(n7075) );
  MUX2_X1 U26031 ( .A(\mem[72][6] ), .B(\mem[73][6] ), .S(n8491), .Z(n7076) );
  MUX2_X1 U26032 ( .A(n7076), .B(n7075), .S(n8333), .Z(n7077) );
  MUX2_X1 U26033 ( .A(n7077), .B(n7074), .S(n8251), .Z(n7078) );
  MUX2_X1 U26034 ( .A(\mem[70][6] ), .B(\mem[71][6] ), .S(n8491), .Z(n7079) );
  MUX2_X1 U26035 ( .A(\mem[68][6] ), .B(\mem[69][6] ), .S(n8491), .Z(n7080) );
  MUX2_X1 U26036 ( .A(n7080), .B(n7079), .S(n8333), .Z(n7081) );
  MUX2_X1 U26037 ( .A(\mem[66][6] ), .B(\mem[67][6] ), .S(n8491), .Z(n7082) );
  MUX2_X1 U26038 ( .A(\mem[64][6] ), .B(\mem[65][6] ), .S(n8491), .Z(n7083) );
  MUX2_X1 U26039 ( .A(n7083), .B(n7082), .S(n8333), .Z(n7084) );
  MUX2_X1 U26040 ( .A(n7084), .B(n7081), .S(n8252), .Z(n7085) );
  MUX2_X1 U26041 ( .A(n7085), .B(n7078), .S(n8213), .Z(n7086) );
  MUX2_X1 U26042 ( .A(n7086), .B(n7071), .S(n8192), .Z(n7087) );
  MUX2_X1 U26043 ( .A(n7087), .B(n7056), .S(n8184), .Z(n7088) );
  MUX2_X1 U26044 ( .A(\mem[62][6] ), .B(\mem[63][6] ), .S(n8491), .Z(n7089) );
  MUX2_X1 U26045 ( .A(\mem[60][6] ), .B(\mem[61][6] ), .S(n8491), .Z(n7090) );
  MUX2_X1 U26046 ( .A(n7090), .B(n7089), .S(n8333), .Z(n7091) );
  MUX2_X1 U26047 ( .A(\mem[58][6] ), .B(\mem[59][6] ), .S(n8491), .Z(n7092) );
  MUX2_X1 U26048 ( .A(\mem[56][6] ), .B(\mem[57][6] ), .S(n8491), .Z(n7093) );
  MUX2_X1 U26049 ( .A(n7093), .B(n7092), .S(n8333), .Z(n7094) );
  MUX2_X1 U26050 ( .A(n7094), .B(n7091), .S(n8259), .Z(n7095) );
  MUX2_X1 U26051 ( .A(\mem[54][6] ), .B(\mem[55][6] ), .S(n8492), .Z(n7096) );
  MUX2_X1 U26052 ( .A(\mem[52][6] ), .B(\mem[53][6] ), .S(n8492), .Z(n7097) );
  MUX2_X1 U26053 ( .A(n7097), .B(n7096), .S(n8333), .Z(n7098) );
  MUX2_X1 U26054 ( .A(\mem[50][6] ), .B(\mem[51][6] ), .S(n8492), .Z(n7099) );
  MUX2_X1 U26055 ( .A(\mem[48][6] ), .B(\mem[49][6] ), .S(n8492), .Z(n7100) );
  MUX2_X1 U26056 ( .A(n7100), .B(n7099), .S(n8333), .Z(n7101) );
  MUX2_X1 U26057 ( .A(n7101), .B(n7098), .S(n8260), .Z(n7102) );
  MUX2_X1 U26058 ( .A(n7102), .B(n7095), .S(n8213), .Z(n7103) );
  MUX2_X1 U26059 ( .A(\mem[46][6] ), .B(\mem[47][6] ), .S(n8492), .Z(n7104) );
  MUX2_X1 U26060 ( .A(\mem[44][6] ), .B(\mem[45][6] ), .S(n8492), .Z(n7105) );
  MUX2_X1 U26061 ( .A(n7105), .B(n7104), .S(n8333), .Z(n7106) );
  MUX2_X1 U26062 ( .A(\mem[42][6] ), .B(\mem[43][6] ), .S(n8492), .Z(n7107) );
  MUX2_X1 U26063 ( .A(\mem[40][6] ), .B(\mem[41][6] ), .S(n8492), .Z(n7108) );
  MUX2_X1 U26064 ( .A(n7108), .B(n7107), .S(n8333), .Z(n7109) );
  MUX2_X1 U26065 ( .A(n7109), .B(n7106), .S(n8261), .Z(n7110) );
  MUX2_X1 U26066 ( .A(\mem[38][6] ), .B(\mem[39][6] ), .S(n8492), .Z(n7111) );
  MUX2_X1 U26067 ( .A(\mem[36][6] ), .B(\mem[37][6] ), .S(n8492), .Z(n7112) );
  MUX2_X1 U26068 ( .A(n7112), .B(n7111), .S(n8333), .Z(n7113) );
  MUX2_X1 U26069 ( .A(\mem[34][6] ), .B(\mem[35][6] ), .S(n8492), .Z(n7114) );
  MUX2_X1 U26070 ( .A(\mem[32][6] ), .B(\mem[33][6] ), .S(n8492), .Z(n7115) );
  MUX2_X1 U26071 ( .A(n7115), .B(n7114), .S(n8333), .Z(n7116) );
  MUX2_X1 U26072 ( .A(n7116), .B(n7113), .S(n8256), .Z(n7117) );
  MUX2_X1 U26073 ( .A(n7117), .B(n7110), .S(n8213), .Z(n7118) );
  MUX2_X1 U26074 ( .A(n7118), .B(n7103), .S(n8192), .Z(n7119) );
  MUX2_X1 U26075 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n8493), .Z(n7120) );
  MUX2_X1 U26076 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n8493), .Z(n7121) );
  MUX2_X1 U26077 ( .A(n7121), .B(n7120), .S(n8334), .Z(n7122) );
  MUX2_X1 U26078 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n8493), .Z(n7123) );
  MUX2_X1 U26079 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n8493), .Z(n7124) );
  MUX2_X1 U26080 ( .A(n7124), .B(n7123), .S(n8334), .Z(n7125) );
  MUX2_X1 U26081 ( .A(n7125), .B(n7122), .S(n8255), .Z(n7126) );
  MUX2_X1 U26082 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n8493), .Z(n7127) );
  MUX2_X1 U26083 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n8493), .Z(n7128) );
  MUX2_X1 U26084 ( .A(n7128), .B(n7127), .S(n8334), .Z(n7129) );
  MUX2_X1 U26085 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n8493), .Z(n7130) );
  MUX2_X1 U26086 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n8493), .Z(n7131) );
  MUX2_X1 U26087 ( .A(n7131), .B(n7130), .S(n8334), .Z(n7132) );
  MUX2_X1 U26088 ( .A(n7132), .B(n7129), .S(n8250), .Z(n7133) );
  MUX2_X1 U26089 ( .A(n7133), .B(n7126), .S(n8213), .Z(n7134) );
  MUX2_X1 U26090 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n8493), .Z(n7135) );
  MUX2_X1 U26091 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n8493), .Z(n7136) );
  MUX2_X1 U26092 ( .A(n7136), .B(n7135), .S(n8334), .Z(n7137) );
  MUX2_X1 U26093 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n8493), .Z(n7138) );
  MUX2_X1 U26094 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n8493), .Z(n7139) );
  MUX2_X1 U26095 ( .A(n7139), .B(n7138), .S(n8334), .Z(n7140) );
  MUX2_X1 U26096 ( .A(n7140), .B(n7137), .S(n8251), .Z(n7141) );
  MUX2_X1 U26097 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n8494), .Z(n7142) );
  MUX2_X1 U26098 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n8494), .Z(n7143) );
  MUX2_X1 U26099 ( .A(n7143), .B(n7142), .S(n8334), .Z(n7144) );
  MUX2_X1 U26100 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n8494), .Z(n7145) );
  MUX2_X1 U26101 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n8494), .Z(n7146) );
  MUX2_X1 U26102 ( .A(n7146), .B(n7145), .S(n8334), .Z(n7147) );
  MUX2_X1 U26103 ( .A(n7147), .B(n7144), .S(n8252), .Z(n7148) );
  MUX2_X1 U26104 ( .A(n7148), .B(n7141), .S(n8213), .Z(n7149) );
  MUX2_X1 U26105 ( .A(n7149), .B(n7134), .S(n8192), .Z(n7150) );
  MUX2_X1 U26106 ( .A(n7150), .B(n7119), .S(n8181), .Z(n7151) );
  MUX2_X1 U26107 ( .A(n7151), .B(n7088), .S(n8180), .Z(n7152) );
  MUX2_X1 U26108 ( .A(n7152), .B(n7025), .S(n8177), .Z(n7153) );
  MUX2_X1 U26109 ( .A(n7153), .B(n6898), .S(N26), .Z(n7154) );
  MUX2_X1 U26110 ( .A(n7154), .B(n6643), .S(N27), .Z(N29) );
  MUX2_X1 U26111 ( .A(\mem[1022][7] ), .B(\mem[1023][7] ), .S(n8494), .Z(n7155) );
  MUX2_X1 U26112 ( .A(\mem[1020][7] ), .B(\mem[1021][7] ), .S(n8494), .Z(n7156) );
  MUX2_X1 U26113 ( .A(n7156), .B(n7155), .S(n8334), .Z(n7157) );
  MUX2_X1 U26114 ( .A(\mem[1018][7] ), .B(\mem[1019][7] ), .S(n8494), .Z(n7158) );
  MUX2_X1 U26115 ( .A(\mem[1016][7] ), .B(\mem[1017][7] ), .S(n8494), .Z(n7159) );
  MUX2_X1 U26116 ( .A(n7159), .B(n7158), .S(n8334), .Z(n7160) );
  MUX2_X1 U26117 ( .A(n7160), .B(n7157), .S(n8259), .Z(n7161) );
  MUX2_X1 U26118 ( .A(\mem[1014][7] ), .B(\mem[1015][7] ), .S(n8494), .Z(n7162) );
  MUX2_X1 U26119 ( .A(\mem[1012][7] ), .B(\mem[1013][7] ), .S(n8494), .Z(n7163) );
  MUX2_X1 U26120 ( .A(n7163), .B(n7162), .S(n8334), .Z(n7164) );
  MUX2_X1 U26121 ( .A(\mem[1010][7] ), .B(\mem[1011][7] ), .S(n8494), .Z(n7165) );
  MUX2_X1 U26122 ( .A(\mem[1008][7] ), .B(\mem[1009][7] ), .S(n8494), .Z(n7166) );
  MUX2_X1 U26123 ( .A(n7166), .B(n7165), .S(n8334), .Z(n7167) );
  MUX2_X1 U26124 ( .A(n7167), .B(n7164), .S(n8260), .Z(n7168) );
  MUX2_X1 U26125 ( .A(n7168), .B(n7161), .S(n8213), .Z(n7169) );
  MUX2_X1 U26126 ( .A(\mem[1006][7] ), .B(\mem[1007][7] ), .S(n8495), .Z(n7170) );
  MUX2_X1 U26127 ( .A(\mem[1004][7] ), .B(\mem[1005][7] ), .S(n8495), .Z(n7171) );
  MUX2_X1 U26128 ( .A(n7171), .B(n7170), .S(n8335), .Z(n7172) );
  MUX2_X1 U26129 ( .A(\mem[1002][7] ), .B(\mem[1003][7] ), .S(n8495), .Z(n7173) );
  MUX2_X1 U26130 ( .A(\mem[1000][7] ), .B(\mem[1001][7] ), .S(n8495), .Z(n7174) );
  MUX2_X1 U26131 ( .A(n7174), .B(n7173), .S(n8335), .Z(n7175) );
  MUX2_X1 U26132 ( .A(n7175), .B(n7172), .S(n8261), .Z(n7176) );
  MUX2_X1 U26133 ( .A(\mem[998][7] ), .B(\mem[999][7] ), .S(n8495), .Z(n7177)
         );
  MUX2_X1 U26134 ( .A(\mem[996][7] ), .B(\mem[997][7] ), .S(n8495), .Z(n7178)
         );
  MUX2_X1 U26135 ( .A(n7178), .B(n7177), .S(n8335), .Z(n7179) );
  MUX2_X1 U26136 ( .A(\mem[994][7] ), .B(\mem[995][7] ), .S(n8495), .Z(n7180)
         );
  MUX2_X1 U26137 ( .A(\mem[992][7] ), .B(\mem[993][7] ), .S(n8495), .Z(n7181)
         );
  MUX2_X1 U26138 ( .A(n7181), .B(n7180), .S(n8335), .Z(n7182) );
  MUX2_X1 U26139 ( .A(n7182), .B(n7179), .S(n8256), .Z(n7183) );
  MUX2_X1 U26140 ( .A(n7183), .B(n7176), .S(n8213), .Z(n7184) );
  MUX2_X1 U26141 ( .A(n7184), .B(n7169), .S(n8192), .Z(n7185) );
  MUX2_X1 U26142 ( .A(\mem[990][7] ), .B(\mem[991][7] ), .S(n8495), .Z(n7186)
         );
  MUX2_X1 U26143 ( .A(\mem[988][7] ), .B(\mem[989][7] ), .S(n8495), .Z(n7187)
         );
  MUX2_X1 U26144 ( .A(n7187), .B(n7186), .S(n8335), .Z(n7188) );
  MUX2_X1 U26145 ( .A(\mem[986][7] ), .B(\mem[987][7] ), .S(n8495), .Z(n7189)
         );
  MUX2_X1 U26146 ( .A(\mem[984][7] ), .B(\mem[985][7] ), .S(n8495), .Z(n7190)
         );
  MUX2_X1 U26147 ( .A(n7190), .B(n7189), .S(n8335), .Z(n7191) );
  MUX2_X1 U26148 ( .A(n7191), .B(n7188), .S(n8257), .Z(n7192) );
  MUX2_X1 U26149 ( .A(\mem[982][7] ), .B(\mem[983][7] ), .S(n8496), .Z(n7193)
         );
  MUX2_X1 U26150 ( .A(\mem[980][7] ), .B(\mem[981][7] ), .S(n8496), .Z(n7194)
         );
  MUX2_X1 U26151 ( .A(n7194), .B(n7193), .S(n8335), .Z(n7195) );
  MUX2_X1 U26152 ( .A(\mem[978][7] ), .B(\mem[979][7] ), .S(n8496), .Z(n7196)
         );
  MUX2_X1 U26153 ( .A(\mem[976][7] ), .B(\mem[977][7] ), .S(n8496), .Z(n7197)
         );
  MUX2_X1 U26154 ( .A(n7197), .B(n7196), .S(n8335), .Z(n7198) );
  MUX2_X1 U26155 ( .A(n7198), .B(n7195), .S(n8258), .Z(n7199) );
  MUX2_X1 U26156 ( .A(n7199), .B(n7192), .S(n8213), .Z(n7200) );
  MUX2_X1 U26157 ( .A(\mem[974][7] ), .B(\mem[975][7] ), .S(n8496), .Z(n7201)
         );
  MUX2_X1 U26158 ( .A(\mem[972][7] ), .B(\mem[973][7] ), .S(n8496), .Z(n7202)
         );
  MUX2_X1 U26159 ( .A(n7202), .B(n7201), .S(n8335), .Z(n7203) );
  MUX2_X1 U26160 ( .A(\mem[970][7] ), .B(\mem[971][7] ), .S(n8496), .Z(n7204)
         );
  MUX2_X1 U26161 ( .A(\mem[968][7] ), .B(\mem[969][7] ), .S(n8496), .Z(n7205)
         );
  MUX2_X1 U26162 ( .A(n7205), .B(n7204), .S(n8335), .Z(n7206) );
  MUX2_X1 U26163 ( .A(n7206), .B(n7203), .S(n8223), .Z(n7207) );
  MUX2_X1 U26164 ( .A(\mem[966][7] ), .B(\mem[967][7] ), .S(n8496), .Z(n7208)
         );
  MUX2_X1 U26165 ( .A(\mem[964][7] ), .B(\mem[965][7] ), .S(n8496), .Z(n7209)
         );
  MUX2_X1 U26166 ( .A(n7209), .B(n7208), .S(n8335), .Z(n7210) );
  MUX2_X1 U26167 ( .A(\mem[962][7] ), .B(\mem[963][7] ), .S(n8496), .Z(n7211)
         );
  MUX2_X1 U26168 ( .A(\mem[960][7] ), .B(\mem[961][7] ), .S(n8496), .Z(n7212)
         );
  MUX2_X1 U26169 ( .A(n7212), .B(n7211), .S(n8335), .Z(n7213) );
  MUX2_X1 U26170 ( .A(n7213), .B(n7210), .S(n8256), .Z(n7214) );
  MUX2_X1 U26171 ( .A(n7214), .B(n7207), .S(n8213), .Z(n7215) );
  MUX2_X1 U26172 ( .A(n7215), .B(n7200), .S(n8192), .Z(n7216) );
  MUX2_X1 U26173 ( .A(n7216), .B(n7185), .S(n8185), .Z(n7217) );
  MUX2_X1 U26174 ( .A(\mem[958][7] ), .B(\mem[959][7] ), .S(n8497), .Z(n7218)
         );
  MUX2_X1 U26175 ( .A(\mem[956][7] ), .B(\mem[957][7] ), .S(n8497), .Z(n7219)
         );
  MUX2_X1 U26176 ( .A(n7219), .B(n7218), .S(n8336), .Z(n7220) );
  MUX2_X1 U26177 ( .A(\mem[954][7] ), .B(\mem[955][7] ), .S(n8497), .Z(n7221)
         );
  MUX2_X1 U26178 ( .A(\mem[952][7] ), .B(\mem[953][7] ), .S(n8497), .Z(n7222)
         );
  MUX2_X1 U26179 ( .A(n7222), .B(n7221), .S(n8336), .Z(n7223) );
  MUX2_X1 U26180 ( .A(n7223), .B(n7220), .S(n8222), .Z(n7224) );
  MUX2_X1 U26181 ( .A(\mem[950][7] ), .B(\mem[951][7] ), .S(n8497), .Z(n7225)
         );
  MUX2_X1 U26182 ( .A(\mem[948][7] ), .B(\mem[949][7] ), .S(n8497), .Z(n7226)
         );
  MUX2_X1 U26183 ( .A(n7226), .B(n7225), .S(n8336), .Z(n7227) );
  MUX2_X1 U26184 ( .A(\mem[946][7] ), .B(\mem[947][7] ), .S(n8497), .Z(n7228)
         );
  MUX2_X1 U26185 ( .A(\mem[944][7] ), .B(\mem[945][7] ), .S(n8497), .Z(n7229)
         );
  MUX2_X1 U26186 ( .A(n7229), .B(n7228), .S(n8336), .Z(n7230) );
  MUX2_X1 U26187 ( .A(n7230), .B(n7227), .S(n8221), .Z(n7231) );
  MUX2_X1 U26188 ( .A(n7231), .B(n7224), .S(n8214), .Z(n7232) );
  MUX2_X1 U26189 ( .A(\mem[942][7] ), .B(\mem[943][7] ), .S(n8497), .Z(n7233)
         );
  MUX2_X1 U26190 ( .A(\mem[940][7] ), .B(\mem[941][7] ), .S(n8497), .Z(n7234)
         );
  MUX2_X1 U26191 ( .A(n7234), .B(n7233), .S(n8336), .Z(n7235) );
  MUX2_X1 U26192 ( .A(\mem[938][7] ), .B(\mem[939][7] ), .S(n8497), .Z(n7236)
         );
  MUX2_X1 U26193 ( .A(\mem[936][7] ), .B(\mem[937][7] ), .S(n8497), .Z(n7237)
         );
  MUX2_X1 U26194 ( .A(n7237), .B(n7236), .S(n8336), .Z(n7238) );
  MUX2_X1 U26195 ( .A(n7238), .B(n7235), .S(n8220), .Z(n7239) );
  MUX2_X1 U26196 ( .A(\mem[934][7] ), .B(\mem[935][7] ), .S(n8498), .Z(n7240)
         );
  MUX2_X1 U26197 ( .A(\mem[932][7] ), .B(\mem[933][7] ), .S(n8498), .Z(n7241)
         );
  MUX2_X1 U26198 ( .A(n7241), .B(n7240), .S(n8336), .Z(n7242) );
  MUX2_X1 U26199 ( .A(\mem[930][7] ), .B(\mem[931][7] ), .S(n8498), .Z(n7243)
         );
  MUX2_X1 U26200 ( .A(\mem[928][7] ), .B(\mem[929][7] ), .S(n8498), .Z(n7244)
         );
  MUX2_X1 U26201 ( .A(n7244), .B(n7243), .S(n8336), .Z(n7245) );
  MUX2_X1 U26202 ( .A(n7245), .B(n7242), .S(n8229), .Z(n7246) );
  MUX2_X1 U26203 ( .A(n7246), .B(n7239), .S(n8214), .Z(n7247) );
  MUX2_X1 U26204 ( .A(n7247), .B(n7232), .S(n8192), .Z(n7248) );
  MUX2_X1 U26205 ( .A(\mem[926][7] ), .B(\mem[927][7] ), .S(n8498), .Z(n7249)
         );
  MUX2_X1 U26206 ( .A(\mem[924][7] ), .B(\mem[925][7] ), .S(n8498), .Z(n7250)
         );
  MUX2_X1 U26207 ( .A(n7250), .B(n7249), .S(n8336), .Z(n7251) );
  MUX2_X1 U26208 ( .A(\mem[922][7] ), .B(\mem[923][7] ), .S(n8498), .Z(n7252)
         );
  MUX2_X1 U26209 ( .A(\mem[920][7] ), .B(\mem[921][7] ), .S(n8498), .Z(n7253)
         );
  MUX2_X1 U26210 ( .A(n7253), .B(n7252), .S(n8336), .Z(n7254) );
  MUX2_X1 U26211 ( .A(n7254), .B(n7251), .S(n8227), .Z(n7255) );
  MUX2_X1 U26212 ( .A(\mem[918][7] ), .B(\mem[919][7] ), .S(n8498), .Z(n7256)
         );
  MUX2_X1 U26213 ( .A(\mem[916][7] ), .B(\mem[917][7] ), .S(n8498), .Z(n7257)
         );
  MUX2_X1 U26214 ( .A(n7257), .B(n7256), .S(n8336), .Z(n7258) );
  MUX2_X1 U26215 ( .A(\mem[914][7] ), .B(\mem[915][7] ), .S(n8498), .Z(n7259)
         );
  MUX2_X1 U26216 ( .A(\mem[912][7] ), .B(\mem[913][7] ), .S(n8498), .Z(n7260)
         );
  MUX2_X1 U26217 ( .A(n7260), .B(n7259), .S(n8336), .Z(n7261) );
  MUX2_X1 U26218 ( .A(n7261), .B(n7258), .S(n8265), .Z(n7262) );
  MUX2_X1 U26219 ( .A(n7262), .B(n7255), .S(n8214), .Z(n7263) );
  MUX2_X1 U26220 ( .A(\mem[910][7] ), .B(\mem[911][7] ), .S(n8499), .Z(n7264)
         );
  MUX2_X1 U26221 ( .A(\mem[908][7] ), .B(\mem[909][7] ), .S(n8499), .Z(n7265)
         );
  MUX2_X1 U26222 ( .A(n7265), .B(n7264), .S(n8337), .Z(n7266) );
  MUX2_X1 U26223 ( .A(\mem[906][7] ), .B(\mem[907][7] ), .S(n8499), .Z(n7267)
         );
  MUX2_X1 U26224 ( .A(\mem[904][7] ), .B(\mem[905][7] ), .S(n8499), .Z(n7268)
         );
  MUX2_X1 U26225 ( .A(n7268), .B(n7267), .S(n8337), .Z(n7269) );
  MUX2_X1 U26226 ( .A(n7269), .B(n7266), .S(n8256), .Z(n7270) );
  MUX2_X1 U26227 ( .A(\mem[902][7] ), .B(\mem[903][7] ), .S(n8499), .Z(n7271)
         );
  MUX2_X1 U26228 ( .A(\mem[900][7] ), .B(\mem[901][7] ), .S(n8499), .Z(n7272)
         );
  MUX2_X1 U26229 ( .A(n7272), .B(n7271), .S(n8337), .Z(n7273) );
  MUX2_X1 U26230 ( .A(\mem[898][7] ), .B(\mem[899][7] ), .S(n8499), .Z(n7274)
         );
  MUX2_X1 U26231 ( .A(\mem[896][7] ), .B(\mem[897][7] ), .S(n8499), .Z(n7275)
         );
  MUX2_X1 U26232 ( .A(n7275), .B(n7274), .S(n8337), .Z(n7276) );
  MUX2_X1 U26233 ( .A(n7276), .B(n7273), .S(n8235), .Z(n7277) );
  MUX2_X1 U26234 ( .A(n7277), .B(n7270), .S(n8214), .Z(n7278) );
  MUX2_X1 U26235 ( .A(n7278), .B(n7263), .S(n8192), .Z(n7279) );
  MUX2_X1 U26236 ( .A(n7279), .B(n7248), .S(N23), .Z(n7280) );
  MUX2_X1 U26237 ( .A(n7280), .B(n7217), .S(n8180), .Z(n7281) );
  MUX2_X1 U26238 ( .A(\mem[894][7] ), .B(\mem[895][7] ), .S(n8499), .Z(n7282)
         );
  MUX2_X1 U26239 ( .A(\mem[892][7] ), .B(\mem[893][7] ), .S(n8499), .Z(n7283)
         );
  MUX2_X1 U26240 ( .A(n7283), .B(n7282), .S(n8337), .Z(n7284) );
  MUX2_X1 U26241 ( .A(\mem[890][7] ), .B(\mem[891][7] ), .S(n8499), .Z(n7285)
         );
  MUX2_X1 U26242 ( .A(\mem[888][7] ), .B(\mem[889][7] ), .S(n8499), .Z(n7286)
         );
  MUX2_X1 U26243 ( .A(n7286), .B(n7285), .S(n8337), .Z(n7287) );
  MUX2_X1 U26244 ( .A(n7287), .B(n7284), .S(n8236), .Z(n7288) );
  MUX2_X1 U26245 ( .A(\mem[886][7] ), .B(\mem[887][7] ), .S(n8500), .Z(n7289)
         );
  MUX2_X1 U26246 ( .A(\mem[884][7] ), .B(\mem[885][7] ), .S(n8500), .Z(n7290)
         );
  MUX2_X1 U26247 ( .A(n7290), .B(n7289), .S(n8337), .Z(n7291) );
  MUX2_X1 U26248 ( .A(\mem[882][7] ), .B(\mem[883][7] ), .S(n8500), .Z(n7292)
         );
  MUX2_X1 U26249 ( .A(\mem[880][7] ), .B(\mem[881][7] ), .S(n8500), .Z(n7293)
         );
  MUX2_X1 U26250 ( .A(n7293), .B(n7292), .S(n8337), .Z(n7294) );
  MUX2_X1 U26251 ( .A(n7294), .B(n7291), .S(n8237), .Z(n7295) );
  MUX2_X1 U26252 ( .A(n7295), .B(n7288), .S(n8214), .Z(n7296) );
  MUX2_X1 U26253 ( .A(\mem[878][7] ), .B(\mem[879][7] ), .S(n8500), .Z(n7297)
         );
  MUX2_X1 U26254 ( .A(\mem[876][7] ), .B(\mem[877][7] ), .S(n8500), .Z(n7298)
         );
  MUX2_X1 U26255 ( .A(n7298), .B(n7297), .S(n8337), .Z(n7299) );
  MUX2_X1 U26256 ( .A(\mem[874][7] ), .B(\mem[875][7] ), .S(n8500), .Z(n7300)
         );
  MUX2_X1 U26257 ( .A(\mem[872][7] ), .B(\mem[873][7] ), .S(n8500), .Z(n7301)
         );
  MUX2_X1 U26258 ( .A(n7301), .B(n7300), .S(n8337), .Z(n7302) );
  MUX2_X1 U26259 ( .A(n7302), .B(n7299), .S(n8232), .Z(n7303) );
  MUX2_X1 U26260 ( .A(\mem[870][7] ), .B(\mem[871][7] ), .S(n8500), .Z(n7304)
         );
  MUX2_X1 U26261 ( .A(\mem[868][7] ), .B(\mem[869][7] ), .S(n8500), .Z(n7305)
         );
  MUX2_X1 U26262 ( .A(n7305), .B(n7304), .S(n8337), .Z(n7306) );
  MUX2_X1 U26263 ( .A(\mem[866][7] ), .B(\mem[867][7] ), .S(n8500), .Z(n7307)
         );
  MUX2_X1 U26264 ( .A(\mem[864][7] ), .B(\mem[865][7] ), .S(n8500), .Z(n7308)
         );
  MUX2_X1 U26265 ( .A(n7308), .B(n7307), .S(n8337), .Z(n7309) );
  MUX2_X1 U26266 ( .A(n7309), .B(n7306), .S(n8233), .Z(n7310) );
  MUX2_X1 U26267 ( .A(n7310), .B(n7303), .S(n8214), .Z(n7311) );
  MUX2_X1 U26268 ( .A(n7311), .B(n7296), .S(n8192), .Z(n7312) );
  MUX2_X1 U26269 ( .A(\mem[862][7] ), .B(\mem[863][7] ), .S(n8501), .Z(n7313)
         );
  MUX2_X1 U26270 ( .A(\mem[860][7] ), .B(\mem[861][7] ), .S(n8501), .Z(n7314)
         );
  MUX2_X1 U26271 ( .A(n7314), .B(n7313), .S(n8338), .Z(n7315) );
  MUX2_X1 U26272 ( .A(\mem[858][7] ), .B(\mem[859][7] ), .S(n8501), .Z(n7316)
         );
  MUX2_X1 U26273 ( .A(\mem[856][7] ), .B(\mem[857][7] ), .S(n8501), .Z(n7317)
         );
  MUX2_X1 U26274 ( .A(n7317), .B(n7316), .S(n8338), .Z(n7318) );
  MUX2_X1 U26275 ( .A(n7318), .B(n7315), .S(n8247), .Z(n7319) );
  MUX2_X1 U26276 ( .A(\mem[854][7] ), .B(\mem[855][7] ), .S(n8501), .Z(n7320)
         );
  MUX2_X1 U26277 ( .A(\mem[852][7] ), .B(\mem[853][7] ), .S(n8501), .Z(n7321)
         );
  MUX2_X1 U26278 ( .A(n7321), .B(n7320), .S(n8338), .Z(n7322) );
  MUX2_X1 U26279 ( .A(\mem[850][7] ), .B(\mem[851][7] ), .S(n8501), .Z(n7323)
         );
  MUX2_X1 U26280 ( .A(\mem[848][7] ), .B(\mem[849][7] ), .S(n8501), .Z(n7324)
         );
  MUX2_X1 U26281 ( .A(n7324), .B(n7323), .S(n8338), .Z(n7325) );
  MUX2_X1 U26282 ( .A(n7325), .B(n7322), .S(n8260), .Z(n7326) );
  MUX2_X1 U26283 ( .A(n7326), .B(n7319), .S(n8214), .Z(n7327) );
  MUX2_X1 U26284 ( .A(\mem[846][7] ), .B(\mem[847][7] ), .S(n8501), .Z(n7328)
         );
  MUX2_X1 U26285 ( .A(\mem[844][7] ), .B(\mem[845][7] ), .S(n8501), .Z(n7329)
         );
  MUX2_X1 U26286 ( .A(n7329), .B(n7328), .S(n8338), .Z(n7330) );
  MUX2_X1 U26287 ( .A(\mem[842][7] ), .B(\mem[843][7] ), .S(n8501), .Z(n7331)
         );
  MUX2_X1 U26288 ( .A(\mem[840][7] ), .B(\mem[841][7] ), .S(n8501), .Z(n7332)
         );
  MUX2_X1 U26289 ( .A(n7332), .B(n7331), .S(n8338), .Z(n7333) );
  MUX2_X1 U26290 ( .A(n7333), .B(n7330), .S(n8259), .Z(n7334) );
  MUX2_X1 U26291 ( .A(\mem[838][7] ), .B(\mem[839][7] ), .S(n8502), .Z(n7335)
         );
  MUX2_X1 U26292 ( .A(\mem[836][7] ), .B(\mem[837][7] ), .S(n8502), .Z(n7336)
         );
  MUX2_X1 U26293 ( .A(n7336), .B(n7335), .S(n8338), .Z(n7337) );
  MUX2_X1 U26294 ( .A(\mem[834][7] ), .B(\mem[835][7] ), .S(n8502), .Z(n7338)
         );
  MUX2_X1 U26295 ( .A(\mem[832][7] ), .B(\mem[833][7] ), .S(n8502), .Z(n7339)
         );
  MUX2_X1 U26296 ( .A(n7339), .B(n7338), .S(n8338), .Z(n7340) );
  MUX2_X1 U26297 ( .A(n7340), .B(n7337), .S(n8221), .Z(n7341) );
  MUX2_X1 U26298 ( .A(n7341), .B(n7334), .S(n8214), .Z(n7342) );
  MUX2_X1 U26299 ( .A(n7342), .B(n7327), .S(n8192), .Z(n7343) );
  MUX2_X1 U26300 ( .A(n7343), .B(n7312), .S(N23), .Z(n7344) );
  MUX2_X1 U26301 ( .A(\mem[830][7] ), .B(\mem[831][7] ), .S(n8502), .Z(n7345)
         );
  MUX2_X1 U26302 ( .A(\mem[828][7] ), .B(\mem[829][7] ), .S(n8502), .Z(n7346)
         );
  MUX2_X1 U26303 ( .A(n7346), .B(n7345), .S(n8338), .Z(n7347) );
  MUX2_X1 U26304 ( .A(\mem[826][7] ), .B(\mem[827][7] ), .S(n8502), .Z(n7348)
         );
  MUX2_X1 U26305 ( .A(\mem[824][7] ), .B(\mem[825][7] ), .S(n8502), .Z(n7349)
         );
  MUX2_X1 U26306 ( .A(n7349), .B(n7348), .S(n8338), .Z(n7350) );
  MUX2_X1 U26307 ( .A(n7350), .B(n7347), .S(n8257), .Z(n7351) );
  MUX2_X1 U26308 ( .A(\mem[822][7] ), .B(\mem[823][7] ), .S(n8502), .Z(n7352)
         );
  MUX2_X1 U26309 ( .A(\mem[820][7] ), .B(\mem[821][7] ), .S(n8502), .Z(n7353)
         );
  MUX2_X1 U26310 ( .A(n7353), .B(n7352), .S(n8338), .Z(n7354) );
  MUX2_X1 U26311 ( .A(\mem[818][7] ), .B(\mem[819][7] ), .S(n8502), .Z(n7355)
         );
  MUX2_X1 U26312 ( .A(\mem[816][7] ), .B(\mem[817][7] ), .S(n8502), .Z(n7356)
         );
  MUX2_X1 U26313 ( .A(n7356), .B(n7355), .S(n8338), .Z(n7357) );
  MUX2_X1 U26314 ( .A(n7357), .B(n7354), .S(n8262), .Z(n7358) );
  MUX2_X1 U26315 ( .A(n7358), .B(n7351), .S(n8214), .Z(n7359) );
  MUX2_X1 U26316 ( .A(\mem[814][7] ), .B(\mem[815][7] ), .S(n8503), .Z(n7360)
         );
  MUX2_X1 U26317 ( .A(\mem[812][7] ), .B(\mem[813][7] ), .S(n8503), .Z(n7361)
         );
  MUX2_X1 U26318 ( .A(n7361), .B(n7360), .S(n8339), .Z(n7362) );
  MUX2_X1 U26319 ( .A(\mem[810][7] ), .B(\mem[811][7] ), .S(n8503), .Z(n7363)
         );
  MUX2_X1 U26320 ( .A(\mem[808][7] ), .B(\mem[809][7] ), .S(n8503), .Z(n7364)
         );
  MUX2_X1 U26321 ( .A(n7364), .B(n7363), .S(n8339), .Z(n7365) );
  MUX2_X1 U26322 ( .A(n7365), .B(n7362), .S(N20), .Z(n7366) );
  MUX2_X1 U26323 ( .A(\mem[806][7] ), .B(\mem[807][7] ), .S(n8503), .Z(n7367)
         );
  MUX2_X1 U26324 ( .A(\mem[804][7] ), .B(\mem[805][7] ), .S(n8503), .Z(n7368)
         );
  MUX2_X1 U26325 ( .A(n7368), .B(n7367), .S(n8339), .Z(n7369) );
  MUX2_X1 U26326 ( .A(\mem[802][7] ), .B(\mem[803][7] ), .S(n8503), .Z(n7370)
         );
  MUX2_X1 U26327 ( .A(\mem[800][7] ), .B(\mem[801][7] ), .S(n8503), .Z(n7371)
         );
  MUX2_X1 U26328 ( .A(n7371), .B(n7370), .S(n8339), .Z(n7372) );
  MUX2_X1 U26329 ( .A(n7372), .B(n7369), .S(n8241), .Z(n7373) );
  MUX2_X1 U26330 ( .A(n7373), .B(n7366), .S(n8214), .Z(n7374) );
  MUX2_X1 U26331 ( .A(n7374), .B(n7359), .S(n8192), .Z(n7375) );
  MUX2_X1 U26332 ( .A(\mem[798][7] ), .B(\mem[799][7] ), .S(n8503), .Z(n7376)
         );
  MUX2_X1 U26333 ( .A(\mem[796][7] ), .B(\mem[797][7] ), .S(n8503), .Z(n7377)
         );
  MUX2_X1 U26334 ( .A(n7377), .B(n7376), .S(n8339), .Z(n7378) );
  MUX2_X1 U26335 ( .A(\mem[794][7] ), .B(\mem[795][7] ), .S(n8503), .Z(n7379)
         );
  MUX2_X1 U26336 ( .A(\mem[792][7] ), .B(\mem[793][7] ), .S(n8503), .Z(n7380)
         );
  MUX2_X1 U26337 ( .A(n7380), .B(n7379), .S(n8339), .Z(n7381) );
  MUX2_X1 U26338 ( .A(n7381), .B(n7378), .S(n8263), .Z(n7382) );
  MUX2_X1 U26339 ( .A(\mem[790][7] ), .B(\mem[791][7] ), .S(n8504), .Z(n7383)
         );
  MUX2_X1 U26340 ( .A(\mem[788][7] ), .B(\mem[789][7] ), .S(n8504), .Z(n7384)
         );
  MUX2_X1 U26341 ( .A(n7384), .B(n7383), .S(n8339), .Z(n7385) );
  MUX2_X1 U26342 ( .A(\mem[786][7] ), .B(\mem[787][7] ), .S(n8504), .Z(n7386)
         );
  MUX2_X1 U26343 ( .A(\mem[784][7] ), .B(\mem[785][7] ), .S(n8504), .Z(n7387)
         );
  MUX2_X1 U26344 ( .A(n7387), .B(n7386), .S(n8339), .Z(n7388) );
  MUX2_X1 U26345 ( .A(n7388), .B(n7385), .S(n8264), .Z(n7389) );
  MUX2_X1 U26346 ( .A(n7389), .B(n7382), .S(n8214), .Z(n7390) );
  MUX2_X1 U26347 ( .A(\mem[782][7] ), .B(\mem[783][7] ), .S(n8504), .Z(n7391)
         );
  MUX2_X1 U26348 ( .A(\mem[780][7] ), .B(\mem[781][7] ), .S(n8504), .Z(n7392)
         );
  MUX2_X1 U26349 ( .A(n7392), .B(n7391), .S(n8339), .Z(n7393) );
  MUX2_X1 U26350 ( .A(\mem[778][7] ), .B(\mem[779][7] ), .S(n8504), .Z(n7394)
         );
  MUX2_X1 U26351 ( .A(\mem[776][7] ), .B(\mem[777][7] ), .S(n8504), .Z(n7395)
         );
  MUX2_X1 U26352 ( .A(n7395), .B(n7394), .S(n8339), .Z(n7396) );
  MUX2_X1 U26353 ( .A(n7396), .B(n7393), .S(n8255), .Z(n7397) );
  MUX2_X1 U26354 ( .A(\mem[774][7] ), .B(\mem[775][7] ), .S(n8504), .Z(n7398)
         );
  MUX2_X1 U26355 ( .A(\mem[772][7] ), .B(\mem[773][7] ), .S(n8504), .Z(n7399)
         );
  MUX2_X1 U26356 ( .A(n7399), .B(n7398), .S(n8339), .Z(n7400) );
  MUX2_X1 U26357 ( .A(\mem[770][7] ), .B(\mem[771][7] ), .S(n8504), .Z(n7401)
         );
  MUX2_X1 U26358 ( .A(\mem[768][7] ), .B(\mem[769][7] ), .S(n8504), .Z(n7402)
         );
  MUX2_X1 U26359 ( .A(n7402), .B(n7401), .S(n8339), .Z(n7403) );
  MUX2_X1 U26360 ( .A(n7403), .B(n7400), .S(n8222), .Z(n7404) );
  MUX2_X1 U26361 ( .A(n7404), .B(n7397), .S(n8214), .Z(n7405) );
  MUX2_X1 U26362 ( .A(n7405), .B(n7390), .S(n8192), .Z(n7406) );
  MUX2_X1 U26363 ( .A(n7406), .B(n7375), .S(N23), .Z(n7407) );
  MUX2_X1 U26364 ( .A(n7407), .B(n7344), .S(n8180), .Z(n7408) );
  MUX2_X1 U26365 ( .A(n7408), .B(n7281), .S(N25), .Z(n7409) );
  MUX2_X1 U26366 ( .A(\mem[766][7] ), .B(\mem[767][7] ), .S(n8505), .Z(n7410)
         );
  MUX2_X1 U26367 ( .A(\mem[764][7] ), .B(\mem[765][7] ), .S(n8505), .Z(n7411)
         );
  MUX2_X1 U26368 ( .A(n7411), .B(n7410), .S(n8340), .Z(n7412) );
  MUX2_X1 U26369 ( .A(\mem[762][7] ), .B(\mem[763][7] ), .S(n8505), .Z(n7413)
         );
  MUX2_X1 U26370 ( .A(\mem[760][7] ), .B(\mem[761][7] ), .S(n8505), .Z(n7414)
         );
  MUX2_X1 U26371 ( .A(n7414), .B(n7413), .S(n8340), .Z(n7415) );
  MUX2_X1 U26372 ( .A(n7415), .B(n7412), .S(n8258), .Z(n7416) );
  MUX2_X1 U26373 ( .A(\mem[758][7] ), .B(\mem[759][7] ), .S(n8505), .Z(n7417)
         );
  MUX2_X1 U26374 ( .A(\mem[756][7] ), .B(\mem[757][7] ), .S(n8505), .Z(n7418)
         );
  MUX2_X1 U26375 ( .A(n7418), .B(n7417), .S(n8340), .Z(n7419) );
  MUX2_X1 U26376 ( .A(\mem[754][7] ), .B(\mem[755][7] ), .S(n8505), .Z(n7420)
         );
  MUX2_X1 U26377 ( .A(\mem[752][7] ), .B(\mem[753][7] ), .S(n8505), .Z(n7421)
         );
  MUX2_X1 U26378 ( .A(n7421), .B(n7420), .S(n8340), .Z(n7422) );
  MUX2_X1 U26379 ( .A(n7422), .B(n7419), .S(n8235), .Z(n7423) );
  MUX2_X1 U26380 ( .A(n7423), .B(n7416), .S(n8215), .Z(n7424) );
  MUX2_X1 U26381 ( .A(\mem[750][7] ), .B(\mem[751][7] ), .S(n8505), .Z(n7425)
         );
  MUX2_X1 U26382 ( .A(\mem[748][7] ), .B(\mem[749][7] ), .S(n8505), .Z(n7426)
         );
  MUX2_X1 U26383 ( .A(n7426), .B(n7425), .S(n8340), .Z(n7427) );
  MUX2_X1 U26384 ( .A(\mem[746][7] ), .B(\mem[747][7] ), .S(n8505), .Z(n7428)
         );
  MUX2_X1 U26385 ( .A(\mem[744][7] ), .B(\mem[745][7] ), .S(n8505), .Z(n7429)
         );
  MUX2_X1 U26386 ( .A(n7429), .B(n7428), .S(n8340), .Z(n7430) );
  MUX2_X1 U26387 ( .A(n7430), .B(n7427), .S(n8236), .Z(n7431) );
  MUX2_X1 U26388 ( .A(\mem[742][7] ), .B(\mem[743][7] ), .S(n8506), .Z(n7432)
         );
  MUX2_X1 U26389 ( .A(\mem[740][7] ), .B(\mem[741][7] ), .S(n8506), .Z(n7433)
         );
  MUX2_X1 U26390 ( .A(n7433), .B(n7432), .S(n8340), .Z(n7434) );
  MUX2_X1 U26391 ( .A(\mem[738][7] ), .B(\mem[739][7] ), .S(n8506), .Z(n7435)
         );
  MUX2_X1 U26392 ( .A(\mem[736][7] ), .B(\mem[737][7] ), .S(n8506), .Z(n7436)
         );
  MUX2_X1 U26393 ( .A(n7436), .B(n7435), .S(n8340), .Z(n7437) );
  MUX2_X1 U26394 ( .A(n7437), .B(n7434), .S(n8237), .Z(n7438) );
  MUX2_X1 U26395 ( .A(n7438), .B(n7431), .S(n8215), .Z(n7439) );
  MUX2_X1 U26396 ( .A(n7439), .B(n7424), .S(n8193), .Z(n7440) );
  MUX2_X1 U26397 ( .A(\mem[734][7] ), .B(\mem[735][7] ), .S(n8506), .Z(n7441)
         );
  MUX2_X1 U26398 ( .A(\mem[732][7] ), .B(\mem[733][7] ), .S(n8506), .Z(n7442)
         );
  MUX2_X1 U26399 ( .A(n7442), .B(n7441), .S(n8340), .Z(n7443) );
  MUX2_X1 U26400 ( .A(\mem[730][7] ), .B(\mem[731][7] ), .S(n8506), .Z(n7444)
         );
  MUX2_X1 U26401 ( .A(\mem[728][7] ), .B(\mem[729][7] ), .S(n8506), .Z(n7445)
         );
  MUX2_X1 U26402 ( .A(n7445), .B(n7444), .S(n8340), .Z(n7446) );
  MUX2_X1 U26403 ( .A(n7446), .B(n7443), .S(n8232), .Z(n7447) );
  MUX2_X1 U26404 ( .A(\mem[726][7] ), .B(\mem[727][7] ), .S(n8506), .Z(n7448)
         );
  MUX2_X1 U26405 ( .A(\mem[724][7] ), .B(\mem[725][7] ), .S(n8506), .Z(n7449)
         );
  MUX2_X1 U26406 ( .A(n7449), .B(n7448), .S(n8340), .Z(n7450) );
  MUX2_X1 U26407 ( .A(\mem[722][7] ), .B(\mem[723][7] ), .S(n8506), .Z(n7451)
         );
  MUX2_X1 U26408 ( .A(\mem[720][7] ), .B(\mem[721][7] ), .S(n8506), .Z(n7452)
         );
  MUX2_X1 U26409 ( .A(n7452), .B(n7451), .S(n8340), .Z(n7453) );
  MUX2_X1 U26410 ( .A(n7453), .B(n7450), .S(n8233), .Z(n7454) );
  MUX2_X1 U26411 ( .A(n7454), .B(n7447), .S(n8215), .Z(n7455) );
  MUX2_X1 U26412 ( .A(\mem[718][7] ), .B(\mem[719][7] ), .S(n8507), .Z(n7456)
         );
  MUX2_X1 U26413 ( .A(\mem[716][7] ), .B(\mem[717][7] ), .S(n8507), .Z(n7457)
         );
  MUX2_X1 U26414 ( .A(n7457), .B(n7456), .S(n8341), .Z(n7458) );
  MUX2_X1 U26415 ( .A(\mem[714][7] ), .B(\mem[715][7] ), .S(n8507), .Z(n7459)
         );
  MUX2_X1 U26416 ( .A(\mem[712][7] ), .B(\mem[713][7] ), .S(n8507), .Z(n7460)
         );
  MUX2_X1 U26417 ( .A(n7460), .B(n7459), .S(n8341), .Z(n7461) );
  MUX2_X1 U26418 ( .A(n7461), .B(n7458), .S(n8234), .Z(n7462) );
  MUX2_X1 U26419 ( .A(\mem[710][7] ), .B(\mem[711][7] ), .S(n8507), .Z(n7463)
         );
  MUX2_X1 U26420 ( .A(\mem[708][7] ), .B(\mem[709][7] ), .S(n8507), .Z(n7464)
         );
  MUX2_X1 U26421 ( .A(n7464), .B(n7463), .S(n8341), .Z(n7465) );
  MUX2_X1 U26422 ( .A(\mem[706][7] ), .B(\mem[707][7] ), .S(n8507), .Z(n7466)
         );
  MUX2_X1 U26423 ( .A(\mem[704][7] ), .B(\mem[705][7] ), .S(n8507), .Z(n7467)
         );
  MUX2_X1 U26424 ( .A(n7467), .B(n7466), .S(n8341), .Z(n7468) );
  MUX2_X1 U26425 ( .A(n7468), .B(n7465), .S(n8230), .Z(n7469) );
  MUX2_X1 U26426 ( .A(n7469), .B(n7462), .S(n8215), .Z(n7470) );
  MUX2_X1 U26427 ( .A(n7470), .B(n7455), .S(n8193), .Z(n7471) );
  MUX2_X1 U26428 ( .A(n7471), .B(n7440), .S(n8183), .Z(n7472) );
  MUX2_X1 U26429 ( .A(\mem[702][7] ), .B(\mem[703][7] ), .S(n8507), .Z(n7473)
         );
  MUX2_X1 U26430 ( .A(\mem[700][7] ), .B(\mem[701][7] ), .S(n8507), .Z(n7474)
         );
  MUX2_X1 U26431 ( .A(n7474), .B(n7473), .S(n8341), .Z(n7475) );
  MUX2_X1 U26432 ( .A(\mem[698][7] ), .B(\mem[699][7] ), .S(n8507), .Z(n7476)
         );
  MUX2_X1 U26433 ( .A(\mem[696][7] ), .B(\mem[697][7] ), .S(n8507), .Z(n7477)
         );
  MUX2_X1 U26434 ( .A(n7477), .B(n7476), .S(n8341), .Z(n7478) );
  MUX2_X1 U26435 ( .A(n7478), .B(n7475), .S(n8231), .Z(n7479) );
  MUX2_X1 U26436 ( .A(\mem[694][7] ), .B(\mem[695][7] ), .S(n8508), .Z(n7480)
         );
  MUX2_X1 U26437 ( .A(\mem[692][7] ), .B(\mem[693][7] ), .S(n8508), .Z(n7481)
         );
  MUX2_X1 U26438 ( .A(n7481), .B(n7480), .S(n8341), .Z(n7482) );
  MUX2_X1 U26439 ( .A(\mem[690][7] ), .B(\mem[691][7] ), .S(n8508), .Z(n7483)
         );
  MUX2_X1 U26440 ( .A(\mem[688][7] ), .B(\mem[689][7] ), .S(n8508), .Z(n7484)
         );
  MUX2_X1 U26441 ( .A(n7484), .B(n7483), .S(n8341), .Z(n7485) );
  MUX2_X1 U26442 ( .A(n7485), .B(n7482), .S(n8227), .Z(n7486) );
  MUX2_X1 U26443 ( .A(n7486), .B(n7479), .S(n8215), .Z(n7487) );
  MUX2_X1 U26444 ( .A(\mem[686][7] ), .B(\mem[687][7] ), .S(n8508), .Z(n7488)
         );
  MUX2_X1 U26445 ( .A(\mem[684][7] ), .B(\mem[685][7] ), .S(n8508), .Z(n7489)
         );
  MUX2_X1 U26446 ( .A(n7489), .B(n7488), .S(n8341), .Z(n7490) );
  MUX2_X1 U26447 ( .A(\mem[682][7] ), .B(\mem[683][7] ), .S(n8508), .Z(n7491)
         );
  MUX2_X1 U26448 ( .A(\mem[680][7] ), .B(\mem[681][7] ), .S(n8508), .Z(n7492)
         );
  MUX2_X1 U26449 ( .A(n7492), .B(n7491), .S(n8341), .Z(n7493) );
  MUX2_X1 U26450 ( .A(n7493), .B(n7490), .S(n8246), .Z(n7494) );
  MUX2_X1 U26451 ( .A(\mem[678][7] ), .B(\mem[679][7] ), .S(n8508), .Z(n7495)
         );
  MUX2_X1 U26452 ( .A(\mem[676][7] ), .B(\mem[677][7] ), .S(n8508), .Z(n7496)
         );
  MUX2_X1 U26453 ( .A(n7496), .B(n7495), .S(n8341), .Z(n7497) );
  MUX2_X1 U26454 ( .A(\mem[674][7] ), .B(\mem[675][7] ), .S(n8508), .Z(n7498)
         );
  MUX2_X1 U26455 ( .A(\mem[672][7] ), .B(\mem[673][7] ), .S(n8508), .Z(n7499)
         );
  MUX2_X1 U26456 ( .A(n7499), .B(n7498), .S(n8341), .Z(n7500) );
  MUX2_X1 U26457 ( .A(n7500), .B(n7497), .S(n8262), .Z(n7501) );
  MUX2_X1 U26458 ( .A(n7501), .B(n7494), .S(n8215), .Z(n7502) );
  MUX2_X1 U26459 ( .A(n7502), .B(n7487), .S(n8193), .Z(n7503) );
  MUX2_X1 U26460 ( .A(\mem[670][7] ), .B(\mem[671][7] ), .S(n8509), .Z(n7504)
         );
  MUX2_X1 U26461 ( .A(\mem[668][7] ), .B(\mem[669][7] ), .S(n8509), .Z(n7505)
         );
  MUX2_X1 U26462 ( .A(n7505), .B(n7504), .S(n8342), .Z(n7506) );
  MUX2_X1 U26463 ( .A(\mem[666][7] ), .B(\mem[667][7] ), .S(n8509), .Z(n7507)
         );
  MUX2_X1 U26464 ( .A(\mem[664][7] ), .B(\mem[665][7] ), .S(n8509), .Z(n7508)
         );
  MUX2_X1 U26465 ( .A(n7508), .B(n7507), .S(n8342), .Z(n7509) );
  MUX2_X1 U26466 ( .A(n7509), .B(n7506), .S(n8235), .Z(n7510) );
  MUX2_X1 U26467 ( .A(\mem[662][7] ), .B(\mem[663][7] ), .S(n8509), .Z(n7511)
         );
  MUX2_X1 U26468 ( .A(\mem[660][7] ), .B(\mem[661][7] ), .S(n8509), .Z(n7512)
         );
  MUX2_X1 U26469 ( .A(n7512), .B(n7511), .S(n8342), .Z(n7513) );
  MUX2_X1 U26470 ( .A(\mem[658][7] ), .B(\mem[659][7] ), .S(n8509), .Z(n7514)
         );
  MUX2_X1 U26471 ( .A(\mem[656][7] ), .B(\mem[657][7] ), .S(n8509), .Z(n7515)
         );
  MUX2_X1 U26472 ( .A(n7515), .B(n7514), .S(n8342), .Z(n7516) );
  MUX2_X1 U26473 ( .A(n7516), .B(n7513), .S(n8247), .Z(n7517) );
  MUX2_X1 U26474 ( .A(n7517), .B(n7510), .S(n8215), .Z(n7518) );
  MUX2_X1 U26475 ( .A(\mem[654][7] ), .B(\mem[655][7] ), .S(n8509), .Z(n7519)
         );
  MUX2_X1 U26476 ( .A(\mem[652][7] ), .B(\mem[653][7] ), .S(n8509), .Z(n7520)
         );
  MUX2_X1 U26477 ( .A(n7520), .B(n7519), .S(n8342), .Z(n7521) );
  MUX2_X1 U26478 ( .A(\mem[650][7] ), .B(\mem[651][7] ), .S(n8509), .Z(n7522)
         );
  MUX2_X1 U26479 ( .A(\mem[648][7] ), .B(\mem[649][7] ), .S(n8509), .Z(n7523)
         );
  MUX2_X1 U26480 ( .A(n7523), .B(n7522), .S(n8342), .Z(n7524) );
  MUX2_X1 U26481 ( .A(n7524), .B(n7521), .S(n8248), .Z(n7525) );
  MUX2_X1 U26482 ( .A(\mem[646][7] ), .B(\mem[647][7] ), .S(n8510), .Z(n7526)
         );
  MUX2_X1 U26483 ( .A(\mem[644][7] ), .B(\mem[645][7] ), .S(n8510), .Z(n7527)
         );
  MUX2_X1 U26484 ( .A(n7527), .B(n7526), .S(n8342), .Z(n7528) );
  MUX2_X1 U26485 ( .A(\mem[642][7] ), .B(\mem[643][7] ), .S(n8510), .Z(n7529)
         );
  MUX2_X1 U26486 ( .A(\mem[640][7] ), .B(\mem[641][7] ), .S(n8510), .Z(n7530)
         );
  MUX2_X1 U26487 ( .A(n7530), .B(n7529), .S(n8342), .Z(n7531) );
  MUX2_X1 U26488 ( .A(n7531), .B(n7528), .S(n8249), .Z(n7532) );
  MUX2_X1 U26489 ( .A(n7532), .B(n7525), .S(n8215), .Z(n7533) );
  MUX2_X1 U26490 ( .A(n7533), .B(n7518), .S(n8193), .Z(n7534) );
  MUX2_X1 U26491 ( .A(n7534), .B(n7503), .S(n8185), .Z(n7535) );
  MUX2_X1 U26492 ( .A(n7535), .B(n7472), .S(n8180), .Z(n7536) );
  MUX2_X1 U26493 ( .A(\mem[638][7] ), .B(\mem[639][7] ), .S(n8510), .Z(n7537)
         );
  MUX2_X1 U26494 ( .A(\mem[636][7] ), .B(\mem[637][7] ), .S(n8510), .Z(n7538)
         );
  MUX2_X1 U26495 ( .A(n7538), .B(n7537), .S(n8342), .Z(n7539) );
  MUX2_X1 U26496 ( .A(\mem[634][7] ), .B(\mem[635][7] ), .S(n8510), .Z(n7540)
         );
  MUX2_X1 U26497 ( .A(\mem[632][7] ), .B(\mem[633][7] ), .S(n8510), .Z(n7541)
         );
  MUX2_X1 U26498 ( .A(n7541), .B(n7540), .S(n8342), .Z(n7542) );
  MUX2_X1 U26499 ( .A(n7542), .B(n7539), .S(n8244), .Z(n7543) );
  MUX2_X1 U26500 ( .A(\mem[630][7] ), .B(\mem[631][7] ), .S(n8510), .Z(n7544)
         );
  MUX2_X1 U26501 ( .A(\mem[628][7] ), .B(\mem[629][7] ), .S(n8510), .Z(n7545)
         );
  MUX2_X1 U26502 ( .A(n7545), .B(n7544), .S(n8342), .Z(n7546) );
  MUX2_X1 U26503 ( .A(\mem[626][7] ), .B(\mem[627][7] ), .S(n8510), .Z(n7547)
         );
  MUX2_X1 U26504 ( .A(\mem[624][7] ), .B(\mem[625][7] ), .S(n8510), .Z(n7548)
         );
  MUX2_X1 U26505 ( .A(n7548), .B(n7547), .S(n8342), .Z(n7549) );
  MUX2_X1 U26506 ( .A(n7549), .B(n7546), .S(n8245), .Z(n7550) );
  MUX2_X1 U26507 ( .A(n7550), .B(n7543), .S(n8215), .Z(n7551) );
  MUX2_X1 U26508 ( .A(\mem[622][7] ), .B(\mem[623][7] ), .S(n8511), .Z(n7552)
         );
  MUX2_X1 U26509 ( .A(\mem[620][7] ), .B(\mem[621][7] ), .S(n8511), .Z(n7553)
         );
  MUX2_X1 U26510 ( .A(n7553), .B(n7552), .S(n8343), .Z(n7554) );
  MUX2_X1 U26511 ( .A(\mem[618][7] ), .B(\mem[619][7] ), .S(n8511), .Z(n7555)
         );
  MUX2_X1 U26512 ( .A(\mem[616][7] ), .B(\mem[617][7] ), .S(n8511), .Z(n7556)
         );
  MUX2_X1 U26513 ( .A(n7556), .B(n7555), .S(n8343), .Z(n7557) );
  MUX2_X1 U26514 ( .A(n7557), .B(n7554), .S(n8246), .Z(n7558) );
  MUX2_X1 U26515 ( .A(\mem[614][7] ), .B(\mem[615][7] ), .S(n8511), .Z(n7559)
         );
  MUX2_X1 U26516 ( .A(\mem[612][7] ), .B(\mem[613][7] ), .S(n8511), .Z(n7560)
         );
  MUX2_X1 U26517 ( .A(n7560), .B(n7559), .S(n8343), .Z(n7561) );
  MUX2_X1 U26518 ( .A(\mem[610][7] ), .B(\mem[611][7] ), .S(n8511), .Z(n7562)
         );
  MUX2_X1 U26519 ( .A(\mem[608][7] ), .B(\mem[609][7] ), .S(n8511), .Z(n7563)
         );
  MUX2_X1 U26520 ( .A(n7563), .B(n7562), .S(n8343), .Z(n7564) );
  MUX2_X1 U26521 ( .A(n7564), .B(n7561), .S(n8253), .Z(n7565) );
  MUX2_X1 U26522 ( .A(n7565), .B(n7558), .S(n8215), .Z(n7566) );
  MUX2_X1 U26523 ( .A(n7566), .B(n7551), .S(n8193), .Z(n7567) );
  MUX2_X1 U26524 ( .A(\mem[606][7] ), .B(\mem[607][7] ), .S(n8511), .Z(n7568)
         );
  MUX2_X1 U26525 ( .A(\mem[604][7] ), .B(\mem[605][7] ), .S(n8511), .Z(n7569)
         );
  MUX2_X1 U26526 ( .A(n7569), .B(n7568), .S(n8343), .Z(n7570) );
  MUX2_X1 U26527 ( .A(\mem[602][7] ), .B(\mem[603][7] ), .S(n8511), .Z(n7571)
         );
  MUX2_X1 U26528 ( .A(\mem[600][7] ), .B(\mem[601][7] ), .S(n8511), .Z(n7572)
         );
  MUX2_X1 U26529 ( .A(n7572), .B(n7571), .S(n8343), .Z(n7573) );
  MUX2_X1 U26530 ( .A(n7573), .B(n7570), .S(n8254), .Z(n7574) );
  MUX2_X1 U26531 ( .A(\mem[598][7] ), .B(\mem[599][7] ), .S(n8512), .Z(n7575)
         );
  MUX2_X1 U26532 ( .A(\mem[596][7] ), .B(\mem[597][7] ), .S(n8512), .Z(n7576)
         );
  MUX2_X1 U26533 ( .A(n7576), .B(n7575), .S(n8343), .Z(n7577) );
  MUX2_X1 U26534 ( .A(\mem[594][7] ), .B(\mem[595][7] ), .S(n8512), .Z(n7578)
         );
  MUX2_X1 U26535 ( .A(\mem[592][7] ), .B(\mem[593][7] ), .S(n8512), .Z(n7579)
         );
  MUX2_X1 U26536 ( .A(n7579), .B(n7578), .S(n8343), .Z(n7580) );
  MUX2_X1 U26537 ( .A(n7580), .B(n7577), .S(n8255), .Z(n7581) );
  MUX2_X1 U26538 ( .A(n7581), .B(n7574), .S(n8215), .Z(n7582) );
  MUX2_X1 U26539 ( .A(\mem[590][7] ), .B(\mem[591][7] ), .S(n8512), .Z(n7583)
         );
  MUX2_X1 U26540 ( .A(\mem[588][7] ), .B(\mem[589][7] ), .S(n8512), .Z(n7584)
         );
  MUX2_X1 U26541 ( .A(n7584), .B(n7583), .S(n8343), .Z(n7585) );
  MUX2_X1 U26542 ( .A(\mem[586][7] ), .B(\mem[587][7] ), .S(n8512), .Z(n7586)
         );
  MUX2_X1 U26543 ( .A(\mem[584][7] ), .B(\mem[585][7] ), .S(n8512), .Z(n7587)
         );
  MUX2_X1 U26544 ( .A(n7587), .B(n7586), .S(n8343), .Z(n7588) );
  MUX2_X1 U26545 ( .A(n7588), .B(n7585), .S(n8250), .Z(n7589) );
  MUX2_X1 U26546 ( .A(\mem[582][7] ), .B(\mem[583][7] ), .S(n8512), .Z(n7590)
         );
  MUX2_X1 U26547 ( .A(\mem[580][7] ), .B(\mem[581][7] ), .S(n8512), .Z(n7591)
         );
  MUX2_X1 U26548 ( .A(n7591), .B(n7590), .S(n8343), .Z(n7592) );
  MUX2_X1 U26549 ( .A(\mem[578][7] ), .B(\mem[579][7] ), .S(n8512), .Z(n7593)
         );
  MUX2_X1 U26550 ( .A(\mem[576][7] ), .B(\mem[577][7] ), .S(n8512), .Z(n7594)
         );
  MUX2_X1 U26551 ( .A(n7594), .B(n7593), .S(n8343), .Z(n7595) );
  MUX2_X1 U26552 ( .A(n7595), .B(n7592), .S(n8251), .Z(n7596) );
  MUX2_X1 U26553 ( .A(n7596), .B(n7589), .S(n8215), .Z(n7597) );
  MUX2_X1 U26554 ( .A(n7597), .B(n7582), .S(n8193), .Z(n7598) );
  MUX2_X1 U26555 ( .A(n7598), .B(n7567), .S(n8185), .Z(n7599) );
  MUX2_X1 U26556 ( .A(\mem[574][7] ), .B(\mem[575][7] ), .S(n8513), .Z(n7600)
         );
  MUX2_X1 U26557 ( .A(\mem[572][7] ), .B(\mem[573][7] ), .S(n8513), .Z(n7601)
         );
  MUX2_X1 U26558 ( .A(n7601), .B(n7600), .S(n8344), .Z(n7602) );
  MUX2_X1 U26559 ( .A(\mem[570][7] ), .B(\mem[571][7] ), .S(n8513), .Z(n7603)
         );
  MUX2_X1 U26560 ( .A(\mem[568][7] ), .B(\mem[569][7] ), .S(n8513), .Z(n7604)
         );
  MUX2_X1 U26561 ( .A(n7604), .B(n7603), .S(n8344), .Z(n7605) );
  MUX2_X1 U26562 ( .A(n7605), .B(n7602), .S(n8224), .Z(n7606) );
  MUX2_X1 U26563 ( .A(\mem[566][7] ), .B(\mem[567][7] ), .S(n8513), .Z(n7607)
         );
  MUX2_X1 U26564 ( .A(\mem[564][7] ), .B(\mem[565][7] ), .S(n8513), .Z(n7608)
         );
  MUX2_X1 U26565 ( .A(n7608), .B(n7607), .S(n8344), .Z(n7609) );
  MUX2_X1 U26566 ( .A(\mem[562][7] ), .B(\mem[563][7] ), .S(n8513), .Z(n7610)
         );
  MUX2_X1 U26567 ( .A(\mem[560][7] ), .B(\mem[561][7] ), .S(n8513), .Z(n7611)
         );
  MUX2_X1 U26568 ( .A(n7611), .B(n7610), .S(n8344), .Z(n7612) );
  MUX2_X1 U26569 ( .A(n7612), .B(n7609), .S(n8238), .Z(n7613) );
  MUX2_X1 U26570 ( .A(n7613), .B(n7606), .S(n8216), .Z(n7614) );
  MUX2_X1 U26571 ( .A(\mem[558][7] ), .B(\mem[559][7] ), .S(n8513), .Z(n7615)
         );
  MUX2_X1 U26572 ( .A(\mem[556][7] ), .B(\mem[557][7] ), .S(n8513), .Z(n7616)
         );
  MUX2_X1 U26573 ( .A(n7616), .B(n7615), .S(n8344), .Z(n7617) );
  MUX2_X1 U26574 ( .A(\mem[554][7] ), .B(\mem[555][7] ), .S(n8513), .Z(n7618)
         );
  MUX2_X1 U26575 ( .A(\mem[552][7] ), .B(\mem[553][7] ), .S(n8513), .Z(n7619)
         );
  MUX2_X1 U26576 ( .A(n7619), .B(n7618), .S(n8344), .Z(n7620) );
  MUX2_X1 U26577 ( .A(n7620), .B(n7617), .S(n8252), .Z(n7621) );
  MUX2_X1 U26578 ( .A(\mem[550][7] ), .B(\mem[551][7] ), .S(n8514), .Z(n7622)
         );
  MUX2_X1 U26579 ( .A(\mem[548][7] ), .B(\mem[549][7] ), .S(n8514), .Z(n7623)
         );
  MUX2_X1 U26580 ( .A(n7623), .B(n7622), .S(n8344), .Z(n7624) );
  MUX2_X1 U26581 ( .A(\mem[546][7] ), .B(\mem[547][7] ), .S(n8514), .Z(n7625)
         );
  MUX2_X1 U26582 ( .A(\mem[544][7] ), .B(\mem[545][7] ), .S(n8514), .Z(n7626)
         );
  MUX2_X1 U26583 ( .A(n7626), .B(n7625), .S(n8344), .Z(n7627) );
  MUX2_X1 U26584 ( .A(n7627), .B(n7624), .S(N20), .Z(n7628) );
  MUX2_X1 U26585 ( .A(n7628), .B(n7621), .S(n8216), .Z(n7629) );
  MUX2_X1 U26586 ( .A(n7629), .B(n7614), .S(n8193), .Z(n7630) );
  MUX2_X1 U26587 ( .A(\mem[542][7] ), .B(\mem[543][7] ), .S(n8514), .Z(n7631)
         );
  MUX2_X1 U26588 ( .A(\mem[540][7] ), .B(\mem[541][7] ), .S(n8514), .Z(n7632)
         );
  MUX2_X1 U26589 ( .A(n7632), .B(n7631), .S(n8344), .Z(n7633) );
  MUX2_X1 U26590 ( .A(\mem[538][7] ), .B(\mem[539][7] ), .S(n8514), .Z(n7634)
         );
  MUX2_X1 U26591 ( .A(\mem[536][7] ), .B(\mem[537][7] ), .S(n8514), .Z(n7635)
         );
  MUX2_X1 U26592 ( .A(n7635), .B(n7634), .S(n8344), .Z(n7636) );
  MUX2_X1 U26593 ( .A(n7636), .B(n7633), .S(n8245), .Z(n7637) );
  MUX2_X1 U26594 ( .A(\mem[534][7] ), .B(\mem[535][7] ), .S(n8514), .Z(n7638)
         );
  MUX2_X1 U26595 ( .A(\mem[532][7] ), .B(\mem[533][7] ), .S(n8514), .Z(n7639)
         );
  MUX2_X1 U26596 ( .A(n7639), .B(n7638), .S(n8344), .Z(n7640) );
  MUX2_X1 U26597 ( .A(\mem[530][7] ), .B(\mem[531][7] ), .S(n8514), .Z(n7641)
         );
  MUX2_X1 U26598 ( .A(\mem[528][7] ), .B(\mem[529][7] ), .S(n8514), .Z(n7642)
         );
  MUX2_X1 U26599 ( .A(n7642), .B(n7641), .S(n8344), .Z(n7643) );
  MUX2_X1 U26600 ( .A(n7643), .B(n7640), .S(n8263), .Z(n7644) );
  MUX2_X1 U26601 ( .A(n7644), .B(n7637), .S(n8216), .Z(n7645) );
  MUX2_X1 U26602 ( .A(\mem[526][7] ), .B(\mem[527][7] ), .S(n8515), .Z(n7646)
         );
  MUX2_X1 U26603 ( .A(\mem[524][7] ), .B(\mem[525][7] ), .S(n8515), .Z(n7647)
         );
  MUX2_X1 U26604 ( .A(n7647), .B(n7646), .S(n8345), .Z(n7648) );
  MUX2_X1 U26605 ( .A(\mem[522][7] ), .B(\mem[523][7] ), .S(n8515), .Z(n7649)
         );
  MUX2_X1 U26606 ( .A(\mem[520][7] ), .B(\mem[521][7] ), .S(n8515), .Z(n7650)
         );
  MUX2_X1 U26607 ( .A(n7650), .B(n7649), .S(n8345), .Z(n7651) );
  MUX2_X1 U26608 ( .A(n7651), .B(n7648), .S(n8229), .Z(n7652) );
  MUX2_X1 U26609 ( .A(\mem[518][7] ), .B(\mem[519][7] ), .S(n8515), .Z(n7653)
         );
  MUX2_X1 U26610 ( .A(\mem[516][7] ), .B(\mem[517][7] ), .S(n8515), .Z(n7654)
         );
  MUX2_X1 U26611 ( .A(n7654), .B(n7653), .S(n8345), .Z(n7655) );
  MUX2_X1 U26612 ( .A(\mem[514][7] ), .B(\mem[515][7] ), .S(n8515), .Z(n7656)
         );
  MUX2_X1 U26613 ( .A(\mem[512][7] ), .B(\mem[513][7] ), .S(n8515), .Z(n7657)
         );
  MUX2_X1 U26614 ( .A(n7657), .B(n7656), .S(n8345), .Z(n7658) );
  MUX2_X1 U26615 ( .A(n7658), .B(n7655), .S(n8223), .Z(n7659) );
  MUX2_X1 U26616 ( .A(n7659), .B(n7652), .S(n8216), .Z(n7660) );
  MUX2_X1 U26617 ( .A(n7660), .B(n7645), .S(n8193), .Z(n7661) );
  MUX2_X1 U26618 ( .A(n7661), .B(n7630), .S(N23), .Z(n7662) );
  MUX2_X1 U26619 ( .A(n7662), .B(n7599), .S(n8180), .Z(n7663) );
  MUX2_X1 U26620 ( .A(n7663), .B(n7536), .S(n8177), .Z(n7664) );
  MUX2_X1 U26621 ( .A(n7664), .B(n7409), .S(N26), .Z(n7665) );
  MUX2_X1 U26622 ( .A(\mem[510][7] ), .B(\mem[511][7] ), .S(n8515), .Z(n7666)
         );
  MUX2_X1 U26623 ( .A(\mem[508][7] ), .B(\mem[509][7] ), .S(n8515), .Z(n7667)
         );
  MUX2_X1 U26624 ( .A(n7667), .B(n7666), .S(n8345), .Z(n7668) );
  MUX2_X1 U26625 ( .A(\mem[506][7] ), .B(\mem[507][7] ), .S(n8515), .Z(n7669)
         );
  MUX2_X1 U26626 ( .A(\mem[504][7] ), .B(\mem[505][7] ), .S(n8515), .Z(n7670)
         );
  MUX2_X1 U26627 ( .A(n7670), .B(n7669), .S(n8345), .Z(n7671) );
  MUX2_X1 U26628 ( .A(n7671), .B(n7668), .S(n8228), .Z(n7672) );
  MUX2_X1 U26629 ( .A(\mem[502][7] ), .B(\mem[503][7] ), .S(n8516), .Z(n7673)
         );
  MUX2_X1 U26630 ( .A(\mem[500][7] ), .B(\mem[501][7] ), .S(n8516), .Z(n7674)
         );
  MUX2_X1 U26631 ( .A(n7674), .B(n7673), .S(n8345), .Z(n7675) );
  MUX2_X1 U26632 ( .A(\mem[498][7] ), .B(\mem[499][7] ), .S(n8516), .Z(n7676)
         );
  MUX2_X1 U26633 ( .A(\mem[496][7] ), .B(\mem[497][7] ), .S(n8516), .Z(n7677)
         );
  MUX2_X1 U26634 ( .A(n7677), .B(n7676), .S(n8345), .Z(n7678) );
  MUX2_X1 U26635 ( .A(n7678), .B(n7675), .S(n8229), .Z(n7679) );
  MUX2_X1 U26636 ( .A(n7679), .B(n7672), .S(n8216), .Z(n7680) );
  MUX2_X1 U26637 ( .A(\mem[494][7] ), .B(\mem[495][7] ), .S(n8516), .Z(n7681)
         );
  MUX2_X1 U26638 ( .A(\mem[492][7] ), .B(\mem[493][7] ), .S(n8516), .Z(n7682)
         );
  MUX2_X1 U26639 ( .A(n7682), .B(n7681), .S(n8345), .Z(n7683) );
  MUX2_X1 U26640 ( .A(\mem[490][7] ), .B(\mem[491][7] ), .S(n8516), .Z(n7684)
         );
  MUX2_X1 U26641 ( .A(\mem[488][7] ), .B(\mem[489][7] ), .S(n8516), .Z(n7685)
         );
  MUX2_X1 U26642 ( .A(n7685), .B(n7684), .S(n8345), .Z(n7686) );
  MUX2_X1 U26643 ( .A(n7686), .B(n7683), .S(n8225), .Z(n7687) );
  MUX2_X1 U26644 ( .A(\mem[486][7] ), .B(\mem[487][7] ), .S(n8516), .Z(n7688)
         );
  MUX2_X1 U26645 ( .A(\mem[484][7] ), .B(\mem[485][7] ), .S(n8516), .Z(n7689)
         );
  MUX2_X1 U26646 ( .A(n7689), .B(n7688), .S(n8345), .Z(n7690) );
  MUX2_X1 U26647 ( .A(\mem[482][7] ), .B(\mem[483][7] ), .S(n8516), .Z(n7691)
         );
  MUX2_X1 U26648 ( .A(\mem[480][7] ), .B(\mem[481][7] ), .S(n8516), .Z(n7692)
         );
  MUX2_X1 U26649 ( .A(n7692), .B(n7691), .S(n8345), .Z(n7693) );
  MUX2_X1 U26650 ( .A(n7693), .B(n7690), .S(n8222), .Z(n7694) );
  MUX2_X1 U26651 ( .A(n7694), .B(n7687), .S(n8216), .Z(n7695) );
  MUX2_X1 U26652 ( .A(n7695), .B(n7680), .S(n8193), .Z(n7696) );
  MUX2_X1 U26653 ( .A(\mem[478][7] ), .B(\mem[479][7] ), .S(n8517), .Z(n7697)
         );
  MUX2_X1 U26654 ( .A(\mem[476][7] ), .B(\mem[477][7] ), .S(n8517), .Z(n7698)
         );
  MUX2_X1 U26655 ( .A(n7698), .B(n7697), .S(n8346), .Z(n7699) );
  MUX2_X1 U26656 ( .A(\mem[474][7] ), .B(\mem[475][7] ), .S(n8517), .Z(n7700)
         );
  MUX2_X1 U26657 ( .A(\mem[472][7] ), .B(\mem[473][7] ), .S(n8517), .Z(n7701)
         );
  MUX2_X1 U26658 ( .A(n7701), .B(n7700), .S(n8346), .Z(n7702) );
  MUX2_X1 U26659 ( .A(n7702), .B(n7699), .S(n8232), .Z(n7703) );
  MUX2_X1 U26660 ( .A(\mem[470][7] ), .B(\mem[471][7] ), .S(n8517), .Z(n7704)
         );
  MUX2_X1 U26661 ( .A(\mem[468][7] ), .B(\mem[469][7] ), .S(n8517), .Z(n7705)
         );
  MUX2_X1 U26662 ( .A(n7705), .B(n7704), .S(n8346), .Z(n7706) );
  MUX2_X1 U26663 ( .A(\mem[466][7] ), .B(\mem[467][7] ), .S(n8517), .Z(n7707)
         );
  MUX2_X1 U26664 ( .A(\mem[464][7] ), .B(\mem[465][7] ), .S(n8517), .Z(n7708)
         );
  MUX2_X1 U26665 ( .A(n7708), .B(n7707), .S(n8346), .Z(n7709) );
  MUX2_X1 U26666 ( .A(n7709), .B(n7706), .S(n8233), .Z(n7710) );
  MUX2_X1 U26667 ( .A(n7710), .B(n7703), .S(n8216), .Z(n7711) );
  MUX2_X1 U26668 ( .A(\mem[462][7] ), .B(\mem[463][7] ), .S(n8517), .Z(n7712)
         );
  MUX2_X1 U26669 ( .A(\mem[460][7] ), .B(\mem[461][7] ), .S(n8517), .Z(n7713)
         );
  MUX2_X1 U26670 ( .A(n7713), .B(n7712), .S(n8346), .Z(n7714) );
  MUX2_X1 U26671 ( .A(\mem[458][7] ), .B(\mem[459][7] ), .S(n8517), .Z(n7715)
         );
  MUX2_X1 U26672 ( .A(\mem[456][7] ), .B(\mem[457][7] ), .S(n8517), .Z(n7716)
         );
  MUX2_X1 U26673 ( .A(n7716), .B(n7715), .S(n8346), .Z(n7717) );
  MUX2_X1 U26674 ( .A(n7717), .B(n7714), .S(n8234), .Z(n7718) );
  MUX2_X1 U26675 ( .A(\mem[454][7] ), .B(\mem[455][7] ), .S(n8518), .Z(n7719)
         );
  MUX2_X1 U26676 ( .A(\mem[452][7] ), .B(\mem[453][7] ), .S(n8518), .Z(n7720)
         );
  MUX2_X1 U26677 ( .A(n7720), .B(n7719), .S(n8346), .Z(n7721) );
  MUX2_X1 U26678 ( .A(\mem[450][7] ), .B(\mem[451][7] ), .S(n8518), .Z(n7722)
         );
  MUX2_X1 U26679 ( .A(\mem[448][7] ), .B(\mem[449][7] ), .S(n8518), .Z(n7723)
         );
  MUX2_X1 U26680 ( .A(n7723), .B(n7722), .S(n8346), .Z(n7724) );
  MUX2_X1 U26681 ( .A(n7724), .B(n7721), .S(n8230), .Z(n7725) );
  MUX2_X1 U26682 ( .A(n7725), .B(n7718), .S(n8216), .Z(n7726) );
  MUX2_X1 U26683 ( .A(n7726), .B(n7711), .S(n8193), .Z(n7727) );
  MUX2_X1 U26684 ( .A(n7727), .B(n7696), .S(n8181), .Z(n7728) );
  MUX2_X1 U26685 ( .A(\mem[446][7] ), .B(\mem[447][7] ), .S(n8518), .Z(n7729)
         );
  MUX2_X1 U26686 ( .A(\mem[444][7] ), .B(\mem[445][7] ), .S(n8518), .Z(n7730)
         );
  MUX2_X1 U26687 ( .A(n7730), .B(n7729), .S(n8346), .Z(n7731) );
  MUX2_X1 U26688 ( .A(\mem[442][7] ), .B(\mem[443][7] ), .S(n8518), .Z(n7732)
         );
  MUX2_X1 U26689 ( .A(\mem[440][7] ), .B(\mem[441][7] ), .S(n8518), .Z(n7733)
         );
  MUX2_X1 U26690 ( .A(n7733), .B(n7732), .S(n8346), .Z(n7734) );
  MUX2_X1 U26691 ( .A(n7734), .B(n7731), .S(n8231), .Z(n7735) );
  MUX2_X1 U26692 ( .A(\mem[438][7] ), .B(\mem[439][7] ), .S(n8518), .Z(n7736)
         );
  MUX2_X1 U26693 ( .A(\mem[436][7] ), .B(\mem[437][7] ), .S(n8518), .Z(n7737)
         );
  MUX2_X1 U26694 ( .A(n7737), .B(n7736), .S(n8346), .Z(n7738) );
  MUX2_X1 U26695 ( .A(\mem[434][7] ), .B(\mem[435][7] ), .S(n8518), .Z(n7739)
         );
  MUX2_X1 U26696 ( .A(\mem[432][7] ), .B(\mem[433][7] ), .S(n8518), .Z(n7740)
         );
  MUX2_X1 U26697 ( .A(n7740), .B(n7739), .S(n8346), .Z(n7741) );
  MUX2_X1 U26698 ( .A(n7741), .B(n7738), .S(n8227), .Z(n7742) );
  MUX2_X1 U26699 ( .A(n7742), .B(n7735), .S(n8216), .Z(n7743) );
  MUX2_X1 U26700 ( .A(\mem[430][7] ), .B(\mem[431][7] ), .S(n8519), .Z(n7744)
         );
  MUX2_X1 U26701 ( .A(\mem[428][7] ), .B(\mem[429][7] ), .S(n8519), .Z(n7745)
         );
  MUX2_X1 U26702 ( .A(n7745), .B(n7744), .S(n8347), .Z(n7746) );
  MUX2_X1 U26703 ( .A(\mem[426][7] ), .B(\mem[427][7] ), .S(n8519), .Z(n7747)
         );
  MUX2_X1 U26704 ( .A(\mem[424][7] ), .B(\mem[425][7] ), .S(n8519), .Z(n7748)
         );
  MUX2_X1 U26705 ( .A(n7748), .B(n7747), .S(n8347), .Z(n7749) );
  MUX2_X1 U26706 ( .A(n7749), .B(n7746), .S(n8227), .Z(n7750) );
  MUX2_X1 U26707 ( .A(\mem[422][7] ), .B(\mem[423][7] ), .S(n8519), .Z(n7751)
         );
  MUX2_X1 U26708 ( .A(\mem[420][7] ), .B(\mem[421][7] ), .S(n8519), .Z(n7752)
         );
  MUX2_X1 U26709 ( .A(n7752), .B(n7751), .S(n8347), .Z(n7753) );
  MUX2_X1 U26710 ( .A(\mem[418][7] ), .B(\mem[419][7] ), .S(n8519), .Z(n7754)
         );
  MUX2_X1 U26711 ( .A(\mem[416][7] ), .B(\mem[417][7] ), .S(n8519), .Z(n7755)
         );
  MUX2_X1 U26712 ( .A(n7755), .B(n7754), .S(n8347), .Z(n7756) );
  MUX2_X1 U26713 ( .A(n7756), .B(n7753), .S(n8262), .Z(n7757) );
  MUX2_X1 U26714 ( .A(n7757), .B(n7750), .S(n8216), .Z(n7758) );
  MUX2_X1 U26715 ( .A(n7758), .B(n7743), .S(n8193), .Z(n7759) );
  MUX2_X1 U26716 ( .A(\mem[414][7] ), .B(\mem[415][7] ), .S(n8519), .Z(n7760)
         );
  MUX2_X1 U26717 ( .A(\mem[412][7] ), .B(\mem[413][7] ), .S(n8519), .Z(n7761)
         );
  MUX2_X1 U26718 ( .A(n7761), .B(n7760), .S(n8347), .Z(n7762) );
  MUX2_X1 U26719 ( .A(\mem[410][7] ), .B(\mem[411][7] ), .S(n8519), .Z(n7763)
         );
  MUX2_X1 U26720 ( .A(\mem[408][7] ), .B(\mem[409][7] ), .S(n8519), .Z(n7764)
         );
  MUX2_X1 U26721 ( .A(n7764), .B(n7763), .S(n8347), .Z(n7765) );
  MUX2_X1 U26722 ( .A(n7765), .B(n7762), .S(n8257), .Z(n7766) );
  MUX2_X1 U26723 ( .A(\mem[406][7] ), .B(\mem[407][7] ), .S(n8520), .Z(n7767)
         );
  MUX2_X1 U26724 ( .A(\mem[404][7] ), .B(\mem[405][7] ), .S(n8520), .Z(n7768)
         );
  MUX2_X1 U26725 ( .A(n7768), .B(n7767), .S(n8347), .Z(n7769) );
  MUX2_X1 U26726 ( .A(\mem[402][7] ), .B(\mem[403][7] ), .S(n8520), .Z(n7770)
         );
  MUX2_X1 U26727 ( .A(\mem[400][7] ), .B(\mem[401][7] ), .S(n8520), .Z(n7771)
         );
  MUX2_X1 U26728 ( .A(n7771), .B(n7770), .S(n8347), .Z(n7772) );
  MUX2_X1 U26729 ( .A(n7772), .B(n7769), .S(n8226), .Z(n7773) );
  MUX2_X1 U26730 ( .A(n7773), .B(n7766), .S(n8216), .Z(n7774) );
  MUX2_X1 U26731 ( .A(\mem[398][7] ), .B(\mem[399][7] ), .S(n8520), .Z(n7775)
         );
  MUX2_X1 U26732 ( .A(\mem[396][7] ), .B(\mem[397][7] ), .S(n8520), .Z(n7776)
         );
  MUX2_X1 U26733 ( .A(n7776), .B(n7775), .S(n8347), .Z(n7777) );
  MUX2_X1 U26734 ( .A(\mem[394][7] ), .B(\mem[395][7] ), .S(n8520), .Z(n7778)
         );
  MUX2_X1 U26735 ( .A(\mem[392][7] ), .B(\mem[393][7] ), .S(n8520), .Z(n7779)
         );
  MUX2_X1 U26736 ( .A(n7779), .B(n7778), .S(n8347), .Z(n7780) );
  MUX2_X1 U26737 ( .A(n7780), .B(n7777), .S(n8241), .Z(n7781) );
  MUX2_X1 U26738 ( .A(\mem[390][7] ), .B(\mem[391][7] ), .S(n8520), .Z(n7782)
         );
  MUX2_X1 U26739 ( .A(\mem[388][7] ), .B(\mem[389][7] ), .S(n8520), .Z(n7783)
         );
  MUX2_X1 U26740 ( .A(n7783), .B(n7782), .S(n8347), .Z(n7784) );
  MUX2_X1 U26741 ( .A(\mem[386][7] ), .B(\mem[387][7] ), .S(n8520), .Z(n7785)
         );
  MUX2_X1 U26742 ( .A(\mem[384][7] ), .B(\mem[385][7] ), .S(n8520), .Z(n7786)
         );
  MUX2_X1 U26743 ( .A(n7786), .B(n7785), .S(n8347), .Z(n7787) );
  MUX2_X1 U26744 ( .A(n7787), .B(n7784), .S(n8242), .Z(n7788) );
  MUX2_X1 U26745 ( .A(n7788), .B(n7781), .S(n8216), .Z(n7789) );
  MUX2_X1 U26746 ( .A(n7789), .B(n7774), .S(n8193), .Z(n7790) );
  MUX2_X1 U26747 ( .A(n7790), .B(n7759), .S(n8181), .Z(n7791) );
  MUX2_X1 U26748 ( .A(n7791), .B(n7728), .S(n8180), .Z(n7792) );
  MUX2_X1 U26749 ( .A(\mem[382][7] ), .B(\mem[383][7] ), .S(n8521), .Z(n7793)
         );
  MUX2_X1 U26750 ( .A(\mem[380][7] ), .B(\mem[381][7] ), .S(n8521), .Z(n7794)
         );
  MUX2_X1 U26751 ( .A(n7794), .B(n7793), .S(n8348), .Z(n7795) );
  MUX2_X1 U26752 ( .A(\mem[378][7] ), .B(\mem[379][7] ), .S(n8521), .Z(n7796)
         );
  MUX2_X1 U26753 ( .A(\mem[376][7] ), .B(\mem[377][7] ), .S(n8521), .Z(n7797)
         );
  MUX2_X1 U26754 ( .A(n7797), .B(n7796), .S(n8348), .Z(n7798) );
  MUX2_X1 U26755 ( .A(n7798), .B(n7795), .S(n8248), .Z(n7799) );
  MUX2_X1 U26756 ( .A(\mem[374][7] ), .B(\mem[375][7] ), .S(n8521), .Z(n7800)
         );
  MUX2_X1 U26757 ( .A(\mem[372][7] ), .B(\mem[373][7] ), .S(n8521), .Z(n7801)
         );
  MUX2_X1 U26758 ( .A(n7801), .B(n7800), .S(n8348), .Z(n7802) );
  MUX2_X1 U26759 ( .A(\mem[370][7] ), .B(\mem[371][7] ), .S(n8521), .Z(n7803)
         );
  MUX2_X1 U26760 ( .A(\mem[368][7] ), .B(\mem[369][7] ), .S(n8521), .Z(n7804)
         );
  MUX2_X1 U26761 ( .A(n7804), .B(n7803), .S(n8348), .Z(n7805) );
  MUX2_X1 U26762 ( .A(n7805), .B(n7802), .S(n8249), .Z(n7806) );
  MUX2_X1 U26763 ( .A(n7806), .B(n7799), .S(n8217), .Z(n7807) );
  MUX2_X1 U26764 ( .A(\mem[366][7] ), .B(\mem[367][7] ), .S(n8521), .Z(n7808)
         );
  MUX2_X1 U26765 ( .A(\mem[364][7] ), .B(\mem[365][7] ), .S(n8521), .Z(n7809)
         );
  MUX2_X1 U26766 ( .A(n7809), .B(n7808), .S(n8348), .Z(n7810) );
  MUX2_X1 U26767 ( .A(\mem[362][7] ), .B(\mem[363][7] ), .S(n8521), .Z(n7811)
         );
  MUX2_X1 U26768 ( .A(\mem[360][7] ), .B(\mem[361][7] ), .S(n8521), .Z(n7812)
         );
  MUX2_X1 U26769 ( .A(n7812), .B(n7811), .S(n8348), .Z(n7813) );
  MUX2_X1 U26770 ( .A(n7813), .B(n7810), .S(n8244), .Z(n7814) );
  MUX2_X1 U26771 ( .A(\mem[358][7] ), .B(\mem[359][7] ), .S(n8522), .Z(n7815)
         );
  MUX2_X1 U26772 ( .A(\mem[356][7] ), .B(\mem[357][7] ), .S(n8522), .Z(n7816)
         );
  MUX2_X1 U26773 ( .A(n7816), .B(n7815), .S(n8348), .Z(n7817) );
  MUX2_X1 U26774 ( .A(\mem[354][7] ), .B(\mem[355][7] ), .S(n8522), .Z(n7818)
         );
  MUX2_X1 U26775 ( .A(\mem[352][7] ), .B(\mem[353][7] ), .S(n8522), .Z(n7819)
         );
  MUX2_X1 U26776 ( .A(n7819), .B(n7818), .S(n8348), .Z(n7820) );
  MUX2_X1 U26777 ( .A(n7820), .B(n7817), .S(n8245), .Z(n7821) );
  MUX2_X1 U26778 ( .A(n7821), .B(n7814), .S(n8217), .Z(n7822) );
  MUX2_X1 U26779 ( .A(n7822), .B(n7807), .S(n8194), .Z(n7823) );
  MUX2_X1 U26780 ( .A(\mem[350][7] ), .B(\mem[351][7] ), .S(n8522), .Z(n7824)
         );
  MUX2_X1 U26781 ( .A(\mem[348][7] ), .B(\mem[349][7] ), .S(n8522), .Z(n7825)
         );
  MUX2_X1 U26782 ( .A(n7825), .B(n7824), .S(n8348), .Z(n7826) );
  MUX2_X1 U26783 ( .A(\mem[346][7] ), .B(\mem[347][7] ), .S(n8522), .Z(n7827)
         );
  MUX2_X1 U26784 ( .A(\mem[344][7] ), .B(\mem[345][7] ), .S(n8522), .Z(n7828)
         );
  MUX2_X1 U26785 ( .A(n7828), .B(n7827), .S(n8348), .Z(n7829) );
  MUX2_X1 U26786 ( .A(n7829), .B(n7826), .S(n8246), .Z(n7830) );
  MUX2_X1 U26787 ( .A(\mem[342][7] ), .B(\mem[343][7] ), .S(n8522), .Z(n7831)
         );
  MUX2_X1 U26788 ( .A(\mem[340][7] ), .B(\mem[341][7] ), .S(n8522), .Z(n7832)
         );
  MUX2_X1 U26789 ( .A(n7832), .B(n7831), .S(n8348), .Z(n7833) );
  MUX2_X1 U26790 ( .A(\mem[338][7] ), .B(\mem[339][7] ), .S(n8522), .Z(n7834)
         );
  MUX2_X1 U26791 ( .A(\mem[336][7] ), .B(\mem[337][7] ), .S(n8522), .Z(n7835)
         );
  MUX2_X1 U26792 ( .A(n7835), .B(n7834), .S(n8348), .Z(n7836) );
  MUX2_X1 U26793 ( .A(n7836), .B(n7833), .S(n8253), .Z(n7837) );
  MUX2_X1 U26794 ( .A(n7837), .B(n7830), .S(n8217), .Z(n7838) );
  MUX2_X1 U26795 ( .A(\mem[334][7] ), .B(\mem[335][7] ), .S(n8523), .Z(n7839)
         );
  MUX2_X1 U26796 ( .A(\mem[332][7] ), .B(\mem[333][7] ), .S(n8523), .Z(n7840)
         );
  MUX2_X1 U26797 ( .A(n7840), .B(n7839), .S(n8349), .Z(n7841) );
  MUX2_X1 U26798 ( .A(\mem[330][7] ), .B(\mem[331][7] ), .S(n8523), .Z(n7842)
         );
  MUX2_X1 U26799 ( .A(\mem[328][7] ), .B(\mem[329][7] ), .S(n8523), .Z(n7843)
         );
  MUX2_X1 U26800 ( .A(n7843), .B(n7842), .S(n8349), .Z(n7844) );
  MUX2_X1 U26801 ( .A(n7844), .B(n7841), .S(n8254), .Z(n7845) );
  MUX2_X1 U26802 ( .A(\mem[326][7] ), .B(\mem[327][7] ), .S(n8523), .Z(n7846)
         );
  MUX2_X1 U26803 ( .A(\mem[324][7] ), .B(\mem[325][7] ), .S(n8523), .Z(n7847)
         );
  MUX2_X1 U26804 ( .A(n7847), .B(n7846), .S(n8349), .Z(n7848) );
  MUX2_X1 U26805 ( .A(\mem[322][7] ), .B(\mem[323][7] ), .S(n8523), .Z(n7849)
         );
  MUX2_X1 U26806 ( .A(\mem[320][7] ), .B(\mem[321][7] ), .S(n8523), .Z(n7850)
         );
  MUX2_X1 U26807 ( .A(n7850), .B(n7849), .S(n8349), .Z(n7851) );
  MUX2_X1 U26808 ( .A(n7851), .B(n7848), .S(n8255), .Z(n7852) );
  MUX2_X1 U26809 ( .A(n7852), .B(n7845), .S(n8217), .Z(n7853) );
  MUX2_X1 U26810 ( .A(n7853), .B(n7838), .S(n8194), .Z(n7854) );
  MUX2_X1 U26811 ( .A(n7854), .B(n7823), .S(n8181), .Z(n7855) );
  MUX2_X1 U26812 ( .A(\mem[318][7] ), .B(\mem[319][7] ), .S(n8523), .Z(n7856)
         );
  MUX2_X1 U26813 ( .A(\mem[316][7] ), .B(\mem[317][7] ), .S(n8523), .Z(n7857)
         );
  MUX2_X1 U26814 ( .A(n7857), .B(n7856), .S(n8349), .Z(n7858) );
  MUX2_X1 U26815 ( .A(\mem[314][7] ), .B(\mem[315][7] ), .S(n8523), .Z(n7859)
         );
  MUX2_X1 U26816 ( .A(\mem[312][7] ), .B(\mem[313][7] ), .S(n8523), .Z(n7860)
         );
  MUX2_X1 U26817 ( .A(n7860), .B(n7859), .S(n8349), .Z(n7861) );
  MUX2_X1 U26818 ( .A(n7861), .B(n7858), .S(n8250), .Z(n7862) );
  MUX2_X1 U26819 ( .A(\mem[310][7] ), .B(\mem[311][7] ), .S(n8524), .Z(n7863)
         );
  MUX2_X1 U26820 ( .A(\mem[308][7] ), .B(\mem[309][7] ), .S(n8524), .Z(n7864)
         );
  MUX2_X1 U26821 ( .A(n7864), .B(n7863), .S(n8349), .Z(n7865) );
  MUX2_X1 U26822 ( .A(\mem[306][7] ), .B(\mem[307][7] ), .S(n8524), .Z(n7866)
         );
  MUX2_X1 U26823 ( .A(\mem[304][7] ), .B(\mem[305][7] ), .S(n8524), .Z(n7867)
         );
  MUX2_X1 U26824 ( .A(n7867), .B(n7866), .S(n8349), .Z(n7868) );
  MUX2_X1 U26825 ( .A(n7868), .B(n7865), .S(n8251), .Z(n7869) );
  MUX2_X1 U26826 ( .A(n7869), .B(n7862), .S(n8217), .Z(n7870) );
  MUX2_X1 U26827 ( .A(\mem[302][7] ), .B(\mem[303][7] ), .S(n8524), .Z(n7871)
         );
  MUX2_X1 U26828 ( .A(\mem[300][7] ), .B(\mem[301][7] ), .S(n8524), .Z(n7872)
         );
  MUX2_X1 U26829 ( .A(n7872), .B(n7871), .S(n8349), .Z(n7873) );
  MUX2_X1 U26830 ( .A(\mem[298][7] ), .B(\mem[299][7] ), .S(n8524), .Z(n7874)
         );
  MUX2_X1 U26831 ( .A(\mem[296][7] ), .B(\mem[297][7] ), .S(n8524), .Z(n7875)
         );
  MUX2_X1 U26832 ( .A(n7875), .B(n7874), .S(n8349), .Z(n7876) );
  MUX2_X1 U26833 ( .A(n7876), .B(n7873), .S(n8252), .Z(n7877) );
  MUX2_X1 U26834 ( .A(\mem[294][7] ), .B(\mem[295][7] ), .S(n8524), .Z(n7878)
         );
  MUX2_X1 U26835 ( .A(\mem[292][7] ), .B(\mem[293][7] ), .S(n8524), .Z(n7879)
         );
  MUX2_X1 U26836 ( .A(n7879), .B(n7878), .S(n8349), .Z(n7880) );
  MUX2_X1 U26837 ( .A(\mem[290][7] ), .B(\mem[291][7] ), .S(n8524), .Z(n7881)
         );
  MUX2_X1 U26838 ( .A(\mem[288][7] ), .B(\mem[289][7] ), .S(n8524), .Z(n7882)
         );
  MUX2_X1 U26839 ( .A(n7882), .B(n7881), .S(n8349), .Z(n7883) );
  MUX2_X1 U26840 ( .A(n7883), .B(n7880), .S(n8259), .Z(n7884) );
  MUX2_X1 U26841 ( .A(n7884), .B(n7877), .S(n8217), .Z(n7885) );
  MUX2_X1 U26842 ( .A(n7885), .B(n7870), .S(n8194), .Z(n7886) );
  MUX2_X1 U26843 ( .A(\mem[286][7] ), .B(\mem[287][7] ), .S(n8525), .Z(n7887)
         );
  MUX2_X1 U26844 ( .A(\mem[284][7] ), .B(\mem[285][7] ), .S(n8525), .Z(n7888)
         );
  MUX2_X1 U26845 ( .A(n7888), .B(n7887), .S(n8350), .Z(n7889) );
  MUX2_X1 U26846 ( .A(\mem[282][7] ), .B(\mem[283][7] ), .S(n8525), .Z(n7890)
         );
  MUX2_X1 U26847 ( .A(\mem[280][7] ), .B(\mem[281][7] ), .S(n8525), .Z(n7891)
         );
  MUX2_X1 U26848 ( .A(n7891), .B(n7890), .S(n8350), .Z(n7892) );
  MUX2_X1 U26849 ( .A(n7892), .B(n7889), .S(n8239), .Z(n7893) );
  MUX2_X1 U26850 ( .A(\mem[278][7] ), .B(\mem[279][7] ), .S(n8525), .Z(n7894)
         );
  MUX2_X1 U26851 ( .A(\mem[276][7] ), .B(\mem[277][7] ), .S(n8525), .Z(n7895)
         );
  MUX2_X1 U26852 ( .A(n7895), .B(n7894), .S(n8350), .Z(n7896) );
  MUX2_X1 U26853 ( .A(\mem[274][7] ), .B(\mem[275][7] ), .S(n8525), .Z(n7897)
         );
  MUX2_X1 U26854 ( .A(\mem[272][7] ), .B(\mem[273][7] ), .S(n8525), .Z(n7898)
         );
  MUX2_X1 U26855 ( .A(n7898), .B(n7897), .S(n8350), .Z(n7899) );
  MUX2_X1 U26856 ( .A(n7899), .B(n7896), .S(n8240), .Z(n7900) );
  MUX2_X1 U26857 ( .A(n7900), .B(n7893), .S(n8217), .Z(n7901) );
  MUX2_X1 U26858 ( .A(\mem[270][7] ), .B(\mem[271][7] ), .S(n8525), .Z(n7902)
         );
  MUX2_X1 U26859 ( .A(\mem[268][7] ), .B(\mem[269][7] ), .S(n8525), .Z(n7903)
         );
  MUX2_X1 U26860 ( .A(n7903), .B(n7902), .S(n8350), .Z(n7904) );
  MUX2_X1 U26861 ( .A(\mem[266][7] ), .B(\mem[267][7] ), .S(n8525), .Z(n7905)
         );
  MUX2_X1 U26862 ( .A(\mem[264][7] ), .B(\mem[265][7] ), .S(n8525), .Z(n7906)
         );
  MUX2_X1 U26863 ( .A(n7906), .B(n7905), .S(n8350), .Z(n7907) );
  MUX2_X1 U26864 ( .A(n7907), .B(n7904), .S(N20), .Z(n7908) );
  MUX2_X1 U26865 ( .A(\mem[262][7] ), .B(\mem[263][7] ), .S(n8526), .Z(n7909)
         );
  MUX2_X1 U26866 ( .A(\mem[260][7] ), .B(\mem[261][7] ), .S(n8526), .Z(n7910)
         );
  MUX2_X1 U26867 ( .A(n7910), .B(n7909), .S(n8350), .Z(n7911) );
  MUX2_X1 U26868 ( .A(\mem[258][7] ), .B(\mem[259][7] ), .S(n8526), .Z(n7912)
         );
  MUX2_X1 U26869 ( .A(\mem[256][7] ), .B(\mem[257][7] ), .S(n8526), .Z(n7913)
         );
  MUX2_X1 U26870 ( .A(n7913), .B(n7912), .S(n8350), .Z(n7914) );
  MUX2_X1 U26871 ( .A(n7914), .B(n7911), .S(n8263), .Z(n7915) );
  MUX2_X1 U26872 ( .A(n7915), .B(n7908), .S(n8217), .Z(n7916) );
  MUX2_X1 U26873 ( .A(n7916), .B(n7901), .S(n8194), .Z(n7917) );
  MUX2_X1 U26874 ( .A(n7917), .B(n7886), .S(n8182), .Z(n7918) );
  MUX2_X1 U26875 ( .A(n7918), .B(n7855), .S(n8180), .Z(n7919) );
  MUX2_X1 U26876 ( .A(n7919), .B(n7792), .S(N25), .Z(n7920) );
  MUX2_X1 U26877 ( .A(\mem[254][7] ), .B(\mem[255][7] ), .S(n8526), .Z(n7921)
         );
  MUX2_X1 U26878 ( .A(\mem[252][7] ), .B(\mem[253][7] ), .S(n8526), .Z(n7922)
         );
  MUX2_X1 U26879 ( .A(n7922), .B(n7921), .S(n8350), .Z(n7923) );
  MUX2_X1 U26880 ( .A(\mem[250][7] ), .B(\mem[251][7] ), .S(n8526), .Z(n7924)
         );
  MUX2_X1 U26881 ( .A(\mem[248][7] ), .B(\mem[249][7] ), .S(n8526), .Z(n7925)
         );
  MUX2_X1 U26882 ( .A(n7925), .B(n7924), .S(n8350), .Z(n7926) );
  MUX2_X1 U26883 ( .A(n7926), .B(n7923), .S(n8228), .Z(n7927) );
  MUX2_X1 U26884 ( .A(\mem[246][7] ), .B(\mem[247][7] ), .S(n8526), .Z(n7928)
         );
  MUX2_X1 U26885 ( .A(\mem[244][7] ), .B(\mem[245][7] ), .S(n8526), .Z(n7929)
         );
  MUX2_X1 U26886 ( .A(n7929), .B(n7928), .S(n8350), .Z(n7930) );
  MUX2_X1 U26887 ( .A(\mem[242][7] ), .B(\mem[243][7] ), .S(n8526), .Z(n7931)
         );
  MUX2_X1 U26888 ( .A(\mem[240][7] ), .B(\mem[241][7] ), .S(n8526), .Z(n7932)
         );
  MUX2_X1 U26889 ( .A(n7932), .B(n7931), .S(n8350), .Z(n7933) );
  MUX2_X1 U26890 ( .A(n7933), .B(n7930), .S(n8248), .Z(n7934) );
  MUX2_X1 U26891 ( .A(n7934), .B(n7927), .S(n8217), .Z(n7935) );
  MUX2_X1 U26892 ( .A(\mem[238][7] ), .B(\mem[239][7] ), .S(n8527), .Z(n7936)
         );
  MUX2_X1 U26893 ( .A(\mem[236][7] ), .B(\mem[237][7] ), .S(n8527), .Z(n7937)
         );
  MUX2_X1 U26894 ( .A(n7937), .B(n7936), .S(n8351), .Z(n7938) );
  MUX2_X1 U26895 ( .A(\mem[234][7] ), .B(\mem[235][7] ), .S(n8527), .Z(n7939)
         );
  MUX2_X1 U26896 ( .A(\mem[232][7] ), .B(\mem[233][7] ), .S(n8527), .Z(n7940)
         );
  MUX2_X1 U26897 ( .A(n7940), .B(n7939), .S(n8351), .Z(n7941) );
  MUX2_X1 U26898 ( .A(n7941), .B(n7938), .S(n8223), .Z(n7942) );
  MUX2_X1 U26899 ( .A(\mem[230][7] ), .B(\mem[231][7] ), .S(n8527), .Z(n7943)
         );
  MUX2_X1 U26900 ( .A(\mem[228][7] ), .B(\mem[229][7] ), .S(n8527), .Z(n7944)
         );
  MUX2_X1 U26901 ( .A(n7944), .B(n7943), .S(n8351), .Z(n7945) );
  MUX2_X1 U26902 ( .A(\mem[226][7] ), .B(\mem[227][7] ), .S(n8527), .Z(n7946)
         );
  MUX2_X1 U26903 ( .A(\mem[224][7] ), .B(\mem[225][7] ), .S(n8527), .Z(n7947)
         );
  MUX2_X1 U26904 ( .A(n7947), .B(n7946), .S(n8351), .Z(n7948) );
  MUX2_X1 U26905 ( .A(n7948), .B(n7945), .S(n8228), .Z(n7949) );
  MUX2_X1 U26906 ( .A(n7949), .B(n7942), .S(n8217), .Z(n7950) );
  MUX2_X1 U26907 ( .A(n7950), .B(n7935), .S(n8194), .Z(n7951) );
  MUX2_X1 U26908 ( .A(\mem[222][7] ), .B(\mem[223][7] ), .S(n8527), .Z(n7952)
         );
  MUX2_X1 U26909 ( .A(\mem[220][7] ), .B(\mem[221][7] ), .S(n8527), .Z(n7953)
         );
  MUX2_X1 U26910 ( .A(n7953), .B(n7952), .S(n8351), .Z(n7954) );
  MUX2_X1 U26911 ( .A(\mem[218][7] ), .B(\mem[219][7] ), .S(n8527), .Z(n7955)
         );
  MUX2_X1 U26912 ( .A(\mem[216][7] ), .B(\mem[217][7] ), .S(n8527), .Z(n7956)
         );
  MUX2_X1 U26913 ( .A(n7956), .B(n7955), .S(n8351), .Z(n7957) );
  MUX2_X1 U26914 ( .A(n7957), .B(n7954), .S(n8229), .Z(n7958) );
  MUX2_X1 U26915 ( .A(\mem[214][7] ), .B(\mem[215][7] ), .S(n8528), .Z(n7959)
         );
  MUX2_X1 U26916 ( .A(\mem[212][7] ), .B(\mem[213][7] ), .S(n8528), .Z(n7960)
         );
  MUX2_X1 U26917 ( .A(n7960), .B(n7959), .S(n8351), .Z(n7961) );
  MUX2_X1 U26918 ( .A(\mem[210][7] ), .B(\mem[211][7] ), .S(n8528), .Z(n7962)
         );
  MUX2_X1 U26919 ( .A(\mem[208][7] ), .B(\mem[209][7] ), .S(n8528), .Z(n7963)
         );
  MUX2_X1 U26920 ( .A(n7963), .B(n7962), .S(n8351), .Z(n7964) );
  MUX2_X1 U26921 ( .A(n7964), .B(n7961), .S(n8225), .Z(n7965) );
  MUX2_X1 U26922 ( .A(n7965), .B(n7958), .S(n8217), .Z(n7966) );
  MUX2_X1 U26923 ( .A(\mem[206][7] ), .B(\mem[207][7] ), .S(n8528), .Z(n7967)
         );
  MUX2_X1 U26924 ( .A(\mem[204][7] ), .B(\mem[205][7] ), .S(n8528), .Z(n7968)
         );
  MUX2_X1 U26925 ( .A(n7968), .B(n7967), .S(n8351), .Z(n7969) );
  MUX2_X1 U26926 ( .A(\mem[202][7] ), .B(\mem[203][7] ), .S(n8528), .Z(n7970)
         );
  MUX2_X1 U26927 ( .A(\mem[200][7] ), .B(\mem[201][7] ), .S(n8528), .Z(n7971)
         );
  MUX2_X1 U26928 ( .A(n7971), .B(n7970), .S(n8351), .Z(n7972) );
  MUX2_X1 U26929 ( .A(n7972), .B(n7969), .S(n8220), .Z(n7973) );
  MUX2_X1 U26930 ( .A(\mem[198][7] ), .B(\mem[199][7] ), .S(n8528), .Z(n7974)
         );
  MUX2_X1 U26931 ( .A(\mem[196][7] ), .B(\mem[197][7] ), .S(n8528), .Z(n7975)
         );
  MUX2_X1 U26932 ( .A(n7975), .B(n7974), .S(n8351), .Z(n7976) );
  MUX2_X1 U26933 ( .A(\mem[194][7] ), .B(\mem[195][7] ), .S(n8528), .Z(n7977)
         );
  MUX2_X1 U26934 ( .A(\mem[192][7] ), .B(\mem[193][7] ), .S(n8528), .Z(n7978)
         );
  MUX2_X1 U26935 ( .A(n7978), .B(n7977), .S(n8351), .Z(n7979) );
  MUX2_X1 U26936 ( .A(n7979), .B(n7976), .S(n8221), .Z(n7980) );
  MUX2_X1 U26937 ( .A(n7980), .B(n7973), .S(n8217), .Z(n7981) );
  MUX2_X1 U26938 ( .A(n7981), .B(n7966), .S(n8194), .Z(n7982) );
  MUX2_X1 U26939 ( .A(n7982), .B(n7951), .S(n8183), .Z(n7983) );
  MUX2_X1 U26940 ( .A(\mem[190][7] ), .B(\mem[191][7] ), .S(n8529), .Z(n7984)
         );
  MUX2_X1 U26941 ( .A(\mem[188][7] ), .B(\mem[189][7] ), .S(n8529), .Z(n7985)
         );
  MUX2_X1 U26942 ( .A(n7985), .B(n7984), .S(n8352), .Z(n7986) );
  MUX2_X1 U26943 ( .A(\mem[186][7] ), .B(\mem[187][7] ), .S(n8529), .Z(n7987)
         );
  MUX2_X1 U26944 ( .A(\mem[184][7] ), .B(\mem[185][7] ), .S(n8529), .Z(n7988)
         );
  MUX2_X1 U26945 ( .A(n7988), .B(n7987), .S(n8352), .Z(n7989) );
  MUX2_X1 U26946 ( .A(n7989), .B(n7986), .S(n8260), .Z(n7990) );
  MUX2_X1 U26947 ( .A(\mem[182][7] ), .B(\mem[183][7] ), .S(n8529), .Z(n7991)
         );
  MUX2_X1 U26948 ( .A(\mem[180][7] ), .B(\mem[181][7] ), .S(n8529), .Z(n7992)
         );
  MUX2_X1 U26949 ( .A(n7992), .B(n7991), .S(n8352), .Z(n7993) );
  MUX2_X1 U26950 ( .A(\mem[178][7] ), .B(\mem[179][7] ), .S(n8529), .Z(n7994)
         );
  MUX2_X1 U26951 ( .A(\mem[176][7] ), .B(\mem[177][7] ), .S(n8529), .Z(n7995)
         );
  MUX2_X1 U26952 ( .A(n7995), .B(n7994), .S(n8352), .Z(n7996) );
  MUX2_X1 U26953 ( .A(n7996), .B(n7993), .S(n8261), .Z(n7997) );
  MUX2_X1 U26954 ( .A(n7997), .B(n7990), .S(n8218), .Z(n7998) );
  MUX2_X1 U26955 ( .A(\mem[174][7] ), .B(\mem[175][7] ), .S(n8529), .Z(n7999)
         );
  MUX2_X1 U26956 ( .A(\mem[172][7] ), .B(\mem[173][7] ), .S(n8529), .Z(n8000)
         );
  MUX2_X1 U26957 ( .A(n8000), .B(n7999), .S(n8352), .Z(n8001) );
  MUX2_X1 U26958 ( .A(\mem[170][7] ), .B(\mem[171][7] ), .S(n8529), .Z(n8002)
         );
  MUX2_X1 U26959 ( .A(\mem[168][7] ), .B(\mem[169][7] ), .S(n8529), .Z(n8003)
         );
  MUX2_X1 U26960 ( .A(n8003), .B(n8002), .S(n8352), .Z(n8004) );
  MUX2_X1 U26961 ( .A(n8004), .B(n8001), .S(n8256), .Z(n8005) );
  MUX2_X1 U26962 ( .A(\mem[166][7] ), .B(\mem[167][7] ), .S(n8530), .Z(n8006)
         );
  MUX2_X1 U26963 ( .A(\mem[164][7] ), .B(\mem[165][7] ), .S(n8530), .Z(n8007)
         );
  MUX2_X1 U26964 ( .A(n8007), .B(n8006), .S(n8352), .Z(n8008) );
  MUX2_X1 U26965 ( .A(\mem[162][7] ), .B(\mem[163][7] ), .S(n8530), .Z(n8009)
         );
  MUX2_X1 U26966 ( .A(\mem[160][7] ), .B(\mem[161][7] ), .S(n8530), .Z(n8010)
         );
  MUX2_X1 U26967 ( .A(n8010), .B(n8009), .S(n8352), .Z(n8011) );
  MUX2_X1 U26968 ( .A(n8011), .B(n8008), .S(n8257), .Z(n8012) );
  MUX2_X1 U26969 ( .A(n8012), .B(n8005), .S(n8218), .Z(n8013) );
  MUX2_X1 U26970 ( .A(n8013), .B(n7998), .S(n8194), .Z(n8014) );
  MUX2_X1 U26971 ( .A(\mem[158][7] ), .B(\mem[159][7] ), .S(n8530), .Z(n8015)
         );
  MUX2_X1 U26972 ( .A(\mem[156][7] ), .B(\mem[157][7] ), .S(n8530), .Z(n8016)
         );
  MUX2_X1 U26973 ( .A(n8016), .B(n8015), .S(n8352), .Z(n8017) );
  MUX2_X1 U26974 ( .A(\mem[154][7] ), .B(\mem[155][7] ), .S(n8530), .Z(n8018)
         );
  MUX2_X1 U26975 ( .A(\mem[152][7] ), .B(\mem[153][7] ), .S(n8530), .Z(n8019)
         );
  MUX2_X1 U26976 ( .A(n8019), .B(n8018), .S(n8352), .Z(n8020) );
  MUX2_X1 U26977 ( .A(n8020), .B(n8017), .S(n8258), .Z(n8021) );
  MUX2_X1 U26978 ( .A(\mem[150][7] ), .B(\mem[151][7] ), .S(n8530), .Z(n8022)
         );
  MUX2_X1 U26979 ( .A(\mem[148][7] ), .B(\mem[149][7] ), .S(n8530), .Z(n8023)
         );
  MUX2_X1 U26980 ( .A(n8023), .B(n8022), .S(n8352), .Z(n8024) );
  MUX2_X1 U26981 ( .A(\mem[146][7] ), .B(\mem[147][7] ), .S(n8530), .Z(n8025)
         );
  MUX2_X1 U26982 ( .A(\mem[144][7] ), .B(\mem[145][7] ), .S(n8530), .Z(n8026)
         );
  MUX2_X1 U26983 ( .A(n8026), .B(n8025), .S(n8352), .Z(n8027) );
  MUX2_X1 U26984 ( .A(n8027), .B(n8024), .S(n8235), .Z(n8028) );
  MUX2_X1 U26985 ( .A(n8028), .B(n8021), .S(n8218), .Z(n8029) );
  MUX2_X1 U26986 ( .A(\mem[142][7] ), .B(\mem[143][7] ), .S(n8531), .Z(n8030)
         );
  MUX2_X1 U26987 ( .A(\mem[140][7] ), .B(\mem[141][7] ), .S(n8531), .Z(n8031)
         );
  MUX2_X1 U26988 ( .A(n8031), .B(n8030), .S(n8353), .Z(n8032) );
  MUX2_X1 U26989 ( .A(\mem[138][7] ), .B(\mem[139][7] ), .S(n8531), .Z(n8033)
         );
  MUX2_X1 U26990 ( .A(\mem[136][7] ), .B(\mem[137][7] ), .S(n8531), .Z(n8034)
         );
  MUX2_X1 U26991 ( .A(n8034), .B(n8033), .S(n8353), .Z(n8035) );
  MUX2_X1 U26992 ( .A(n8035), .B(n8032), .S(n8236), .Z(n8036) );
  MUX2_X1 U26993 ( .A(\mem[134][7] ), .B(\mem[135][7] ), .S(n8531), .Z(n8037)
         );
  MUX2_X1 U26994 ( .A(\mem[132][7] ), .B(\mem[133][7] ), .S(n8531), .Z(n8038)
         );
  MUX2_X1 U26995 ( .A(n8038), .B(n8037), .S(n8353), .Z(n8039) );
  MUX2_X1 U26996 ( .A(\mem[130][7] ), .B(\mem[131][7] ), .S(n8531), .Z(n8040)
         );
  MUX2_X1 U26997 ( .A(\mem[128][7] ), .B(\mem[129][7] ), .S(n8531), .Z(n8041)
         );
  MUX2_X1 U26998 ( .A(n8041), .B(n8040), .S(n8353), .Z(n8042) );
  MUX2_X1 U26999 ( .A(n8042), .B(n8039), .S(n8237), .Z(n8043) );
  MUX2_X1 U27000 ( .A(n8043), .B(n8036), .S(n8218), .Z(n8044) );
  MUX2_X1 U27001 ( .A(n8044), .B(n8029), .S(n8194), .Z(n8045) );
  MUX2_X1 U27002 ( .A(n8045), .B(n8014), .S(n8184), .Z(n8046) );
  MUX2_X1 U27003 ( .A(n8046), .B(n7983), .S(n8180), .Z(n8047) );
  MUX2_X1 U27004 ( .A(\mem[126][7] ), .B(\mem[127][7] ), .S(n8531), .Z(n8048)
         );
  MUX2_X1 U27005 ( .A(\mem[124][7] ), .B(\mem[125][7] ), .S(n8531), .Z(n8049)
         );
  MUX2_X1 U27006 ( .A(n8049), .B(n8048), .S(n8353), .Z(n8050) );
  MUX2_X1 U27007 ( .A(\mem[122][7] ), .B(\mem[123][7] ), .S(n8531), .Z(n8051)
         );
  MUX2_X1 U27008 ( .A(\mem[120][7] ), .B(\mem[121][7] ), .S(n8531), .Z(n8052)
         );
  MUX2_X1 U27009 ( .A(n8052), .B(n8051), .S(n8353), .Z(n8053) );
  MUX2_X1 U27010 ( .A(n8053), .B(n8050), .S(n8232), .Z(n8054) );
  MUX2_X1 U27011 ( .A(\mem[118][7] ), .B(\mem[119][7] ), .S(n8532), .Z(n8055)
         );
  MUX2_X1 U27012 ( .A(\mem[116][7] ), .B(\mem[117][7] ), .S(n8532), .Z(n8056)
         );
  MUX2_X1 U27013 ( .A(n8056), .B(n8055), .S(n8353), .Z(n8057) );
  MUX2_X1 U27014 ( .A(\mem[114][7] ), .B(\mem[115][7] ), .S(n8532), .Z(n8058)
         );
  MUX2_X1 U27015 ( .A(\mem[112][7] ), .B(\mem[113][7] ), .S(n8532), .Z(n8059)
         );
  MUX2_X1 U27016 ( .A(n8059), .B(n8058), .S(n8353), .Z(n8060) );
  MUX2_X1 U27017 ( .A(n8060), .B(n8057), .S(n8233), .Z(n8061) );
  MUX2_X1 U27018 ( .A(n8061), .B(n8054), .S(n8218), .Z(n8062) );
  MUX2_X1 U27019 ( .A(\mem[110][7] ), .B(\mem[111][7] ), .S(n8532), .Z(n8063)
         );
  MUX2_X1 U27020 ( .A(\mem[108][7] ), .B(\mem[109][7] ), .S(n8532), .Z(n8064)
         );
  MUX2_X1 U27021 ( .A(n8064), .B(n8063), .S(n8353), .Z(n8065) );
  MUX2_X1 U27022 ( .A(\mem[106][7] ), .B(\mem[107][7] ), .S(n8532), .Z(n8066)
         );
  MUX2_X1 U27023 ( .A(\mem[104][7] ), .B(\mem[105][7] ), .S(n8532), .Z(n8067)
         );
  MUX2_X1 U27024 ( .A(n8067), .B(n8066), .S(n8353), .Z(n8068) );
  MUX2_X1 U27025 ( .A(n8068), .B(n8065), .S(n8234), .Z(n8069) );
  MUX2_X1 U27026 ( .A(\mem[102][7] ), .B(\mem[103][7] ), .S(n8532), .Z(n8070)
         );
  MUX2_X1 U27027 ( .A(\mem[100][7] ), .B(\mem[101][7] ), .S(n8532), .Z(n8071)
         );
  MUX2_X1 U27028 ( .A(n8071), .B(n8070), .S(n8353), .Z(n8072) );
  MUX2_X1 U27029 ( .A(\mem[98][7] ), .B(\mem[99][7] ), .S(n8532), .Z(n8073) );
  MUX2_X1 U27030 ( .A(\mem[96][7] ), .B(\mem[97][7] ), .S(n8532), .Z(n8074) );
  MUX2_X1 U27031 ( .A(n8074), .B(n8073), .S(n8353), .Z(n8075) );
  MUX2_X1 U27032 ( .A(n8075), .B(n8072), .S(n8230), .Z(n8076) );
  MUX2_X1 U27033 ( .A(n8076), .B(n8069), .S(n8218), .Z(n8077) );
  MUX2_X1 U27034 ( .A(n8077), .B(n8062), .S(n8194), .Z(n8078) );
  MUX2_X1 U27035 ( .A(\mem[94][7] ), .B(\mem[95][7] ), .S(n8533), .Z(n8079) );
  MUX2_X1 U27036 ( .A(\mem[92][7] ), .B(\mem[93][7] ), .S(n8533), .Z(n8080) );
  MUX2_X1 U27037 ( .A(n8080), .B(n8079), .S(n8354), .Z(n8081) );
  MUX2_X1 U27038 ( .A(\mem[90][7] ), .B(\mem[91][7] ), .S(n8533), .Z(n8082) );
  MUX2_X1 U27039 ( .A(\mem[88][7] ), .B(\mem[89][7] ), .S(n8533), .Z(n8083) );
  MUX2_X1 U27040 ( .A(n8083), .B(n8082), .S(n8354), .Z(n8084) );
  MUX2_X1 U27041 ( .A(n8084), .B(n8081), .S(n8262), .Z(n8085) );
  MUX2_X1 U27042 ( .A(\mem[86][7] ), .B(\mem[87][7] ), .S(n8533), .Z(n8086) );
  MUX2_X1 U27043 ( .A(\mem[84][7] ), .B(\mem[85][7] ), .S(n8533), .Z(n8087) );
  MUX2_X1 U27044 ( .A(n8087), .B(n8086), .S(n8354), .Z(n8088) );
  MUX2_X1 U27045 ( .A(\mem[82][7] ), .B(\mem[83][7] ), .S(n8533), .Z(n8089) );
  MUX2_X1 U27046 ( .A(\mem[80][7] ), .B(\mem[81][7] ), .S(n8533), .Z(n8090) );
  MUX2_X1 U27047 ( .A(n8090), .B(n8089), .S(n8354), .Z(n8091) );
  MUX2_X1 U27048 ( .A(n8091), .B(n8088), .S(n8262), .Z(n8092) );
  MUX2_X1 U27049 ( .A(n8092), .B(n8085), .S(n8218), .Z(n8093) );
  MUX2_X1 U27050 ( .A(\mem[78][7] ), .B(\mem[79][7] ), .S(n8533), .Z(n8094) );
  MUX2_X1 U27051 ( .A(\mem[76][7] ), .B(\mem[77][7] ), .S(n8533), .Z(n8095) );
  MUX2_X1 U27052 ( .A(n8095), .B(n8094), .S(n8354), .Z(n8096) );
  MUX2_X1 U27053 ( .A(\mem[74][7] ), .B(\mem[75][7] ), .S(n8533), .Z(n8097) );
  MUX2_X1 U27054 ( .A(\mem[72][7] ), .B(\mem[73][7] ), .S(n8533), .Z(n8098) );
  MUX2_X1 U27055 ( .A(n8098), .B(n8097), .S(n8354), .Z(n8099) );
  MUX2_X1 U27056 ( .A(n8099), .B(n8096), .S(n8262), .Z(n8100) );
  MUX2_X1 U27057 ( .A(\mem[70][7] ), .B(\mem[71][7] ), .S(n8534), .Z(n8101) );
  MUX2_X1 U27058 ( .A(\mem[68][7] ), .B(\mem[69][7] ), .S(n8534), .Z(n8102) );
  MUX2_X1 U27059 ( .A(n8102), .B(n8101), .S(n8354), .Z(n8103) );
  MUX2_X1 U27060 ( .A(\mem[66][7] ), .B(\mem[67][7] ), .S(n8534), .Z(n8104) );
  MUX2_X1 U27061 ( .A(\mem[64][7] ), .B(\mem[65][7] ), .S(n8534), .Z(n8105) );
  MUX2_X1 U27062 ( .A(n8105), .B(n8104), .S(n8354), .Z(n8106) );
  MUX2_X1 U27063 ( .A(n8106), .B(n8103), .S(n8262), .Z(n8107) );
  MUX2_X1 U27064 ( .A(n8107), .B(n8100), .S(n8218), .Z(n8108) );
  MUX2_X1 U27065 ( .A(n8108), .B(n8093), .S(n8194), .Z(n8109) );
  MUX2_X1 U27066 ( .A(n8109), .B(n8078), .S(n8182), .Z(n8110) );
  MUX2_X1 U27067 ( .A(\mem[62][7] ), .B(\mem[63][7] ), .S(n8534), .Z(n8111) );
  MUX2_X1 U27068 ( .A(\mem[60][7] ), .B(\mem[61][7] ), .S(n8534), .Z(n8112) );
  MUX2_X1 U27069 ( .A(n8112), .B(n8111), .S(n8354), .Z(n8113) );
  MUX2_X1 U27070 ( .A(\mem[58][7] ), .B(\mem[59][7] ), .S(n8534), .Z(n8114) );
  MUX2_X1 U27071 ( .A(\mem[56][7] ), .B(\mem[57][7] ), .S(n8534), .Z(n8115) );
  MUX2_X1 U27072 ( .A(n8115), .B(n8114), .S(n8354), .Z(n8116) );
  MUX2_X1 U27073 ( .A(n8116), .B(n8113), .S(n8262), .Z(n8117) );
  MUX2_X1 U27074 ( .A(\mem[54][7] ), .B(\mem[55][7] ), .S(n8534), .Z(n8118) );
  MUX2_X1 U27075 ( .A(\mem[52][7] ), .B(\mem[53][7] ), .S(n8534), .Z(n8119) );
  MUX2_X1 U27076 ( .A(n8119), .B(n8118), .S(n8354), .Z(n8120) );
  MUX2_X1 U27077 ( .A(\mem[50][7] ), .B(\mem[51][7] ), .S(n8534), .Z(n8121) );
  MUX2_X1 U27078 ( .A(\mem[48][7] ), .B(\mem[49][7] ), .S(n8534), .Z(n8122) );
  MUX2_X1 U27079 ( .A(n8122), .B(n8121), .S(n8354), .Z(n8123) );
  MUX2_X1 U27080 ( .A(n8123), .B(n8120), .S(n8262), .Z(n8124) );
  MUX2_X1 U27081 ( .A(n8124), .B(n8117), .S(n8218), .Z(n8125) );
  MUX2_X1 U27082 ( .A(\mem[46][7] ), .B(\mem[47][7] ), .S(n8535), .Z(n8126) );
  MUX2_X1 U27083 ( .A(\mem[44][7] ), .B(\mem[45][7] ), .S(n8535), .Z(n8127) );
  MUX2_X1 U27084 ( .A(n8127), .B(n8126), .S(n8355), .Z(n8128) );
  MUX2_X1 U27085 ( .A(\mem[42][7] ), .B(\mem[43][7] ), .S(n8535), .Z(n8129) );
  MUX2_X1 U27086 ( .A(\mem[40][7] ), .B(\mem[41][7] ), .S(n8535), .Z(n8130) );
  MUX2_X1 U27087 ( .A(n8130), .B(n8129), .S(n8355), .Z(n8131) );
  MUX2_X1 U27088 ( .A(n8131), .B(n8128), .S(n8262), .Z(n8132) );
  MUX2_X1 U27089 ( .A(\mem[38][7] ), .B(\mem[39][7] ), .S(n8535), .Z(n8133) );
  MUX2_X1 U27090 ( .A(\mem[36][7] ), .B(\mem[37][7] ), .S(n8535), .Z(n8134) );
  MUX2_X1 U27091 ( .A(n8134), .B(n8133), .S(n8355), .Z(n8135) );
  MUX2_X1 U27092 ( .A(\mem[34][7] ), .B(\mem[35][7] ), .S(n8535), .Z(n8136) );
  MUX2_X1 U27093 ( .A(\mem[32][7] ), .B(\mem[33][7] ), .S(n8535), .Z(n8137) );
  MUX2_X1 U27094 ( .A(n8137), .B(n8136), .S(n8355), .Z(n8138) );
  MUX2_X1 U27095 ( .A(n8138), .B(n8135), .S(n8262), .Z(n8139) );
  MUX2_X1 U27096 ( .A(n8139), .B(n8132), .S(n8218), .Z(n8140) );
  MUX2_X1 U27097 ( .A(n8140), .B(n8125), .S(n8194), .Z(n8141) );
  MUX2_X1 U27098 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n8535), .Z(n8142) );
  MUX2_X1 U27099 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n8535), .Z(n8143) );
  MUX2_X1 U27100 ( .A(n8143), .B(n8142), .S(n8355), .Z(n8144) );
  MUX2_X1 U27101 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n8535), .Z(n8145) );
  MUX2_X1 U27102 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n8535), .Z(n8146) );
  MUX2_X1 U27103 ( .A(n8146), .B(n8145), .S(n8355), .Z(n8147) );
  MUX2_X1 U27104 ( .A(n8147), .B(n8144), .S(n8262), .Z(n8148) );
  MUX2_X1 U27105 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n8536), .Z(n8149) );
  MUX2_X1 U27106 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n8536), .Z(n8150) );
  MUX2_X1 U27107 ( .A(n8150), .B(n8149), .S(n8355), .Z(n8151) );
  MUX2_X1 U27108 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n8536), .Z(n8152) );
  MUX2_X1 U27109 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n8536), .Z(n8153) );
  MUX2_X1 U27110 ( .A(n8153), .B(n8152), .S(n8355), .Z(n8154) );
  MUX2_X1 U27111 ( .A(n8154), .B(n8151), .S(n8262), .Z(n8155) );
  MUX2_X1 U27112 ( .A(n8155), .B(n8148), .S(n8218), .Z(n8156) );
  MUX2_X1 U27113 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n8536), .Z(n8157) );
  MUX2_X1 U27114 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n8536), .Z(n8158) );
  MUX2_X1 U27115 ( .A(n8158), .B(n8157), .S(n8355), .Z(n8159) );
  MUX2_X1 U27116 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n8536), .Z(n8160) );
  MUX2_X1 U27117 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n8536), .Z(n8161) );
  MUX2_X1 U27118 ( .A(n8161), .B(n8160), .S(n8355), .Z(n8162) );
  MUX2_X1 U27119 ( .A(n8162), .B(n8159), .S(n8262), .Z(n8163) );
  MUX2_X1 U27120 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n8536), .Z(n8164) );
  MUX2_X1 U27121 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n8536), .Z(n8165) );
  MUX2_X1 U27122 ( .A(n8165), .B(n8164), .S(n8355), .Z(n8166) );
  MUX2_X1 U27123 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n8536), .Z(n8167) );
  MUX2_X1 U27124 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n8536), .Z(n8168) );
  MUX2_X1 U27125 ( .A(n8168), .B(n8167), .S(n8355), .Z(n8169) );
  MUX2_X1 U27126 ( .A(n8169), .B(n8166), .S(n8262), .Z(n8170) );
  MUX2_X1 U27127 ( .A(n8170), .B(n8163), .S(n8218), .Z(n8171) );
  MUX2_X1 U27128 ( .A(n8171), .B(n8156), .S(n8194), .Z(n8172) );
  MUX2_X1 U27129 ( .A(n8172), .B(n8141), .S(n8185), .Z(n8173) );
  MUX2_X1 U27130 ( .A(n8173), .B(n8110), .S(n8180), .Z(n8174) );
  MUX2_X1 U27131 ( .A(n8174), .B(n8047), .S(n8177), .Z(n8175) );
  MUX2_X1 U27132 ( .A(n8175), .B(n7920), .S(N26), .Z(n8176) );
  MUX2_X1 U27133 ( .A(n8176), .B(n7665), .S(N27), .Z(N28) );
  CLKBUF_X1 U27134 ( .A(N24), .Z(n8178) );
  CLKBUF_X1 U27135 ( .A(n8225), .Z(n8226) );
  CLKBUF_X1 U27136 ( .A(n8388), .Z(n8389) );
  INV_X1 U27137 ( .A(N18), .ZN(n8604) );
  INV_X1 U27138 ( .A(N19), .ZN(n8605) );
  INV_X1 U27139 ( .A(N21), .ZN(n8606) );
  INV_X1 U27140 ( .A(N23), .ZN(n8607) );
  INV_X1 U27141 ( .A(N24), .ZN(n8608) );
endmodule


module memory_WIDTH16_SIZE32_LOGSIZE6 ( clk, data_in, data_out, addr, wr_en );
  input [15:0] data_in;
  output [15:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][15] , \mem[31][14] , \mem[31][13] ,
         \mem[31][12] , \mem[31][11] , \mem[31][10] , \mem[31][9] ,
         \mem[31][8] , \mem[31][7] , \mem[31][6] , \mem[31][5] , \mem[31][4] ,
         \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] , \mem[30][15] ,
         \mem[30][14] , \mem[30][13] , \mem[30][12] , \mem[30][11] ,
         \mem[30][10] , \mem[30][9] , \mem[30][8] , \mem[30][7] , \mem[30][6] ,
         \mem[30][5] , \mem[30][4] , \mem[30][3] , \mem[30][2] , \mem[30][1] ,
         \mem[30][0] , \mem[29][15] , \mem[29][14] , \mem[29][13] ,
         \mem[29][12] , \mem[29][11] , \mem[29][10] , \mem[29][9] ,
         \mem[29][8] , \mem[29][7] , \mem[29][6] , \mem[29][5] , \mem[29][4] ,
         \mem[29][3] , \mem[29][2] , \mem[29][1] , \mem[29][0] , \mem[28][15] ,
         \mem[28][14] , \mem[28][13] , \mem[28][12] , \mem[28][11] ,
         \mem[28][10] , \mem[28][9] , \mem[28][8] , \mem[28][7] , \mem[28][6] ,
         \mem[28][5] , \mem[28][4] , \mem[28][3] , \mem[28][2] , \mem[28][1] ,
         \mem[28][0] , \mem[27][15] , \mem[27][14] , \mem[27][13] ,
         \mem[27][12] , \mem[27][11] , \mem[27][10] , \mem[27][9] ,
         \mem[27][8] , \mem[27][7] , \mem[27][6] , \mem[27][5] , \mem[27][4] ,
         \mem[27][3] , \mem[27][2] , \mem[27][1] , \mem[27][0] , \mem[26][15] ,
         \mem[26][14] , \mem[26][13] , \mem[26][12] , \mem[26][11] ,
         \mem[26][10] , \mem[26][9] , \mem[26][8] , \mem[26][7] , \mem[26][6] ,
         \mem[26][5] , \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] ,
         \mem[26][0] , \mem[25][15] , \mem[25][14] , \mem[25][13] ,
         \mem[25][12] , \mem[25][11] , \mem[25][10] , \mem[25][9] ,
         \mem[25][8] , \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] ,
         \mem[25][3] , \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][15] ,
         \mem[24][14] , \mem[24][13] , \mem[24][12] , \mem[24][11] ,
         \mem[24][10] , \mem[24][9] , \mem[24][8] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][15] , \mem[23][14] , \mem[23][13] ,
         \mem[23][12] , \mem[23][11] , \mem[23][10] , \mem[23][9] ,
         \mem[23][8] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][15] ,
         \mem[22][14] , \mem[22][13] , \mem[22][12] , \mem[22][11] ,
         \mem[22][10] , \mem[22][9] , \mem[22][8] , \mem[22][7] , \mem[22][6] ,
         \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] , \mem[22][1] ,
         \mem[22][0] , \mem[21][15] , \mem[21][14] , \mem[21][13] ,
         \mem[21][12] , \mem[21][11] , \mem[21][10] , \mem[21][9] ,
         \mem[21][8] , \mem[21][7] , \mem[21][6] , \mem[21][5] , \mem[21][4] ,
         \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] , \mem[20][15] ,
         \mem[20][14] , \mem[20][13] , \mem[20][12] , \mem[20][11] ,
         \mem[20][10] , \mem[20][9] , \mem[20][8] , \mem[20][7] , \mem[20][6] ,
         \mem[20][5] , \mem[20][4] , \mem[20][3] , \mem[20][2] , \mem[20][1] ,
         \mem[20][0] , \mem[19][15] , \mem[19][14] , \mem[19][13] ,
         \mem[19][12] , \mem[19][11] , \mem[19][10] , \mem[19][9] ,
         \mem[19][8] , \mem[19][7] , \mem[19][6] , \mem[19][5] , \mem[19][4] ,
         \mem[19][3] , \mem[19][2] , \mem[19][1] , \mem[19][0] , \mem[18][15] ,
         \mem[18][14] , \mem[18][13] , \mem[18][12] , \mem[18][11] ,
         \mem[18][10] , \mem[18][9] , \mem[18][8] , \mem[18][7] , \mem[18][6] ,
         \mem[18][5] , \mem[18][4] , \mem[18][3] , \mem[18][2] , \mem[18][1] ,
         \mem[18][0] , \mem[17][15] , \mem[17][14] , \mem[17][13] ,
         \mem[17][12] , \mem[17][11] , \mem[17][10] , \mem[17][9] ,
         \mem[17][8] , \mem[17][7] , \mem[17][6] , \mem[17][5] , \mem[17][4] ,
         \mem[17][3] , \mem[17][2] , \mem[17][1] , \mem[17][0] , \mem[16][15] ,
         \mem[16][14] , \mem[16][13] , \mem[16][12] , \mem[16][11] ,
         \mem[16][10] , \mem[16][9] , \mem[16][8] , \mem[16][7] , \mem[16][6] ,
         \mem[16][5] , \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] ,
         \mem[16][0] , \mem[15][15] , \mem[15][14] , \mem[15][13] ,
         \mem[15][12] , \mem[15][11] , \mem[15][10] , \mem[15][9] ,
         \mem[15][8] , \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] ,
         \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][15] ,
         \mem[14][14] , \mem[14][13] , \mem[14][12] , \mem[14][11] ,
         \mem[14][10] , \mem[14][9] , \mem[14][8] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][15] , \mem[13][14] , \mem[13][13] ,
         \mem[13][12] , \mem[13][11] , \mem[13][10] , \mem[13][9] ,
         \mem[13][8] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][15] ,
         \mem[12][14] , \mem[12][13] , \mem[12][12] , \mem[12][11] ,
         \mem[12][10] , \mem[12][9] , \mem[12][8] , \mem[12][7] , \mem[12][6] ,
         \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] , \mem[12][1] ,
         \mem[12][0] , \mem[11][15] , \mem[11][14] , \mem[11][13] ,
         \mem[11][12] , \mem[11][11] , \mem[11][10] , \mem[11][9] ,
         \mem[11][8] , \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] ,
         \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[10][15] ,
         \mem[10][14] , \mem[10][13] , \mem[10][12] , \mem[10][11] ,
         \mem[10][10] , \mem[10][9] , \mem[10][8] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[9][15] , \mem[9][14] , \mem[9][13] , \mem[9][12] ,
         \mem[9][11] , \mem[9][10] , \mem[9][9] , \mem[9][8] , \mem[9][7] ,
         \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] ,
         \mem[9][1] , \mem[9][0] , \mem[8][15] , \mem[8][14] , \mem[8][13] ,
         \mem[8][12] , \mem[8][11] , \mem[8][10] , \mem[8][9] , \mem[8][8] ,
         \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] , \mem[8][3] ,
         \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][15] , \mem[7][14] ,
         \mem[7][13] , \mem[7][12] , \mem[7][11] , \mem[7][10] , \mem[7][9] ,
         \mem[7][8] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][15] ,
         \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] ,
         \mem[4][11] , \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] ,
         \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] ,
         \mem[4][1] , \mem[4][0] , \mem[3][15] , \mem[3][14] , \mem[3][13] ,
         \mem[3][12] , \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] ,
         \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] ,
         \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][15] ,
         \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[15]  ( .D(N15), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N16), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N17), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N18), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N19), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N20), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N21), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N22), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N23), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N24), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N25), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N26), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N27), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N28), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N29), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N30), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][15]  ( .D(n1090), .CK(clk), .Q(\mem[31][15] ) );
  DFF_X1 \mem_reg[31][14]  ( .D(n1089), .CK(clk), .Q(\mem[31][14] ) );
  DFF_X1 \mem_reg[31][13]  ( .D(n1088), .CK(clk), .Q(\mem[31][13] ) );
  DFF_X1 \mem_reg[31][12]  ( .D(n1087), .CK(clk), .Q(\mem[31][12] ) );
  DFF_X1 \mem_reg[31][11]  ( .D(n1086), .CK(clk), .Q(\mem[31][11] ) );
  DFF_X1 \mem_reg[31][10]  ( .D(n1085), .CK(clk), .Q(\mem[31][10] ) );
  DFF_X1 \mem_reg[31][9]  ( .D(n1084), .CK(clk), .Q(\mem[31][9] ) );
  DFF_X1 \mem_reg[31][8]  ( .D(n1083), .CK(clk), .Q(\mem[31][8] ) );
  DFF_X1 \mem_reg[31][7]  ( .D(n1082), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n1081), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n1080), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n1079), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n1078), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n1077), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n1076), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n1075), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][15]  ( .D(n1074), .CK(clk), .Q(\mem[30][15] ) );
  DFF_X1 \mem_reg[30][14]  ( .D(n1073), .CK(clk), .Q(\mem[30][14] ) );
  DFF_X1 \mem_reg[30][13]  ( .D(n1072), .CK(clk), .Q(\mem[30][13] ) );
  DFF_X1 \mem_reg[30][12]  ( .D(n1071), .CK(clk), .Q(\mem[30][12] ) );
  DFF_X1 \mem_reg[30][11]  ( .D(n1070), .CK(clk), .Q(\mem[30][11] ) );
  DFF_X1 \mem_reg[30][10]  ( .D(n1069), .CK(clk), .Q(\mem[30][10] ) );
  DFF_X1 \mem_reg[30][9]  ( .D(n1068), .CK(clk), .Q(\mem[30][9] ) );
  DFF_X1 \mem_reg[30][8]  ( .D(n1067), .CK(clk), .Q(\mem[30][8] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n1066), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n1065), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n1064), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n1063), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n1062), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n1061), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n1060), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n1059), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][15]  ( .D(n1058), .CK(clk), .Q(\mem[29][15] ) );
  DFF_X1 \mem_reg[29][14]  ( .D(n1057), .CK(clk), .Q(\mem[29][14] ) );
  DFF_X1 \mem_reg[29][13]  ( .D(n1056), .CK(clk), .Q(\mem[29][13] ) );
  DFF_X1 \mem_reg[29][12]  ( .D(n1055), .CK(clk), .Q(\mem[29][12] ) );
  DFF_X1 \mem_reg[29][11]  ( .D(n1054), .CK(clk), .Q(\mem[29][11] ) );
  DFF_X1 \mem_reg[29][10]  ( .D(n1053), .CK(clk), .Q(\mem[29][10] ) );
  DFF_X1 \mem_reg[29][9]  ( .D(n1052), .CK(clk), .Q(\mem[29][9] ) );
  DFF_X1 \mem_reg[29][8]  ( .D(n1051), .CK(clk), .Q(\mem[29][8] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n1050), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n1049), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n1048), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n1047), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n1046), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n1045), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n1044), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n1043), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][15]  ( .D(n1042), .CK(clk), .Q(\mem[28][15] ) );
  DFF_X1 \mem_reg[28][14]  ( .D(n1041), .CK(clk), .Q(\mem[28][14] ) );
  DFF_X1 \mem_reg[28][13]  ( .D(n1040), .CK(clk), .Q(\mem[28][13] ) );
  DFF_X1 \mem_reg[28][12]  ( .D(n1039), .CK(clk), .Q(\mem[28][12] ) );
  DFF_X1 \mem_reg[28][11]  ( .D(n1038), .CK(clk), .Q(\mem[28][11] ) );
  DFF_X1 \mem_reg[28][10]  ( .D(n1037), .CK(clk), .Q(\mem[28][10] ) );
  DFF_X1 \mem_reg[28][9]  ( .D(n1036), .CK(clk), .Q(\mem[28][9] ) );
  DFF_X1 \mem_reg[28][8]  ( .D(n1035), .CK(clk), .Q(\mem[28][8] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n1034), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n1033), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n1032), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n1031), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n1030), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n1029), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n1028), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n1027), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][15]  ( .D(n1026), .CK(clk), .Q(\mem[27][15] ) );
  DFF_X1 \mem_reg[27][14]  ( .D(n1025), .CK(clk), .Q(\mem[27][14] ) );
  DFF_X1 \mem_reg[27][13]  ( .D(n1024), .CK(clk), .Q(\mem[27][13] ) );
  DFF_X1 \mem_reg[27][12]  ( .D(n1023), .CK(clk), .Q(\mem[27][12] ) );
  DFF_X1 \mem_reg[27][11]  ( .D(n1022), .CK(clk), .Q(\mem[27][11] ) );
  DFF_X1 \mem_reg[27][10]  ( .D(n1021), .CK(clk), .Q(\mem[27][10] ) );
  DFF_X1 \mem_reg[27][9]  ( .D(n1020), .CK(clk), .Q(\mem[27][9] ) );
  DFF_X1 \mem_reg[27][8]  ( .D(n1019), .CK(clk), .Q(\mem[27][8] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n1018), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n1017), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n1016), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n1015), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n1014), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n1013), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n1012), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n1011), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][15]  ( .D(n1010), .CK(clk), .Q(\mem[26][15] ) );
  DFF_X1 \mem_reg[26][14]  ( .D(n1009), .CK(clk), .Q(\mem[26][14] ) );
  DFF_X1 \mem_reg[26][13]  ( .D(n1008), .CK(clk), .Q(\mem[26][13] ) );
  DFF_X1 \mem_reg[26][12]  ( .D(n1007), .CK(clk), .Q(\mem[26][12] ) );
  DFF_X1 \mem_reg[26][11]  ( .D(n1006), .CK(clk), .Q(\mem[26][11] ) );
  DFF_X1 \mem_reg[26][10]  ( .D(n1005), .CK(clk), .Q(\mem[26][10] ) );
  DFF_X1 \mem_reg[26][9]  ( .D(n1004), .CK(clk), .Q(\mem[26][9] ) );
  DFF_X1 \mem_reg[26][8]  ( .D(n1003), .CK(clk), .Q(\mem[26][8] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n1002), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n1001), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n1000), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n999), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n998), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n997), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n996), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n995), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][15]  ( .D(n994), .CK(clk), .Q(\mem[25][15] ) );
  DFF_X1 \mem_reg[25][14]  ( .D(n993), .CK(clk), .Q(\mem[25][14] ) );
  DFF_X1 \mem_reg[25][13]  ( .D(n992), .CK(clk), .Q(\mem[25][13] ) );
  DFF_X1 \mem_reg[25][12]  ( .D(n991), .CK(clk), .Q(\mem[25][12] ) );
  DFF_X1 \mem_reg[25][11]  ( .D(n990), .CK(clk), .Q(\mem[25][11] ) );
  DFF_X1 \mem_reg[25][10]  ( .D(n989), .CK(clk), .Q(\mem[25][10] ) );
  DFF_X1 \mem_reg[25][9]  ( .D(n988), .CK(clk), .Q(\mem[25][9] ) );
  DFF_X1 \mem_reg[25][8]  ( .D(n987), .CK(clk), .Q(\mem[25][8] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n986), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n985), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n984), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n983), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n982), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n981), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n980), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n979), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][15]  ( .D(n978), .CK(clk), .Q(\mem[24][15] ) );
  DFF_X1 \mem_reg[24][14]  ( .D(n977), .CK(clk), .Q(\mem[24][14] ) );
  DFF_X1 \mem_reg[24][13]  ( .D(n976), .CK(clk), .Q(\mem[24][13] ) );
  DFF_X1 \mem_reg[24][12]  ( .D(n975), .CK(clk), .Q(\mem[24][12] ) );
  DFF_X1 \mem_reg[24][11]  ( .D(n974), .CK(clk), .Q(\mem[24][11] ) );
  DFF_X1 \mem_reg[24][10]  ( .D(n973), .CK(clk), .Q(\mem[24][10] ) );
  DFF_X1 \mem_reg[24][9]  ( .D(n972), .CK(clk), .Q(\mem[24][9] ) );
  DFF_X1 \mem_reg[24][8]  ( .D(n971), .CK(clk), .Q(\mem[24][8] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n970), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n969), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n968), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n967), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n966), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n965), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n964), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n963), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][15]  ( .D(n962), .CK(clk), .Q(\mem[23][15] ) );
  DFF_X1 \mem_reg[23][14]  ( .D(n961), .CK(clk), .Q(\mem[23][14] ) );
  DFF_X1 \mem_reg[23][13]  ( .D(n960), .CK(clk), .Q(\mem[23][13] ) );
  DFF_X1 \mem_reg[23][12]  ( .D(n959), .CK(clk), .Q(\mem[23][12] ) );
  DFF_X1 \mem_reg[23][11]  ( .D(n958), .CK(clk), .Q(\mem[23][11] ) );
  DFF_X1 \mem_reg[23][10]  ( .D(n957), .CK(clk), .Q(\mem[23][10] ) );
  DFF_X1 \mem_reg[23][9]  ( .D(n956), .CK(clk), .Q(\mem[23][9] ) );
  DFF_X1 \mem_reg[23][8]  ( .D(n955), .CK(clk), .Q(\mem[23][8] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n954), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n953), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n952), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n951), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n950), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n949), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n948), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n947), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][15]  ( .D(n946), .CK(clk), .Q(\mem[22][15] ) );
  DFF_X1 \mem_reg[22][14]  ( .D(n945), .CK(clk), .Q(\mem[22][14] ) );
  DFF_X1 \mem_reg[22][13]  ( .D(n944), .CK(clk), .Q(\mem[22][13] ) );
  DFF_X1 \mem_reg[22][12]  ( .D(n943), .CK(clk), .Q(\mem[22][12] ) );
  DFF_X1 \mem_reg[22][11]  ( .D(n942), .CK(clk), .Q(\mem[22][11] ) );
  DFF_X1 \mem_reg[22][10]  ( .D(n941), .CK(clk), .Q(\mem[22][10] ) );
  DFF_X1 \mem_reg[22][9]  ( .D(n940), .CK(clk), .Q(\mem[22][9] ) );
  DFF_X1 \mem_reg[22][8]  ( .D(n939), .CK(clk), .Q(\mem[22][8] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n938), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n937), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n936), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n935), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n934), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n933), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n932), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n931), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][15]  ( .D(n930), .CK(clk), .Q(\mem[21][15] ) );
  DFF_X1 \mem_reg[21][14]  ( .D(n929), .CK(clk), .Q(\mem[21][14] ) );
  DFF_X1 \mem_reg[21][13]  ( .D(n928), .CK(clk), .Q(\mem[21][13] ) );
  DFF_X1 \mem_reg[21][12]  ( .D(n927), .CK(clk), .Q(\mem[21][12] ) );
  DFF_X1 \mem_reg[21][11]  ( .D(n926), .CK(clk), .Q(\mem[21][11] ) );
  DFF_X1 \mem_reg[21][10]  ( .D(n925), .CK(clk), .Q(\mem[21][10] ) );
  DFF_X1 \mem_reg[21][9]  ( .D(n924), .CK(clk), .Q(\mem[21][9] ) );
  DFF_X1 \mem_reg[21][8]  ( .D(n923), .CK(clk), .Q(\mem[21][8] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n922), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n921), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n920), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n919), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n918), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n917), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n916), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n915), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][15]  ( .D(n914), .CK(clk), .Q(\mem[20][15] ) );
  DFF_X1 \mem_reg[20][14]  ( .D(n913), .CK(clk), .Q(\mem[20][14] ) );
  DFF_X1 \mem_reg[20][13]  ( .D(n912), .CK(clk), .Q(\mem[20][13] ) );
  DFF_X1 \mem_reg[20][12]  ( .D(n911), .CK(clk), .Q(\mem[20][12] ) );
  DFF_X1 \mem_reg[20][11]  ( .D(n910), .CK(clk), .Q(\mem[20][11] ) );
  DFF_X1 \mem_reg[20][10]  ( .D(n909), .CK(clk), .Q(\mem[20][10] ) );
  DFF_X1 \mem_reg[20][9]  ( .D(n908), .CK(clk), .Q(\mem[20][9] ) );
  DFF_X1 \mem_reg[20][8]  ( .D(n907), .CK(clk), .Q(\mem[20][8] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n906), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n905), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n904), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n903), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n902), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n901), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n900), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n899), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][15]  ( .D(n898), .CK(clk), .Q(\mem[19][15] ) );
  DFF_X1 \mem_reg[19][14]  ( .D(n897), .CK(clk), .Q(\mem[19][14] ) );
  DFF_X1 \mem_reg[19][13]  ( .D(n896), .CK(clk), .Q(\mem[19][13] ) );
  DFF_X1 \mem_reg[19][12]  ( .D(n895), .CK(clk), .Q(\mem[19][12] ) );
  DFF_X1 \mem_reg[19][11]  ( .D(n894), .CK(clk), .Q(\mem[19][11] ) );
  DFF_X1 \mem_reg[19][10]  ( .D(n893), .CK(clk), .Q(\mem[19][10] ) );
  DFF_X1 \mem_reg[19][9]  ( .D(n892), .CK(clk), .Q(\mem[19][9] ) );
  DFF_X1 \mem_reg[19][8]  ( .D(n891), .CK(clk), .Q(\mem[19][8] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n890), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n889), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n888), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n887), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n886), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n885), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n884), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n883), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][15]  ( .D(n882), .CK(clk), .Q(\mem[18][15] ) );
  DFF_X1 \mem_reg[18][14]  ( .D(n881), .CK(clk), .Q(\mem[18][14] ) );
  DFF_X1 \mem_reg[18][13]  ( .D(n880), .CK(clk), .Q(\mem[18][13] ) );
  DFF_X1 \mem_reg[18][12]  ( .D(n879), .CK(clk), .Q(\mem[18][12] ) );
  DFF_X1 \mem_reg[18][11]  ( .D(n878), .CK(clk), .Q(\mem[18][11] ) );
  DFF_X1 \mem_reg[18][10]  ( .D(n877), .CK(clk), .Q(\mem[18][10] ) );
  DFF_X1 \mem_reg[18][9]  ( .D(n876), .CK(clk), .Q(\mem[18][9] ) );
  DFF_X1 \mem_reg[18][8]  ( .D(n875), .CK(clk), .Q(\mem[18][8] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n874), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n873), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n872), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n871), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n870), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n869), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n868), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n867), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][15]  ( .D(n866), .CK(clk), .Q(\mem[17][15] ) );
  DFF_X1 \mem_reg[17][14]  ( .D(n865), .CK(clk), .Q(\mem[17][14] ) );
  DFF_X1 \mem_reg[17][13]  ( .D(n864), .CK(clk), .Q(\mem[17][13] ) );
  DFF_X1 \mem_reg[17][12]  ( .D(n863), .CK(clk), .Q(\mem[17][12] ) );
  DFF_X1 \mem_reg[17][11]  ( .D(n862), .CK(clk), .Q(\mem[17][11] ) );
  DFF_X1 \mem_reg[17][10]  ( .D(n861), .CK(clk), .Q(\mem[17][10] ) );
  DFF_X1 \mem_reg[17][9]  ( .D(n860), .CK(clk), .Q(\mem[17][9] ) );
  DFF_X1 \mem_reg[17][8]  ( .D(n859), .CK(clk), .Q(\mem[17][8] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n858), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n857), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n856), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n855), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n854), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n853), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n852), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n851), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][15]  ( .D(n850), .CK(clk), .Q(\mem[16][15] ) );
  DFF_X1 \mem_reg[16][14]  ( .D(n849), .CK(clk), .Q(\mem[16][14] ) );
  DFF_X1 \mem_reg[16][13]  ( .D(n848), .CK(clk), .Q(\mem[16][13] ) );
  DFF_X1 \mem_reg[16][12]  ( .D(n847), .CK(clk), .Q(\mem[16][12] ) );
  DFF_X1 \mem_reg[16][11]  ( .D(n846), .CK(clk), .Q(\mem[16][11] ) );
  DFF_X1 \mem_reg[16][10]  ( .D(n845), .CK(clk), .Q(\mem[16][10] ) );
  DFF_X1 \mem_reg[16][9]  ( .D(n844), .CK(clk), .Q(\mem[16][9] ) );
  DFF_X1 \mem_reg[16][8]  ( .D(n843), .CK(clk), .Q(\mem[16][8] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n842), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n841), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n840), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n839), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n838), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n837), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n836), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n835), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][15]  ( .D(n834), .CK(clk), .Q(\mem[15][15] ) );
  DFF_X1 \mem_reg[15][14]  ( .D(n833), .CK(clk), .Q(\mem[15][14] ) );
  DFF_X1 \mem_reg[15][13]  ( .D(n832), .CK(clk), .Q(\mem[15][13] ) );
  DFF_X1 \mem_reg[15][12]  ( .D(n831), .CK(clk), .Q(\mem[15][12] ) );
  DFF_X1 \mem_reg[15][11]  ( .D(n830), .CK(clk), .Q(\mem[15][11] ) );
  DFF_X1 \mem_reg[15][10]  ( .D(n829), .CK(clk), .Q(\mem[15][10] ) );
  DFF_X1 \mem_reg[15][9]  ( .D(n828), .CK(clk), .Q(\mem[15][9] ) );
  DFF_X1 \mem_reg[15][8]  ( .D(n827), .CK(clk), .Q(\mem[15][8] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n826), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n825), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n824), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n823), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n822), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n821), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n820), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n819), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][15]  ( .D(n818), .CK(clk), .Q(\mem[14][15] ) );
  DFF_X1 \mem_reg[14][14]  ( .D(n817), .CK(clk), .Q(\mem[14][14] ) );
  DFF_X1 \mem_reg[14][13]  ( .D(n816), .CK(clk), .Q(\mem[14][13] ) );
  DFF_X1 \mem_reg[14][12]  ( .D(n815), .CK(clk), .Q(\mem[14][12] ) );
  DFF_X1 \mem_reg[14][11]  ( .D(n814), .CK(clk), .Q(\mem[14][11] ) );
  DFF_X1 \mem_reg[14][10]  ( .D(n813), .CK(clk), .Q(\mem[14][10] ) );
  DFF_X1 \mem_reg[14][9]  ( .D(n812), .CK(clk), .Q(\mem[14][9] ) );
  DFF_X1 \mem_reg[14][8]  ( .D(n811), .CK(clk), .Q(\mem[14][8] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n810), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n809), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n808), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n807), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n806), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n805), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n804), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n803), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][15]  ( .D(n802), .CK(clk), .Q(\mem[13][15] ) );
  DFF_X1 \mem_reg[13][14]  ( .D(n801), .CK(clk), .Q(\mem[13][14] ) );
  DFF_X1 \mem_reg[13][13]  ( .D(n800), .CK(clk), .Q(\mem[13][13] ) );
  DFF_X1 \mem_reg[13][12]  ( .D(n799), .CK(clk), .Q(\mem[13][12] ) );
  DFF_X1 \mem_reg[13][11]  ( .D(n798), .CK(clk), .Q(\mem[13][11] ) );
  DFF_X1 \mem_reg[13][10]  ( .D(n797), .CK(clk), .Q(\mem[13][10] ) );
  DFF_X1 \mem_reg[13][9]  ( .D(n796), .CK(clk), .Q(\mem[13][9] ) );
  DFF_X1 \mem_reg[13][8]  ( .D(n795), .CK(clk), .Q(\mem[13][8] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n794), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n793), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n792), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n791), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n790), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n789), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n788), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n787), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][15]  ( .D(n786), .CK(clk), .Q(\mem[12][15] ) );
  DFF_X1 \mem_reg[12][14]  ( .D(n785), .CK(clk), .Q(\mem[12][14] ) );
  DFF_X1 \mem_reg[12][13]  ( .D(n784), .CK(clk), .Q(\mem[12][13] ) );
  DFF_X1 \mem_reg[12][12]  ( .D(n783), .CK(clk), .Q(\mem[12][12] ) );
  DFF_X1 \mem_reg[12][11]  ( .D(n782), .CK(clk), .Q(\mem[12][11] ) );
  DFF_X1 \mem_reg[12][10]  ( .D(n781), .CK(clk), .Q(\mem[12][10] ) );
  DFF_X1 \mem_reg[12][9]  ( .D(n780), .CK(clk), .Q(\mem[12][9] ) );
  DFF_X1 \mem_reg[12][8]  ( .D(n779), .CK(clk), .Q(\mem[12][8] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n778), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n777), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n776), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n775), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n774), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n773), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n772), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n771), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][15]  ( .D(n770), .CK(clk), .Q(\mem[11][15] ) );
  DFF_X1 \mem_reg[11][14]  ( .D(n769), .CK(clk), .Q(\mem[11][14] ) );
  DFF_X1 \mem_reg[11][13]  ( .D(n768), .CK(clk), .Q(\mem[11][13] ) );
  DFF_X1 \mem_reg[11][12]  ( .D(n767), .CK(clk), .Q(\mem[11][12] ) );
  DFF_X1 \mem_reg[11][11]  ( .D(n766), .CK(clk), .Q(\mem[11][11] ) );
  DFF_X1 \mem_reg[11][10]  ( .D(n765), .CK(clk), .Q(\mem[11][10] ) );
  DFF_X1 \mem_reg[11][9]  ( .D(n764), .CK(clk), .Q(\mem[11][9] ) );
  DFF_X1 \mem_reg[11][8]  ( .D(n763), .CK(clk), .Q(\mem[11][8] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n762), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n761), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n760), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n759), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n758), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n757), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n756), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n755), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][15]  ( .D(n754), .CK(clk), .Q(\mem[10][15] ) );
  DFF_X1 \mem_reg[10][14]  ( .D(n753), .CK(clk), .Q(\mem[10][14] ) );
  DFF_X1 \mem_reg[10][13]  ( .D(n752), .CK(clk), .Q(\mem[10][13] ) );
  DFF_X1 \mem_reg[10][12]  ( .D(n751), .CK(clk), .Q(\mem[10][12] ) );
  DFF_X1 \mem_reg[10][11]  ( .D(n750), .CK(clk), .Q(\mem[10][11] ) );
  DFF_X1 \mem_reg[10][10]  ( .D(n749), .CK(clk), .Q(\mem[10][10] ) );
  DFF_X1 \mem_reg[10][9]  ( .D(n748), .CK(clk), .Q(\mem[10][9] ) );
  DFF_X1 \mem_reg[10][8]  ( .D(n747), .CK(clk), .Q(\mem[10][8] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n746), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n745), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n744), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n743), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n742), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n741), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n740), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n739), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][15]  ( .D(n738), .CK(clk), .Q(\mem[9][15] ) );
  DFF_X1 \mem_reg[9][14]  ( .D(n737), .CK(clk), .Q(\mem[9][14] ) );
  DFF_X1 \mem_reg[9][13]  ( .D(n736), .CK(clk), .Q(\mem[9][13] ) );
  DFF_X1 \mem_reg[9][12]  ( .D(n735), .CK(clk), .Q(\mem[9][12] ) );
  DFF_X1 \mem_reg[9][11]  ( .D(n734), .CK(clk), .Q(\mem[9][11] ) );
  DFF_X1 \mem_reg[9][10]  ( .D(n733), .CK(clk), .Q(\mem[9][10] ) );
  DFF_X1 \mem_reg[9][9]  ( .D(n732), .CK(clk), .Q(\mem[9][9] ) );
  DFF_X1 \mem_reg[9][8]  ( .D(n731), .CK(clk), .Q(\mem[9][8] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n729), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n728), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n727), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n726), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n725), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n724), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n723), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][15]  ( .D(n722), .CK(clk), .Q(\mem[8][15] ) );
  DFF_X1 \mem_reg[8][14]  ( .D(n721), .CK(clk), .Q(\mem[8][14] ) );
  DFF_X1 \mem_reg[8][13]  ( .D(n720), .CK(clk), .Q(\mem[8][13] ) );
  DFF_X1 \mem_reg[8][12]  ( .D(n719), .CK(clk), .Q(\mem[8][12] ) );
  DFF_X1 \mem_reg[8][11]  ( .D(n718), .CK(clk), .Q(\mem[8][11] ) );
  DFF_X1 \mem_reg[8][10]  ( .D(n717), .CK(clk), .Q(\mem[8][10] ) );
  DFF_X1 \mem_reg[8][9]  ( .D(n716), .CK(clk), .Q(\mem[8][9] ) );
  DFF_X1 \mem_reg[8][8]  ( .D(n715), .CK(clk), .Q(\mem[8][8] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n714), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n713), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n712), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n711), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n710), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n709), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n708), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n707), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n706), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n705), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n704), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n703), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n702), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n701), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n700), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n699), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n698), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n697), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n696), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n695), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n694), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n693), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n692), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n691), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n690), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n689), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n688), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n687), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n686), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n685), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n684), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n683), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n682), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n681), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n680), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n679), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n678), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n677), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n676), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n675), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n674), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n673), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n672), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n671), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n670), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n669), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n668), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n667), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n666), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n665), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n664), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n663), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n662), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n661), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n660), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n659), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n658), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n657), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n656), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n655), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n654), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n653), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n652), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n651), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n650), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n649), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n648), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n647), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n646), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n645), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n644), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n643), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n642), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n641), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n640), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n639), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n638), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n637), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n636), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n635), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n634), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n633), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n632), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n631), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n630), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n629), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n628), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n627), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n626), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n625), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n624), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n623), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n622), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n621), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n620), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n619), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n618), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n617), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n616), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n615), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n614), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n613), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n612), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n611), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n610), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n609), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n608), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n607), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n606), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n605), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n604), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n603), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n602), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n601), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n600), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n599), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n598), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n597), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n596), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n595), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n594), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n593), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n592), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n591), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n590), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n589), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n588), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n587), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n586), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n585), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n584), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n583), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n582), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n581), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n580), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n579), .CK(clk), .Q(\mem[0][0] ) );
  BUF_X1 U3 ( .A(N10), .Z(n1561) );
  CLKBUF_X1 U4 ( .A(N11), .Z(n1557) );
  CLKBUF_X1 U5 ( .A(n1560), .Z(n1558) );
  CLKBUF_X1 U6 ( .A(n1560), .Z(n1559) );
  BUF_X1 U7 ( .A(n1572), .Z(n1568) );
  BUF_X1 U8 ( .A(n1572), .Z(n1569) );
  BUF_X1 U9 ( .A(n1572), .Z(n1570) );
  BUF_X1 U10 ( .A(n1571), .Z(n1564) );
  BUF_X1 U11 ( .A(n1572), .Z(n1565) );
  BUF_X1 U12 ( .A(n1572), .Z(n1566) );
  BUF_X1 U13 ( .A(n1572), .Z(n1567) );
  BUF_X1 U14 ( .A(n1571), .Z(n1562) );
  BUF_X1 U15 ( .A(n1571), .Z(n1563) );
  BUF_X1 U16 ( .A(n1560), .Z(n1556) );
  BUF_X1 U17 ( .A(n1571), .Z(n1572) );
  BUF_X1 U18 ( .A(n22), .Z(n1620) );
  BUF_X1 U19 ( .A(n168), .Z(n1612) );
  BUF_X1 U20 ( .A(n186), .Z(n1611) );
  BUF_X1 U21 ( .A(n203), .Z(n1610) );
  BUF_X1 U22 ( .A(n305), .Z(n1604) );
  BUF_X1 U23 ( .A(n340), .Z(n1602) );
  BUF_X1 U24 ( .A(n357), .Z(n1601) );
  BUF_X1 U25 ( .A(n460), .Z(n1595) );
  BUF_X1 U26 ( .A(n477), .Z(n1594) );
  BUF_X1 U27 ( .A(n494), .Z(n1593) );
  BUF_X1 U28 ( .A(n41), .Z(n1619) );
  BUF_X1 U29 ( .A(n59), .Z(n1618) );
  BUF_X1 U30 ( .A(n77), .Z(n1617) );
  BUF_X1 U31 ( .A(n95), .Z(n1616) );
  BUF_X1 U32 ( .A(n113), .Z(n1615) );
  BUF_X1 U33 ( .A(n149), .Z(n1613) );
  BUF_X1 U34 ( .A(n237), .Z(n1608) );
  BUF_X1 U35 ( .A(n271), .Z(n1606) );
  BUF_X1 U36 ( .A(n288), .Z(n1605) );
  BUF_X1 U37 ( .A(n391), .Z(n1599) );
  BUF_X1 U38 ( .A(n408), .Z(n1598) );
  BUF_X1 U39 ( .A(n425), .Z(n1597) );
  BUF_X1 U40 ( .A(n511), .Z(n1592) );
  BUF_X1 U41 ( .A(n528), .Z(n1591) );
  BUF_X1 U42 ( .A(n545), .Z(n1590) );
  BUF_X1 U43 ( .A(n562), .Z(n1589) );
  BUF_X1 U44 ( .A(n220), .Z(n1609) );
  BUF_X1 U45 ( .A(n442), .Z(n1596) );
  BUF_X1 U46 ( .A(n254), .Z(n1607) );
  BUF_X1 U47 ( .A(n323), .Z(n1603) );
  BUF_X1 U48 ( .A(n131), .Z(n1614) );
  BUF_X1 U49 ( .A(n374), .Z(n1600) );
  BUF_X1 U50 ( .A(N11), .Z(n1560) );
  BUF_X1 U51 ( .A(N10), .Z(n1571) );
  BUF_X1 U52 ( .A(N13), .Z(n1550) );
  BUF_X1 U53 ( .A(N13), .Z(n1551) );
  NAND2_X1 U54 ( .A1(n39), .A2(n40), .ZN(n22) );
  NAND2_X1 U55 ( .A1(n58), .A2(n40), .ZN(n41) );
  NAND2_X1 U56 ( .A1(n76), .A2(n40), .ZN(n59) );
  NAND2_X1 U57 ( .A1(n94), .A2(n40), .ZN(n77) );
  NAND2_X1 U58 ( .A1(n185), .A2(n39), .ZN(n168) );
  NAND2_X1 U59 ( .A1(n185), .A2(n58), .ZN(n186) );
  NAND2_X1 U60 ( .A1(n185), .A2(n76), .ZN(n203) );
  NAND2_X1 U61 ( .A1(n185), .A2(n94), .ZN(n220) );
  NAND2_X1 U62 ( .A1(n322), .A2(n39), .ZN(n305) );
  NAND2_X1 U63 ( .A1(n322), .A2(n58), .ZN(n323) );
  NAND2_X1 U64 ( .A1(n322), .A2(n76), .ZN(n340) );
  NAND2_X1 U65 ( .A1(n322), .A2(n94), .ZN(n357) );
  NAND2_X1 U66 ( .A1(n459), .A2(n39), .ZN(n442) );
  NAND2_X1 U67 ( .A1(n459), .A2(n58), .ZN(n460) );
  NAND2_X1 U68 ( .A1(n459), .A2(n76), .ZN(n477) );
  NAND2_X1 U69 ( .A1(n459), .A2(n94), .ZN(n494) );
  NAND2_X1 U70 ( .A1(n322), .A2(n112), .ZN(n374) );
  NAND2_X1 U71 ( .A1(n322), .A2(n130), .ZN(n391) );
  NAND2_X1 U72 ( .A1(n322), .A2(n148), .ZN(n408) );
  NAND2_X1 U73 ( .A1(n322), .A2(n166), .ZN(n425) );
  NAND2_X1 U74 ( .A1(n459), .A2(n112), .ZN(n511) );
  NAND2_X1 U75 ( .A1(n459), .A2(n130), .ZN(n528) );
  NAND2_X1 U76 ( .A1(n459), .A2(n148), .ZN(n545) );
  NAND2_X1 U77 ( .A1(n459), .A2(n166), .ZN(n562) );
  NAND2_X1 U78 ( .A1(n112), .A2(n40), .ZN(n95) );
  NAND2_X1 U79 ( .A1(n130), .A2(n40), .ZN(n113) );
  NAND2_X1 U80 ( .A1(n148), .A2(n40), .ZN(n131) );
  NAND2_X1 U81 ( .A1(n166), .A2(n40), .ZN(n149) );
  NAND2_X1 U82 ( .A1(n185), .A2(n112), .ZN(n237) );
  NAND2_X1 U83 ( .A1(n185), .A2(n130), .ZN(n254) );
  NAND2_X1 U84 ( .A1(n185), .A2(n148), .ZN(n271) );
  NAND2_X1 U85 ( .A1(n185), .A2(n166), .ZN(n288) );
  NOR3_X1 U86 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n39) );
  NOR3_X1 U87 ( .A1(N11), .A2(N12), .A3(n1621), .ZN(n58) );
  NOR3_X1 U88 ( .A1(N10), .A2(N12), .A3(n1622), .ZN(n76) );
  NOR3_X1 U89 ( .A1(n1621), .A2(N12), .A3(n1622), .ZN(n94) );
  AND3_X1 U90 ( .A1(n1623), .A2(n1640), .A3(n167), .ZN(n40) );
  AND3_X1 U91 ( .A1(n167), .A2(n1623), .A3(N14), .ZN(n322) );
  AND3_X1 U92 ( .A1(N13), .A2(n167), .A3(N14), .ZN(n459) );
  AND3_X1 U93 ( .A1(n167), .A2(n1640), .A3(N13), .ZN(n185) );
  INV_X1 U94 ( .A(N14), .ZN(n1640) );
  AND3_X1 U95 ( .A1(n1621), .A2(n1622), .A3(N12), .ZN(n112) );
  AND3_X1 U96 ( .A1(N10), .A2(n1622), .A3(N12), .ZN(n130) );
  AND3_X1 U97 ( .A1(N11), .A2(n1621), .A3(N12), .ZN(n148) );
  AND3_X1 U98 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n166) );
  BUF_X1 U99 ( .A(n1638), .Z(n1587) );
  BUF_X1 U100 ( .A(n1636), .Z(n1585) );
  BUF_X1 U101 ( .A(n1635), .Z(n1584) );
  BUF_X1 U102 ( .A(n1634), .Z(n1583) );
  BUF_X1 U103 ( .A(n1633), .Z(n1582) );
  BUF_X1 U104 ( .A(n1632), .Z(n1581) );
  BUF_X1 U105 ( .A(n1630), .Z(n1579) );
  BUF_X1 U106 ( .A(n1629), .Z(n1578) );
  BUF_X1 U107 ( .A(n1628), .Z(n1577) );
  BUF_X1 U108 ( .A(n1627), .Z(n1576) );
  BUF_X1 U109 ( .A(n1625), .Z(n1574) );
  BUF_X1 U110 ( .A(n1624), .Z(n1573) );
  BUF_X1 U111 ( .A(n1639), .Z(n1588) );
  BUF_X1 U112 ( .A(n1631), .Z(n1580) );
  BUF_X1 U113 ( .A(n1626), .Z(n1575) );
  BUF_X1 U114 ( .A(n1637), .Z(n1586) );
  NOR2_X1 U115 ( .A1(n1641), .A2(addr[5]), .ZN(n167) );
  INV_X1 U116 ( .A(wr_en), .ZN(n1641) );
  OAI21_X1 U117 ( .B1(n1581), .B2(n41), .A(n49), .ZN(n602) );
  NAND2_X1 U118 ( .A1(\mem[1][7] ), .A2(n41), .ZN(n49) );
  OAI21_X1 U119 ( .B1(n1631), .B2(n41), .A(n50), .ZN(n603) );
  NAND2_X1 U120 ( .A1(\mem[1][8] ), .A2(n1619), .ZN(n50) );
  OAI21_X1 U121 ( .B1(n1579), .B2(n41), .A(n51), .ZN(n604) );
  NAND2_X1 U122 ( .A1(\mem[1][9] ), .A2(n1619), .ZN(n51) );
  OAI21_X1 U123 ( .B1(n1578), .B2(n41), .A(n52), .ZN(n605) );
  NAND2_X1 U124 ( .A1(\mem[1][10] ), .A2(n1619), .ZN(n52) );
  OAI21_X1 U125 ( .B1(n1577), .B2(n41), .A(n53), .ZN(n606) );
  NAND2_X1 U126 ( .A1(\mem[1][11] ), .A2(n1619), .ZN(n53) );
  OAI21_X1 U127 ( .B1(n1576), .B2(n41), .A(n54), .ZN(n607) );
  NAND2_X1 U128 ( .A1(\mem[1][12] ), .A2(n1619), .ZN(n54) );
  OAI21_X1 U129 ( .B1(n1626), .B2(n41), .A(n55), .ZN(n608) );
  NAND2_X1 U130 ( .A1(\mem[1][13] ), .A2(n1619), .ZN(n55) );
  OAI21_X1 U131 ( .B1(n1574), .B2(n41), .A(n56), .ZN(n609) );
  NAND2_X1 U132 ( .A1(\mem[1][14] ), .A2(n1619), .ZN(n56) );
  OAI21_X1 U133 ( .B1(n1581), .B2(n59), .A(n67), .ZN(n618) );
  NAND2_X1 U134 ( .A1(\mem[2][7] ), .A2(n59), .ZN(n67) );
  OAI21_X1 U135 ( .B1(n1631), .B2(n59), .A(n68), .ZN(n619) );
  NAND2_X1 U136 ( .A1(\mem[2][8] ), .A2(n1618), .ZN(n68) );
  OAI21_X1 U137 ( .B1(n1579), .B2(n59), .A(n69), .ZN(n620) );
  NAND2_X1 U138 ( .A1(\mem[2][9] ), .A2(n1618), .ZN(n69) );
  OAI21_X1 U139 ( .B1(n1578), .B2(n59), .A(n70), .ZN(n621) );
  NAND2_X1 U140 ( .A1(\mem[2][10] ), .A2(n1618), .ZN(n70) );
  OAI21_X1 U141 ( .B1(n1577), .B2(n59), .A(n71), .ZN(n622) );
  NAND2_X1 U142 ( .A1(\mem[2][11] ), .A2(n1618), .ZN(n71) );
  OAI21_X1 U143 ( .B1(n1576), .B2(n59), .A(n72), .ZN(n623) );
  NAND2_X1 U144 ( .A1(\mem[2][12] ), .A2(n1618), .ZN(n72) );
  OAI21_X1 U145 ( .B1(n1626), .B2(n59), .A(n73), .ZN(n624) );
  NAND2_X1 U146 ( .A1(\mem[2][13] ), .A2(n1618), .ZN(n73) );
  OAI21_X1 U147 ( .B1(n1574), .B2(n59), .A(n74), .ZN(n625) );
  NAND2_X1 U148 ( .A1(\mem[2][14] ), .A2(n1618), .ZN(n74) );
  OAI21_X1 U149 ( .B1(n1581), .B2(n77), .A(n85), .ZN(n634) );
  NAND2_X1 U150 ( .A1(\mem[3][7] ), .A2(n77), .ZN(n85) );
  OAI21_X1 U151 ( .B1(n1631), .B2(n77), .A(n86), .ZN(n635) );
  NAND2_X1 U152 ( .A1(\mem[3][8] ), .A2(n1617), .ZN(n86) );
  OAI21_X1 U153 ( .B1(n1579), .B2(n77), .A(n87), .ZN(n636) );
  NAND2_X1 U154 ( .A1(\mem[3][9] ), .A2(n1617), .ZN(n87) );
  OAI21_X1 U155 ( .B1(n1578), .B2(n77), .A(n88), .ZN(n637) );
  NAND2_X1 U156 ( .A1(\mem[3][10] ), .A2(n1617), .ZN(n88) );
  OAI21_X1 U157 ( .B1(n1577), .B2(n77), .A(n89), .ZN(n638) );
  NAND2_X1 U158 ( .A1(\mem[3][11] ), .A2(n1617), .ZN(n89) );
  OAI21_X1 U159 ( .B1(n1576), .B2(n77), .A(n90), .ZN(n639) );
  NAND2_X1 U160 ( .A1(\mem[3][12] ), .A2(n1617), .ZN(n90) );
  OAI21_X1 U161 ( .B1(n1626), .B2(n77), .A(n91), .ZN(n640) );
  NAND2_X1 U162 ( .A1(\mem[3][13] ), .A2(n1617), .ZN(n91) );
  OAI21_X1 U163 ( .B1(n1574), .B2(n77), .A(n92), .ZN(n641) );
  NAND2_X1 U164 ( .A1(\mem[3][14] ), .A2(n1617), .ZN(n92) );
  OAI21_X1 U165 ( .B1(n1632), .B2(n305), .A(n313), .ZN(n842) );
  NAND2_X1 U166 ( .A1(\mem[16][7] ), .A2(n1604), .ZN(n313) );
  OAI21_X1 U167 ( .B1(n1580), .B2(n1604), .A(n314), .ZN(n843) );
  NAND2_X1 U168 ( .A1(\mem[16][8] ), .A2(n1604), .ZN(n314) );
  OAI21_X1 U169 ( .B1(n1630), .B2(n305), .A(n315), .ZN(n844) );
  NAND2_X1 U170 ( .A1(\mem[16][9] ), .A2(n1604), .ZN(n315) );
  OAI21_X1 U171 ( .B1(n1629), .B2(n305), .A(n316), .ZN(n845) );
  NAND2_X1 U172 ( .A1(\mem[16][10] ), .A2(n1604), .ZN(n316) );
  OAI21_X1 U173 ( .B1(n1628), .B2(n305), .A(n317), .ZN(n846) );
  NAND2_X1 U174 ( .A1(\mem[16][11] ), .A2(n1604), .ZN(n317) );
  OAI21_X1 U175 ( .B1(n1627), .B2(n305), .A(n318), .ZN(n847) );
  NAND2_X1 U176 ( .A1(\mem[16][12] ), .A2(n1604), .ZN(n318) );
  OAI21_X1 U177 ( .B1(n1575), .B2(n305), .A(n319), .ZN(n848) );
  NAND2_X1 U178 ( .A1(\mem[16][13] ), .A2(n1604), .ZN(n319) );
  OAI21_X1 U179 ( .B1(n1625), .B2(n305), .A(n320), .ZN(n849) );
  NAND2_X1 U180 ( .A1(\mem[16][14] ), .A2(n1604), .ZN(n320) );
  OAI21_X1 U181 ( .B1(n1632), .B2(n1603), .A(n331), .ZN(n858) );
  NAND2_X1 U182 ( .A1(\mem[17][7] ), .A2(n1603), .ZN(n331) );
  OAI21_X1 U183 ( .B1(n1580), .B2(n1603), .A(n332), .ZN(n859) );
  NAND2_X1 U184 ( .A1(\mem[17][8] ), .A2(n323), .ZN(n332) );
  OAI21_X1 U185 ( .B1(n1630), .B2(n1603), .A(n333), .ZN(n860) );
  NAND2_X1 U186 ( .A1(\mem[17][9] ), .A2(n323), .ZN(n333) );
  OAI21_X1 U187 ( .B1(n1629), .B2(n1603), .A(n334), .ZN(n861) );
  NAND2_X1 U188 ( .A1(\mem[17][10] ), .A2(n323), .ZN(n334) );
  OAI21_X1 U189 ( .B1(n1628), .B2(n1603), .A(n335), .ZN(n862) );
  NAND2_X1 U190 ( .A1(\mem[17][11] ), .A2(n323), .ZN(n335) );
  OAI21_X1 U191 ( .B1(n1627), .B2(n1603), .A(n336), .ZN(n863) );
  NAND2_X1 U192 ( .A1(\mem[17][12] ), .A2(n323), .ZN(n336) );
  OAI21_X1 U193 ( .B1(n1575), .B2(n1603), .A(n337), .ZN(n864) );
  NAND2_X1 U194 ( .A1(\mem[17][13] ), .A2(n323), .ZN(n337) );
  OAI21_X1 U195 ( .B1(n1625), .B2(n1603), .A(n338), .ZN(n865) );
  NAND2_X1 U196 ( .A1(\mem[17][14] ), .A2(n323), .ZN(n338) );
  OAI21_X1 U197 ( .B1(n1632), .B2(n340), .A(n348), .ZN(n874) );
  NAND2_X1 U198 ( .A1(\mem[18][7] ), .A2(n1602), .ZN(n348) );
  OAI21_X1 U199 ( .B1(n1580), .B2(n1602), .A(n349), .ZN(n875) );
  NAND2_X1 U200 ( .A1(\mem[18][8] ), .A2(n1602), .ZN(n349) );
  OAI21_X1 U201 ( .B1(n1630), .B2(n340), .A(n350), .ZN(n876) );
  NAND2_X1 U202 ( .A1(\mem[18][9] ), .A2(n1602), .ZN(n350) );
  OAI21_X1 U203 ( .B1(n1629), .B2(n340), .A(n351), .ZN(n877) );
  NAND2_X1 U204 ( .A1(\mem[18][10] ), .A2(n1602), .ZN(n351) );
  OAI21_X1 U205 ( .B1(n1628), .B2(n340), .A(n352), .ZN(n878) );
  NAND2_X1 U206 ( .A1(\mem[18][11] ), .A2(n1602), .ZN(n352) );
  OAI21_X1 U207 ( .B1(n1627), .B2(n340), .A(n353), .ZN(n879) );
  NAND2_X1 U208 ( .A1(\mem[18][12] ), .A2(n1602), .ZN(n353) );
  OAI21_X1 U209 ( .B1(n1575), .B2(n340), .A(n354), .ZN(n880) );
  NAND2_X1 U210 ( .A1(\mem[18][13] ), .A2(n1602), .ZN(n354) );
  OAI21_X1 U211 ( .B1(n1625), .B2(n340), .A(n355), .ZN(n881) );
  NAND2_X1 U212 ( .A1(\mem[18][14] ), .A2(n1602), .ZN(n355) );
  OAI21_X1 U213 ( .B1(n1632), .B2(n357), .A(n365), .ZN(n890) );
  NAND2_X1 U214 ( .A1(\mem[19][7] ), .A2(n1601), .ZN(n365) );
  OAI21_X1 U215 ( .B1(n1580), .B2(n1601), .A(n366), .ZN(n891) );
  NAND2_X1 U216 ( .A1(\mem[19][8] ), .A2(n1601), .ZN(n366) );
  OAI21_X1 U217 ( .B1(n1630), .B2(n357), .A(n367), .ZN(n892) );
  NAND2_X1 U218 ( .A1(\mem[19][9] ), .A2(n1601), .ZN(n367) );
  OAI21_X1 U219 ( .B1(n1629), .B2(n357), .A(n368), .ZN(n893) );
  NAND2_X1 U220 ( .A1(\mem[19][10] ), .A2(n1601), .ZN(n368) );
  OAI21_X1 U221 ( .B1(n1628), .B2(n357), .A(n369), .ZN(n894) );
  NAND2_X1 U222 ( .A1(\mem[19][11] ), .A2(n1601), .ZN(n369) );
  OAI21_X1 U223 ( .B1(n1627), .B2(n357), .A(n370), .ZN(n895) );
  NAND2_X1 U224 ( .A1(\mem[19][12] ), .A2(n1601), .ZN(n370) );
  OAI21_X1 U225 ( .B1(n1575), .B2(n357), .A(n371), .ZN(n896) );
  NAND2_X1 U226 ( .A1(\mem[19][13] ), .A2(n1601), .ZN(n371) );
  OAI21_X1 U227 ( .B1(n1625), .B2(n357), .A(n372), .ZN(n897) );
  NAND2_X1 U228 ( .A1(\mem[19][14] ), .A2(n1601), .ZN(n372) );
  OAI21_X1 U229 ( .B1(n1632), .B2(n442), .A(n450), .ZN(n970) );
  NAND2_X1 U230 ( .A1(\mem[24][7] ), .A2(n1596), .ZN(n450) );
  OAI21_X1 U231 ( .B1(n1580), .B2(n442), .A(n451), .ZN(n971) );
  NAND2_X1 U232 ( .A1(\mem[24][8] ), .A2(n1596), .ZN(n451) );
  OAI21_X1 U233 ( .B1(n1630), .B2(n442), .A(n452), .ZN(n972) );
  NAND2_X1 U234 ( .A1(\mem[24][9] ), .A2(n442), .ZN(n452) );
  OAI21_X1 U235 ( .B1(n1629), .B2(n442), .A(n453), .ZN(n973) );
  NAND2_X1 U236 ( .A1(\mem[24][10] ), .A2(n442), .ZN(n453) );
  OAI21_X1 U237 ( .B1(n1628), .B2(n442), .A(n454), .ZN(n974) );
  NAND2_X1 U238 ( .A1(\mem[24][11] ), .A2(n442), .ZN(n454) );
  OAI21_X1 U239 ( .B1(n1627), .B2(n442), .A(n455), .ZN(n975) );
  NAND2_X1 U240 ( .A1(\mem[24][12] ), .A2(n1596), .ZN(n455) );
  OAI21_X1 U241 ( .B1(n1575), .B2(n442), .A(n456), .ZN(n976) );
  NAND2_X1 U242 ( .A1(\mem[24][13] ), .A2(n442), .ZN(n456) );
  OAI21_X1 U243 ( .B1(n1625), .B2(n442), .A(n457), .ZN(n977) );
  NAND2_X1 U244 ( .A1(\mem[24][14] ), .A2(n442), .ZN(n457) );
  OAI21_X1 U245 ( .B1(n1632), .B2(n460), .A(n468), .ZN(n986) );
  NAND2_X1 U246 ( .A1(\mem[25][7] ), .A2(n1595), .ZN(n468) );
  OAI21_X1 U247 ( .B1(n1580), .B2(n1595), .A(n469), .ZN(n987) );
  NAND2_X1 U248 ( .A1(\mem[25][8] ), .A2(n1595), .ZN(n469) );
  OAI21_X1 U249 ( .B1(n1630), .B2(n460), .A(n470), .ZN(n988) );
  NAND2_X1 U250 ( .A1(\mem[25][9] ), .A2(n1595), .ZN(n470) );
  OAI21_X1 U251 ( .B1(n1629), .B2(n460), .A(n471), .ZN(n989) );
  NAND2_X1 U252 ( .A1(\mem[25][10] ), .A2(n1595), .ZN(n471) );
  OAI21_X1 U253 ( .B1(n1628), .B2(n460), .A(n472), .ZN(n990) );
  NAND2_X1 U254 ( .A1(\mem[25][11] ), .A2(n1595), .ZN(n472) );
  OAI21_X1 U255 ( .B1(n1627), .B2(n460), .A(n473), .ZN(n991) );
  NAND2_X1 U256 ( .A1(\mem[25][12] ), .A2(n1595), .ZN(n473) );
  OAI21_X1 U257 ( .B1(n1575), .B2(n460), .A(n474), .ZN(n992) );
  NAND2_X1 U258 ( .A1(\mem[25][13] ), .A2(n1595), .ZN(n474) );
  OAI21_X1 U259 ( .B1(n1625), .B2(n460), .A(n475), .ZN(n993) );
  NAND2_X1 U260 ( .A1(\mem[25][14] ), .A2(n1595), .ZN(n475) );
  OAI21_X1 U261 ( .B1(n1632), .B2(n477), .A(n485), .ZN(n1002) );
  NAND2_X1 U262 ( .A1(\mem[26][7] ), .A2(n1594), .ZN(n485) );
  OAI21_X1 U263 ( .B1(n1631), .B2(n1594), .A(n486), .ZN(n1003) );
  NAND2_X1 U264 ( .A1(\mem[26][8] ), .A2(n1594), .ZN(n486) );
  OAI21_X1 U265 ( .B1(n1630), .B2(n477), .A(n487), .ZN(n1004) );
  NAND2_X1 U266 ( .A1(\mem[26][9] ), .A2(n1594), .ZN(n487) );
  OAI21_X1 U267 ( .B1(n1629), .B2(n477), .A(n488), .ZN(n1005) );
  NAND2_X1 U268 ( .A1(\mem[26][10] ), .A2(n1594), .ZN(n488) );
  OAI21_X1 U269 ( .B1(n1628), .B2(n477), .A(n489), .ZN(n1006) );
  NAND2_X1 U270 ( .A1(\mem[26][11] ), .A2(n1594), .ZN(n489) );
  OAI21_X1 U271 ( .B1(n1627), .B2(n477), .A(n490), .ZN(n1007) );
  NAND2_X1 U272 ( .A1(\mem[26][12] ), .A2(n1594), .ZN(n490) );
  OAI21_X1 U273 ( .B1(n1626), .B2(n477), .A(n491), .ZN(n1008) );
  NAND2_X1 U274 ( .A1(\mem[26][13] ), .A2(n1594), .ZN(n491) );
  OAI21_X1 U275 ( .B1(n1625), .B2(n477), .A(n492), .ZN(n1009) );
  NAND2_X1 U276 ( .A1(\mem[26][14] ), .A2(n1594), .ZN(n492) );
  OAI21_X1 U277 ( .B1(n1632), .B2(n494), .A(n502), .ZN(n1018) );
  NAND2_X1 U278 ( .A1(\mem[27][7] ), .A2(n1593), .ZN(n502) );
  OAI21_X1 U279 ( .B1(n1631), .B2(n1593), .A(n503), .ZN(n1019) );
  NAND2_X1 U280 ( .A1(\mem[27][8] ), .A2(n1593), .ZN(n503) );
  OAI21_X1 U281 ( .B1(n1630), .B2(n494), .A(n504), .ZN(n1020) );
  NAND2_X1 U282 ( .A1(\mem[27][9] ), .A2(n1593), .ZN(n504) );
  OAI21_X1 U283 ( .B1(n1629), .B2(n494), .A(n505), .ZN(n1021) );
  NAND2_X1 U284 ( .A1(\mem[27][10] ), .A2(n1593), .ZN(n505) );
  OAI21_X1 U285 ( .B1(n1628), .B2(n494), .A(n506), .ZN(n1022) );
  NAND2_X1 U286 ( .A1(\mem[27][11] ), .A2(n1593), .ZN(n506) );
  OAI21_X1 U287 ( .B1(n1627), .B2(n494), .A(n507), .ZN(n1023) );
  NAND2_X1 U288 ( .A1(\mem[27][12] ), .A2(n1593), .ZN(n507) );
  OAI21_X1 U289 ( .B1(n1626), .B2(n494), .A(n508), .ZN(n1024) );
  NAND2_X1 U290 ( .A1(\mem[27][13] ), .A2(n1593), .ZN(n508) );
  OAI21_X1 U291 ( .B1(n1625), .B2(n494), .A(n509), .ZN(n1025) );
  NAND2_X1 U292 ( .A1(\mem[27][14] ), .A2(n1593), .ZN(n509) );
  OAI21_X1 U293 ( .B1(n1581), .B2(n95), .A(n103), .ZN(n650) );
  NAND2_X1 U294 ( .A1(\mem[4][7] ), .A2(n95), .ZN(n103) );
  OAI21_X1 U295 ( .B1(n1631), .B2(n95), .A(n104), .ZN(n651) );
  NAND2_X1 U296 ( .A1(\mem[4][8] ), .A2(n1616), .ZN(n104) );
  OAI21_X1 U297 ( .B1(n1579), .B2(n95), .A(n105), .ZN(n652) );
  NAND2_X1 U298 ( .A1(\mem[4][9] ), .A2(n1616), .ZN(n105) );
  OAI21_X1 U299 ( .B1(n1578), .B2(n95), .A(n106), .ZN(n653) );
  NAND2_X1 U300 ( .A1(\mem[4][10] ), .A2(n1616), .ZN(n106) );
  OAI21_X1 U301 ( .B1(n1577), .B2(n95), .A(n107), .ZN(n654) );
  NAND2_X1 U302 ( .A1(\mem[4][11] ), .A2(n1616), .ZN(n107) );
  OAI21_X1 U303 ( .B1(n1576), .B2(n95), .A(n108), .ZN(n655) );
  NAND2_X1 U304 ( .A1(\mem[4][12] ), .A2(n1616), .ZN(n108) );
  OAI21_X1 U305 ( .B1(n1626), .B2(n95), .A(n109), .ZN(n656) );
  NAND2_X1 U306 ( .A1(\mem[4][13] ), .A2(n1616), .ZN(n109) );
  OAI21_X1 U307 ( .B1(n1574), .B2(n95), .A(n110), .ZN(n657) );
  NAND2_X1 U308 ( .A1(\mem[4][14] ), .A2(n1616), .ZN(n110) );
  OAI21_X1 U309 ( .B1(n1581), .B2(n113), .A(n121), .ZN(n666) );
  NAND2_X1 U310 ( .A1(\mem[5][7] ), .A2(n113), .ZN(n121) );
  OAI21_X1 U311 ( .B1(n1631), .B2(n113), .A(n122), .ZN(n667) );
  NAND2_X1 U312 ( .A1(\mem[5][8] ), .A2(n1615), .ZN(n122) );
  OAI21_X1 U313 ( .B1(n1579), .B2(n113), .A(n123), .ZN(n668) );
  NAND2_X1 U314 ( .A1(\mem[5][9] ), .A2(n1615), .ZN(n123) );
  OAI21_X1 U315 ( .B1(n1578), .B2(n113), .A(n124), .ZN(n669) );
  NAND2_X1 U316 ( .A1(\mem[5][10] ), .A2(n1615), .ZN(n124) );
  OAI21_X1 U317 ( .B1(n1577), .B2(n113), .A(n125), .ZN(n670) );
  NAND2_X1 U318 ( .A1(\mem[5][11] ), .A2(n1615), .ZN(n125) );
  OAI21_X1 U319 ( .B1(n1576), .B2(n113), .A(n126), .ZN(n671) );
  NAND2_X1 U320 ( .A1(\mem[5][12] ), .A2(n1615), .ZN(n126) );
  OAI21_X1 U321 ( .B1(n1626), .B2(n113), .A(n127), .ZN(n672) );
  NAND2_X1 U322 ( .A1(\mem[5][13] ), .A2(n1615), .ZN(n127) );
  OAI21_X1 U323 ( .B1(n1574), .B2(n113), .A(n128), .ZN(n673) );
  NAND2_X1 U324 ( .A1(\mem[5][14] ), .A2(n1615), .ZN(n128) );
  OAI21_X1 U325 ( .B1(n1581), .B2(n1614), .A(n139), .ZN(n682) );
  NAND2_X1 U326 ( .A1(\mem[6][7] ), .A2(n1614), .ZN(n139) );
  OAI21_X1 U327 ( .B1(n1631), .B2(n1614), .A(n140), .ZN(n683) );
  NAND2_X1 U328 ( .A1(\mem[6][8] ), .A2(n131), .ZN(n140) );
  OAI21_X1 U329 ( .B1(n1579), .B2(n1614), .A(n141), .ZN(n684) );
  NAND2_X1 U330 ( .A1(\mem[6][9] ), .A2(n131), .ZN(n141) );
  OAI21_X1 U331 ( .B1(n1578), .B2(n1614), .A(n142), .ZN(n685) );
  NAND2_X1 U332 ( .A1(\mem[6][10] ), .A2(n131), .ZN(n142) );
  OAI21_X1 U333 ( .B1(n1577), .B2(n1614), .A(n143), .ZN(n686) );
  NAND2_X1 U334 ( .A1(\mem[6][11] ), .A2(n131), .ZN(n143) );
  OAI21_X1 U335 ( .B1(n1576), .B2(n1614), .A(n144), .ZN(n687) );
  NAND2_X1 U336 ( .A1(\mem[6][12] ), .A2(n131), .ZN(n144) );
  OAI21_X1 U337 ( .B1(n1626), .B2(n1614), .A(n145), .ZN(n688) );
  NAND2_X1 U338 ( .A1(\mem[6][13] ), .A2(n131), .ZN(n145) );
  OAI21_X1 U339 ( .B1(n1574), .B2(n1614), .A(n146), .ZN(n689) );
  NAND2_X1 U340 ( .A1(\mem[6][14] ), .A2(n131), .ZN(n146) );
  OAI21_X1 U341 ( .B1(n1581), .B2(n149), .A(n157), .ZN(n698) );
  NAND2_X1 U342 ( .A1(\mem[7][7] ), .A2(n149), .ZN(n157) );
  OAI21_X1 U343 ( .B1(n1631), .B2(n149), .A(n158), .ZN(n699) );
  NAND2_X1 U344 ( .A1(\mem[7][8] ), .A2(n1613), .ZN(n158) );
  OAI21_X1 U345 ( .B1(n1579), .B2(n149), .A(n159), .ZN(n700) );
  NAND2_X1 U346 ( .A1(\mem[7][9] ), .A2(n1613), .ZN(n159) );
  OAI21_X1 U347 ( .B1(n1578), .B2(n149), .A(n160), .ZN(n701) );
  NAND2_X1 U348 ( .A1(\mem[7][10] ), .A2(n1613), .ZN(n160) );
  OAI21_X1 U349 ( .B1(n1577), .B2(n149), .A(n161), .ZN(n702) );
  NAND2_X1 U350 ( .A1(\mem[7][11] ), .A2(n1613), .ZN(n161) );
  OAI21_X1 U351 ( .B1(n1576), .B2(n149), .A(n162), .ZN(n703) );
  NAND2_X1 U352 ( .A1(\mem[7][12] ), .A2(n1613), .ZN(n162) );
  OAI21_X1 U353 ( .B1(n1626), .B2(n149), .A(n163), .ZN(n704) );
  NAND2_X1 U354 ( .A1(\mem[7][13] ), .A2(n1613), .ZN(n163) );
  OAI21_X1 U355 ( .B1(n1574), .B2(n149), .A(n164), .ZN(n705) );
  NAND2_X1 U356 ( .A1(\mem[7][14] ), .A2(n1613), .ZN(n164) );
  OAI21_X1 U357 ( .B1(n1581), .B2(n237), .A(n245), .ZN(n778) );
  NAND2_X1 U358 ( .A1(\mem[12][7] ), .A2(n237), .ZN(n245) );
  OAI21_X1 U359 ( .B1(n1631), .B2(n237), .A(n246), .ZN(n779) );
  NAND2_X1 U360 ( .A1(\mem[12][8] ), .A2(n1608), .ZN(n246) );
  OAI21_X1 U361 ( .B1(n1579), .B2(n237), .A(n247), .ZN(n780) );
  NAND2_X1 U362 ( .A1(\mem[12][9] ), .A2(n1608), .ZN(n247) );
  OAI21_X1 U363 ( .B1(n1578), .B2(n237), .A(n248), .ZN(n781) );
  NAND2_X1 U364 ( .A1(\mem[12][10] ), .A2(n1608), .ZN(n248) );
  OAI21_X1 U365 ( .B1(n1577), .B2(n237), .A(n249), .ZN(n782) );
  NAND2_X1 U366 ( .A1(\mem[12][11] ), .A2(n1608), .ZN(n249) );
  OAI21_X1 U367 ( .B1(n1576), .B2(n237), .A(n250), .ZN(n783) );
  NAND2_X1 U368 ( .A1(\mem[12][12] ), .A2(n1608), .ZN(n250) );
  OAI21_X1 U369 ( .B1(n1626), .B2(n237), .A(n251), .ZN(n784) );
  NAND2_X1 U370 ( .A1(\mem[12][13] ), .A2(n1608), .ZN(n251) );
  OAI21_X1 U371 ( .B1(n1574), .B2(n237), .A(n252), .ZN(n785) );
  NAND2_X1 U372 ( .A1(\mem[12][14] ), .A2(n1608), .ZN(n252) );
  OAI21_X1 U373 ( .B1(n1632), .B2(n254), .A(n262), .ZN(n794) );
  NAND2_X1 U374 ( .A1(\mem[13][7] ), .A2(n1607), .ZN(n262) );
  OAI21_X1 U375 ( .B1(n1580), .B2(n254), .A(n263), .ZN(n795) );
  NAND2_X1 U376 ( .A1(\mem[13][8] ), .A2(n254), .ZN(n263) );
  OAI21_X1 U377 ( .B1(n1630), .B2(n254), .A(n264), .ZN(n796) );
  NAND2_X1 U378 ( .A1(\mem[13][9] ), .A2(n254), .ZN(n264) );
  OAI21_X1 U379 ( .B1(n1629), .B2(n254), .A(n265), .ZN(n797) );
  NAND2_X1 U380 ( .A1(\mem[13][10] ), .A2(n254), .ZN(n265) );
  OAI21_X1 U381 ( .B1(n1628), .B2(n254), .A(n266), .ZN(n798) );
  NAND2_X1 U382 ( .A1(\mem[13][11] ), .A2(n254), .ZN(n266) );
  OAI21_X1 U383 ( .B1(n1627), .B2(n254), .A(n267), .ZN(n799) );
  NAND2_X1 U384 ( .A1(\mem[13][12] ), .A2(n254), .ZN(n267) );
  OAI21_X1 U385 ( .B1(n1575), .B2(n254), .A(n268), .ZN(n800) );
  NAND2_X1 U386 ( .A1(\mem[13][13] ), .A2(n254), .ZN(n268) );
  OAI21_X1 U387 ( .B1(n1625), .B2(n254), .A(n269), .ZN(n801) );
  NAND2_X1 U388 ( .A1(\mem[13][14] ), .A2(n254), .ZN(n269) );
  OAI21_X1 U389 ( .B1(n1632), .B2(n271), .A(n279), .ZN(n810) );
  NAND2_X1 U390 ( .A1(\mem[14][7] ), .A2(n271), .ZN(n279) );
  OAI21_X1 U391 ( .B1(n1580), .B2(n271), .A(n280), .ZN(n811) );
  NAND2_X1 U392 ( .A1(\mem[14][8] ), .A2(n1606), .ZN(n280) );
  OAI21_X1 U393 ( .B1(n1630), .B2(n271), .A(n281), .ZN(n812) );
  NAND2_X1 U394 ( .A1(\mem[14][9] ), .A2(n1606), .ZN(n281) );
  OAI21_X1 U395 ( .B1(n1629), .B2(n271), .A(n282), .ZN(n813) );
  NAND2_X1 U396 ( .A1(\mem[14][10] ), .A2(n1606), .ZN(n282) );
  OAI21_X1 U397 ( .B1(n1628), .B2(n271), .A(n283), .ZN(n814) );
  NAND2_X1 U398 ( .A1(\mem[14][11] ), .A2(n1606), .ZN(n283) );
  OAI21_X1 U399 ( .B1(n1627), .B2(n271), .A(n284), .ZN(n815) );
  NAND2_X1 U400 ( .A1(\mem[14][12] ), .A2(n1606), .ZN(n284) );
  OAI21_X1 U401 ( .B1(n1575), .B2(n271), .A(n285), .ZN(n816) );
  NAND2_X1 U402 ( .A1(\mem[14][13] ), .A2(n1606), .ZN(n285) );
  OAI21_X1 U403 ( .B1(n1625), .B2(n271), .A(n286), .ZN(n817) );
  NAND2_X1 U404 ( .A1(\mem[14][14] ), .A2(n1606), .ZN(n286) );
  OAI21_X1 U405 ( .B1(n1632), .B2(n288), .A(n296), .ZN(n826) );
  NAND2_X1 U406 ( .A1(\mem[15][7] ), .A2(n288), .ZN(n296) );
  OAI21_X1 U407 ( .B1(n1580), .B2(n288), .A(n297), .ZN(n827) );
  NAND2_X1 U408 ( .A1(\mem[15][8] ), .A2(n1605), .ZN(n297) );
  OAI21_X1 U409 ( .B1(n1630), .B2(n288), .A(n298), .ZN(n828) );
  NAND2_X1 U410 ( .A1(\mem[15][9] ), .A2(n1605), .ZN(n298) );
  OAI21_X1 U411 ( .B1(n1629), .B2(n288), .A(n299), .ZN(n829) );
  NAND2_X1 U412 ( .A1(\mem[15][10] ), .A2(n1605), .ZN(n299) );
  OAI21_X1 U413 ( .B1(n1628), .B2(n288), .A(n300), .ZN(n830) );
  NAND2_X1 U414 ( .A1(\mem[15][11] ), .A2(n1605), .ZN(n300) );
  OAI21_X1 U415 ( .B1(n1627), .B2(n288), .A(n301), .ZN(n831) );
  NAND2_X1 U416 ( .A1(\mem[15][12] ), .A2(n1605), .ZN(n301) );
  OAI21_X1 U417 ( .B1(n1575), .B2(n288), .A(n302), .ZN(n832) );
  NAND2_X1 U418 ( .A1(\mem[15][13] ), .A2(n1605), .ZN(n302) );
  OAI21_X1 U419 ( .B1(n1625), .B2(n288), .A(n303), .ZN(n833) );
  NAND2_X1 U420 ( .A1(\mem[15][14] ), .A2(n1605), .ZN(n303) );
  OAI21_X1 U421 ( .B1(n1632), .B2(n1600), .A(n382), .ZN(n906) );
  NAND2_X1 U422 ( .A1(\mem[20][7] ), .A2(n1600), .ZN(n382) );
  OAI21_X1 U423 ( .B1(n1580), .B2(n1600), .A(n383), .ZN(n907) );
  NAND2_X1 U424 ( .A1(\mem[20][8] ), .A2(n374), .ZN(n383) );
  OAI21_X1 U425 ( .B1(n1630), .B2(n1600), .A(n384), .ZN(n908) );
  NAND2_X1 U426 ( .A1(\mem[20][9] ), .A2(n374), .ZN(n384) );
  OAI21_X1 U427 ( .B1(n1629), .B2(n1600), .A(n385), .ZN(n909) );
  NAND2_X1 U428 ( .A1(\mem[20][10] ), .A2(n374), .ZN(n385) );
  OAI21_X1 U429 ( .B1(n1628), .B2(n1600), .A(n386), .ZN(n910) );
  NAND2_X1 U430 ( .A1(\mem[20][11] ), .A2(n374), .ZN(n386) );
  OAI21_X1 U431 ( .B1(n1627), .B2(n1600), .A(n387), .ZN(n911) );
  NAND2_X1 U432 ( .A1(\mem[20][12] ), .A2(n374), .ZN(n387) );
  OAI21_X1 U433 ( .B1(n1575), .B2(n1600), .A(n388), .ZN(n912) );
  NAND2_X1 U434 ( .A1(\mem[20][13] ), .A2(n374), .ZN(n388) );
  OAI21_X1 U435 ( .B1(n1625), .B2(n1600), .A(n389), .ZN(n913) );
  NAND2_X1 U436 ( .A1(\mem[20][14] ), .A2(n374), .ZN(n389) );
  OAI21_X1 U437 ( .B1(n1632), .B2(n391), .A(n399), .ZN(n922) );
  NAND2_X1 U438 ( .A1(\mem[21][7] ), .A2(n1599), .ZN(n399) );
  OAI21_X1 U439 ( .B1(n1580), .B2(n1599), .A(n400), .ZN(n923) );
  NAND2_X1 U440 ( .A1(\mem[21][8] ), .A2(n1599), .ZN(n400) );
  OAI21_X1 U441 ( .B1(n1630), .B2(n391), .A(n401), .ZN(n924) );
  NAND2_X1 U442 ( .A1(\mem[21][9] ), .A2(n1599), .ZN(n401) );
  OAI21_X1 U443 ( .B1(n1629), .B2(n391), .A(n402), .ZN(n925) );
  NAND2_X1 U444 ( .A1(\mem[21][10] ), .A2(n1599), .ZN(n402) );
  OAI21_X1 U445 ( .B1(n1628), .B2(n391), .A(n403), .ZN(n926) );
  NAND2_X1 U446 ( .A1(\mem[21][11] ), .A2(n1599), .ZN(n403) );
  OAI21_X1 U447 ( .B1(n1627), .B2(n391), .A(n404), .ZN(n927) );
  NAND2_X1 U448 ( .A1(\mem[21][12] ), .A2(n1599), .ZN(n404) );
  OAI21_X1 U449 ( .B1(n1575), .B2(n391), .A(n405), .ZN(n928) );
  NAND2_X1 U450 ( .A1(\mem[21][13] ), .A2(n1599), .ZN(n405) );
  OAI21_X1 U451 ( .B1(n1625), .B2(n391), .A(n406), .ZN(n929) );
  NAND2_X1 U452 ( .A1(\mem[21][14] ), .A2(n1599), .ZN(n406) );
  OAI21_X1 U453 ( .B1(n1632), .B2(n408), .A(n416), .ZN(n938) );
  NAND2_X1 U454 ( .A1(\mem[22][7] ), .A2(n1598), .ZN(n416) );
  OAI21_X1 U455 ( .B1(n1580), .B2(n1598), .A(n417), .ZN(n939) );
  NAND2_X1 U456 ( .A1(\mem[22][8] ), .A2(n1598), .ZN(n417) );
  OAI21_X1 U457 ( .B1(n1630), .B2(n408), .A(n418), .ZN(n940) );
  NAND2_X1 U458 ( .A1(\mem[22][9] ), .A2(n1598), .ZN(n418) );
  OAI21_X1 U459 ( .B1(n1629), .B2(n408), .A(n419), .ZN(n941) );
  NAND2_X1 U460 ( .A1(\mem[22][10] ), .A2(n1598), .ZN(n419) );
  OAI21_X1 U461 ( .B1(n1628), .B2(n408), .A(n420), .ZN(n942) );
  NAND2_X1 U462 ( .A1(\mem[22][11] ), .A2(n1598), .ZN(n420) );
  OAI21_X1 U463 ( .B1(n1627), .B2(n408), .A(n421), .ZN(n943) );
  NAND2_X1 U464 ( .A1(\mem[22][12] ), .A2(n1598), .ZN(n421) );
  OAI21_X1 U465 ( .B1(n1575), .B2(n408), .A(n422), .ZN(n944) );
  NAND2_X1 U466 ( .A1(\mem[22][13] ), .A2(n1598), .ZN(n422) );
  OAI21_X1 U467 ( .B1(n1625), .B2(n408), .A(n423), .ZN(n945) );
  NAND2_X1 U468 ( .A1(\mem[22][14] ), .A2(n1598), .ZN(n423) );
  OAI21_X1 U469 ( .B1(n1632), .B2(n425), .A(n433), .ZN(n954) );
  NAND2_X1 U470 ( .A1(\mem[23][7] ), .A2(n1597), .ZN(n433) );
  OAI21_X1 U471 ( .B1(n1580), .B2(n1597), .A(n434), .ZN(n955) );
  NAND2_X1 U472 ( .A1(\mem[23][8] ), .A2(n1597), .ZN(n434) );
  OAI21_X1 U473 ( .B1(n1630), .B2(n425), .A(n435), .ZN(n956) );
  NAND2_X1 U474 ( .A1(\mem[23][9] ), .A2(n1597), .ZN(n435) );
  OAI21_X1 U475 ( .B1(n1629), .B2(n425), .A(n436), .ZN(n957) );
  NAND2_X1 U476 ( .A1(\mem[23][10] ), .A2(n1597), .ZN(n436) );
  OAI21_X1 U477 ( .B1(n1628), .B2(n425), .A(n437), .ZN(n958) );
  NAND2_X1 U478 ( .A1(\mem[23][11] ), .A2(n1597), .ZN(n437) );
  OAI21_X1 U479 ( .B1(n1627), .B2(n425), .A(n438), .ZN(n959) );
  NAND2_X1 U480 ( .A1(\mem[23][12] ), .A2(n1597), .ZN(n438) );
  OAI21_X1 U481 ( .B1(n1575), .B2(n425), .A(n439), .ZN(n960) );
  NAND2_X1 U482 ( .A1(\mem[23][13] ), .A2(n1597), .ZN(n439) );
  OAI21_X1 U483 ( .B1(n1625), .B2(n425), .A(n440), .ZN(n961) );
  NAND2_X1 U484 ( .A1(\mem[23][14] ), .A2(n1597), .ZN(n440) );
  OAI21_X1 U485 ( .B1(n1632), .B2(n511), .A(n519), .ZN(n1034) );
  NAND2_X1 U486 ( .A1(\mem[28][7] ), .A2(n1592), .ZN(n519) );
  OAI21_X1 U487 ( .B1(n1631), .B2(n1592), .A(n520), .ZN(n1035) );
  NAND2_X1 U488 ( .A1(\mem[28][8] ), .A2(n1592), .ZN(n520) );
  OAI21_X1 U489 ( .B1(n1630), .B2(n511), .A(n521), .ZN(n1036) );
  NAND2_X1 U490 ( .A1(\mem[28][9] ), .A2(n1592), .ZN(n521) );
  OAI21_X1 U491 ( .B1(n1629), .B2(n511), .A(n522), .ZN(n1037) );
  NAND2_X1 U492 ( .A1(\mem[28][10] ), .A2(n1592), .ZN(n522) );
  OAI21_X1 U493 ( .B1(n1628), .B2(n511), .A(n523), .ZN(n1038) );
  NAND2_X1 U494 ( .A1(\mem[28][11] ), .A2(n1592), .ZN(n523) );
  OAI21_X1 U495 ( .B1(n1627), .B2(n511), .A(n524), .ZN(n1039) );
  NAND2_X1 U496 ( .A1(\mem[28][12] ), .A2(n1592), .ZN(n524) );
  OAI21_X1 U497 ( .B1(n1626), .B2(n511), .A(n525), .ZN(n1040) );
  NAND2_X1 U498 ( .A1(\mem[28][13] ), .A2(n1592), .ZN(n525) );
  OAI21_X1 U499 ( .B1(n1625), .B2(n511), .A(n526), .ZN(n1041) );
  NAND2_X1 U500 ( .A1(\mem[28][14] ), .A2(n1592), .ZN(n526) );
  OAI21_X1 U501 ( .B1(n1632), .B2(n528), .A(n536), .ZN(n1050) );
  NAND2_X1 U502 ( .A1(\mem[29][7] ), .A2(n1591), .ZN(n536) );
  OAI21_X1 U503 ( .B1(n1631), .B2(n1591), .A(n537), .ZN(n1051) );
  NAND2_X1 U504 ( .A1(\mem[29][8] ), .A2(n1591), .ZN(n537) );
  OAI21_X1 U505 ( .B1(n1630), .B2(n528), .A(n538), .ZN(n1052) );
  NAND2_X1 U506 ( .A1(\mem[29][9] ), .A2(n1591), .ZN(n538) );
  OAI21_X1 U507 ( .B1(n1629), .B2(n528), .A(n539), .ZN(n1053) );
  NAND2_X1 U508 ( .A1(\mem[29][10] ), .A2(n1591), .ZN(n539) );
  OAI21_X1 U509 ( .B1(n1628), .B2(n528), .A(n540), .ZN(n1054) );
  NAND2_X1 U510 ( .A1(\mem[29][11] ), .A2(n1591), .ZN(n540) );
  OAI21_X1 U511 ( .B1(n1627), .B2(n528), .A(n541), .ZN(n1055) );
  NAND2_X1 U512 ( .A1(\mem[29][12] ), .A2(n1591), .ZN(n541) );
  OAI21_X1 U513 ( .B1(n1626), .B2(n528), .A(n542), .ZN(n1056) );
  NAND2_X1 U514 ( .A1(\mem[29][13] ), .A2(n1591), .ZN(n542) );
  OAI21_X1 U515 ( .B1(n1625), .B2(n528), .A(n543), .ZN(n1057) );
  NAND2_X1 U516 ( .A1(\mem[29][14] ), .A2(n1591), .ZN(n543) );
  OAI21_X1 U517 ( .B1(n1632), .B2(n545), .A(n553), .ZN(n1066) );
  NAND2_X1 U518 ( .A1(\mem[30][7] ), .A2(n1590), .ZN(n553) );
  OAI21_X1 U519 ( .B1(n1631), .B2(n1590), .A(n554), .ZN(n1067) );
  NAND2_X1 U520 ( .A1(\mem[30][8] ), .A2(n1590), .ZN(n554) );
  OAI21_X1 U521 ( .B1(n1630), .B2(n545), .A(n555), .ZN(n1068) );
  NAND2_X1 U522 ( .A1(\mem[30][9] ), .A2(n1590), .ZN(n555) );
  OAI21_X1 U523 ( .B1(n1629), .B2(n545), .A(n556), .ZN(n1069) );
  NAND2_X1 U524 ( .A1(\mem[30][10] ), .A2(n1590), .ZN(n556) );
  OAI21_X1 U525 ( .B1(n1628), .B2(n545), .A(n557), .ZN(n1070) );
  NAND2_X1 U526 ( .A1(\mem[30][11] ), .A2(n1590), .ZN(n557) );
  OAI21_X1 U527 ( .B1(n1627), .B2(n545), .A(n558), .ZN(n1071) );
  NAND2_X1 U528 ( .A1(\mem[30][12] ), .A2(n1590), .ZN(n558) );
  OAI21_X1 U529 ( .B1(n1626), .B2(n545), .A(n559), .ZN(n1072) );
  NAND2_X1 U530 ( .A1(\mem[30][13] ), .A2(n1590), .ZN(n559) );
  OAI21_X1 U531 ( .B1(n1625), .B2(n545), .A(n560), .ZN(n1073) );
  NAND2_X1 U532 ( .A1(\mem[30][14] ), .A2(n1590), .ZN(n560) );
  OAI21_X1 U533 ( .B1(n1632), .B2(n562), .A(n570), .ZN(n1082) );
  NAND2_X1 U534 ( .A1(\mem[31][7] ), .A2(n1589), .ZN(n570) );
  OAI21_X1 U535 ( .B1(n1631), .B2(n1589), .A(n571), .ZN(n1083) );
  NAND2_X1 U536 ( .A1(\mem[31][8] ), .A2(n1589), .ZN(n571) );
  OAI21_X1 U537 ( .B1(n1630), .B2(n562), .A(n572), .ZN(n1084) );
  NAND2_X1 U538 ( .A1(\mem[31][9] ), .A2(n1589), .ZN(n572) );
  OAI21_X1 U539 ( .B1(n1629), .B2(n562), .A(n573), .ZN(n1085) );
  NAND2_X1 U540 ( .A1(\mem[31][10] ), .A2(n1589), .ZN(n573) );
  OAI21_X1 U541 ( .B1(n1628), .B2(n562), .A(n574), .ZN(n1086) );
  NAND2_X1 U542 ( .A1(\mem[31][11] ), .A2(n1589), .ZN(n574) );
  OAI21_X1 U543 ( .B1(n1627), .B2(n562), .A(n575), .ZN(n1087) );
  NAND2_X1 U544 ( .A1(\mem[31][12] ), .A2(n1589), .ZN(n575) );
  OAI21_X1 U545 ( .B1(n1626), .B2(n562), .A(n576), .ZN(n1088) );
  NAND2_X1 U546 ( .A1(\mem[31][13] ), .A2(n1589), .ZN(n576) );
  OAI21_X1 U547 ( .B1(n1625), .B2(n562), .A(n577), .ZN(n1089) );
  NAND2_X1 U548 ( .A1(\mem[31][14] ), .A2(n1589), .ZN(n577) );
  OAI21_X1 U549 ( .B1(n22), .B2(n1631), .A(n31), .ZN(n587) );
  NAND2_X1 U550 ( .A1(\mem[0][8] ), .A2(n22), .ZN(n31) );
  OAI21_X1 U551 ( .B1(n22), .B2(n1579), .A(n32), .ZN(n588) );
  NAND2_X1 U552 ( .A1(\mem[0][9] ), .A2(n22), .ZN(n32) );
  OAI21_X1 U553 ( .B1(n22), .B2(n1578), .A(n33), .ZN(n589) );
  NAND2_X1 U554 ( .A1(\mem[0][10] ), .A2(n22), .ZN(n33) );
  OAI21_X1 U555 ( .B1(n22), .B2(n1577), .A(n34), .ZN(n590) );
  NAND2_X1 U556 ( .A1(\mem[0][11] ), .A2(n22), .ZN(n34) );
  OAI21_X1 U557 ( .B1(n22), .B2(n1576), .A(n35), .ZN(n591) );
  NAND2_X1 U558 ( .A1(\mem[0][12] ), .A2(n22), .ZN(n35) );
  OAI21_X1 U559 ( .B1(n22), .B2(n1626), .A(n36), .ZN(n592) );
  NAND2_X1 U560 ( .A1(\mem[0][13] ), .A2(n22), .ZN(n36) );
  OAI21_X1 U561 ( .B1(n22), .B2(n1574), .A(n37), .ZN(n593) );
  NAND2_X1 U562 ( .A1(\mem[0][14] ), .A2(n22), .ZN(n37) );
  OAI21_X1 U563 ( .B1(n1639), .B2(n477), .A(n478), .ZN(n995) );
  NAND2_X1 U564 ( .A1(\mem[26][0] ), .A2(n1594), .ZN(n478) );
  OAI21_X1 U565 ( .B1(n1624), .B2(n477), .A(n493), .ZN(n1010) );
  NAND2_X1 U566 ( .A1(\mem[26][15] ), .A2(n1594), .ZN(n493) );
  OAI21_X1 U567 ( .B1(n1639), .B2(n494), .A(n495), .ZN(n1011) );
  NAND2_X1 U568 ( .A1(\mem[27][0] ), .A2(n1593), .ZN(n495) );
  OAI21_X1 U569 ( .B1(n1624), .B2(n494), .A(n510), .ZN(n1026) );
  NAND2_X1 U570 ( .A1(\mem[27][15] ), .A2(n1593), .ZN(n510) );
  OAI21_X1 U571 ( .B1(n1639), .B2(n511), .A(n512), .ZN(n1027) );
  NAND2_X1 U572 ( .A1(\mem[28][0] ), .A2(n1592), .ZN(n512) );
  OAI21_X1 U573 ( .B1(n1624), .B2(n511), .A(n527), .ZN(n1042) );
  NAND2_X1 U574 ( .A1(\mem[28][15] ), .A2(n1592), .ZN(n527) );
  OAI21_X1 U575 ( .B1(n1639), .B2(n528), .A(n529), .ZN(n1043) );
  NAND2_X1 U576 ( .A1(\mem[29][0] ), .A2(n1591), .ZN(n529) );
  OAI21_X1 U577 ( .B1(n1624), .B2(n528), .A(n544), .ZN(n1058) );
  NAND2_X1 U578 ( .A1(\mem[29][15] ), .A2(n1591), .ZN(n544) );
  OAI21_X1 U579 ( .B1(n1639), .B2(n545), .A(n546), .ZN(n1059) );
  NAND2_X1 U580 ( .A1(\mem[30][0] ), .A2(n1590), .ZN(n546) );
  OAI21_X1 U581 ( .B1(n1624), .B2(n545), .A(n561), .ZN(n1074) );
  NAND2_X1 U582 ( .A1(\mem[30][15] ), .A2(n1590), .ZN(n561) );
  OAI21_X1 U583 ( .B1(n1639), .B2(n562), .A(n563), .ZN(n1075) );
  NAND2_X1 U584 ( .A1(\mem[31][0] ), .A2(n1589), .ZN(n563) );
  OAI21_X1 U585 ( .B1(n1624), .B2(n562), .A(n578), .ZN(n1090) );
  NAND2_X1 U586 ( .A1(\mem[31][15] ), .A2(n1589), .ZN(n578) );
  OAI21_X1 U587 ( .B1(n1638), .B2(n477), .A(n479), .ZN(n996) );
  NAND2_X1 U588 ( .A1(\mem[26][1] ), .A2(n1594), .ZN(n479) );
  OAI21_X1 U589 ( .B1(n1586), .B2(n477), .A(n480), .ZN(n997) );
  NAND2_X1 U590 ( .A1(\mem[26][2] ), .A2(n1594), .ZN(n480) );
  OAI21_X1 U591 ( .B1(n1636), .B2(n477), .A(n481), .ZN(n998) );
  NAND2_X1 U592 ( .A1(\mem[26][3] ), .A2(n1594), .ZN(n481) );
  OAI21_X1 U593 ( .B1(n1635), .B2(n477), .A(n482), .ZN(n999) );
  NAND2_X1 U594 ( .A1(\mem[26][4] ), .A2(n477), .ZN(n482) );
  OAI21_X1 U595 ( .B1(n1634), .B2(n477), .A(n483), .ZN(n1000) );
  NAND2_X1 U596 ( .A1(\mem[26][5] ), .A2(n477), .ZN(n483) );
  OAI21_X1 U597 ( .B1(n1633), .B2(n477), .A(n484), .ZN(n1001) );
  NAND2_X1 U598 ( .A1(\mem[26][6] ), .A2(n477), .ZN(n484) );
  OAI21_X1 U599 ( .B1(n1638), .B2(n494), .A(n496), .ZN(n1012) );
  NAND2_X1 U600 ( .A1(\mem[27][1] ), .A2(n1593), .ZN(n496) );
  OAI21_X1 U601 ( .B1(n1586), .B2(n494), .A(n497), .ZN(n1013) );
  NAND2_X1 U602 ( .A1(\mem[27][2] ), .A2(n1593), .ZN(n497) );
  OAI21_X1 U603 ( .B1(n1636), .B2(n494), .A(n498), .ZN(n1014) );
  NAND2_X1 U604 ( .A1(\mem[27][3] ), .A2(n1593), .ZN(n498) );
  OAI21_X1 U605 ( .B1(n1635), .B2(n494), .A(n499), .ZN(n1015) );
  NAND2_X1 U606 ( .A1(\mem[27][4] ), .A2(n494), .ZN(n499) );
  OAI21_X1 U607 ( .B1(n1634), .B2(n494), .A(n500), .ZN(n1016) );
  NAND2_X1 U608 ( .A1(\mem[27][5] ), .A2(n494), .ZN(n500) );
  OAI21_X1 U609 ( .B1(n1633), .B2(n494), .A(n501), .ZN(n1017) );
  NAND2_X1 U610 ( .A1(\mem[27][6] ), .A2(n494), .ZN(n501) );
  OAI21_X1 U611 ( .B1(n1638), .B2(n511), .A(n513), .ZN(n1028) );
  NAND2_X1 U612 ( .A1(\mem[28][1] ), .A2(n1592), .ZN(n513) );
  OAI21_X1 U613 ( .B1(n1586), .B2(n511), .A(n514), .ZN(n1029) );
  NAND2_X1 U614 ( .A1(\mem[28][2] ), .A2(n1592), .ZN(n514) );
  OAI21_X1 U615 ( .B1(n1636), .B2(n511), .A(n515), .ZN(n1030) );
  NAND2_X1 U616 ( .A1(\mem[28][3] ), .A2(n1592), .ZN(n515) );
  OAI21_X1 U617 ( .B1(n1635), .B2(n511), .A(n516), .ZN(n1031) );
  NAND2_X1 U618 ( .A1(\mem[28][4] ), .A2(n511), .ZN(n516) );
  OAI21_X1 U619 ( .B1(n1634), .B2(n511), .A(n517), .ZN(n1032) );
  NAND2_X1 U620 ( .A1(\mem[28][5] ), .A2(n511), .ZN(n517) );
  OAI21_X1 U621 ( .B1(n1633), .B2(n511), .A(n518), .ZN(n1033) );
  NAND2_X1 U622 ( .A1(\mem[28][6] ), .A2(n511), .ZN(n518) );
  OAI21_X1 U623 ( .B1(n1638), .B2(n528), .A(n530), .ZN(n1044) );
  NAND2_X1 U624 ( .A1(\mem[29][1] ), .A2(n1591), .ZN(n530) );
  OAI21_X1 U625 ( .B1(n1586), .B2(n528), .A(n531), .ZN(n1045) );
  NAND2_X1 U626 ( .A1(\mem[29][2] ), .A2(n1591), .ZN(n531) );
  OAI21_X1 U627 ( .B1(n1636), .B2(n528), .A(n532), .ZN(n1046) );
  NAND2_X1 U628 ( .A1(\mem[29][3] ), .A2(n1591), .ZN(n532) );
  OAI21_X1 U629 ( .B1(n1635), .B2(n528), .A(n533), .ZN(n1047) );
  NAND2_X1 U630 ( .A1(\mem[29][4] ), .A2(n528), .ZN(n533) );
  OAI21_X1 U631 ( .B1(n1634), .B2(n528), .A(n534), .ZN(n1048) );
  NAND2_X1 U632 ( .A1(\mem[29][5] ), .A2(n528), .ZN(n534) );
  OAI21_X1 U633 ( .B1(n1633), .B2(n528), .A(n535), .ZN(n1049) );
  NAND2_X1 U634 ( .A1(\mem[29][6] ), .A2(n528), .ZN(n535) );
  OAI21_X1 U635 ( .B1(n1638), .B2(n545), .A(n547), .ZN(n1060) );
  NAND2_X1 U636 ( .A1(\mem[30][1] ), .A2(n1590), .ZN(n547) );
  OAI21_X1 U637 ( .B1(n1586), .B2(n545), .A(n548), .ZN(n1061) );
  NAND2_X1 U638 ( .A1(\mem[30][2] ), .A2(n1590), .ZN(n548) );
  OAI21_X1 U639 ( .B1(n1636), .B2(n545), .A(n549), .ZN(n1062) );
  NAND2_X1 U640 ( .A1(\mem[30][3] ), .A2(n1590), .ZN(n549) );
  OAI21_X1 U641 ( .B1(n1635), .B2(n545), .A(n550), .ZN(n1063) );
  NAND2_X1 U642 ( .A1(\mem[30][4] ), .A2(n545), .ZN(n550) );
  OAI21_X1 U643 ( .B1(n1634), .B2(n545), .A(n551), .ZN(n1064) );
  NAND2_X1 U644 ( .A1(\mem[30][5] ), .A2(n545), .ZN(n551) );
  OAI21_X1 U645 ( .B1(n1633), .B2(n545), .A(n552), .ZN(n1065) );
  NAND2_X1 U646 ( .A1(\mem[30][6] ), .A2(n545), .ZN(n552) );
  OAI21_X1 U647 ( .B1(n1638), .B2(n562), .A(n564), .ZN(n1076) );
  NAND2_X1 U648 ( .A1(\mem[31][1] ), .A2(n1589), .ZN(n564) );
  OAI21_X1 U649 ( .B1(n1586), .B2(n562), .A(n565), .ZN(n1077) );
  NAND2_X1 U650 ( .A1(\mem[31][2] ), .A2(n1589), .ZN(n565) );
  OAI21_X1 U651 ( .B1(n1636), .B2(n562), .A(n566), .ZN(n1078) );
  NAND2_X1 U652 ( .A1(\mem[31][3] ), .A2(n1589), .ZN(n566) );
  OAI21_X1 U653 ( .B1(n1635), .B2(n562), .A(n567), .ZN(n1079) );
  NAND2_X1 U654 ( .A1(\mem[31][4] ), .A2(n562), .ZN(n567) );
  OAI21_X1 U655 ( .B1(n1634), .B2(n562), .A(n568), .ZN(n1080) );
  NAND2_X1 U656 ( .A1(\mem[31][5] ), .A2(n562), .ZN(n568) );
  OAI21_X1 U657 ( .B1(n1633), .B2(n562), .A(n569), .ZN(n1081) );
  NAND2_X1 U658 ( .A1(\mem[31][6] ), .A2(n562), .ZN(n569) );
  OAI21_X1 U659 ( .B1(n1620), .B2(n1639), .A(n23), .ZN(n579) );
  NAND2_X1 U660 ( .A1(\mem[0][0] ), .A2(n22), .ZN(n23) );
  OAI21_X1 U661 ( .B1(n1620), .B2(n1587), .A(n24), .ZN(n580) );
  NAND2_X1 U662 ( .A1(\mem[0][1] ), .A2(n22), .ZN(n24) );
  OAI21_X1 U663 ( .B1(n1620), .B2(n1637), .A(n25), .ZN(n581) );
  NAND2_X1 U664 ( .A1(\mem[0][2] ), .A2(n22), .ZN(n25) );
  OAI21_X1 U665 ( .B1(n1620), .B2(n1585), .A(n26), .ZN(n582) );
  NAND2_X1 U666 ( .A1(\mem[0][3] ), .A2(n22), .ZN(n26) );
  OAI21_X1 U667 ( .B1(n1620), .B2(n1584), .A(n27), .ZN(n583) );
  NAND2_X1 U668 ( .A1(\mem[0][4] ), .A2(n1620), .ZN(n27) );
  OAI21_X1 U669 ( .B1(n1620), .B2(n1583), .A(n28), .ZN(n584) );
  NAND2_X1 U670 ( .A1(\mem[0][5] ), .A2(n1620), .ZN(n28) );
  OAI21_X1 U671 ( .B1(n1620), .B2(n1582), .A(n29), .ZN(n585) );
  NAND2_X1 U672 ( .A1(\mem[0][6] ), .A2(n1620), .ZN(n29) );
  OAI21_X1 U673 ( .B1(n1620), .B2(n1581), .A(n30), .ZN(n586) );
  NAND2_X1 U674 ( .A1(\mem[0][7] ), .A2(n1620), .ZN(n30) );
  OAI21_X1 U675 ( .B1(n1620), .B2(n1624), .A(n38), .ZN(n594) );
  NAND2_X1 U676 ( .A1(\mem[0][15] ), .A2(n22), .ZN(n38) );
  OAI21_X1 U677 ( .B1(n1639), .B2(n41), .A(n42), .ZN(n595) );
  NAND2_X1 U678 ( .A1(\mem[1][0] ), .A2(n1619), .ZN(n42) );
  OAI21_X1 U679 ( .B1(n1587), .B2(n41), .A(n43), .ZN(n596) );
  NAND2_X1 U680 ( .A1(\mem[1][1] ), .A2(n1619), .ZN(n43) );
  OAI21_X1 U681 ( .B1(n1637), .B2(n41), .A(n44), .ZN(n597) );
  NAND2_X1 U682 ( .A1(\mem[1][2] ), .A2(n1619), .ZN(n44) );
  OAI21_X1 U683 ( .B1(n1585), .B2(n41), .A(n45), .ZN(n598) );
  NAND2_X1 U684 ( .A1(\mem[1][3] ), .A2(n1619), .ZN(n45) );
  OAI21_X1 U685 ( .B1(n1584), .B2(n41), .A(n46), .ZN(n599) );
  NAND2_X1 U686 ( .A1(\mem[1][4] ), .A2(n41), .ZN(n46) );
  OAI21_X1 U687 ( .B1(n1583), .B2(n41), .A(n47), .ZN(n600) );
  NAND2_X1 U688 ( .A1(\mem[1][5] ), .A2(n41), .ZN(n47) );
  OAI21_X1 U689 ( .B1(n1582), .B2(n41), .A(n48), .ZN(n601) );
  NAND2_X1 U690 ( .A1(\mem[1][6] ), .A2(n41), .ZN(n48) );
  OAI21_X1 U691 ( .B1(n1624), .B2(n41), .A(n57), .ZN(n610) );
  NAND2_X1 U692 ( .A1(\mem[1][15] ), .A2(n1619), .ZN(n57) );
  OAI21_X1 U693 ( .B1(n1639), .B2(n59), .A(n60), .ZN(n611) );
  NAND2_X1 U694 ( .A1(\mem[2][0] ), .A2(n1618), .ZN(n60) );
  OAI21_X1 U695 ( .B1(n1587), .B2(n59), .A(n61), .ZN(n612) );
  NAND2_X1 U696 ( .A1(\mem[2][1] ), .A2(n1618), .ZN(n61) );
  OAI21_X1 U697 ( .B1(n1637), .B2(n59), .A(n62), .ZN(n613) );
  NAND2_X1 U698 ( .A1(\mem[2][2] ), .A2(n1618), .ZN(n62) );
  OAI21_X1 U699 ( .B1(n1585), .B2(n59), .A(n63), .ZN(n614) );
  NAND2_X1 U700 ( .A1(\mem[2][3] ), .A2(n1618), .ZN(n63) );
  OAI21_X1 U701 ( .B1(n1584), .B2(n59), .A(n64), .ZN(n615) );
  NAND2_X1 U702 ( .A1(\mem[2][4] ), .A2(n59), .ZN(n64) );
  OAI21_X1 U703 ( .B1(n1583), .B2(n59), .A(n65), .ZN(n616) );
  NAND2_X1 U704 ( .A1(\mem[2][5] ), .A2(n59), .ZN(n65) );
  OAI21_X1 U705 ( .B1(n1582), .B2(n59), .A(n66), .ZN(n617) );
  NAND2_X1 U706 ( .A1(\mem[2][6] ), .A2(n59), .ZN(n66) );
  OAI21_X1 U707 ( .B1(n1624), .B2(n59), .A(n75), .ZN(n626) );
  NAND2_X1 U708 ( .A1(\mem[2][15] ), .A2(n1618), .ZN(n75) );
  OAI21_X1 U709 ( .B1(n1639), .B2(n77), .A(n78), .ZN(n627) );
  NAND2_X1 U710 ( .A1(\mem[3][0] ), .A2(n1617), .ZN(n78) );
  OAI21_X1 U711 ( .B1(n1587), .B2(n77), .A(n79), .ZN(n628) );
  NAND2_X1 U712 ( .A1(\mem[3][1] ), .A2(n1617), .ZN(n79) );
  OAI21_X1 U713 ( .B1(n1637), .B2(n77), .A(n80), .ZN(n629) );
  NAND2_X1 U714 ( .A1(\mem[3][2] ), .A2(n1617), .ZN(n80) );
  OAI21_X1 U715 ( .B1(n1585), .B2(n77), .A(n81), .ZN(n630) );
  NAND2_X1 U716 ( .A1(\mem[3][3] ), .A2(n1617), .ZN(n81) );
  OAI21_X1 U717 ( .B1(n1584), .B2(n77), .A(n82), .ZN(n631) );
  NAND2_X1 U718 ( .A1(\mem[3][4] ), .A2(n77), .ZN(n82) );
  OAI21_X1 U719 ( .B1(n1583), .B2(n77), .A(n83), .ZN(n632) );
  NAND2_X1 U720 ( .A1(\mem[3][5] ), .A2(n77), .ZN(n83) );
  OAI21_X1 U721 ( .B1(n1582), .B2(n77), .A(n84), .ZN(n633) );
  NAND2_X1 U722 ( .A1(\mem[3][6] ), .A2(n77), .ZN(n84) );
  OAI21_X1 U723 ( .B1(n1624), .B2(n77), .A(n93), .ZN(n642) );
  NAND2_X1 U724 ( .A1(\mem[3][15] ), .A2(n1617), .ZN(n93) );
  OAI21_X1 U725 ( .B1(n1639), .B2(n95), .A(n96), .ZN(n643) );
  NAND2_X1 U726 ( .A1(\mem[4][0] ), .A2(n1616), .ZN(n96) );
  OAI21_X1 U727 ( .B1(n1587), .B2(n95), .A(n97), .ZN(n644) );
  NAND2_X1 U728 ( .A1(\mem[4][1] ), .A2(n1616), .ZN(n97) );
  OAI21_X1 U729 ( .B1(n1637), .B2(n95), .A(n98), .ZN(n645) );
  NAND2_X1 U730 ( .A1(\mem[4][2] ), .A2(n1616), .ZN(n98) );
  OAI21_X1 U731 ( .B1(n1585), .B2(n95), .A(n99), .ZN(n646) );
  NAND2_X1 U732 ( .A1(\mem[4][3] ), .A2(n1616), .ZN(n99) );
  OAI21_X1 U733 ( .B1(n1584), .B2(n95), .A(n100), .ZN(n647) );
  NAND2_X1 U734 ( .A1(\mem[4][4] ), .A2(n95), .ZN(n100) );
  OAI21_X1 U735 ( .B1(n1583), .B2(n95), .A(n101), .ZN(n648) );
  NAND2_X1 U736 ( .A1(\mem[4][5] ), .A2(n95), .ZN(n101) );
  OAI21_X1 U737 ( .B1(n1582), .B2(n95), .A(n102), .ZN(n649) );
  NAND2_X1 U738 ( .A1(\mem[4][6] ), .A2(n95), .ZN(n102) );
  OAI21_X1 U739 ( .B1(n1624), .B2(n95), .A(n111), .ZN(n658) );
  NAND2_X1 U740 ( .A1(\mem[4][15] ), .A2(n1616), .ZN(n111) );
  OAI21_X1 U741 ( .B1(n1639), .B2(n113), .A(n114), .ZN(n659) );
  NAND2_X1 U742 ( .A1(\mem[5][0] ), .A2(n1615), .ZN(n114) );
  OAI21_X1 U743 ( .B1(n1587), .B2(n113), .A(n115), .ZN(n660) );
  NAND2_X1 U744 ( .A1(\mem[5][1] ), .A2(n1615), .ZN(n115) );
  OAI21_X1 U745 ( .B1(n1637), .B2(n113), .A(n116), .ZN(n661) );
  NAND2_X1 U746 ( .A1(\mem[5][2] ), .A2(n1615), .ZN(n116) );
  OAI21_X1 U747 ( .B1(n1585), .B2(n113), .A(n117), .ZN(n662) );
  NAND2_X1 U748 ( .A1(\mem[5][3] ), .A2(n1615), .ZN(n117) );
  OAI21_X1 U749 ( .B1(n1584), .B2(n113), .A(n118), .ZN(n663) );
  NAND2_X1 U750 ( .A1(\mem[5][4] ), .A2(n113), .ZN(n118) );
  OAI21_X1 U751 ( .B1(n1583), .B2(n113), .A(n119), .ZN(n664) );
  NAND2_X1 U752 ( .A1(\mem[5][5] ), .A2(n113), .ZN(n119) );
  OAI21_X1 U753 ( .B1(n1582), .B2(n113), .A(n120), .ZN(n665) );
  NAND2_X1 U754 ( .A1(\mem[5][6] ), .A2(n113), .ZN(n120) );
  OAI21_X1 U755 ( .B1(n1624), .B2(n113), .A(n129), .ZN(n674) );
  NAND2_X1 U756 ( .A1(\mem[5][15] ), .A2(n1615), .ZN(n129) );
  OAI21_X1 U757 ( .B1(n1639), .B2(n1614), .A(n132), .ZN(n675) );
  NAND2_X1 U758 ( .A1(\mem[6][0] ), .A2(n131), .ZN(n132) );
  OAI21_X1 U759 ( .B1(n1587), .B2(n131), .A(n133), .ZN(n676) );
  NAND2_X1 U760 ( .A1(\mem[6][1] ), .A2(n131), .ZN(n133) );
  OAI21_X1 U761 ( .B1(n1637), .B2(n131), .A(n134), .ZN(n677) );
  NAND2_X1 U762 ( .A1(\mem[6][2] ), .A2(n131), .ZN(n134) );
  OAI21_X1 U763 ( .B1(n1585), .B2(n131), .A(n135), .ZN(n678) );
  NAND2_X1 U764 ( .A1(\mem[6][3] ), .A2(n131), .ZN(n135) );
  OAI21_X1 U765 ( .B1(n1584), .B2(n131), .A(n136), .ZN(n679) );
  NAND2_X1 U766 ( .A1(\mem[6][4] ), .A2(n1614), .ZN(n136) );
  OAI21_X1 U767 ( .B1(n1583), .B2(n131), .A(n137), .ZN(n680) );
  NAND2_X1 U768 ( .A1(\mem[6][5] ), .A2(n1614), .ZN(n137) );
  OAI21_X1 U769 ( .B1(n1582), .B2(n131), .A(n138), .ZN(n681) );
  NAND2_X1 U770 ( .A1(\mem[6][6] ), .A2(n1614), .ZN(n138) );
  OAI21_X1 U771 ( .B1(n1624), .B2(n131), .A(n147), .ZN(n690) );
  NAND2_X1 U772 ( .A1(\mem[6][15] ), .A2(n131), .ZN(n147) );
  OAI21_X1 U773 ( .B1(n1639), .B2(n149), .A(n150), .ZN(n691) );
  NAND2_X1 U774 ( .A1(\mem[7][0] ), .A2(n1613), .ZN(n150) );
  OAI21_X1 U775 ( .B1(n1587), .B2(n149), .A(n151), .ZN(n692) );
  NAND2_X1 U776 ( .A1(\mem[7][1] ), .A2(n1613), .ZN(n151) );
  OAI21_X1 U777 ( .B1(n1637), .B2(n149), .A(n152), .ZN(n693) );
  NAND2_X1 U778 ( .A1(\mem[7][2] ), .A2(n1613), .ZN(n152) );
  OAI21_X1 U779 ( .B1(n1585), .B2(n149), .A(n153), .ZN(n694) );
  NAND2_X1 U780 ( .A1(\mem[7][3] ), .A2(n1613), .ZN(n153) );
  OAI21_X1 U781 ( .B1(n1584), .B2(n149), .A(n154), .ZN(n695) );
  NAND2_X1 U782 ( .A1(\mem[7][4] ), .A2(n149), .ZN(n154) );
  OAI21_X1 U783 ( .B1(n1583), .B2(n149), .A(n155), .ZN(n696) );
  NAND2_X1 U784 ( .A1(\mem[7][5] ), .A2(n149), .ZN(n155) );
  OAI21_X1 U785 ( .B1(n1582), .B2(n149), .A(n156), .ZN(n697) );
  NAND2_X1 U786 ( .A1(\mem[7][6] ), .A2(n149), .ZN(n156) );
  OAI21_X1 U787 ( .B1(n1624), .B2(n149), .A(n165), .ZN(n706) );
  NAND2_X1 U788 ( .A1(\mem[7][15] ), .A2(n1613), .ZN(n165) );
  OAI21_X1 U789 ( .B1(n1639), .B2(n237), .A(n238), .ZN(n771) );
  NAND2_X1 U790 ( .A1(\mem[12][0] ), .A2(n1608), .ZN(n238) );
  OAI21_X1 U791 ( .B1(n1587), .B2(n237), .A(n239), .ZN(n772) );
  NAND2_X1 U792 ( .A1(\mem[12][1] ), .A2(n1608), .ZN(n239) );
  OAI21_X1 U793 ( .B1(n1637), .B2(n237), .A(n240), .ZN(n773) );
  NAND2_X1 U794 ( .A1(\mem[12][2] ), .A2(n1608), .ZN(n240) );
  OAI21_X1 U795 ( .B1(n1585), .B2(n237), .A(n241), .ZN(n774) );
  NAND2_X1 U796 ( .A1(\mem[12][3] ), .A2(n1608), .ZN(n241) );
  OAI21_X1 U797 ( .B1(n1584), .B2(n237), .A(n242), .ZN(n775) );
  NAND2_X1 U798 ( .A1(\mem[12][4] ), .A2(n237), .ZN(n242) );
  OAI21_X1 U799 ( .B1(n1583), .B2(n237), .A(n243), .ZN(n776) );
  NAND2_X1 U800 ( .A1(\mem[12][5] ), .A2(n237), .ZN(n243) );
  OAI21_X1 U801 ( .B1(n1582), .B2(n237), .A(n244), .ZN(n777) );
  NAND2_X1 U802 ( .A1(\mem[12][6] ), .A2(n237), .ZN(n244) );
  OAI21_X1 U803 ( .B1(n1624), .B2(n237), .A(n253), .ZN(n786) );
  NAND2_X1 U804 ( .A1(\mem[12][15] ), .A2(n1608), .ZN(n253) );
  OAI21_X1 U805 ( .B1(n1588), .B2(n1607), .A(n255), .ZN(n787) );
  NAND2_X1 U806 ( .A1(\mem[13][0] ), .A2(n254), .ZN(n255) );
  OAI21_X1 U807 ( .B1(n1638), .B2(n1607), .A(n256), .ZN(n788) );
  NAND2_X1 U808 ( .A1(\mem[13][1] ), .A2(n254), .ZN(n256) );
  OAI21_X1 U809 ( .B1(n1586), .B2(n1607), .A(n257), .ZN(n789) );
  NAND2_X1 U810 ( .A1(\mem[13][2] ), .A2(n254), .ZN(n257) );
  OAI21_X1 U811 ( .B1(n1636), .B2(n1607), .A(n258), .ZN(n790) );
  NAND2_X1 U812 ( .A1(\mem[13][3] ), .A2(n254), .ZN(n258) );
  OAI21_X1 U813 ( .B1(n1635), .B2(n1607), .A(n259), .ZN(n791) );
  NAND2_X1 U814 ( .A1(\mem[13][4] ), .A2(n1607), .ZN(n259) );
  OAI21_X1 U815 ( .B1(n1634), .B2(n1607), .A(n260), .ZN(n792) );
  NAND2_X1 U816 ( .A1(\mem[13][5] ), .A2(n1607), .ZN(n260) );
  OAI21_X1 U817 ( .B1(n1633), .B2(n1607), .A(n261), .ZN(n793) );
  NAND2_X1 U818 ( .A1(\mem[13][6] ), .A2(n1607), .ZN(n261) );
  OAI21_X1 U819 ( .B1(n1573), .B2(n1607), .A(n270), .ZN(n802) );
  NAND2_X1 U820 ( .A1(\mem[13][15] ), .A2(n254), .ZN(n270) );
  OAI21_X1 U821 ( .B1(n1588), .B2(n271), .A(n272), .ZN(n803) );
  NAND2_X1 U822 ( .A1(\mem[14][0] ), .A2(n1606), .ZN(n272) );
  OAI21_X1 U823 ( .B1(n1638), .B2(n271), .A(n273), .ZN(n804) );
  NAND2_X1 U824 ( .A1(\mem[14][1] ), .A2(n1606), .ZN(n273) );
  OAI21_X1 U825 ( .B1(n1586), .B2(n271), .A(n274), .ZN(n805) );
  NAND2_X1 U826 ( .A1(\mem[14][2] ), .A2(n1606), .ZN(n274) );
  OAI21_X1 U827 ( .B1(n1636), .B2(n271), .A(n275), .ZN(n806) );
  NAND2_X1 U828 ( .A1(\mem[14][3] ), .A2(n1606), .ZN(n275) );
  OAI21_X1 U829 ( .B1(n1635), .B2(n271), .A(n276), .ZN(n807) );
  NAND2_X1 U830 ( .A1(\mem[14][4] ), .A2(n271), .ZN(n276) );
  OAI21_X1 U831 ( .B1(n1634), .B2(n271), .A(n277), .ZN(n808) );
  NAND2_X1 U832 ( .A1(\mem[14][5] ), .A2(n271), .ZN(n277) );
  OAI21_X1 U833 ( .B1(n1633), .B2(n271), .A(n278), .ZN(n809) );
  NAND2_X1 U834 ( .A1(\mem[14][6] ), .A2(n271), .ZN(n278) );
  OAI21_X1 U835 ( .B1(n1573), .B2(n271), .A(n287), .ZN(n818) );
  NAND2_X1 U836 ( .A1(\mem[14][15] ), .A2(n1606), .ZN(n287) );
  OAI21_X1 U837 ( .B1(n1588), .B2(n288), .A(n289), .ZN(n819) );
  NAND2_X1 U838 ( .A1(\mem[15][0] ), .A2(n1605), .ZN(n289) );
  OAI21_X1 U839 ( .B1(n1638), .B2(n288), .A(n290), .ZN(n820) );
  NAND2_X1 U840 ( .A1(\mem[15][1] ), .A2(n1605), .ZN(n290) );
  OAI21_X1 U841 ( .B1(n1586), .B2(n288), .A(n291), .ZN(n821) );
  NAND2_X1 U842 ( .A1(\mem[15][2] ), .A2(n1605), .ZN(n291) );
  OAI21_X1 U843 ( .B1(n1636), .B2(n288), .A(n292), .ZN(n822) );
  NAND2_X1 U844 ( .A1(\mem[15][3] ), .A2(n1605), .ZN(n292) );
  OAI21_X1 U845 ( .B1(n1635), .B2(n288), .A(n293), .ZN(n823) );
  NAND2_X1 U846 ( .A1(\mem[15][4] ), .A2(n288), .ZN(n293) );
  OAI21_X1 U847 ( .B1(n1634), .B2(n288), .A(n294), .ZN(n824) );
  NAND2_X1 U848 ( .A1(\mem[15][5] ), .A2(n288), .ZN(n294) );
  OAI21_X1 U849 ( .B1(n1633), .B2(n288), .A(n295), .ZN(n825) );
  NAND2_X1 U850 ( .A1(\mem[15][6] ), .A2(n288), .ZN(n295) );
  OAI21_X1 U851 ( .B1(n1573), .B2(n288), .A(n304), .ZN(n834) );
  NAND2_X1 U852 ( .A1(\mem[15][15] ), .A2(n1605), .ZN(n304) );
  OAI21_X1 U853 ( .B1(n1588), .B2(n305), .A(n306), .ZN(n835) );
  NAND2_X1 U854 ( .A1(\mem[16][0] ), .A2(n1604), .ZN(n306) );
  OAI21_X1 U855 ( .B1(n1638), .B2(n305), .A(n307), .ZN(n836) );
  NAND2_X1 U856 ( .A1(\mem[16][1] ), .A2(n1604), .ZN(n307) );
  OAI21_X1 U857 ( .B1(n1586), .B2(n305), .A(n308), .ZN(n837) );
  NAND2_X1 U858 ( .A1(\mem[16][2] ), .A2(n1604), .ZN(n308) );
  OAI21_X1 U859 ( .B1(n1636), .B2(n305), .A(n309), .ZN(n838) );
  NAND2_X1 U860 ( .A1(\mem[16][3] ), .A2(n1604), .ZN(n309) );
  OAI21_X1 U861 ( .B1(n1635), .B2(n305), .A(n310), .ZN(n839) );
  NAND2_X1 U862 ( .A1(\mem[16][4] ), .A2(n305), .ZN(n310) );
  OAI21_X1 U863 ( .B1(n1634), .B2(n305), .A(n311), .ZN(n840) );
  NAND2_X1 U864 ( .A1(\mem[16][5] ), .A2(n305), .ZN(n311) );
  OAI21_X1 U865 ( .B1(n1633), .B2(n305), .A(n312), .ZN(n841) );
  NAND2_X1 U866 ( .A1(\mem[16][6] ), .A2(n305), .ZN(n312) );
  OAI21_X1 U867 ( .B1(n1573), .B2(n305), .A(n321), .ZN(n850) );
  NAND2_X1 U868 ( .A1(\mem[16][15] ), .A2(n1604), .ZN(n321) );
  OAI21_X1 U869 ( .B1(n1588), .B2(n323), .A(n324), .ZN(n851) );
  NAND2_X1 U870 ( .A1(\mem[17][0] ), .A2(n1603), .ZN(n324) );
  OAI21_X1 U871 ( .B1(n1638), .B2(n323), .A(n325), .ZN(n852) );
  NAND2_X1 U872 ( .A1(\mem[17][1] ), .A2(n323), .ZN(n325) );
  OAI21_X1 U873 ( .B1(n1586), .B2(n1603), .A(n326), .ZN(n853) );
  NAND2_X1 U874 ( .A1(\mem[17][2] ), .A2(n323), .ZN(n326) );
  OAI21_X1 U875 ( .B1(n1636), .B2(n323), .A(n327), .ZN(n854) );
  NAND2_X1 U876 ( .A1(\mem[17][3] ), .A2(n323), .ZN(n327) );
  OAI21_X1 U877 ( .B1(n1635), .B2(n323), .A(n328), .ZN(n855) );
  NAND2_X1 U878 ( .A1(\mem[17][4] ), .A2(n1603), .ZN(n328) );
  OAI21_X1 U879 ( .B1(n1634), .B2(n323), .A(n329), .ZN(n856) );
  NAND2_X1 U880 ( .A1(\mem[17][5] ), .A2(n1603), .ZN(n329) );
  OAI21_X1 U881 ( .B1(n1633), .B2(n323), .A(n330), .ZN(n857) );
  NAND2_X1 U882 ( .A1(\mem[17][6] ), .A2(n1603), .ZN(n330) );
  OAI21_X1 U883 ( .B1(n1573), .B2(n323), .A(n339), .ZN(n866) );
  NAND2_X1 U884 ( .A1(\mem[17][15] ), .A2(n323), .ZN(n339) );
  OAI21_X1 U885 ( .B1(n1588), .B2(n340), .A(n341), .ZN(n867) );
  NAND2_X1 U886 ( .A1(\mem[18][0] ), .A2(n1602), .ZN(n341) );
  OAI21_X1 U887 ( .B1(n1638), .B2(n340), .A(n342), .ZN(n868) );
  NAND2_X1 U888 ( .A1(\mem[18][1] ), .A2(n1602), .ZN(n342) );
  OAI21_X1 U889 ( .B1(n1586), .B2(n340), .A(n343), .ZN(n869) );
  NAND2_X1 U890 ( .A1(\mem[18][2] ), .A2(n1602), .ZN(n343) );
  OAI21_X1 U891 ( .B1(n1636), .B2(n340), .A(n344), .ZN(n870) );
  NAND2_X1 U892 ( .A1(\mem[18][3] ), .A2(n1602), .ZN(n344) );
  OAI21_X1 U893 ( .B1(n1635), .B2(n340), .A(n345), .ZN(n871) );
  NAND2_X1 U894 ( .A1(\mem[18][4] ), .A2(n340), .ZN(n345) );
  OAI21_X1 U895 ( .B1(n1634), .B2(n340), .A(n346), .ZN(n872) );
  NAND2_X1 U896 ( .A1(\mem[18][5] ), .A2(n340), .ZN(n346) );
  OAI21_X1 U897 ( .B1(n1633), .B2(n340), .A(n347), .ZN(n873) );
  NAND2_X1 U898 ( .A1(\mem[18][6] ), .A2(n340), .ZN(n347) );
  OAI21_X1 U899 ( .B1(n1573), .B2(n340), .A(n356), .ZN(n882) );
  NAND2_X1 U900 ( .A1(\mem[18][15] ), .A2(n1602), .ZN(n356) );
  OAI21_X1 U901 ( .B1(n1588), .B2(n357), .A(n358), .ZN(n883) );
  NAND2_X1 U902 ( .A1(\mem[19][0] ), .A2(n1601), .ZN(n358) );
  OAI21_X1 U903 ( .B1(n1638), .B2(n357), .A(n359), .ZN(n884) );
  NAND2_X1 U904 ( .A1(\mem[19][1] ), .A2(n1601), .ZN(n359) );
  OAI21_X1 U905 ( .B1(n1586), .B2(n357), .A(n360), .ZN(n885) );
  NAND2_X1 U906 ( .A1(\mem[19][2] ), .A2(n1601), .ZN(n360) );
  OAI21_X1 U907 ( .B1(n1636), .B2(n357), .A(n361), .ZN(n886) );
  NAND2_X1 U908 ( .A1(\mem[19][3] ), .A2(n1601), .ZN(n361) );
  OAI21_X1 U909 ( .B1(n1635), .B2(n357), .A(n362), .ZN(n887) );
  NAND2_X1 U910 ( .A1(\mem[19][4] ), .A2(n357), .ZN(n362) );
  OAI21_X1 U911 ( .B1(n1634), .B2(n357), .A(n363), .ZN(n888) );
  NAND2_X1 U912 ( .A1(\mem[19][5] ), .A2(n357), .ZN(n363) );
  OAI21_X1 U913 ( .B1(n1633), .B2(n357), .A(n364), .ZN(n889) );
  NAND2_X1 U914 ( .A1(\mem[19][6] ), .A2(n357), .ZN(n364) );
  OAI21_X1 U915 ( .B1(n1573), .B2(n357), .A(n373), .ZN(n898) );
  NAND2_X1 U916 ( .A1(\mem[19][15] ), .A2(n1601), .ZN(n373) );
  OAI21_X1 U917 ( .B1(n1588), .B2(n374), .A(n375), .ZN(n899) );
  NAND2_X1 U918 ( .A1(\mem[20][0] ), .A2(n1600), .ZN(n375) );
  OAI21_X1 U919 ( .B1(n1638), .B2(n374), .A(n376), .ZN(n900) );
  NAND2_X1 U920 ( .A1(\mem[20][1] ), .A2(n374), .ZN(n376) );
  OAI21_X1 U921 ( .B1(n1586), .B2(n1600), .A(n377), .ZN(n901) );
  NAND2_X1 U922 ( .A1(\mem[20][2] ), .A2(n374), .ZN(n377) );
  OAI21_X1 U923 ( .B1(n1636), .B2(n374), .A(n378), .ZN(n902) );
  NAND2_X1 U924 ( .A1(\mem[20][3] ), .A2(n374), .ZN(n378) );
  OAI21_X1 U925 ( .B1(n1635), .B2(n374), .A(n379), .ZN(n903) );
  NAND2_X1 U926 ( .A1(\mem[20][4] ), .A2(n1600), .ZN(n379) );
  OAI21_X1 U927 ( .B1(n1634), .B2(n374), .A(n380), .ZN(n904) );
  NAND2_X1 U928 ( .A1(\mem[20][5] ), .A2(n1600), .ZN(n380) );
  OAI21_X1 U929 ( .B1(n1633), .B2(n374), .A(n381), .ZN(n905) );
  NAND2_X1 U930 ( .A1(\mem[20][6] ), .A2(n1600), .ZN(n381) );
  OAI21_X1 U931 ( .B1(n1573), .B2(n374), .A(n390), .ZN(n914) );
  NAND2_X1 U932 ( .A1(\mem[20][15] ), .A2(n374), .ZN(n390) );
  OAI21_X1 U933 ( .B1(n1588), .B2(n391), .A(n392), .ZN(n915) );
  NAND2_X1 U934 ( .A1(\mem[21][0] ), .A2(n1599), .ZN(n392) );
  OAI21_X1 U935 ( .B1(n1638), .B2(n391), .A(n393), .ZN(n916) );
  NAND2_X1 U936 ( .A1(\mem[21][1] ), .A2(n1599), .ZN(n393) );
  OAI21_X1 U937 ( .B1(n1637), .B2(n391), .A(n394), .ZN(n917) );
  NAND2_X1 U938 ( .A1(\mem[21][2] ), .A2(n1599), .ZN(n394) );
  OAI21_X1 U939 ( .B1(n1636), .B2(n391), .A(n395), .ZN(n918) );
  NAND2_X1 U940 ( .A1(\mem[21][3] ), .A2(n1599), .ZN(n395) );
  OAI21_X1 U941 ( .B1(n1635), .B2(n391), .A(n396), .ZN(n919) );
  NAND2_X1 U942 ( .A1(\mem[21][4] ), .A2(n391), .ZN(n396) );
  OAI21_X1 U943 ( .B1(n1634), .B2(n391), .A(n397), .ZN(n920) );
  NAND2_X1 U944 ( .A1(\mem[21][5] ), .A2(n391), .ZN(n397) );
  OAI21_X1 U945 ( .B1(n1633), .B2(n391), .A(n398), .ZN(n921) );
  NAND2_X1 U946 ( .A1(\mem[21][6] ), .A2(n391), .ZN(n398) );
  OAI21_X1 U947 ( .B1(n1573), .B2(n391), .A(n407), .ZN(n930) );
  NAND2_X1 U948 ( .A1(\mem[21][15] ), .A2(n1599), .ZN(n407) );
  OAI21_X1 U949 ( .B1(n1588), .B2(n408), .A(n409), .ZN(n931) );
  NAND2_X1 U950 ( .A1(\mem[22][0] ), .A2(n1598), .ZN(n409) );
  OAI21_X1 U951 ( .B1(n1638), .B2(n408), .A(n410), .ZN(n932) );
  NAND2_X1 U952 ( .A1(\mem[22][1] ), .A2(n1598), .ZN(n410) );
  OAI21_X1 U953 ( .B1(n1637), .B2(n408), .A(n411), .ZN(n933) );
  NAND2_X1 U954 ( .A1(\mem[22][2] ), .A2(n1598), .ZN(n411) );
  OAI21_X1 U955 ( .B1(n1636), .B2(n408), .A(n412), .ZN(n934) );
  NAND2_X1 U956 ( .A1(\mem[22][3] ), .A2(n1598), .ZN(n412) );
  OAI21_X1 U957 ( .B1(n1635), .B2(n408), .A(n413), .ZN(n935) );
  NAND2_X1 U958 ( .A1(\mem[22][4] ), .A2(n408), .ZN(n413) );
  OAI21_X1 U959 ( .B1(n1634), .B2(n408), .A(n414), .ZN(n936) );
  NAND2_X1 U960 ( .A1(\mem[22][5] ), .A2(n408), .ZN(n414) );
  OAI21_X1 U961 ( .B1(n1633), .B2(n408), .A(n415), .ZN(n937) );
  NAND2_X1 U962 ( .A1(\mem[22][6] ), .A2(n408), .ZN(n415) );
  OAI21_X1 U963 ( .B1(n1573), .B2(n408), .A(n424), .ZN(n946) );
  NAND2_X1 U964 ( .A1(\mem[22][15] ), .A2(n1598), .ZN(n424) );
  OAI21_X1 U965 ( .B1(n1588), .B2(n425), .A(n426), .ZN(n947) );
  NAND2_X1 U966 ( .A1(\mem[23][0] ), .A2(n1597), .ZN(n426) );
  OAI21_X1 U967 ( .B1(n1638), .B2(n425), .A(n427), .ZN(n948) );
  NAND2_X1 U968 ( .A1(\mem[23][1] ), .A2(n1597), .ZN(n427) );
  OAI21_X1 U969 ( .B1(n1637), .B2(n425), .A(n428), .ZN(n949) );
  NAND2_X1 U970 ( .A1(\mem[23][2] ), .A2(n1597), .ZN(n428) );
  OAI21_X1 U971 ( .B1(n1636), .B2(n425), .A(n429), .ZN(n950) );
  NAND2_X1 U972 ( .A1(\mem[23][3] ), .A2(n1597), .ZN(n429) );
  OAI21_X1 U973 ( .B1(n1635), .B2(n425), .A(n430), .ZN(n951) );
  NAND2_X1 U974 ( .A1(\mem[23][4] ), .A2(n425), .ZN(n430) );
  OAI21_X1 U975 ( .B1(n1634), .B2(n425), .A(n431), .ZN(n952) );
  NAND2_X1 U976 ( .A1(\mem[23][5] ), .A2(n425), .ZN(n431) );
  OAI21_X1 U977 ( .B1(n1633), .B2(n425), .A(n432), .ZN(n953) );
  NAND2_X1 U978 ( .A1(\mem[23][6] ), .A2(n425), .ZN(n432) );
  OAI21_X1 U979 ( .B1(n1573), .B2(n425), .A(n441), .ZN(n962) );
  NAND2_X1 U980 ( .A1(\mem[23][15] ), .A2(n1597), .ZN(n441) );
  OAI21_X1 U981 ( .B1(n1588), .B2(n1596), .A(n443), .ZN(n963) );
  NAND2_X1 U982 ( .A1(\mem[24][0] ), .A2(n442), .ZN(n443) );
  OAI21_X1 U983 ( .B1(n1638), .B2(n1596), .A(n444), .ZN(n964) );
  NAND2_X1 U984 ( .A1(\mem[24][1] ), .A2(n442), .ZN(n444) );
  OAI21_X1 U985 ( .B1(n1637), .B2(n1596), .A(n445), .ZN(n965) );
  NAND2_X1 U986 ( .A1(\mem[24][2] ), .A2(n442), .ZN(n445) );
  OAI21_X1 U987 ( .B1(n1636), .B2(n1596), .A(n446), .ZN(n966) );
  NAND2_X1 U988 ( .A1(\mem[24][3] ), .A2(n442), .ZN(n446) );
  OAI21_X1 U989 ( .B1(n1635), .B2(n1596), .A(n447), .ZN(n967) );
  NAND2_X1 U990 ( .A1(\mem[24][4] ), .A2(n1596), .ZN(n447) );
  OAI21_X1 U991 ( .B1(n1634), .B2(n1596), .A(n448), .ZN(n968) );
  NAND2_X1 U992 ( .A1(\mem[24][5] ), .A2(n1596), .ZN(n448) );
  OAI21_X1 U993 ( .B1(n1633), .B2(n1596), .A(n449), .ZN(n969) );
  NAND2_X1 U994 ( .A1(\mem[24][6] ), .A2(n1596), .ZN(n449) );
  OAI21_X1 U995 ( .B1(n1573), .B2(n1596), .A(n458), .ZN(n978) );
  NAND2_X1 U996 ( .A1(\mem[24][15] ), .A2(n442), .ZN(n458) );
  OAI21_X1 U997 ( .B1(n1588), .B2(n460), .A(n461), .ZN(n979) );
  NAND2_X1 U998 ( .A1(\mem[25][0] ), .A2(n1595), .ZN(n461) );
  OAI21_X1 U999 ( .B1(n1638), .B2(n460), .A(n462), .ZN(n980) );
  NAND2_X1 U1000 ( .A1(\mem[25][1] ), .A2(n1595), .ZN(n462) );
  OAI21_X1 U1001 ( .B1(n1637), .B2(n460), .A(n463), .ZN(n981) );
  NAND2_X1 U1002 ( .A1(\mem[25][2] ), .A2(n1595), .ZN(n463) );
  OAI21_X1 U1003 ( .B1(n1636), .B2(n460), .A(n464), .ZN(n982) );
  NAND2_X1 U1004 ( .A1(\mem[25][3] ), .A2(n1595), .ZN(n464) );
  OAI21_X1 U1005 ( .B1(n1635), .B2(n460), .A(n465), .ZN(n983) );
  NAND2_X1 U1006 ( .A1(\mem[25][4] ), .A2(n460), .ZN(n465) );
  OAI21_X1 U1007 ( .B1(n1634), .B2(n460), .A(n466), .ZN(n984) );
  NAND2_X1 U1008 ( .A1(\mem[25][5] ), .A2(n460), .ZN(n466) );
  OAI21_X1 U1009 ( .B1(n1633), .B2(n460), .A(n467), .ZN(n985) );
  NAND2_X1 U1010 ( .A1(\mem[25][6] ), .A2(n460), .ZN(n467) );
  OAI21_X1 U1011 ( .B1(n1573), .B2(n460), .A(n476), .ZN(n994) );
  NAND2_X1 U1012 ( .A1(\mem[25][15] ), .A2(n1595), .ZN(n476) );
  OAI21_X1 U1013 ( .B1(n1584), .B2(n168), .A(n173), .ZN(n711) );
  NAND2_X1 U1014 ( .A1(\mem[8][4] ), .A2(n168), .ZN(n173) );
  OAI21_X1 U1015 ( .B1(n1583), .B2(n168), .A(n174), .ZN(n712) );
  NAND2_X1 U1016 ( .A1(\mem[8][5] ), .A2(n168), .ZN(n174) );
  OAI21_X1 U1017 ( .B1(n1582), .B2(n168), .A(n175), .ZN(n713) );
  NAND2_X1 U1018 ( .A1(\mem[8][6] ), .A2(n168), .ZN(n175) );
  OAI21_X1 U1019 ( .B1(n1581), .B2(n168), .A(n176), .ZN(n714) );
  NAND2_X1 U1020 ( .A1(\mem[8][7] ), .A2(n168), .ZN(n176) );
  OAI21_X1 U1021 ( .B1(n1584), .B2(n186), .A(n191), .ZN(n727) );
  NAND2_X1 U1022 ( .A1(\mem[9][4] ), .A2(n186), .ZN(n191) );
  OAI21_X1 U1023 ( .B1(n1583), .B2(n186), .A(n192), .ZN(n728) );
  NAND2_X1 U1024 ( .A1(\mem[9][5] ), .A2(n186), .ZN(n192) );
  OAI21_X1 U1025 ( .B1(n1582), .B2(n186), .A(n193), .ZN(n729) );
  NAND2_X1 U1026 ( .A1(\mem[9][6] ), .A2(n186), .ZN(n193) );
  OAI21_X1 U1027 ( .B1(n1581), .B2(n186), .A(n194), .ZN(n730) );
  NAND2_X1 U1028 ( .A1(\mem[9][7] ), .A2(n186), .ZN(n194) );
  OAI21_X1 U1029 ( .B1(n1584), .B2(n203), .A(n208), .ZN(n743) );
  NAND2_X1 U1030 ( .A1(\mem[10][4] ), .A2(n203), .ZN(n208) );
  OAI21_X1 U1031 ( .B1(n1583), .B2(n203), .A(n209), .ZN(n744) );
  NAND2_X1 U1032 ( .A1(\mem[10][5] ), .A2(n203), .ZN(n209) );
  OAI21_X1 U1033 ( .B1(n1582), .B2(n203), .A(n210), .ZN(n745) );
  NAND2_X1 U1034 ( .A1(\mem[10][6] ), .A2(n203), .ZN(n210) );
  OAI21_X1 U1035 ( .B1(n1581), .B2(n203), .A(n211), .ZN(n746) );
  NAND2_X1 U1036 ( .A1(\mem[10][7] ), .A2(n203), .ZN(n211) );
  OAI21_X1 U1037 ( .B1(n1584), .B2(n1609), .A(n225), .ZN(n759) );
  NAND2_X1 U1038 ( .A1(\mem[11][4] ), .A2(n1609), .ZN(n225) );
  OAI21_X1 U1039 ( .B1(n1583), .B2(n1609), .A(n226), .ZN(n760) );
  NAND2_X1 U1040 ( .A1(\mem[11][5] ), .A2(n1609), .ZN(n226) );
  OAI21_X1 U1041 ( .B1(n1582), .B2(n1609), .A(n227), .ZN(n761) );
  NAND2_X1 U1042 ( .A1(\mem[11][6] ), .A2(n1609), .ZN(n227) );
  OAI21_X1 U1043 ( .B1(n1581), .B2(n220), .A(n228), .ZN(n762) );
  NAND2_X1 U1044 ( .A1(\mem[11][7] ), .A2(n1609), .ZN(n228) );
  OAI21_X1 U1045 ( .B1(n1639), .B2(n168), .A(n169), .ZN(n707) );
  NAND2_X1 U1046 ( .A1(\mem[8][0] ), .A2(n1612), .ZN(n169) );
  OAI21_X1 U1047 ( .B1(n1587), .B2(n168), .A(n170), .ZN(n708) );
  NAND2_X1 U1048 ( .A1(\mem[8][1] ), .A2(n1612), .ZN(n170) );
  OAI21_X1 U1049 ( .B1(n1637), .B2(n168), .A(n171), .ZN(n709) );
  NAND2_X1 U1050 ( .A1(\mem[8][2] ), .A2(n1612), .ZN(n171) );
  OAI21_X1 U1051 ( .B1(n1585), .B2(n168), .A(n172), .ZN(n710) );
  NAND2_X1 U1052 ( .A1(\mem[8][3] ), .A2(n1612), .ZN(n172) );
  OAI21_X1 U1053 ( .B1(n1631), .B2(n168), .A(n177), .ZN(n715) );
  NAND2_X1 U1054 ( .A1(\mem[8][8] ), .A2(n1612), .ZN(n177) );
  OAI21_X1 U1055 ( .B1(n1579), .B2(n168), .A(n178), .ZN(n716) );
  NAND2_X1 U1056 ( .A1(\mem[8][9] ), .A2(n1612), .ZN(n178) );
  OAI21_X1 U1057 ( .B1(n1578), .B2(n168), .A(n179), .ZN(n717) );
  NAND2_X1 U1058 ( .A1(\mem[8][10] ), .A2(n1612), .ZN(n179) );
  OAI21_X1 U1059 ( .B1(n1577), .B2(n168), .A(n180), .ZN(n718) );
  NAND2_X1 U1060 ( .A1(\mem[8][11] ), .A2(n1612), .ZN(n180) );
  OAI21_X1 U1061 ( .B1(n1576), .B2(n168), .A(n181), .ZN(n719) );
  NAND2_X1 U1062 ( .A1(\mem[8][12] ), .A2(n1612), .ZN(n181) );
  OAI21_X1 U1063 ( .B1(n1626), .B2(n168), .A(n182), .ZN(n720) );
  NAND2_X1 U1064 ( .A1(\mem[8][13] ), .A2(n1612), .ZN(n182) );
  OAI21_X1 U1065 ( .B1(n1574), .B2(n168), .A(n183), .ZN(n721) );
  NAND2_X1 U1066 ( .A1(\mem[8][14] ), .A2(n1612), .ZN(n183) );
  OAI21_X1 U1067 ( .B1(n1624), .B2(n168), .A(n184), .ZN(n722) );
  NAND2_X1 U1068 ( .A1(\mem[8][15] ), .A2(n1612), .ZN(n184) );
  OAI21_X1 U1069 ( .B1(n1639), .B2(n186), .A(n187), .ZN(n723) );
  NAND2_X1 U1070 ( .A1(\mem[9][0] ), .A2(n1611), .ZN(n187) );
  OAI21_X1 U1071 ( .B1(n1587), .B2(n186), .A(n188), .ZN(n724) );
  NAND2_X1 U1072 ( .A1(\mem[9][1] ), .A2(n1611), .ZN(n188) );
  OAI21_X1 U1073 ( .B1(n1637), .B2(n186), .A(n189), .ZN(n725) );
  NAND2_X1 U1074 ( .A1(\mem[9][2] ), .A2(n1611), .ZN(n189) );
  OAI21_X1 U1075 ( .B1(n1585), .B2(n186), .A(n190), .ZN(n726) );
  NAND2_X1 U1076 ( .A1(\mem[9][3] ), .A2(n1611), .ZN(n190) );
  OAI21_X1 U1077 ( .B1(n1631), .B2(n186), .A(n195), .ZN(n731) );
  NAND2_X1 U1078 ( .A1(\mem[9][8] ), .A2(n1611), .ZN(n195) );
  OAI21_X1 U1079 ( .B1(n1579), .B2(n186), .A(n196), .ZN(n732) );
  NAND2_X1 U1080 ( .A1(\mem[9][9] ), .A2(n1611), .ZN(n196) );
  OAI21_X1 U1081 ( .B1(n1578), .B2(n186), .A(n197), .ZN(n733) );
  NAND2_X1 U1082 ( .A1(\mem[9][10] ), .A2(n1611), .ZN(n197) );
  OAI21_X1 U1083 ( .B1(n1577), .B2(n186), .A(n198), .ZN(n734) );
  NAND2_X1 U1084 ( .A1(\mem[9][11] ), .A2(n1611), .ZN(n198) );
  OAI21_X1 U1085 ( .B1(n1576), .B2(n186), .A(n199), .ZN(n735) );
  NAND2_X1 U1086 ( .A1(\mem[9][12] ), .A2(n1611), .ZN(n199) );
  OAI21_X1 U1087 ( .B1(n1626), .B2(n186), .A(n200), .ZN(n736) );
  NAND2_X1 U1088 ( .A1(\mem[9][13] ), .A2(n1611), .ZN(n200) );
  OAI21_X1 U1089 ( .B1(n1574), .B2(n186), .A(n201), .ZN(n737) );
  NAND2_X1 U1090 ( .A1(\mem[9][14] ), .A2(n1611), .ZN(n201) );
  OAI21_X1 U1091 ( .B1(n1624), .B2(n186), .A(n202), .ZN(n738) );
  NAND2_X1 U1092 ( .A1(\mem[9][15] ), .A2(n1611), .ZN(n202) );
  OAI21_X1 U1093 ( .B1(n1639), .B2(n203), .A(n204), .ZN(n739) );
  NAND2_X1 U1094 ( .A1(\mem[10][0] ), .A2(n1610), .ZN(n204) );
  OAI21_X1 U1095 ( .B1(n1587), .B2(n203), .A(n205), .ZN(n740) );
  NAND2_X1 U1096 ( .A1(\mem[10][1] ), .A2(n1610), .ZN(n205) );
  OAI21_X1 U1097 ( .B1(n1637), .B2(n203), .A(n206), .ZN(n741) );
  NAND2_X1 U1098 ( .A1(\mem[10][2] ), .A2(n1610), .ZN(n206) );
  OAI21_X1 U1099 ( .B1(n1585), .B2(n203), .A(n207), .ZN(n742) );
  NAND2_X1 U1100 ( .A1(\mem[10][3] ), .A2(n1610), .ZN(n207) );
  OAI21_X1 U1101 ( .B1(n1631), .B2(n203), .A(n212), .ZN(n747) );
  NAND2_X1 U1102 ( .A1(\mem[10][8] ), .A2(n1610), .ZN(n212) );
  OAI21_X1 U1103 ( .B1(n1579), .B2(n203), .A(n213), .ZN(n748) );
  NAND2_X1 U1104 ( .A1(\mem[10][9] ), .A2(n1610), .ZN(n213) );
  OAI21_X1 U1105 ( .B1(n1578), .B2(n203), .A(n214), .ZN(n749) );
  NAND2_X1 U1106 ( .A1(\mem[10][10] ), .A2(n1610), .ZN(n214) );
  OAI21_X1 U1107 ( .B1(n1577), .B2(n203), .A(n215), .ZN(n750) );
  NAND2_X1 U1108 ( .A1(\mem[10][11] ), .A2(n1610), .ZN(n215) );
  OAI21_X1 U1109 ( .B1(n1576), .B2(n203), .A(n216), .ZN(n751) );
  NAND2_X1 U1110 ( .A1(\mem[10][12] ), .A2(n1610), .ZN(n216) );
  OAI21_X1 U1111 ( .B1(n1626), .B2(n203), .A(n217), .ZN(n752) );
  NAND2_X1 U1112 ( .A1(\mem[10][13] ), .A2(n1610), .ZN(n217) );
  OAI21_X1 U1113 ( .B1(n1574), .B2(n203), .A(n218), .ZN(n753) );
  NAND2_X1 U1114 ( .A1(\mem[10][14] ), .A2(n1610), .ZN(n218) );
  OAI21_X1 U1115 ( .B1(n1624), .B2(n203), .A(n219), .ZN(n754) );
  NAND2_X1 U1116 ( .A1(\mem[10][15] ), .A2(n1610), .ZN(n219) );
  OAI21_X1 U1117 ( .B1(n1639), .B2(n1609), .A(n221), .ZN(n755) );
  NAND2_X1 U1118 ( .A1(\mem[11][0] ), .A2(n220), .ZN(n221) );
  OAI21_X1 U1119 ( .B1(n1587), .B2(n1609), .A(n222), .ZN(n756) );
  NAND2_X1 U1120 ( .A1(\mem[11][1] ), .A2(n220), .ZN(n222) );
  OAI21_X1 U1121 ( .B1(n1637), .B2(n1609), .A(n223), .ZN(n757) );
  NAND2_X1 U1122 ( .A1(\mem[11][2] ), .A2(n220), .ZN(n223) );
  OAI21_X1 U1123 ( .B1(n1585), .B2(n1609), .A(n224), .ZN(n758) );
  NAND2_X1 U1124 ( .A1(\mem[11][3] ), .A2(n220), .ZN(n224) );
  OAI21_X1 U1125 ( .B1(n1631), .B2(n220), .A(n229), .ZN(n763) );
  NAND2_X1 U1126 ( .A1(\mem[11][8] ), .A2(n220), .ZN(n229) );
  OAI21_X1 U1127 ( .B1(n1579), .B2(n220), .A(n230), .ZN(n764) );
  NAND2_X1 U1128 ( .A1(\mem[11][9] ), .A2(n220), .ZN(n230) );
  OAI21_X1 U1129 ( .B1(n1578), .B2(n220), .A(n231), .ZN(n765) );
  NAND2_X1 U1130 ( .A1(\mem[11][10] ), .A2(n220), .ZN(n231) );
  OAI21_X1 U1131 ( .B1(n1577), .B2(n220), .A(n232), .ZN(n766) );
  NAND2_X1 U1132 ( .A1(\mem[11][11] ), .A2(n220), .ZN(n232) );
  OAI21_X1 U1133 ( .B1(n1576), .B2(n220), .A(n233), .ZN(n767) );
  NAND2_X1 U1134 ( .A1(\mem[11][12] ), .A2(n220), .ZN(n233) );
  OAI21_X1 U1135 ( .B1(n1626), .B2(n220), .A(n234), .ZN(n768) );
  NAND2_X1 U1136 ( .A1(\mem[11][13] ), .A2(n220), .ZN(n234) );
  OAI21_X1 U1137 ( .B1(n1574), .B2(n220), .A(n235), .ZN(n769) );
  NAND2_X1 U1138 ( .A1(\mem[11][14] ), .A2(n220), .ZN(n235) );
  OAI21_X1 U1139 ( .B1(n1624), .B2(n1609), .A(n236), .ZN(n770) );
  NAND2_X1 U1140 ( .A1(\mem[11][15] ), .A2(n220), .ZN(n236) );
  INV_X1 U1141 ( .A(data_in[0]), .ZN(n1639) );
  INV_X1 U1142 ( .A(data_in[1]), .ZN(n1638) );
  INV_X1 U1143 ( .A(data_in[2]), .ZN(n1637) );
  INV_X1 U1144 ( .A(data_in[3]), .ZN(n1636) );
  INV_X1 U1145 ( .A(data_in[4]), .ZN(n1635) );
  INV_X1 U1146 ( .A(data_in[5]), .ZN(n1634) );
  INV_X1 U1147 ( .A(data_in[6]), .ZN(n1633) );
  INV_X1 U1148 ( .A(data_in[7]), .ZN(n1632) );
  INV_X1 U1149 ( .A(data_in[8]), .ZN(n1631) );
  INV_X1 U1150 ( .A(data_in[9]), .ZN(n1630) );
  INV_X1 U1151 ( .A(data_in[10]), .ZN(n1629) );
  INV_X1 U1152 ( .A(data_in[11]), .ZN(n1628) );
  INV_X1 U1153 ( .A(data_in[12]), .ZN(n1627) );
  INV_X1 U1154 ( .A(data_in[13]), .ZN(n1626) );
  INV_X1 U1155 ( .A(data_in[14]), .ZN(n1625) );
  INV_X1 U1156 ( .A(data_in[15]), .ZN(n1624) );
  MUX2_X1 U1157 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n1561), .Z(n1) );
  MUX2_X1 U1158 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n1561), .Z(n2) );
  MUX2_X1 U1159 ( .A(n2), .B(n1), .S(n1555), .Z(n3) );
  MUX2_X1 U1160 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n1561), .Z(n4) );
  MUX2_X1 U1161 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n1561), .Z(n5) );
  MUX2_X1 U1162 ( .A(n5), .B(n4), .S(n1555), .Z(n6) );
  MUX2_X1 U1163 ( .A(n6), .B(n3), .S(n1552), .Z(n7) );
  MUX2_X1 U1164 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n1561), .Z(n8) );
  MUX2_X1 U1165 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n1561), .Z(n9) );
  MUX2_X1 U1166 ( .A(n9), .B(n8), .S(n1555), .Z(n10) );
  MUX2_X1 U1167 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n1561), .Z(n11) );
  MUX2_X1 U1168 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n1571), .Z(n12) );
  MUX2_X1 U1169 ( .A(n12), .B(n11), .S(n1555), .Z(n13) );
  MUX2_X1 U1170 ( .A(n13), .B(n10), .S(n1552), .Z(n14) );
  MUX2_X1 U1171 ( .A(n14), .B(n7), .S(n1550), .Z(n15) );
  MUX2_X1 U1172 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n1561), .Z(n16) );
  MUX2_X1 U1173 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n1561), .Z(n17) );
  MUX2_X1 U1174 ( .A(n17), .B(n16), .S(n1555), .Z(n18) );
  MUX2_X1 U1175 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n1561), .Z(n19) );
  MUX2_X1 U1176 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n1568), .Z(n20) );
  MUX2_X1 U1177 ( .A(n20), .B(n19), .S(n1555), .Z(n21) );
  MUX2_X1 U1178 ( .A(n21), .B(n18), .S(n1552), .Z(n1091) );
  MUX2_X1 U1179 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n1561), .Z(n1092) );
  MUX2_X1 U1180 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n1572), .Z(n1093) );
  MUX2_X1 U1181 ( .A(n1093), .B(n1092), .S(n1555), .Z(n1094) );
  MUX2_X1 U1182 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n1572), .Z(n1095) );
  MUX2_X1 U1183 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n1571), .Z(n1096) );
  MUX2_X1 U1184 ( .A(n1096), .B(n1095), .S(n1555), .Z(n1097) );
  MUX2_X1 U1185 ( .A(n1097), .B(n1094), .S(n1552), .Z(n1098) );
  MUX2_X1 U1186 ( .A(n1098), .B(n1091), .S(n1550), .Z(n1099) );
  MUX2_X1 U1187 ( .A(n1099), .B(n15), .S(N14), .Z(N30) );
  MUX2_X1 U1188 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n1562), .Z(n1100) );
  MUX2_X1 U1189 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n1562), .Z(n1101) );
  MUX2_X1 U1190 ( .A(n1101), .B(n1100), .S(N11), .Z(n1102) );
  MUX2_X1 U1191 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n1562), .Z(n1103) );
  MUX2_X1 U1192 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n1562), .Z(n1104) );
  MUX2_X1 U1193 ( .A(n1104), .B(n1103), .S(n1560), .Z(n1105) );
  MUX2_X1 U1194 ( .A(n1105), .B(n1102), .S(n1553), .Z(n1106) );
  MUX2_X1 U1195 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n1562), .Z(n1107) );
  MUX2_X1 U1196 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n1562), .Z(n1108) );
  MUX2_X1 U1197 ( .A(n1108), .B(n1107), .S(N11), .Z(n1109) );
  MUX2_X1 U1198 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n1562), .Z(n1110) );
  MUX2_X1 U1199 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n1562), .Z(n1111) );
  MUX2_X1 U1200 ( .A(n1111), .B(n1110), .S(n1560), .Z(n1112) );
  MUX2_X1 U1201 ( .A(n1112), .B(n1109), .S(n1553), .Z(n1113) );
  MUX2_X1 U1202 ( .A(n1113), .B(n1106), .S(n1551), .Z(n1114) );
  MUX2_X1 U1203 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n1562), .Z(n1115) );
  MUX2_X1 U1204 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n1562), .Z(n1116) );
  MUX2_X1 U1205 ( .A(n1116), .B(n1115), .S(n1560), .Z(n1117) );
  MUX2_X1 U1206 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n1562), .Z(n1118) );
  MUX2_X1 U1207 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n1562), .Z(n1119) );
  MUX2_X1 U1208 ( .A(n1119), .B(n1118), .S(n1560), .Z(n1120) );
  MUX2_X1 U1209 ( .A(n1120), .B(n1117), .S(n1553), .Z(n1121) );
  MUX2_X1 U1210 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n1563), .Z(n1122) );
  MUX2_X1 U1211 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n1563), .Z(n1123) );
  MUX2_X1 U1212 ( .A(n1123), .B(n1122), .S(n1560), .Z(n1124) );
  MUX2_X1 U1213 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n1563), .Z(n1125) );
  MUX2_X1 U1214 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n1563), .Z(n1126) );
  MUX2_X1 U1215 ( .A(n1126), .B(n1125), .S(N11), .Z(n1127) );
  MUX2_X1 U1216 ( .A(n1127), .B(n1124), .S(n1553), .Z(n1128) );
  MUX2_X1 U1217 ( .A(n1128), .B(n1121), .S(n1551), .Z(n1129) );
  MUX2_X1 U1218 ( .A(n1129), .B(n1114), .S(N14), .Z(N29) );
  MUX2_X1 U1219 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n1563), .Z(n1130) );
  MUX2_X1 U1220 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n1563), .Z(n1131) );
  MUX2_X1 U1221 ( .A(n1131), .B(n1130), .S(n1560), .Z(n1132) );
  MUX2_X1 U1222 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n1563), .Z(n1133) );
  MUX2_X1 U1223 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n1563), .Z(n1134) );
  MUX2_X1 U1224 ( .A(n1134), .B(n1133), .S(n1560), .Z(n1135) );
  MUX2_X1 U1225 ( .A(n1135), .B(n1132), .S(n1553), .Z(n1136) );
  MUX2_X1 U1226 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n1563), .Z(n1137) );
  MUX2_X1 U1227 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n1563), .Z(n1138) );
  MUX2_X1 U1228 ( .A(n1138), .B(n1137), .S(n1560), .Z(n1139) );
  MUX2_X1 U1229 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n1563), .Z(n1140) );
  MUX2_X1 U1230 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n1563), .Z(n1141) );
  MUX2_X1 U1231 ( .A(n1141), .B(n1140), .S(n1560), .Z(n1142) );
  MUX2_X1 U1232 ( .A(n1142), .B(n1139), .S(n1553), .Z(n1143) );
  MUX2_X1 U1233 ( .A(n1143), .B(n1136), .S(n1550), .Z(n1144) );
  MUX2_X1 U1234 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n1567), .Z(n1145) );
  MUX2_X1 U1235 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n1565), .Z(n1146) );
  MUX2_X1 U1236 ( .A(n1146), .B(n1145), .S(n1555), .Z(n1147) );
  MUX2_X1 U1237 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n1570), .Z(n1148) );
  MUX2_X1 U1238 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n1567), .Z(n1149) );
  MUX2_X1 U1239 ( .A(n1149), .B(n1148), .S(n1560), .Z(n1150) );
  MUX2_X1 U1240 ( .A(n1150), .B(n1147), .S(n1553), .Z(n1151) );
  MUX2_X1 U1241 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n1572), .Z(n1152) );
  MUX2_X1 U1242 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n1571), .Z(n1153) );
  MUX2_X1 U1243 ( .A(n1153), .B(n1152), .S(n1560), .Z(n1154) );
  MUX2_X1 U1244 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n1572), .Z(n1155) );
  MUX2_X1 U1245 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n1571), .Z(n1156) );
  MUX2_X1 U1246 ( .A(n1156), .B(n1155), .S(n1560), .Z(n1157) );
  MUX2_X1 U1247 ( .A(n1157), .B(n1154), .S(n1553), .Z(n1158) );
  MUX2_X1 U1248 ( .A(n1158), .B(n1151), .S(n1550), .Z(n1159) );
  MUX2_X1 U1249 ( .A(n1159), .B(n1144), .S(N14), .Z(N28) );
  MUX2_X1 U1250 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n1571), .Z(n1160) );
  MUX2_X1 U1251 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n1563), .Z(n1161) );
  MUX2_X1 U1252 ( .A(n1161), .B(n1160), .S(n1555), .Z(n1162) );
  MUX2_X1 U1253 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n1563), .Z(n1163) );
  MUX2_X1 U1254 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n1571), .Z(n1164) );
  MUX2_X1 U1255 ( .A(n1164), .B(n1163), .S(n1560), .Z(n1165) );
  MUX2_X1 U1256 ( .A(n1165), .B(n1162), .S(n1553), .Z(n1166) );
  MUX2_X1 U1257 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n1568), .Z(n1167) );
  MUX2_X1 U1258 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n1571), .Z(n1168) );
  MUX2_X1 U1259 ( .A(n1168), .B(n1167), .S(n1555), .Z(n1169) );
  MUX2_X1 U1260 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n1572), .Z(n1170) );
  MUX2_X1 U1261 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n1571), .Z(n1171) );
  MUX2_X1 U1262 ( .A(n1171), .B(n1170), .S(n1560), .Z(n1172) );
  MUX2_X1 U1263 ( .A(n1172), .B(n1169), .S(n1553), .Z(n1173) );
  MUX2_X1 U1264 ( .A(n1173), .B(n1166), .S(n1551), .Z(n1174) );
  MUX2_X1 U1265 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n1561), .Z(n1175) );
  MUX2_X1 U1266 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n1571), .Z(n1176) );
  MUX2_X1 U1267 ( .A(n1176), .B(n1175), .S(n1560), .Z(n1177) );
  MUX2_X1 U1268 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n1572), .Z(n1178) );
  MUX2_X1 U1269 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n1571), .Z(n1179) );
  MUX2_X1 U1270 ( .A(n1179), .B(n1178), .S(n1560), .Z(n1180) );
  MUX2_X1 U1271 ( .A(n1180), .B(n1177), .S(n1553), .Z(n1181) );
  MUX2_X1 U1272 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n1571), .Z(n1182) );
  MUX2_X1 U1273 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n1572), .Z(n1183) );
  MUX2_X1 U1274 ( .A(n1183), .B(n1182), .S(n1560), .Z(n1184) );
  MUX2_X1 U1275 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n1565), .Z(n1185) );
  MUX2_X1 U1276 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n1572), .Z(n1186) );
  MUX2_X1 U1277 ( .A(n1186), .B(n1185), .S(n1560), .Z(n1187) );
  MUX2_X1 U1278 ( .A(n1187), .B(n1184), .S(n1553), .Z(n1188) );
  MUX2_X1 U1279 ( .A(n1188), .B(n1181), .S(n1551), .Z(n1189) );
  MUX2_X1 U1280 ( .A(n1189), .B(n1174), .S(N14), .Z(N27) );
  MUX2_X1 U1281 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n1562), .Z(n1190) );
  MUX2_X1 U1282 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n1568), .Z(n1191) );
  MUX2_X1 U1283 ( .A(n1191), .B(n1190), .S(n1556), .Z(n1192) );
  MUX2_X1 U1284 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n1565), .Z(n1193) );
  MUX2_X1 U1285 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n1194) );
  MUX2_X1 U1286 ( .A(n1194), .B(n1193), .S(n1556), .Z(n1195) );
  MUX2_X1 U1287 ( .A(n1195), .B(n1192), .S(n1552), .Z(n1196) );
  MUX2_X1 U1288 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n1563), .Z(n1197) );
  MUX2_X1 U1289 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n1571), .Z(n1198) );
  MUX2_X1 U1290 ( .A(n1198), .B(n1197), .S(n1556), .Z(n1199) );
  MUX2_X1 U1291 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n1571), .Z(n1200) );
  MUX2_X1 U1292 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(N10), .Z(n1201) );
  MUX2_X1 U1293 ( .A(n1201), .B(n1200), .S(n1556), .Z(n1202) );
  MUX2_X1 U1294 ( .A(n1202), .B(n1199), .S(n1552), .Z(n1203) );
  MUX2_X1 U1295 ( .A(n1203), .B(n1196), .S(n1550), .Z(n1204) );
  MUX2_X1 U1296 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n1567), .Z(n1205) );
  MUX2_X1 U1297 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(N10), .Z(n1206) );
  MUX2_X1 U1298 ( .A(n1206), .B(n1205), .S(n1556), .Z(n1207) );
  MUX2_X1 U1299 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n1569), .Z(n1208) );
  MUX2_X1 U1300 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n1209) );
  MUX2_X1 U1301 ( .A(n1209), .B(n1208), .S(n1556), .Z(n1210) );
  MUX2_X1 U1302 ( .A(n1210), .B(n1207), .S(n1552), .Z(n1211) );
  MUX2_X1 U1303 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n1561), .Z(n1212) );
  MUX2_X1 U1304 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n1561), .Z(n1213) );
  MUX2_X1 U1305 ( .A(n1213), .B(n1212), .S(n1556), .Z(n1214) );
  MUX2_X1 U1306 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n1561), .Z(n1215) );
  MUX2_X1 U1307 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n1562), .Z(n1216) );
  MUX2_X1 U1308 ( .A(n1216), .B(n1215), .S(n1556), .Z(n1217) );
  MUX2_X1 U1309 ( .A(n1217), .B(n1214), .S(n1554), .Z(n1218) );
  MUX2_X1 U1310 ( .A(n1218), .B(n1211), .S(n1550), .Z(n1219) );
  MUX2_X1 U1311 ( .A(n1219), .B(n1204), .S(N14), .Z(N26) );
  MUX2_X1 U1312 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n1561), .Z(n1220) );
  MUX2_X1 U1313 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n1562), .Z(n1221) );
  MUX2_X1 U1314 ( .A(n1221), .B(n1220), .S(n1556), .Z(n1222) );
  MUX2_X1 U1315 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n1561), .Z(n1223) );
  MUX2_X1 U1316 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n1563), .Z(n1224) );
  MUX2_X1 U1317 ( .A(n1224), .B(n1223), .S(n1556), .Z(n1225) );
  MUX2_X1 U1318 ( .A(n1225), .B(n1222), .S(n1552), .Z(n1226) );
  MUX2_X1 U1319 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n1562), .Z(n1227) );
  MUX2_X1 U1320 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n1562), .Z(n1228) );
  MUX2_X1 U1321 ( .A(n1228), .B(n1227), .S(n1556), .Z(n1229) );
  MUX2_X1 U1322 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n1563), .Z(n1230) );
  MUX2_X1 U1323 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n1563), .Z(n1231) );
  MUX2_X1 U1324 ( .A(n1231), .B(n1230), .S(n1556), .Z(n1232) );
  MUX2_X1 U1325 ( .A(n1232), .B(n1229), .S(n1552), .Z(n1233) );
  MUX2_X1 U1326 ( .A(n1233), .B(n1226), .S(n1550), .Z(n1234) );
  MUX2_X1 U1327 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n1562), .Z(n1235) );
  MUX2_X1 U1328 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n1566), .Z(n1236) );
  MUX2_X1 U1329 ( .A(n1236), .B(n1235), .S(n1557), .Z(n1237) );
  MUX2_X1 U1330 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n1572), .Z(n1238) );
  MUX2_X1 U1331 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n1567), .Z(n1239) );
  MUX2_X1 U1332 ( .A(n1239), .B(n1238), .S(n1557), .Z(n1240) );
  MUX2_X1 U1333 ( .A(n1240), .B(n1237), .S(n1552), .Z(n1241) );
  MUX2_X1 U1334 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n1572), .Z(n1242) );
  MUX2_X1 U1335 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n1568), .Z(n1243) );
  MUX2_X1 U1336 ( .A(n1243), .B(n1242), .S(n1557), .Z(n1244) );
  MUX2_X1 U1337 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n1562), .Z(n1245) );
  MUX2_X1 U1338 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n1571), .Z(n1246) );
  MUX2_X1 U1339 ( .A(n1246), .B(n1245), .S(n1557), .Z(n1247) );
  MUX2_X1 U1340 ( .A(n1247), .B(n1244), .S(N12), .Z(n1248) );
  MUX2_X1 U1341 ( .A(n1248), .B(n1241), .S(n1550), .Z(n1249) );
  MUX2_X1 U1342 ( .A(n1249), .B(n1234), .S(N14), .Z(N25) );
  MUX2_X1 U1343 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n1563), .Z(n1250) );
  MUX2_X1 U1344 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n1572), .Z(n1251) );
  MUX2_X1 U1345 ( .A(n1251), .B(n1250), .S(n1557), .Z(n1252) );
  MUX2_X1 U1346 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n1572), .Z(n1253) );
  MUX2_X1 U1347 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n1571), .Z(n1254) );
  MUX2_X1 U1348 ( .A(n1254), .B(n1253), .S(n1557), .Z(n1255) );
  MUX2_X1 U1349 ( .A(n1255), .B(n1252), .S(n1552), .Z(n1256) );
  MUX2_X1 U1350 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n1562), .Z(n1257) );
  MUX2_X1 U1351 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n1571), .Z(n1258) );
  MUX2_X1 U1352 ( .A(n1258), .B(n1257), .S(n1557), .Z(n1259) );
  MUX2_X1 U1353 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n1572), .Z(n1260) );
  MUX2_X1 U1354 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n1572), .Z(n1261) );
  MUX2_X1 U1355 ( .A(n1261), .B(n1260), .S(n1557), .Z(n1262) );
  MUX2_X1 U1356 ( .A(n1262), .B(n1259), .S(n1553), .Z(n1263) );
  MUX2_X1 U1357 ( .A(n1263), .B(n1256), .S(n1550), .Z(n1264) );
  MUX2_X1 U1358 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n1565), .Z(n1265) );
  MUX2_X1 U1359 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n1572), .Z(n1266) );
  MUX2_X1 U1360 ( .A(n1266), .B(n1265), .S(n1557), .Z(n1267) );
  MUX2_X1 U1361 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n1569), .Z(n1268) );
  MUX2_X1 U1362 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n1571), .Z(n1269) );
  MUX2_X1 U1363 ( .A(n1269), .B(n1268), .S(n1557), .Z(n1270) );
  MUX2_X1 U1364 ( .A(n1270), .B(n1267), .S(n1552), .Z(n1271) );
  MUX2_X1 U1365 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n1571), .Z(n1272) );
  MUX2_X1 U1366 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n1572), .Z(n1273) );
  MUX2_X1 U1367 ( .A(n1273), .B(n1272), .S(n1557), .Z(n1274) );
  MUX2_X1 U1368 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n1571), .Z(n1275) );
  MUX2_X1 U1369 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n1571), .Z(n1276) );
  MUX2_X1 U1370 ( .A(n1276), .B(n1275), .S(n1557), .Z(n1277) );
  MUX2_X1 U1371 ( .A(n1277), .B(n1274), .S(n1552), .Z(n1278) );
  MUX2_X1 U1372 ( .A(n1278), .B(n1271), .S(n1550), .Z(n1279) );
  MUX2_X1 U1373 ( .A(n1279), .B(n1264), .S(N14), .Z(N24) );
  MUX2_X1 U1374 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n1566), .Z(n1280) );
  MUX2_X1 U1375 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n1572), .Z(n1281) );
  MUX2_X1 U1376 ( .A(n1281), .B(n1280), .S(n1560), .Z(n1282) );
  MUX2_X1 U1377 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n1572), .Z(n1283) );
  MUX2_X1 U1378 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n1570), .Z(n1284) );
  MUX2_X1 U1379 ( .A(n1284), .B(n1283), .S(n1556), .Z(n1285) );
  MUX2_X1 U1380 ( .A(n1285), .B(n1282), .S(n1552), .Z(n1286) );
  MUX2_X1 U1381 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n1566), .Z(n1287) );
  MUX2_X1 U1382 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n1564), .Z(n1288) );
  MUX2_X1 U1383 ( .A(n1288), .B(n1287), .S(n1556), .Z(n1289) );
  MUX2_X1 U1384 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n1563), .Z(n1290) );
  MUX2_X1 U1385 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n1569), .Z(n1291) );
  MUX2_X1 U1386 ( .A(n1291), .B(n1290), .S(n1559), .Z(n1292) );
  MUX2_X1 U1387 ( .A(n1292), .B(n1289), .S(n1554), .Z(n1293) );
  MUX2_X1 U1388 ( .A(n1293), .B(n1286), .S(n1550), .Z(n1294) );
  MUX2_X1 U1389 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n1564), .Z(n1295) );
  MUX2_X1 U1390 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n1569), .Z(n1296) );
  MUX2_X1 U1391 ( .A(n1296), .B(n1295), .S(n1556), .Z(n1297) );
  MUX2_X1 U1392 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n1570), .Z(n1298) );
  MUX2_X1 U1393 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n1572), .Z(n1299) );
  MUX2_X1 U1394 ( .A(n1299), .B(n1298), .S(n1558), .Z(n1300) );
  MUX2_X1 U1395 ( .A(n1300), .B(n1297), .S(n1553), .Z(n1301) );
  MUX2_X1 U1396 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n1561), .Z(n1302) );
  MUX2_X1 U1397 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n1563), .Z(n1303) );
  MUX2_X1 U1398 ( .A(n1303), .B(n1302), .S(n1559), .Z(n1304) );
  MUX2_X1 U1399 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n1562), .Z(n1305) );
  MUX2_X1 U1400 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n1562), .Z(n1306) );
  MUX2_X1 U1401 ( .A(n1306), .B(n1305), .S(n1559), .Z(n1307) );
  MUX2_X1 U1402 ( .A(n1307), .B(n1304), .S(n1553), .Z(n1308) );
  MUX2_X1 U1403 ( .A(n1308), .B(n1301), .S(n1550), .Z(n1309) );
  MUX2_X1 U1404 ( .A(n1309), .B(n1294), .S(N14), .Z(N23) );
  MUX2_X1 U1405 ( .A(\mem[30][8] ), .B(\mem[31][8] ), .S(n1561), .Z(n1310) );
  MUX2_X1 U1406 ( .A(\mem[28][8] ), .B(\mem[29][8] ), .S(n1561), .Z(n1311) );
  MUX2_X1 U1407 ( .A(n1311), .B(n1310), .S(n1558), .Z(n1312) );
  MUX2_X1 U1408 ( .A(\mem[26][8] ), .B(\mem[27][8] ), .S(n1561), .Z(n1313) );
  MUX2_X1 U1409 ( .A(\mem[24][8] ), .B(\mem[25][8] ), .S(n1563), .Z(n1314) );
  MUX2_X1 U1410 ( .A(n1314), .B(n1313), .S(n1558), .Z(n1315) );
  MUX2_X1 U1411 ( .A(n1315), .B(n1312), .S(n1554), .Z(n1316) );
  MUX2_X1 U1412 ( .A(\mem[22][8] ), .B(\mem[23][8] ), .S(n1561), .Z(n1317) );
  MUX2_X1 U1413 ( .A(\mem[20][8] ), .B(\mem[21][8] ), .S(n1561), .Z(n1318) );
  MUX2_X1 U1414 ( .A(n1318), .B(n1317), .S(n1559), .Z(n1319) );
  MUX2_X1 U1415 ( .A(\mem[18][8] ), .B(\mem[19][8] ), .S(n1563), .Z(n1320) );
  MUX2_X1 U1416 ( .A(\mem[16][8] ), .B(\mem[17][8] ), .S(n1562), .Z(n1321) );
  MUX2_X1 U1417 ( .A(n1321), .B(n1320), .S(n1556), .Z(n1322) );
  MUX2_X1 U1418 ( .A(n1322), .B(n1319), .S(n1552), .Z(n1323) );
  MUX2_X1 U1419 ( .A(n1323), .B(n1316), .S(n1550), .Z(n1324) );
  MUX2_X1 U1420 ( .A(\mem[14][8] ), .B(\mem[15][8] ), .S(n1564), .Z(n1325) );
  MUX2_X1 U1421 ( .A(\mem[12][8] ), .B(\mem[13][8] ), .S(n1564), .Z(n1326) );
  MUX2_X1 U1422 ( .A(n1326), .B(n1325), .S(n1555), .Z(n1327) );
  MUX2_X1 U1423 ( .A(\mem[10][8] ), .B(\mem[11][8] ), .S(n1564), .Z(n1328) );
  MUX2_X1 U1424 ( .A(\mem[8][8] ), .B(\mem[9][8] ), .S(n1564), .Z(n1329) );
  MUX2_X1 U1425 ( .A(n1329), .B(n1328), .S(n1557), .Z(n1330) );
  MUX2_X1 U1426 ( .A(n1330), .B(n1327), .S(n1552), .Z(n1331) );
  MUX2_X1 U1427 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n1564), .Z(n1332) );
  MUX2_X1 U1428 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n1564), .Z(n1333) );
  MUX2_X1 U1429 ( .A(n1333), .B(n1332), .S(n1555), .Z(n1334) );
  MUX2_X1 U1430 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n1564), .Z(n1335) );
  MUX2_X1 U1431 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n1564), .Z(n1336) );
  MUX2_X1 U1432 ( .A(n1336), .B(n1335), .S(n1557), .Z(n1337) );
  MUX2_X1 U1433 ( .A(n1337), .B(n1334), .S(n1554), .Z(n1338) );
  MUX2_X1 U1434 ( .A(n1338), .B(n1331), .S(n1550), .Z(n1339) );
  MUX2_X1 U1435 ( .A(n1339), .B(n1324), .S(N14), .Z(N22) );
  MUX2_X1 U1436 ( .A(\mem[30][9] ), .B(\mem[31][9] ), .S(n1564), .Z(n1340) );
  MUX2_X1 U1437 ( .A(\mem[28][9] ), .B(\mem[29][9] ), .S(n1564), .Z(n1341) );
  MUX2_X1 U1438 ( .A(n1341), .B(n1340), .S(n1555), .Z(n1342) );
  MUX2_X1 U1439 ( .A(\mem[26][9] ), .B(\mem[27][9] ), .S(n1564), .Z(n1343) );
  MUX2_X1 U1440 ( .A(\mem[24][9] ), .B(\mem[25][9] ), .S(n1564), .Z(n1344) );
  MUX2_X1 U1441 ( .A(n1344), .B(n1343), .S(n1557), .Z(n1345) );
  MUX2_X1 U1442 ( .A(n1345), .B(n1342), .S(n1554), .Z(n1346) );
  MUX2_X1 U1443 ( .A(\mem[22][9] ), .B(\mem[23][9] ), .S(n1564), .Z(n1347) );
  MUX2_X1 U1444 ( .A(\mem[20][9] ), .B(\mem[21][9] ), .S(n1564), .Z(n1348) );
  MUX2_X1 U1445 ( .A(n1348), .B(n1347), .S(n1555), .Z(n1349) );
  MUX2_X1 U1446 ( .A(\mem[18][9] ), .B(\mem[19][9] ), .S(n1567), .Z(n1350) );
  MUX2_X1 U1447 ( .A(\mem[16][9] ), .B(\mem[17][9] ), .S(n1566), .Z(n1351) );
  MUX2_X1 U1448 ( .A(n1351), .B(n1350), .S(n1555), .Z(n1352) );
  MUX2_X1 U1449 ( .A(n1352), .B(n1349), .S(n1552), .Z(n1353) );
  MUX2_X1 U1450 ( .A(n1353), .B(n1346), .S(n1550), .Z(n1354) );
  MUX2_X1 U1451 ( .A(\mem[14][9] ), .B(\mem[15][9] ), .S(n1566), .Z(n1355) );
  MUX2_X1 U1452 ( .A(\mem[12][9] ), .B(\mem[13][9] ), .S(n1570), .Z(n1356) );
  MUX2_X1 U1453 ( .A(n1356), .B(n1355), .S(n1555), .Z(n1357) );
  MUX2_X1 U1454 ( .A(\mem[10][9] ), .B(\mem[11][9] ), .S(n1565), .Z(n1358) );
  MUX2_X1 U1455 ( .A(\mem[8][9] ), .B(\mem[9][9] ), .S(n1567), .Z(n1359) );
  MUX2_X1 U1456 ( .A(n1359), .B(n1358), .S(n1555), .Z(n1360) );
  MUX2_X1 U1457 ( .A(n1360), .B(n1357), .S(n1553), .Z(n1361) );
  MUX2_X1 U1458 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n1568), .Z(n1362) );
  MUX2_X1 U1459 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n1568), .Z(n1363) );
  MUX2_X1 U1460 ( .A(n1363), .B(n1362), .S(n1557), .Z(n1364) );
  MUX2_X1 U1461 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n1570), .Z(n1365) );
  MUX2_X1 U1462 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n1569), .Z(n1366) );
  MUX2_X1 U1463 ( .A(n1366), .B(n1365), .S(n1560), .Z(n1367) );
  MUX2_X1 U1464 ( .A(n1367), .B(n1364), .S(n1553), .Z(n1368) );
  MUX2_X1 U1465 ( .A(n1368), .B(n1361), .S(n1550), .Z(n1369) );
  MUX2_X1 U1466 ( .A(n1369), .B(n1354), .S(N14), .Z(N21) );
  MUX2_X1 U1467 ( .A(\mem[30][10] ), .B(\mem[31][10] ), .S(n1568), .Z(n1370)
         );
  MUX2_X1 U1468 ( .A(\mem[28][10] ), .B(\mem[29][10] ), .S(n1566), .Z(n1371)
         );
  MUX2_X1 U1469 ( .A(n1371), .B(n1370), .S(n1557), .Z(n1372) );
  MUX2_X1 U1470 ( .A(\mem[26][10] ), .B(\mem[27][10] ), .S(n1565), .Z(n1373)
         );
  MUX2_X1 U1471 ( .A(\mem[24][10] ), .B(\mem[25][10] ), .S(n1567), .Z(n1374)
         );
  MUX2_X1 U1472 ( .A(n1374), .B(n1373), .S(n1557), .Z(n1375) );
  MUX2_X1 U1473 ( .A(n1375), .B(n1372), .S(n1554), .Z(n1376) );
  MUX2_X1 U1474 ( .A(\mem[22][10] ), .B(\mem[23][10] ), .S(n1567), .Z(n1377)
         );
  MUX2_X1 U1475 ( .A(\mem[20][10] ), .B(\mem[21][10] ), .S(n1565), .Z(n1378)
         );
  MUX2_X1 U1476 ( .A(n1378), .B(n1377), .S(n1555), .Z(n1379) );
  MUX2_X1 U1477 ( .A(\mem[18][10] ), .B(\mem[19][10] ), .S(n1569), .Z(n1380)
         );
  MUX2_X1 U1478 ( .A(\mem[16][10] ), .B(\mem[17][10] ), .S(n1564), .Z(n1381)
         );
  MUX2_X1 U1479 ( .A(n1381), .B(n1380), .S(n1555), .Z(n1382) );
  MUX2_X1 U1480 ( .A(n1382), .B(n1379), .S(n1552), .Z(n1383) );
  MUX2_X1 U1481 ( .A(n1383), .B(n1376), .S(n1551), .Z(n1384) );
  MUX2_X1 U1482 ( .A(\mem[14][10] ), .B(\mem[15][10] ), .S(n1570), .Z(n1385)
         );
  MUX2_X1 U1483 ( .A(\mem[12][10] ), .B(\mem[13][10] ), .S(n1568), .Z(n1386)
         );
  MUX2_X1 U1484 ( .A(n1386), .B(n1385), .S(n1555), .Z(n1387) );
  MUX2_X1 U1485 ( .A(\mem[10][10] ), .B(\mem[11][10] ), .S(n1570), .Z(n1388)
         );
  MUX2_X1 U1486 ( .A(\mem[8][10] ), .B(\mem[9][10] ), .S(n1565), .Z(n1389) );
  MUX2_X1 U1487 ( .A(n1389), .B(n1388), .S(n1555), .Z(n1390) );
  MUX2_X1 U1488 ( .A(n1390), .B(n1387), .S(n1552), .Z(n1391) );
  MUX2_X1 U1489 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n1569), .Z(n1392) );
  MUX2_X1 U1490 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n1569), .Z(n1393) );
  MUX2_X1 U1491 ( .A(n1393), .B(n1392), .S(n1557), .Z(n1394) );
  MUX2_X1 U1492 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n1569), .Z(n1395) );
  MUX2_X1 U1493 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n1566), .Z(n1396) );
  MUX2_X1 U1494 ( .A(n1396), .B(n1395), .S(n1557), .Z(n1397) );
  MUX2_X1 U1495 ( .A(n1397), .B(n1394), .S(n1553), .Z(n1398) );
  MUX2_X1 U1496 ( .A(n1398), .B(n1391), .S(n1551), .Z(n1399) );
  MUX2_X1 U1497 ( .A(n1399), .B(n1384), .S(N14), .Z(N20) );
  MUX2_X1 U1498 ( .A(\mem[30][11] ), .B(\mem[31][11] ), .S(n1566), .Z(n1400)
         );
  MUX2_X1 U1499 ( .A(\mem[28][11] ), .B(\mem[29][11] ), .S(n1567), .Z(n1401)
         );
  MUX2_X1 U1500 ( .A(n1401), .B(n1400), .S(n1557), .Z(n1402) );
  MUX2_X1 U1501 ( .A(\mem[26][11] ), .B(\mem[27][11] ), .S(n1568), .Z(n1403)
         );
  MUX2_X1 U1502 ( .A(\mem[24][11] ), .B(\mem[25][11] ), .S(n1570), .Z(n1404)
         );
  MUX2_X1 U1503 ( .A(n1404), .B(n1403), .S(n1555), .Z(n1405) );
  MUX2_X1 U1504 ( .A(n1405), .B(n1402), .S(n1552), .Z(n1406) );
  MUX2_X1 U1505 ( .A(\mem[22][11] ), .B(\mem[23][11] ), .S(n1565), .Z(n1407)
         );
  MUX2_X1 U1506 ( .A(\mem[20][11] ), .B(\mem[21][11] ), .S(n1564), .Z(n1408)
         );
  MUX2_X1 U1507 ( .A(n1408), .B(n1407), .S(n1557), .Z(n1409) );
  MUX2_X1 U1508 ( .A(\mem[18][11] ), .B(\mem[19][11] ), .S(n1566), .Z(n1410)
         );
  MUX2_X1 U1509 ( .A(\mem[16][11] ), .B(\mem[17][11] ), .S(n1570), .Z(n1411)
         );
  MUX2_X1 U1510 ( .A(n1411), .B(n1410), .S(n1557), .Z(n1412) );
  MUX2_X1 U1511 ( .A(n1412), .B(n1409), .S(n1553), .Z(n1413) );
  MUX2_X1 U1512 ( .A(n1413), .B(n1406), .S(n1551), .Z(n1414) );
  MUX2_X1 U1513 ( .A(\mem[14][11] ), .B(\mem[15][11] ), .S(n1565), .Z(n1415)
         );
  MUX2_X1 U1514 ( .A(\mem[12][11] ), .B(\mem[13][11] ), .S(n1565), .Z(n1416)
         );
  MUX2_X1 U1515 ( .A(n1416), .B(n1415), .S(n1558), .Z(n1417) );
  MUX2_X1 U1516 ( .A(\mem[10][11] ), .B(\mem[11][11] ), .S(n1565), .Z(n1418)
         );
  MUX2_X1 U1517 ( .A(\mem[8][11] ), .B(\mem[9][11] ), .S(n1565), .Z(n1419) );
  MUX2_X1 U1518 ( .A(n1419), .B(n1418), .S(n1558), .Z(n1420) );
  MUX2_X1 U1519 ( .A(n1420), .B(n1417), .S(n1553), .Z(n1421) );
  MUX2_X1 U1520 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n1565), .Z(n1422) );
  MUX2_X1 U1521 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n1565), .Z(n1423) );
  MUX2_X1 U1522 ( .A(n1423), .B(n1422), .S(n1558), .Z(n1424) );
  MUX2_X1 U1523 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n1565), .Z(n1425) );
  MUX2_X1 U1524 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n1565), .Z(n1426) );
  MUX2_X1 U1525 ( .A(n1426), .B(n1425), .S(n1558), .Z(n1427) );
  MUX2_X1 U1526 ( .A(n1427), .B(n1424), .S(n1554), .Z(n1428) );
  MUX2_X1 U1527 ( .A(n1428), .B(n1421), .S(n1551), .Z(n1429) );
  MUX2_X1 U1528 ( .A(n1429), .B(n1414), .S(N14), .Z(N19) );
  MUX2_X1 U1529 ( .A(\mem[30][12] ), .B(\mem[31][12] ), .S(n1565), .Z(n1430)
         );
  MUX2_X1 U1530 ( .A(\mem[28][12] ), .B(\mem[29][12] ), .S(n1565), .Z(n1431)
         );
  MUX2_X1 U1531 ( .A(n1431), .B(n1430), .S(n1558), .Z(n1432) );
  MUX2_X1 U1532 ( .A(\mem[26][12] ), .B(\mem[27][12] ), .S(n1565), .Z(n1433)
         );
  MUX2_X1 U1533 ( .A(\mem[24][12] ), .B(\mem[25][12] ), .S(n1565), .Z(n1434)
         );
  MUX2_X1 U1534 ( .A(n1434), .B(n1433), .S(n1558), .Z(n1435) );
  MUX2_X1 U1535 ( .A(n1435), .B(n1432), .S(n1553), .Z(n1436) );
  MUX2_X1 U1536 ( .A(\mem[22][12] ), .B(\mem[23][12] ), .S(n1566), .Z(n1437)
         );
  MUX2_X1 U1537 ( .A(\mem[20][12] ), .B(\mem[21][12] ), .S(n1566), .Z(n1438)
         );
  MUX2_X1 U1538 ( .A(n1438), .B(n1437), .S(n1558), .Z(n1439) );
  MUX2_X1 U1539 ( .A(\mem[18][12] ), .B(\mem[19][12] ), .S(n1566), .Z(n1440)
         );
  MUX2_X1 U1540 ( .A(\mem[16][12] ), .B(\mem[17][12] ), .S(n1566), .Z(n1441)
         );
  MUX2_X1 U1541 ( .A(n1441), .B(n1440), .S(n1558), .Z(n1442) );
  MUX2_X1 U1542 ( .A(n1442), .B(n1439), .S(n1554), .Z(n1443) );
  MUX2_X1 U1543 ( .A(n1443), .B(n1436), .S(n1551), .Z(n1444) );
  MUX2_X1 U1544 ( .A(\mem[14][12] ), .B(\mem[15][12] ), .S(n1566), .Z(n1445)
         );
  MUX2_X1 U1545 ( .A(\mem[12][12] ), .B(\mem[13][12] ), .S(n1566), .Z(n1446)
         );
  MUX2_X1 U1546 ( .A(n1446), .B(n1445), .S(n1558), .Z(n1447) );
  MUX2_X1 U1547 ( .A(\mem[10][12] ), .B(\mem[11][12] ), .S(n1566), .Z(n1448)
         );
  MUX2_X1 U1548 ( .A(\mem[8][12] ), .B(\mem[9][12] ), .S(n1566), .Z(n1449) );
  MUX2_X1 U1549 ( .A(n1449), .B(n1448), .S(n1558), .Z(n1450) );
  MUX2_X1 U1550 ( .A(n1450), .B(n1447), .S(n1554), .Z(n1451) );
  MUX2_X1 U1551 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n1566), .Z(n1452) );
  MUX2_X1 U1552 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n1566), .Z(n1453) );
  MUX2_X1 U1553 ( .A(n1453), .B(n1452), .S(n1558), .Z(n1454) );
  MUX2_X1 U1554 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n1566), .Z(n1455) );
  MUX2_X1 U1555 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n1566), .Z(n1456) );
  MUX2_X1 U1556 ( .A(n1456), .B(n1455), .S(n1558), .Z(n1457) );
  MUX2_X1 U1557 ( .A(n1457), .B(n1454), .S(n1552), .Z(n1458) );
  MUX2_X1 U1558 ( .A(n1458), .B(n1451), .S(n1551), .Z(n1459) );
  MUX2_X1 U1559 ( .A(n1459), .B(n1444), .S(N14), .Z(N18) );
  MUX2_X1 U1560 ( .A(\mem[30][13] ), .B(\mem[31][13] ), .S(n1567), .Z(n1460)
         );
  MUX2_X1 U1561 ( .A(\mem[28][13] ), .B(\mem[29][13] ), .S(n1567), .Z(n1461)
         );
  MUX2_X1 U1562 ( .A(n1461), .B(n1460), .S(n1559), .Z(n1462) );
  MUX2_X1 U1563 ( .A(\mem[26][13] ), .B(\mem[27][13] ), .S(n1567), .Z(n1463)
         );
  MUX2_X1 U1564 ( .A(\mem[24][13] ), .B(\mem[25][13] ), .S(n1567), .Z(n1464)
         );
  MUX2_X1 U1565 ( .A(n1464), .B(n1463), .S(n1559), .Z(n1465) );
  MUX2_X1 U1566 ( .A(n1465), .B(n1462), .S(n1554), .Z(n1466) );
  MUX2_X1 U1567 ( .A(\mem[22][13] ), .B(\mem[23][13] ), .S(n1567), .Z(n1467)
         );
  MUX2_X1 U1568 ( .A(\mem[20][13] ), .B(\mem[21][13] ), .S(n1567), .Z(n1468)
         );
  MUX2_X1 U1569 ( .A(n1468), .B(n1467), .S(n1559), .Z(n1469) );
  MUX2_X1 U1570 ( .A(\mem[18][13] ), .B(\mem[19][13] ), .S(n1567), .Z(n1470)
         );
  MUX2_X1 U1571 ( .A(\mem[16][13] ), .B(\mem[17][13] ), .S(n1567), .Z(n1471)
         );
  MUX2_X1 U1572 ( .A(n1471), .B(n1470), .S(n1559), .Z(n1472) );
  MUX2_X1 U1573 ( .A(n1472), .B(n1469), .S(n1554), .Z(n1473) );
  MUX2_X1 U1574 ( .A(n1473), .B(n1466), .S(n1551), .Z(n1474) );
  MUX2_X1 U1575 ( .A(\mem[14][13] ), .B(\mem[15][13] ), .S(n1567), .Z(n1475)
         );
  MUX2_X1 U1576 ( .A(\mem[12][13] ), .B(\mem[13][13] ), .S(n1567), .Z(n1476)
         );
  MUX2_X1 U1577 ( .A(n1476), .B(n1475), .S(n1559), .Z(n1477) );
  MUX2_X1 U1578 ( .A(\mem[10][13] ), .B(\mem[11][13] ), .S(n1567), .Z(n1478)
         );
  MUX2_X1 U1579 ( .A(\mem[8][13] ), .B(\mem[9][13] ), .S(n1567), .Z(n1479) );
  MUX2_X1 U1580 ( .A(n1479), .B(n1478), .S(n1559), .Z(n1480) );
  MUX2_X1 U1581 ( .A(n1480), .B(n1477), .S(n1554), .Z(n1481) );
  MUX2_X1 U1582 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n1568), .Z(n1482) );
  MUX2_X1 U1583 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n1568), .Z(n1483) );
  MUX2_X1 U1584 ( .A(n1483), .B(n1482), .S(n1559), .Z(n1484) );
  MUX2_X1 U1585 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n1568), .Z(n1485) );
  MUX2_X1 U1586 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n1568), .Z(n1486) );
  MUX2_X1 U1587 ( .A(n1486), .B(n1485), .S(n1559), .Z(n1487) );
  MUX2_X1 U1588 ( .A(n1487), .B(n1484), .S(n1554), .Z(n1488) );
  MUX2_X1 U1589 ( .A(n1488), .B(n1481), .S(n1551), .Z(n1489) );
  MUX2_X1 U1590 ( .A(n1489), .B(n1474), .S(N14), .Z(N17) );
  MUX2_X1 U1591 ( .A(\mem[30][14] ), .B(\mem[31][14] ), .S(n1568), .Z(n1490)
         );
  MUX2_X1 U1592 ( .A(\mem[28][14] ), .B(\mem[29][14] ), .S(n1568), .Z(n1491)
         );
  MUX2_X1 U1593 ( .A(n1491), .B(n1490), .S(n1559), .Z(n1492) );
  MUX2_X1 U1594 ( .A(\mem[26][14] ), .B(\mem[27][14] ), .S(n1568), .Z(n1493)
         );
  MUX2_X1 U1595 ( .A(\mem[24][14] ), .B(\mem[25][14] ), .S(n1568), .Z(n1494)
         );
  MUX2_X1 U1596 ( .A(n1494), .B(n1493), .S(n1559), .Z(n1495) );
  MUX2_X1 U1597 ( .A(n1495), .B(n1492), .S(n1554), .Z(n1496) );
  MUX2_X1 U1598 ( .A(\mem[22][14] ), .B(\mem[23][14] ), .S(n1568), .Z(n1497)
         );
  MUX2_X1 U1599 ( .A(\mem[20][14] ), .B(\mem[21][14] ), .S(n1568), .Z(n1498)
         );
  MUX2_X1 U1600 ( .A(n1498), .B(n1497), .S(n1559), .Z(n1499) );
  MUX2_X1 U1601 ( .A(\mem[18][14] ), .B(\mem[19][14] ), .S(n1568), .Z(n1500)
         );
  MUX2_X1 U1602 ( .A(\mem[16][14] ), .B(\mem[17][14] ), .S(n1568), .Z(n1501)
         );
  MUX2_X1 U1603 ( .A(n1501), .B(n1500), .S(n1559), .Z(n1502) );
  MUX2_X1 U1604 ( .A(n1502), .B(n1499), .S(n1554), .Z(n1503) );
  MUX2_X1 U1605 ( .A(n1503), .B(n1496), .S(n1551), .Z(n1504) );
  MUX2_X1 U1606 ( .A(\mem[14][14] ), .B(\mem[15][14] ), .S(n1569), .Z(n1505)
         );
  MUX2_X1 U1607 ( .A(\mem[12][14] ), .B(\mem[13][14] ), .S(n1569), .Z(n1506)
         );
  MUX2_X1 U1608 ( .A(n1506), .B(n1505), .S(n1558), .Z(n1507) );
  MUX2_X1 U1609 ( .A(\mem[10][14] ), .B(\mem[11][14] ), .S(n1569), .Z(n1508)
         );
  MUX2_X1 U1610 ( .A(\mem[8][14] ), .B(\mem[9][14] ), .S(n1569), .Z(n1509) );
  MUX2_X1 U1611 ( .A(n1509), .B(n1508), .S(n1556), .Z(n1510) );
  MUX2_X1 U1612 ( .A(n1510), .B(n1507), .S(n1554), .Z(n1511) );
  MUX2_X1 U1613 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n1569), .Z(n1512) );
  MUX2_X1 U1614 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n1569), .Z(n1513) );
  MUX2_X1 U1615 ( .A(n1513), .B(n1512), .S(n1559), .Z(n1514) );
  MUX2_X1 U1616 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n1569), .Z(n1515) );
  MUX2_X1 U1617 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n1569), .Z(n1516) );
  MUX2_X1 U1618 ( .A(n1516), .B(n1515), .S(n1559), .Z(n1517) );
  MUX2_X1 U1619 ( .A(n1517), .B(n1514), .S(n1554), .Z(n1518) );
  MUX2_X1 U1620 ( .A(n1518), .B(n1511), .S(n1551), .Z(n1519) );
  MUX2_X1 U1621 ( .A(n1519), .B(n1504), .S(N14), .Z(N16) );
  MUX2_X1 U1622 ( .A(\mem[30][15] ), .B(\mem[31][15] ), .S(n1569), .Z(n1520)
         );
  MUX2_X1 U1623 ( .A(\mem[28][15] ), .B(\mem[29][15] ), .S(n1569), .Z(n1521)
         );
  MUX2_X1 U1624 ( .A(n1521), .B(n1520), .S(n1560), .Z(n1522) );
  MUX2_X1 U1625 ( .A(\mem[26][15] ), .B(\mem[27][15] ), .S(n1569), .Z(n1523)
         );
  MUX2_X1 U1626 ( .A(\mem[24][15] ), .B(\mem[25][15] ), .S(n1569), .Z(n1524)
         );
  MUX2_X1 U1627 ( .A(n1524), .B(n1523), .S(n1558), .Z(n1525) );
  MUX2_X1 U1628 ( .A(n1525), .B(n1522), .S(n1554), .Z(n1526) );
  MUX2_X1 U1629 ( .A(\mem[22][15] ), .B(\mem[23][15] ), .S(n1570), .Z(n1527)
         );
  MUX2_X1 U1630 ( .A(\mem[20][15] ), .B(\mem[21][15] ), .S(n1570), .Z(n1528)
         );
  MUX2_X1 U1631 ( .A(n1528), .B(n1527), .S(n1556), .Z(n1529) );
  MUX2_X1 U1632 ( .A(\mem[18][15] ), .B(\mem[19][15] ), .S(n1570), .Z(n1530)
         );
  MUX2_X1 U1633 ( .A(\mem[16][15] ), .B(\mem[17][15] ), .S(n1570), .Z(n1531)
         );
  MUX2_X1 U1634 ( .A(n1531), .B(n1530), .S(n1558), .Z(n1532) );
  MUX2_X1 U1635 ( .A(n1532), .B(n1529), .S(n1554), .Z(n1533) );
  MUX2_X1 U1636 ( .A(n1533), .B(n1526), .S(n1551), .Z(n1534) );
  MUX2_X1 U1637 ( .A(\mem[14][15] ), .B(\mem[15][15] ), .S(n1570), .Z(n1535)
         );
  MUX2_X1 U1638 ( .A(\mem[12][15] ), .B(\mem[13][15] ), .S(n1570), .Z(n1536)
         );
  MUX2_X1 U1639 ( .A(n1536), .B(n1535), .S(n1559), .Z(n1537) );
  MUX2_X1 U1640 ( .A(\mem[10][15] ), .B(\mem[11][15] ), .S(n1570), .Z(n1538)
         );
  MUX2_X1 U1641 ( .A(\mem[8][15] ), .B(\mem[9][15] ), .S(n1570), .Z(n1539) );
  MUX2_X1 U1642 ( .A(n1539), .B(n1538), .S(n1558), .Z(n1540) );
  MUX2_X1 U1643 ( .A(n1540), .B(n1537), .S(n1554), .Z(n1541) );
  MUX2_X1 U1644 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n1570), .Z(n1542) );
  MUX2_X1 U1645 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n1570), .Z(n1543) );
  MUX2_X1 U1646 ( .A(n1543), .B(n1542), .S(n1556), .Z(n1544) );
  MUX2_X1 U1647 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n1570), .Z(n1545) );
  MUX2_X1 U1648 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n1570), .Z(n1546) );
  MUX2_X1 U1649 ( .A(n1546), .B(n1545), .S(n1556), .Z(n1547) );
  MUX2_X1 U1650 ( .A(n1547), .B(n1544), .S(n1554), .Z(n1548) );
  MUX2_X1 U1651 ( .A(n1548), .B(n1541), .S(n1551), .Z(n1549) );
  MUX2_X1 U1652 ( .A(n1549), .B(n1534), .S(N14), .Z(N15) );
  CLKBUF_X1 U1653 ( .A(N12), .Z(n1552) );
  CLKBUF_X1 U1654 ( .A(N12), .Z(n1553) );
  CLKBUF_X1 U1655 ( .A(N12), .Z(n1554) );
  CLKBUF_X1 U1656 ( .A(N11), .Z(n1555) );
  INV_X1 U1657 ( .A(N10), .ZN(n1621) );
  INV_X1 U1658 ( .A(N11), .ZN(n1622) );
  INV_X1 U1659 ( .A(N13), .ZN(n1623) );
endmodule


module datapath_K32_logK6_b8_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357;

  FA_X1 U12 ( .A(n12), .B(n55), .CI(n54), .CO(n11), .S(product[4]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n299), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n298), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n297), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n296), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n295), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n79), .B(n69), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n92), .CI(n80), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n94), .B(n88), .CI(n101), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  INV_X1 U157 ( .A(n304), .ZN(n206) );
  INV_X1 U158 ( .A(n306), .ZN(n288) );
  BUF_X1 U159 ( .A(n325), .Z(n291) );
  NAND3_X1 U160 ( .A1(n282), .A2(n283), .A3(n284), .ZN(n49) );
  INV_X1 U161 ( .A(n15), .ZN(n300) );
  XOR2_X1 U162 ( .A(n95), .B(n102), .Z(n207) );
  AND3_X1 U163 ( .A1(n274), .A2(n275), .A3(n276), .ZN(product[15]) );
  XNOR2_X2 U164 ( .A(a[6]), .B(a[5]), .ZN(n334) );
  NAND2_X1 U165 ( .A1(n253), .A2(n34), .ZN(n209) );
  XOR2_X1 U166 ( .A(n305), .B(b[0]), .Z(n314) );
  CLKBUF_X1 U167 ( .A(n351), .Z(n210) );
  XOR2_X1 U168 ( .A(n211), .B(n212), .Z(product[6]) );
  AND3_X1 U169 ( .A1(n241), .A2(n240), .A3(n242), .ZN(n211) );
  XNOR2_X1 U170 ( .A(n46), .B(n49), .ZN(n212) );
  NAND3_X1 U171 ( .A1(n216), .A2(n217), .A3(n218), .ZN(n213) );
  NAND3_X1 U172 ( .A1(n241), .A2(n240), .A3(n242), .ZN(n214) );
  AND2_X1 U173 ( .A1(n104), .A2(n72), .ZN(n215) );
  NAND2_X1 U174 ( .A1(n214), .A2(n46), .ZN(n216) );
  NAND2_X1 U175 ( .A1(n10), .A2(n49), .ZN(n217) );
  NAND2_X1 U176 ( .A1(n46), .A2(n49), .ZN(n218) );
  NAND3_X1 U177 ( .A1(n216), .A2(n217), .A3(n218), .ZN(n9) );
  NAND3_X1 U178 ( .A1(n271), .A2(n272), .A3(n270), .ZN(n219) );
  NAND3_X1 U179 ( .A1(n271), .A2(n272), .A3(n270), .ZN(n220) );
  NAND3_X1 U180 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n221) );
  NAND3_X1 U181 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n222) );
  XNOR2_X1 U182 ( .A(n223), .B(n215), .ZN(product[2]) );
  XNOR2_X1 U183 ( .A(n103), .B(n96), .ZN(n223) );
  XNOR2_X1 U184 ( .A(n224), .B(n226), .ZN(product[3]) );
  XNOR2_X1 U185 ( .A(n207), .B(n71), .ZN(n224) );
  NAND2_X1 U186 ( .A1(n334), .A2(n353), .ZN(n336) );
  NAND3_X1 U187 ( .A1(n229), .A2(n228), .A3(n227), .ZN(n225) );
  NAND3_X1 U188 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n226) );
  NAND2_X1 U189 ( .A1(n103), .A2(n96), .ZN(n227) );
  NAND2_X1 U190 ( .A1(n103), .A2(n215), .ZN(n228) );
  NAND2_X1 U191 ( .A1(n96), .A2(n14), .ZN(n229) );
  NAND3_X1 U192 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n13) );
  NAND2_X1 U193 ( .A1(n207), .A2(n71), .ZN(n230) );
  NAND2_X1 U194 ( .A1(n56), .A2(n225), .ZN(n231) );
  NAND2_X1 U195 ( .A1(n71), .A2(n13), .ZN(n232) );
  NAND3_X1 U196 ( .A1(n230), .A2(n231), .A3(n232), .ZN(n12) );
  XNOR2_X1 U197 ( .A(n233), .B(n255), .ZN(product[13]) );
  AND3_X1 U198 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n233) );
  XOR2_X1 U199 ( .A(n87), .B(n70), .Z(n234) );
  BUF_X2 U200 ( .A(n323), .Z(n235) );
  XOR2_X1 U201 ( .A(a[4]), .B(n305), .Z(n323) );
  NAND3_X1 U202 ( .A1(n257), .A2(n256), .A3(n258), .ZN(n236) );
  XNOR2_X1 U203 ( .A(n237), .B(n273), .ZN(product[14]) );
  AND3_X1 U204 ( .A1(n257), .A2(n256), .A3(n258), .ZN(n237) );
  XNOR2_X1 U205 ( .A(n213), .B(n238), .ZN(product[7]) );
  XNOR2_X1 U206 ( .A(n40), .B(n45), .ZN(n238) );
  XNOR2_X1 U207 ( .A(n11), .B(n239), .ZN(product[5]) );
  XNOR2_X1 U208 ( .A(n50), .B(n53), .ZN(n239) );
  NAND2_X1 U209 ( .A1(n11), .A2(n50), .ZN(n240) );
  NAND2_X1 U210 ( .A1(n11), .A2(n53), .ZN(n241) );
  NAND2_X1 U211 ( .A1(n50), .A2(n53), .ZN(n242) );
  NAND3_X1 U212 ( .A1(n241), .A2(n240), .A3(n242), .ZN(n10) );
  NAND3_X1 U213 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n243) );
  NAND3_X1 U214 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n244) );
  XOR2_X1 U215 ( .A(n27), .B(n24), .Z(n245) );
  XOR2_X1 U216 ( .A(n220), .B(n245), .Z(product[10]) );
  NAND2_X1 U217 ( .A1(n219), .A2(n27), .ZN(n246) );
  NAND2_X1 U218 ( .A1(n6), .A2(n24), .ZN(n247) );
  NAND2_X1 U219 ( .A1(n27), .A2(n24), .ZN(n248) );
  NAND3_X1 U220 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n5) );
  XOR2_X1 U221 ( .A(n18), .B(n19), .Z(n249) );
  XOR2_X1 U222 ( .A(n222), .B(n249), .Z(product[12]) );
  NAND2_X1 U223 ( .A1(n221), .A2(n18), .ZN(n250) );
  NAND2_X1 U224 ( .A1(n4), .A2(n19), .ZN(n251) );
  NAND2_X1 U225 ( .A1(n18), .A2(n19), .ZN(n252) );
  NAND3_X1 U226 ( .A1(n285), .A2(n287), .A3(n286), .ZN(n253) );
  NAND3_X1 U227 ( .A1(n285), .A2(n286), .A3(n287), .ZN(n254) );
  XOR2_X1 U228 ( .A(n17), .B(n300), .Z(n255) );
  NAND2_X1 U229 ( .A1(n243), .A2(n17), .ZN(n256) );
  NAND2_X1 U230 ( .A1(n243), .A2(n300), .ZN(n257) );
  NAND2_X1 U231 ( .A1(n17), .A2(n300), .ZN(n258) );
  NAND3_X1 U232 ( .A1(n257), .A2(n256), .A3(n258), .ZN(n2) );
  XOR2_X1 U233 ( .A(n23), .B(n20), .Z(n259) );
  XOR2_X1 U234 ( .A(n244), .B(n259), .Z(product[11]) );
  NAND2_X1 U235 ( .A1(n244), .A2(n23), .ZN(n260) );
  NAND2_X1 U236 ( .A1(n5), .A2(n20), .ZN(n261) );
  NAND2_X1 U237 ( .A1(n23), .A2(n20), .ZN(n262) );
  NAND3_X1 U238 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n4) );
  NAND3_X1 U239 ( .A1(n209), .A2(n266), .A3(n268), .ZN(n263) );
  NAND3_X1 U240 ( .A1(n266), .A2(n209), .A3(n268), .ZN(n264) );
  XOR2_X1 U241 ( .A(n34), .B(n39), .Z(n265) );
  XOR2_X1 U242 ( .A(n265), .B(n254), .Z(product[8]) );
  NAND2_X1 U243 ( .A1(n34), .A2(n39), .ZN(n266) );
  NAND2_X1 U244 ( .A1(n253), .A2(n34), .ZN(n267) );
  NAND2_X1 U245 ( .A1(n8), .A2(n39), .ZN(n268) );
  NAND3_X1 U246 ( .A1(n268), .A2(n266), .A3(n267), .ZN(n7) );
  XOR2_X1 U247 ( .A(n28), .B(n33), .Z(n269) );
  XOR2_X1 U248 ( .A(n269), .B(n264), .Z(product[9]) );
  NAND2_X1 U249 ( .A1(n28), .A2(n33), .ZN(n270) );
  NAND2_X1 U250 ( .A1(n263), .A2(n28), .ZN(n271) );
  NAND2_X1 U251 ( .A1(n7), .A2(n33), .ZN(n272) );
  NAND3_X1 U252 ( .A1(n271), .A2(n272), .A3(n270), .ZN(n6) );
  XOR2_X1 U253 ( .A(n301), .B(n15), .Z(n273) );
  NAND2_X1 U254 ( .A1(n236), .A2(n301), .ZN(n274) );
  NAND2_X1 U255 ( .A1(n2), .A2(n15), .ZN(n275) );
  NAND2_X1 U256 ( .A1(n301), .A2(n15), .ZN(n276) );
  XOR2_X1 U257 ( .A(a[2]), .B(a[3]), .Z(n351) );
  CLKBUF_X1 U258 ( .A(n309), .Z(n280) );
  INV_X1 U259 ( .A(n289), .ZN(n277) );
  INV_X1 U260 ( .A(n289), .ZN(n290) );
  BUF_X1 U261 ( .A(a[1]), .Z(n279) );
  INV_X1 U262 ( .A(n31), .ZN(n296) );
  INV_X1 U263 ( .A(n332), .ZN(n299) );
  XNOR2_X1 U264 ( .A(n52), .B(n278), .ZN(n50) );
  XNOR2_X1 U265 ( .A(n93), .B(n100), .ZN(n278) );
  INV_X1 U266 ( .A(n21), .ZN(n298) );
  INV_X1 U267 ( .A(n343), .ZN(n301) );
  INV_X1 U268 ( .A(n312), .ZN(n295) );
  INV_X1 U269 ( .A(n321), .ZN(n297) );
  INV_X1 U270 ( .A(a[5]), .ZN(n304) );
  INV_X1 U271 ( .A(a[7]), .ZN(n303) );
  INV_X1 U272 ( .A(b[0]), .ZN(n302) );
  INV_X1 U273 ( .A(a[0]), .ZN(n281) );
  INV_X1 U274 ( .A(a[0]), .ZN(n307) );
  XNOR2_X2 U275 ( .A(a[1]), .B(a[2]), .ZN(n294) );
  NAND2_X1 U276 ( .A1(n234), .A2(n93), .ZN(n282) );
  NAND2_X1 U277 ( .A1(n234), .A2(n100), .ZN(n283) );
  NAND2_X1 U278 ( .A1(n93), .A2(n100), .ZN(n284) );
  NAND2_X1 U279 ( .A1(n9), .A2(n40), .ZN(n285) );
  NAND2_X1 U280 ( .A1(n9), .A2(n45), .ZN(n286) );
  NAND2_X1 U281 ( .A1(n40), .A2(n45), .ZN(n287) );
  NAND3_X1 U282 ( .A1(n286), .A2(n287), .A3(n285), .ZN(n8) );
  NAND2_X1 U283 ( .A1(a[1]), .A2(n307), .ZN(n309) );
  XNOR2_X1 U284 ( .A(a[1]), .B(a[2]), .ZN(n313) );
  INV_X1 U285 ( .A(a[3]), .ZN(n289) );
  NAND2_X1 U286 ( .A1(n323), .A2(n352), .ZN(n325) );
  NAND2_X1 U287 ( .A1(n351), .A2(n313), .ZN(n292) );
  NAND2_X1 U288 ( .A1(n294), .A2(n210), .ZN(n293) );
  NAND2_X1 U289 ( .A1(n351), .A2(n313), .ZN(n315) );
  INV_X1 U290 ( .A(a[3]), .ZN(n305) );
  INV_X1 U291 ( .A(a[1]), .ZN(n306) );
  NOR2_X1 U292 ( .A1(n281), .A2(n302), .ZN(product[0]) );
  OAI22_X1 U293 ( .A1(n308), .A2(n280), .B1(n310), .B2(n281), .ZN(n99) );
  OAI22_X1 U294 ( .A1(n310), .A2(n280), .B1(n311), .B2(n281), .ZN(n98) );
  XNOR2_X1 U295 ( .A(b[6]), .B(n288), .ZN(n310) );
  OAI22_X1 U296 ( .A1(n281), .A2(n311), .B1(n280), .B2(n311), .ZN(n312) );
  XNOR2_X1 U297 ( .A(b[7]), .B(n288), .ZN(n311) );
  NOR2_X1 U298 ( .A1(n294), .A2(n302), .ZN(n96) );
  OAI22_X1 U299 ( .A1(n314), .A2(n315), .B1(n294), .B2(n316), .ZN(n95) );
  OAI22_X1 U300 ( .A1(n316), .A2(n292), .B1(n294), .B2(n317), .ZN(n94) );
  XNOR2_X1 U301 ( .A(b[1]), .B(n290), .ZN(n316) );
  OAI22_X1 U302 ( .A1(n317), .A2(n293), .B1(n294), .B2(n318), .ZN(n93) );
  XNOR2_X1 U303 ( .A(b[2]), .B(n277), .ZN(n317) );
  OAI22_X1 U304 ( .A1(n318), .A2(n292), .B1(n294), .B2(n319), .ZN(n92) );
  XNOR2_X1 U305 ( .A(b[3]), .B(n277), .ZN(n318) );
  OAI22_X1 U306 ( .A1(n319), .A2(n292), .B1(n294), .B2(n320), .ZN(n91) );
  XNOR2_X1 U307 ( .A(b[4]), .B(n277), .ZN(n319) );
  OAI22_X1 U308 ( .A1(n322), .A2(n294), .B1(n292), .B2(n322), .ZN(n321) );
  NOR2_X1 U309 ( .A1(n323), .A2(n302), .ZN(n88) );
  OAI22_X1 U310 ( .A1(n324), .A2(n325), .B1(n235), .B2(n326), .ZN(n87) );
  XNOR2_X1 U311 ( .A(a[5]), .B(b[0]), .ZN(n324) );
  OAI22_X1 U312 ( .A1(n326), .A2(n291), .B1(n235), .B2(n327), .ZN(n86) );
  XNOR2_X1 U313 ( .A(b[1]), .B(a[5]), .ZN(n326) );
  OAI22_X1 U314 ( .A1(n327), .A2(n291), .B1(n235), .B2(n328), .ZN(n85) );
  XNOR2_X1 U315 ( .A(b[2]), .B(a[5]), .ZN(n327) );
  OAI22_X1 U316 ( .A1(n328), .A2(n291), .B1(n235), .B2(n329), .ZN(n84) );
  XNOR2_X1 U317 ( .A(b[3]), .B(a[5]), .ZN(n328) );
  OAI22_X1 U318 ( .A1(n329), .A2(n291), .B1(n235), .B2(n330), .ZN(n83) );
  XNOR2_X1 U319 ( .A(b[4]), .B(n206), .ZN(n329) );
  OAI22_X1 U320 ( .A1(n330), .A2(n291), .B1(n235), .B2(n331), .ZN(n82) );
  XNOR2_X1 U321 ( .A(b[5]), .B(n206), .ZN(n330) );
  OAI22_X1 U322 ( .A1(n333), .A2(n235), .B1(n291), .B2(n333), .ZN(n332) );
  NOR2_X1 U323 ( .A1(n334), .A2(n302), .ZN(n80) );
  OAI22_X1 U324 ( .A1(n335), .A2(n336), .B1(n334), .B2(n337), .ZN(n79) );
  XNOR2_X1 U325 ( .A(a[7]), .B(b[0]), .ZN(n335) );
  OAI22_X1 U326 ( .A1(n338), .A2(n336), .B1(n334), .B2(n339), .ZN(n77) );
  OAI22_X1 U327 ( .A1(n339), .A2(n336), .B1(n334), .B2(n340), .ZN(n76) );
  XNOR2_X1 U328 ( .A(b[3]), .B(a[7]), .ZN(n339) );
  OAI22_X1 U329 ( .A1(n340), .A2(n336), .B1(n334), .B2(n341), .ZN(n75) );
  XNOR2_X1 U330 ( .A(b[4]), .B(a[7]), .ZN(n340) );
  OAI22_X1 U331 ( .A1(n341), .A2(n336), .B1(n334), .B2(n342), .ZN(n74) );
  XNOR2_X1 U332 ( .A(b[5]), .B(a[7]), .ZN(n341) );
  OAI22_X1 U333 ( .A1(n344), .A2(n334), .B1(n336), .B2(n344), .ZN(n343) );
  OAI21_X1 U334 ( .B1(b[0]), .B2(n306), .A(n309), .ZN(n72) );
  OAI21_X1 U335 ( .B1(n305), .B2(n293), .A(n345), .ZN(n71) );
  OR3_X1 U336 ( .A1(n294), .A2(b[0]), .A3(n305), .ZN(n345) );
  OAI21_X1 U337 ( .B1(n304), .B2(n325), .A(n346), .ZN(n70) );
  OR3_X1 U338 ( .A1(n323), .A2(b[0]), .A3(n304), .ZN(n346) );
  OAI21_X1 U339 ( .B1(n303), .B2(n336), .A(n347), .ZN(n69) );
  OR3_X1 U340 ( .A1(n334), .A2(b[0]), .A3(n303), .ZN(n347) );
  XNOR2_X1 U341 ( .A(n348), .B(n349), .ZN(n38) );
  OR2_X1 U342 ( .A1(n348), .A2(n349), .ZN(n37) );
  OAI22_X1 U343 ( .A1(n320), .A2(n293), .B1(n294), .B2(n350), .ZN(n349) );
  XNOR2_X1 U344 ( .A(b[5]), .B(n277), .ZN(n320) );
  OAI22_X1 U345 ( .A1(n337), .A2(n336), .B1(n334), .B2(n338), .ZN(n348) );
  XNOR2_X1 U346 ( .A(b[2]), .B(a[7]), .ZN(n338) );
  XNOR2_X1 U347 ( .A(b[1]), .B(a[7]), .ZN(n337) );
  OAI22_X1 U348 ( .A1(n350), .A2(n293), .B1(n294), .B2(n322), .ZN(n31) );
  XNOR2_X1 U349 ( .A(b[7]), .B(n277), .ZN(n322) );
  XNOR2_X1 U350 ( .A(b[6]), .B(n290), .ZN(n350) );
  OAI22_X1 U351 ( .A1(n331), .A2(n291), .B1(n235), .B2(n333), .ZN(n21) );
  XNOR2_X1 U352 ( .A(b[7]), .B(n206), .ZN(n333) );
  XNOR2_X1 U353 ( .A(n304), .B(a[4]), .ZN(n352) );
  XNOR2_X1 U354 ( .A(b[6]), .B(n206), .ZN(n331) );
  OAI22_X1 U355 ( .A1(n342), .A2(n336), .B1(n334), .B2(n344), .ZN(n15) );
  XNOR2_X1 U356 ( .A(b[7]), .B(a[7]), .ZN(n344) );
  XNOR2_X1 U357 ( .A(n303), .B(a[6]), .ZN(n353) );
  XNOR2_X1 U358 ( .A(b[6]), .B(a[7]), .ZN(n342) );
  OAI22_X1 U359 ( .A1(b[0]), .A2(n309), .B1(n354), .B2(n281), .ZN(n104) );
  OAI22_X1 U360 ( .A1(n354), .A2(n309), .B1(n355), .B2(n307), .ZN(n103) );
  XNOR2_X1 U361 ( .A(a[1]), .B(b[1]), .ZN(n354) );
  OAI22_X1 U362 ( .A1(n355), .A2(n309), .B1(n356), .B2(n281), .ZN(n102) );
  XNOR2_X1 U363 ( .A(n279), .B(b[2]), .ZN(n355) );
  OAI22_X1 U364 ( .A1(n356), .A2(n280), .B1(n357), .B2(n307), .ZN(n101) );
  XNOR2_X1 U365 ( .A(n279), .B(b[3]), .ZN(n356) );
  OAI22_X1 U366 ( .A1(n357), .A2(n280), .B1(n308), .B2(n281), .ZN(n100) );
  XNOR2_X1 U367 ( .A(b[5]), .B(n288), .ZN(n308) );
  XNOR2_X1 U368 ( .A(b[4]), .B(n288), .ZN(n357) );
endmodule


module datapath_K32_logK6_b8_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(n83), .B(B[1]), .CI(A[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(A[7]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(A[11]), .Z(n2) );
  CLKBUF_X1 U3 ( .A(n70), .Z(n3) );
  CLKBUF_X1 U4 ( .A(A[12]), .Z(n4) );
  CLKBUF_X1 U5 ( .A(n77), .Z(n5) );
  NAND3_X1 U6 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n6) );
  NAND3_X1 U7 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n7) );
  NAND3_X1 U8 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n8) );
  CLKBUF_X1 U9 ( .A(n42), .Z(n9) );
  NAND3_X1 U10 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n10) );
  XNOR2_X1 U11 ( .A(A[15]), .B(B[15]), .ZN(n78) );
  CLKBUF_X1 U12 ( .A(n20), .Z(n11) );
  NAND3_X1 U13 ( .A1(n42), .A2(n44), .A3(n43), .ZN(n12) );
  NAND3_X1 U14 ( .A1(n9), .A2(n44), .A3(n43), .ZN(n13) );
  NAND3_X1 U15 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n14) );
  CLKBUF_X1 U16 ( .A(carry[10]), .Z(n15) );
  XOR2_X1 U17 ( .A(carry[2]), .B(B[2]), .Z(n16) );
  XOR2_X1 U18 ( .A(A[2]), .B(n16), .Z(SUM[2]) );
  NAND2_X1 U19 ( .A1(A[2]), .A2(carry[2]), .ZN(n17) );
  NAND2_X1 U20 ( .A1(A[2]), .A2(B[2]), .ZN(n18) );
  NAND2_X1 U21 ( .A1(carry[2]), .A2(B[2]), .ZN(n19) );
  NAND3_X1 U22 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[3]) );
  NAND3_X1 U23 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n20) );
  CLKBUF_X1 U24 ( .A(n14), .Z(n21) );
  NAND3_X1 U25 ( .A1(n27), .A2(n26), .A3(n25), .ZN(n22) );
  NAND3_X1 U26 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n23) );
  XOR2_X1 U27 ( .A(A[3]), .B(B[3]), .Z(n24) );
  XOR2_X1 U28 ( .A(n24), .B(n10), .Z(SUM[3]) );
  NAND2_X1 U29 ( .A1(A[3]), .A2(B[3]), .ZN(n25) );
  NAND2_X1 U30 ( .A1(A[3]), .A2(n10), .ZN(n26) );
  NAND2_X1 U31 ( .A1(B[3]), .A2(carry[3]), .ZN(n27) );
  NAND3_X1 U32 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[4]) );
  XOR2_X1 U33 ( .A(A[4]), .B(B[4]), .Z(n28) );
  XOR2_X1 U34 ( .A(n28), .B(n23), .Z(SUM[4]) );
  NAND2_X1 U35 ( .A1(A[4]), .A2(B[4]), .ZN(n29) );
  NAND2_X1 U36 ( .A1(A[4]), .A2(n22), .ZN(n30) );
  NAND2_X1 U37 ( .A1(B[4]), .A2(carry[4]), .ZN(n31) );
  NAND3_X1 U38 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[5]) );
  XOR2_X1 U39 ( .A(A[5]), .B(B[5]), .Z(n32) );
  XOR2_X1 U40 ( .A(n7), .B(n32), .Z(SUM[5]) );
  NAND2_X1 U41 ( .A1(n6), .A2(A[5]), .ZN(n33) );
  NAND2_X1 U42 ( .A1(carry[5]), .A2(B[5]), .ZN(n34) );
  NAND2_X1 U43 ( .A1(A[5]), .A2(B[5]), .ZN(n35) );
  NAND3_X1 U44 ( .A1(n34), .A2(n33), .A3(n35), .ZN(carry[6]) );
  XOR2_X1 U45 ( .A(n21), .B(B[6]), .Z(n36) );
  XOR2_X1 U46 ( .A(A[6]), .B(n36), .Z(SUM[6]) );
  NAND2_X1 U47 ( .A1(n14), .A2(A[6]), .ZN(n37) );
  NAND2_X1 U48 ( .A1(A[6]), .A2(B[6]), .ZN(n38) );
  NAND2_X1 U49 ( .A1(carry[6]), .A2(B[6]), .ZN(n39) );
  NAND3_X1 U50 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[7]) );
  CLKBUF_X1 U51 ( .A(n50), .Z(n40) );
  XOR2_X1 U52 ( .A(n1), .B(B[7]), .Z(n41) );
  XOR2_X1 U53 ( .A(n11), .B(n41), .Z(SUM[7]) );
  NAND2_X1 U54 ( .A1(n20), .A2(A[7]), .ZN(n42) );
  NAND2_X1 U55 ( .A1(carry[7]), .A2(B[7]), .ZN(n43) );
  NAND2_X1 U56 ( .A1(A[7]), .A2(B[7]), .ZN(n44) );
  NAND3_X1 U57 ( .A1(n42), .A2(n44), .A3(n43), .ZN(carry[8]) );
  NAND3_X1 U58 ( .A1(n75), .A2(n76), .A3(n77), .ZN(n45) );
  NAND3_X1 U59 ( .A1(n49), .A2(n40), .A3(n51), .ZN(n46) );
  NAND2_X1 U60 ( .A1(carry[11]), .A2(B[11]), .ZN(n47) );
  XOR2_X1 U61 ( .A(A[8]), .B(B[8]), .Z(n48) );
  XOR2_X1 U62 ( .A(n13), .B(n48), .Z(SUM[8]) );
  NAND2_X1 U63 ( .A1(n12), .A2(A[8]), .ZN(n49) );
  NAND2_X1 U64 ( .A1(carry[8]), .A2(B[8]), .ZN(n50) );
  NAND2_X1 U65 ( .A1(A[8]), .A2(B[8]), .ZN(n51) );
  NAND3_X1 U66 ( .A1(n49), .A2(n50), .A3(n51), .ZN(carry[9]) );
  NAND3_X1 U67 ( .A1(n56), .A2(n55), .A3(n57), .ZN(n52) );
  CLKBUF_X1 U68 ( .A(n47), .Z(n53) );
  XOR2_X1 U69 ( .A(A[9]), .B(B[9]), .Z(n54) );
  XOR2_X1 U70 ( .A(n46), .B(n54), .Z(SUM[9]) );
  NAND2_X1 U71 ( .A1(n8), .A2(A[9]), .ZN(n55) );
  NAND2_X1 U72 ( .A1(carry[9]), .A2(B[9]), .ZN(n56) );
  NAND2_X1 U73 ( .A1(A[9]), .A2(B[9]), .ZN(n57) );
  NAND3_X1 U74 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[10]) );
  NAND3_X1 U75 ( .A1(n47), .A2(n70), .A3(n72), .ZN(n58) );
  NAND3_X1 U76 ( .A1(n53), .A2(n3), .A3(n72), .ZN(n59) );
  NAND3_X1 U77 ( .A1(n67), .A2(n66), .A3(n68), .ZN(n60) );
  CLKBUF_X1 U78 ( .A(n75), .Z(n61) );
  CLKBUF_X1 U79 ( .A(n76), .Z(n62) );
  CLKBUF_X1 U80 ( .A(carry[11]), .Z(n63) );
  NAND3_X1 U81 ( .A1(n61), .A2(n62), .A3(n5), .ZN(n64) );
  XOR2_X1 U82 ( .A(A[10]), .B(B[10]), .Z(n65) );
  XOR2_X1 U83 ( .A(n15), .B(n65), .Z(SUM[10]) );
  NAND2_X1 U84 ( .A1(n52), .A2(A[10]), .ZN(n66) );
  NAND2_X1 U85 ( .A1(carry[10]), .A2(B[10]), .ZN(n67) );
  NAND2_X1 U86 ( .A1(A[10]), .A2(B[10]), .ZN(n68) );
  NAND3_X1 U87 ( .A1(n67), .A2(n66), .A3(n68), .ZN(carry[11]) );
  XOR2_X1 U88 ( .A(n2), .B(B[11]), .Z(n69) );
  XOR2_X1 U89 ( .A(n63), .B(n69), .Z(SUM[11]) );
  NAND2_X1 U90 ( .A1(n60), .A2(A[11]), .ZN(n70) );
  NAND2_X1 U91 ( .A1(carry[11]), .A2(B[11]), .ZN(n71) );
  NAND2_X1 U92 ( .A1(A[11]), .A2(B[11]), .ZN(n72) );
  NAND3_X1 U93 ( .A1(n70), .A2(n71), .A3(n72), .ZN(carry[12]) );
  NAND3_X1 U94 ( .A1(n75), .A2(n76), .A3(n77), .ZN(n73) );
  XOR2_X1 U95 ( .A(n4), .B(B[12]), .Z(n74) );
  XOR2_X1 U96 ( .A(n59), .B(n74), .Z(SUM[12]) );
  NAND2_X1 U97 ( .A1(n58), .A2(A[12]), .ZN(n75) );
  NAND2_X1 U98 ( .A1(carry[12]), .A2(B[12]), .ZN(n76) );
  NAND2_X1 U99 ( .A1(A[12]), .A2(B[12]), .ZN(n77) );
  XNOR2_X1 U100 ( .A(carry[15]), .B(n78), .ZN(SUM[15]) );
  XOR2_X1 U101 ( .A(A[13]), .B(B[13]), .Z(n79) );
  XOR2_X1 U102 ( .A(n64), .B(n79), .Z(SUM[13]) );
  NAND2_X1 U103 ( .A1(A[13]), .A2(n45), .ZN(n80) );
  NAND2_X1 U104 ( .A1(n73), .A2(B[13]), .ZN(n81) );
  NAND2_X1 U105 ( .A1(A[13]), .A2(B[13]), .ZN(n82) );
  NAND3_X1 U106 ( .A1(n80), .A2(n81), .A3(n82), .ZN(carry[14]) );
  AND2_X1 U107 ( .A1(B[0]), .A2(A[0]), .ZN(n83) );
  XOR2_X1 U108 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module datapath_K32_logK6_b8 ( clk, addr_x, wr_en_x, data_in, addr_a, wr_en_a, 
        clear_acc, addr_y, wr_en_y, data_out );
  input [5:0] addr_x;
  input [7:0] data_in;
  input [11:0] addr_a;
  input [5:0] addr_y;
  output [15:0] data_out;
  input clk, wr_en_x, wr_en_a, clear_acc, wr_en_y;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, \mul[9] , \mul[8] , \mul[7] , \mul[6] , \mul[5] , \mul[4] ,
         \mul[3] , \mul[2] , \mul[1] , \mul[15] , \mul[14] , \mul[13] ,
         \mul[12] , \mul[11] , \mul[10] , \mul[0] , n1;
  wire   [7:0] xout;
  wire   [7:0] aout;
  wire   [15:0] mac;
  wire   [15:0] sum;

  DFF_X1 \mac_reg[14]  ( .D(N17), .CK(clk), .Q(mac[14]) );
  DFF_X1 \mac_reg[13]  ( .D(N16), .CK(clk), .Q(mac[13]) );
  DFF_X1 \mac_reg[12]  ( .D(N15), .CK(clk), .Q(mac[12]) );
  DFF_X1 \mac_reg[11]  ( .D(N14), .CK(clk), .Q(mac[11]) );
  DFF_X1 \mac_reg[10]  ( .D(N13), .CK(clk), .Q(mac[10]) );
  DFF_X1 \mac_reg[9]  ( .D(N12), .CK(clk), .Q(mac[9]) );
  DFF_X1 \mac_reg[8]  ( .D(N11), .CK(clk), .Q(mac[8]) );
  DFF_X1 \mac_reg[7]  ( .D(N10), .CK(clk), .Q(mac[7]) );
  DFF_X1 \mac_reg[6]  ( .D(N9), .CK(clk), .Q(mac[6]) );
  DFF_X1 \mac_reg[5]  ( .D(N8), .CK(clk), .Q(mac[5]) );
  DFF_X1 \mac_reg[4]  ( .D(N7), .CK(clk), .Q(mac[4]) );
  DFF_X1 \mac_reg[3]  ( .D(N6), .CK(clk), .Q(mac[3]) );
  DFF_X1 \mac_reg[2]  ( .D(N5), .CK(clk), .Q(mac[2]) );
  DFF_X1 \mac_reg[1]  ( .D(N4), .CK(clk), .Q(mac[1]) );
  DFF_X1 \mac_reg[0]  ( .D(N3), .CK(clk), .Q(mac[0]) );
  memory_WIDTH8_SIZE32_LOGSIZE6 x ( .clk(clk), .data_in(data_in), .data_out(
        xout), .addr(addr_x), .wr_en(wr_en_x) );
  memory_WIDTH8_SIZE1024_LOGSIZE12 a ( .clk(clk), .data_in(data_in), 
        .data_out(aout), .addr(addr_a), .wr_en(wr_en_a) );
  memory_WIDTH16_SIZE32_LOGSIZE6 y ( .clk(clk), .data_in(mac), .data_out(
        data_out), .addr(addr_y), .wr_en(wr_en_y) );
  datapath_K32_logK6_b8_DW_mult_tc_0 mult_258 ( .a(xout), .b(aout), .product({
        \mul[15] , \mul[14] , \mul[13] , \mul[12] , \mul[11] , \mul[10] , 
        \mul[9] , \mul[8] , \mul[7] , \mul[6] , \mul[5] , \mul[4] , \mul[3] , 
        \mul[2] , \mul[1] , \mul[0] }) );
  datapath_K32_logK6_b8_DW01_add_0 add_259 ( .A({\mul[15] , \mul[14] , 
        \mul[13] , \mul[12] , \mul[11] , \mul[10] , \mul[9] , \mul[8] , 
        \mul[7] , \mul[6] , \mul[5] , \mul[4] , \mul[3] , \mul[2] , \mul[1] , 
        \mul[0] }), .B(mac), .CI(1'b0), .SUM(sum) );
  DFF_X1 \mac_reg[15]  ( .D(N18), .CK(clk), .Q(mac[15]) );
  AND2_X1 U3 ( .A1(sum[0]), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(clear_acc), .ZN(n1) );
  AND2_X1 U5 ( .A1(sum[10]), .A2(n1), .ZN(N13) );
  AND2_X1 U6 ( .A1(sum[11]), .A2(n1), .ZN(N14) );
  AND2_X1 U7 ( .A1(sum[14]), .A2(n1), .ZN(N17) );
  AND2_X1 U8 ( .A1(sum[13]), .A2(n1), .ZN(N16) );
  AND2_X1 U9 ( .A1(sum[12]), .A2(n1), .ZN(N15) );
  AND2_X1 U10 ( .A1(sum[1]), .A2(n1), .ZN(N4) );
  AND2_X1 U11 ( .A1(sum[2]), .A2(n1), .ZN(N5) );
  AND2_X1 U12 ( .A1(sum[3]), .A2(n1), .ZN(N6) );
  AND2_X1 U13 ( .A1(sum[4]), .A2(n1), .ZN(N7) );
  AND2_X1 U14 ( .A1(sum[5]), .A2(n1), .ZN(N8) );
  AND2_X1 U15 ( .A1(sum[6]), .A2(n1), .ZN(N9) );
  AND2_X1 U16 ( .A1(sum[7]), .A2(n1), .ZN(N10) );
  AND2_X1 U17 ( .A1(sum[8]), .A2(n1), .ZN(N11) );
  AND2_X1 U18 ( .A1(sum[9]), .A2(n1), .ZN(N12) );
  AND2_X1 U19 ( .A1(sum[15]), .A2(n1), .ZN(N18) );
endmodule


module mvm_32_1_8_0 ( clk, reset, loadMatrix, loadVector, start, done, data_in, 
        data_out );
  input [7:0] data_in;
  output [15:0] data_out;
  input clk, reset, loadMatrix, loadVector, start;
  output done;
  wire   wr_en_x, wr_en_a, clear_acc, wr_en_y;
  wire   [5:0] addr_x;
  wire   [11:0] addr_a;
  wire   [5:0] addr_y;
  wire   SYNOPSYS_UNCONNECTED__0;

  control_K32_logK6 ctl ( .clk(clk), .start(start), .reset(reset), 
        .loadMatrix(loadMatrix), .loadVector(loadVector), .addr_x({
        SYNOPSYS_UNCONNECTED__0, addr_x[4:0]}), .wr_en_x(wr_en_x), .addr_a(
        addr_a), .wr_en_a(wr_en_a), .clear_acc(clear_acc), .addr_y(addr_y), 
        .wr_en_y(wr_en_y), .done(done) );
  datapath_K32_logK6_b8 dtpth ( .clk(clk), .addr_x({1'b0, addr_x[4:0]}), 
        .wr_en_x(wr_en_x), .data_in(data_in), .addr_a(addr_a), .wr_en_a(
        wr_en_a), .clear_acc(clear_acc), .addr_y(addr_y), .wr_en_y(wr_en_y), 
        .data_out(data_out) );
endmodule

